magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal1 >>
rect 1500 1959 1530 2011
rect 1702 1959 1732 2011
rect 3996 1959 4026 2011
rect 4198 1959 4228 2011
rect 6492 1959 6522 2011
rect 6694 1959 6724 2011
rect 8988 1959 9018 2011
rect 9190 1959 9220 2011
rect 11484 1959 11514 2011
rect 11686 1959 11716 2011
rect 13980 1959 14010 2011
rect 14182 1959 14212 2011
rect 16476 1959 16506 2011
rect 16678 1959 16708 2011
rect 18972 1959 19002 2011
rect 19174 1959 19204 2011
rect 21468 1959 21498 2011
rect 21670 1959 21700 2011
rect 23964 1959 23994 2011
rect 24166 1959 24196 2011
rect 26460 1959 26490 2011
rect 26662 1959 26692 2011
rect 28956 1959 28986 2011
rect 29158 1959 29188 2011
rect 31452 1959 31482 2011
rect 31654 1959 31684 2011
rect 33948 1959 33978 2011
rect 34150 1959 34180 2011
rect 36444 1959 36474 2011
rect 36646 1959 36676 2011
rect 38940 1959 38970 2011
rect 39142 1959 39172 2011
rect 41436 1959 41466 2011
rect 41638 1959 41668 2011
rect 43932 1959 43962 2011
rect 44134 1959 44164 2011
rect 46428 1959 46458 2011
rect 46630 1959 46660 2011
rect 48924 1959 48954 2011
rect 49126 1959 49156 2011
rect 51420 1959 51450 2011
rect 51622 1959 51652 2011
rect 53916 1959 53946 2011
rect 54118 1959 54148 2011
rect 56412 1959 56442 2011
rect 56614 1959 56644 2011
rect 58908 1959 58938 2011
rect 59110 1959 59140 2011
rect 61404 1959 61434 2011
rect 61606 1959 61636 2011
rect 63900 1959 63930 2011
rect 64102 1959 64132 2011
rect 66396 1959 66426 2011
rect 66598 1959 66628 2011
rect 68892 1959 68922 2011
rect 69094 1959 69124 2011
rect 71388 1959 71418 2011
rect 71590 1959 71620 2011
rect 73884 1959 73914 2011
rect 74086 1959 74116 2011
rect 76380 1959 76410 2011
rect 76582 1959 76612 2011
rect 78876 1959 78906 2011
rect 79078 1959 79108 2011
rect 1615 1604 1667 1610
rect 1615 1546 1667 1552
rect 4111 1604 4163 1610
rect 4111 1546 4163 1552
rect 6607 1604 6659 1610
rect 6607 1546 6659 1552
rect 9103 1604 9155 1610
rect 9103 1546 9155 1552
rect 11599 1604 11651 1610
rect 11599 1546 11651 1552
rect 14095 1604 14147 1610
rect 14095 1546 14147 1552
rect 16591 1604 16643 1610
rect 16591 1546 16643 1552
rect 19087 1604 19139 1610
rect 19087 1546 19139 1552
rect 21583 1604 21635 1610
rect 21583 1546 21635 1552
rect 24079 1604 24131 1610
rect 24079 1546 24131 1552
rect 26575 1604 26627 1610
rect 26575 1546 26627 1552
rect 29071 1604 29123 1610
rect 29071 1546 29123 1552
rect 31567 1604 31619 1610
rect 31567 1546 31619 1552
rect 34063 1604 34115 1610
rect 34063 1546 34115 1552
rect 36559 1604 36611 1610
rect 36559 1546 36611 1552
rect 39055 1604 39107 1610
rect 39055 1546 39107 1552
rect 41551 1604 41603 1610
rect 41551 1546 41603 1552
rect 44047 1604 44099 1610
rect 44047 1546 44099 1552
rect 46543 1604 46595 1610
rect 46543 1546 46595 1552
rect 49039 1604 49091 1610
rect 49039 1546 49091 1552
rect 51535 1604 51587 1610
rect 51535 1546 51587 1552
rect 54031 1604 54083 1610
rect 54031 1546 54083 1552
rect 56527 1604 56579 1610
rect 56527 1546 56579 1552
rect 59023 1604 59075 1610
rect 59023 1546 59075 1552
rect 61519 1604 61571 1610
rect 61519 1546 61571 1552
rect 64015 1604 64067 1610
rect 64015 1546 64067 1552
rect 66511 1604 66563 1610
rect 66511 1546 66563 1552
rect 69007 1604 69059 1610
rect 69007 1546 69059 1552
rect 71503 1604 71555 1610
rect 71503 1546 71555 1552
rect 73999 1604 74051 1610
rect 73999 1546 74051 1552
rect 76495 1604 76547 1610
rect 76495 1546 76547 1552
rect 78991 1604 79043 1610
rect 78991 1546 79043 1552
rect 1604 1167 1656 1173
rect 1604 1109 1656 1115
rect 4100 1167 4152 1173
rect 4100 1109 4152 1115
rect 6596 1167 6648 1173
rect 6596 1109 6648 1115
rect 9092 1167 9144 1173
rect 9092 1109 9144 1115
rect 11588 1167 11640 1173
rect 11588 1109 11640 1115
rect 14084 1167 14136 1173
rect 14084 1109 14136 1115
rect 16580 1167 16632 1173
rect 16580 1109 16632 1115
rect 19076 1167 19128 1173
rect 19076 1109 19128 1115
rect 21572 1167 21624 1173
rect 21572 1109 21624 1115
rect 24068 1167 24120 1173
rect 24068 1109 24120 1115
rect 26564 1167 26616 1173
rect 26564 1109 26616 1115
rect 29060 1167 29112 1173
rect 29060 1109 29112 1115
rect 31556 1167 31608 1173
rect 31556 1109 31608 1115
rect 34052 1167 34104 1173
rect 34052 1109 34104 1115
rect 36548 1167 36600 1173
rect 36548 1109 36600 1115
rect 39044 1167 39096 1173
rect 39044 1109 39096 1115
rect 41540 1167 41592 1173
rect 41540 1109 41592 1115
rect 44036 1167 44088 1173
rect 44036 1109 44088 1115
rect 46532 1167 46584 1173
rect 46532 1109 46584 1115
rect 49028 1167 49080 1173
rect 49028 1109 49080 1115
rect 51524 1167 51576 1173
rect 51524 1109 51576 1115
rect 54020 1167 54072 1173
rect 54020 1109 54072 1115
rect 56516 1167 56568 1173
rect 56516 1109 56568 1115
rect 59012 1167 59064 1173
rect 59012 1109 59064 1115
rect 61508 1167 61560 1173
rect 61508 1109 61560 1115
rect 64004 1167 64056 1173
rect 64004 1109 64056 1115
rect 66500 1167 66552 1173
rect 66500 1109 66552 1115
rect 68996 1167 69048 1173
rect 68996 1109 69048 1115
rect 71492 1167 71544 1173
rect 71492 1109 71544 1115
rect 73988 1167 74040 1173
rect 73988 1109 74040 1115
rect 76484 1167 76536 1173
rect 76484 1109 76536 1115
rect 78980 1167 79032 1173
rect 78980 1109 79032 1115
rect 1725 836 1777 842
rect 1725 778 1777 784
rect 4221 836 4273 842
rect 4221 778 4273 784
rect 6717 836 6769 842
rect 6717 778 6769 784
rect 9213 836 9265 842
rect 9213 778 9265 784
rect 11709 836 11761 842
rect 11709 778 11761 784
rect 14205 836 14257 842
rect 14205 778 14257 784
rect 16701 836 16753 842
rect 16701 778 16753 784
rect 19197 836 19249 842
rect 19197 778 19249 784
rect 21693 836 21745 842
rect 21693 778 21745 784
rect 24189 836 24241 842
rect 24189 778 24241 784
rect 26685 836 26737 842
rect 26685 778 26737 784
rect 29181 836 29233 842
rect 29181 778 29233 784
rect 31677 836 31729 842
rect 31677 778 31729 784
rect 34173 836 34225 842
rect 34173 778 34225 784
rect 36669 836 36721 842
rect 36669 778 36721 784
rect 39165 836 39217 842
rect 39165 778 39217 784
rect 41661 836 41713 842
rect 41661 778 41713 784
rect 44157 836 44209 842
rect 44157 778 44209 784
rect 46653 836 46705 842
rect 46653 778 46705 784
rect 49149 836 49201 842
rect 49149 778 49201 784
rect 51645 836 51697 842
rect 51645 778 51697 784
rect 54141 836 54193 842
rect 54141 778 54193 784
rect 56637 836 56689 842
rect 56637 778 56689 784
rect 59133 836 59185 842
rect 59133 778 59185 784
rect 61629 836 61681 842
rect 61629 778 61681 784
rect 64125 836 64177 842
rect 64125 778 64177 784
rect 66621 836 66673 842
rect 66621 778 66673 784
rect 69117 836 69169 842
rect 69117 778 69169 784
rect 71613 836 71665 842
rect 71613 778 71665 784
rect 74109 836 74161 842
rect 74109 778 74161 784
rect 76605 836 76657 842
rect 76605 778 76657 784
rect 79101 836 79153 842
rect 79101 778 79153 784
rect 1610 633 1662 639
rect 1610 575 1662 581
rect 4106 633 4158 639
rect 4106 575 4158 581
rect 6602 633 6654 639
rect 6602 575 6654 581
rect 9098 633 9150 639
rect 9098 575 9150 581
rect 11594 633 11646 639
rect 11594 575 11646 581
rect 14090 633 14142 639
rect 14090 575 14142 581
rect 16586 633 16638 639
rect 16586 575 16638 581
rect 19082 633 19134 639
rect 19082 575 19134 581
rect 21578 633 21630 639
rect 21578 575 21630 581
rect 24074 633 24126 639
rect 24074 575 24126 581
rect 26570 633 26622 639
rect 26570 575 26622 581
rect 29066 633 29118 639
rect 29066 575 29118 581
rect 31562 633 31614 639
rect 31562 575 31614 581
rect 34058 633 34110 639
rect 34058 575 34110 581
rect 36554 633 36606 639
rect 36554 575 36606 581
rect 39050 633 39102 639
rect 39050 575 39102 581
rect 41546 633 41598 639
rect 41546 575 41598 581
rect 44042 633 44094 639
rect 44042 575 44094 581
rect 46538 633 46590 639
rect 46538 575 46590 581
rect 49034 633 49086 639
rect 49034 575 49086 581
rect 51530 633 51582 639
rect 51530 575 51582 581
rect 54026 633 54078 639
rect 54026 575 54078 581
rect 56522 633 56574 639
rect 56522 575 56574 581
rect 59018 633 59070 639
rect 59018 575 59070 581
rect 61514 633 61566 639
rect 61514 575 61566 581
rect 64010 633 64062 639
rect 64010 575 64062 581
rect 66506 633 66558 639
rect 66506 575 66558 581
rect 69002 633 69054 639
rect 69002 575 69054 581
rect 71498 633 71550 639
rect 71498 575 71550 581
rect 73994 633 74046 639
rect 73994 575 74046 581
rect 76490 633 76542 639
rect 76490 575 76542 581
rect 78986 633 79038 639
rect 78986 575 79038 581
rect 1624 217 1676 223
rect 1624 159 1676 165
rect 4120 217 4172 223
rect 4120 159 4172 165
rect 6616 217 6668 223
rect 6616 159 6668 165
rect 9112 217 9164 223
rect 9112 159 9164 165
rect 11608 217 11660 223
rect 11608 159 11660 165
rect 14104 217 14156 223
rect 14104 159 14156 165
rect 16600 217 16652 223
rect 16600 159 16652 165
rect 19096 217 19148 223
rect 19096 159 19148 165
rect 21592 217 21644 223
rect 21592 159 21644 165
rect 24088 217 24140 223
rect 24088 159 24140 165
rect 26584 217 26636 223
rect 26584 159 26636 165
rect 29080 217 29132 223
rect 29080 159 29132 165
rect 31576 217 31628 223
rect 31576 159 31628 165
rect 34072 217 34124 223
rect 34072 159 34124 165
rect 36568 217 36620 223
rect 36568 159 36620 165
rect 39064 217 39116 223
rect 39064 159 39116 165
rect 41560 217 41612 223
rect 41560 159 41612 165
rect 44056 217 44108 223
rect 44056 159 44108 165
rect 46552 217 46604 223
rect 46552 159 46604 165
rect 49048 217 49100 223
rect 49048 159 49100 165
rect 51544 217 51596 223
rect 51544 159 51596 165
rect 54040 217 54092 223
rect 54040 159 54092 165
rect 56536 217 56588 223
rect 56536 159 56588 165
rect 59032 217 59084 223
rect 59032 159 59084 165
rect 61528 217 61580 223
rect 61528 159 61580 165
rect 64024 217 64076 223
rect 64024 159 64076 165
rect 66520 217 66572 223
rect 66520 159 66572 165
rect 69016 217 69068 223
rect 69016 159 69068 165
rect 71512 217 71564 223
rect 71512 159 71564 165
rect 74008 217 74060 223
rect 74008 159 74060 165
rect 76504 217 76556 223
rect 76504 159 76556 165
rect 79000 217 79052 223
rect 79000 159 79052 165
rect 1473 94 20817 128
rect 21441 94 40785 128
rect 41409 94 60753 128
rect 61377 94 80721 128
rect 1629 4 1689 60
rect 4125 4 4185 60
rect 6621 4 6681 60
rect 9117 4 9177 60
rect 11613 4 11673 60
rect 14109 4 14169 60
rect 16605 4 16665 60
rect 19101 4 19161 60
rect 21597 4 21657 60
rect 24093 4 24153 60
rect 26589 4 26649 60
rect 29085 4 29145 60
rect 31581 4 31641 60
rect 34077 4 34137 60
rect 36573 4 36633 60
rect 39069 4 39129 60
rect 41565 4 41625 60
rect 44061 4 44121 60
rect 46557 4 46617 60
rect 49053 4 49113 60
rect 51549 4 51609 60
rect 54045 4 54105 60
rect 56541 4 56601 60
rect 59037 4 59097 60
rect 61533 4 61593 60
rect 64029 4 64089 60
rect 66525 4 66585 60
rect 69021 4 69081 60
rect 71517 4 71577 60
rect 74013 4 74073 60
rect 76509 4 76569 60
rect 79005 4 79065 60
<< via1 >>
rect 1615 1552 1667 1604
rect 4111 1552 4163 1604
rect 6607 1552 6659 1604
rect 9103 1552 9155 1604
rect 11599 1552 11651 1604
rect 14095 1552 14147 1604
rect 16591 1552 16643 1604
rect 19087 1552 19139 1604
rect 21583 1552 21635 1604
rect 24079 1552 24131 1604
rect 26575 1552 26627 1604
rect 29071 1552 29123 1604
rect 31567 1552 31619 1604
rect 34063 1552 34115 1604
rect 36559 1552 36611 1604
rect 39055 1552 39107 1604
rect 41551 1552 41603 1604
rect 44047 1552 44099 1604
rect 46543 1552 46595 1604
rect 49039 1552 49091 1604
rect 51535 1552 51587 1604
rect 54031 1552 54083 1604
rect 56527 1552 56579 1604
rect 59023 1552 59075 1604
rect 61519 1552 61571 1604
rect 64015 1552 64067 1604
rect 66511 1552 66563 1604
rect 69007 1552 69059 1604
rect 71503 1552 71555 1604
rect 73999 1552 74051 1604
rect 76495 1552 76547 1604
rect 78991 1552 79043 1604
rect 1604 1115 1656 1167
rect 4100 1115 4152 1167
rect 6596 1115 6648 1167
rect 9092 1115 9144 1167
rect 11588 1115 11640 1167
rect 14084 1115 14136 1167
rect 16580 1115 16632 1167
rect 19076 1115 19128 1167
rect 21572 1115 21624 1167
rect 24068 1115 24120 1167
rect 26564 1115 26616 1167
rect 29060 1115 29112 1167
rect 31556 1115 31608 1167
rect 34052 1115 34104 1167
rect 36548 1115 36600 1167
rect 39044 1115 39096 1167
rect 41540 1115 41592 1167
rect 44036 1115 44088 1167
rect 46532 1115 46584 1167
rect 49028 1115 49080 1167
rect 51524 1115 51576 1167
rect 54020 1115 54072 1167
rect 56516 1115 56568 1167
rect 59012 1115 59064 1167
rect 61508 1115 61560 1167
rect 64004 1115 64056 1167
rect 66500 1115 66552 1167
rect 68996 1115 69048 1167
rect 71492 1115 71544 1167
rect 73988 1115 74040 1167
rect 76484 1115 76536 1167
rect 78980 1115 79032 1167
rect 1725 784 1777 836
rect 4221 784 4273 836
rect 6717 784 6769 836
rect 9213 784 9265 836
rect 11709 784 11761 836
rect 14205 784 14257 836
rect 16701 784 16753 836
rect 19197 784 19249 836
rect 21693 784 21745 836
rect 24189 784 24241 836
rect 26685 784 26737 836
rect 29181 784 29233 836
rect 31677 784 31729 836
rect 34173 784 34225 836
rect 36669 784 36721 836
rect 39165 784 39217 836
rect 41661 784 41713 836
rect 44157 784 44209 836
rect 46653 784 46705 836
rect 49149 784 49201 836
rect 51645 784 51697 836
rect 54141 784 54193 836
rect 56637 784 56689 836
rect 59133 784 59185 836
rect 61629 784 61681 836
rect 64125 784 64177 836
rect 66621 784 66673 836
rect 69117 784 69169 836
rect 71613 784 71665 836
rect 74109 784 74161 836
rect 76605 784 76657 836
rect 79101 784 79153 836
rect 1610 581 1662 633
rect 4106 581 4158 633
rect 6602 581 6654 633
rect 9098 581 9150 633
rect 11594 581 11646 633
rect 14090 581 14142 633
rect 16586 581 16638 633
rect 19082 581 19134 633
rect 21578 581 21630 633
rect 24074 581 24126 633
rect 26570 581 26622 633
rect 29066 581 29118 633
rect 31562 581 31614 633
rect 34058 581 34110 633
rect 36554 581 36606 633
rect 39050 581 39102 633
rect 41546 581 41598 633
rect 44042 581 44094 633
rect 46538 581 46590 633
rect 49034 581 49086 633
rect 51530 581 51582 633
rect 54026 581 54078 633
rect 56522 581 56574 633
rect 59018 581 59070 633
rect 61514 581 61566 633
rect 64010 581 64062 633
rect 66506 581 66558 633
rect 69002 581 69054 633
rect 71498 581 71550 633
rect 73994 581 74046 633
rect 76490 581 76542 633
rect 78986 581 79038 633
rect 1624 165 1676 217
rect 4120 165 4172 217
rect 6616 165 6668 217
rect 9112 165 9164 217
rect 11608 165 11660 217
rect 14104 165 14156 217
rect 16600 165 16652 217
rect 19096 165 19148 217
rect 21592 165 21644 217
rect 24088 165 24140 217
rect 26584 165 26636 217
rect 29080 165 29132 217
rect 31576 165 31628 217
rect 34072 165 34124 217
rect 36568 165 36620 217
rect 39064 165 39116 217
rect 41560 165 41612 217
rect 44056 165 44108 217
rect 46552 165 46604 217
rect 49048 165 49100 217
rect 51544 165 51596 217
rect 54040 165 54092 217
rect 56536 165 56588 217
rect 59032 165 59084 217
rect 61528 165 61580 217
rect 64024 165 64076 217
rect 66520 165 66572 217
rect 69016 165 69068 217
rect 71512 165 71564 217
rect 74008 165 74060 217
rect 76504 165 76556 217
rect 79000 165 79052 217
<< metal2 >>
rect 1613 1606 1669 1615
rect 1613 1541 1669 1550
rect 4109 1606 4165 1615
rect 4109 1541 4165 1550
rect 6605 1606 6661 1615
rect 6605 1541 6661 1550
rect 9101 1606 9157 1615
rect 9101 1541 9157 1550
rect 11597 1606 11653 1615
rect 11597 1541 11653 1550
rect 14093 1606 14149 1615
rect 14093 1541 14149 1550
rect 16589 1606 16645 1615
rect 16589 1541 16645 1550
rect 19085 1606 19141 1615
rect 19085 1541 19141 1550
rect 21581 1606 21637 1615
rect 21581 1541 21637 1550
rect 24077 1606 24133 1615
rect 24077 1541 24133 1550
rect 26573 1606 26629 1615
rect 26573 1541 26629 1550
rect 29069 1606 29125 1615
rect 29069 1541 29125 1550
rect 31565 1606 31621 1615
rect 31565 1541 31621 1550
rect 34061 1606 34117 1615
rect 34061 1541 34117 1550
rect 36557 1606 36613 1615
rect 36557 1541 36613 1550
rect 39053 1606 39109 1615
rect 39053 1541 39109 1550
rect 41549 1606 41605 1615
rect 41549 1541 41605 1550
rect 44045 1606 44101 1615
rect 44045 1541 44101 1550
rect 46541 1606 46597 1615
rect 46541 1541 46597 1550
rect 49037 1606 49093 1615
rect 49037 1541 49093 1550
rect 51533 1606 51589 1615
rect 51533 1541 51589 1550
rect 54029 1606 54085 1615
rect 54029 1541 54085 1550
rect 56525 1606 56581 1615
rect 56525 1541 56581 1550
rect 59021 1606 59077 1615
rect 59021 1541 59077 1550
rect 61517 1606 61573 1615
rect 61517 1541 61573 1550
rect 64013 1606 64069 1615
rect 64013 1541 64069 1550
rect 66509 1606 66565 1615
rect 66509 1541 66565 1550
rect 69005 1606 69061 1615
rect 69005 1541 69061 1550
rect 71501 1606 71557 1615
rect 71501 1541 71557 1550
rect 73997 1606 74053 1615
rect 73997 1541 74053 1550
rect 76493 1606 76549 1615
rect 76493 1541 76549 1550
rect 78989 1606 79045 1615
rect 78989 1541 79045 1550
rect 1602 1169 1658 1178
rect 1602 1104 1658 1113
rect 4098 1169 4154 1178
rect 4098 1104 4154 1113
rect 6594 1169 6650 1178
rect 6594 1104 6650 1113
rect 9090 1169 9146 1178
rect 9090 1104 9146 1113
rect 11586 1169 11642 1178
rect 11586 1104 11642 1113
rect 14082 1169 14138 1178
rect 14082 1104 14138 1113
rect 16578 1169 16634 1178
rect 16578 1104 16634 1113
rect 19074 1169 19130 1178
rect 19074 1104 19130 1113
rect 21570 1169 21626 1178
rect 21570 1104 21626 1113
rect 24066 1169 24122 1178
rect 24066 1104 24122 1113
rect 26562 1169 26618 1178
rect 26562 1104 26618 1113
rect 29058 1169 29114 1178
rect 29058 1104 29114 1113
rect 31554 1169 31610 1178
rect 31554 1104 31610 1113
rect 34050 1169 34106 1178
rect 34050 1104 34106 1113
rect 36546 1169 36602 1178
rect 36546 1104 36602 1113
rect 39042 1169 39098 1178
rect 39042 1104 39098 1113
rect 41538 1169 41594 1178
rect 41538 1104 41594 1113
rect 44034 1169 44090 1178
rect 44034 1104 44090 1113
rect 46530 1169 46586 1178
rect 46530 1104 46586 1113
rect 49026 1169 49082 1178
rect 49026 1104 49082 1113
rect 51522 1169 51578 1178
rect 51522 1104 51578 1113
rect 54018 1169 54074 1178
rect 54018 1104 54074 1113
rect 56514 1169 56570 1178
rect 56514 1104 56570 1113
rect 59010 1169 59066 1178
rect 59010 1104 59066 1113
rect 61506 1169 61562 1178
rect 61506 1104 61562 1113
rect 64002 1169 64058 1178
rect 64002 1104 64058 1113
rect 66498 1169 66554 1178
rect 66498 1104 66554 1113
rect 68994 1169 69050 1178
rect 68994 1104 69050 1113
rect 71490 1169 71546 1178
rect 71490 1104 71546 1113
rect 73986 1169 74042 1178
rect 73986 1104 74042 1113
rect 76482 1169 76538 1178
rect 76482 1104 76538 1113
rect 78978 1169 79034 1178
rect 78978 1104 79034 1113
rect 1723 837 1779 846
rect 1723 772 1779 781
rect 4219 837 4275 846
rect 4219 772 4275 781
rect 6715 837 6771 846
rect 6715 772 6771 781
rect 9211 837 9267 846
rect 9211 772 9267 781
rect 11707 837 11763 846
rect 11707 772 11763 781
rect 14203 837 14259 846
rect 14203 772 14259 781
rect 16699 837 16755 846
rect 16699 772 16755 781
rect 19195 837 19251 846
rect 19195 772 19251 781
rect 21691 837 21747 846
rect 21691 772 21747 781
rect 24187 837 24243 846
rect 24187 772 24243 781
rect 26683 837 26739 846
rect 26683 772 26739 781
rect 29179 837 29235 846
rect 29179 772 29235 781
rect 31675 837 31731 846
rect 31675 772 31731 781
rect 34171 837 34227 846
rect 34171 772 34227 781
rect 36667 837 36723 846
rect 36667 772 36723 781
rect 39163 837 39219 846
rect 39163 772 39219 781
rect 41659 837 41715 846
rect 41659 772 41715 781
rect 44155 837 44211 846
rect 44155 772 44211 781
rect 46651 837 46707 846
rect 46651 772 46707 781
rect 49147 837 49203 846
rect 49147 772 49203 781
rect 51643 837 51699 846
rect 51643 772 51699 781
rect 54139 837 54195 846
rect 54139 772 54195 781
rect 56635 837 56691 846
rect 56635 772 56691 781
rect 59131 837 59187 846
rect 59131 772 59187 781
rect 61627 837 61683 846
rect 61627 772 61683 781
rect 64123 837 64179 846
rect 64123 772 64179 781
rect 66619 837 66675 846
rect 66619 772 66675 781
rect 69115 837 69171 846
rect 69115 772 69171 781
rect 71611 837 71667 846
rect 71611 772 71667 781
rect 74107 837 74163 846
rect 74107 772 74163 781
rect 76603 837 76659 846
rect 76603 772 76659 781
rect 79099 837 79155 846
rect 79099 772 79155 781
rect 1608 635 1664 644
rect 1608 570 1664 579
rect 4104 635 4160 644
rect 4104 570 4160 579
rect 6600 635 6656 644
rect 6600 570 6656 579
rect 9096 635 9152 644
rect 9096 570 9152 579
rect 11592 635 11648 644
rect 11592 570 11648 579
rect 14088 635 14144 644
rect 14088 570 14144 579
rect 16584 635 16640 644
rect 16584 570 16640 579
rect 19080 635 19136 644
rect 19080 570 19136 579
rect 21576 635 21632 644
rect 21576 570 21632 579
rect 24072 635 24128 644
rect 24072 570 24128 579
rect 26568 635 26624 644
rect 26568 570 26624 579
rect 29064 635 29120 644
rect 29064 570 29120 579
rect 31560 635 31616 644
rect 31560 570 31616 579
rect 34056 635 34112 644
rect 34056 570 34112 579
rect 36552 635 36608 644
rect 36552 570 36608 579
rect 39048 635 39104 644
rect 39048 570 39104 579
rect 41544 635 41600 644
rect 41544 570 41600 579
rect 44040 635 44096 644
rect 44040 570 44096 579
rect 46536 635 46592 644
rect 46536 570 46592 579
rect 49032 635 49088 644
rect 49032 570 49088 579
rect 51528 635 51584 644
rect 51528 570 51584 579
rect 54024 635 54080 644
rect 54024 570 54080 579
rect 56520 635 56576 644
rect 56520 570 56576 579
rect 59016 635 59072 644
rect 59016 570 59072 579
rect 61512 635 61568 644
rect 61512 570 61568 579
rect 64008 635 64064 644
rect 64008 570 64064 579
rect 66504 635 66560 644
rect 66504 570 66560 579
rect 69000 635 69056 644
rect 69000 570 69056 579
rect 71496 635 71552 644
rect 71496 570 71552 579
rect 73992 635 74048 644
rect 73992 570 74048 579
rect 76488 635 76544 644
rect 76488 570 76544 579
rect 78984 635 79040 644
rect 78984 570 79040 579
rect 1622 219 1678 228
rect 1622 154 1678 163
rect 4118 219 4174 228
rect 4118 154 4174 163
rect 6614 219 6670 228
rect 6614 154 6670 163
rect 9110 219 9166 228
rect 9110 154 9166 163
rect 11606 219 11662 228
rect 11606 154 11662 163
rect 14102 219 14158 228
rect 14102 154 14158 163
rect 16598 219 16654 228
rect 16598 154 16654 163
rect 19094 219 19150 228
rect 19094 154 19150 163
rect 21590 219 21646 228
rect 21590 154 21646 163
rect 24086 219 24142 228
rect 24086 154 24142 163
rect 26582 219 26638 228
rect 26582 154 26638 163
rect 29078 219 29134 228
rect 29078 154 29134 163
rect 31574 219 31630 228
rect 31574 154 31630 163
rect 34070 219 34126 228
rect 34070 154 34126 163
rect 36566 219 36622 228
rect 36566 154 36622 163
rect 39062 219 39118 228
rect 39062 154 39118 163
rect 41558 219 41614 228
rect 41558 154 41614 163
rect 44054 219 44110 228
rect 44054 154 44110 163
rect 46550 219 46606 228
rect 46550 154 46606 163
rect 49046 219 49102 228
rect 49046 154 49102 163
rect 51542 219 51598 228
rect 51542 154 51598 163
rect 54038 219 54094 228
rect 54038 154 54094 163
rect 56534 219 56590 228
rect 56534 154 56590 163
rect 59030 219 59086 228
rect 59030 154 59086 163
rect 61526 219 61582 228
rect 61526 154 61582 163
rect 64022 219 64078 228
rect 64022 154 64078 163
rect 66518 219 66574 228
rect 66518 154 66574 163
rect 69014 219 69070 228
rect 69014 154 69070 163
rect 71510 219 71566 228
rect 71510 154 71566 163
rect 74006 219 74062 228
rect 74006 154 74062 163
rect 76502 219 76558 228
rect 76502 154 76558 163
rect 78998 219 79054 228
rect 78998 154 79054 163
<< via2 >>
rect 1613 1604 1669 1606
rect 1613 1552 1615 1604
rect 1615 1552 1667 1604
rect 1667 1552 1669 1604
rect 1613 1550 1669 1552
rect 4109 1604 4165 1606
rect 4109 1552 4111 1604
rect 4111 1552 4163 1604
rect 4163 1552 4165 1604
rect 4109 1550 4165 1552
rect 6605 1604 6661 1606
rect 6605 1552 6607 1604
rect 6607 1552 6659 1604
rect 6659 1552 6661 1604
rect 6605 1550 6661 1552
rect 9101 1604 9157 1606
rect 9101 1552 9103 1604
rect 9103 1552 9155 1604
rect 9155 1552 9157 1604
rect 9101 1550 9157 1552
rect 11597 1604 11653 1606
rect 11597 1552 11599 1604
rect 11599 1552 11651 1604
rect 11651 1552 11653 1604
rect 11597 1550 11653 1552
rect 14093 1604 14149 1606
rect 14093 1552 14095 1604
rect 14095 1552 14147 1604
rect 14147 1552 14149 1604
rect 14093 1550 14149 1552
rect 16589 1604 16645 1606
rect 16589 1552 16591 1604
rect 16591 1552 16643 1604
rect 16643 1552 16645 1604
rect 16589 1550 16645 1552
rect 19085 1604 19141 1606
rect 19085 1552 19087 1604
rect 19087 1552 19139 1604
rect 19139 1552 19141 1604
rect 19085 1550 19141 1552
rect 21581 1604 21637 1606
rect 21581 1552 21583 1604
rect 21583 1552 21635 1604
rect 21635 1552 21637 1604
rect 21581 1550 21637 1552
rect 24077 1604 24133 1606
rect 24077 1552 24079 1604
rect 24079 1552 24131 1604
rect 24131 1552 24133 1604
rect 24077 1550 24133 1552
rect 26573 1604 26629 1606
rect 26573 1552 26575 1604
rect 26575 1552 26627 1604
rect 26627 1552 26629 1604
rect 26573 1550 26629 1552
rect 29069 1604 29125 1606
rect 29069 1552 29071 1604
rect 29071 1552 29123 1604
rect 29123 1552 29125 1604
rect 29069 1550 29125 1552
rect 31565 1604 31621 1606
rect 31565 1552 31567 1604
rect 31567 1552 31619 1604
rect 31619 1552 31621 1604
rect 31565 1550 31621 1552
rect 34061 1604 34117 1606
rect 34061 1552 34063 1604
rect 34063 1552 34115 1604
rect 34115 1552 34117 1604
rect 34061 1550 34117 1552
rect 36557 1604 36613 1606
rect 36557 1552 36559 1604
rect 36559 1552 36611 1604
rect 36611 1552 36613 1604
rect 36557 1550 36613 1552
rect 39053 1604 39109 1606
rect 39053 1552 39055 1604
rect 39055 1552 39107 1604
rect 39107 1552 39109 1604
rect 39053 1550 39109 1552
rect 41549 1604 41605 1606
rect 41549 1552 41551 1604
rect 41551 1552 41603 1604
rect 41603 1552 41605 1604
rect 41549 1550 41605 1552
rect 44045 1604 44101 1606
rect 44045 1552 44047 1604
rect 44047 1552 44099 1604
rect 44099 1552 44101 1604
rect 44045 1550 44101 1552
rect 46541 1604 46597 1606
rect 46541 1552 46543 1604
rect 46543 1552 46595 1604
rect 46595 1552 46597 1604
rect 46541 1550 46597 1552
rect 49037 1604 49093 1606
rect 49037 1552 49039 1604
rect 49039 1552 49091 1604
rect 49091 1552 49093 1604
rect 49037 1550 49093 1552
rect 51533 1604 51589 1606
rect 51533 1552 51535 1604
rect 51535 1552 51587 1604
rect 51587 1552 51589 1604
rect 51533 1550 51589 1552
rect 54029 1604 54085 1606
rect 54029 1552 54031 1604
rect 54031 1552 54083 1604
rect 54083 1552 54085 1604
rect 54029 1550 54085 1552
rect 56525 1604 56581 1606
rect 56525 1552 56527 1604
rect 56527 1552 56579 1604
rect 56579 1552 56581 1604
rect 56525 1550 56581 1552
rect 59021 1604 59077 1606
rect 59021 1552 59023 1604
rect 59023 1552 59075 1604
rect 59075 1552 59077 1604
rect 59021 1550 59077 1552
rect 61517 1604 61573 1606
rect 61517 1552 61519 1604
rect 61519 1552 61571 1604
rect 61571 1552 61573 1604
rect 61517 1550 61573 1552
rect 64013 1604 64069 1606
rect 64013 1552 64015 1604
rect 64015 1552 64067 1604
rect 64067 1552 64069 1604
rect 64013 1550 64069 1552
rect 66509 1604 66565 1606
rect 66509 1552 66511 1604
rect 66511 1552 66563 1604
rect 66563 1552 66565 1604
rect 66509 1550 66565 1552
rect 69005 1604 69061 1606
rect 69005 1552 69007 1604
rect 69007 1552 69059 1604
rect 69059 1552 69061 1604
rect 69005 1550 69061 1552
rect 71501 1604 71557 1606
rect 71501 1552 71503 1604
rect 71503 1552 71555 1604
rect 71555 1552 71557 1604
rect 71501 1550 71557 1552
rect 73997 1604 74053 1606
rect 73997 1552 73999 1604
rect 73999 1552 74051 1604
rect 74051 1552 74053 1604
rect 73997 1550 74053 1552
rect 76493 1604 76549 1606
rect 76493 1552 76495 1604
rect 76495 1552 76547 1604
rect 76547 1552 76549 1604
rect 76493 1550 76549 1552
rect 78989 1604 79045 1606
rect 78989 1552 78991 1604
rect 78991 1552 79043 1604
rect 79043 1552 79045 1604
rect 78989 1550 79045 1552
rect 1602 1167 1658 1169
rect 1602 1115 1604 1167
rect 1604 1115 1656 1167
rect 1656 1115 1658 1167
rect 1602 1113 1658 1115
rect 4098 1167 4154 1169
rect 4098 1115 4100 1167
rect 4100 1115 4152 1167
rect 4152 1115 4154 1167
rect 4098 1113 4154 1115
rect 6594 1167 6650 1169
rect 6594 1115 6596 1167
rect 6596 1115 6648 1167
rect 6648 1115 6650 1167
rect 6594 1113 6650 1115
rect 9090 1167 9146 1169
rect 9090 1115 9092 1167
rect 9092 1115 9144 1167
rect 9144 1115 9146 1167
rect 9090 1113 9146 1115
rect 11586 1167 11642 1169
rect 11586 1115 11588 1167
rect 11588 1115 11640 1167
rect 11640 1115 11642 1167
rect 11586 1113 11642 1115
rect 14082 1167 14138 1169
rect 14082 1115 14084 1167
rect 14084 1115 14136 1167
rect 14136 1115 14138 1167
rect 14082 1113 14138 1115
rect 16578 1167 16634 1169
rect 16578 1115 16580 1167
rect 16580 1115 16632 1167
rect 16632 1115 16634 1167
rect 16578 1113 16634 1115
rect 19074 1167 19130 1169
rect 19074 1115 19076 1167
rect 19076 1115 19128 1167
rect 19128 1115 19130 1167
rect 19074 1113 19130 1115
rect 21570 1167 21626 1169
rect 21570 1115 21572 1167
rect 21572 1115 21624 1167
rect 21624 1115 21626 1167
rect 21570 1113 21626 1115
rect 24066 1167 24122 1169
rect 24066 1115 24068 1167
rect 24068 1115 24120 1167
rect 24120 1115 24122 1167
rect 24066 1113 24122 1115
rect 26562 1167 26618 1169
rect 26562 1115 26564 1167
rect 26564 1115 26616 1167
rect 26616 1115 26618 1167
rect 26562 1113 26618 1115
rect 29058 1167 29114 1169
rect 29058 1115 29060 1167
rect 29060 1115 29112 1167
rect 29112 1115 29114 1167
rect 29058 1113 29114 1115
rect 31554 1167 31610 1169
rect 31554 1115 31556 1167
rect 31556 1115 31608 1167
rect 31608 1115 31610 1167
rect 31554 1113 31610 1115
rect 34050 1167 34106 1169
rect 34050 1115 34052 1167
rect 34052 1115 34104 1167
rect 34104 1115 34106 1167
rect 34050 1113 34106 1115
rect 36546 1167 36602 1169
rect 36546 1115 36548 1167
rect 36548 1115 36600 1167
rect 36600 1115 36602 1167
rect 36546 1113 36602 1115
rect 39042 1167 39098 1169
rect 39042 1115 39044 1167
rect 39044 1115 39096 1167
rect 39096 1115 39098 1167
rect 39042 1113 39098 1115
rect 41538 1167 41594 1169
rect 41538 1115 41540 1167
rect 41540 1115 41592 1167
rect 41592 1115 41594 1167
rect 41538 1113 41594 1115
rect 44034 1167 44090 1169
rect 44034 1115 44036 1167
rect 44036 1115 44088 1167
rect 44088 1115 44090 1167
rect 44034 1113 44090 1115
rect 46530 1167 46586 1169
rect 46530 1115 46532 1167
rect 46532 1115 46584 1167
rect 46584 1115 46586 1167
rect 46530 1113 46586 1115
rect 49026 1167 49082 1169
rect 49026 1115 49028 1167
rect 49028 1115 49080 1167
rect 49080 1115 49082 1167
rect 49026 1113 49082 1115
rect 51522 1167 51578 1169
rect 51522 1115 51524 1167
rect 51524 1115 51576 1167
rect 51576 1115 51578 1167
rect 51522 1113 51578 1115
rect 54018 1167 54074 1169
rect 54018 1115 54020 1167
rect 54020 1115 54072 1167
rect 54072 1115 54074 1167
rect 54018 1113 54074 1115
rect 56514 1167 56570 1169
rect 56514 1115 56516 1167
rect 56516 1115 56568 1167
rect 56568 1115 56570 1167
rect 56514 1113 56570 1115
rect 59010 1167 59066 1169
rect 59010 1115 59012 1167
rect 59012 1115 59064 1167
rect 59064 1115 59066 1167
rect 59010 1113 59066 1115
rect 61506 1167 61562 1169
rect 61506 1115 61508 1167
rect 61508 1115 61560 1167
rect 61560 1115 61562 1167
rect 61506 1113 61562 1115
rect 64002 1167 64058 1169
rect 64002 1115 64004 1167
rect 64004 1115 64056 1167
rect 64056 1115 64058 1167
rect 64002 1113 64058 1115
rect 66498 1167 66554 1169
rect 66498 1115 66500 1167
rect 66500 1115 66552 1167
rect 66552 1115 66554 1167
rect 66498 1113 66554 1115
rect 68994 1167 69050 1169
rect 68994 1115 68996 1167
rect 68996 1115 69048 1167
rect 69048 1115 69050 1167
rect 68994 1113 69050 1115
rect 71490 1167 71546 1169
rect 71490 1115 71492 1167
rect 71492 1115 71544 1167
rect 71544 1115 71546 1167
rect 71490 1113 71546 1115
rect 73986 1167 74042 1169
rect 73986 1115 73988 1167
rect 73988 1115 74040 1167
rect 74040 1115 74042 1167
rect 73986 1113 74042 1115
rect 76482 1167 76538 1169
rect 76482 1115 76484 1167
rect 76484 1115 76536 1167
rect 76536 1115 76538 1167
rect 76482 1113 76538 1115
rect 78978 1167 79034 1169
rect 78978 1115 78980 1167
rect 78980 1115 79032 1167
rect 79032 1115 79034 1167
rect 78978 1113 79034 1115
rect 1723 836 1779 837
rect 1723 784 1725 836
rect 1725 784 1777 836
rect 1777 784 1779 836
rect 1723 781 1779 784
rect 4219 836 4275 837
rect 4219 784 4221 836
rect 4221 784 4273 836
rect 4273 784 4275 836
rect 4219 781 4275 784
rect 6715 836 6771 837
rect 6715 784 6717 836
rect 6717 784 6769 836
rect 6769 784 6771 836
rect 6715 781 6771 784
rect 9211 836 9267 837
rect 9211 784 9213 836
rect 9213 784 9265 836
rect 9265 784 9267 836
rect 9211 781 9267 784
rect 11707 836 11763 837
rect 11707 784 11709 836
rect 11709 784 11761 836
rect 11761 784 11763 836
rect 11707 781 11763 784
rect 14203 836 14259 837
rect 14203 784 14205 836
rect 14205 784 14257 836
rect 14257 784 14259 836
rect 14203 781 14259 784
rect 16699 836 16755 837
rect 16699 784 16701 836
rect 16701 784 16753 836
rect 16753 784 16755 836
rect 16699 781 16755 784
rect 19195 836 19251 837
rect 19195 784 19197 836
rect 19197 784 19249 836
rect 19249 784 19251 836
rect 19195 781 19251 784
rect 21691 836 21747 837
rect 21691 784 21693 836
rect 21693 784 21745 836
rect 21745 784 21747 836
rect 21691 781 21747 784
rect 24187 836 24243 837
rect 24187 784 24189 836
rect 24189 784 24241 836
rect 24241 784 24243 836
rect 24187 781 24243 784
rect 26683 836 26739 837
rect 26683 784 26685 836
rect 26685 784 26737 836
rect 26737 784 26739 836
rect 26683 781 26739 784
rect 29179 836 29235 837
rect 29179 784 29181 836
rect 29181 784 29233 836
rect 29233 784 29235 836
rect 29179 781 29235 784
rect 31675 836 31731 837
rect 31675 784 31677 836
rect 31677 784 31729 836
rect 31729 784 31731 836
rect 31675 781 31731 784
rect 34171 836 34227 837
rect 34171 784 34173 836
rect 34173 784 34225 836
rect 34225 784 34227 836
rect 34171 781 34227 784
rect 36667 836 36723 837
rect 36667 784 36669 836
rect 36669 784 36721 836
rect 36721 784 36723 836
rect 36667 781 36723 784
rect 39163 836 39219 837
rect 39163 784 39165 836
rect 39165 784 39217 836
rect 39217 784 39219 836
rect 39163 781 39219 784
rect 41659 836 41715 837
rect 41659 784 41661 836
rect 41661 784 41713 836
rect 41713 784 41715 836
rect 41659 781 41715 784
rect 44155 836 44211 837
rect 44155 784 44157 836
rect 44157 784 44209 836
rect 44209 784 44211 836
rect 44155 781 44211 784
rect 46651 836 46707 837
rect 46651 784 46653 836
rect 46653 784 46705 836
rect 46705 784 46707 836
rect 46651 781 46707 784
rect 49147 836 49203 837
rect 49147 784 49149 836
rect 49149 784 49201 836
rect 49201 784 49203 836
rect 49147 781 49203 784
rect 51643 836 51699 837
rect 51643 784 51645 836
rect 51645 784 51697 836
rect 51697 784 51699 836
rect 51643 781 51699 784
rect 54139 836 54195 837
rect 54139 784 54141 836
rect 54141 784 54193 836
rect 54193 784 54195 836
rect 54139 781 54195 784
rect 56635 836 56691 837
rect 56635 784 56637 836
rect 56637 784 56689 836
rect 56689 784 56691 836
rect 56635 781 56691 784
rect 59131 836 59187 837
rect 59131 784 59133 836
rect 59133 784 59185 836
rect 59185 784 59187 836
rect 59131 781 59187 784
rect 61627 836 61683 837
rect 61627 784 61629 836
rect 61629 784 61681 836
rect 61681 784 61683 836
rect 61627 781 61683 784
rect 64123 836 64179 837
rect 64123 784 64125 836
rect 64125 784 64177 836
rect 64177 784 64179 836
rect 64123 781 64179 784
rect 66619 836 66675 837
rect 66619 784 66621 836
rect 66621 784 66673 836
rect 66673 784 66675 836
rect 66619 781 66675 784
rect 69115 836 69171 837
rect 69115 784 69117 836
rect 69117 784 69169 836
rect 69169 784 69171 836
rect 69115 781 69171 784
rect 71611 836 71667 837
rect 71611 784 71613 836
rect 71613 784 71665 836
rect 71665 784 71667 836
rect 71611 781 71667 784
rect 74107 836 74163 837
rect 74107 784 74109 836
rect 74109 784 74161 836
rect 74161 784 74163 836
rect 74107 781 74163 784
rect 76603 836 76659 837
rect 76603 784 76605 836
rect 76605 784 76657 836
rect 76657 784 76659 836
rect 76603 781 76659 784
rect 79099 836 79155 837
rect 79099 784 79101 836
rect 79101 784 79153 836
rect 79153 784 79155 836
rect 79099 781 79155 784
rect 1608 633 1664 635
rect 1608 581 1610 633
rect 1610 581 1662 633
rect 1662 581 1664 633
rect 1608 579 1664 581
rect 4104 633 4160 635
rect 4104 581 4106 633
rect 4106 581 4158 633
rect 4158 581 4160 633
rect 4104 579 4160 581
rect 6600 633 6656 635
rect 6600 581 6602 633
rect 6602 581 6654 633
rect 6654 581 6656 633
rect 6600 579 6656 581
rect 9096 633 9152 635
rect 9096 581 9098 633
rect 9098 581 9150 633
rect 9150 581 9152 633
rect 9096 579 9152 581
rect 11592 633 11648 635
rect 11592 581 11594 633
rect 11594 581 11646 633
rect 11646 581 11648 633
rect 11592 579 11648 581
rect 14088 633 14144 635
rect 14088 581 14090 633
rect 14090 581 14142 633
rect 14142 581 14144 633
rect 14088 579 14144 581
rect 16584 633 16640 635
rect 16584 581 16586 633
rect 16586 581 16638 633
rect 16638 581 16640 633
rect 16584 579 16640 581
rect 19080 633 19136 635
rect 19080 581 19082 633
rect 19082 581 19134 633
rect 19134 581 19136 633
rect 19080 579 19136 581
rect 21576 633 21632 635
rect 21576 581 21578 633
rect 21578 581 21630 633
rect 21630 581 21632 633
rect 21576 579 21632 581
rect 24072 633 24128 635
rect 24072 581 24074 633
rect 24074 581 24126 633
rect 24126 581 24128 633
rect 24072 579 24128 581
rect 26568 633 26624 635
rect 26568 581 26570 633
rect 26570 581 26622 633
rect 26622 581 26624 633
rect 26568 579 26624 581
rect 29064 633 29120 635
rect 29064 581 29066 633
rect 29066 581 29118 633
rect 29118 581 29120 633
rect 29064 579 29120 581
rect 31560 633 31616 635
rect 31560 581 31562 633
rect 31562 581 31614 633
rect 31614 581 31616 633
rect 31560 579 31616 581
rect 34056 633 34112 635
rect 34056 581 34058 633
rect 34058 581 34110 633
rect 34110 581 34112 633
rect 34056 579 34112 581
rect 36552 633 36608 635
rect 36552 581 36554 633
rect 36554 581 36606 633
rect 36606 581 36608 633
rect 36552 579 36608 581
rect 39048 633 39104 635
rect 39048 581 39050 633
rect 39050 581 39102 633
rect 39102 581 39104 633
rect 39048 579 39104 581
rect 41544 633 41600 635
rect 41544 581 41546 633
rect 41546 581 41598 633
rect 41598 581 41600 633
rect 41544 579 41600 581
rect 44040 633 44096 635
rect 44040 581 44042 633
rect 44042 581 44094 633
rect 44094 581 44096 633
rect 44040 579 44096 581
rect 46536 633 46592 635
rect 46536 581 46538 633
rect 46538 581 46590 633
rect 46590 581 46592 633
rect 46536 579 46592 581
rect 49032 633 49088 635
rect 49032 581 49034 633
rect 49034 581 49086 633
rect 49086 581 49088 633
rect 49032 579 49088 581
rect 51528 633 51584 635
rect 51528 581 51530 633
rect 51530 581 51582 633
rect 51582 581 51584 633
rect 51528 579 51584 581
rect 54024 633 54080 635
rect 54024 581 54026 633
rect 54026 581 54078 633
rect 54078 581 54080 633
rect 54024 579 54080 581
rect 56520 633 56576 635
rect 56520 581 56522 633
rect 56522 581 56574 633
rect 56574 581 56576 633
rect 56520 579 56576 581
rect 59016 633 59072 635
rect 59016 581 59018 633
rect 59018 581 59070 633
rect 59070 581 59072 633
rect 59016 579 59072 581
rect 61512 633 61568 635
rect 61512 581 61514 633
rect 61514 581 61566 633
rect 61566 581 61568 633
rect 61512 579 61568 581
rect 64008 633 64064 635
rect 64008 581 64010 633
rect 64010 581 64062 633
rect 64062 581 64064 633
rect 64008 579 64064 581
rect 66504 633 66560 635
rect 66504 581 66506 633
rect 66506 581 66558 633
rect 66558 581 66560 633
rect 66504 579 66560 581
rect 69000 633 69056 635
rect 69000 581 69002 633
rect 69002 581 69054 633
rect 69054 581 69056 633
rect 69000 579 69056 581
rect 71496 633 71552 635
rect 71496 581 71498 633
rect 71498 581 71550 633
rect 71550 581 71552 633
rect 71496 579 71552 581
rect 73992 633 74048 635
rect 73992 581 73994 633
rect 73994 581 74046 633
rect 74046 581 74048 633
rect 73992 579 74048 581
rect 76488 633 76544 635
rect 76488 581 76490 633
rect 76490 581 76542 633
rect 76542 581 76544 633
rect 76488 579 76544 581
rect 78984 633 79040 635
rect 78984 581 78986 633
rect 78986 581 79038 633
rect 79038 581 79040 633
rect 78984 579 79040 581
rect 1622 217 1678 219
rect 1622 165 1624 217
rect 1624 165 1676 217
rect 1676 165 1678 217
rect 1622 163 1678 165
rect 4118 217 4174 219
rect 4118 165 4120 217
rect 4120 165 4172 217
rect 4172 165 4174 217
rect 4118 163 4174 165
rect 6614 217 6670 219
rect 6614 165 6616 217
rect 6616 165 6668 217
rect 6668 165 6670 217
rect 6614 163 6670 165
rect 9110 217 9166 219
rect 9110 165 9112 217
rect 9112 165 9164 217
rect 9164 165 9166 217
rect 9110 163 9166 165
rect 11606 217 11662 219
rect 11606 165 11608 217
rect 11608 165 11660 217
rect 11660 165 11662 217
rect 11606 163 11662 165
rect 14102 217 14158 219
rect 14102 165 14104 217
rect 14104 165 14156 217
rect 14156 165 14158 217
rect 14102 163 14158 165
rect 16598 217 16654 219
rect 16598 165 16600 217
rect 16600 165 16652 217
rect 16652 165 16654 217
rect 16598 163 16654 165
rect 19094 217 19150 219
rect 19094 165 19096 217
rect 19096 165 19148 217
rect 19148 165 19150 217
rect 19094 163 19150 165
rect 21590 217 21646 219
rect 21590 165 21592 217
rect 21592 165 21644 217
rect 21644 165 21646 217
rect 21590 163 21646 165
rect 24086 217 24142 219
rect 24086 165 24088 217
rect 24088 165 24140 217
rect 24140 165 24142 217
rect 24086 163 24142 165
rect 26582 217 26638 219
rect 26582 165 26584 217
rect 26584 165 26636 217
rect 26636 165 26638 217
rect 26582 163 26638 165
rect 29078 217 29134 219
rect 29078 165 29080 217
rect 29080 165 29132 217
rect 29132 165 29134 217
rect 29078 163 29134 165
rect 31574 217 31630 219
rect 31574 165 31576 217
rect 31576 165 31628 217
rect 31628 165 31630 217
rect 31574 163 31630 165
rect 34070 217 34126 219
rect 34070 165 34072 217
rect 34072 165 34124 217
rect 34124 165 34126 217
rect 34070 163 34126 165
rect 36566 217 36622 219
rect 36566 165 36568 217
rect 36568 165 36620 217
rect 36620 165 36622 217
rect 36566 163 36622 165
rect 39062 217 39118 219
rect 39062 165 39064 217
rect 39064 165 39116 217
rect 39116 165 39118 217
rect 39062 163 39118 165
rect 41558 217 41614 219
rect 41558 165 41560 217
rect 41560 165 41612 217
rect 41612 165 41614 217
rect 41558 163 41614 165
rect 44054 217 44110 219
rect 44054 165 44056 217
rect 44056 165 44108 217
rect 44108 165 44110 217
rect 44054 163 44110 165
rect 46550 217 46606 219
rect 46550 165 46552 217
rect 46552 165 46604 217
rect 46604 165 46606 217
rect 46550 163 46606 165
rect 49046 217 49102 219
rect 49046 165 49048 217
rect 49048 165 49100 217
rect 49100 165 49102 217
rect 49046 163 49102 165
rect 51542 217 51598 219
rect 51542 165 51544 217
rect 51544 165 51596 217
rect 51596 165 51598 217
rect 51542 163 51598 165
rect 54038 217 54094 219
rect 54038 165 54040 217
rect 54040 165 54092 217
rect 54092 165 54094 217
rect 54038 163 54094 165
rect 56534 217 56590 219
rect 56534 165 56536 217
rect 56536 165 56588 217
rect 56588 165 56590 217
rect 56534 163 56590 165
rect 59030 217 59086 219
rect 59030 165 59032 217
rect 59032 165 59084 217
rect 59084 165 59086 217
rect 59030 163 59086 165
rect 61526 217 61582 219
rect 61526 165 61528 217
rect 61528 165 61580 217
rect 61580 165 61582 217
rect 61526 163 61582 165
rect 64022 217 64078 219
rect 64022 165 64024 217
rect 64024 165 64076 217
rect 64076 165 64078 217
rect 64022 163 64078 165
rect 66518 217 66574 219
rect 66518 165 66520 217
rect 66520 165 66572 217
rect 66572 165 66574 217
rect 66518 163 66574 165
rect 69014 217 69070 219
rect 69014 165 69016 217
rect 69016 165 69068 217
rect 69068 165 69070 217
rect 69014 163 69070 165
rect 71510 217 71566 219
rect 71510 165 71512 217
rect 71512 165 71564 217
rect 71564 165 71566 217
rect 71510 163 71566 165
rect 74006 217 74062 219
rect 74006 165 74008 217
rect 74008 165 74060 217
rect 74060 165 74062 217
rect 74006 163 74062 165
rect 76502 217 76558 219
rect 76502 165 76504 217
rect 76504 165 76556 217
rect 76556 165 76558 217
rect 76502 163 76558 165
rect 78998 217 79054 219
rect 78998 165 79000 217
rect 79000 165 79052 217
rect 79052 165 79054 217
rect 78998 163 79054 165
<< metal3 >>
rect 1592 1606 1690 1627
rect 1592 1550 1613 1606
rect 1669 1550 1690 1606
rect 1592 1529 1690 1550
rect 4088 1606 4186 1627
rect 4088 1550 4109 1606
rect 4165 1550 4186 1606
rect 4088 1529 4186 1550
rect 6584 1606 6682 1627
rect 6584 1550 6605 1606
rect 6661 1550 6682 1606
rect 6584 1529 6682 1550
rect 9080 1606 9178 1627
rect 9080 1550 9101 1606
rect 9157 1550 9178 1606
rect 9080 1529 9178 1550
rect 11576 1606 11674 1627
rect 11576 1550 11597 1606
rect 11653 1550 11674 1606
rect 11576 1529 11674 1550
rect 14072 1606 14170 1627
rect 14072 1550 14093 1606
rect 14149 1550 14170 1606
rect 14072 1529 14170 1550
rect 16568 1606 16666 1627
rect 16568 1550 16589 1606
rect 16645 1550 16666 1606
rect 16568 1529 16666 1550
rect 19064 1606 19162 1627
rect 19064 1550 19085 1606
rect 19141 1550 19162 1606
rect 19064 1529 19162 1550
rect 21560 1606 21658 1627
rect 21560 1550 21581 1606
rect 21637 1550 21658 1606
rect 21560 1529 21658 1550
rect 24056 1606 24154 1627
rect 24056 1550 24077 1606
rect 24133 1550 24154 1606
rect 24056 1529 24154 1550
rect 26552 1606 26650 1627
rect 26552 1550 26573 1606
rect 26629 1550 26650 1606
rect 26552 1529 26650 1550
rect 29048 1606 29146 1627
rect 29048 1550 29069 1606
rect 29125 1550 29146 1606
rect 29048 1529 29146 1550
rect 31544 1606 31642 1627
rect 31544 1550 31565 1606
rect 31621 1550 31642 1606
rect 31544 1529 31642 1550
rect 34040 1606 34138 1627
rect 34040 1550 34061 1606
rect 34117 1550 34138 1606
rect 34040 1529 34138 1550
rect 36536 1606 36634 1627
rect 36536 1550 36557 1606
rect 36613 1550 36634 1606
rect 36536 1529 36634 1550
rect 39032 1606 39130 1627
rect 39032 1550 39053 1606
rect 39109 1550 39130 1606
rect 39032 1529 39130 1550
rect 41528 1606 41626 1627
rect 41528 1550 41549 1606
rect 41605 1550 41626 1606
rect 41528 1529 41626 1550
rect 44024 1606 44122 1627
rect 44024 1550 44045 1606
rect 44101 1550 44122 1606
rect 44024 1529 44122 1550
rect 46520 1606 46618 1627
rect 46520 1550 46541 1606
rect 46597 1550 46618 1606
rect 46520 1529 46618 1550
rect 49016 1606 49114 1627
rect 49016 1550 49037 1606
rect 49093 1550 49114 1606
rect 49016 1529 49114 1550
rect 51512 1606 51610 1627
rect 51512 1550 51533 1606
rect 51589 1550 51610 1606
rect 51512 1529 51610 1550
rect 54008 1606 54106 1627
rect 54008 1550 54029 1606
rect 54085 1550 54106 1606
rect 54008 1529 54106 1550
rect 56504 1606 56602 1627
rect 56504 1550 56525 1606
rect 56581 1550 56602 1606
rect 56504 1529 56602 1550
rect 59000 1606 59098 1627
rect 59000 1550 59021 1606
rect 59077 1550 59098 1606
rect 59000 1529 59098 1550
rect 61496 1606 61594 1627
rect 61496 1550 61517 1606
rect 61573 1550 61594 1606
rect 61496 1529 61594 1550
rect 63992 1606 64090 1627
rect 63992 1550 64013 1606
rect 64069 1550 64090 1606
rect 63992 1529 64090 1550
rect 66488 1606 66586 1627
rect 66488 1550 66509 1606
rect 66565 1550 66586 1606
rect 66488 1529 66586 1550
rect 68984 1606 69082 1627
rect 68984 1550 69005 1606
rect 69061 1550 69082 1606
rect 68984 1529 69082 1550
rect 71480 1606 71578 1627
rect 71480 1550 71501 1606
rect 71557 1550 71578 1606
rect 71480 1529 71578 1550
rect 73976 1606 74074 1627
rect 73976 1550 73997 1606
rect 74053 1550 74074 1606
rect 73976 1529 74074 1550
rect 76472 1606 76570 1627
rect 76472 1550 76493 1606
rect 76549 1550 76570 1606
rect 76472 1529 76570 1550
rect 78968 1606 79066 1627
rect 78968 1550 78989 1606
rect 79045 1550 79066 1606
rect 78968 1529 79066 1550
rect 1581 1169 1679 1190
rect 1581 1113 1602 1169
rect 1658 1113 1679 1169
rect 1581 1092 1679 1113
rect 4077 1169 4175 1190
rect 4077 1113 4098 1169
rect 4154 1113 4175 1169
rect 4077 1092 4175 1113
rect 6573 1169 6671 1190
rect 6573 1113 6594 1169
rect 6650 1113 6671 1169
rect 6573 1092 6671 1113
rect 9069 1169 9167 1190
rect 9069 1113 9090 1169
rect 9146 1113 9167 1169
rect 9069 1092 9167 1113
rect 11565 1169 11663 1190
rect 11565 1113 11586 1169
rect 11642 1113 11663 1169
rect 11565 1092 11663 1113
rect 14061 1169 14159 1190
rect 14061 1113 14082 1169
rect 14138 1113 14159 1169
rect 14061 1092 14159 1113
rect 16557 1169 16655 1190
rect 16557 1113 16578 1169
rect 16634 1113 16655 1169
rect 16557 1092 16655 1113
rect 19053 1169 19151 1190
rect 19053 1113 19074 1169
rect 19130 1113 19151 1169
rect 19053 1092 19151 1113
rect 21549 1169 21647 1190
rect 21549 1113 21570 1169
rect 21626 1113 21647 1169
rect 21549 1092 21647 1113
rect 24045 1169 24143 1190
rect 24045 1113 24066 1169
rect 24122 1113 24143 1169
rect 24045 1092 24143 1113
rect 26541 1169 26639 1190
rect 26541 1113 26562 1169
rect 26618 1113 26639 1169
rect 26541 1092 26639 1113
rect 29037 1169 29135 1190
rect 29037 1113 29058 1169
rect 29114 1113 29135 1169
rect 29037 1092 29135 1113
rect 31533 1169 31631 1190
rect 31533 1113 31554 1169
rect 31610 1113 31631 1169
rect 31533 1092 31631 1113
rect 34029 1169 34127 1190
rect 34029 1113 34050 1169
rect 34106 1113 34127 1169
rect 34029 1092 34127 1113
rect 36525 1169 36623 1190
rect 36525 1113 36546 1169
rect 36602 1113 36623 1169
rect 36525 1092 36623 1113
rect 39021 1169 39119 1190
rect 39021 1113 39042 1169
rect 39098 1113 39119 1169
rect 39021 1092 39119 1113
rect 41517 1169 41615 1190
rect 41517 1113 41538 1169
rect 41594 1113 41615 1169
rect 41517 1092 41615 1113
rect 44013 1169 44111 1190
rect 44013 1113 44034 1169
rect 44090 1113 44111 1169
rect 44013 1092 44111 1113
rect 46509 1169 46607 1190
rect 46509 1113 46530 1169
rect 46586 1113 46607 1169
rect 46509 1092 46607 1113
rect 49005 1169 49103 1190
rect 49005 1113 49026 1169
rect 49082 1113 49103 1169
rect 49005 1092 49103 1113
rect 51501 1169 51599 1190
rect 51501 1113 51522 1169
rect 51578 1113 51599 1169
rect 51501 1092 51599 1113
rect 53997 1169 54095 1190
rect 53997 1113 54018 1169
rect 54074 1113 54095 1169
rect 53997 1092 54095 1113
rect 56493 1169 56591 1190
rect 56493 1113 56514 1169
rect 56570 1113 56591 1169
rect 56493 1092 56591 1113
rect 58989 1169 59087 1190
rect 58989 1113 59010 1169
rect 59066 1113 59087 1169
rect 58989 1092 59087 1113
rect 61485 1169 61583 1190
rect 61485 1113 61506 1169
rect 61562 1113 61583 1169
rect 61485 1092 61583 1113
rect 63981 1169 64079 1190
rect 63981 1113 64002 1169
rect 64058 1113 64079 1169
rect 63981 1092 64079 1113
rect 66477 1169 66575 1190
rect 66477 1113 66498 1169
rect 66554 1113 66575 1169
rect 66477 1092 66575 1113
rect 68973 1169 69071 1190
rect 68973 1113 68994 1169
rect 69050 1113 69071 1169
rect 68973 1092 69071 1113
rect 71469 1169 71567 1190
rect 71469 1113 71490 1169
rect 71546 1113 71567 1169
rect 71469 1092 71567 1113
rect 73965 1169 74063 1190
rect 73965 1113 73986 1169
rect 74042 1113 74063 1169
rect 73965 1092 74063 1113
rect 76461 1169 76559 1190
rect 76461 1113 76482 1169
rect 76538 1113 76559 1169
rect 76461 1092 76559 1113
rect 78957 1169 79055 1190
rect 78957 1113 78978 1169
rect 79034 1113 79055 1169
rect 78957 1092 79055 1113
rect 1702 837 1800 858
rect 1702 781 1723 837
rect 1779 781 1800 837
rect 1702 760 1800 781
rect 4198 837 4296 858
rect 4198 781 4219 837
rect 4275 781 4296 837
rect 4198 760 4296 781
rect 6694 837 6792 858
rect 6694 781 6715 837
rect 6771 781 6792 837
rect 6694 760 6792 781
rect 9190 837 9288 858
rect 9190 781 9211 837
rect 9267 781 9288 837
rect 9190 760 9288 781
rect 11686 837 11784 858
rect 11686 781 11707 837
rect 11763 781 11784 837
rect 11686 760 11784 781
rect 14182 837 14280 858
rect 14182 781 14203 837
rect 14259 781 14280 837
rect 14182 760 14280 781
rect 16678 837 16776 858
rect 16678 781 16699 837
rect 16755 781 16776 837
rect 16678 760 16776 781
rect 19174 837 19272 858
rect 19174 781 19195 837
rect 19251 781 19272 837
rect 19174 760 19272 781
rect 21670 837 21768 858
rect 21670 781 21691 837
rect 21747 781 21768 837
rect 21670 760 21768 781
rect 24166 837 24264 858
rect 24166 781 24187 837
rect 24243 781 24264 837
rect 24166 760 24264 781
rect 26662 837 26760 858
rect 26662 781 26683 837
rect 26739 781 26760 837
rect 26662 760 26760 781
rect 29158 837 29256 858
rect 29158 781 29179 837
rect 29235 781 29256 837
rect 29158 760 29256 781
rect 31654 837 31752 858
rect 31654 781 31675 837
rect 31731 781 31752 837
rect 31654 760 31752 781
rect 34150 837 34248 858
rect 34150 781 34171 837
rect 34227 781 34248 837
rect 34150 760 34248 781
rect 36646 837 36744 858
rect 36646 781 36667 837
rect 36723 781 36744 837
rect 36646 760 36744 781
rect 39142 837 39240 858
rect 39142 781 39163 837
rect 39219 781 39240 837
rect 39142 760 39240 781
rect 41638 837 41736 858
rect 41638 781 41659 837
rect 41715 781 41736 837
rect 41638 760 41736 781
rect 44134 837 44232 858
rect 44134 781 44155 837
rect 44211 781 44232 837
rect 44134 760 44232 781
rect 46630 837 46728 858
rect 46630 781 46651 837
rect 46707 781 46728 837
rect 46630 760 46728 781
rect 49126 837 49224 858
rect 49126 781 49147 837
rect 49203 781 49224 837
rect 49126 760 49224 781
rect 51622 837 51720 858
rect 51622 781 51643 837
rect 51699 781 51720 837
rect 51622 760 51720 781
rect 54118 837 54216 858
rect 54118 781 54139 837
rect 54195 781 54216 837
rect 54118 760 54216 781
rect 56614 837 56712 858
rect 56614 781 56635 837
rect 56691 781 56712 837
rect 56614 760 56712 781
rect 59110 837 59208 858
rect 59110 781 59131 837
rect 59187 781 59208 837
rect 59110 760 59208 781
rect 61606 837 61704 858
rect 61606 781 61627 837
rect 61683 781 61704 837
rect 61606 760 61704 781
rect 64102 837 64200 858
rect 64102 781 64123 837
rect 64179 781 64200 837
rect 64102 760 64200 781
rect 66598 837 66696 858
rect 66598 781 66619 837
rect 66675 781 66696 837
rect 66598 760 66696 781
rect 69094 837 69192 858
rect 69094 781 69115 837
rect 69171 781 69192 837
rect 69094 760 69192 781
rect 71590 837 71688 858
rect 71590 781 71611 837
rect 71667 781 71688 837
rect 71590 760 71688 781
rect 74086 837 74184 858
rect 74086 781 74107 837
rect 74163 781 74184 837
rect 74086 760 74184 781
rect 76582 837 76680 858
rect 76582 781 76603 837
rect 76659 781 76680 837
rect 76582 760 76680 781
rect 79078 837 79176 858
rect 79078 781 79099 837
rect 79155 781 79176 837
rect 79078 760 79176 781
rect 1587 635 1685 656
rect 1587 579 1608 635
rect 1664 579 1685 635
rect 1587 558 1685 579
rect 4083 635 4181 656
rect 4083 579 4104 635
rect 4160 579 4181 635
rect 4083 558 4181 579
rect 6579 635 6677 656
rect 6579 579 6600 635
rect 6656 579 6677 635
rect 6579 558 6677 579
rect 9075 635 9173 656
rect 9075 579 9096 635
rect 9152 579 9173 635
rect 9075 558 9173 579
rect 11571 635 11669 656
rect 11571 579 11592 635
rect 11648 579 11669 635
rect 11571 558 11669 579
rect 14067 635 14165 656
rect 14067 579 14088 635
rect 14144 579 14165 635
rect 14067 558 14165 579
rect 16563 635 16661 656
rect 16563 579 16584 635
rect 16640 579 16661 635
rect 16563 558 16661 579
rect 19059 635 19157 656
rect 19059 579 19080 635
rect 19136 579 19157 635
rect 19059 558 19157 579
rect 21555 635 21653 656
rect 21555 579 21576 635
rect 21632 579 21653 635
rect 21555 558 21653 579
rect 24051 635 24149 656
rect 24051 579 24072 635
rect 24128 579 24149 635
rect 24051 558 24149 579
rect 26547 635 26645 656
rect 26547 579 26568 635
rect 26624 579 26645 635
rect 26547 558 26645 579
rect 29043 635 29141 656
rect 29043 579 29064 635
rect 29120 579 29141 635
rect 29043 558 29141 579
rect 31539 635 31637 656
rect 31539 579 31560 635
rect 31616 579 31637 635
rect 31539 558 31637 579
rect 34035 635 34133 656
rect 34035 579 34056 635
rect 34112 579 34133 635
rect 34035 558 34133 579
rect 36531 635 36629 656
rect 36531 579 36552 635
rect 36608 579 36629 635
rect 36531 558 36629 579
rect 39027 635 39125 656
rect 39027 579 39048 635
rect 39104 579 39125 635
rect 39027 558 39125 579
rect 41523 635 41621 656
rect 41523 579 41544 635
rect 41600 579 41621 635
rect 41523 558 41621 579
rect 44019 635 44117 656
rect 44019 579 44040 635
rect 44096 579 44117 635
rect 44019 558 44117 579
rect 46515 635 46613 656
rect 46515 579 46536 635
rect 46592 579 46613 635
rect 46515 558 46613 579
rect 49011 635 49109 656
rect 49011 579 49032 635
rect 49088 579 49109 635
rect 49011 558 49109 579
rect 51507 635 51605 656
rect 51507 579 51528 635
rect 51584 579 51605 635
rect 51507 558 51605 579
rect 54003 635 54101 656
rect 54003 579 54024 635
rect 54080 579 54101 635
rect 54003 558 54101 579
rect 56499 635 56597 656
rect 56499 579 56520 635
rect 56576 579 56597 635
rect 56499 558 56597 579
rect 58995 635 59093 656
rect 58995 579 59016 635
rect 59072 579 59093 635
rect 58995 558 59093 579
rect 61491 635 61589 656
rect 61491 579 61512 635
rect 61568 579 61589 635
rect 61491 558 61589 579
rect 63987 635 64085 656
rect 63987 579 64008 635
rect 64064 579 64085 635
rect 63987 558 64085 579
rect 66483 635 66581 656
rect 66483 579 66504 635
rect 66560 579 66581 635
rect 66483 558 66581 579
rect 68979 635 69077 656
rect 68979 579 69000 635
rect 69056 579 69077 635
rect 68979 558 69077 579
rect 71475 635 71573 656
rect 71475 579 71496 635
rect 71552 579 71573 635
rect 71475 558 71573 579
rect 73971 635 74069 656
rect 73971 579 73992 635
rect 74048 579 74069 635
rect 73971 558 74069 579
rect 76467 635 76565 656
rect 76467 579 76488 635
rect 76544 579 76565 635
rect 76467 558 76565 579
rect 78963 635 79061 656
rect 78963 579 78984 635
rect 79040 579 79061 635
rect 78963 558 79061 579
rect 1601 219 1699 240
rect 1601 163 1622 219
rect 1678 163 1699 219
rect 1601 142 1699 163
rect 4097 219 4195 240
rect 4097 163 4118 219
rect 4174 163 4195 219
rect 4097 142 4195 163
rect 6593 219 6691 240
rect 6593 163 6614 219
rect 6670 163 6691 219
rect 6593 142 6691 163
rect 9089 219 9187 240
rect 9089 163 9110 219
rect 9166 163 9187 219
rect 9089 142 9187 163
rect 11585 219 11683 240
rect 11585 163 11606 219
rect 11662 163 11683 219
rect 11585 142 11683 163
rect 14081 219 14179 240
rect 14081 163 14102 219
rect 14158 163 14179 219
rect 14081 142 14179 163
rect 16577 219 16675 240
rect 16577 163 16598 219
rect 16654 163 16675 219
rect 16577 142 16675 163
rect 19073 219 19171 240
rect 19073 163 19094 219
rect 19150 163 19171 219
rect 19073 142 19171 163
rect 21569 219 21667 240
rect 21569 163 21590 219
rect 21646 163 21667 219
rect 21569 142 21667 163
rect 24065 219 24163 240
rect 24065 163 24086 219
rect 24142 163 24163 219
rect 24065 142 24163 163
rect 26561 219 26659 240
rect 26561 163 26582 219
rect 26638 163 26659 219
rect 26561 142 26659 163
rect 29057 219 29155 240
rect 29057 163 29078 219
rect 29134 163 29155 219
rect 29057 142 29155 163
rect 31553 219 31651 240
rect 31553 163 31574 219
rect 31630 163 31651 219
rect 31553 142 31651 163
rect 34049 219 34147 240
rect 34049 163 34070 219
rect 34126 163 34147 219
rect 34049 142 34147 163
rect 36545 219 36643 240
rect 36545 163 36566 219
rect 36622 163 36643 219
rect 36545 142 36643 163
rect 39041 219 39139 240
rect 39041 163 39062 219
rect 39118 163 39139 219
rect 39041 142 39139 163
rect 41537 219 41635 240
rect 41537 163 41558 219
rect 41614 163 41635 219
rect 41537 142 41635 163
rect 44033 219 44131 240
rect 44033 163 44054 219
rect 44110 163 44131 219
rect 44033 142 44131 163
rect 46529 219 46627 240
rect 46529 163 46550 219
rect 46606 163 46627 219
rect 46529 142 46627 163
rect 49025 219 49123 240
rect 49025 163 49046 219
rect 49102 163 49123 219
rect 49025 142 49123 163
rect 51521 219 51619 240
rect 51521 163 51542 219
rect 51598 163 51619 219
rect 51521 142 51619 163
rect 54017 219 54115 240
rect 54017 163 54038 219
rect 54094 163 54115 219
rect 54017 142 54115 163
rect 56513 219 56611 240
rect 56513 163 56534 219
rect 56590 163 56611 219
rect 56513 142 56611 163
rect 59009 219 59107 240
rect 59009 163 59030 219
rect 59086 163 59107 219
rect 59009 142 59107 163
rect 61505 219 61603 240
rect 61505 163 61526 219
rect 61582 163 61603 219
rect 61505 142 61603 163
rect 64001 219 64099 240
rect 64001 163 64022 219
rect 64078 163 64099 219
rect 64001 142 64099 163
rect 66497 219 66595 240
rect 66497 163 66518 219
rect 66574 163 66595 219
rect 66497 142 66595 163
rect 68993 219 69091 240
rect 68993 163 69014 219
rect 69070 163 69091 219
rect 68993 142 69091 163
rect 71489 219 71587 240
rect 71489 163 71510 219
rect 71566 163 71587 219
rect 71489 142 71587 163
rect 73985 219 74083 240
rect 73985 163 74006 219
rect 74062 163 74083 219
rect 73985 142 74083 163
rect 76481 219 76579 240
rect 76481 163 76502 219
rect 76558 163 76579 219
rect 76481 142 76579 163
rect 78977 219 79075 240
rect 78977 163 78998 219
rect 79054 163 79075 219
rect 78977 142 79075 163
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_0
timestamp 1701704242
transform 1 0 18846 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_1
timestamp 1701704242
transform 1 0 16350 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_2
timestamp 1701704242
transform 1 0 13854 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_3
timestamp 1701704242
transform 1 0 11358 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_4
timestamp 1701704242
transform 1 0 8862 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_5
timestamp 1701704242
transform 1 0 6366 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_6
timestamp 1701704242
transform 1 0 3870 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_7
timestamp 1701704242
transform 1 0 1374 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_8
timestamp 1701704242
transform 1 0 38814 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_9
timestamp 1701704242
transform 1 0 36318 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_10
timestamp 1701704242
transform 1 0 33822 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_11
timestamp 1701704242
transform 1 0 31326 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_12
timestamp 1701704242
transform 1 0 28830 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_13
timestamp 1701704242
transform 1 0 26334 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_14
timestamp 1701704242
transform 1 0 23838 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_15
timestamp 1701704242
transform 1 0 21342 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_16
timestamp 1701704242
transform 1 0 58782 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_17
timestamp 1701704242
transform 1 0 56286 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_18
timestamp 1701704242
transform 1 0 53790 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_19
timestamp 1701704242
transform 1 0 51294 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_20
timestamp 1701704242
transform 1 0 48798 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_21
timestamp 1701704242
transform 1 0 46302 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_22
timestamp 1701704242
transform 1 0 43806 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_23
timestamp 1701704242
transform 1 0 41310 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_24
timestamp 1701704242
transform 1 0 78750 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_25
timestamp 1701704242
transform 1 0 76254 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_26
timestamp 1701704242
transform 1 0 73758 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_27
timestamp 1701704242
transform 1 0 71262 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_28
timestamp 1701704242
transform 1 0 68766 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_29
timestamp 1701704242
transform 1 0 66270 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_30
timestamp 1701704242
transform 1 0 63774 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_2  sky130_fd_bd_sram__openram_write_driver_31
timestamp 1701704242
transform 1 0 61278 0 1 0
box -376 4 880 2011
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_0
timestamp 1701704242
transform 1 0 14090 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_1
timestamp 1701704242
transform 1 0 14084 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_2
timestamp 1701704242
transform 1 0 14104 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_3
timestamp 1701704242
transform 1 0 11599 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_4
timestamp 1701704242
transform 1 0 11709 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_5
timestamp 1701704242
transform 1 0 11594 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_6
timestamp 1701704242
transform 1 0 11588 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_7
timestamp 1701704242
transform 1 0 11608 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_8
timestamp 1701704242
transform 1 0 9103 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_9
timestamp 1701704242
transform 1 0 9213 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_10
timestamp 1701704242
transform 1 0 9098 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_11
timestamp 1701704242
transform 1 0 9092 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_12
timestamp 1701704242
transform 1 0 9112 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_13
timestamp 1701704242
transform 1 0 6607 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_14
timestamp 1701704242
transform 1 0 6717 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_15
timestamp 1701704242
transform 1 0 6602 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_16
timestamp 1701704242
transform 1 0 6596 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_17
timestamp 1701704242
transform 1 0 6616 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_18
timestamp 1701704242
transform 1 0 4111 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_19
timestamp 1701704242
transform 1 0 4221 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_20
timestamp 1701704242
transform 1 0 4106 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_21
timestamp 1701704242
transform 1 0 4100 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_22
timestamp 1701704242
transform 1 0 4120 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_23
timestamp 1701704242
transform 1 0 1615 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_24
timestamp 1701704242
transform 1 0 1725 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_25
timestamp 1701704242
transform 1 0 1610 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_26
timestamp 1701704242
transform 1 0 1604 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_27
timestamp 1701704242
transform 1 0 1624 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_28
timestamp 1701704242
transform 1 0 19087 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_29
timestamp 1701704242
transform 1 0 19197 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_30
timestamp 1701704242
transform 1 0 19082 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_31
timestamp 1701704242
transform 1 0 19076 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_32
timestamp 1701704242
transform 1 0 19096 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_33
timestamp 1701704242
transform 1 0 16591 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_34
timestamp 1701704242
transform 1 0 16701 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_35
timestamp 1701704242
transform 1 0 16586 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_36
timestamp 1701704242
transform 1 0 16580 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_37
timestamp 1701704242
transform 1 0 16600 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_38
timestamp 1701704242
transform 1 0 14095 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_39
timestamp 1701704242
transform 1 0 14205 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_40
timestamp 1701704242
transform 1 0 36548 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_41
timestamp 1701704242
transform 1 0 36568 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_42
timestamp 1701704242
transform 1 0 34063 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_43
timestamp 1701704242
transform 1 0 34173 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_44
timestamp 1701704242
transform 1 0 34058 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_45
timestamp 1701704242
transform 1 0 34052 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_46
timestamp 1701704242
transform 1 0 34072 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_47
timestamp 1701704242
transform 1 0 31567 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_48
timestamp 1701704242
transform 1 0 31677 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_49
timestamp 1701704242
transform 1 0 31562 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_50
timestamp 1701704242
transform 1 0 31556 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_51
timestamp 1701704242
transform 1 0 31576 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_52
timestamp 1701704242
transform 1 0 29071 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_53
timestamp 1701704242
transform 1 0 29181 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_54
timestamp 1701704242
transform 1 0 29066 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_55
timestamp 1701704242
transform 1 0 29060 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_56
timestamp 1701704242
transform 1 0 29080 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_57
timestamp 1701704242
transform 1 0 26575 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_58
timestamp 1701704242
transform 1 0 26685 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_59
timestamp 1701704242
transform 1 0 26570 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_60
timestamp 1701704242
transform 1 0 26564 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_61
timestamp 1701704242
transform 1 0 26584 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_62
timestamp 1701704242
transform 1 0 24079 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_63
timestamp 1701704242
transform 1 0 24189 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_64
timestamp 1701704242
transform 1 0 24074 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_65
timestamp 1701704242
transform 1 0 24068 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_66
timestamp 1701704242
transform 1 0 24088 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_67
timestamp 1701704242
transform 1 0 21583 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_68
timestamp 1701704242
transform 1 0 21693 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_69
timestamp 1701704242
transform 1 0 21578 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_70
timestamp 1701704242
transform 1 0 21572 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_71
timestamp 1701704242
transform 1 0 21592 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_72
timestamp 1701704242
transform 1 0 39055 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_73
timestamp 1701704242
transform 1 0 39165 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_74
timestamp 1701704242
transform 1 0 39050 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_75
timestamp 1701704242
transform 1 0 39044 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_76
timestamp 1701704242
transform 1 0 39064 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_77
timestamp 1701704242
transform 1 0 36559 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_78
timestamp 1701704242
transform 1 0 36669 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_79
timestamp 1701704242
transform 1 0 36554 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_80
timestamp 1701704242
transform 1 0 59032 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_81
timestamp 1701704242
transform 1 0 56527 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_82
timestamp 1701704242
transform 1 0 56637 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_83
timestamp 1701704242
transform 1 0 56522 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_84
timestamp 1701704242
transform 1 0 56516 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_85
timestamp 1701704242
transform 1 0 56536 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_86
timestamp 1701704242
transform 1 0 54031 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_87
timestamp 1701704242
transform 1 0 54141 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_88
timestamp 1701704242
transform 1 0 54026 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_89
timestamp 1701704242
transform 1 0 54020 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_90
timestamp 1701704242
transform 1 0 54040 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_91
timestamp 1701704242
transform 1 0 51535 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_92
timestamp 1701704242
transform 1 0 51645 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_93
timestamp 1701704242
transform 1 0 51530 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_94
timestamp 1701704242
transform 1 0 51524 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_95
timestamp 1701704242
transform 1 0 51544 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_96
timestamp 1701704242
transform 1 0 49039 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_97
timestamp 1701704242
transform 1 0 49149 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_98
timestamp 1701704242
transform 1 0 49034 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_99
timestamp 1701704242
transform 1 0 49028 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_100
timestamp 1701704242
transform 1 0 49048 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_101
timestamp 1701704242
transform 1 0 46543 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_102
timestamp 1701704242
transform 1 0 46653 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_103
timestamp 1701704242
transform 1 0 46538 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_104
timestamp 1701704242
transform 1 0 46532 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_105
timestamp 1701704242
transform 1 0 46552 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_106
timestamp 1701704242
transform 1 0 44047 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_107
timestamp 1701704242
transform 1 0 44157 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_108
timestamp 1701704242
transform 1 0 44042 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_109
timestamp 1701704242
transform 1 0 44036 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_110
timestamp 1701704242
transform 1 0 44056 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_111
timestamp 1701704242
transform 1 0 41551 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_112
timestamp 1701704242
transform 1 0 41661 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_113
timestamp 1701704242
transform 1 0 41546 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_114
timestamp 1701704242
transform 1 0 41540 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_115
timestamp 1701704242
transform 1 0 41560 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_116
timestamp 1701704242
transform 1 0 59023 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_117
timestamp 1701704242
transform 1 0 59133 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_118
timestamp 1701704242
transform 1 0 59018 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_119
timestamp 1701704242
transform 1 0 59012 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_120
timestamp 1701704242
transform 1 0 78991 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_121
timestamp 1701704242
transform 1 0 79101 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_122
timestamp 1701704242
transform 1 0 78986 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_123
timestamp 1701704242
transform 1 0 78980 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_124
timestamp 1701704242
transform 1 0 79000 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_125
timestamp 1701704242
transform 1 0 76495 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_126
timestamp 1701704242
transform 1 0 76605 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_127
timestamp 1701704242
transform 1 0 76490 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_128
timestamp 1701704242
transform 1 0 76484 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_129
timestamp 1701704242
transform 1 0 76504 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_130
timestamp 1701704242
transform 1 0 73999 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_131
timestamp 1701704242
transform 1 0 74109 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_132
timestamp 1701704242
transform 1 0 73994 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_133
timestamp 1701704242
transform 1 0 73988 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_134
timestamp 1701704242
transform 1 0 74008 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_135
timestamp 1701704242
transform 1 0 71503 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_136
timestamp 1701704242
transform 1 0 71613 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_137
timestamp 1701704242
transform 1 0 71498 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_138
timestamp 1701704242
transform 1 0 71492 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_139
timestamp 1701704242
transform 1 0 71512 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_140
timestamp 1701704242
transform 1 0 69007 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_141
timestamp 1701704242
transform 1 0 69117 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_142
timestamp 1701704242
transform 1 0 69002 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_143
timestamp 1701704242
transform 1 0 68996 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_144
timestamp 1701704242
transform 1 0 69016 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_145
timestamp 1701704242
transform 1 0 66511 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_146
timestamp 1701704242
transform 1 0 66621 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_147
timestamp 1701704242
transform 1 0 66506 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_148
timestamp 1701704242
transform 1 0 66500 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_149
timestamp 1701704242
transform 1 0 66520 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_150
timestamp 1701704242
transform 1 0 64015 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_151
timestamp 1701704242
transform 1 0 64125 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_152
timestamp 1701704242
transform 1 0 64010 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_153
timestamp 1701704242
transform 1 0 64004 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_154
timestamp 1701704242
transform 1 0 64024 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_155
timestamp 1701704242
transform 1 0 61519 0 1 1546
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_156
timestamp 1701704242
transform 1 0 61629 0 1 778
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_157
timestamp 1701704242
transform 1 0 61514 0 1 575
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_158
timestamp 1701704242
transform 1 0 61508 0 1 1109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_21  sky130_sram_2kbyte_1rw1r_32x512_8_contact_21_159
timestamp 1701704242
transform 1 0 61528 0 1 159
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_0
timestamp 1701704242
transform 1 0 14083 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_1
timestamp 1701704242
transform 1 0 14077 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_2
timestamp 1701704242
transform 1 0 14097 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_3
timestamp 1701704242
transform 1 0 11592 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_4
timestamp 1701704242
transform 1 0 11702 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_5
timestamp 1701704242
transform 1 0 11587 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_6
timestamp 1701704242
transform 1 0 11581 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_7
timestamp 1701704242
transform 1 0 11601 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_8
timestamp 1701704242
transform 1 0 9096 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_9
timestamp 1701704242
transform 1 0 9206 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_10
timestamp 1701704242
transform 1 0 9091 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_11
timestamp 1701704242
transform 1 0 9085 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_12
timestamp 1701704242
transform 1 0 9105 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_13
timestamp 1701704242
transform 1 0 6600 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_14
timestamp 1701704242
transform 1 0 6710 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_15
timestamp 1701704242
transform 1 0 6595 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_16
timestamp 1701704242
transform 1 0 6589 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_17
timestamp 1701704242
transform 1 0 6609 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_18
timestamp 1701704242
transform 1 0 4104 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_19
timestamp 1701704242
transform 1 0 4214 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_20
timestamp 1701704242
transform 1 0 4099 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_21
timestamp 1701704242
transform 1 0 4093 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_22
timestamp 1701704242
transform 1 0 4113 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_23
timestamp 1701704242
transform 1 0 1608 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_24
timestamp 1701704242
transform 1 0 1718 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_25
timestamp 1701704242
transform 1 0 1603 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_26
timestamp 1701704242
transform 1 0 1597 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_27
timestamp 1701704242
transform 1 0 1617 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_28
timestamp 1701704242
transform 1 0 19080 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_29
timestamp 1701704242
transform 1 0 19190 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_30
timestamp 1701704242
transform 1 0 19075 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_31
timestamp 1701704242
transform 1 0 19069 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_32
timestamp 1701704242
transform 1 0 19089 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_33
timestamp 1701704242
transform 1 0 16584 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_34
timestamp 1701704242
transform 1 0 16694 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_35
timestamp 1701704242
transform 1 0 16579 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_36
timestamp 1701704242
transform 1 0 16573 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_37
timestamp 1701704242
transform 1 0 16593 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_38
timestamp 1701704242
transform 1 0 14088 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_39
timestamp 1701704242
transform 1 0 14198 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_40
timestamp 1701704242
transform 1 0 36541 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_41
timestamp 1701704242
transform 1 0 36561 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_42
timestamp 1701704242
transform 1 0 34056 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_43
timestamp 1701704242
transform 1 0 34166 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_44
timestamp 1701704242
transform 1 0 34051 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_45
timestamp 1701704242
transform 1 0 34045 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_46
timestamp 1701704242
transform 1 0 34065 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_47
timestamp 1701704242
transform 1 0 31560 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_48
timestamp 1701704242
transform 1 0 31670 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_49
timestamp 1701704242
transform 1 0 31555 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_50
timestamp 1701704242
transform 1 0 31549 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_51
timestamp 1701704242
transform 1 0 31569 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_52
timestamp 1701704242
transform 1 0 29064 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_53
timestamp 1701704242
transform 1 0 29174 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_54
timestamp 1701704242
transform 1 0 29059 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_55
timestamp 1701704242
transform 1 0 29053 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_56
timestamp 1701704242
transform 1 0 29073 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_57
timestamp 1701704242
transform 1 0 26568 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_58
timestamp 1701704242
transform 1 0 26678 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_59
timestamp 1701704242
transform 1 0 26563 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_60
timestamp 1701704242
transform 1 0 26557 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_61
timestamp 1701704242
transform 1 0 26577 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_62
timestamp 1701704242
transform 1 0 24072 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_63
timestamp 1701704242
transform 1 0 24182 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_64
timestamp 1701704242
transform 1 0 24067 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_65
timestamp 1701704242
transform 1 0 24061 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_66
timestamp 1701704242
transform 1 0 24081 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_67
timestamp 1701704242
transform 1 0 21576 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_68
timestamp 1701704242
transform 1 0 21686 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_69
timestamp 1701704242
transform 1 0 21571 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_70
timestamp 1701704242
transform 1 0 21565 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_71
timestamp 1701704242
transform 1 0 21585 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_72
timestamp 1701704242
transform 1 0 39048 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_73
timestamp 1701704242
transform 1 0 39158 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_74
timestamp 1701704242
transform 1 0 39043 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_75
timestamp 1701704242
transform 1 0 39037 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_76
timestamp 1701704242
transform 1 0 39057 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_77
timestamp 1701704242
transform 1 0 36552 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_78
timestamp 1701704242
transform 1 0 36662 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_79
timestamp 1701704242
transform 1 0 36547 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_80
timestamp 1701704242
transform 1 0 59025 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_81
timestamp 1701704242
transform 1 0 56520 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_82
timestamp 1701704242
transform 1 0 56630 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_83
timestamp 1701704242
transform 1 0 56515 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_84
timestamp 1701704242
transform 1 0 56509 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_85
timestamp 1701704242
transform 1 0 56529 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_86
timestamp 1701704242
transform 1 0 54024 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_87
timestamp 1701704242
transform 1 0 54134 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_88
timestamp 1701704242
transform 1 0 54019 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_89
timestamp 1701704242
transform 1 0 54013 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_90
timestamp 1701704242
transform 1 0 54033 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_91
timestamp 1701704242
transform 1 0 51528 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_92
timestamp 1701704242
transform 1 0 51638 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_93
timestamp 1701704242
transform 1 0 51523 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_94
timestamp 1701704242
transform 1 0 51517 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_95
timestamp 1701704242
transform 1 0 51537 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_96
timestamp 1701704242
transform 1 0 49032 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_97
timestamp 1701704242
transform 1 0 49142 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_98
timestamp 1701704242
transform 1 0 49027 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_99
timestamp 1701704242
transform 1 0 49021 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_100
timestamp 1701704242
transform 1 0 49041 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_101
timestamp 1701704242
transform 1 0 46536 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_102
timestamp 1701704242
transform 1 0 46646 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_103
timestamp 1701704242
transform 1 0 46531 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_104
timestamp 1701704242
transform 1 0 46525 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_105
timestamp 1701704242
transform 1 0 46545 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_106
timestamp 1701704242
transform 1 0 44040 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_107
timestamp 1701704242
transform 1 0 44150 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_108
timestamp 1701704242
transform 1 0 44035 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_109
timestamp 1701704242
transform 1 0 44029 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_110
timestamp 1701704242
transform 1 0 44049 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_111
timestamp 1701704242
transform 1 0 41544 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_112
timestamp 1701704242
transform 1 0 41654 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_113
timestamp 1701704242
transform 1 0 41539 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_114
timestamp 1701704242
transform 1 0 41533 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_115
timestamp 1701704242
transform 1 0 41553 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_116
timestamp 1701704242
transform 1 0 59016 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_117
timestamp 1701704242
transform 1 0 59126 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_118
timestamp 1701704242
transform 1 0 59011 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_119
timestamp 1701704242
transform 1 0 59005 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_120
timestamp 1701704242
transform 1 0 78984 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_121
timestamp 1701704242
transform 1 0 79094 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_122
timestamp 1701704242
transform 1 0 78979 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_123
timestamp 1701704242
transform 1 0 78973 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_124
timestamp 1701704242
transform 1 0 78993 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_125
timestamp 1701704242
transform 1 0 76488 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_126
timestamp 1701704242
transform 1 0 76598 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_127
timestamp 1701704242
transform 1 0 76483 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_128
timestamp 1701704242
transform 1 0 76477 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_129
timestamp 1701704242
transform 1 0 76497 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_130
timestamp 1701704242
transform 1 0 73992 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_131
timestamp 1701704242
transform 1 0 74102 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_132
timestamp 1701704242
transform 1 0 73987 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_133
timestamp 1701704242
transform 1 0 73981 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_134
timestamp 1701704242
transform 1 0 74001 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_135
timestamp 1701704242
transform 1 0 71496 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_136
timestamp 1701704242
transform 1 0 71606 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_137
timestamp 1701704242
transform 1 0 71491 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_138
timestamp 1701704242
transform 1 0 71485 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_139
timestamp 1701704242
transform 1 0 71505 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_140
timestamp 1701704242
transform 1 0 69000 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_141
timestamp 1701704242
transform 1 0 69110 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_142
timestamp 1701704242
transform 1 0 68995 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_143
timestamp 1701704242
transform 1 0 68989 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_144
timestamp 1701704242
transform 1 0 69009 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_145
timestamp 1701704242
transform 1 0 66504 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_146
timestamp 1701704242
transform 1 0 66614 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_147
timestamp 1701704242
transform 1 0 66499 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_148
timestamp 1701704242
transform 1 0 66493 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_149
timestamp 1701704242
transform 1 0 66513 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_150
timestamp 1701704242
transform 1 0 64008 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_151
timestamp 1701704242
transform 1 0 64118 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_152
timestamp 1701704242
transform 1 0 64003 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_153
timestamp 1701704242
transform 1 0 63997 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_154
timestamp 1701704242
transform 1 0 64017 0 1 154
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_155
timestamp 1701704242
transform 1 0 61512 0 1 1541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_156
timestamp 1701704242
transform 1 0 61622 0 1 772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_157
timestamp 1701704242
transform 1 0 61507 0 1 570
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_158
timestamp 1701704242
transform 1 0 61501 0 1 1104
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_22  sky130_sram_2kbyte_1rw1r_32x512_8_contact_22_159
timestamp 1701704242
transform 1 0 61521 0 1 154
box 0 0 1 1
<< labels >>
rlabel metal3 s 46509 1092 46607 1190 4 vdd
port 1 nsew
rlabel metal3 s 49005 1092 49103 1190 4 vdd
port 1 nsew
rlabel metal3 s 71469 1092 71567 1190 4 vdd
port 1 nsew
rlabel metal3 s 68973 1092 69071 1190 4 vdd
port 1 nsew
rlabel metal3 s 53997 1092 54095 1190 4 vdd
port 1 nsew
rlabel metal3 s 66477 1092 66575 1190 4 vdd
port 1 nsew
rlabel metal3 s 51501 1092 51599 1190 4 vdd
port 1 nsew
rlabel metal3 s 73965 1092 74063 1190 4 vdd
port 1 nsew
rlabel metal3 s 41517 1092 41615 1190 4 vdd
port 1 nsew
rlabel metal3 s 58989 1092 59087 1190 4 vdd
port 1 nsew
rlabel metal3 s 61485 1092 61583 1190 4 vdd
port 1 nsew
rlabel metal3 s 78957 1092 79055 1190 4 vdd
port 1 nsew
rlabel metal3 s 44013 1092 44111 1190 4 vdd
port 1 nsew
rlabel metal3 s 56493 1092 56591 1190 4 vdd
port 1 nsew
rlabel metal3 s 63981 1092 64079 1190 4 vdd
port 1 nsew
rlabel metal3 s 76461 1092 76559 1190 4 vdd
port 1 nsew
rlabel metal3 s 49126 760 49224 858 4 gnd
port 2 nsew
rlabel metal3 s 61606 760 61704 858 4 gnd
port 2 nsew
rlabel metal3 s 79078 760 79176 858 4 gnd
port 2 nsew
rlabel metal3 s 59000 1529 59098 1627 4 gnd
port 2 nsew
rlabel metal3 s 69094 760 69192 858 4 gnd
port 2 nsew
rlabel metal3 s 41523 558 41621 656 4 gnd
port 2 nsew
rlabel metal3 s 66483 558 66581 656 4 gnd
port 2 nsew
rlabel metal3 s 76582 760 76680 858 4 gnd
port 2 nsew
rlabel metal3 s 63987 558 64085 656 4 gnd
port 2 nsew
rlabel metal3 s 71590 760 71688 858 4 gnd
port 2 nsew
rlabel metal3 s 51622 760 51720 858 4 gnd
port 2 nsew
rlabel metal3 s 51512 1529 51610 1627 4 gnd
port 2 nsew
rlabel metal3 s 68979 558 69077 656 4 gnd
port 2 nsew
rlabel metal3 s 54008 1529 54106 1627 4 gnd
port 2 nsew
rlabel metal3 s 66598 760 66696 858 4 gnd
port 2 nsew
rlabel metal3 s 76472 1529 76570 1627 4 gnd
port 2 nsew
rlabel metal3 s 56504 1529 56602 1627 4 gnd
port 2 nsew
rlabel metal3 s 41528 1529 41626 1627 4 gnd
port 2 nsew
rlabel metal3 s 54118 760 54216 858 4 gnd
port 2 nsew
rlabel metal3 s 73976 1529 74074 1627 4 gnd
port 2 nsew
rlabel metal3 s 49011 558 49109 656 4 gnd
port 2 nsew
rlabel metal3 s 59110 760 59208 858 4 gnd
port 2 nsew
rlabel metal3 s 64102 760 64200 858 4 gnd
port 2 nsew
rlabel metal3 s 74086 760 74184 858 4 gnd
port 2 nsew
rlabel metal3 s 68984 1529 69082 1627 4 gnd
port 2 nsew
rlabel metal3 s 58995 558 59093 656 4 gnd
port 2 nsew
rlabel metal3 s 46515 558 46613 656 4 gnd
port 2 nsew
rlabel metal3 s 49016 1529 49114 1627 4 gnd
port 2 nsew
rlabel metal3 s 73971 558 74069 656 4 gnd
port 2 nsew
rlabel metal3 s 44019 558 44117 656 4 gnd
port 2 nsew
rlabel metal3 s 71480 1529 71578 1627 4 gnd
port 2 nsew
rlabel metal3 s 61496 1529 61594 1627 4 gnd
port 2 nsew
rlabel metal3 s 76467 558 76565 656 4 gnd
port 2 nsew
rlabel metal3 s 63992 1529 64090 1627 4 gnd
port 2 nsew
rlabel metal3 s 78968 1529 79066 1627 4 gnd
port 2 nsew
rlabel metal3 s 44134 760 44232 858 4 gnd
port 2 nsew
rlabel metal3 s 78963 558 79061 656 4 gnd
port 2 nsew
rlabel metal3 s 46630 760 46728 858 4 gnd
port 2 nsew
rlabel metal3 s 46520 1529 46618 1627 4 gnd
port 2 nsew
rlabel metal3 s 66488 1529 66586 1627 4 gnd
port 2 nsew
rlabel metal3 s 61491 558 61589 656 4 gnd
port 2 nsew
rlabel metal3 s 56614 760 56712 858 4 gnd
port 2 nsew
rlabel metal3 s 54003 558 54101 656 4 gnd
port 2 nsew
rlabel metal3 s 56499 558 56597 656 4 gnd
port 2 nsew
rlabel metal3 s 41638 760 41736 858 4 gnd
port 2 nsew
rlabel metal3 s 44024 1529 44122 1627 4 gnd
port 2 nsew
rlabel metal3 s 51507 558 51605 656 4 gnd
port 2 nsew
rlabel metal3 s 71475 558 71573 656 4 gnd
port 2 nsew
rlabel metal3 s 34040 1529 34138 1627 4 gnd
port 2 nsew
rlabel metal3 s 1581 1092 1679 1190 4 vdd
port 1 nsew
rlabel metal3 s 16557 1092 16655 1190 4 vdd
port 1 nsew
rlabel metal3 s 16563 558 16661 656 4 gnd
port 2 nsew
rlabel metal3 s 31654 760 31752 858 4 gnd
port 2 nsew
rlabel metal3 s 29158 760 29256 858 4 gnd
port 2 nsew
rlabel metal3 s 4088 1529 4186 1627 4 gnd
port 2 nsew
rlabel metal3 s 14182 760 14280 858 4 gnd
port 2 nsew
rlabel metal3 s 6579 558 6677 656 4 gnd
port 2 nsew
rlabel metal3 s 11565 1092 11663 1190 4 vdd
port 1 nsew
rlabel metal3 s 14061 1092 14159 1190 4 vdd
port 1 nsew
rlabel metal3 s 6573 1092 6671 1190 4 vdd
port 1 nsew
rlabel metal3 s 26552 1529 26650 1627 4 gnd
port 2 nsew
rlabel metal3 s 1592 1529 1690 1627 4 gnd
port 2 nsew
rlabel metal3 s 16568 1529 16666 1627 4 gnd
port 2 nsew
rlabel metal3 s 11576 1529 11674 1627 4 gnd
port 2 nsew
rlabel metal3 s 36531 558 36629 656 4 gnd
port 2 nsew
rlabel metal3 s 36525 1092 36623 1190 4 vdd
port 1 nsew
rlabel metal3 s 9080 1529 9178 1627 4 gnd
port 2 nsew
rlabel metal3 s 16678 760 16776 858 4 gnd
port 2 nsew
rlabel metal3 s 39027 558 39125 656 4 gnd
port 2 nsew
rlabel metal3 s 24166 760 24264 858 4 gnd
port 2 nsew
rlabel metal3 s 21670 760 21768 858 4 gnd
port 2 nsew
rlabel metal3 s 29037 1092 29135 1190 4 vdd
port 1 nsew
rlabel metal3 s 4077 1092 4175 1190 4 vdd
port 1 nsew
rlabel metal3 s 9075 558 9173 656 4 gnd
port 2 nsew
rlabel metal3 s 24045 1092 24143 1190 4 vdd
port 1 nsew
rlabel metal3 s 14072 1529 14170 1627 4 gnd
port 2 nsew
rlabel metal3 s 4198 760 4296 858 4 gnd
port 2 nsew
rlabel metal3 s 39021 1092 39119 1190 4 vdd
port 1 nsew
rlabel metal3 s 21560 1529 21658 1627 4 gnd
port 2 nsew
rlabel metal3 s 31544 1529 31642 1627 4 gnd
port 2 nsew
rlabel metal3 s 19053 1092 19151 1190 4 vdd
port 1 nsew
rlabel metal3 s 39142 760 39240 858 4 gnd
port 2 nsew
rlabel metal3 s 21549 1092 21647 1190 4 vdd
port 1 nsew
rlabel metal3 s 34035 558 34133 656 4 gnd
port 2 nsew
rlabel metal3 s 11571 558 11669 656 4 gnd
port 2 nsew
rlabel metal3 s 31539 558 31637 656 4 gnd
port 2 nsew
rlabel metal3 s 31533 1092 31631 1190 4 vdd
port 1 nsew
rlabel metal3 s 26541 1092 26639 1190 4 vdd
port 1 nsew
rlabel metal3 s 24051 558 24149 656 4 gnd
port 2 nsew
rlabel metal3 s 36646 760 36744 858 4 gnd
port 2 nsew
rlabel metal3 s 11686 760 11784 858 4 gnd
port 2 nsew
rlabel metal3 s 4083 558 4181 656 4 gnd
port 2 nsew
rlabel metal3 s 19174 760 19272 858 4 gnd
port 2 nsew
rlabel metal3 s 9069 1092 9167 1190 4 vdd
port 1 nsew
rlabel metal3 s 9190 760 9288 858 4 gnd
port 2 nsew
rlabel metal3 s 21555 558 21653 656 4 gnd
port 2 nsew
rlabel metal3 s 6694 760 6792 858 4 gnd
port 2 nsew
rlabel metal3 s 19059 558 19157 656 4 gnd
port 2 nsew
rlabel metal3 s 6584 1529 6682 1627 4 gnd
port 2 nsew
rlabel metal3 s 1587 558 1685 656 4 gnd
port 2 nsew
rlabel metal3 s 26662 760 26760 858 4 gnd
port 2 nsew
rlabel metal3 s 14067 558 14165 656 4 gnd
port 2 nsew
rlabel metal3 s 1702 760 1800 858 4 gnd
port 2 nsew
rlabel metal3 s 36536 1529 36634 1627 4 gnd
port 2 nsew
rlabel metal3 s 29048 1529 29146 1627 4 gnd
port 2 nsew
rlabel metal3 s 34150 760 34248 858 4 gnd
port 2 nsew
rlabel metal3 s 24056 1529 24154 1627 4 gnd
port 2 nsew
rlabel metal3 s 29043 558 29141 656 4 gnd
port 2 nsew
rlabel metal3 s 34029 1092 34127 1190 4 vdd
port 1 nsew
rlabel metal3 s 26547 558 26645 656 4 gnd
port 2 nsew
rlabel metal3 s 39032 1529 39130 1627 4 gnd
port 2 nsew
rlabel metal3 s 19064 1529 19162 1627 4 gnd
port 2 nsew
rlabel metal3 s 34049 142 34147 240 4 vdd
port 1 nsew
rlabel metal3 s 16577 142 16675 240 4 vdd
port 1 nsew
rlabel metal3 s 14081 142 14179 240 4 vdd
port 1 nsew
rlabel metal3 s 1601 142 1699 240 4 vdd
port 1 nsew
rlabel metal3 s 39041 142 39139 240 4 vdd
port 1 nsew
rlabel metal3 s 21569 142 21667 240 4 vdd
port 1 nsew
rlabel metal3 s 36545 142 36643 240 4 vdd
port 1 nsew
rlabel metal3 s 26561 142 26659 240 4 vdd
port 1 nsew
rlabel metal3 s 9089 142 9187 240 4 vdd
port 1 nsew
rlabel metal3 s 19073 142 19171 240 4 vdd
port 1 nsew
rlabel metal3 s 31553 142 31651 240 4 vdd
port 1 nsew
rlabel metal3 s 29057 142 29155 240 4 vdd
port 1 nsew
rlabel metal3 s 11585 142 11683 240 4 vdd
port 1 nsew
rlabel metal3 s 4097 142 4195 240 4 vdd
port 1 nsew
rlabel metal3 s 24065 142 24163 240 4 vdd
port 1 nsew
rlabel metal3 s 6593 142 6691 240 4 vdd
port 1 nsew
rlabel metal3 s 46529 142 46627 240 4 vdd
port 1 nsew
rlabel metal3 s 71489 142 71587 240 4 vdd
port 1 nsew
rlabel metal3 s 41537 142 41635 240 4 vdd
port 1 nsew
rlabel metal3 s 76481 142 76579 240 4 vdd
port 1 nsew
rlabel metal3 s 68993 142 69091 240 4 vdd
port 1 nsew
rlabel metal3 s 73985 142 74083 240 4 vdd
port 1 nsew
rlabel metal3 s 61505 142 61603 240 4 vdd
port 1 nsew
rlabel metal3 s 56513 142 56611 240 4 vdd
port 1 nsew
rlabel metal3 s 66497 142 66595 240 4 vdd
port 1 nsew
rlabel metal3 s 51521 142 51619 240 4 vdd
port 1 nsew
rlabel metal3 s 64001 142 64099 240 4 vdd
port 1 nsew
rlabel metal3 s 49025 142 49123 240 4 vdd
port 1 nsew
rlabel metal3 s 78977 142 79075 240 4 vdd
port 1 nsew
rlabel metal3 s 44033 142 44131 240 4 vdd
port 1 nsew
rlabel metal3 s 54017 142 54115 240 4 vdd
port 1 nsew
rlabel metal3 s 59009 142 59107 240 4 vdd
port 1 nsew
rlabel metal1 s 1629 4 1689 60 4 data_0
port 3 nsew
rlabel metal1 s 1500 1959 1530 2011 4 bl_0
port 4 nsew
rlabel metal1 s 1702 1959 1732 2011 4 br_0
port 5 nsew
rlabel metal1 s 4125 4 4185 60 4 data_1
port 6 nsew
rlabel metal1 s 3996 1959 4026 2011 4 bl_1
port 7 nsew
rlabel metal1 s 4198 1959 4228 2011 4 br_1
port 8 nsew
rlabel metal1 s 6621 4 6681 60 4 data_2
port 9 nsew
rlabel metal1 s 6492 1959 6522 2011 4 bl_2
port 10 nsew
rlabel metal1 s 6694 1959 6724 2011 4 br_2
port 11 nsew
rlabel metal1 s 9117 4 9177 60 4 data_3
port 12 nsew
rlabel metal1 s 8988 1959 9018 2011 4 bl_3
port 13 nsew
rlabel metal1 s 9190 1959 9220 2011 4 br_3
port 14 nsew
rlabel metal1 s 11613 4 11673 60 4 data_4
port 15 nsew
rlabel metal1 s 11484 1959 11514 2011 4 bl_4
port 16 nsew
rlabel metal1 s 11686 1959 11716 2011 4 br_4
port 17 nsew
rlabel metal1 s 14109 4 14169 60 4 data_5
port 18 nsew
rlabel metal1 s 13980 1959 14010 2011 4 bl_5
port 19 nsew
rlabel metal1 s 14182 1959 14212 2011 4 br_5
port 20 nsew
rlabel metal1 s 16605 4 16665 60 4 data_6
port 21 nsew
rlabel metal1 s 16476 1959 16506 2011 4 bl_6
port 22 nsew
rlabel metal1 s 16678 1959 16708 2011 4 br_6
port 23 nsew
rlabel metal1 s 19101 4 19161 60 4 data_7
port 24 nsew
rlabel metal1 s 18972 1959 19002 2011 4 bl_7
port 25 nsew
rlabel metal1 s 19174 1959 19204 2011 4 br_7
port 26 nsew
rlabel metal1 s 21597 4 21657 60 4 data_8
port 27 nsew
rlabel metal1 s 21468 1959 21498 2011 4 bl_8
port 28 nsew
rlabel metal1 s 21670 1959 21700 2011 4 br_8
port 29 nsew
rlabel metal1 s 24093 4 24153 60 4 data_9
port 30 nsew
rlabel metal1 s 23964 1959 23994 2011 4 bl_9
port 31 nsew
rlabel metal1 s 24166 1959 24196 2011 4 br_9
port 32 nsew
rlabel metal1 s 26589 4 26649 60 4 data_10
port 33 nsew
rlabel metal1 s 26460 1959 26490 2011 4 bl_10
port 34 nsew
rlabel metal1 s 26662 1959 26692 2011 4 br_10
port 35 nsew
rlabel metal1 s 29085 4 29145 60 4 data_11
port 36 nsew
rlabel metal1 s 28956 1959 28986 2011 4 bl_11
port 37 nsew
rlabel metal1 s 29158 1959 29188 2011 4 br_11
port 38 nsew
rlabel metal1 s 31581 4 31641 60 4 data_12
port 39 nsew
rlabel metal1 s 31452 1959 31482 2011 4 bl_12
port 40 nsew
rlabel metal1 s 31654 1959 31684 2011 4 br_12
port 41 nsew
rlabel metal1 s 34077 4 34137 60 4 data_13
port 42 nsew
rlabel metal1 s 33948 1959 33978 2011 4 bl_13
port 43 nsew
rlabel metal1 s 34150 1959 34180 2011 4 br_13
port 44 nsew
rlabel metal1 s 36573 4 36633 60 4 data_14
port 45 nsew
rlabel metal1 s 36444 1959 36474 2011 4 bl_14
port 46 nsew
rlabel metal1 s 36646 1959 36676 2011 4 br_14
port 47 nsew
rlabel metal1 s 39069 4 39129 60 4 data_15
port 48 nsew
rlabel metal1 s 38940 1959 38970 2011 4 bl_15
port 49 nsew
rlabel metal1 s 39142 1959 39172 2011 4 br_15
port 50 nsew
rlabel metal1 s 41565 4 41625 60 4 data_16
port 51 nsew
rlabel metal1 s 41436 1959 41466 2011 4 bl_16
port 52 nsew
rlabel metal1 s 41638 1959 41668 2011 4 br_16
port 53 nsew
rlabel metal1 s 44061 4 44121 60 4 data_17
port 54 nsew
rlabel metal1 s 43932 1959 43962 2011 4 bl_17
port 55 nsew
rlabel metal1 s 44134 1959 44164 2011 4 br_17
port 56 nsew
rlabel metal1 s 46557 4 46617 60 4 data_18
port 57 nsew
rlabel metal1 s 46428 1959 46458 2011 4 bl_18
port 58 nsew
rlabel metal1 s 46630 1959 46660 2011 4 br_18
port 59 nsew
rlabel metal1 s 49053 4 49113 60 4 data_19
port 60 nsew
rlabel metal1 s 48924 1959 48954 2011 4 bl_19
port 61 nsew
rlabel metal1 s 49126 1959 49156 2011 4 br_19
port 62 nsew
rlabel metal1 s 51549 4 51609 60 4 data_20
port 63 nsew
rlabel metal1 s 51420 1959 51450 2011 4 bl_20
port 64 nsew
rlabel metal1 s 51622 1959 51652 2011 4 br_20
port 65 nsew
rlabel metal1 s 54045 4 54105 60 4 data_21
port 66 nsew
rlabel metal1 s 53916 1959 53946 2011 4 bl_21
port 67 nsew
rlabel metal1 s 54118 1959 54148 2011 4 br_21
port 68 nsew
rlabel metal1 s 56541 4 56601 60 4 data_22
port 69 nsew
rlabel metal1 s 56412 1959 56442 2011 4 bl_22
port 70 nsew
rlabel metal1 s 56614 1959 56644 2011 4 br_22
port 71 nsew
rlabel metal1 s 59037 4 59097 60 4 data_23
port 72 nsew
rlabel metal1 s 58908 1959 58938 2011 4 bl_23
port 73 nsew
rlabel metal1 s 59110 1959 59140 2011 4 br_23
port 74 nsew
rlabel metal1 s 61533 4 61593 60 4 data_24
port 75 nsew
rlabel metal1 s 61404 1959 61434 2011 4 bl_24
port 76 nsew
rlabel metal1 s 61606 1959 61636 2011 4 br_24
port 77 nsew
rlabel metal1 s 64029 4 64089 60 4 data_25
port 78 nsew
rlabel metal1 s 63900 1959 63930 2011 4 bl_25
port 79 nsew
rlabel metal1 s 64102 1959 64132 2011 4 br_25
port 80 nsew
rlabel metal1 s 66525 4 66585 60 4 data_26
port 81 nsew
rlabel metal1 s 66396 1959 66426 2011 4 bl_26
port 82 nsew
rlabel metal1 s 66598 1959 66628 2011 4 br_26
port 83 nsew
rlabel metal1 s 69021 4 69081 60 4 data_27
port 84 nsew
rlabel metal1 s 68892 1959 68922 2011 4 bl_27
port 85 nsew
rlabel metal1 s 69094 1959 69124 2011 4 br_27
port 86 nsew
rlabel metal1 s 71517 4 71577 60 4 data_28
port 87 nsew
rlabel metal1 s 71388 1959 71418 2011 4 bl_28
port 88 nsew
rlabel metal1 s 71590 1959 71620 2011 4 br_28
port 89 nsew
rlabel metal1 s 74013 4 74073 60 4 data_29
port 90 nsew
rlabel metal1 s 73884 1959 73914 2011 4 bl_29
port 91 nsew
rlabel metal1 s 74086 1959 74116 2011 4 br_29
port 92 nsew
rlabel metal1 s 76509 4 76569 60 4 data_30
port 93 nsew
rlabel metal1 s 76380 1959 76410 2011 4 bl_30
port 94 nsew
rlabel metal1 s 76582 1959 76612 2011 4 br_30
port 95 nsew
rlabel metal1 s 79005 4 79065 60 4 data_31
port 96 nsew
rlabel metal1 s 78876 1959 78906 2011 4 bl_31
port 97 nsew
rlabel metal1 s 79078 1959 79108 2011 4 br_31
port 98 nsew
rlabel metal1 s 1473 94 20817 128 4 en_0
port 99 nsew
rlabel metal1 s 21441 94 40785 128 4 en_1
port 100 nsew
rlabel metal1 s 41409 94 60753 128 4 en_2
port 101 nsew
rlabel metal1 s 61377 94 80721 128 4 en_3
port 102 nsew
<< properties >>
string FIXED_BBOX 0 0 79250 2011
string GDS_END 1446436
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 1364708
<< end >>
