magic
tech sky130B
timestamp 1701704242
<< pwell >>
rect -13 -13 38 688
<< ndiff >>
rect 0 669 25 675
rect 0 652 4 669
rect 21 652 25 669
rect 0 635 25 652
rect 0 618 4 635
rect 21 618 25 635
rect 0 601 25 618
rect 0 584 4 601
rect 21 584 25 601
rect 0 567 25 584
rect 0 550 4 567
rect 21 550 25 567
rect 0 533 25 550
rect 0 516 4 533
rect 21 516 25 533
rect 0 499 25 516
rect 0 482 4 499
rect 21 482 25 499
rect 0 465 25 482
rect 0 448 4 465
rect 21 448 25 465
rect 0 431 25 448
rect 0 414 4 431
rect 21 414 25 431
rect 0 397 25 414
rect 0 380 4 397
rect 21 380 25 397
rect 0 363 25 380
rect 0 346 4 363
rect 21 346 25 363
rect 0 329 25 346
rect 0 312 4 329
rect 21 312 25 329
rect 0 295 25 312
rect 0 278 4 295
rect 21 278 25 295
rect 0 261 25 278
rect 0 244 4 261
rect 21 244 25 261
rect 0 227 25 244
rect 0 210 4 227
rect 21 210 25 227
rect 0 193 25 210
rect 0 176 4 193
rect 21 176 25 193
rect 0 159 25 176
rect 0 142 4 159
rect 21 142 25 159
rect 0 125 25 142
rect 0 108 4 125
rect 21 108 25 125
rect 0 91 25 108
rect 0 74 4 91
rect 21 74 25 91
rect 0 57 25 74
rect 0 40 4 57
rect 21 40 25 57
rect 0 23 25 40
rect 0 6 4 23
rect 21 6 25 23
rect 0 0 25 6
<< ndiffc >>
rect 4 652 21 669
rect 4 618 21 635
rect 4 584 21 601
rect 4 550 21 567
rect 4 516 21 533
rect 4 482 21 499
rect 4 448 21 465
rect 4 414 21 431
rect 4 380 21 397
rect 4 346 21 363
rect 4 312 21 329
rect 4 278 21 295
rect 4 244 21 261
rect 4 210 21 227
rect 4 176 21 193
rect 4 142 21 159
rect 4 108 21 125
rect 4 74 21 91
rect 4 40 21 57
rect 4 6 21 23
<< locali >>
rect 4 669 21 677
rect 4 635 21 652
rect 4 601 21 618
rect 4 567 21 584
rect 4 533 21 550
rect 4 499 21 516
rect 4 465 21 482
rect 4 431 21 448
rect 4 397 21 414
rect 4 363 21 380
rect 4 329 21 346
rect 4 295 21 312
rect 4 261 21 278
rect 4 227 21 244
rect 4 193 21 210
rect 4 159 21 176
rect 4 125 21 142
rect 4 91 21 108
rect 4 57 21 74
rect 4 23 21 40
rect 4 -2 21 6
<< properties >>
string GDS_END 2730086
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2728610
<< end >>
