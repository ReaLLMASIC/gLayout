magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -154 -66 222 366
<< mvpmos >>
rect 0 0 100 300
<< mvpdiff >>
rect -88 250 0 300
rect -88 216 -77 250
rect -43 216 0 250
rect -88 182 0 216
rect -88 148 -77 182
rect -43 148 0 182
rect -88 114 0 148
rect -88 80 -77 114
rect -43 80 0 114
rect -88 46 0 80
rect -88 12 -77 46
rect -43 12 0 46
rect -88 0 0 12
rect 100 250 156 300
rect 100 216 111 250
rect 145 216 156 250
rect 100 182 156 216
rect 100 148 111 182
rect 145 148 156 182
rect 100 114 156 148
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
<< mvpdiffc >>
rect -77 216 -43 250
rect -77 148 -43 182
rect -77 80 -43 114
rect -77 12 -43 46
rect 111 216 145 250
rect 111 148 145 182
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 300 100 326
rect 0 -26 100 0
<< locali >>
rect -77 250 -43 266
rect -77 182 -43 216
rect -77 114 -43 148
rect -77 46 -43 80
rect -77 -4 -43 12
rect 111 250 145 266
rect 111 182 145 216
rect 111 114 145 148
rect 111 46 145 80
rect 111 -4 145 12
use DFL1sd2_CDNS_52468879185253  DFL1sd2_CDNS_52468879185253_0
timestamp 1701704242
transform -1 0 -32 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_52468879185253  DFL1sd2_CDNS_52468879185253_1
timestamp 1701704242
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -60 131 -60 131 0 FreeSans 300 0 0 0 S
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 70892850
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70891768
<< end >>
