magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 53 161
<< metal1 >>
rect -6 161 59 164
rect -6 0 0 161
rect 53 0 59 161
rect -6 -3 59 0
<< properties >>
string GDS_END 97530284
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97529512
<< end >>
