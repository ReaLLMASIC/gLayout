magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1027 203
rect 30 -17 64 21
<< locali >>
rect 28 215 248 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 323 85 493
rect 119 367 153 527
rect 187 323 253 493
rect 287 367 321 527
rect 371 323 405 493
rect 439 367 505 527
rect 539 323 573 493
rect 607 367 673 527
rect 707 323 741 493
rect 775 367 841 527
rect 875 323 909 493
rect 19 289 319 323
rect 371 289 909 323
rect 943 297 1009 527
rect 284 249 319 289
rect 858 263 909 289
rect 284 215 809 249
rect 284 181 319 215
rect 858 211 977 263
rect 858 181 909 211
rect 35 147 319 181
rect 371 147 909 181
rect 35 51 69 147
rect 103 17 169 113
rect 203 52 237 147
rect 271 17 337 113
rect 371 51 405 147
rect 439 17 505 113
rect 539 51 573 147
rect 607 17 673 113
rect 707 51 741 147
rect 775 17 841 113
rect 875 51 909 147
rect 943 17 1009 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< obsm1 >>
rect 693 261 821 264
rect 693 215 982 261
rect 693 212 821 215
<< obsm2 >>
rect 689 201 825 275
<< metal3 >>
rect 679 270 835 271
rect 679 206 685 270
rect 749 206 765 270
rect 829 206 835 270
rect 679 205 835 206
<< via3 >>
rect 685 206 749 270
rect 765 206 829 270
<< metal4 >>
rect 274 136 594 372
<< via4 >>
rect 594 270 830 372
rect 594 206 685 270
rect 685 206 749 270
rect 749 206 765 270
rect 765 206 829 270
rect 829 206 830 270
rect 594 136 830 206
<< metal5 >>
rect 250 390 854 432
rect 250 372 854 389
rect 250 136 594 372
rect 830 136 854 372
rect 250 112 854 136
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 1027 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal5 s 250 390 854 432 6 X
port 6 nsew signal output
rlabel metal5 s 250 112 854 389 6 X
port 6 nsew signal output
rlabel via4 s 594 136 830 372 6 X
port 6 nsew signal output
rlabel metal4 s 274 136 830 372 6 X
port 6 nsew signal output
rlabel via3 s 765 206 829 270 6 X
port 6 nsew signal output
rlabel via3 s 685 206 749 270 6 X
port 6 nsew signal output
rlabel metal3 s 679 205 835 271 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 18906
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 8946
<< end >>
