magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -36 -36 161 636
<< pdiff >>
rect 0 522 60 600
rect 0 488 11 522
rect 45 488 60 522
rect 0 454 60 488
rect 0 420 11 454
rect 45 420 60 454
rect 0 386 60 420
rect 0 352 11 386
rect 45 352 60 386
rect 0 318 60 352
rect 0 284 11 318
rect 45 284 60 318
rect 0 250 60 284
rect 0 216 11 250
rect 45 216 60 250
rect 0 182 60 216
rect 0 148 11 182
rect 45 148 60 182
rect 0 114 60 148
rect 0 80 11 114
rect 45 80 60 114
rect 0 46 60 80
rect 0 12 11 46
rect 45 12 60 46
rect 0 0 60 12
<< pdiffc >>
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< nsubdiff >>
rect 60 522 125 600
rect 60 488 79 522
rect 113 488 125 522
rect 60 454 125 488
rect 60 420 79 454
rect 113 420 125 454
rect 60 386 125 420
rect 60 352 79 386
rect 113 352 125 386
rect 60 318 125 352
rect 60 284 79 318
rect 113 284 125 318
rect 60 250 125 284
rect 60 216 79 250
rect 113 216 125 250
rect 60 182 125 216
rect 60 148 79 182
rect 113 148 125 182
rect 60 114 125 148
rect 60 80 79 114
rect 113 80 125 114
rect 60 46 125 80
rect 60 12 79 46
rect 113 12 125 46
rect 60 0 125 12
<< nsubdiffcont >>
rect 79 488 113 522
rect 79 420 113 454
rect 79 352 113 386
rect 79 284 113 318
rect 79 216 113 250
rect 79 148 113 182
rect 79 80 113 114
rect 79 12 113 46
<< locali >>
rect 11 534 113 538
rect 45 522 113 534
rect 45 488 79 522
rect 11 462 113 488
rect 45 454 113 462
rect 45 420 79 454
rect 11 390 113 420
rect 45 386 113 390
rect 45 352 79 386
rect 11 318 113 352
rect 45 284 79 318
rect 11 250 113 284
rect 45 216 79 250
rect 45 212 113 216
rect 11 182 113 212
rect 45 148 79 182
rect 45 140 113 148
rect 11 114 113 140
rect 45 80 79 114
rect 45 68 113 80
rect 11 46 113 68
rect 45 12 79 46
rect 45 -4 113 12
<< viali >>
rect 11 522 45 534
rect 11 500 45 522
rect 11 454 45 462
rect 11 428 45 454
rect 11 386 45 390
rect 11 356 45 386
rect 11 284 45 318
rect 11 216 45 246
rect 11 212 45 216
rect 11 148 45 174
rect 11 140 45 148
rect 11 80 45 102
rect 11 68 45 80
rect 11 12 45 30
rect 11 -4 45 12
<< metal1 >>
rect 5 534 51 546
rect 5 500 11 534
rect 45 500 51 534
rect 5 462 51 500
rect 5 428 11 462
rect 45 428 51 462
rect 5 390 51 428
rect 5 356 11 390
rect 45 356 51 390
rect 5 318 51 356
rect 5 284 11 318
rect 45 284 51 318
rect 5 246 51 284
rect 5 212 11 246
rect 45 212 51 246
rect 5 174 51 212
rect 5 140 11 174
rect 45 140 51 174
rect 5 102 51 140
rect 5 68 11 102
rect 45 68 51 102
rect 5 30 51 68
rect 5 -4 11 30
rect 45 -4 51 30
rect 5 -16 51 -4
<< properties >>
string GDS_END 86601078
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86599026
<< end >>
