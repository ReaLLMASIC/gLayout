magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 1123 3235 1676 3296
rect 832 3193 1676 3235
rect 802 3061 1676 3193
rect 832 3019 1676 3061
rect 1123 2564 1676 3019
<< mvnsubdiff >>
rect 838 3144 1121 3157
rect 838 3110 862 3144
rect 896 3110 930 3144
rect 964 3110 998 3144
rect 1032 3110 1121 3144
rect 838 3097 1121 3110
<< mvnsubdiffcont >>
rect 862 3110 896 3144
rect 930 3110 964 3144
rect 998 3110 1032 3144
<< poly >>
rect 403 3251 537 3267
rect 403 3217 419 3251
rect 453 3217 487 3251
rect 521 3217 537 3251
rect 403 3201 537 3217
rect 593 3037 727 3053
rect 593 3003 609 3037
rect 643 3003 677 3037
rect 711 3003 727 3037
rect 593 2987 727 3003
rect 1942 2582 2238 2598
rect 1942 2548 1958 2582
rect 1992 2548 2034 2582
rect 2068 2548 2111 2582
rect 2145 2548 2188 2582
rect 2222 2548 2238 2582
rect 1942 2532 2238 2548
rect 107 1118 403 1134
rect 107 1084 123 1118
rect 157 1084 200 1118
rect 234 1084 277 1118
rect 311 1084 353 1118
rect 387 1084 403 1118
rect 107 1068 403 1084
rect 459 1118 755 1134
rect 459 1084 475 1118
rect 509 1084 552 1118
rect 586 1084 629 1118
rect 663 1084 705 1118
rect 739 1084 755 1118
rect 459 1068 755 1084
rect 1930 718 2064 734
rect 1930 684 1946 718
rect 1980 684 2014 718
rect 2048 684 2064 718
rect 1930 668 2064 684
<< polycont >>
rect 419 3217 453 3251
rect 487 3217 521 3251
rect 609 3003 643 3037
rect 677 3003 711 3037
rect 1958 2548 1992 2582
rect 2034 2548 2068 2582
rect 2111 2548 2145 2582
rect 2188 2548 2222 2582
rect 123 1084 157 1118
rect 200 1084 234 1118
rect 277 1084 311 1118
rect 353 1084 387 1118
rect 475 1084 509 1118
rect 552 1084 586 1118
rect 629 1084 663 1118
rect 705 1084 739 1118
rect 1946 684 1980 718
rect 2014 684 2048 718
<< locali >>
rect 403 3257 793 3287
rect 403 3223 404 3257
rect 438 3251 476 3257
rect 510 3251 793 3257
rect 453 3223 476 3251
rect 403 3217 419 3223
rect 453 3217 487 3223
rect 521 3217 793 3251
rect 341 3130 432 3147
rect 341 3096 357 3130
rect 391 3096 432 3130
rect 341 3058 432 3096
rect 548 3108 582 3146
rect 686 3081 793 3217
rect 1776 3200 1820 3234
rect 1854 3200 1898 3234
rect 1742 3162 1932 3200
rect 838 3144 1121 3157
rect 896 3110 921 3144
rect 964 3110 998 3144
rect 1038 3110 1087 3144
rect 838 3097 1121 3110
rect 1776 3128 1820 3162
rect 1854 3128 1898 3162
rect 1742 3090 1932 3128
rect 341 3024 357 3058
rect 391 3037 432 3058
rect 1776 3056 1820 3090
rect 1854 3056 1898 3090
rect 391 3024 609 3037
rect 341 3003 609 3024
rect 643 3003 677 3037
rect 711 3003 727 3037
rect 1742 3018 1932 3056
rect 1776 2984 1820 3018
rect 1854 2984 1898 3018
rect 2249 3162 2283 3200
rect 2249 3090 2283 3128
rect 2249 3018 2283 3056
rect 2073 2726 2107 2764
rect 1935 2548 1958 2582
rect 2007 2548 2034 2582
rect 2068 2548 2111 2582
rect 2145 2548 2188 2582
rect 2222 2548 2238 2582
rect 107 1174 660 1208
rect 694 1174 732 1208
rect 107 1118 403 1174
rect 107 1084 123 1118
rect 157 1084 200 1118
rect 234 1084 277 1118
rect 311 1084 353 1118
rect 387 1084 403 1118
rect 459 1084 475 1118
rect 509 1084 552 1118
rect 586 1084 629 1118
rect 671 1084 705 1118
rect 743 1084 755 1118
rect 238 769 272 811
rect 238 693 272 735
rect 238 617 272 659
rect 238 541 272 583
rect 590 766 624 811
rect 590 687 624 732
rect 1586 718 1620 734
rect 1586 696 1946 718
rect 1620 684 1946 696
rect 1980 684 2014 718
rect 2048 684 2064 718
rect 590 607 624 653
rect 238 464 272 507
rect 2073 502 2107 540
rect 62 210 96 248
rect 62 138 96 176
rect 62 66 96 104
rect 414 210 448 248
rect 414 138 448 176
rect 414 66 448 104
rect 766 210 800 248
rect 766 138 800 176
rect 766 66 800 104
rect 1821 248 1897 282
rect 1787 210 1931 248
rect 1821 176 1897 210
rect 1787 138 1931 176
rect 1821 104 1897 138
rect 1787 66 1931 104
rect 1821 32 1897 66
<< viali >>
rect 404 3251 438 3257
rect 476 3251 510 3257
rect 404 3223 419 3251
rect 419 3223 438 3251
rect 476 3223 487 3251
rect 487 3223 510 3251
rect 357 3096 391 3130
rect 548 3146 582 3180
rect 548 3074 582 3108
rect 1742 3200 1776 3234
rect 1820 3200 1854 3234
rect 1898 3200 1932 3234
rect 838 3110 862 3144
rect 862 3110 872 3144
rect 921 3110 930 3144
rect 930 3110 955 3144
rect 1004 3110 1032 3144
rect 1032 3110 1038 3144
rect 1087 3110 1121 3144
rect 1742 3128 1776 3162
rect 1820 3128 1854 3162
rect 1898 3128 1932 3162
rect 357 3024 391 3058
rect 1742 3056 1776 3090
rect 1820 3056 1854 3090
rect 1898 3056 1932 3090
rect 1742 2984 1776 3018
rect 1820 2984 1854 3018
rect 1898 2984 1932 3018
rect 2249 3200 2283 3234
rect 2249 3128 2283 3162
rect 2249 3056 2283 3090
rect 2249 2984 2283 3018
rect 2073 2764 2107 2798
rect 2073 2692 2107 2726
rect 1901 2548 1935 2582
rect 1973 2548 1992 2582
rect 1992 2548 2007 2582
rect 660 1174 694 1208
rect 732 1174 766 1208
rect 637 1084 663 1118
rect 663 1084 671 1118
rect 709 1084 739 1118
rect 739 1084 743 1118
rect 238 811 272 845
rect 238 735 272 769
rect 238 659 272 693
rect 238 583 272 617
rect 590 811 624 845
rect 590 732 624 766
rect 590 653 624 687
rect 1586 734 1620 768
rect 1586 662 1620 696
rect 590 573 624 607
rect 238 507 272 541
rect 2073 540 2107 574
rect 2073 468 2107 502
rect 238 430 272 464
rect 62 248 96 282
rect 62 176 96 210
rect 62 104 96 138
rect 62 32 96 66
rect 414 248 448 282
rect 414 176 448 210
rect 414 104 448 138
rect 414 32 448 66
rect 766 248 800 282
rect 766 176 800 210
rect 766 104 800 138
rect 766 32 800 66
rect 1787 248 1821 282
rect 1897 248 1931 282
rect 1787 176 1821 210
rect 1897 176 1931 210
rect 1787 104 1821 138
rect 1897 104 1931 138
rect 1787 32 1821 66
rect 1897 32 1931 66
<< metal1 >>
rect 392 3257 522 3263
rect 392 3223 404 3257
rect 438 3223 476 3257
rect 510 3223 522 3257
tri 1184 3234 1196 3246 se
rect 1196 3234 2289 3246
rect 392 3217 522 3223
tri 1167 3217 1184 3234 se
rect 1184 3217 1742 3234
rect 351 3130 397 3144
rect 351 3096 357 3130
rect 391 3096 397 3130
rect 351 3058 397 3096
rect 351 3024 357 3058
rect 391 3024 397 3058
rect 351 1866 397 3024
rect 464 2172 510 3217
tri 1150 3200 1167 3217 se
rect 1167 3200 1742 3217
rect 1776 3200 1820 3234
rect 1854 3200 1898 3234
rect 1932 3200 2249 3234
rect 2283 3200 2289 3234
tri 1142 3192 1150 3200 se
rect 1150 3192 2289 3200
rect 542 3180 2289 3192
rect 542 3146 548 3180
rect 582 3162 2289 3180
rect 582 3146 1742 3162
rect 542 3144 1742 3146
rect 542 3110 838 3144
rect 872 3110 921 3144
rect 955 3110 1004 3144
rect 1038 3110 1087 3144
rect 1121 3128 1742 3144
rect 1776 3128 1820 3162
rect 1854 3128 1898 3162
rect 1932 3128 2249 3162
rect 2283 3128 2289 3162
rect 1121 3110 2289 3128
rect 542 3108 2289 3110
rect 542 3074 548 3108
rect 582 3090 2289 3108
rect 582 3074 1742 3090
rect 542 3062 1742 3074
tri 1106 3056 1112 3062 ne
rect 1112 3056 1742 3062
rect 1776 3056 1820 3090
rect 1854 3056 1898 3090
rect 1932 3056 2249 3090
rect 2283 3056 2289 3090
tri 1112 3018 1150 3056 ne
rect 1150 3018 2289 3056
tri 1150 2984 1184 3018 ne
rect 1184 2984 1742 3018
rect 1776 2984 1820 3018
rect 1854 2984 1898 3018
rect 1932 2984 2249 3018
rect 2283 2984 2289 3018
tri 1184 2972 1196 2984 ne
rect 1196 2972 2289 2984
rect 2067 2798 2113 2810
rect 2067 2764 2073 2798
rect 2107 2764 2113 2798
rect 2067 2726 2113 2764
rect 2067 2692 2073 2726
rect 2107 2692 2113 2726
tri 1658 2582 1664 2588 se
rect 1664 2582 2019 2588
tri 1624 2548 1658 2582 se
rect 1658 2548 1901 2582
rect 1935 2548 1973 2582
rect 2007 2548 2019 2582
tri 1598 2522 1624 2548 se
rect 1624 2542 2019 2548
rect 1624 2522 1664 2542
tri 1664 2522 1684 2542 nw
tri 1580 2504 1598 2522 se
rect 1598 2504 1646 2522
tri 1646 2504 1664 2522 nw
tri 510 2172 530 2192 sw
tri 464 2106 530 2172 ne
tri 530 2106 596 2172 sw
tri 530 2040 596 2106 ne
tri 596 2040 662 2106 sw
tri 596 1974 662 2040 ne
tri 662 1974 728 2040 sw
tri 662 1908 728 1974 ne
tri 728 1908 794 1974 sw
tri 728 1886 750 1908 ne
rect 750 1886 794 1908
tri 794 1886 816 1908 sw
tri 351 1846 371 1866 ne
rect 371 1846 397 1866
tri 397 1846 437 1886 sw
tri 750 1846 790 1886 ne
rect 790 1846 816 1886
tri 816 1846 856 1886 sw
tri 371 1820 397 1846 ne
rect 397 1820 437 1846
tri 397 1780 437 1820 ne
tri 437 1780 503 1846 sw
tri 790 1842 794 1846 ne
rect 794 1842 856 1846
tri 856 1842 860 1846 sw
tri 794 1780 856 1842 ne
rect 856 1780 860 1842
tri 860 1780 922 1842 sw
tri 437 1714 503 1780 ne
tri 503 1714 569 1780 sw
tri 856 1776 860 1780 ne
rect 860 1776 922 1780
tri 922 1776 926 1780 sw
tri 503 1694 523 1714 ne
tri 495 1208 523 1236 se
rect 523 1216 569 1714
tri 860 1710 926 1776 ne
tri 926 1710 992 1776 sw
tri 926 1644 992 1710 ne
tri 992 1644 1058 1710 sw
tri 992 1624 1012 1644 ne
rect 523 1208 561 1216
tri 561 1208 569 1216 nw
rect 648 1208 778 1214
tri 461 1174 495 1208 se
rect 495 1174 527 1208
tri 527 1174 561 1208 nw
rect 648 1174 660 1208
rect 694 1174 732 1208
rect 766 1174 778 1208
tri 457 1170 461 1174 se
rect 461 1170 523 1174
tri 523 1170 527 1174 nw
tri 405 1118 457 1170 se
rect 457 1118 471 1170
tri 471 1118 523 1170 nw
rect 648 1168 778 1174
rect 625 1118 755 1124
tri 391 1104 405 1118 se
rect 405 1104 457 1118
tri 457 1104 471 1118 nw
tri 371 1084 391 1104 se
rect 391 1084 437 1104
tri 437 1084 457 1104 nw
rect 625 1084 637 1118
rect 671 1084 709 1118
rect 743 1084 755 1118
tri 325 1038 371 1084 se
rect 371 1038 391 1084
tri 391 1038 437 1084 nw
rect 625 1078 755 1084
tri 259 972 325 1038 se
tri 325 972 391 1038 nw
tri 232 945 259 972 se
rect 259 945 298 972
tri 298 945 325 972 nw
rect 232 845 278 945
tri 278 925 298 945 nw
rect 232 811 238 845
rect 272 811 278 845
rect 232 769 278 811
rect 232 735 238 769
rect 272 735 278 769
rect 232 693 278 735
rect 232 659 238 693
rect 272 659 278 693
rect 232 617 278 659
rect 232 583 238 617
rect 272 583 278 617
rect 232 541 278 583
rect 584 845 630 857
rect 584 811 590 845
rect 624 811 630 845
rect 584 766 630 811
rect 584 732 590 766
rect 624 732 630 766
rect 584 724 630 732
rect 1012 724 1058 1644
rect 584 687 1058 724
rect 584 653 590 687
rect 624 678 1058 687
rect 1580 768 1626 2504
tri 1626 2484 1646 2504 nw
rect 1580 734 1586 768
rect 1620 734 1626 768
rect 1580 696 1626 734
rect 624 653 630 678
rect 584 607 630 653
rect 584 573 590 607
rect 624 573 630 607
rect 584 561 630 573
rect 1580 662 1586 696
rect 1620 662 1626 696
rect 232 507 238 541
rect 272 507 278 541
rect 232 464 278 507
tri 1551 468 1580 497 se
rect 1580 477 1626 662
rect 1580 468 1617 477
tri 1617 468 1626 477 nw
rect 2067 574 2113 2692
rect 2067 540 2073 574
rect 2107 540 2113 574
rect 2067 502 2113 540
rect 2067 468 2073 502
rect 2107 468 2113 502
rect 232 430 238 464
rect 272 430 278 464
tri 1514 431 1551 468 se
rect 1551 431 1580 468
tri 1580 431 1617 468 nw
rect 2067 456 2113 468
rect 232 419 278 430
tri 1502 419 1514 431 se
rect 1514 419 1568 431
tri 1568 419 1580 431 nw
rect 232 373 1522 419
tri 1522 373 1568 419 nw
rect 48 282 1937 294
rect 48 248 62 282
rect 96 248 414 282
rect 448 248 766 282
rect 800 248 1787 282
rect 1821 248 1897 282
rect 1931 248 1937 282
rect 48 210 1937 248
rect 48 176 62 210
rect 96 176 414 210
rect 448 176 766 210
rect 800 176 1787 210
rect 1821 176 1897 210
rect 1931 176 1937 210
rect 48 138 1937 176
rect 48 104 62 138
rect 96 104 414 138
rect 448 104 766 138
rect 800 104 1787 138
rect 1821 104 1897 138
rect 1931 104 1937 138
rect 48 66 1937 104
rect 48 32 62 66
rect 96 32 414 66
rect 448 32 766 66
rect 800 32 1787 66
rect 1821 32 1897 66
rect 1931 32 1937 66
rect 48 20 1937 32
use nfet_CDNS_52468879185919  nfet_CDNS_52468879185919_0
timestamp 1701704242
transform 1 0 459 0 1 36
box -79 -32 522 1032
use nfet_CDNS_52468879185921  nfet_CDNS_52468879185921_0
timestamp 1701704242
transform 1 0 107 0 1 36
box -79 -32 375 1032
use nfet_CDNS_52468879185922  nfet_CDNS_52468879185922_0
timestamp 1701704242
transform -1 0 2062 0 1 36
box -79 -32 346 632
use pfet_CDNS_52468879185918  pfet_CDNS_52468879185918_0
timestamp 1701704242
transform -1 0 537 0 1 3085
box -119 -66 239 150
use pfet_CDNS_52468879185918  pfet_CDNS_52468879185918_1
timestamp 1701704242
transform 1 0 593 0 1 3085
box -119 -66 239 150
use pfet_CDNS_52468879185920  pfet_CDNS_52468879185920_0
timestamp 1701704242
transform -1 0 2238 0 -1 3230
box -119 -66 562 666
<< labels >>
flabel metal1 s 1721 3077 1857 3198 0 FreeSans 200 0 0 0 vswitch
port 1 nsew
flabel metal1 s 695 123 766 209 0 FreeSans 200 0 0 0 vssa
port 2 nsew
flabel metal1 s 2072 628 2109 697 0 FreeSans 200 270 0 0 out_h
port 3 nsew
<< properties >>
string GDS_END 80519252
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80508348
string path 20.300 78.175 28.675 78.175 
<< end >>
