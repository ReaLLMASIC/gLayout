magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -77 435 645 797
<< pwell >>
rect -67 347 635 435
rect -55 93 623 347
<< nmos >>
rect 58 119 108 319
rect 176 119 226 319
rect 342 119 392 319
rect 460 119 510 319
<< pmoshvt >>
rect 58 561 108 761
rect 176 561 226 761
rect 342 561 392 761
rect 460 561 510 761
<< ndiff >>
rect -29 307 58 319
rect -29 273 -17 307
rect 17 273 58 307
rect -29 239 58 273
rect -29 205 -17 239
rect 17 205 58 239
rect -29 171 58 205
rect -29 137 -17 171
rect 17 137 58 171
rect -29 119 58 137
rect 108 307 176 319
rect 108 273 125 307
rect 159 273 176 307
rect 108 239 176 273
rect 108 205 125 239
rect 159 205 176 239
rect 108 171 176 205
rect 108 137 125 171
rect 159 137 176 171
rect 108 119 176 137
rect 226 307 342 319
rect 226 273 267 307
rect 301 273 342 307
rect 226 239 342 273
rect 226 205 267 239
rect 301 205 342 239
rect 226 171 342 205
rect 226 137 267 171
rect 301 137 342 171
rect 226 119 342 137
rect 392 307 460 319
rect 392 273 409 307
rect 443 273 460 307
rect 392 239 460 273
rect 392 205 409 239
rect 443 205 460 239
rect 392 171 460 205
rect 392 137 409 171
rect 443 137 460 171
rect 392 119 460 137
rect 510 307 597 319
rect 510 273 551 307
rect 585 273 597 307
rect 510 239 597 273
rect 510 205 551 239
rect 585 205 597 239
rect 510 171 597 205
rect 510 137 551 171
rect 585 137 597 171
rect 510 119 597 137
<< pdiff >>
rect -29 743 58 761
rect -29 709 -17 743
rect 17 709 58 743
rect -29 675 58 709
rect -29 641 -17 675
rect 17 641 58 675
rect -29 607 58 641
rect -29 573 -17 607
rect 17 573 58 607
rect -29 561 58 573
rect 108 743 176 761
rect 108 709 125 743
rect 159 709 176 743
rect 108 675 176 709
rect 108 641 125 675
rect 159 641 176 675
rect 108 607 176 641
rect 108 573 125 607
rect 159 573 176 607
rect 108 561 176 573
rect 226 743 342 761
rect 226 709 267 743
rect 301 709 342 743
rect 226 675 342 709
rect 226 641 267 675
rect 301 641 342 675
rect 226 607 342 641
rect 226 573 267 607
rect 301 573 342 607
rect 226 561 342 573
rect 392 743 460 761
rect 392 709 409 743
rect 443 709 460 743
rect 392 675 460 709
rect 392 641 409 675
rect 443 641 460 675
rect 392 607 460 641
rect 392 573 409 607
rect 443 573 460 607
rect 392 561 460 573
rect 510 743 597 761
rect 510 709 551 743
rect 585 709 597 743
rect 510 675 597 709
rect 510 641 551 675
rect 585 641 597 675
rect 510 607 597 641
rect 510 573 551 607
rect 585 573 597 607
rect 510 561 597 573
<< ndiffc >>
rect -17 273 17 307
rect -17 205 17 239
rect -17 137 17 171
rect 125 273 159 307
rect 125 205 159 239
rect 125 137 159 171
rect 267 273 301 307
rect 267 205 301 239
rect 267 137 301 171
rect 409 273 443 307
rect 409 205 443 239
rect 409 137 443 171
rect 551 273 585 307
rect 551 205 585 239
rect 551 137 585 171
<< pdiffc >>
rect -17 709 17 743
rect -17 641 17 675
rect -17 573 17 607
rect 125 709 159 743
rect 125 641 159 675
rect 125 573 159 607
rect 267 709 301 743
rect 267 641 301 675
rect 267 573 301 607
rect 409 709 443 743
rect 409 641 443 675
rect 409 573 443 607
rect 551 709 585 743
rect 551 641 585 675
rect 551 573 585 607
<< psubdiff >>
rect -41 407 41 409
rect -41 373 -17 407
rect 17 373 41 407
rect 243 407 325 409
rect 243 373 267 407
rect 301 373 325 407
rect 527 407 609 409
rect 527 373 551 407
rect 585 373 609 407
<< nsubdiff >>
rect -41 473 -17 507
rect 17 473 41 507
rect -41 471 41 473
rect 243 473 267 507
rect 301 473 325 507
rect 243 471 325 473
rect 527 473 551 507
rect 585 473 609 507
rect 527 471 609 473
<< psubdiffcont >>
rect -17 373 17 407
rect 267 373 301 407
rect 551 373 585 407
<< nsubdiffcont >>
rect -17 473 17 507
rect 267 473 301 507
rect 551 473 585 507
<< poly >>
rect 35 843 533 859
rect 35 809 51 843
rect 85 809 199 843
rect 233 809 335 843
rect 369 809 483 843
rect 517 809 533 843
rect 35 793 533 809
rect 58 761 108 793
rect 176 761 226 793
rect 342 761 392 793
rect 460 761 510 793
rect 58 319 108 561
rect 176 319 226 561
rect 342 319 392 561
rect 460 319 510 561
rect 58 87 108 119
rect 176 87 226 119
rect 342 87 392 119
rect 460 87 510 119
rect 35 71 533 87
rect 35 37 51 71
rect 85 37 199 71
rect 233 37 335 71
rect 369 37 483 71
rect 517 37 533 71
rect 35 21 533 37
<< polycont >>
rect 51 809 85 843
rect 199 809 233 843
rect 335 809 369 843
rect 483 809 517 843
rect 51 37 85 71
rect 199 37 233 71
rect 335 37 369 71
rect 483 37 517 71
<< locali >>
rect 51 843 85 859
rect -17 743 17 759
rect -17 675 17 709
rect -17 607 17 629
rect -17 507 17 523
rect -17 457 17 460
rect -17 420 17 423
rect -17 357 17 373
rect -17 251 17 273
rect -17 171 17 205
rect -17 121 17 137
rect 51 71 85 809
rect 51 21 85 37
rect 125 743 159 859
rect 125 675 159 709
rect 125 607 159 641
rect 125 307 159 573
rect 125 239 159 273
rect 125 171 159 205
rect 125 99 159 137
rect 125 21 159 65
rect 199 843 369 859
rect 233 809 335 843
rect 199 793 369 809
rect 199 87 233 793
rect 267 743 301 759
rect 267 675 301 709
rect 267 607 301 629
rect 267 507 301 523
rect 267 457 301 460
rect 267 420 301 423
rect 267 357 301 373
rect 267 251 301 273
rect 267 171 301 205
rect 267 121 301 137
rect 335 87 369 793
rect 199 71 369 87
rect 233 37 335 71
rect 199 21 369 37
rect 409 743 443 859
rect 409 675 443 709
rect 409 607 443 641
rect 409 307 443 573
rect 409 239 443 273
rect 409 171 443 205
rect 409 99 443 137
rect 409 21 443 65
rect 483 843 517 859
rect 483 71 517 809
rect 551 743 585 759
rect 551 675 585 709
rect 551 607 585 629
rect 551 507 585 523
rect 551 457 585 460
rect 551 420 585 423
rect 551 357 585 373
rect 551 251 585 273
rect 551 171 585 205
rect 551 121 585 137
rect 483 21 517 37
<< viali >>
rect -17 641 17 663
rect -17 629 17 641
rect -17 573 17 591
rect -17 557 17 573
rect -17 473 17 494
rect -17 460 17 473
rect -17 407 17 420
rect -17 386 17 407
rect -17 307 17 323
rect -17 289 17 307
rect -17 239 17 251
rect -17 217 17 239
rect 125 137 159 171
rect 125 65 159 99
rect 267 641 301 663
rect 267 629 301 641
rect 267 573 301 591
rect 267 557 301 573
rect 267 473 301 494
rect 267 460 301 473
rect 267 407 301 420
rect 267 386 301 407
rect 267 307 301 323
rect 267 289 301 307
rect 267 239 301 251
rect 267 217 301 239
rect 409 137 443 171
rect 409 65 443 99
rect 551 641 585 663
rect 551 629 585 641
rect 551 573 585 591
rect 551 557 585 573
rect 551 473 585 494
rect 551 460 585 473
rect 551 407 585 420
rect 551 386 585 407
rect 551 307 585 323
rect 551 289 585 307
rect 551 239 585 251
rect 551 217 585 239
<< metal1 >>
rect -29 663 597 669
rect -29 629 -17 663
rect 17 629 267 663
rect 301 629 551 663
rect 585 629 597 663
rect -29 591 597 629
rect -29 557 -17 591
rect 17 557 267 591
rect 301 557 551 591
rect 585 557 597 591
rect -29 535 597 557
rect -29 494 597 500
rect -29 460 -17 494
rect 17 460 267 494
rect 301 460 551 494
rect 585 460 597 494
rect -29 454 597 460
rect -29 420 597 426
rect -29 386 -17 420
rect 17 386 267 420
rect 301 386 551 420
rect 585 386 597 420
rect -29 380 597 386
rect -29 323 597 346
rect -29 289 -17 323
rect 17 289 267 323
rect 301 289 551 323
rect 585 289 597 323
rect -29 251 597 289
rect -29 217 -17 251
rect 17 217 267 251
rect 301 217 551 251
rect 585 217 597 251
rect -29 211 597 217
rect 119 171 449 183
rect 119 137 125 171
rect 159 155 409 171
rect 159 137 172 155
tri 172 137 190 155 nw
tri 378 137 396 155 ne
rect 396 137 409 155
rect 443 137 449 171
rect 119 99 165 137
tri 165 130 172 137 nw
tri 396 130 403 137 ne
rect 119 65 125 99
rect 159 65 165 99
rect 119 53 165 65
rect 403 99 449 137
rect 403 65 409 99
rect 443 65 449 99
rect 403 53 449 65
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1701704242
transform -1 0 585 0 -1 494
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1701704242
transform -1 0 301 0 -1 494
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1701704242
transform -1 0 17 0 -1 494
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1701704242
transform 1 0 -17 0 1 386
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1701704242
transform 1 0 267 0 1 386
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1701704242
transform 1 0 551 0 1 386
box 0 0 1 1
<< labels >>
flabel comment s 385 32 385 32 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 385 850 385 850 0 FreeSans 100 0 0 0 no_jumper_check
flabel metal1 s -29 211 0 346 0 FreeSans 200 0 0 0 vgnd
port 4 nsew
flabel metal1 s -29 535 0 669 0 FreeSans 200 0 0 0 vpwr
port 3 nsew
flabel metal1 s 568 211 597 346 0 FreeSans 200 0 0 0 vgnd
port 4 nsew
flabel metal1 s 568 535 597 669 0 FreeSans 200 0 0 0 vpwr
port 3 nsew
flabel metal1 s 119 53 165 155 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel metal1 s 403 53 449 155 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel metal1 s 119 155 449 183 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel metal1 s -29 380 0 426 3 FreeSans 400 0 0 0 vnb
port 1 nsew
flabel metal1 s 568 380 597 426 3 FreeSans 400 0 0 0 vnb
port 1 nsew
flabel metal1 s 568 454 597 500 3 FreeSans 400 0 0 0 vpb
port 2 nsew
flabel metal1 s -29 454 0 500 3 FreeSans 400 0 0 0 vpb
port 2 nsew
flabel locali s 51 809 85 859 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel locali s 51 21 85 71 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel locali s 199 21 369 71 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel locali s 483 21 517 71 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel locali s 409 21 443 71 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel locali s 125 21 159 71 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel locali s 125 809 159 859 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel locali s 483 809 517 859 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel locali s 199 809 369 859 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel locali s 409 809 443 859 0 FreeSans 200 0 0 0 out
port 5 nsew
flabel poly s 35 809 533 859 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel poly s 35 21 533 71 0 FreeSans 200 0 0 0 in
port 7 nsew
<< properties >>
string GDS_END 79656178
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79645312
<< end >>
