magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal1 >>
rect 126 1959 156 2011
rect 328 1959 358 2011
rect 1374 1959 1404 2011
rect 1576 1959 1606 2011
rect 2622 1959 2652 2011
rect 2824 1959 2854 2011
rect 3870 1959 3900 2011
rect 4072 1959 4102 2011
rect 5118 1959 5148 2011
rect 5320 1959 5350 2011
rect 6366 1959 6396 2011
rect 6568 1959 6598 2011
rect 7614 1959 7644 2011
rect 7816 1959 7846 2011
rect 8862 1959 8892 2011
rect 9064 1959 9094 2011
rect 10110 1959 10140 2011
rect 10312 1959 10342 2011
rect 11358 1959 11388 2011
rect 11560 1959 11590 2011
rect 12606 1959 12636 2011
rect 12808 1959 12838 2011
rect 13854 1959 13884 2011
rect 14056 1959 14086 2011
rect 15102 1959 15132 2011
rect 15304 1959 15334 2011
rect 16350 1959 16380 2011
rect 16552 1959 16582 2011
rect 17598 1959 17628 2011
rect 17800 1959 17830 2011
rect 18846 1959 18876 2011
rect 19048 1959 19078 2011
rect 20094 1959 20124 2011
rect 20296 1959 20326 2011
rect 21342 1959 21372 2011
rect 21544 1959 21574 2011
rect 22590 1959 22620 2011
rect 22792 1959 22822 2011
rect 23838 1959 23868 2011
rect 24040 1959 24070 2011
rect 25086 1959 25116 2011
rect 25288 1959 25318 2011
rect 26334 1959 26364 2011
rect 26536 1959 26566 2011
rect 27582 1959 27612 2011
rect 27784 1959 27814 2011
rect 28830 1959 28860 2011
rect 29032 1959 29062 2011
rect 30078 1959 30108 2011
rect 30280 1959 30310 2011
rect 31326 1959 31356 2011
rect 31528 1959 31558 2011
rect 32574 1959 32604 2011
rect 32776 1959 32806 2011
rect 33822 1959 33852 2011
rect 34024 1959 34054 2011
rect 35070 1959 35100 2011
rect 35272 1959 35302 2011
rect 36318 1959 36348 2011
rect 36520 1959 36550 2011
rect 37566 1959 37596 2011
rect 37768 1959 37798 2011
rect 38814 1959 38844 2011
rect 39016 1959 39046 2011
rect 241 1604 293 1610
rect 241 1546 293 1552
rect 1489 1604 1541 1610
rect 1489 1546 1541 1552
rect 2737 1604 2789 1610
rect 2737 1546 2789 1552
rect 3985 1604 4037 1610
rect 3985 1546 4037 1552
rect 5233 1604 5285 1610
rect 5233 1546 5285 1552
rect 6481 1604 6533 1610
rect 6481 1546 6533 1552
rect 7729 1604 7781 1610
rect 7729 1546 7781 1552
rect 8977 1604 9029 1610
rect 8977 1546 9029 1552
rect 10225 1604 10277 1610
rect 10225 1546 10277 1552
rect 11473 1604 11525 1610
rect 11473 1546 11525 1552
rect 12721 1604 12773 1610
rect 12721 1546 12773 1552
rect 13969 1604 14021 1610
rect 13969 1546 14021 1552
rect 15217 1604 15269 1610
rect 15217 1546 15269 1552
rect 16465 1604 16517 1610
rect 16465 1546 16517 1552
rect 17713 1604 17765 1610
rect 17713 1546 17765 1552
rect 18961 1604 19013 1610
rect 18961 1546 19013 1552
rect 20209 1604 20261 1610
rect 20209 1546 20261 1552
rect 21457 1604 21509 1610
rect 21457 1546 21509 1552
rect 22705 1604 22757 1610
rect 22705 1546 22757 1552
rect 23953 1604 24005 1610
rect 23953 1546 24005 1552
rect 25201 1604 25253 1610
rect 25201 1546 25253 1552
rect 26449 1604 26501 1610
rect 26449 1546 26501 1552
rect 27697 1604 27749 1610
rect 27697 1546 27749 1552
rect 28945 1604 28997 1610
rect 28945 1546 28997 1552
rect 30193 1604 30245 1610
rect 30193 1546 30245 1552
rect 31441 1604 31493 1610
rect 31441 1546 31493 1552
rect 32689 1604 32741 1610
rect 32689 1546 32741 1552
rect 33937 1604 33989 1610
rect 33937 1546 33989 1552
rect 35185 1604 35237 1610
rect 35185 1546 35237 1552
rect 36433 1604 36485 1610
rect 36433 1546 36485 1552
rect 37681 1604 37733 1610
rect 37681 1546 37733 1552
rect 38929 1604 38981 1610
rect 38929 1546 38981 1552
rect 230 1167 282 1173
rect 230 1109 282 1115
rect 1478 1167 1530 1173
rect 1478 1109 1530 1115
rect 2726 1167 2778 1173
rect 2726 1109 2778 1115
rect 3974 1167 4026 1173
rect 3974 1109 4026 1115
rect 5222 1167 5274 1173
rect 5222 1109 5274 1115
rect 6470 1167 6522 1173
rect 6470 1109 6522 1115
rect 7718 1167 7770 1173
rect 7718 1109 7770 1115
rect 8966 1167 9018 1173
rect 8966 1109 9018 1115
rect 10214 1167 10266 1173
rect 10214 1109 10266 1115
rect 11462 1167 11514 1173
rect 11462 1109 11514 1115
rect 12710 1167 12762 1173
rect 12710 1109 12762 1115
rect 13958 1167 14010 1173
rect 13958 1109 14010 1115
rect 15206 1167 15258 1173
rect 15206 1109 15258 1115
rect 16454 1167 16506 1173
rect 16454 1109 16506 1115
rect 17702 1167 17754 1173
rect 17702 1109 17754 1115
rect 18950 1167 19002 1173
rect 18950 1109 19002 1115
rect 20198 1167 20250 1173
rect 20198 1109 20250 1115
rect 21446 1167 21498 1173
rect 21446 1109 21498 1115
rect 22694 1167 22746 1173
rect 22694 1109 22746 1115
rect 23942 1167 23994 1173
rect 23942 1109 23994 1115
rect 25190 1167 25242 1173
rect 25190 1109 25242 1115
rect 26438 1167 26490 1173
rect 26438 1109 26490 1115
rect 27686 1167 27738 1173
rect 27686 1109 27738 1115
rect 28934 1167 28986 1173
rect 28934 1109 28986 1115
rect 30182 1167 30234 1173
rect 30182 1109 30234 1115
rect 31430 1167 31482 1173
rect 31430 1109 31482 1115
rect 32678 1167 32730 1173
rect 32678 1109 32730 1115
rect 33926 1167 33978 1173
rect 33926 1109 33978 1115
rect 35174 1167 35226 1173
rect 35174 1109 35226 1115
rect 36422 1167 36474 1173
rect 36422 1109 36474 1115
rect 37670 1167 37722 1173
rect 37670 1109 37722 1115
rect 38918 1167 38970 1173
rect 38918 1109 38970 1115
rect 351 836 403 842
rect 351 778 403 784
rect 1599 836 1651 842
rect 1599 778 1651 784
rect 2847 836 2899 842
rect 2847 778 2899 784
rect 4095 836 4147 842
rect 4095 778 4147 784
rect 5343 836 5395 842
rect 5343 778 5395 784
rect 6591 836 6643 842
rect 6591 778 6643 784
rect 7839 836 7891 842
rect 7839 778 7891 784
rect 9087 836 9139 842
rect 9087 778 9139 784
rect 10335 836 10387 842
rect 10335 778 10387 784
rect 11583 836 11635 842
rect 11583 778 11635 784
rect 12831 836 12883 842
rect 12831 778 12883 784
rect 14079 836 14131 842
rect 14079 778 14131 784
rect 15327 836 15379 842
rect 15327 778 15379 784
rect 16575 836 16627 842
rect 16575 778 16627 784
rect 17823 836 17875 842
rect 17823 778 17875 784
rect 19071 836 19123 842
rect 19071 778 19123 784
rect 20319 836 20371 842
rect 20319 778 20371 784
rect 21567 836 21619 842
rect 21567 778 21619 784
rect 22815 836 22867 842
rect 22815 778 22867 784
rect 24063 836 24115 842
rect 24063 778 24115 784
rect 25311 836 25363 842
rect 25311 778 25363 784
rect 26559 836 26611 842
rect 26559 778 26611 784
rect 27807 836 27859 842
rect 27807 778 27859 784
rect 29055 836 29107 842
rect 29055 778 29107 784
rect 30303 836 30355 842
rect 30303 778 30355 784
rect 31551 836 31603 842
rect 31551 778 31603 784
rect 32799 836 32851 842
rect 32799 778 32851 784
rect 34047 836 34099 842
rect 34047 778 34099 784
rect 35295 836 35347 842
rect 35295 778 35347 784
rect 36543 836 36595 842
rect 36543 778 36595 784
rect 37791 836 37843 842
rect 37791 778 37843 784
rect 39039 836 39091 842
rect 39039 778 39091 784
rect 236 633 288 639
rect 236 575 288 581
rect 1484 633 1536 639
rect 1484 575 1536 581
rect 2732 633 2784 639
rect 2732 575 2784 581
rect 3980 633 4032 639
rect 3980 575 4032 581
rect 5228 633 5280 639
rect 5228 575 5280 581
rect 6476 633 6528 639
rect 6476 575 6528 581
rect 7724 633 7776 639
rect 7724 575 7776 581
rect 8972 633 9024 639
rect 8972 575 9024 581
rect 10220 633 10272 639
rect 10220 575 10272 581
rect 11468 633 11520 639
rect 11468 575 11520 581
rect 12716 633 12768 639
rect 12716 575 12768 581
rect 13964 633 14016 639
rect 13964 575 14016 581
rect 15212 633 15264 639
rect 15212 575 15264 581
rect 16460 633 16512 639
rect 16460 575 16512 581
rect 17708 633 17760 639
rect 17708 575 17760 581
rect 18956 633 19008 639
rect 18956 575 19008 581
rect 20204 633 20256 639
rect 20204 575 20256 581
rect 21452 633 21504 639
rect 21452 575 21504 581
rect 22700 633 22752 639
rect 22700 575 22752 581
rect 23948 633 24000 639
rect 23948 575 24000 581
rect 25196 633 25248 639
rect 25196 575 25248 581
rect 26444 633 26496 639
rect 26444 575 26496 581
rect 27692 633 27744 639
rect 27692 575 27744 581
rect 28940 633 28992 639
rect 28940 575 28992 581
rect 30188 633 30240 639
rect 30188 575 30240 581
rect 31436 633 31488 639
rect 31436 575 31488 581
rect 32684 633 32736 639
rect 32684 575 32736 581
rect 33932 633 33984 639
rect 33932 575 33984 581
rect 35180 633 35232 639
rect 35180 575 35232 581
rect 36428 633 36480 639
rect 36428 575 36480 581
rect 37676 633 37728 639
rect 37676 575 37728 581
rect 38924 633 38976 639
rect 38924 575 38976 581
rect 250 217 302 223
rect 250 159 302 165
rect 1498 217 1550 223
rect 1498 159 1550 165
rect 2746 217 2798 223
rect 2746 159 2798 165
rect 3994 217 4046 223
rect 3994 159 4046 165
rect 5242 217 5294 223
rect 5242 159 5294 165
rect 6490 217 6542 223
rect 6490 159 6542 165
rect 7738 217 7790 223
rect 7738 159 7790 165
rect 8986 217 9038 223
rect 8986 159 9038 165
rect 10234 217 10286 223
rect 10234 159 10286 165
rect 11482 217 11534 223
rect 11482 159 11534 165
rect 12730 217 12782 223
rect 12730 159 12782 165
rect 13978 217 14030 223
rect 13978 159 14030 165
rect 15226 217 15278 223
rect 15226 159 15278 165
rect 16474 217 16526 223
rect 16474 159 16526 165
rect 17722 217 17774 223
rect 17722 159 17774 165
rect 18970 217 19022 223
rect 18970 159 19022 165
rect 20218 217 20270 223
rect 20218 159 20270 165
rect 21466 217 21518 223
rect 21466 159 21518 165
rect 22714 217 22766 223
rect 22714 159 22766 165
rect 23962 217 24014 223
rect 23962 159 24014 165
rect 25210 217 25262 223
rect 25210 159 25262 165
rect 26458 217 26510 223
rect 26458 159 26510 165
rect 27706 217 27758 223
rect 27706 159 27758 165
rect 28954 217 29006 223
rect 28954 159 29006 165
rect 30202 217 30254 223
rect 30202 159 30254 165
rect 31450 217 31502 223
rect 31450 159 31502 165
rect 32698 217 32750 223
rect 32698 159 32750 165
rect 33946 217 33998 223
rect 33946 159 33998 165
rect 35194 217 35246 223
rect 35194 159 35246 165
rect 36442 217 36494 223
rect 36442 159 36494 165
rect 37690 217 37742 223
rect 37690 159 37742 165
rect 38938 217 38990 223
rect 38938 159 38990 165
rect 99 94 9459 128
rect 10083 94 19443 128
rect 20067 94 29427 128
rect 30051 94 39411 128
rect 255 4 315 60
rect 1503 4 1563 60
rect 2751 4 2811 60
rect 3999 4 4059 60
rect 5247 4 5307 60
rect 6495 4 6555 60
rect 7743 4 7803 60
rect 8991 4 9051 60
rect 10239 4 10299 60
rect 11487 4 11547 60
rect 12735 4 12795 60
rect 13983 4 14043 60
rect 15231 4 15291 60
rect 16479 4 16539 60
rect 17727 4 17787 60
rect 18975 4 19035 60
rect 20223 4 20283 60
rect 21471 4 21531 60
rect 22719 4 22779 60
rect 23967 4 24027 60
rect 25215 4 25275 60
rect 26463 4 26523 60
rect 27711 4 27771 60
rect 28959 4 29019 60
rect 30207 4 30267 60
rect 31455 4 31515 60
rect 32703 4 32763 60
rect 33951 4 34011 60
rect 35199 4 35259 60
rect 36447 4 36507 60
rect 37695 4 37755 60
rect 38943 4 39003 60
<< via1 >>
rect 241 1552 293 1604
rect 1489 1552 1541 1604
rect 2737 1552 2789 1604
rect 3985 1552 4037 1604
rect 5233 1552 5285 1604
rect 6481 1552 6533 1604
rect 7729 1552 7781 1604
rect 8977 1552 9029 1604
rect 10225 1552 10277 1604
rect 11473 1552 11525 1604
rect 12721 1552 12773 1604
rect 13969 1552 14021 1604
rect 15217 1552 15269 1604
rect 16465 1552 16517 1604
rect 17713 1552 17765 1604
rect 18961 1552 19013 1604
rect 20209 1552 20261 1604
rect 21457 1552 21509 1604
rect 22705 1552 22757 1604
rect 23953 1552 24005 1604
rect 25201 1552 25253 1604
rect 26449 1552 26501 1604
rect 27697 1552 27749 1604
rect 28945 1552 28997 1604
rect 30193 1552 30245 1604
rect 31441 1552 31493 1604
rect 32689 1552 32741 1604
rect 33937 1552 33989 1604
rect 35185 1552 35237 1604
rect 36433 1552 36485 1604
rect 37681 1552 37733 1604
rect 38929 1552 38981 1604
rect 230 1115 282 1167
rect 1478 1115 1530 1167
rect 2726 1115 2778 1167
rect 3974 1115 4026 1167
rect 5222 1115 5274 1167
rect 6470 1115 6522 1167
rect 7718 1115 7770 1167
rect 8966 1115 9018 1167
rect 10214 1115 10266 1167
rect 11462 1115 11514 1167
rect 12710 1115 12762 1167
rect 13958 1115 14010 1167
rect 15206 1115 15258 1167
rect 16454 1115 16506 1167
rect 17702 1115 17754 1167
rect 18950 1115 19002 1167
rect 20198 1115 20250 1167
rect 21446 1115 21498 1167
rect 22694 1115 22746 1167
rect 23942 1115 23994 1167
rect 25190 1115 25242 1167
rect 26438 1115 26490 1167
rect 27686 1115 27738 1167
rect 28934 1115 28986 1167
rect 30182 1115 30234 1167
rect 31430 1115 31482 1167
rect 32678 1115 32730 1167
rect 33926 1115 33978 1167
rect 35174 1115 35226 1167
rect 36422 1115 36474 1167
rect 37670 1115 37722 1167
rect 38918 1115 38970 1167
rect 351 784 403 836
rect 1599 784 1651 836
rect 2847 784 2899 836
rect 4095 784 4147 836
rect 5343 784 5395 836
rect 6591 784 6643 836
rect 7839 784 7891 836
rect 9087 784 9139 836
rect 10335 784 10387 836
rect 11583 784 11635 836
rect 12831 784 12883 836
rect 14079 784 14131 836
rect 15327 784 15379 836
rect 16575 784 16627 836
rect 17823 784 17875 836
rect 19071 784 19123 836
rect 20319 784 20371 836
rect 21567 784 21619 836
rect 22815 784 22867 836
rect 24063 784 24115 836
rect 25311 784 25363 836
rect 26559 784 26611 836
rect 27807 784 27859 836
rect 29055 784 29107 836
rect 30303 784 30355 836
rect 31551 784 31603 836
rect 32799 784 32851 836
rect 34047 784 34099 836
rect 35295 784 35347 836
rect 36543 784 36595 836
rect 37791 784 37843 836
rect 39039 784 39091 836
rect 236 581 288 633
rect 1484 581 1536 633
rect 2732 581 2784 633
rect 3980 581 4032 633
rect 5228 581 5280 633
rect 6476 581 6528 633
rect 7724 581 7776 633
rect 8972 581 9024 633
rect 10220 581 10272 633
rect 11468 581 11520 633
rect 12716 581 12768 633
rect 13964 581 14016 633
rect 15212 581 15264 633
rect 16460 581 16512 633
rect 17708 581 17760 633
rect 18956 581 19008 633
rect 20204 581 20256 633
rect 21452 581 21504 633
rect 22700 581 22752 633
rect 23948 581 24000 633
rect 25196 581 25248 633
rect 26444 581 26496 633
rect 27692 581 27744 633
rect 28940 581 28992 633
rect 30188 581 30240 633
rect 31436 581 31488 633
rect 32684 581 32736 633
rect 33932 581 33984 633
rect 35180 581 35232 633
rect 36428 581 36480 633
rect 37676 581 37728 633
rect 38924 581 38976 633
rect 250 165 302 217
rect 1498 165 1550 217
rect 2746 165 2798 217
rect 3994 165 4046 217
rect 5242 165 5294 217
rect 6490 165 6542 217
rect 7738 165 7790 217
rect 8986 165 9038 217
rect 10234 165 10286 217
rect 11482 165 11534 217
rect 12730 165 12782 217
rect 13978 165 14030 217
rect 15226 165 15278 217
rect 16474 165 16526 217
rect 17722 165 17774 217
rect 18970 165 19022 217
rect 20218 165 20270 217
rect 21466 165 21518 217
rect 22714 165 22766 217
rect 23962 165 24014 217
rect 25210 165 25262 217
rect 26458 165 26510 217
rect 27706 165 27758 217
rect 28954 165 29006 217
rect 30202 165 30254 217
rect 31450 165 31502 217
rect 32698 165 32750 217
rect 33946 165 33998 217
rect 35194 165 35246 217
rect 36442 165 36494 217
rect 37690 165 37742 217
rect 38938 165 38990 217
<< metal2 >>
rect 239 1606 295 1615
rect 239 1541 295 1550
rect 1487 1606 1543 1615
rect 1487 1541 1543 1550
rect 2735 1606 2791 1615
rect 2735 1541 2791 1550
rect 3983 1606 4039 1615
rect 3983 1541 4039 1550
rect 5231 1606 5287 1615
rect 5231 1541 5287 1550
rect 6479 1606 6535 1615
rect 6479 1541 6535 1550
rect 7727 1606 7783 1615
rect 7727 1541 7783 1550
rect 8975 1606 9031 1615
rect 8975 1541 9031 1550
rect 10223 1606 10279 1615
rect 10223 1541 10279 1550
rect 11471 1606 11527 1615
rect 11471 1541 11527 1550
rect 12719 1606 12775 1615
rect 12719 1541 12775 1550
rect 13967 1606 14023 1615
rect 13967 1541 14023 1550
rect 15215 1606 15271 1615
rect 15215 1541 15271 1550
rect 16463 1606 16519 1615
rect 16463 1541 16519 1550
rect 17711 1606 17767 1615
rect 17711 1541 17767 1550
rect 18959 1606 19015 1615
rect 18959 1541 19015 1550
rect 20207 1606 20263 1615
rect 20207 1541 20263 1550
rect 21455 1606 21511 1615
rect 21455 1541 21511 1550
rect 22703 1606 22759 1615
rect 22703 1541 22759 1550
rect 23951 1606 24007 1615
rect 23951 1541 24007 1550
rect 25199 1606 25255 1615
rect 25199 1541 25255 1550
rect 26447 1606 26503 1615
rect 26447 1541 26503 1550
rect 27695 1606 27751 1615
rect 27695 1541 27751 1550
rect 28943 1606 28999 1615
rect 28943 1541 28999 1550
rect 30191 1606 30247 1615
rect 30191 1541 30247 1550
rect 31439 1606 31495 1615
rect 31439 1541 31495 1550
rect 32687 1606 32743 1615
rect 32687 1541 32743 1550
rect 33935 1606 33991 1615
rect 33935 1541 33991 1550
rect 35183 1606 35239 1615
rect 35183 1541 35239 1550
rect 36431 1606 36487 1615
rect 36431 1541 36487 1550
rect 37679 1606 37735 1615
rect 37679 1541 37735 1550
rect 38927 1606 38983 1615
rect 38927 1541 38983 1550
rect 228 1169 284 1178
rect 228 1104 284 1113
rect 1476 1169 1532 1178
rect 1476 1104 1532 1113
rect 2724 1169 2780 1178
rect 2724 1104 2780 1113
rect 3972 1169 4028 1178
rect 3972 1104 4028 1113
rect 5220 1169 5276 1178
rect 5220 1104 5276 1113
rect 6468 1169 6524 1178
rect 6468 1104 6524 1113
rect 7716 1169 7772 1178
rect 7716 1104 7772 1113
rect 8964 1169 9020 1178
rect 8964 1104 9020 1113
rect 10212 1169 10268 1178
rect 10212 1104 10268 1113
rect 11460 1169 11516 1178
rect 11460 1104 11516 1113
rect 12708 1169 12764 1178
rect 12708 1104 12764 1113
rect 13956 1169 14012 1178
rect 13956 1104 14012 1113
rect 15204 1169 15260 1178
rect 15204 1104 15260 1113
rect 16452 1169 16508 1178
rect 16452 1104 16508 1113
rect 17700 1169 17756 1178
rect 17700 1104 17756 1113
rect 18948 1169 19004 1178
rect 18948 1104 19004 1113
rect 20196 1169 20252 1178
rect 20196 1104 20252 1113
rect 21444 1169 21500 1178
rect 21444 1104 21500 1113
rect 22692 1169 22748 1178
rect 22692 1104 22748 1113
rect 23940 1169 23996 1178
rect 23940 1104 23996 1113
rect 25188 1169 25244 1178
rect 25188 1104 25244 1113
rect 26436 1169 26492 1178
rect 26436 1104 26492 1113
rect 27684 1169 27740 1178
rect 27684 1104 27740 1113
rect 28932 1169 28988 1178
rect 28932 1104 28988 1113
rect 30180 1169 30236 1178
rect 30180 1104 30236 1113
rect 31428 1169 31484 1178
rect 31428 1104 31484 1113
rect 32676 1169 32732 1178
rect 32676 1104 32732 1113
rect 33924 1169 33980 1178
rect 33924 1104 33980 1113
rect 35172 1169 35228 1178
rect 35172 1104 35228 1113
rect 36420 1169 36476 1178
rect 36420 1104 36476 1113
rect 37668 1169 37724 1178
rect 37668 1104 37724 1113
rect 38916 1169 38972 1178
rect 38916 1104 38972 1113
rect 349 837 405 846
rect 349 772 405 781
rect 1597 837 1653 846
rect 1597 772 1653 781
rect 2845 837 2901 846
rect 2845 772 2901 781
rect 4093 837 4149 846
rect 4093 772 4149 781
rect 5341 837 5397 846
rect 5341 772 5397 781
rect 6589 837 6645 846
rect 6589 772 6645 781
rect 7837 837 7893 846
rect 7837 772 7893 781
rect 9085 837 9141 846
rect 9085 772 9141 781
rect 10333 837 10389 846
rect 10333 772 10389 781
rect 11581 837 11637 846
rect 11581 772 11637 781
rect 12829 837 12885 846
rect 12829 772 12885 781
rect 14077 837 14133 846
rect 14077 772 14133 781
rect 15325 837 15381 846
rect 15325 772 15381 781
rect 16573 837 16629 846
rect 16573 772 16629 781
rect 17821 837 17877 846
rect 17821 772 17877 781
rect 19069 837 19125 846
rect 19069 772 19125 781
rect 20317 837 20373 846
rect 20317 772 20373 781
rect 21565 837 21621 846
rect 21565 772 21621 781
rect 22813 837 22869 846
rect 22813 772 22869 781
rect 24061 837 24117 846
rect 24061 772 24117 781
rect 25309 837 25365 846
rect 25309 772 25365 781
rect 26557 837 26613 846
rect 26557 772 26613 781
rect 27805 837 27861 846
rect 27805 772 27861 781
rect 29053 837 29109 846
rect 29053 772 29109 781
rect 30301 837 30357 846
rect 30301 772 30357 781
rect 31549 837 31605 846
rect 31549 772 31605 781
rect 32797 837 32853 846
rect 32797 772 32853 781
rect 34045 837 34101 846
rect 34045 772 34101 781
rect 35293 837 35349 846
rect 35293 772 35349 781
rect 36541 837 36597 846
rect 36541 772 36597 781
rect 37789 837 37845 846
rect 37789 772 37845 781
rect 39037 837 39093 846
rect 39037 772 39093 781
rect 234 635 290 644
rect 234 570 290 579
rect 1482 635 1538 644
rect 1482 570 1538 579
rect 2730 635 2786 644
rect 2730 570 2786 579
rect 3978 635 4034 644
rect 3978 570 4034 579
rect 5226 635 5282 644
rect 5226 570 5282 579
rect 6474 635 6530 644
rect 6474 570 6530 579
rect 7722 635 7778 644
rect 7722 570 7778 579
rect 8970 635 9026 644
rect 8970 570 9026 579
rect 10218 635 10274 644
rect 10218 570 10274 579
rect 11466 635 11522 644
rect 11466 570 11522 579
rect 12714 635 12770 644
rect 12714 570 12770 579
rect 13962 635 14018 644
rect 13962 570 14018 579
rect 15210 635 15266 644
rect 15210 570 15266 579
rect 16458 635 16514 644
rect 16458 570 16514 579
rect 17706 635 17762 644
rect 17706 570 17762 579
rect 18954 635 19010 644
rect 18954 570 19010 579
rect 20202 635 20258 644
rect 20202 570 20258 579
rect 21450 635 21506 644
rect 21450 570 21506 579
rect 22698 635 22754 644
rect 22698 570 22754 579
rect 23946 635 24002 644
rect 23946 570 24002 579
rect 25194 635 25250 644
rect 25194 570 25250 579
rect 26442 635 26498 644
rect 26442 570 26498 579
rect 27690 635 27746 644
rect 27690 570 27746 579
rect 28938 635 28994 644
rect 28938 570 28994 579
rect 30186 635 30242 644
rect 30186 570 30242 579
rect 31434 635 31490 644
rect 31434 570 31490 579
rect 32682 635 32738 644
rect 32682 570 32738 579
rect 33930 635 33986 644
rect 33930 570 33986 579
rect 35178 635 35234 644
rect 35178 570 35234 579
rect 36426 635 36482 644
rect 36426 570 36482 579
rect 37674 635 37730 644
rect 37674 570 37730 579
rect 38922 635 38978 644
rect 38922 570 38978 579
rect 248 219 304 228
rect 248 154 304 163
rect 1496 219 1552 228
rect 1496 154 1552 163
rect 2744 219 2800 228
rect 2744 154 2800 163
rect 3992 219 4048 228
rect 3992 154 4048 163
rect 5240 219 5296 228
rect 5240 154 5296 163
rect 6488 219 6544 228
rect 6488 154 6544 163
rect 7736 219 7792 228
rect 7736 154 7792 163
rect 8984 219 9040 228
rect 8984 154 9040 163
rect 10232 219 10288 228
rect 10232 154 10288 163
rect 11480 219 11536 228
rect 11480 154 11536 163
rect 12728 219 12784 228
rect 12728 154 12784 163
rect 13976 219 14032 228
rect 13976 154 14032 163
rect 15224 219 15280 228
rect 15224 154 15280 163
rect 16472 219 16528 228
rect 16472 154 16528 163
rect 17720 219 17776 228
rect 17720 154 17776 163
rect 18968 219 19024 228
rect 18968 154 19024 163
rect 20216 219 20272 228
rect 20216 154 20272 163
rect 21464 219 21520 228
rect 21464 154 21520 163
rect 22712 219 22768 228
rect 22712 154 22768 163
rect 23960 219 24016 228
rect 23960 154 24016 163
rect 25208 219 25264 228
rect 25208 154 25264 163
rect 26456 219 26512 228
rect 26456 154 26512 163
rect 27704 219 27760 228
rect 27704 154 27760 163
rect 28952 219 29008 228
rect 28952 154 29008 163
rect 30200 219 30256 228
rect 30200 154 30256 163
rect 31448 219 31504 228
rect 31448 154 31504 163
rect 32696 219 32752 228
rect 32696 154 32752 163
rect 33944 219 34000 228
rect 33944 154 34000 163
rect 35192 219 35248 228
rect 35192 154 35248 163
rect 36440 219 36496 228
rect 36440 154 36496 163
rect 37688 219 37744 228
rect 37688 154 37744 163
rect 38936 219 38992 228
rect 38936 154 38992 163
<< via2 >>
rect 239 1604 295 1606
rect 239 1552 241 1604
rect 241 1552 293 1604
rect 293 1552 295 1604
rect 239 1550 295 1552
rect 1487 1604 1543 1606
rect 1487 1552 1489 1604
rect 1489 1552 1541 1604
rect 1541 1552 1543 1604
rect 1487 1550 1543 1552
rect 2735 1604 2791 1606
rect 2735 1552 2737 1604
rect 2737 1552 2789 1604
rect 2789 1552 2791 1604
rect 2735 1550 2791 1552
rect 3983 1604 4039 1606
rect 3983 1552 3985 1604
rect 3985 1552 4037 1604
rect 4037 1552 4039 1604
rect 3983 1550 4039 1552
rect 5231 1604 5287 1606
rect 5231 1552 5233 1604
rect 5233 1552 5285 1604
rect 5285 1552 5287 1604
rect 5231 1550 5287 1552
rect 6479 1604 6535 1606
rect 6479 1552 6481 1604
rect 6481 1552 6533 1604
rect 6533 1552 6535 1604
rect 6479 1550 6535 1552
rect 7727 1604 7783 1606
rect 7727 1552 7729 1604
rect 7729 1552 7781 1604
rect 7781 1552 7783 1604
rect 7727 1550 7783 1552
rect 8975 1604 9031 1606
rect 8975 1552 8977 1604
rect 8977 1552 9029 1604
rect 9029 1552 9031 1604
rect 8975 1550 9031 1552
rect 10223 1604 10279 1606
rect 10223 1552 10225 1604
rect 10225 1552 10277 1604
rect 10277 1552 10279 1604
rect 10223 1550 10279 1552
rect 11471 1604 11527 1606
rect 11471 1552 11473 1604
rect 11473 1552 11525 1604
rect 11525 1552 11527 1604
rect 11471 1550 11527 1552
rect 12719 1604 12775 1606
rect 12719 1552 12721 1604
rect 12721 1552 12773 1604
rect 12773 1552 12775 1604
rect 12719 1550 12775 1552
rect 13967 1604 14023 1606
rect 13967 1552 13969 1604
rect 13969 1552 14021 1604
rect 14021 1552 14023 1604
rect 13967 1550 14023 1552
rect 15215 1604 15271 1606
rect 15215 1552 15217 1604
rect 15217 1552 15269 1604
rect 15269 1552 15271 1604
rect 15215 1550 15271 1552
rect 16463 1604 16519 1606
rect 16463 1552 16465 1604
rect 16465 1552 16517 1604
rect 16517 1552 16519 1604
rect 16463 1550 16519 1552
rect 17711 1604 17767 1606
rect 17711 1552 17713 1604
rect 17713 1552 17765 1604
rect 17765 1552 17767 1604
rect 17711 1550 17767 1552
rect 18959 1604 19015 1606
rect 18959 1552 18961 1604
rect 18961 1552 19013 1604
rect 19013 1552 19015 1604
rect 18959 1550 19015 1552
rect 20207 1604 20263 1606
rect 20207 1552 20209 1604
rect 20209 1552 20261 1604
rect 20261 1552 20263 1604
rect 20207 1550 20263 1552
rect 21455 1604 21511 1606
rect 21455 1552 21457 1604
rect 21457 1552 21509 1604
rect 21509 1552 21511 1604
rect 21455 1550 21511 1552
rect 22703 1604 22759 1606
rect 22703 1552 22705 1604
rect 22705 1552 22757 1604
rect 22757 1552 22759 1604
rect 22703 1550 22759 1552
rect 23951 1604 24007 1606
rect 23951 1552 23953 1604
rect 23953 1552 24005 1604
rect 24005 1552 24007 1604
rect 23951 1550 24007 1552
rect 25199 1604 25255 1606
rect 25199 1552 25201 1604
rect 25201 1552 25253 1604
rect 25253 1552 25255 1604
rect 25199 1550 25255 1552
rect 26447 1604 26503 1606
rect 26447 1552 26449 1604
rect 26449 1552 26501 1604
rect 26501 1552 26503 1604
rect 26447 1550 26503 1552
rect 27695 1604 27751 1606
rect 27695 1552 27697 1604
rect 27697 1552 27749 1604
rect 27749 1552 27751 1604
rect 27695 1550 27751 1552
rect 28943 1604 28999 1606
rect 28943 1552 28945 1604
rect 28945 1552 28997 1604
rect 28997 1552 28999 1604
rect 28943 1550 28999 1552
rect 30191 1604 30247 1606
rect 30191 1552 30193 1604
rect 30193 1552 30245 1604
rect 30245 1552 30247 1604
rect 30191 1550 30247 1552
rect 31439 1604 31495 1606
rect 31439 1552 31441 1604
rect 31441 1552 31493 1604
rect 31493 1552 31495 1604
rect 31439 1550 31495 1552
rect 32687 1604 32743 1606
rect 32687 1552 32689 1604
rect 32689 1552 32741 1604
rect 32741 1552 32743 1604
rect 32687 1550 32743 1552
rect 33935 1604 33991 1606
rect 33935 1552 33937 1604
rect 33937 1552 33989 1604
rect 33989 1552 33991 1604
rect 33935 1550 33991 1552
rect 35183 1604 35239 1606
rect 35183 1552 35185 1604
rect 35185 1552 35237 1604
rect 35237 1552 35239 1604
rect 35183 1550 35239 1552
rect 36431 1604 36487 1606
rect 36431 1552 36433 1604
rect 36433 1552 36485 1604
rect 36485 1552 36487 1604
rect 36431 1550 36487 1552
rect 37679 1604 37735 1606
rect 37679 1552 37681 1604
rect 37681 1552 37733 1604
rect 37733 1552 37735 1604
rect 37679 1550 37735 1552
rect 38927 1604 38983 1606
rect 38927 1552 38929 1604
rect 38929 1552 38981 1604
rect 38981 1552 38983 1604
rect 38927 1550 38983 1552
rect 228 1167 284 1169
rect 228 1115 230 1167
rect 230 1115 282 1167
rect 282 1115 284 1167
rect 228 1113 284 1115
rect 1476 1167 1532 1169
rect 1476 1115 1478 1167
rect 1478 1115 1530 1167
rect 1530 1115 1532 1167
rect 1476 1113 1532 1115
rect 2724 1167 2780 1169
rect 2724 1115 2726 1167
rect 2726 1115 2778 1167
rect 2778 1115 2780 1167
rect 2724 1113 2780 1115
rect 3972 1167 4028 1169
rect 3972 1115 3974 1167
rect 3974 1115 4026 1167
rect 4026 1115 4028 1167
rect 3972 1113 4028 1115
rect 5220 1167 5276 1169
rect 5220 1115 5222 1167
rect 5222 1115 5274 1167
rect 5274 1115 5276 1167
rect 5220 1113 5276 1115
rect 6468 1167 6524 1169
rect 6468 1115 6470 1167
rect 6470 1115 6522 1167
rect 6522 1115 6524 1167
rect 6468 1113 6524 1115
rect 7716 1167 7772 1169
rect 7716 1115 7718 1167
rect 7718 1115 7770 1167
rect 7770 1115 7772 1167
rect 7716 1113 7772 1115
rect 8964 1167 9020 1169
rect 8964 1115 8966 1167
rect 8966 1115 9018 1167
rect 9018 1115 9020 1167
rect 8964 1113 9020 1115
rect 10212 1167 10268 1169
rect 10212 1115 10214 1167
rect 10214 1115 10266 1167
rect 10266 1115 10268 1167
rect 10212 1113 10268 1115
rect 11460 1167 11516 1169
rect 11460 1115 11462 1167
rect 11462 1115 11514 1167
rect 11514 1115 11516 1167
rect 11460 1113 11516 1115
rect 12708 1167 12764 1169
rect 12708 1115 12710 1167
rect 12710 1115 12762 1167
rect 12762 1115 12764 1167
rect 12708 1113 12764 1115
rect 13956 1167 14012 1169
rect 13956 1115 13958 1167
rect 13958 1115 14010 1167
rect 14010 1115 14012 1167
rect 13956 1113 14012 1115
rect 15204 1167 15260 1169
rect 15204 1115 15206 1167
rect 15206 1115 15258 1167
rect 15258 1115 15260 1167
rect 15204 1113 15260 1115
rect 16452 1167 16508 1169
rect 16452 1115 16454 1167
rect 16454 1115 16506 1167
rect 16506 1115 16508 1167
rect 16452 1113 16508 1115
rect 17700 1167 17756 1169
rect 17700 1115 17702 1167
rect 17702 1115 17754 1167
rect 17754 1115 17756 1167
rect 17700 1113 17756 1115
rect 18948 1167 19004 1169
rect 18948 1115 18950 1167
rect 18950 1115 19002 1167
rect 19002 1115 19004 1167
rect 18948 1113 19004 1115
rect 20196 1167 20252 1169
rect 20196 1115 20198 1167
rect 20198 1115 20250 1167
rect 20250 1115 20252 1167
rect 20196 1113 20252 1115
rect 21444 1167 21500 1169
rect 21444 1115 21446 1167
rect 21446 1115 21498 1167
rect 21498 1115 21500 1167
rect 21444 1113 21500 1115
rect 22692 1167 22748 1169
rect 22692 1115 22694 1167
rect 22694 1115 22746 1167
rect 22746 1115 22748 1167
rect 22692 1113 22748 1115
rect 23940 1167 23996 1169
rect 23940 1115 23942 1167
rect 23942 1115 23994 1167
rect 23994 1115 23996 1167
rect 23940 1113 23996 1115
rect 25188 1167 25244 1169
rect 25188 1115 25190 1167
rect 25190 1115 25242 1167
rect 25242 1115 25244 1167
rect 25188 1113 25244 1115
rect 26436 1167 26492 1169
rect 26436 1115 26438 1167
rect 26438 1115 26490 1167
rect 26490 1115 26492 1167
rect 26436 1113 26492 1115
rect 27684 1167 27740 1169
rect 27684 1115 27686 1167
rect 27686 1115 27738 1167
rect 27738 1115 27740 1167
rect 27684 1113 27740 1115
rect 28932 1167 28988 1169
rect 28932 1115 28934 1167
rect 28934 1115 28986 1167
rect 28986 1115 28988 1167
rect 28932 1113 28988 1115
rect 30180 1167 30236 1169
rect 30180 1115 30182 1167
rect 30182 1115 30234 1167
rect 30234 1115 30236 1167
rect 30180 1113 30236 1115
rect 31428 1167 31484 1169
rect 31428 1115 31430 1167
rect 31430 1115 31482 1167
rect 31482 1115 31484 1167
rect 31428 1113 31484 1115
rect 32676 1167 32732 1169
rect 32676 1115 32678 1167
rect 32678 1115 32730 1167
rect 32730 1115 32732 1167
rect 32676 1113 32732 1115
rect 33924 1167 33980 1169
rect 33924 1115 33926 1167
rect 33926 1115 33978 1167
rect 33978 1115 33980 1167
rect 33924 1113 33980 1115
rect 35172 1167 35228 1169
rect 35172 1115 35174 1167
rect 35174 1115 35226 1167
rect 35226 1115 35228 1167
rect 35172 1113 35228 1115
rect 36420 1167 36476 1169
rect 36420 1115 36422 1167
rect 36422 1115 36474 1167
rect 36474 1115 36476 1167
rect 36420 1113 36476 1115
rect 37668 1167 37724 1169
rect 37668 1115 37670 1167
rect 37670 1115 37722 1167
rect 37722 1115 37724 1167
rect 37668 1113 37724 1115
rect 38916 1167 38972 1169
rect 38916 1115 38918 1167
rect 38918 1115 38970 1167
rect 38970 1115 38972 1167
rect 38916 1113 38972 1115
rect 349 836 405 837
rect 349 784 351 836
rect 351 784 403 836
rect 403 784 405 836
rect 349 781 405 784
rect 1597 836 1653 837
rect 1597 784 1599 836
rect 1599 784 1651 836
rect 1651 784 1653 836
rect 1597 781 1653 784
rect 2845 836 2901 837
rect 2845 784 2847 836
rect 2847 784 2899 836
rect 2899 784 2901 836
rect 2845 781 2901 784
rect 4093 836 4149 837
rect 4093 784 4095 836
rect 4095 784 4147 836
rect 4147 784 4149 836
rect 4093 781 4149 784
rect 5341 836 5397 837
rect 5341 784 5343 836
rect 5343 784 5395 836
rect 5395 784 5397 836
rect 5341 781 5397 784
rect 6589 836 6645 837
rect 6589 784 6591 836
rect 6591 784 6643 836
rect 6643 784 6645 836
rect 6589 781 6645 784
rect 7837 836 7893 837
rect 7837 784 7839 836
rect 7839 784 7891 836
rect 7891 784 7893 836
rect 7837 781 7893 784
rect 9085 836 9141 837
rect 9085 784 9087 836
rect 9087 784 9139 836
rect 9139 784 9141 836
rect 9085 781 9141 784
rect 10333 836 10389 837
rect 10333 784 10335 836
rect 10335 784 10387 836
rect 10387 784 10389 836
rect 10333 781 10389 784
rect 11581 836 11637 837
rect 11581 784 11583 836
rect 11583 784 11635 836
rect 11635 784 11637 836
rect 11581 781 11637 784
rect 12829 836 12885 837
rect 12829 784 12831 836
rect 12831 784 12883 836
rect 12883 784 12885 836
rect 12829 781 12885 784
rect 14077 836 14133 837
rect 14077 784 14079 836
rect 14079 784 14131 836
rect 14131 784 14133 836
rect 14077 781 14133 784
rect 15325 836 15381 837
rect 15325 784 15327 836
rect 15327 784 15379 836
rect 15379 784 15381 836
rect 15325 781 15381 784
rect 16573 836 16629 837
rect 16573 784 16575 836
rect 16575 784 16627 836
rect 16627 784 16629 836
rect 16573 781 16629 784
rect 17821 836 17877 837
rect 17821 784 17823 836
rect 17823 784 17875 836
rect 17875 784 17877 836
rect 17821 781 17877 784
rect 19069 836 19125 837
rect 19069 784 19071 836
rect 19071 784 19123 836
rect 19123 784 19125 836
rect 19069 781 19125 784
rect 20317 836 20373 837
rect 20317 784 20319 836
rect 20319 784 20371 836
rect 20371 784 20373 836
rect 20317 781 20373 784
rect 21565 836 21621 837
rect 21565 784 21567 836
rect 21567 784 21619 836
rect 21619 784 21621 836
rect 21565 781 21621 784
rect 22813 836 22869 837
rect 22813 784 22815 836
rect 22815 784 22867 836
rect 22867 784 22869 836
rect 22813 781 22869 784
rect 24061 836 24117 837
rect 24061 784 24063 836
rect 24063 784 24115 836
rect 24115 784 24117 836
rect 24061 781 24117 784
rect 25309 836 25365 837
rect 25309 784 25311 836
rect 25311 784 25363 836
rect 25363 784 25365 836
rect 25309 781 25365 784
rect 26557 836 26613 837
rect 26557 784 26559 836
rect 26559 784 26611 836
rect 26611 784 26613 836
rect 26557 781 26613 784
rect 27805 836 27861 837
rect 27805 784 27807 836
rect 27807 784 27859 836
rect 27859 784 27861 836
rect 27805 781 27861 784
rect 29053 836 29109 837
rect 29053 784 29055 836
rect 29055 784 29107 836
rect 29107 784 29109 836
rect 29053 781 29109 784
rect 30301 836 30357 837
rect 30301 784 30303 836
rect 30303 784 30355 836
rect 30355 784 30357 836
rect 30301 781 30357 784
rect 31549 836 31605 837
rect 31549 784 31551 836
rect 31551 784 31603 836
rect 31603 784 31605 836
rect 31549 781 31605 784
rect 32797 836 32853 837
rect 32797 784 32799 836
rect 32799 784 32851 836
rect 32851 784 32853 836
rect 32797 781 32853 784
rect 34045 836 34101 837
rect 34045 784 34047 836
rect 34047 784 34099 836
rect 34099 784 34101 836
rect 34045 781 34101 784
rect 35293 836 35349 837
rect 35293 784 35295 836
rect 35295 784 35347 836
rect 35347 784 35349 836
rect 35293 781 35349 784
rect 36541 836 36597 837
rect 36541 784 36543 836
rect 36543 784 36595 836
rect 36595 784 36597 836
rect 36541 781 36597 784
rect 37789 836 37845 837
rect 37789 784 37791 836
rect 37791 784 37843 836
rect 37843 784 37845 836
rect 37789 781 37845 784
rect 39037 836 39093 837
rect 39037 784 39039 836
rect 39039 784 39091 836
rect 39091 784 39093 836
rect 39037 781 39093 784
rect 234 633 290 635
rect 234 581 236 633
rect 236 581 288 633
rect 288 581 290 633
rect 234 579 290 581
rect 1482 633 1538 635
rect 1482 581 1484 633
rect 1484 581 1536 633
rect 1536 581 1538 633
rect 1482 579 1538 581
rect 2730 633 2786 635
rect 2730 581 2732 633
rect 2732 581 2784 633
rect 2784 581 2786 633
rect 2730 579 2786 581
rect 3978 633 4034 635
rect 3978 581 3980 633
rect 3980 581 4032 633
rect 4032 581 4034 633
rect 3978 579 4034 581
rect 5226 633 5282 635
rect 5226 581 5228 633
rect 5228 581 5280 633
rect 5280 581 5282 633
rect 5226 579 5282 581
rect 6474 633 6530 635
rect 6474 581 6476 633
rect 6476 581 6528 633
rect 6528 581 6530 633
rect 6474 579 6530 581
rect 7722 633 7778 635
rect 7722 581 7724 633
rect 7724 581 7776 633
rect 7776 581 7778 633
rect 7722 579 7778 581
rect 8970 633 9026 635
rect 8970 581 8972 633
rect 8972 581 9024 633
rect 9024 581 9026 633
rect 8970 579 9026 581
rect 10218 633 10274 635
rect 10218 581 10220 633
rect 10220 581 10272 633
rect 10272 581 10274 633
rect 10218 579 10274 581
rect 11466 633 11522 635
rect 11466 581 11468 633
rect 11468 581 11520 633
rect 11520 581 11522 633
rect 11466 579 11522 581
rect 12714 633 12770 635
rect 12714 581 12716 633
rect 12716 581 12768 633
rect 12768 581 12770 633
rect 12714 579 12770 581
rect 13962 633 14018 635
rect 13962 581 13964 633
rect 13964 581 14016 633
rect 14016 581 14018 633
rect 13962 579 14018 581
rect 15210 633 15266 635
rect 15210 581 15212 633
rect 15212 581 15264 633
rect 15264 581 15266 633
rect 15210 579 15266 581
rect 16458 633 16514 635
rect 16458 581 16460 633
rect 16460 581 16512 633
rect 16512 581 16514 633
rect 16458 579 16514 581
rect 17706 633 17762 635
rect 17706 581 17708 633
rect 17708 581 17760 633
rect 17760 581 17762 633
rect 17706 579 17762 581
rect 18954 633 19010 635
rect 18954 581 18956 633
rect 18956 581 19008 633
rect 19008 581 19010 633
rect 18954 579 19010 581
rect 20202 633 20258 635
rect 20202 581 20204 633
rect 20204 581 20256 633
rect 20256 581 20258 633
rect 20202 579 20258 581
rect 21450 633 21506 635
rect 21450 581 21452 633
rect 21452 581 21504 633
rect 21504 581 21506 633
rect 21450 579 21506 581
rect 22698 633 22754 635
rect 22698 581 22700 633
rect 22700 581 22752 633
rect 22752 581 22754 633
rect 22698 579 22754 581
rect 23946 633 24002 635
rect 23946 581 23948 633
rect 23948 581 24000 633
rect 24000 581 24002 633
rect 23946 579 24002 581
rect 25194 633 25250 635
rect 25194 581 25196 633
rect 25196 581 25248 633
rect 25248 581 25250 633
rect 25194 579 25250 581
rect 26442 633 26498 635
rect 26442 581 26444 633
rect 26444 581 26496 633
rect 26496 581 26498 633
rect 26442 579 26498 581
rect 27690 633 27746 635
rect 27690 581 27692 633
rect 27692 581 27744 633
rect 27744 581 27746 633
rect 27690 579 27746 581
rect 28938 633 28994 635
rect 28938 581 28940 633
rect 28940 581 28992 633
rect 28992 581 28994 633
rect 28938 579 28994 581
rect 30186 633 30242 635
rect 30186 581 30188 633
rect 30188 581 30240 633
rect 30240 581 30242 633
rect 30186 579 30242 581
rect 31434 633 31490 635
rect 31434 581 31436 633
rect 31436 581 31488 633
rect 31488 581 31490 633
rect 31434 579 31490 581
rect 32682 633 32738 635
rect 32682 581 32684 633
rect 32684 581 32736 633
rect 32736 581 32738 633
rect 32682 579 32738 581
rect 33930 633 33986 635
rect 33930 581 33932 633
rect 33932 581 33984 633
rect 33984 581 33986 633
rect 33930 579 33986 581
rect 35178 633 35234 635
rect 35178 581 35180 633
rect 35180 581 35232 633
rect 35232 581 35234 633
rect 35178 579 35234 581
rect 36426 633 36482 635
rect 36426 581 36428 633
rect 36428 581 36480 633
rect 36480 581 36482 633
rect 36426 579 36482 581
rect 37674 633 37730 635
rect 37674 581 37676 633
rect 37676 581 37728 633
rect 37728 581 37730 633
rect 37674 579 37730 581
rect 38922 633 38978 635
rect 38922 581 38924 633
rect 38924 581 38976 633
rect 38976 581 38978 633
rect 38922 579 38978 581
rect 248 217 304 219
rect 248 165 250 217
rect 250 165 302 217
rect 302 165 304 217
rect 248 163 304 165
rect 1496 217 1552 219
rect 1496 165 1498 217
rect 1498 165 1550 217
rect 1550 165 1552 217
rect 1496 163 1552 165
rect 2744 217 2800 219
rect 2744 165 2746 217
rect 2746 165 2798 217
rect 2798 165 2800 217
rect 2744 163 2800 165
rect 3992 217 4048 219
rect 3992 165 3994 217
rect 3994 165 4046 217
rect 4046 165 4048 217
rect 3992 163 4048 165
rect 5240 217 5296 219
rect 5240 165 5242 217
rect 5242 165 5294 217
rect 5294 165 5296 217
rect 5240 163 5296 165
rect 6488 217 6544 219
rect 6488 165 6490 217
rect 6490 165 6542 217
rect 6542 165 6544 217
rect 6488 163 6544 165
rect 7736 217 7792 219
rect 7736 165 7738 217
rect 7738 165 7790 217
rect 7790 165 7792 217
rect 7736 163 7792 165
rect 8984 217 9040 219
rect 8984 165 8986 217
rect 8986 165 9038 217
rect 9038 165 9040 217
rect 8984 163 9040 165
rect 10232 217 10288 219
rect 10232 165 10234 217
rect 10234 165 10286 217
rect 10286 165 10288 217
rect 10232 163 10288 165
rect 11480 217 11536 219
rect 11480 165 11482 217
rect 11482 165 11534 217
rect 11534 165 11536 217
rect 11480 163 11536 165
rect 12728 217 12784 219
rect 12728 165 12730 217
rect 12730 165 12782 217
rect 12782 165 12784 217
rect 12728 163 12784 165
rect 13976 217 14032 219
rect 13976 165 13978 217
rect 13978 165 14030 217
rect 14030 165 14032 217
rect 13976 163 14032 165
rect 15224 217 15280 219
rect 15224 165 15226 217
rect 15226 165 15278 217
rect 15278 165 15280 217
rect 15224 163 15280 165
rect 16472 217 16528 219
rect 16472 165 16474 217
rect 16474 165 16526 217
rect 16526 165 16528 217
rect 16472 163 16528 165
rect 17720 217 17776 219
rect 17720 165 17722 217
rect 17722 165 17774 217
rect 17774 165 17776 217
rect 17720 163 17776 165
rect 18968 217 19024 219
rect 18968 165 18970 217
rect 18970 165 19022 217
rect 19022 165 19024 217
rect 18968 163 19024 165
rect 20216 217 20272 219
rect 20216 165 20218 217
rect 20218 165 20270 217
rect 20270 165 20272 217
rect 20216 163 20272 165
rect 21464 217 21520 219
rect 21464 165 21466 217
rect 21466 165 21518 217
rect 21518 165 21520 217
rect 21464 163 21520 165
rect 22712 217 22768 219
rect 22712 165 22714 217
rect 22714 165 22766 217
rect 22766 165 22768 217
rect 22712 163 22768 165
rect 23960 217 24016 219
rect 23960 165 23962 217
rect 23962 165 24014 217
rect 24014 165 24016 217
rect 23960 163 24016 165
rect 25208 217 25264 219
rect 25208 165 25210 217
rect 25210 165 25262 217
rect 25262 165 25264 217
rect 25208 163 25264 165
rect 26456 217 26512 219
rect 26456 165 26458 217
rect 26458 165 26510 217
rect 26510 165 26512 217
rect 26456 163 26512 165
rect 27704 217 27760 219
rect 27704 165 27706 217
rect 27706 165 27758 217
rect 27758 165 27760 217
rect 27704 163 27760 165
rect 28952 217 29008 219
rect 28952 165 28954 217
rect 28954 165 29006 217
rect 29006 165 29008 217
rect 28952 163 29008 165
rect 30200 217 30256 219
rect 30200 165 30202 217
rect 30202 165 30254 217
rect 30254 165 30256 217
rect 30200 163 30256 165
rect 31448 217 31504 219
rect 31448 165 31450 217
rect 31450 165 31502 217
rect 31502 165 31504 217
rect 31448 163 31504 165
rect 32696 217 32752 219
rect 32696 165 32698 217
rect 32698 165 32750 217
rect 32750 165 32752 217
rect 32696 163 32752 165
rect 33944 217 34000 219
rect 33944 165 33946 217
rect 33946 165 33998 217
rect 33998 165 34000 217
rect 33944 163 34000 165
rect 35192 217 35248 219
rect 35192 165 35194 217
rect 35194 165 35246 217
rect 35246 165 35248 217
rect 35192 163 35248 165
rect 36440 217 36496 219
rect 36440 165 36442 217
rect 36442 165 36494 217
rect 36494 165 36496 217
rect 36440 163 36496 165
rect 37688 217 37744 219
rect 37688 165 37690 217
rect 37690 165 37742 217
rect 37742 165 37744 217
rect 37688 163 37744 165
rect 38936 217 38992 219
rect 38936 165 38938 217
rect 38938 165 38990 217
rect 38990 165 38992 217
rect 38936 163 38992 165
<< metal3 >>
rect 218 1606 316 1627
rect 218 1550 239 1606
rect 295 1550 316 1606
rect 218 1529 316 1550
rect 1466 1606 1564 1627
rect 1466 1550 1487 1606
rect 1543 1550 1564 1606
rect 1466 1529 1564 1550
rect 2714 1606 2812 1627
rect 2714 1550 2735 1606
rect 2791 1550 2812 1606
rect 2714 1529 2812 1550
rect 3962 1606 4060 1627
rect 3962 1550 3983 1606
rect 4039 1550 4060 1606
rect 3962 1529 4060 1550
rect 5210 1606 5308 1627
rect 5210 1550 5231 1606
rect 5287 1550 5308 1606
rect 5210 1529 5308 1550
rect 6458 1606 6556 1627
rect 6458 1550 6479 1606
rect 6535 1550 6556 1606
rect 6458 1529 6556 1550
rect 7706 1606 7804 1627
rect 7706 1550 7727 1606
rect 7783 1550 7804 1606
rect 7706 1529 7804 1550
rect 8954 1606 9052 1627
rect 8954 1550 8975 1606
rect 9031 1550 9052 1606
rect 8954 1529 9052 1550
rect 10202 1606 10300 1627
rect 10202 1550 10223 1606
rect 10279 1550 10300 1606
rect 10202 1529 10300 1550
rect 11450 1606 11548 1627
rect 11450 1550 11471 1606
rect 11527 1550 11548 1606
rect 11450 1529 11548 1550
rect 12698 1606 12796 1627
rect 12698 1550 12719 1606
rect 12775 1550 12796 1606
rect 12698 1529 12796 1550
rect 13946 1606 14044 1627
rect 13946 1550 13967 1606
rect 14023 1550 14044 1606
rect 13946 1529 14044 1550
rect 15194 1606 15292 1627
rect 15194 1550 15215 1606
rect 15271 1550 15292 1606
rect 15194 1529 15292 1550
rect 16442 1606 16540 1627
rect 16442 1550 16463 1606
rect 16519 1550 16540 1606
rect 16442 1529 16540 1550
rect 17690 1606 17788 1627
rect 17690 1550 17711 1606
rect 17767 1550 17788 1606
rect 17690 1529 17788 1550
rect 18938 1606 19036 1627
rect 18938 1550 18959 1606
rect 19015 1550 19036 1606
rect 18938 1529 19036 1550
rect 20186 1606 20284 1627
rect 20186 1550 20207 1606
rect 20263 1550 20284 1606
rect 20186 1529 20284 1550
rect 21434 1606 21532 1627
rect 21434 1550 21455 1606
rect 21511 1550 21532 1606
rect 21434 1529 21532 1550
rect 22682 1606 22780 1627
rect 22682 1550 22703 1606
rect 22759 1550 22780 1606
rect 22682 1529 22780 1550
rect 23930 1606 24028 1627
rect 23930 1550 23951 1606
rect 24007 1550 24028 1606
rect 23930 1529 24028 1550
rect 25178 1606 25276 1627
rect 25178 1550 25199 1606
rect 25255 1550 25276 1606
rect 25178 1529 25276 1550
rect 26426 1606 26524 1627
rect 26426 1550 26447 1606
rect 26503 1550 26524 1606
rect 26426 1529 26524 1550
rect 27674 1606 27772 1627
rect 27674 1550 27695 1606
rect 27751 1550 27772 1606
rect 27674 1529 27772 1550
rect 28922 1606 29020 1627
rect 28922 1550 28943 1606
rect 28999 1550 29020 1606
rect 28922 1529 29020 1550
rect 30170 1606 30268 1627
rect 30170 1550 30191 1606
rect 30247 1550 30268 1606
rect 30170 1529 30268 1550
rect 31418 1606 31516 1627
rect 31418 1550 31439 1606
rect 31495 1550 31516 1606
rect 31418 1529 31516 1550
rect 32666 1606 32764 1627
rect 32666 1550 32687 1606
rect 32743 1550 32764 1606
rect 32666 1529 32764 1550
rect 33914 1606 34012 1627
rect 33914 1550 33935 1606
rect 33991 1550 34012 1606
rect 33914 1529 34012 1550
rect 35162 1606 35260 1627
rect 35162 1550 35183 1606
rect 35239 1550 35260 1606
rect 35162 1529 35260 1550
rect 36410 1606 36508 1627
rect 36410 1550 36431 1606
rect 36487 1550 36508 1606
rect 36410 1529 36508 1550
rect 37658 1606 37756 1627
rect 37658 1550 37679 1606
rect 37735 1550 37756 1606
rect 37658 1529 37756 1550
rect 38906 1606 39004 1627
rect 38906 1550 38927 1606
rect 38983 1550 39004 1606
rect 38906 1529 39004 1550
rect 207 1169 305 1190
rect 207 1113 228 1169
rect 284 1113 305 1169
rect 207 1092 305 1113
rect 1455 1169 1553 1190
rect 1455 1113 1476 1169
rect 1532 1113 1553 1169
rect 1455 1092 1553 1113
rect 2703 1169 2801 1190
rect 2703 1113 2724 1169
rect 2780 1113 2801 1169
rect 2703 1092 2801 1113
rect 3951 1169 4049 1190
rect 3951 1113 3972 1169
rect 4028 1113 4049 1169
rect 3951 1092 4049 1113
rect 5199 1169 5297 1190
rect 5199 1113 5220 1169
rect 5276 1113 5297 1169
rect 5199 1092 5297 1113
rect 6447 1169 6545 1190
rect 6447 1113 6468 1169
rect 6524 1113 6545 1169
rect 6447 1092 6545 1113
rect 7695 1169 7793 1190
rect 7695 1113 7716 1169
rect 7772 1113 7793 1169
rect 7695 1092 7793 1113
rect 8943 1169 9041 1190
rect 8943 1113 8964 1169
rect 9020 1113 9041 1169
rect 8943 1092 9041 1113
rect 10191 1169 10289 1190
rect 10191 1113 10212 1169
rect 10268 1113 10289 1169
rect 10191 1092 10289 1113
rect 11439 1169 11537 1190
rect 11439 1113 11460 1169
rect 11516 1113 11537 1169
rect 11439 1092 11537 1113
rect 12687 1169 12785 1190
rect 12687 1113 12708 1169
rect 12764 1113 12785 1169
rect 12687 1092 12785 1113
rect 13935 1169 14033 1190
rect 13935 1113 13956 1169
rect 14012 1113 14033 1169
rect 13935 1092 14033 1113
rect 15183 1169 15281 1190
rect 15183 1113 15204 1169
rect 15260 1113 15281 1169
rect 15183 1092 15281 1113
rect 16431 1169 16529 1190
rect 16431 1113 16452 1169
rect 16508 1113 16529 1169
rect 16431 1092 16529 1113
rect 17679 1169 17777 1190
rect 17679 1113 17700 1169
rect 17756 1113 17777 1169
rect 17679 1092 17777 1113
rect 18927 1169 19025 1190
rect 18927 1113 18948 1169
rect 19004 1113 19025 1169
rect 18927 1092 19025 1113
rect 20175 1169 20273 1190
rect 20175 1113 20196 1169
rect 20252 1113 20273 1169
rect 20175 1092 20273 1113
rect 21423 1169 21521 1190
rect 21423 1113 21444 1169
rect 21500 1113 21521 1169
rect 21423 1092 21521 1113
rect 22671 1169 22769 1190
rect 22671 1113 22692 1169
rect 22748 1113 22769 1169
rect 22671 1092 22769 1113
rect 23919 1169 24017 1190
rect 23919 1113 23940 1169
rect 23996 1113 24017 1169
rect 23919 1092 24017 1113
rect 25167 1169 25265 1190
rect 25167 1113 25188 1169
rect 25244 1113 25265 1169
rect 25167 1092 25265 1113
rect 26415 1169 26513 1190
rect 26415 1113 26436 1169
rect 26492 1113 26513 1169
rect 26415 1092 26513 1113
rect 27663 1169 27761 1190
rect 27663 1113 27684 1169
rect 27740 1113 27761 1169
rect 27663 1092 27761 1113
rect 28911 1169 29009 1190
rect 28911 1113 28932 1169
rect 28988 1113 29009 1169
rect 28911 1092 29009 1113
rect 30159 1169 30257 1190
rect 30159 1113 30180 1169
rect 30236 1113 30257 1169
rect 30159 1092 30257 1113
rect 31407 1169 31505 1190
rect 31407 1113 31428 1169
rect 31484 1113 31505 1169
rect 31407 1092 31505 1113
rect 32655 1169 32753 1190
rect 32655 1113 32676 1169
rect 32732 1113 32753 1169
rect 32655 1092 32753 1113
rect 33903 1169 34001 1190
rect 33903 1113 33924 1169
rect 33980 1113 34001 1169
rect 33903 1092 34001 1113
rect 35151 1169 35249 1190
rect 35151 1113 35172 1169
rect 35228 1113 35249 1169
rect 35151 1092 35249 1113
rect 36399 1169 36497 1190
rect 36399 1113 36420 1169
rect 36476 1113 36497 1169
rect 36399 1092 36497 1113
rect 37647 1169 37745 1190
rect 37647 1113 37668 1169
rect 37724 1113 37745 1169
rect 37647 1092 37745 1113
rect 38895 1169 38993 1190
rect 38895 1113 38916 1169
rect 38972 1113 38993 1169
rect 38895 1092 38993 1113
rect 328 837 426 858
rect 328 781 349 837
rect 405 781 426 837
rect 328 760 426 781
rect 1576 837 1674 858
rect 1576 781 1597 837
rect 1653 781 1674 837
rect 1576 760 1674 781
rect 2824 837 2922 858
rect 2824 781 2845 837
rect 2901 781 2922 837
rect 2824 760 2922 781
rect 4072 837 4170 858
rect 4072 781 4093 837
rect 4149 781 4170 837
rect 4072 760 4170 781
rect 5320 837 5418 858
rect 5320 781 5341 837
rect 5397 781 5418 837
rect 5320 760 5418 781
rect 6568 837 6666 858
rect 6568 781 6589 837
rect 6645 781 6666 837
rect 6568 760 6666 781
rect 7816 837 7914 858
rect 7816 781 7837 837
rect 7893 781 7914 837
rect 7816 760 7914 781
rect 9064 837 9162 858
rect 9064 781 9085 837
rect 9141 781 9162 837
rect 9064 760 9162 781
rect 10312 837 10410 858
rect 10312 781 10333 837
rect 10389 781 10410 837
rect 10312 760 10410 781
rect 11560 837 11658 858
rect 11560 781 11581 837
rect 11637 781 11658 837
rect 11560 760 11658 781
rect 12808 837 12906 858
rect 12808 781 12829 837
rect 12885 781 12906 837
rect 12808 760 12906 781
rect 14056 837 14154 858
rect 14056 781 14077 837
rect 14133 781 14154 837
rect 14056 760 14154 781
rect 15304 837 15402 858
rect 15304 781 15325 837
rect 15381 781 15402 837
rect 15304 760 15402 781
rect 16552 837 16650 858
rect 16552 781 16573 837
rect 16629 781 16650 837
rect 16552 760 16650 781
rect 17800 837 17898 858
rect 17800 781 17821 837
rect 17877 781 17898 837
rect 17800 760 17898 781
rect 19048 837 19146 858
rect 19048 781 19069 837
rect 19125 781 19146 837
rect 19048 760 19146 781
rect 20296 837 20394 858
rect 20296 781 20317 837
rect 20373 781 20394 837
rect 20296 760 20394 781
rect 21544 837 21642 858
rect 21544 781 21565 837
rect 21621 781 21642 837
rect 21544 760 21642 781
rect 22792 837 22890 858
rect 22792 781 22813 837
rect 22869 781 22890 837
rect 22792 760 22890 781
rect 24040 837 24138 858
rect 24040 781 24061 837
rect 24117 781 24138 837
rect 24040 760 24138 781
rect 25288 837 25386 858
rect 25288 781 25309 837
rect 25365 781 25386 837
rect 25288 760 25386 781
rect 26536 837 26634 858
rect 26536 781 26557 837
rect 26613 781 26634 837
rect 26536 760 26634 781
rect 27784 837 27882 858
rect 27784 781 27805 837
rect 27861 781 27882 837
rect 27784 760 27882 781
rect 29032 837 29130 858
rect 29032 781 29053 837
rect 29109 781 29130 837
rect 29032 760 29130 781
rect 30280 837 30378 858
rect 30280 781 30301 837
rect 30357 781 30378 837
rect 30280 760 30378 781
rect 31528 837 31626 858
rect 31528 781 31549 837
rect 31605 781 31626 837
rect 31528 760 31626 781
rect 32776 837 32874 858
rect 32776 781 32797 837
rect 32853 781 32874 837
rect 32776 760 32874 781
rect 34024 837 34122 858
rect 34024 781 34045 837
rect 34101 781 34122 837
rect 34024 760 34122 781
rect 35272 837 35370 858
rect 35272 781 35293 837
rect 35349 781 35370 837
rect 35272 760 35370 781
rect 36520 837 36618 858
rect 36520 781 36541 837
rect 36597 781 36618 837
rect 36520 760 36618 781
rect 37768 837 37866 858
rect 37768 781 37789 837
rect 37845 781 37866 837
rect 37768 760 37866 781
rect 39016 837 39114 858
rect 39016 781 39037 837
rect 39093 781 39114 837
rect 39016 760 39114 781
rect 213 635 311 656
rect 213 579 234 635
rect 290 579 311 635
rect 213 558 311 579
rect 1461 635 1559 656
rect 1461 579 1482 635
rect 1538 579 1559 635
rect 1461 558 1559 579
rect 2709 635 2807 656
rect 2709 579 2730 635
rect 2786 579 2807 635
rect 2709 558 2807 579
rect 3957 635 4055 656
rect 3957 579 3978 635
rect 4034 579 4055 635
rect 3957 558 4055 579
rect 5205 635 5303 656
rect 5205 579 5226 635
rect 5282 579 5303 635
rect 5205 558 5303 579
rect 6453 635 6551 656
rect 6453 579 6474 635
rect 6530 579 6551 635
rect 6453 558 6551 579
rect 7701 635 7799 656
rect 7701 579 7722 635
rect 7778 579 7799 635
rect 7701 558 7799 579
rect 8949 635 9047 656
rect 8949 579 8970 635
rect 9026 579 9047 635
rect 8949 558 9047 579
rect 10197 635 10295 656
rect 10197 579 10218 635
rect 10274 579 10295 635
rect 10197 558 10295 579
rect 11445 635 11543 656
rect 11445 579 11466 635
rect 11522 579 11543 635
rect 11445 558 11543 579
rect 12693 635 12791 656
rect 12693 579 12714 635
rect 12770 579 12791 635
rect 12693 558 12791 579
rect 13941 635 14039 656
rect 13941 579 13962 635
rect 14018 579 14039 635
rect 13941 558 14039 579
rect 15189 635 15287 656
rect 15189 579 15210 635
rect 15266 579 15287 635
rect 15189 558 15287 579
rect 16437 635 16535 656
rect 16437 579 16458 635
rect 16514 579 16535 635
rect 16437 558 16535 579
rect 17685 635 17783 656
rect 17685 579 17706 635
rect 17762 579 17783 635
rect 17685 558 17783 579
rect 18933 635 19031 656
rect 18933 579 18954 635
rect 19010 579 19031 635
rect 18933 558 19031 579
rect 20181 635 20279 656
rect 20181 579 20202 635
rect 20258 579 20279 635
rect 20181 558 20279 579
rect 21429 635 21527 656
rect 21429 579 21450 635
rect 21506 579 21527 635
rect 21429 558 21527 579
rect 22677 635 22775 656
rect 22677 579 22698 635
rect 22754 579 22775 635
rect 22677 558 22775 579
rect 23925 635 24023 656
rect 23925 579 23946 635
rect 24002 579 24023 635
rect 23925 558 24023 579
rect 25173 635 25271 656
rect 25173 579 25194 635
rect 25250 579 25271 635
rect 25173 558 25271 579
rect 26421 635 26519 656
rect 26421 579 26442 635
rect 26498 579 26519 635
rect 26421 558 26519 579
rect 27669 635 27767 656
rect 27669 579 27690 635
rect 27746 579 27767 635
rect 27669 558 27767 579
rect 28917 635 29015 656
rect 28917 579 28938 635
rect 28994 579 29015 635
rect 28917 558 29015 579
rect 30165 635 30263 656
rect 30165 579 30186 635
rect 30242 579 30263 635
rect 30165 558 30263 579
rect 31413 635 31511 656
rect 31413 579 31434 635
rect 31490 579 31511 635
rect 31413 558 31511 579
rect 32661 635 32759 656
rect 32661 579 32682 635
rect 32738 579 32759 635
rect 32661 558 32759 579
rect 33909 635 34007 656
rect 33909 579 33930 635
rect 33986 579 34007 635
rect 33909 558 34007 579
rect 35157 635 35255 656
rect 35157 579 35178 635
rect 35234 579 35255 635
rect 35157 558 35255 579
rect 36405 635 36503 656
rect 36405 579 36426 635
rect 36482 579 36503 635
rect 36405 558 36503 579
rect 37653 635 37751 656
rect 37653 579 37674 635
rect 37730 579 37751 635
rect 37653 558 37751 579
rect 38901 635 38999 656
rect 38901 579 38922 635
rect 38978 579 38999 635
rect 38901 558 38999 579
rect 227 219 325 240
rect 227 163 248 219
rect 304 163 325 219
rect 227 142 325 163
rect 1475 219 1573 240
rect 1475 163 1496 219
rect 1552 163 1573 219
rect 1475 142 1573 163
rect 2723 219 2821 240
rect 2723 163 2744 219
rect 2800 163 2821 219
rect 2723 142 2821 163
rect 3971 219 4069 240
rect 3971 163 3992 219
rect 4048 163 4069 219
rect 3971 142 4069 163
rect 5219 219 5317 240
rect 5219 163 5240 219
rect 5296 163 5317 219
rect 5219 142 5317 163
rect 6467 219 6565 240
rect 6467 163 6488 219
rect 6544 163 6565 219
rect 6467 142 6565 163
rect 7715 219 7813 240
rect 7715 163 7736 219
rect 7792 163 7813 219
rect 7715 142 7813 163
rect 8963 219 9061 240
rect 8963 163 8984 219
rect 9040 163 9061 219
rect 8963 142 9061 163
rect 10211 219 10309 240
rect 10211 163 10232 219
rect 10288 163 10309 219
rect 10211 142 10309 163
rect 11459 219 11557 240
rect 11459 163 11480 219
rect 11536 163 11557 219
rect 11459 142 11557 163
rect 12707 219 12805 240
rect 12707 163 12728 219
rect 12784 163 12805 219
rect 12707 142 12805 163
rect 13955 219 14053 240
rect 13955 163 13976 219
rect 14032 163 14053 219
rect 13955 142 14053 163
rect 15203 219 15301 240
rect 15203 163 15224 219
rect 15280 163 15301 219
rect 15203 142 15301 163
rect 16451 219 16549 240
rect 16451 163 16472 219
rect 16528 163 16549 219
rect 16451 142 16549 163
rect 17699 219 17797 240
rect 17699 163 17720 219
rect 17776 163 17797 219
rect 17699 142 17797 163
rect 18947 219 19045 240
rect 18947 163 18968 219
rect 19024 163 19045 219
rect 18947 142 19045 163
rect 20195 219 20293 240
rect 20195 163 20216 219
rect 20272 163 20293 219
rect 20195 142 20293 163
rect 21443 219 21541 240
rect 21443 163 21464 219
rect 21520 163 21541 219
rect 21443 142 21541 163
rect 22691 219 22789 240
rect 22691 163 22712 219
rect 22768 163 22789 219
rect 22691 142 22789 163
rect 23939 219 24037 240
rect 23939 163 23960 219
rect 24016 163 24037 219
rect 23939 142 24037 163
rect 25187 219 25285 240
rect 25187 163 25208 219
rect 25264 163 25285 219
rect 25187 142 25285 163
rect 26435 219 26533 240
rect 26435 163 26456 219
rect 26512 163 26533 219
rect 26435 142 26533 163
rect 27683 219 27781 240
rect 27683 163 27704 219
rect 27760 163 27781 219
rect 27683 142 27781 163
rect 28931 219 29029 240
rect 28931 163 28952 219
rect 29008 163 29029 219
rect 28931 142 29029 163
rect 30179 219 30277 240
rect 30179 163 30200 219
rect 30256 163 30277 219
rect 30179 142 30277 163
rect 31427 219 31525 240
rect 31427 163 31448 219
rect 31504 163 31525 219
rect 31427 142 31525 163
rect 32675 219 32773 240
rect 32675 163 32696 219
rect 32752 163 32773 219
rect 32675 142 32773 163
rect 33923 219 34021 240
rect 33923 163 33944 219
rect 34000 163 34021 219
rect 33923 142 34021 163
rect 35171 219 35269 240
rect 35171 163 35192 219
rect 35248 163 35269 219
rect 35171 142 35269 163
rect 36419 219 36517 240
rect 36419 163 36440 219
rect 36496 163 36517 219
rect 36419 142 36517 163
rect 37667 219 37765 240
rect 37667 163 37688 219
rect 37744 163 37765 219
rect 37667 142 37765 163
rect 38915 219 39013 240
rect 38915 163 38936 219
rect 38992 163 39013 219
rect 38915 142 39013 163
use contact_14  contact_14_0
timestamp 1701704242
transform 1 0 6591 0 1 778
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1701704242
transform 1 0 6476 0 1 575
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1701704242
transform 1 0 2746 0 1 159
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1701704242
transform 1 0 6490 0 1 159
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1701704242
transform 1 0 2732 0 1 575
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1701704242
transform 1 0 7738 0 1 159
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1701704242
transform 1 0 351 0 1 778
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1701704242
transform 1 0 236 0 1 575
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1701704242
transform 1 0 5343 0 1 778
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1701704242
transform 1 0 250 0 1 159
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1701704242
transform 1 0 3994 0 1 159
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1701704242
transform 1 0 5228 0 1 575
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1701704242
transform 1 0 9087 0 1 778
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1701704242
transform 1 0 1599 0 1 778
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1701704242
transform 1 0 8972 0 1 575
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1701704242
transform 1 0 1498 0 1 159
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1701704242
transform 1 0 5242 0 1 159
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1701704242
transform 1 0 8986 0 1 159
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1701704242
transform 1 0 1484 0 1 575
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1701704242
transform 1 0 2847 0 1 778
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1701704242
transform 1 0 8977 0 1 1546
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1701704242
transform 1 0 8966 0 1 1109
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1701704242
transform 1 0 7729 0 1 1546
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1701704242
transform 1 0 7718 0 1 1109
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1701704242
transform 1 0 6481 0 1 1546
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1701704242
transform 1 0 6470 0 1 1109
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1701704242
transform 1 0 5233 0 1 1546
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1701704242
transform 1 0 5222 0 1 1109
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1701704242
transform 1 0 3985 0 1 1546
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1701704242
transform 1 0 3974 0 1 1109
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1701704242
transform 1 0 2737 0 1 1546
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1701704242
transform 1 0 2726 0 1 1109
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1701704242
transform 1 0 1489 0 1 1546
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1701704242
transform 1 0 1478 0 1 1109
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1701704242
transform 1 0 241 0 1 1546
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1701704242
transform 1 0 230 0 1 1109
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1701704242
transform 1 0 7839 0 1 778
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1701704242
transform 1 0 4095 0 1 778
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1701704242
transform 1 0 7724 0 1 575
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1701704242
transform 1 0 3980 0 1 575
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1701704242
transform 1 0 17722 0 1 159
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1701704242
transform 1 0 16575 0 1 778
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1701704242
transform 1 0 16460 0 1 575
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1701704242
transform 1 0 16474 0 1 159
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1701704242
transform 1 0 18961 0 1 1546
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1701704242
transform 1 0 18950 0 1 1109
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1701704242
transform 1 0 17713 0 1 1546
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1701704242
transform 1 0 17702 0 1 1109
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1701704242
transform 1 0 16465 0 1 1546
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1701704242
transform 1 0 16454 0 1 1109
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1701704242
transform 1 0 15217 0 1 1546
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1701704242
transform 1 0 15206 0 1 1109
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1701704242
transform 1 0 13969 0 1 1546
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1701704242
transform 1 0 13958 0 1 1109
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1701704242
transform 1 0 12721 0 1 1546
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1701704242
transform 1 0 12710 0 1 1109
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1701704242
transform 1 0 11473 0 1 1546
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1701704242
transform 1 0 11462 0 1 1109
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1701704242
transform 1 0 10225 0 1 1546
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1701704242
transform 1 0 10214 0 1 1109
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1701704242
transform 1 0 15327 0 1 778
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1701704242
transform 1 0 15212 0 1 575
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1701704242
transform 1 0 15226 0 1 159
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1701704242
transform 1 0 14079 0 1 778
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1701704242
transform 1 0 13964 0 1 575
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1701704242
transform 1 0 13978 0 1 159
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1701704242
transform 1 0 12831 0 1 778
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1701704242
transform 1 0 12716 0 1 575
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1701704242
transform 1 0 12730 0 1 159
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1701704242
transform 1 0 11583 0 1 778
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1701704242
transform 1 0 11468 0 1 575
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1701704242
transform 1 0 11482 0 1 159
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1701704242
transform 1 0 10335 0 1 778
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1701704242
transform 1 0 10220 0 1 575
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1701704242
transform 1 0 10234 0 1 159
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1701704242
transform 1 0 19071 0 1 778
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1701704242
transform 1 0 18956 0 1 575
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1701704242
transform 1 0 18970 0 1 159
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1701704242
transform 1 0 17823 0 1 778
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1701704242
transform 1 0 17708 0 1 575
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1701704242
transform 1 0 22700 0 1 575
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1701704242
transform 1 0 28954 0 1 159
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1701704242
transform 1 0 22815 0 1 778
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1701704242
transform 1 0 27706 0 1 159
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1701704242
transform 1 0 27807 0 1 778
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1701704242
transform 1 0 20218 0 1 159
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1701704242
transform 1 0 27692 0 1 575
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1701704242
transform 1 0 26449 0 1 1546
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1701704242
transform 1 0 26559 0 1 778
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1701704242
transform 1 0 26438 0 1 1109
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1701704242
transform 1 0 26444 0 1 575
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1701704242
transform 1 0 25201 0 1 1546
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1701704242
transform 1 0 25190 0 1 1109
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1701704242
transform 1 0 22714 0 1 159
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1701704242
transform 1 0 23953 0 1 1546
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1701704242
transform 1 0 26458 0 1 159
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1701704242
transform 1 0 23942 0 1 1109
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1701704242
transform 1 0 22705 0 1 1546
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1701704242
transform 1 0 20319 0 1 778
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1701704242
transform 1 0 22694 0 1 1109
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1701704242
transform 1 0 25311 0 1 778
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1701704242
transform 1 0 21457 0 1 1546
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1701704242
transform 1 0 21446 0 1 1109
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1701704242
transform 1 0 25196 0 1 575
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1701704242
transform 1 0 20209 0 1 1546
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1701704242
transform 1 0 21567 0 1 778
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1701704242
transform 1 0 20198 0 1 1109
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1701704242
transform 1 0 25210 0 1 159
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1701704242
transform 1 0 21452 0 1 575
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1701704242
transform 1 0 24063 0 1 778
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1701704242
transform 1 0 28945 0 1 1546
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1701704242
transform 1 0 23948 0 1 575
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1701704242
transform 1 0 28934 0 1 1109
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1701704242
transform 1 0 27697 0 1 1546
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1701704242
transform 1 0 20204 0 1 575
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1701704242
transform 1 0 27686 0 1 1109
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1701704242
transform 1 0 23962 0 1 159
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1701704242
transform 1 0 29055 0 1 778
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1701704242
transform 1 0 28940 0 1 575
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1701704242
transform 1 0 21466 0 1 159
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1701704242
transform 1 0 39039 0 1 778
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1701704242
transform 1 0 38924 0 1 575
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1701704242
transform 1 0 38938 0 1 159
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1701704242
transform 1 0 37791 0 1 778
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1701704242
transform 1 0 37676 0 1 575
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1701704242
transform 1 0 37690 0 1 159
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1701704242
transform 1 0 36543 0 1 778
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1701704242
transform 1 0 36428 0 1 575
box 0 0 1 1
use contact_14  contact_14_128
timestamp 1701704242
transform 1 0 36442 0 1 159
box 0 0 1 1
use contact_14  contact_14_129
timestamp 1701704242
transform 1 0 35295 0 1 778
box 0 0 1 1
use contact_14  contact_14_130
timestamp 1701704242
transform 1 0 35180 0 1 575
box 0 0 1 1
use contact_14  contact_14_131
timestamp 1701704242
transform 1 0 35194 0 1 159
box 0 0 1 1
use contact_14  contact_14_132
timestamp 1701704242
transform 1 0 34047 0 1 778
box 0 0 1 1
use contact_14  contact_14_133
timestamp 1701704242
transform 1 0 33932 0 1 575
box 0 0 1 1
use contact_14  contact_14_134
timestamp 1701704242
transform 1 0 33946 0 1 159
box 0 0 1 1
use contact_14  contact_14_135
timestamp 1701704242
transform 1 0 32799 0 1 778
box 0 0 1 1
use contact_14  contact_14_136
timestamp 1701704242
transform 1 0 32684 0 1 575
box 0 0 1 1
use contact_14  contact_14_137
timestamp 1701704242
transform 1 0 32698 0 1 159
box 0 0 1 1
use contact_14  contact_14_138
timestamp 1701704242
transform 1 0 31551 0 1 778
box 0 0 1 1
use contact_14  contact_14_139
timestamp 1701704242
transform 1 0 31436 0 1 575
box 0 0 1 1
use contact_14  contact_14_140
timestamp 1701704242
transform 1 0 31450 0 1 159
box 0 0 1 1
use contact_14  contact_14_141
timestamp 1701704242
transform 1 0 30303 0 1 778
box 0 0 1 1
use contact_14  contact_14_142
timestamp 1701704242
transform 1 0 30188 0 1 575
box 0 0 1 1
use contact_14  contact_14_143
timestamp 1701704242
transform 1 0 30202 0 1 159
box 0 0 1 1
use contact_14  contact_14_144
timestamp 1701704242
transform 1 0 38929 0 1 1546
box 0 0 1 1
use contact_14  contact_14_145
timestamp 1701704242
transform 1 0 38918 0 1 1109
box 0 0 1 1
use contact_14  contact_14_146
timestamp 1701704242
transform 1 0 37681 0 1 1546
box 0 0 1 1
use contact_14  contact_14_147
timestamp 1701704242
transform 1 0 37670 0 1 1109
box 0 0 1 1
use contact_14  contact_14_148
timestamp 1701704242
transform 1 0 36433 0 1 1546
box 0 0 1 1
use contact_14  contact_14_149
timestamp 1701704242
transform 1 0 36422 0 1 1109
box 0 0 1 1
use contact_14  contact_14_150
timestamp 1701704242
transform 1 0 35185 0 1 1546
box 0 0 1 1
use contact_14  contact_14_151
timestamp 1701704242
transform 1 0 35174 0 1 1109
box 0 0 1 1
use contact_14  contact_14_152
timestamp 1701704242
transform 1 0 33937 0 1 1546
box 0 0 1 1
use contact_14  contact_14_153
timestamp 1701704242
transform 1 0 33926 0 1 1109
box 0 0 1 1
use contact_14  contact_14_154
timestamp 1701704242
transform 1 0 32689 0 1 1546
box 0 0 1 1
use contact_14  contact_14_155
timestamp 1701704242
transform 1 0 32678 0 1 1109
box 0 0 1 1
use contact_14  contact_14_156
timestamp 1701704242
transform 1 0 31441 0 1 1546
box 0 0 1 1
use contact_14  contact_14_157
timestamp 1701704242
transform 1 0 31430 0 1 1109
box 0 0 1 1
use contact_14  contact_14_158
timestamp 1701704242
transform 1 0 30193 0 1 1546
box 0 0 1 1
use contact_14  contact_14_159
timestamp 1701704242
transform 1 0 30182 0 1 1109
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1701704242
transform 1 0 6584 0 1 772
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1701704242
transform 1 0 6469 0 1 570
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1701704242
transform 1 0 2739 0 1 154
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1701704242
transform 1 0 6483 0 1 154
box 0 0 1 1
use contact_15  contact_15_4
timestamp 1701704242
transform 1 0 2725 0 1 570
box 0 0 1 1
use contact_15  contact_15_5
timestamp 1701704242
transform 1 0 7731 0 1 154
box 0 0 1 1
use contact_15  contact_15_6
timestamp 1701704242
transform 1 0 344 0 1 772
box 0 0 1 1
use contact_15  contact_15_7
timestamp 1701704242
transform 1 0 229 0 1 570
box 0 0 1 1
use contact_15  contact_15_8
timestamp 1701704242
transform 1 0 5336 0 1 772
box 0 0 1 1
use contact_15  contact_15_9
timestamp 1701704242
transform 1 0 243 0 1 154
box 0 0 1 1
use contact_15  contact_15_10
timestamp 1701704242
transform 1 0 3987 0 1 154
box 0 0 1 1
use contact_15  contact_15_11
timestamp 1701704242
transform 1 0 5221 0 1 570
box 0 0 1 1
use contact_15  contact_15_12
timestamp 1701704242
transform 1 0 9080 0 1 772
box 0 0 1 1
use contact_15  contact_15_13
timestamp 1701704242
transform 1 0 1592 0 1 772
box 0 0 1 1
use contact_15  contact_15_14
timestamp 1701704242
transform 1 0 8965 0 1 570
box 0 0 1 1
use contact_15  contact_15_15
timestamp 1701704242
transform 1 0 1491 0 1 154
box 0 0 1 1
use contact_15  contact_15_16
timestamp 1701704242
transform 1 0 5235 0 1 154
box 0 0 1 1
use contact_15  contact_15_17
timestamp 1701704242
transform 1 0 8979 0 1 154
box 0 0 1 1
use contact_15  contact_15_18
timestamp 1701704242
transform 1 0 1477 0 1 570
box 0 0 1 1
use contact_15  contact_15_19
timestamp 1701704242
transform 1 0 2840 0 1 772
box 0 0 1 1
use contact_15  contact_15_20
timestamp 1701704242
transform 1 0 8970 0 1 1541
box 0 0 1 1
use contact_15  contact_15_21
timestamp 1701704242
transform 1 0 8959 0 1 1104
box 0 0 1 1
use contact_15  contact_15_22
timestamp 1701704242
transform 1 0 7722 0 1 1541
box 0 0 1 1
use contact_15  contact_15_23
timestamp 1701704242
transform 1 0 7711 0 1 1104
box 0 0 1 1
use contact_15  contact_15_24
timestamp 1701704242
transform 1 0 6474 0 1 1541
box 0 0 1 1
use contact_15  contact_15_25
timestamp 1701704242
transform 1 0 6463 0 1 1104
box 0 0 1 1
use contact_15  contact_15_26
timestamp 1701704242
transform 1 0 5226 0 1 1541
box 0 0 1 1
use contact_15  contact_15_27
timestamp 1701704242
transform 1 0 5215 0 1 1104
box 0 0 1 1
use contact_15  contact_15_28
timestamp 1701704242
transform 1 0 3978 0 1 1541
box 0 0 1 1
use contact_15  contact_15_29
timestamp 1701704242
transform 1 0 3967 0 1 1104
box 0 0 1 1
use contact_15  contact_15_30
timestamp 1701704242
transform 1 0 2730 0 1 1541
box 0 0 1 1
use contact_15  contact_15_31
timestamp 1701704242
transform 1 0 2719 0 1 1104
box 0 0 1 1
use contact_15  contact_15_32
timestamp 1701704242
transform 1 0 1482 0 1 1541
box 0 0 1 1
use contact_15  contact_15_33
timestamp 1701704242
transform 1 0 1471 0 1 1104
box 0 0 1 1
use contact_15  contact_15_34
timestamp 1701704242
transform 1 0 234 0 1 1541
box 0 0 1 1
use contact_15  contact_15_35
timestamp 1701704242
transform 1 0 223 0 1 1104
box 0 0 1 1
use contact_15  contact_15_36
timestamp 1701704242
transform 1 0 7832 0 1 772
box 0 0 1 1
use contact_15  contact_15_37
timestamp 1701704242
transform 1 0 4088 0 1 772
box 0 0 1 1
use contact_15  contact_15_38
timestamp 1701704242
transform 1 0 7717 0 1 570
box 0 0 1 1
use contact_15  contact_15_39
timestamp 1701704242
transform 1 0 3973 0 1 570
box 0 0 1 1
use contact_15  contact_15_40
timestamp 1701704242
transform 1 0 17715 0 1 154
box 0 0 1 1
use contact_15  contact_15_41
timestamp 1701704242
transform 1 0 16568 0 1 772
box 0 0 1 1
use contact_15  contact_15_42
timestamp 1701704242
transform 1 0 16453 0 1 570
box 0 0 1 1
use contact_15  contact_15_43
timestamp 1701704242
transform 1 0 16467 0 1 154
box 0 0 1 1
use contact_15  contact_15_44
timestamp 1701704242
transform 1 0 18954 0 1 1541
box 0 0 1 1
use contact_15  contact_15_45
timestamp 1701704242
transform 1 0 18943 0 1 1104
box 0 0 1 1
use contact_15  contact_15_46
timestamp 1701704242
transform 1 0 17706 0 1 1541
box 0 0 1 1
use contact_15  contact_15_47
timestamp 1701704242
transform 1 0 17695 0 1 1104
box 0 0 1 1
use contact_15  contact_15_48
timestamp 1701704242
transform 1 0 16458 0 1 1541
box 0 0 1 1
use contact_15  contact_15_49
timestamp 1701704242
transform 1 0 16447 0 1 1104
box 0 0 1 1
use contact_15  contact_15_50
timestamp 1701704242
transform 1 0 15210 0 1 1541
box 0 0 1 1
use contact_15  contact_15_51
timestamp 1701704242
transform 1 0 15199 0 1 1104
box 0 0 1 1
use contact_15  contact_15_52
timestamp 1701704242
transform 1 0 13962 0 1 1541
box 0 0 1 1
use contact_15  contact_15_53
timestamp 1701704242
transform 1 0 13951 0 1 1104
box 0 0 1 1
use contact_15  contact_15_54
timestamp 1701704242
transform 1 0 12714 0 1 1541
box 0 0 1 1
use contact_15  contact_15_55
timestamp 1701704242
transform 1 0 12703 0 1 1104
box 0 0 1 1
use contact_15  contact_15_56
timestamp 1701704242
transform 1 0 11466 0 1 1541
box 0 0 1 1
use contact_15  contact_15_57
timestamp 1701704242
transform 1 0 11455 0 1 1104
box 0 0 1 1
use contact_15  contact_15_58
timestamp 1701704242
transform 1 0 10218 0 1 1541
box 0 0 1 1
use contact_15  contact_15_59
timestamp 1701704242
transform 1 0 10207 0 1 1104
box 0 0 1 1
use contact_15  contact_15_60
timestamp 1701704242
transform 1 0 15320 0 1 772
box 0 0 1 1
use contact_15  contact_15_61
timestamp 1701704242
transform 1 0 15205 0 1 570
box 0 0 1 1
use contact_15  contact_15_62
timestamp 1701704242
transform 1 0 15219 0 1 154
box 0 0 1 1
use contact_15  contact_15_63
timestamp 1701704242
transform 1 0 14072 0 1 772
box 0 0 1 1
use contact_15  contact_15_64
timestamp 1701704242
transform 1 0 13957 0 1 570
box 0 0 1 1
use contact_15  contact_15_65
timestamp 1701704242
transform 1 0 13971 0 1 154
box 0 0 1 1
use contact_15  contact_15_66
timestamp 1701704242
transform 1 0 12824 0 1 772
box 0 0 1 1
use contact_15  contact_15_67
timestamp 1701704242
transform 1 0 12709 0 1 570
box 0 0 1 1
use contact_15  contact_15_68
timestamp 1701704242
transform 1 0 12723 0 1 154
box 0 0 1 1
use contact_15  contact_15_69
timestamp 1701704242
transform 1 0 11576 0 1 772
box 0 0 1 1
use contact_15  contact_15_70
timestamp 1701704242
transform 1 0 11461 0 1 570
box 0 0 1 1
use contact_15  contact_15_71
timestamp 1701704242
transform 1 0 11475 0 1 154
box 0 0 1 1
use contact_15  contact_15_72
timestamp 1701704242
transform 1 0 10328 0 1 772
box 0 0 1 1
use contact_15  contact_15_73
timestamp 1701704242
transform 1 0 10213 0 1 570
box 0 0 1 1
use contact_15  contact_15_74
timestamp 1701704242
transform 1 0 10227 0 1 154
box 0 0 1 1
use contact_15  contact_15_75
timestamp 1701704242
transform 1 0 19064 0 1 772
box 0 0 1 1
use contact_15  contact_15_76
timestamp 1701704242
transform 1 0 18949 0 1 570
box 0 0 1 1
use contact_15  contact_15_77
timestamp 1701704242
transform 1 0 18963 0 1 154
box 0 0 1 1
use contact_15  contact_15_78
timestamp 1701704242
transform 1 0 17816 0 1 772
box 0 0 1 1
use contact_15  contact_15_79
timestamp 1701704242
transform 1 0 17701 0 1 570
box 0 0 1 1
use contact_15  contact_15_80
timestamp 1701704242
transform 1 0 22693 0 1 570
box 0 0 1 1
use contact_15  contact_15_81
timestamp 1701704242
transform 1 0 28947 0 1 154
box 0 0 1 1
use contact_15  contact_15_82
timestamp 1701704242
transform 1 0 22808 0 1 772
box 0 0 1 1
use contact_15  contact_15_83
timestamp 1701704242
transform 1 0 27699 0 1 154
box 0 0 1 1
use contact_15  contact_15_84
timestamp 1701704242
transform 1 0 27800 0 1 772
box 0 0 1 1
use contact_15  contact_15_85
timestamp 1701704242
transform 1 0 20211 0 1 154
box 0 0 1 1
use contact_15  contact_15_86
timestamp 1701704242
transform 1 0 27685 0 1 570
box 0 0 1 1
use contact_15  contact_15_87
timestamp 1701704242
transform 1 0 26442 0 1 1541
box 0 0 1 1
use contact_15  contact_15_88
timestamp 1701704242
transform 1 0 26552 0 1 772
box 0 0 1 1
use contact_15  contact_15_89
timestamp 1701704242
transform 1 0 26431 0 1 1104
box 0 0 1 1
use contact_15  contact_15_90
timestamp 1701704242
transform 1 0 26437 0 1 570
box 0 0 1 1
use contact_15  contact_15_91
timestamp 1701704242
transform 1 0 25194 0 1 1541
box 0 0 1 1
use contact_15  contact_15_92
timestamp 1701704242
transform 1 0 25183 0 1 1104
box 0 0 1 1
use contact_15  contact_15_93
timestamp 1701704242
transform 1 0 22707 0 1 154
box 0 0 1 1
use contact_15  contact_15_94
timestamp 1701704242
transform 1 0 23946 0 1 1541
box 0 0 1 1
use contact_15  contact_15_95
timestamp 1701704242
transform 1 0 26451 0 1 154
box 0 0 1 1
use contact_15  contact_15_96
timestamp 1701704242
transform 1 0 23935 0 1 1104
box 0 0 1 1
use contact_15  contact_15_97
timestamp 1701704242
transform 1 0 22698 0 1 1541
box 0 0 1 1
use contact_15  contact_15_98
timestamp 1701704242
transform 1 0 20312 0 1 772
box 0 0 1 1
use contact_15  contact_15_99
timestamp 1701704242
transform 1 0 22687 0 1 1104
box 0 0 1 1
use contact_15  contact_15_100
timestamp 1701704242
transform 1 0 25304 0 1 772
box 0 0 1 1
use contact_15  contact_15_101
timestamp 1701704242
transform 1 0 21450 0 1 1541
box 0 0 1 1
use contact_15  contact_15_102
timestamp 1701704242
transform 1 0 21439 0 1 1104
box 0 0 1 1
use contact_15  contact_15_103
timestamp 1701704242
transform 1 0 25189 0 1 570
box 0 0 1 1
use contact_15  contact_15_104
timestamp 1701704242
transform 1 0 20202 0 1 1541
box 0 0 1 1
use contact_15  contact_15_105
timestamp 1701704242
transform 1 0 21560 0 1 772
box 0 0 1 1
use contact_15  contact_15_106
timestamp 1701704242
transform 1 0 20191 0 1 1104
box 0 0 1 1
use contact_15  contact_15_107
timestamp 1701704242
transform 1 0 25203 0 1 154
box 0 0 1 1
use contact_15  contact_15_108
timestamp 1701704242
transform 1 0 21445 0 1 570
box 0 0 1 1
use contact_15  contact_15_109
timestamp 1701704242
transform 1 0 24056 0 1 772
box 0 0 1 1
use contact_15  contact_15_110
timestamp 1701704242
transform 1 0 28938 0 1 1541
box 0 0 1 1
use contact_15  contact_15_111
timestamp 1701704242
transform 1 0 23941 0 1 570
box 0 0 1 1
use contact_15  contact_15_112
timestamp 1701704242
transform 1 0 28927 0 1 1104
box 0 0 1 1
use contact_15  contact_15_113
timestamp 1701704242
transform 1 0 27690 0 1 1541
box 0 0 1 1
use contact_15  contact_15_114
timestamp 1701704242
transform 1 0 20197 0 1 570
box 0 0 1 1
use contact_15  contact_15_115
timestamp 1701704242
transform 1 0 27679 0 1 1104
box 0 0 1 1
use contact_15  contact_15_116
timestamp 1701704242
transform 1 0 23955 0 1 154
box 0 0 1 1
use contact_15  contact_15_117
timestamp 1701704242
transform 1 0 29048 0 1 772
box 0 0 1 1
use contact_15  contact_15_118
timestamp 1701704242
transform 1 0 28933 0 1 570
box 0 0 1 1
use contact_15  contact_15_119
timestamp 1701704242
transform 1 0 21459 0 1 154
box 0 0 1 1
use contact_15  contact_15_120
timestamp 1701704242
transform 1 0 39032 0 1 772
box 0 0 1 1
use contact_15  contact_15_121
timestamp 1701704242
transform 1 0 38917 0 1 570
box 0 0 1 1
use contact_15  contact_15_122
timestamp 1701704242
transform 1 0 38931 0 1 154
box 0 0 1 1
use contact_15  contact_15_123
timestamp 1701704242
transform 1 0 37784 0 1 772
box 0 0 1 1
use contact_15  contact_15_124
timestamp 1701704242
transform 1 0 37669 0 1 570
box 0 0 1 1
use contact_15  contact_15_125
timestamp 1701704242
transform 1 0 37683 0 1 154
box 0 0 1 1
use contact_15  contact_15_126
timestamp 1701704242
transform 1 0 36536 0 1 772
box 0 0 1 1
use contact_15  contact_15_127
timestamp 1701704242
transform 1 0 36421 0 1 570
box 0 0 1 1
use contact_15  contact_15_128
timestamp 1701704242
transform 1 0 36435 0 1 154
box 0 0 1 1
use contact_15  contact_15_129
timestamp 1701704242
transform 1 0 35288 0 1 772
box 0 0 1 1
use contact_15  contact_15_130
timestamp 1701704242
transform 1 0 35173 0 1 570
box 0 0 1 1
use contact_15  contact_15_131
timestamp 1701704242
transform 1 0 35187 0 1 154
box 0 0 1 1
use contact_15  contact_15_132
timestamp 1701704242
transform 1 0 34040 0 1 772
box 0 0 1 1
use contact_15  contact_15_133
timestamp 1701704242
transform 1 0 33925 0 1 570
box 0 0 1 1
use contact_15  contact_15_134
timestamp 1701704242
transform 1 0 33939 0 1 154
box 0 0 1 1
use contact_15  contact_15_135
timestamp 1701704242
transform 1 0 32792 0 1 772
box 0 0 1 1
use contact_15  contact_15_136
timestamp 1701704242
transform 1 0 32677 0 1 570
box 0 0 1 1
use contact_15  contact_15_137
timestamp 1701704242
transform 1 0 32691 0 1 154
box 0 0 1 1
use contact_15  contact_15_138
timestamp 1701704242
transform 1 0 31544 0 1 772
box 0 0 1 1
use contact_15  contact_15_139
timestamp 1701704242
transform 1 0 31429 0 1 570
box 0 0 1 1
use contact_15  contact_15_140
timestamp 1701704242
transform 1 0 31443 0 1 154
box 0 0 1 1
use contact_15  contact_15_141
timestamp 1701704242
transform 1 0 30296 0 1 772
box 0 0 1 1
use contact_15  contact_15_142
timestamp 1701704242
transform 1 0 30181 0 1 570
box 0 0 1 1
use contact_15  contact_15_143
timestamp 1701704242
transform 1 0 30195 0 1 154
box 0 0 1 1
use contact_15  contact_15_144
timestamp 1701704242
transform 1 0 38922 0 1 1541
box 0 0 1 1
use contact_15  contact_15_145
timestamp 1701704242
transform 1 0 38911 0 1 1104
box 0 0 1 1
use contact_15  contact_15_146
timestamp 1701704242
transform 1 0 37674 0 1 1541
box 0 0 1 1
use contact_15  contact_15_147
timestamp 1701704242
transform 1 0 37663 0 1 1104
box 0 0 1 1
use contact_15  contact_15_148
timestamp 1701704242
transform 1 0 36426 0 1 1541
box 0 0 1 1
use contact_15  contact_15_149
timestamp 1701704242
transform 1 0 36415 0 1 1104
box 0 0 1 1
use contact_15  contact_15_150
timestamp 1701704242
transform 1 0 35178 0 1 1541
box 0 0 1 1
use contact_15  contact_15_151
timestamp 1701704242
transform 1 0 35167 0 1 1104
box 0 0 1 1
use contact_15  contact_15_152
timestamp 1701704242
transform 1 0 33930 0 1 1541
box 0 0 1 1
use contact_15  contact_15_153
timestamp 1701704242
transform 1 0 33919 0 1 1104
box 0 0 1 1
use contact_15  contact_15_154
timestamp 1701704242
transform 1 0 32682 0 1 1541
box 0 0 1 1
use contact_15  contact_15_155
timestamp 1701704242
transform 1 0 32671 0 1 1104
box 0 0 1 1
use contact_15  contact_15_156
timestamp 1701704242
transform 1 0 31434 0 1 1541
box 0 0 1 1
use contact_15  contact_15_157
timestamp 1701704242
transform 1 0 31423 0 1 1104
box 0 0 1 1
use contact_15  contact_15_158
timestamp 1701704242
transform 1 0 30186 0 1 1541
box 0 0 1 1
use contact_15  contact_15_159
timestamp 1701704242
transform 1 0 30175 0 1 1104
box 0 0 1 1
use write_driver  write_driver_0
timestamp 1701704242
transform 1 0 8736 0 1 0
box -152 4 656 2011
use write_driver  write_driver_1
timestamp 1701704242
transform 1 0 7488 0 1 0
box -152 4 656 2011
use write_driver  write_driver_2
timestamp 1701704242
transform 1 0 6240 0 1 0
box -152 4 656 2011
use write_driver  write_driver_3
timestamp 1701704242
transform 1 0 4992 0 1 0
box -152 4 656 2011
use write_driver  write_driver_4
timestamp 1701704242
transform 1 0 3744 0 1 0
box -152 4 656 2011
use write_driver  write_driver_5
timestamp 1701704242
transform 1 0 2496 0 1 0
box -152 4 656 2011
use write_driver  write_driver_6
timestamp 1701704242
transform 1 0 1248 0 1 0
box -152 4 656 2011
use write_driver  write_driver_7
timestamp 1701704242
transform 1 0 0 0 1 0
box -152 4 656 2011
use write_driver  write_driver_8
timestamp 1701704242
transform 1 0 18720 0 1 0
box -152 4 656 2011
use write_driver  write_driver_9
timestamp 1701704242
transform 1 0 17472 0 1 0
box -152 4 656 2011
use write_driver  write_driver_10
timestamp 1701704242
transform 1 0 16224 0 1 0
box -152 4 656 2011
use write_driver  write_driver_11
timestamp 1701704242
transform 1 0 14976 0 1 0
box -152 4 656 2011
use write_driver  write_driver_12
timestamp 1701704242
transform 1 0 13728 0 1 0
box -152 4 656 2011
use write_driver  write_driver_13
timestamp 1701704242
transform 1 0 12480 0 1 0
box -152 4 656 2011
use write_driver  write_driver_14
timestamp 1701704242
transform 1 0 11232 0 1 0
box -152 4 656 2011
use write_driver  write_driver_15
timestamp 1701704242
transform 1 0 9984 0 1 0
box -152 4 656 2011
use write_driver  write_driver_16
timestamp 1701704242
transform 1 0 28704 0 1 0
box -152 4 656 2011
use write_driver  write_driver_17
timestamp 1701704242
transform 1 0 27456 0 1 0
box -152 4 656 2011
use write_driver  write_driver_18
timestamp 1701704242
transform 1 0 26208 0 1 0
box -152 4 656 2011
use write_driver  write_driver_19
timestamp 1701704242
transform 1 0 24960 0 1 0
box -152 4 656 2011
use write_driver  write_driver_20
timestamp 1701704242
transform 1 0 23712 0 1 0
box -152 4 656 2011
use write_driver  write_driver_21
timestamp 1701704242
transform 1 0 22464 0 1 0
box -152 4 656 2011
use write_driver  write_driver_22
timestamp 1701704242
transform 1 0 21216 0 1 0
box -152 4 656 2011
use write_driver  write_driver_23
timestamp 1701704242
transform 1 0 19968 0 1 0
box -152 4 656 2011
use write_driver  write_driver_24
timestamp 1701704242
transform 1 0 38688 0 1 0
box -152 4 656 2011
use write_driver  write_driver_25
timestamp 1701704242
transform 1 0 37440 0 1 0
box -152 4 656 2011
use write_driver  write_driver_26
timestamp 1701704242
transform 1 0 36192 0 1 0
box -152 4 656 2011
use write_driver  write_driver_27
timestamp 1701704242
transform 1 0 34944 0 1 0
box -152 4 656 2011
use write_driver  write_driver_28
timestamp 1701704242
transform 1 0 33696 0 1 0
box -152 4 656 2011
use write_driver  write_driver_29
timestamp 1701704242
transform 1 0 32448 0 1 0
box -152 4 656 2011
use write_driver  write_driver_30
timestamp 1701704242
transform 1 0 31200 0 1 0
box -152 4 656 2011
use write_driver  write_driver_31
timestamp 1701704242
transform 1 0 29952 0 1 0
box -152 4 656 2011
<< labels >>
rlabel metal1 s 28845 1985 28845 1985 4 bl_23
port 79 nsew
rlabel metal1 s 14071 1985 14071 1985 4 br_11
port 56 nsew
rlabel metal1 s 1591 1985 1591 1985 4 br_1
port 36 nsew
rlabel metal1 s 2637 1985 2637 1985 4 bl_2
port 37 nsew
rlabel metal1 s 15319 1985 15319 1985 4 br_12
port 58 nsew
rlabel metal1 s 21501 32 21501 32 4 data_17
port 18 nsew
rlabel metal1 s 141 1985 141 1985 4 bl_0
port 33 nsew
rlabel metal1 s 29047 1985 29047 1985 4 br_23
port 80 nsew
rlabel metal1 s 17757 32 17757 32 4 data_14
port 15 nsew
rlabel metal1 s 4779 111 4779 111 4 en_0
port 97 nsew
rlabel metal1 s 14763 111 14763 111 4 en_1
port 98 nsew
rlabel metal1 s 19005 32 19005 32 4 data_15
port 16 nsew
rlabel metal1 s 35287 1985 35287 1985 4 br_28
port 90 nsew
rlabel metal1 s 32589 1985 32589 1985 4 bl_26
port 85 nsew
rlabel metal1 s 22749 32 22749 32 4 data_18
port 19 nsew
rlabel metal1 s 5335 1985 5335 1985 4 br_4
port 42 nsew
rlabel metal1 s 36477 32 36477 32 4 data_29
port 30 nsew
rlabel metal1 s 17613 1985 17613 1985 4 bl_14
port 61 nsew
rlabel metal1 s 12621 1985 12621 1985 4 bl_10
port 53 nsew
rlabel metal1 s 20109 1985 20109 1985 4 bl_16
port 65 nsew
rlabel metal1 s 31485 32 31485 32 4 data_25
port 26 nsew
rlabel metal1 s 38829 1985 38829 1985 4 bl_31
port 95 nsew
rlabel metal1 s 37581 1985 37581 1985 4 bl_30
port 93 nsew
rlabel metal1 s 6525 32 6525 32 4 data_5
port 6 nsew
rlabel metal1 s 32733 32 32733 32 4 data_26
port 27 nsew
rlabel metal1 s 3885 1985 3885 1985 4 bl_3
port 39 nsew
rlabel metal1 s 343 1985 343 1985 4 br_0
port 34 nsew
rlabel metal1 s 22605 1985 22605 1985 4 bl_18
port 69 nsew
rlabel metal1 s 15117 1985 15117 1985 4 bl_12
port 57 nsew
rlabel metal1 s 16567 1985 16567 1985 4 br_13
port 60 nsew
rlabel metal1 s 35229 32 35229 32 4 data_28
port 29 nsew
rlabel metal1 s 27799 1985 27799 1985 4 br_22
port 78 nsew
rlabel metal1 s 24747 111 24747 111 4 en_2
port 99 nsew
rlabel metal1 s 33837 1985 33837 1985 4 bl_27
port 87 nsew
rlabel metal1 s 1533 32 1533 32 4 data_1
port 2 nsew
rlabel metal1 s 20311 1985 20311 1985 4 br_16
port 66 nsew
rlabel metal1 s 4087 1985 4087 1985 4 br_3
port 40 nsew
rlabel metal1 s 23853 1985 23853 1985 4 bl_19
port 71 nsew
rlabel metal1 s 9021 32 9021 32 4 data_7
port 8 nsew
rlabel metal1 s 27741 32 27741 32 4 data_22
port 23 nsew
rlabel metal1 s 27597 1985 27597 1985 4 bl_22
port 77 nsew
rlabel metal1 s 21357 1985 21357 1985 4 bl_17
port 67 nsew
rlabel metal1 s 7629 1985 7629 1985 4 bl_6
port 45 nsew
rlabel metal1 s 39031 1985 39031 1985 4 br_31
port 96 nsew
rlabel metal1 s 26349 1985 26349 1985 4 bl_21
port 75 nsew
rlabel metal1 s 285 32 285 32 4 data_0
port 1 nsew
rlabel metal1 s 16509 32 16509 32 4 data_13
port 14 nsew
rlabel metal1 s 34731 111 34731 111 4 en_3
port 100 nsew
rlabel metal1 s 12823 1985 12823 1985 4 br_10
port 54 nsew
rlabel metal1 s 15261 32 15261 32 4 data_12
port 13 nsew
rlabel metal1 s 32791 1985 32791 1985 4 br_26
port 86 nsew
rlabel metal1 s 22807 1985 22807 1985 4 br_18
port 70 nsew
rlabel metal1 s 1389 1985 1389 1985 4 bl_1
port 35 nsew
rlabel metal1 s 36535 1985 36535 1985 4 br_29
port 92 nsew
rlabel metal1 s 28989 32 28989 32 4 data_23
port 24 nsew
rlabel metal1 s 36333 1985 36333 1985 4 bl_29
port 91 nsew
rlabel metal1 s 30093 1985 30093 1985 4 bl_24
port 81 nsew
rlabel metal1 s 12765 32 12765 32 4 data_10
port 11 nsew
rlabel metal1 s 37783 1985 37783 1985 4 br_30
port 94 nsew
rlabel metal1 s 6381 1985 6381 1985 4 bl_5
port 43 nsew
rlabel metal1 s 21559 1985 21559 1985 4 br_17
port 68 nsew
rlabel metal1 s 25101 1985 25101 1985 4 bl_20
port 73 nsew
rlabel metal1 s 8877 1985 8877 1985 4 bl_7
port 47 nsew
rlabel metal1 s 11575 1985 11575 1985 4 br_9
port 52 nsew
rlabel metal1 s 26551 1985 26551 1985 4 br_21
port 76 nsew
rlabel metal1 s 7773 32 7773 32 4 data_6
port 7 nsew
rlabel metal1 s 20253 32 20253 32 4 data_16
port 17 nsew
rlabel metal1 s 11517 32 11517 32 4 data_9
port 10 nsew
rlabel metal1 s 7831 1985 7831 1985 4 br_6
port 46 nsew
rlabel metal1 s 31341 1985 31341 1985 4 bl_25
port 83 nsew
rlabel metal1 s 13869 1985 13869 1985 4 bl_11
port 55 nsew
rlabel metal1 s 25303 1985 25303 1985 4 br_20
port 74 nsew
rlabel metal1 s 5277 32 5277 32 4 data_4
port 5 nsew
rlabel metal1 s 31543 1985 31543 1985 4 br_25
port 84 nsew
rlabel metal1 s 2781 32 2781 32 4 data_2
port 3 nsew
rlabel metal1 s 25245 32 25245 32 4 data_20
port 21 nsew
rlabel metal1 s 38973 32 38973 32 4 data_31
port 32 nsew
rlabel metal1 s 19063 1985 19063 1985 4 br_15
port 64 nsew
rlabel metal1 s 6583 1985 6583 1985 4 br_5
port 44 nsew
rlabel metal1 s 24055 1985 24055 1985 4 br_19
port 72 nsew
rlabel metal1 s 18861 1985 18861 1985 4 bl_15
port 63 nsew
rlabel metal1 s 16365 1985 16365 1985 4 bl_13
port 59 nsew
rlabel metal1 s 34039 1985 34039 1985 4 br_27
port 88 nsew
rlabel metal1 s 10125 1985 10125 1985 4 bl_8
port 49 nsew
rlabel metal1 s 10269 32 10269 32 4 data_8
port 9 nsew
rlabel metal1 s 23997 32 23997 32 4 data_19
port 20 nsew
rlabel metal1 s 2839 1985 2839 1985 4 br_2
port 38 nsew
rlabel metal1 s 9079 1985 9079 1985 4 br_7
port 48 nsew
rlabel metal1 s 10327 1985 10327 1985 4 br_8
port 50 nsew
rlabel metal1 s 30295 1985 30295 1985 4 br_24
port 82 nsew
rlabel metal1 s 11373 1985 11373 1985 4 bl_9
port 51 nsew
rlabel metal1 s 4029 32 4029 32 4 data_3
port 4 nsew
rlabel metal1 s 33981 32 33981 32 4 data_27
port 28 nsew
rlabel metal1 s 35085 1985 35085 1985 4 bl_28
port 89 nsew
rlabel metal1 s 14013 32 14013 32 4 data_11
port 12 nsew
rlabel metal1 s 26493 32 26493 32 4 data_21
port 22 nsew
rlabel metal1 s 37725 32 37725 32 4 data_30
port 31 nsew
rlabel metal1 s 17815 1985 17815 1985 4 br_14
port 62 nsew
rlabel metal1 s 5133 1985 5133 1985 4 bl_4
port 41 nsew
rlabel metal1 s 30237 32 30237 32 4 data_24
port 25 nsew
rlabel metal3 s 21472 1141 21472 1141 4 vdd
port 101 nsew
rlabel metal3 s 22720 1141 22720 1141 4 vdd
port 101 nsew
rlabel metal3 s 28960 1141 28960 1141 4 vdd
port 101 nsew
rlabel metal3 s 36448 1141 36448 1141 4 vdd
port 101 nsew
rlabel metal3 s 35200 1141 35200 1141 4 vdd
port 101 nsew
rlabel metal3 s 30208 1141 30208 1141 4 vdd
port 101 nsew
rlabel metal3 s 37696 1141 37696 1141 4 vdd
port 101 nsew
rlabel metal3 s 33952 1141 33952 1141 4 vdd
port 101 nsew
rlabel metal3 s 26464 1141 26464 1141 4 vdd
port 101 nsew
rlabel metal3 s 25216 1141 25216 1141 4 vdd
port 101 nsew
rlabel metal3 s 38944 1141 38944 1141 4 vdd
port 101 nsew
rlabel metal3 s 31456 1141 31456 1141 4 vdd
port 101 nsew
rlabel metal3 s 23968 1141 23968 1141 4 vdd
port 101 nsew
rlabel metal3 s 32704 1141 32704 1141 4 vdd
port 101 nsew
rlabel metal3 s 20224 1141 20224 1141 4 vdd
port 101 nsew
rlabel metal3 s 27712 1141 27712 1141 4 vdd
port 101 nsew
rlabel metal3 s 21483 1578 21483 1578 4 gnd
port 102 nsew
rlabel metal3 s 30219 1578 30219 1578 4 gnd
port 102 nsew
rlabel metal3 s 27723 1578 27723 1578 4 gnd
port 102 nsew
rlabel metal3 s 32715 1578 32715 1578 4 gnd
port 102 nsew
rlabel metal3 s 28971 1578 28971 1578 4 gnd
port 102 nsew
rlabel metal3 s 23979 1578 23979 1578 4 gnd
port 102 nsew
rlabel metal3 s 33963 1578 33963 1578 4 gnd
port 102 nsew
rlabel metal3 s 20235 1578 20235 1578 4 gnd
port 102 nsew
rlabel metal3 s 22731 1578 22731 1578 4 gnd
port 102 nsew
rlabel metal3 s 25227 1578 25227 1578 4 gnd
port 102 nsew
rlabel metal3 s 31467 1578 31467 1578 4 gnd
port 102 nsew
rlabel metal3 s 38955 1578 38955 1578 4 gnd
port 102 nsew
rlabel metal3 s 26475 1578 26475 1578 4 gnd
port 102 nsew
rlabel metal3 s 35211 1578 35211 1578 4 gnd
port 102 nsew
rlabel metal3 s 36459 1578 36459 1578 4 gnd
port 102 nsew
rlabel metal3 s 37707 1578 37707 1578 4 gnd
port 102 nsew
rlabel metal3 s 27718 607 27718 607 4 gnd
port 102 nsew
rlabel metal3 s 37702 607 37702 607 4 gnd
port 102 nsew
rlabel metal3 s 36454 607 36454 607 4 gnd
port 102 nsew
rlabel metal3 s 35206 607 35206 607 4 gnd
port 102 nsew
rlabel metal3 s 32710 607 32710 607 4 gnd
port 102 nsew
rlabel metal3 s 33958 607 33958 607 4 gnd
port 102 nsew
rlabel metal3 s 28966 607 28966 607 4 gnd
port 102 nsew
rlabel metal3 s 26585 809 26585 809 4 gnd
port 102 nsew
rlabel metal3 s 39065 809 39065 809 4 gnd
port 102 nsew
rlabel metal3 s 37817 809 37817 809 4 gnd
port 102 nsew
rlabel metal3 s 32825 809 32825 809 4 gnd
port 102 nsew
rlabel metal3 s 22841 809 22841 809 4 gnd
port 102 nsew
rlabel metal3 s 36569 809 36569 809 4 gnd
port 102 nsew
rlabel metal3 s 23974 607 23974 607 4 gnd
port 102 nsew
rlabel metal3 s 21593 809 21593 809 4 gnd
port 102 nsew
rlabel metal3 s 34073 809 34073 809 4 gnd
port 102 nsew
rlabel metal3 s 22726 607 22726 607 4 gnd
port 102 nsew
rlabel metal3 s 25337 809 25337 809 4 gnd
port 102 nsew
rlabel metal3 s 30214 607 30214 607 4 gnd
port 102 nsew
rlabel metal3 s 27833 809 27833 809 4 gnd
port 102 nsew
rlabel metal3 s 31462 607 31462 607 4 gnd
port 102 nsew
rlabel metal3 s 24089 809 24089 809 4 gnd
port 102 nsew
rlabel metal3 s 25222 607 25222 607 4 gnd
port 102 nsew
rlabel metal3 s 20345 809 20345 809 4 gnd
port 102 nsew
rlabel metal3 s 26470 607 26470 607 4 gnd
port 102 nsew
rlabel metal3 s 30329 809 30329 809 4 gnd
port 102 nsew
rlabel metal3 s 38950 607 38950 607 4 gnd
port 102 nsew
rlabel metal3 s 31577 809 31577 809 4 gnd
port 102 nsew
rlabel metal3 s 29081 809 29081 809 4 gnd
port 102 nsew
rlabel metal3 s 35321 809 35321 809 4 gnd
port 102 nsew
rlabel metal3 s 20230 607 20230 607 4 gnd
port 102 nsew
rlabel metal3 s 21478 607 21478 607 4 gnd
port 102 nsew
rlabel metal3 s 7750 607 7750 607 4 gnd
port 102 nsew
rlabel metal3 s 1625 809 1625 809 4 gnd
port 102 nsew
rlabel metal3 s 13990 607 13990 607 4 gnd
port 102 nsew
rlabel metal3 s 2758 607 2758 607 4 gnd
port 102 nsew
rlabel metal3 s 8998 607 8998 607 4 gnd
port 102 nsew
rlabel metal3 s 2873 809 2873 809 4 gnd
port 102 nsew
rlabel metal3 s 12742 607 12742 607 4 gnd
port 102 nsew
rlabel metal3 s 377 809 377 809 4 gnd
port 102 nsew
rlabel metal3 s 17734 607 17734 607 4 gnd
port 102 nsew
rlabel metal3 s 14105 809 14105 809 4 gnd
port 102 nsew
rlabel metal3 s 6617 809 6617 809 4 gnd
port 102 nsew
rlabel metal3 s 15238 607 15238 607 4 gnd
port 102 nsew
rlabel metal3 s 18982 607 18982 607 4 gnd
port 102 nsew
rlabel metal3 s 12857 809 12857 809 4 gnd
port 102 nsew
rlabel metal3 s 9113 809 9113 809 4 gnd
port 102 nsew
rlabel metal3 s 10246 607 10246 607 4 gnd
port 102 nsew
rlabel metal3 s 4006 607 4006 607 4 gnd
port 102 nsew
rlabel metal3 s 262 607 262 607 4 gnd
port 102 nsew
rlabel metal3 s 5369 809 5369 809 4 gnd
port 102 nsew
rlabel metal3 s 16601 809 16601 809 4 gnd
port 102 nsew
rlabel metal3 s 7865 809 7865 809 4 gnd
port 102 nsew
rlabel metal3 s 11494 607 11494 607 4 gnd
port 102 nsew
rlabel metal3 s 4121 809 4121 809 4 gnd
port 102 nsew
rlabel metal3 s 6502 607 6502 607 4 gnd
port 102 nsew
rlabel metal3 s 1510 607 1510 607 4 gnd
port 102 nsew
rlabel metal3 s 15353 809 15353 809 4 gnd
port 102 nsew
rlabel metal3 s 11609 809 11609 809 4 gnd
port 102 nsew
rlabel metal3 s 16486 607 16486 607 4 gnd
port 102 nsew
rlabel metal3 s 10361 809 10361 809 4 gnd
port 102 nsew
rlabel metal3 s 17849 809 17849 809 4 gnd
port 102 nsew
rlabel metal3 s 19097 809 19097 809 4 gnd
port 102 nsew
rlabel metal3 s 5254 607 5254 607 4 gnd
port 102 nsew
rlabel metal3 s 267 1578 267 1578 4 gnd
port 102 nsew
rlabel metal3 s 8992 1141 8992 1141 4 vdd
port 101 nsew
rlabel metal3 s 6507 1578 6507 1578 4 gnd
port 102 nsew
rlabel metal3 s 18987 1578 18987 1578 4 gnd
port 102 nsew
rlabel metal3 s 13984 1141 13984 1141 4 vdd
port 101 nsew
rlabel metal3 s 11499 1578 11499 1578 4 gnd
port 102 nsew
rlabel metal3 s 2763 1578 2763 1578 4 gnd
port 102 nsew
rlabel metal3 s 2752 1141 2752 1141 4 vdd
port 101 nsew
rlabel metal3 s 13995 1578 13995 1578 4 gnd
port 102 nsew
rlabel metal3 s 17728 1141 17728 1141 4 vdd
port 101 nsew
rlabel metal3 s 15243 1578 15243 1578 4 gnd
port 102 nsew
rlabel metal3 s 18976 1141 18976 1141 4 vdd
port 101 nsew
rlabel metal3 s 256 1141 256 1141 4 vdd
port 101 nsew
rlabel metal3 s 11488 1141 11488 1141 4 vdd
port 101 nsew
rlabel metal3 s 12736 1141 12736 1141 4 vdd
port 101 nsew
rlabel metal3 s 1515 1578 1515 1578 4 gnd
port 102 nsew
rlabel metal3 s 6496 1141 6496 1141 4 vdd
port 101 nsew
rlabel metal3 s 17739 1578 17739 1578 4 gnd
port 102 nsew
rlabel metal3 s 16491 1578 16491 1578 4 gnd
port 102 nsew
rlabel metal3 s 12747 1578 12747 1578 4 gnd
port 102 nsew
rlabel metal3 s 7744 1141 7744 1141 4 vdd
port 101 nsew
rlabel metal3 s 10251 1578 10251 1578 4 gnd
port 102 nsew
rlabel metal3 s 16480 1141 16480 1141 4 vdd
port 101 nsew
rlabel metal3 s 4000 1141 4000 1141 4 vdd
port 101 nsew
rlabel metal3 s 5248 1141 5248 1141 4 vdd
port 101 nsew
rlabel metal3 s 9003 1578 9003 1578 4 gnd
port 102 nsew
rlabel metal3 s 15232 1141 15232 1141 4 vdd
port 101 nsew
rlabel metal3 s 7755 1578 7755 1578 4 gnd
port 102 nsew
rlabel metal3 s 10240 1141 10240 1141 4 vdd
port 101 nsew
rlabel metal3 s 1504 1141 1504 1141 4 vdd
port 101 nsew
rlabel metal3 s 4011 1578 4011 1578 4 gnd
port 102 nsew
rlabel metal3 s 5259 1578 5259 1578 4 gnd
port 102 nsew
rlabel metal3 s 17748 191 17748 191 4 vdd
port 101 nsew
rlabel metal3 s 14004 191 14004 191 4 vdd
port 101 nsew
rlabel metal3 s 10260 191 10260 191 4 vdd
port 101 nsew
rlabel metal3 s 4020 191 4020 191 4 vdd
port 101 nsew
rlabel metal3 s 11508 191 11508 191 4 vdd
port 101 nsew
rlabel metal3 s 16500 191 16500 191 4 vdd
port 101 nsew
rlabel metal3 s 12756 191 12756 191 4 vdd
port 101 nsew
rlabel metal3 s 276 191 276 191 4 vdd
port 101 nsew
rlabel metal3 s 5268 191 5268 191 4 vdd
port 101 nsew
rlabel metal3 s 7764 191 7764 191 4 vdd
port 101 nsew
rlabel metal3 s 9012 191 9012 191 4 vdd
port 101 nsew
rlabel metal3 s 1524 191 1524 191 4 vdd
port 101 nsew
rlabel metal3 s 2772 191 2772 191 4 vdd
port 101 nsew
rlabel metal3 s 15252 191 15252 191 4 vdd
port 101 nsew
rlabel metal3 s 18996 191 18996 191 4 vdd
port 101 nsew
rlabel metal3 s 6516 191 6516 191 4 vdd
port 101 nsew
rlabel metal3 s 32724 191 32724 191 4 vdd
port 101 nsew
rlabel metal3 s 33972 191 33972 191 4 vdd
port 101 nsew
rlabel metal3 s 22740 191 22740 191 4 vdd
port 101 nsew
rlabel metal3 s 35220 191 35220 191 4 vdd
port 101 nsew
rlabel metal3 s 28980 191 28980 191 4 vdd
port 101 nsew
rlabel metal3 s 38964 191 38964 191 4 vdd
port 101 nsew
rlabel metal3 s 20244 191 20244 191 4 vdd
port 101 nsew
rlabel metal3 s 26484 191 26484 191 4 vdd
port 101 nsew
rlabel metal3 s 23988 191 23988 191 4 vdd
port 101 nsew
rlabel metal3 s 25236 191 25236 191 4 vdd
port 101 nsew
rlabel metal3 s 31476 191 31476 191 4 vdd
port 101 nsew
rlabel metal3 s 27732 191 27732 191 4 vdd
port 101 nsew
rlabel metal3 s 37716 191 37716 191 4 vdd
port 101 nsew
rlabel metal3 s 36468 191 36468 191 4 vdd
port 101 nsew
rlabel metal3 s 21492 191 21492 191 4 vdd
port 101 nsew
rlabel metal3 s 30228 191 30228 191 4 vdd
port 101 nsew
<< properties >>
string FIXED_BBOX 0 0 39936 2011
string GDS_END 3507640
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3453320
<< end >>
