magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -17 25533 15032 27476
<< pwell >>
rect 33 27537 14908 28315
rect 27 25206 8330 25471
rect 12382 25206 14908 25471
rect 27 24622 14908 25206
rect 27 24437 14900 24622
rect 27 19920 287 24437
rect 27 19304 14900 19920
rect 27 18941 11773 19304
rect 14434 18941 14900 19304
rect 27 18595 14900 18941
rect 171 17829 14798 18595
<< mvpsubdiff >>
rect 59 28283 14882 28289
rect 59 28249 121 28283
rect 155 28249 190 28283
rect 224 28249 259 28283
rect 293 28249 328 28283
rect 362 28249 397 28283
rect 431 28249 466 28283
rect 500 28249 535 28283
rect 569 28249 604 28283
rect 638 28249 673 28283
rect 707 28249 742 28283
rect 776 28249 811 28283
rect 845 28249 880 28283
rect 914 28249 949 28283
rect 983 28249 1018 28283
rect 1052 28249 1087 28283
rect 1121 28249 1156 28283
rect 59 28215 1156 28249
rect 59 28181 121 28215
rect 155 28181 190 28215
rect 224 28181 259 28215
rect 293 28181 328 28215
rect 362 28181 397 28215
rect 431 28181 466 28215
rect 500 28181 535 28215
rect 569 28181 604 28215
rect 638 28181 673 28215
rect 707 28181 742 28215
rect 776 28181 811 28215
rect 845 28181 880 28215
rect 914 28181 949 28215
rect 983 28181 1018 28215
rect 1052 28181 1087 28215
rect 1121 28181 1156 28215
rect 59 28147 1156 28181
rect 59 28113 121 28147
rect 155 28113 190 28147
rect 224 28113 259 28147
rect 293 28113 328 28147
rect 362 28113 397 28147
rect 431 28113 466 28147
rect 500 28113 535 28147
rect 569 28113 604 28147
rect 638 28113 673 28147
rect 707 28113 742 28147
rect 776 28113 811 28147
rect 845 28113 880 28147
rect 914 28113 949 28147
rect 983 28113 1018 28147
rect 1052 28113 1087 28147
rect 1121 28113 1156 28147
rect 59 28079 1156 28113
rect 59 28045 121 28079
rect 155 28045 190 28079
rect 224 28045 259 28079
rect 293 28045 328 28079
rect 362 28045 397 28079
rect 431 28045 466 28079
rect 500 28045 535 28079
rect 569 28045 604 28079
rect 638 28045 673 28079
rect 707 28045 742 28079
rect 776 28045 811 28079
rect 845 28045 880 28079
rect 914 28045 949 28079
rect 983 28045 1018 28079
rect 1052 28045 1087 28079
rect 1121 28045 1156 28079
rect 59 28011 1156 28045
rect 59 27977 121 28011
rect 155 27977 190 28011
rect 224 27977 259 28011
rect 293 27977 328 28011
rect 362 27977 397 28011
rect 431 27977 466 28011
rect 500 27977 535 28011
rect 569 27977 604 28011
rect 638 27977 673 28011
rect 707 27977 742 28011
rect 776 27977 811 28011
rect 845 27977 880 28011
rect 914 27977 949 28011
rect 983 27977 1018 28011
rect 1052 27977 1087 28011
rect 1121 27977 1156 28011
rect 59 27943 1156 27977
rect 59 27909 121 27943
rect 155 27909 190 27943
rect 224 27909 259 27943
rect 293 27909 328 27943
rect 362 27909 397 27943
rect 431 27909 466 27943
rect 500 27909 535 27943
rect 569 27909 604 27943
rect 638 27909 673 27943
rect 707 27909 742 27943
rect 776 27909 811 27943
rect 845 27909 880 27943
rect 914 27909 949 27943
rect 983 27909 1018 27943
rect 1052 27909 1087 27943
rect 1121 27909 1156 27943
rect 59 27875 1156 27909
rect 59 27841 121 27875
rect 155 27841 190 27875
rect 224 27841 259 27875
rect 293 27841 328 27875
rect 362 27841 397 27875
rect 431 27841 466 27875
rect 500 27841 535 27875
rect 569 27841 604 27875
rect 638 27841 673 27875
rect 707 27841 742 27875
rect 776 27841 811 27875
rect 845 27841 880 27875
rect 914 27841 949 27875
rect 983 27841 1018 27875
rect 1052 27841 1087 27875
rect 1121 27841 1156 27875
rect 59 27807 1156 27841
rect 59 27773 121 27807
rect 155 27773 190 27807
rect 224 27773 259 27807
rect 293 27773 328 27807
rect 362 27773 397 27807
rect 431 27773 466 27807
rect 500 27773 535 27807
rect 569 27773 604 27807
rect 638 27773 673 27807
rect 707 27773 742 27807
rect 776 27773 811 27807
rect 845 27773 880 27807
rect 914 27773 949 27807
rect 983 27773 1018 27807
rect 1052 27773 1087 27807
rect 1121 27773 1156 27807
rect 59 27739 1156 27773
rect 59 27705 121 27739
rect 155 27705 190 27739
rect 224 27705 259 27739
rect 293 27705 328 27739
rect 362 27705 397 27739
rect 431 27705 466 27739
rect 500 27705 535 27739
rect 569 27705 604 27739
rect 638 27705 673 27739
rect 707 27705 742 27739
rect 776 27705 811 27739
rect 845 27705 880 27739
rect 914 27705 949 27739
rect 983 27705 1018 27739
rect 1052 27705 1087 27739
rect 1121 27705 1156 27739
rect 59 27671 1156 27705
rect 59 27637 121 27671
rect 155 27637 190 27671
rect 224 27637 259 27671
rect 293 27637 328 27671
rect 362 27637 397 27671
rect 431 27637 466 27671
rect 500 27637 535 27671
rect 569 27637 604 27671
rect 638 27637 673 27671
rect 707 27637 742 27671
rect 776 27637 811 27671
rect 845 27637 880 27671
rect 914 27637 949 27671
rect 983 27637 1018 27671
rect 1052 27637 1087 27671
rect 1121 27637 1156 27671
rect 59 27603 1156 27637
rect 59 27569 121 27603
rect 155 27569 190 27603
rect 224 27569 259 27603
rect 293 27569 328 27603
rect 362 27569 397 27603
rect 431 27569 466 27603
rect 500 27569 535 27603
rect 569 27569 604 27603
rect 638 27569 673 27603
rect 707 27569 742 27603
rect 776 27569 811 27603
rect 845 27569 880 27603
rect 914 27569 949 27603
rect 983 27569 1018 27603
rect 1052 27569 1087 27603
rect 1121 27569 1156 27603
rect 14858 27569 14882 28283
rect 59 27563 14882 27569
rect 53 25444 8304 25445
rect 53 25410 77 25444
rect 111 25410 146 25444
rect 180 25410 215 25444
rect 249 25410 284 25444
rect 318 25410 353 25444
rect 387 25410 422 25444
rect 456 25410 491 25444
rect 525 25410 560 25444
rect 594 25410 629 25444
rect 663 25410 698 25444
rect 732 25410 766 25444
rect 800 25410 834 25444
rect 868 25410 902 25444
rect 936 25410 970 25444
rect 1004 25410 1038 25444
rect 1072 25410 1106 25444
rect 1140 25410 1174 25444
rect 1208 25410 1242 25444
rect 1276 25410 1310 25444
rect 1344 25410 1378 25444
rect 1412 25410 1446 25444
rect 1480 25410 1514 25444
rect 1548 25410 1582 25444
rect 1616 25410 1650 25444
rect 1684 25410 1718 25444
rect 1752 25410 1786 25444
rect 1820 25410 1854 25444
rect 1888 25410 1922 25444
rect 1956 25410 1990 25444
rect 2024 25410 2058 25444
rect 2092 25410 2126 25444
rect 2160 25410 2194 25444
rect 2228 25410 2262 25444
rect 2296 25410 2330 25444
rect 2364 25410 2398 25444
rect 2432 25410 2466 25444
rect 2500 25410 2534 25444
rect 2568 25410 2602 25444
rect 2636 25410 2670 25444
rect 2704 25410 2738 25444
rect 2772 25410 2806 25444
rect 2840 25410 2874 25444
rect 2908 25410 2942 25444
rect 2976 25410 3010 25444
rect 3044 25410 3078 25444
rect 3112 25410 3146 25444
rect 3180 25410 3214 25444
rect 3248 25410 3282 25444
rect 3316 25410 3350 25444
rect 3384 25410 3418 25444
rect 3452 25410 3486 25444
rect 3520 25410 3554 25444
rect 3588 25410 3622 25444
rect 3656 25410 3690 25444
rect 3724 25410 3758 25444
rect 3792 25410 3826 25444
rect 3860 25410 3894 25444
rect 3928 25410 3962 25444
rect 3996 25410 4030 25444
rect 4064 25410 4098 25444
rect 4132 25410 4166 25444
rect 4200 25410 4234 25444
rect 4268 25410 4302 25444
rect 4336 25410 4370 25444
rect 4404 25410 4438 25444
rect 4472 25410 4506 25444
rect 4540 25410 4574 25444
rect 4608 25410 4642 25444
rect 4676 25410 4710 25444
rect 4744 25410 4778 25444
rect 4812 25410 4846 25444
rect 4880 25410 4914 25444
rect 4948 25410 4982 25444
rect 5016 25410 5050 25444
rect 5084 25410 5118 25444
rect 5152 25410 5186 25444
rect 5220 25410 5254 25444
rect 5288 25410 5322 25444
rect 5356 25410 5390 25444
rect 5424 25410 5458 25444
rect 5492 25410 5526 25444
rect 5560 25410 5594 25444
rect 5628 25410 5662 25444
rect 5696 25410 5730 25444
rect 5764 25410 5798 25444
rect 5832 25410 5866 25444
rect 5900 25410 5934 25444
rect 5968 25410 6002 25444
rect 6036 25410 6070 25444
rect 6104 25410 6138 25444
rect 6172 25410 6206 25444
rect 6240 25410 6274 25444
rect 6308 25410 6342 25444
rect 6376 25410 6410 25444
rect 6444 25410 6478 25444
rect 6512 25410 6546 25444
rect 6580 25410 6614 25444
rect 6648 25410 6682 25444
rect 6716 25410 6750 25444
rect 6784 25410 6818 25444
rect 6852 25410 6886 25444
rect 6920 25410 6954 25444
rect 6988 25410 7022 25444
rect 7056 25410 7090 25444
rect 7124 25410 7158 25444
rect 7192 25410 7226 25444
rect 7260 25410 7294 25444
rect 7328 25410 7362 25444
rect 7396 25410 7430 25444
rect 7464 25410 7498 25444
rect 7532 25410 7566 25444
rect 7600 25410 7634 25444
rect 7668 25410 7702 25444
rect 7736 25410 7770 25444
rect 7804 25410 7838 25444
rect 7872 25410 7906 25444
rect 7940 25410 7974 25444
rect 8008 25410 8042 25444
rect 8076 25410 8110 25444
rect 8144 25410 8178 25444
rect 8212 25410 8246 25444
rect 8280 25410 8304 25444
rect 53 25358 8304 25410
rect 53 25324 77 25358
rect 111 25324 146 25358
rect 180 25324 215 25358
rect 249 25324 284 25358
rect 318 25324 353 25358
rect 387 25324 422 25358
rect 456 25324 491 25358
rect 525 25324 560 25358
rect 594 25324 629 25358
rect 663 25324 698 25358
rect 732 25324 766 25358
rect 800 25324 834 25358
rect 868 25324 902 25358
rect 936 25324 970 25358
rect 1004 25324 1038 25358
rect 1072 25324 1106 25358
rect 1140 25324 1174 25358
rect 1208 25324 1242 25358
rect 1276 25324 1310 25358
rect 1344 25324 1378 25358
rect 1412 25324 1446 25358
rect 1480 25324 1514 25358
rect 1548 25324 1582 25358
rect 1616 25324 1650 25358
rect 1684 25324 1718 25358
rect 1752 25324 1786 25358
rect 1820 25324 1854 25358
rect 1888 25324 1922 25358
rect 1956 25324 1990 25358
rect 2024 25324 2058 25358
rect 2092 25324 2126 25358
rect 2160 25324 2194 25358
rect 2228 25324 2262 25358
rect 2296 25324 2330 25358
rect 2364 25324 2398 25358
rect 2432 25324 2466 25358
rect 2500 25324 2534 25358
rect 2568 25324 2602 25358
rect 2636 25324 2670 25358
rect 2704 25324 2738 25358
rect 2772 25324 2806 25358
rect 2840 25324 2874 25358
rect 2908 25324 2942 25358
rect 2976 25324 3010 25358
rect 3044 25324 3078 25358
rect 3112 25324 3146 25358
rect 3180 25324 3214 25358
rect 3248 25324 3282 25358
rect 3316 25324 3350 25358
rect 3384 25324 3418 25358
rect 3452 25324 3486 25358
rect 3520 25324 3554 25358
rect 3588 25324 3622 25358
rect 3656 25324 3690 25358
rect 3724 25324 3758 25358
rect 3792 25324 3826 25358
rect 3860 25324 3894 25358
rect 3928 25324 3962 25358
rect 3996 25324 4030 25358
rect 4064 25324 4098 25358
rect 4132 25324 4166 25358
rect 4200 25324 4234 25358
rect 4268 25324 4302 25358
rect 4336 25324 4370 25358
rect 4404 25324 4438 25358
rect 4472 25324 4506 25358
rect 4540 25324 4574 25358
rect 4608 25324 4642 25358
rect 4676 25324 4710 25358
rect 4744 25324 4778 25358
rect 4812 25324 4846 25358
rect 4880 25324 4914 25358
rect 4948 25324 4982 25358
rect 5016 25324 5050 25358
rect 5084 25324 5118 25358
rect 5152 25324 5186 25358
rect 5220 25324 5254 25358
rect 5288 25324 5322 25358
rect 5356 25324 5390 25358
rect 5424 25324 5458 25358
rect 5492 25324 5526 25358
rect 5560 25324 5594 25358
rect 5628 25324 5662 25358
rect 5696 25324 5730 25358
rect 5764 25324 5798 25358
rect 5832 25324 5866 25358
rect 5900 25324 5934 25358
rect 5968 25324 6002 25358
rect 6036 25324 6070 25358
rect 6104 25324 6138 25358
rect 6172 25324 6206 25358
rect 6240 25324 6274 25358
rect 6308 25324 6342 25358
rect 6376 25324 6410 25358
rect 6444 25324 6478 25358
rect 6512 25324 6546 25358
rect 6580 25324 6614 25358
rect 6648 25324 6682 25358
rect 6716 25324 6750 25358
rect 6784 25324 6818 25358
rect 6852 25324 6886 25358
rect 6920 25324 6954 25358
rect 6988 25324 7022 25358
rect 7056 25324 7090 25358
rect 7124 25324 7158 25358
rect 7192 25324 7226 25358
rect 7260 25324 7294 25358
rect 7328 25324 7362 25358
rect 7396 25324 7430 25358
rect 7464 25324 7498 25358
rect 7532 25324 7566 25358
rect 7600 25324 7634 25358
rect 7668 25324 7702 25358
rect 7736 25324 7770 25358
rect 7804 25324 7838 25358
rect 7872 25324 7906 25358
rect 7940 25324 7974 25358
rect 8008 25324 8042 25358
rect 8076 25324 8110 25358
rect 8144 25324 8178 25358
rect 8212 25324 8246 25358
rect 8280 25324 8304 25358
rect 53 25272 8304 25324
rect 53 25238 77 25272
rect 111 25238 146 25272
rect 180 25238 215 25272
rect 249 25238 284 25272
rect 318 25238 353 25272
rect 387 25238 422 25272
rect 456 25238 491 25272
rect 525 25238 560 25272
rect 594 25238 629 25272
rect 663 25238 698 25272
rect 732 25238 766 25272
rect 800 25238 834 25272
rect 868 25238 902 25272
rect 936 25238 970 25272
rect 1004 25238 1038 25272
rect 1072 25238 1106 25272
rect 1140 25238 1174 25272
rect 1208 25238 1242 25272
rect 1276 25238 1310 25272
rect 1344 25238 1378 25272
rect 1412 25238 1446 25272
rect 1480 25238 1514 25272
rect 1548 25238 1582 25272
rect 1616 25238 1650 25272
rect 1684 25238 1718 25272
rect 1752 25238 1786 25272
rect 1820 25238 1854 25272
rect 1888 25238 1922 25272
rect 1956 25238 1990 25272
rect 2024 25238 2058 25272
rect 2092 25238 2126 25272
rect 2160 25238 2194 25272
rect 2228 25238 2262 25272
rect 2296 25238 2330 25272
rect 2364 25238 2398 25272
rect 2432 25238 2466 25272
rect 2500 25238 2534 25272
rect 2568 25238 2602 25272
rect 2636 25238 2670 25272
rect 2704 25238 2738 25272
rect 2772 25238 2806 25272
rect 2840 25238 2874 25272
rect 2908 25238 2942 25272
rect 2976 25238 3010 25272
rect 3044 25238 3078 25272
rect 3112 25238 3146 25272
rect 3180 25238 3214 25272
rect 3248 25238 3282 25272
rect 3316 25238 3350 25272
rect 3384 25238 3418 25272
rect 3452 25238 3486 25272
rect 3520 25238 3554 25272
rect 3588 25238 3622 25272
rect 3656 25238 3690 25272
rect 3724 25238 3758 25272
rect 3792 25238 3826 25272
rect 3860 25238 3894 25272
rect 3928 25238 3962 25272
rect 3996 25238 4030 25272
rect 4064 25238 4098 25272
rect 4132 25238 4166 25272
rect 4200 25238 4234 25272
rect 4268 25238 4302 25272
rect 4336 25238 4370 25272
rect 4404 25238 4438 25272
rect 4472 25238 4506 25272
rect 4540 25238 4574 25272
rect 4608 25238 4642 25272
rect 4676 25238 4710 25272
rect 4744 25238 4778 25272
rect 4812 25238 4846 25272
rect 4880 25238 4914 25272
rect 4948 25238 4982 25272
rect 5016 25238 5050 25272
rect 5084 25238 5118 25272
rect 5152 25238 5186 25272
rect 5220 25238 5254 25272
rect 5288 25238 5322 25272
rect 5356 25238 5390 25272
rect 5424 25238 5458 25272
rect 5492 25238 5526 25272
rect 5560 25238 5594 25272
rect 5628 25238 5662 25272
rect 5696 25238 5730 25272
rect 5764 25238 5798 25272
rect 5832 25238 5866 25272
rect 5900 25238 5934 25272
rect 5968 25238 6002 25272
rect 6036 25238 6070 25272
rect 6104 25238 6138 25272
rect 6172 25238 6206 25272
rect 6240 25238 6274 25272
rect 6308 25238 6342 25272
rect 6376 25238 6410 25272
rect 6444 25238 6478 25272
rect 6512 25238 6546 25272
rect 6580 25238 6614 25272
rect 6648 25238 6682 25272
rect 6716 25238 6750 25272
rect 6784 25238 6818 25272
rect 6852 25238 6886 25272
rect 6920 25238 6954 25272
rect 6988 25238 7022 25272
rect 7056 25238 7090 25272
rect 7124 25238 7158 25272
rect 7192 25238 7226 25272
rect 7260 25238 7294 25272
rect 7328 25238 7362 25272
rect 7396 25238 7430 25272
rect 7464 25238 7498 25272
rect 7532 25238 7566 25272
rect 7600 25238 7634 25272
rect 7668 25238 7702 25272
rect 7736 25238 7770 25272
rect 7804 25238 7838 25272
rect 7872 25238 7906 25272
rect 7940 25238 7974 25272
rect 8008 25238 8042 25272
rect 8076 25238 8110 25272
rect 8144 25238 8178 25272
rect 8212 25238 8246 25272
rect 8280 25238 8304 25272
rect 53 25180 8304 25238
rect 12408 25444 14882 25445
rect 12408 25410 12432 25444
rect 12466 25410 12501 25444
rect 12535 25410 12570 25444
rect 12604 25410 12639 25444
rect 12673 25410 12708 25444
rect 12742 25410 12777 25444
rect 12811 25410 12846 25444
rect 12880 25410 12915 25444
rect 12949 25410 12984 25444
rect 13018 25410 13053 25444
rect 13087 25410 13122 25444
rect 13156 25410 13191 25444
rect 13225 25410 13260 25444
rect 13294 25410 13328 25444
rect 13362 25410 13396 25444
rect 13430 25410 13464 25444
rect 13498 25410 13532 25444
rect 13566 25410 13600 25444
rect 13634 25410 13668 25444
rect 13702 25410 13736 25444
rect 13770 25410 13804 25444
rect 13838 25410 13872 25444
rect 13906 25410 13940 25444
rect 13974 25410 14008 25444
rect 14042 25410 14076 25444
rect 14110 25410 14144 25444
rect 14178 25410 14212 25444
rect 14246 25410 14280 25444
rect 14314 25410 14348 25444
rect 14382 25410 14416 25444
rect 14450 25410 14484 25444
rect 14518 25410 14552 25444
rect 14586 25410 14620 25444
rect 14654 25410 14688 25444
rect 14722 25410 14756 25444
rect 14790 25410 14824 25444
rect 14858 25410 14882 25444
rect 12408 25358 14882 25410
rect 12408 25324 12432 25358
rect 12466 25324 12501 25358
rect 12535 25324 12570 25358
rect 12604 25324 12639 25358
rect 12673 25324 12708 25358
rect 12742 25324 12777 25358
rect 12811 25324 12846 25358
rect 12880 25324 12915 25358
rect 12949 25324 12984 25358
rect 13018 25324 13053 25358
rect 13087 25324 13122 25358
rect 13156 25324 13191 25358
rect 13225 25324 13260 25358
rect 13294 25324 13328 25358
rect 13362 25324 13396 25358
rect 13430 25324 13464 25358
rect 13498 25324 13532 25358
rect 13566 25324 13600 25358
rect 13634 25324 13668 25358
rect 13702 25324 13736 25358
rect 13770 25324 13804 25358
rect 13838 25324 13872 25358
rect 13906 25324 13940 25358
rect 13974 25324 14008 25358
rect 14042 25324 14076 25358
rect 14110 25324 14144 25358
rect 14178 25324 14212 25358
rect 14246 25324 14280 25358
rect 14314 25324 14348 25358
rect 14382 25324 14416 25358
rect 14450 25324 14484 25358
rect 14518 25324 14552 25358
rect 14586 25324 14620 25358
rect 14654 25324 14688 25358
rect 14722 25324 14756 25358
rect 14790 25324 14824 25358
rect 14858 25324 14882 25358
rect 12408 25272 14882 25324
rect 12408 25238 12432 25272
rect 12466 25238 12501 25272
rect 12535 25238 12570 25272
rect 12604 25238 12639 25272
rect 12673 25238 12708 25272
rect 12742 25238 12777 25272
rect 12811 25238 12846 25272
rect 12880 25238 12915 25272
rect 12949 25238 12984 25272
rect 13018 25238 13053 25272
rect 13087 25238 13122 25272
rect 13156 25238 13191 25272
rect 13225 25238 13260 25272
rect 13294 25238 13328 25272
rect 13362 25238 13396 25272
rect 13430 25238 13464 25272
rect 13498 25238 13532 25272
rect 13566 25238 13600 25272
rect 13634 25238 13668 25272
rect 13702 25238 13736 25272
rect 13770 25238 13804 25272
rect 13838 25238 13872 25272
rect 13906 25238 13940 25272
rect 13974 25238 14008 25272
rect 14042 25238 14076 25272
rect 14110 25238 14144 25272
rect 14178 25238 14212 25272
rect 14246 25238 14280 25272
rect 14314 25238 14348 25272
rect 14382 25238 14416 25272
rect 14450 25238 14484 25272
rect 14518 25238 14552 25272
rect 14586 25238 14620 25272
rect 14654 25238 14688 25272
rect 14722 25238 14756 25272
rect 14790 25238 14824 25272
rect 14858 25238 14882 25272
rect 12408 25180 14882 25238
rect 53 25178 14882 25180
rect 53 25144 124 25178
rect 158 25144 193 25178
rect 227 25144 262 25178
rect 296 25144 331 25178
rect 365 25144 400 25178
rect 434 25144 469 25178
rect 503 25144 538 25178
rect 572 25144 607 25178
rect 641 25144 676 25178
rect 710 25144 745 25178
rect 779 25144 814 25178
rect 848 25144 883 25178
rect 917 25144 952 25178
rect 986 25144 1020 25178
rect 1054 25144 1088 25178
rect 1122 25144 1156 25178
rect 1190 25144 1224 25178
rect 1258 25144 1292 25178
rect 1326 25144 1360 25178
rect 1394 25144 1428 25178
rect 1462 25144 1496 25178
rect 1530 25144 1564 25178
rect 1598 25144 1632 25178
rect 1666 25144 1700 25178
rect 1734 25144 1768 25178
rect 1802 25144 1836 25178
rect 1870 25144 1904 25178
rect 1938 25144 1972 25178
rect 2006 25144 2040 25178
rect 2074 25144 2108 25178
rect 2142 25144 2176 25178
rect 2210 25144 2244 25178
rect 2278 25144 2312 25178
rect 2346 25144 2380 25178
rect 2414 25144 2448 25178
rect 2482 25144 2516 25178
rect 2550 25144 2584 25178
rect 2618 25144 2652 25178
rect 2686 25144 2720 25178
rect 2754 25144 2788 25178
rect 2822 25144 2856 25178
rect 2890 25144 2924 25178
rect 2958 25144 2992 25178
rect 3026 25144 3060 25178
rect 3094 25144 3128 25178
rect 3162 25144 3196 25178
rect 3230 25144 3264 25178
rect 3298 25144 3332 25178
rect 3366 25144 3400 25178
rect 3434 25144 3468 25178
rect 3502 25144 3536 25178
rect 3570 25144 3604 25178
rect 3638 25144 3672 25178
rect 3706 25144 3740 25178
rect 3774 25144 3808 25178
rect 3842 25144 3876 25178
rect 3910 25144 3944 25178
rect 3978 25144 4012 25178
rect 4046 25144 4080 25178
rect 4114 25144 4148 25178
rect 4182 25144 4216 25178
rect 4250 25144 4284 25178
rect 4318 25144 4352 25178
rect 4386 25144 4420 25178
rect 4454 25144 4488 25178
rect 4522 25144 4556 25178
rect 4590 25144 4624 25178
rect 4658 25144 4692 25178
rect 4726 25144 4760 25178
rect 4794 25144 4828 25178
rect 4862 25144 4896 25178
rect 4930 25144 4964 25178
rect 4998 25144 5032 25178
rect 5066 25144 5100 25178
rect 5134 25144 5168 25178
rect 5202 25144 5236 25178
rect 5270 25144 5304 25178
rect 5338 25144 5372 25178
rect 5406 25144 5440 25178
rect 5474 25144 5508 25178
rect 5542 25144 5576 25178
rect 5610 25144 5644 25178
rect 5678 25144 5712 25178
rect 5746 25144 5780 25178
rect 5814 25144 5848 25178
rect 5882 25144 5916 25178
rect 5950 25144 5984 25178
rect 6018 25144 6052 25178
rect 6086 25144 6120 25178
rect 6154 25144 6188 25178
rect 6222 25144 6256 25178
rect 6290 25144 6324 25178
rect 6358 25144 6392 25178
rect 6426 25144 6460 25178
rect 6494 25144 6528 25178
rect 6562 25144 6596 25178
rect 6630 25144 6664 25178
rect 6698 25144 6732 25178
rect 6766 25144 6800 25178
rect 6834 25144 6868 25178
rect 6902 25144 6936 25178
rect 6970 25144 7004 25178
rect 7038 25144 7072 25178
rect 7106 25144 7140 25178
rect 7174 25144 7208 25178
rect 7242 25144 7276 25178
rect 7310 25144 7344 25178
rect 7378 25144 7412 25178
rect 7446 25144 7480 25178
rect 7514 25144 7548 25178
rect 7582 25144 7616 25178
rect 7650 25144 7684 25178
rect 7718 25144 7752 25178
rect 7786 25144 7820 25178
rect 7854 25144 7888 25178
rect 7922 25144 7956 25178
rect 7990 25144 8024 25178
rect 8058 25144 8092 25178
rect 8126 25144 8160 25178
rect 8194 25144 8228 25178
rect 8262 25144 8296 25178
rect 8330 25144 8364 25178
rect 8398 25144 8432 25178
rect 8466 25144 8500 25178
rect 8534 25144 8568 25178
rect 8602 25144 8636 25178
rect 8670 25144 8704 25178
rect 8738 25144 8772 25178
rect 8806 25144 8840 25178
rect 8874 25144 8908 25178
rect 8942 25144 8976 25178
rect 9010 25144 9044 25178
rect 9078 25144 9112 25178
rect 9146 25144 9180 25178
rect 9214 25144 9248 25178
rect 9282 25144 9316 25178
rect 9350 25144 9384 25178
rect 9418 25144 9452 25178
rect 9486 25144 9520 25178
rect 9554 25144 9588 25178
rect 9622 25144 9656 25178
rect 9690 25144 9724 25178
rect 9758 25144 9792 25178
rect 9826 25144 9860 25178
rect 9894 25144 9928 25178
rect 9962 25144 9996 25178
rect 10030 25144 10064 25178
rect 10098 25144 10132 25178
rect 10166 25144 10200 25178
rect 10234 25144 10268 25178
rect 10302 25144 10336 25178
rect 10370 25144 10404 25178
rect 10438 25144 10472 25178
rect 10506 25144 10540 25178
rect 10574 25144 10608 25178
rect 10642 25144 10676 25178
rect 10710 25144 10744 25178
rect 10778 25144 10812 25178
rect 10846 25144 10880 25178
rect 10914 25144 10948 25178
rect 10982 25144 11016 25178
rect 11050 25144 11084 25178
rect 11118 25144 11152 25178
rect 11186 25144 11220 25178
rect 11254 25144 11288 25178
rect 11322 25144 11356 25178
rect 11390 25144 11424 25178
rect 11458 25144 11492 25178
rect 11526 25144 11560 25178
rect 11594 25144 11628 25178
rect 11662 25144 11696 25178
rect 11730 25144 11764 25178
rect 11798 25144 11832 25178
rect 11866 25144 11900 25178
rect 11934 25144 11968 25178
rect 12002 25144 12036 25178
rect 12070 25144 12104 25178
rect 12138 25144 12172 25178
rect 12206 25144 12240 25178
rect 12274 25144 12308 25178
rect 12342 25144 12376 25178
rect 12410 25144 12444 25178
rect 12478 25144 12512 25178
rect 12546 25144 12580 25178
rect 12614 25144 12648 25178
rect 12682 25144 12716 25178
rect 12750 25144 12784 25178
rect 12818 25144 12852 25178
rect 12886 25144 12920 25178
rect 12954 25144 12988 25178
rect 13022 25144 13056 25178
rect 13090 25144 13124 25178
rect 13158 25144 13192 25178
rect 13226 25144 13260 25178
rect 13294 25144 13328 25178
rect 13362 25144 13396 25178
rect 13430 25144 13464 25178
rect 13498 25144 13532 25178
rect 13566 25144 13600 25178
rect 13634 25144 13668 25178
rect 13702 25144 13736 25178
rect 13770 25144 13804 25178
rect 13838 25144 13872 25178
rect 13906 25144 13940 25178
rect 13974 25144 14008 25178
rect 14042 25144 14076 25178
rect 14110 25144 14144 25178
rect 14178 25144 14212 25178
rect 14246 25144 14280 25178
rect 14314 25144 14348 25178
rect 14382 25144 14416 25178
rect 14450 25144 14484 25178
rect 14518 25144 14552 25178
rect 14586 25144 14620 25178
rect 14654 25144 14688 25178
rect 14722 25144 14756 25178
rect 14790 25144 14824 25178
rect 14858 25144 14882 25178
rect 53 25106 14882 25144
rect 53 25072 124 25106
rect 158 25072 193 25106
rect 227 25072 262 25106
rect 296 25072 331 25106
rect 365 25072 400 25106
rect 434 25072 469 25106
rect 503 25072 538 25106
rect 572 25072 607 25106
rect 641 25072 676 25106
rect 710 25072 745 25106
rect 779 25072 814 25106
rect 848 25072 883 25106
rect 917 25072 952 25106
rect 986 25072 1020 25106
rect 1054 25072 1088 25106
rect 1122 25072 1156 25106
rect 1190 25072 1224 25106
rect 1258 25072 1292 25106
rect 1326 25072 1360 25106
rect 1394 25072 1428 25106
rect 1462 25072 1496 25106
rect 1530 25072 1564 25106
rect 1598 25072 1632 25106
rect 1666 25072 1700 25106
rect 1734 25072 1768 25106
rect 1802 25072 1836 25106
rect 1870 25072 1904 25106
rect 1938 25072 1972 25106
rect 2006 25072 2040 25106
rect 2074 25072 2108 25106
rect 2142 25072 2176 25106
rect 2210 25072 2244 25106
rect 2278 25072 2312 25106
rect 2346 25072 2380 25106
rect 2414 25072 2448 25106
rect 2482 25072 2516 25106
rect 2550 25072 2584 25106
rect 2618 25072 2652 25106
rect 2686 25072 2720 25106
rect 2754 25072 2788 25106
rect 2822 25072 2856 25106
rect 2890 25072 2924 25106
rect 2958 25072 2992 25106
rect 3026 25072 3060 25106
rect 3094 25072 3128 25106
rect 3162 25072 3196 25106
rect 3230 25072 3264 25106
rect 3298 25072 3332 25106
rect 3366 25072 3400 25106
rect 3434 25072 3468 25106
rect 3502 25072 3536 25106
rect 3570 25072 3604 25106
rect 3638 25072 3672 25106
rect 3706 25072 3740 25106
rect 3774 25072 3808 25106
rect 3842 25072 3876 25106
rect 3910 25072 3944 25106
rect 3978 25072 4012 25106
rect 4046 25072 4080 25106
rect 4114 25072 4148 25106
rect 4182 25072 4216 25106
rect 4250 25072 4284 25106
rect 4318 25072 4352 25106
rect 4386 25072 4420 25106
rect 4454 25072 4488 25106
rect 4522 25072 4556 25106
rect 4590 25072 4624 25106
rect 4658 25072 4692 25106
rect 4726 25072 4760 25106
rect 4794 25072 4828 25106
rect 4862 25072 4896 25106
rect 4930 25072 4964 25106
rect 4998 25072 5032 25106
rect 5066 25072 5100 25106
rect 5134 25072 5168 25106
rect 5202 25072 5236 25106
rect 5270 25072 5304 25106
rect 5338 25072 5372 25106
rect 5406 25072 5440 25106
rect 5474 25072 5508 25106
rect 5542 25072 5576 25106
rect 5610 25072 5644 25106
rect 5678 25072 5712 25106
rect 5746 25072 5780 25106
rect 5814 25072 5848 25106
rect 5882 25072 5916 25106
rect 5950 25072 5984 25106
rect 6018 25072 6052 25106
rect 6086 25072 6120 25106
rect 6154 25072 6188 25106
rect 6222 25072 6256 25106
rect 6290 25072 6324 25106
rect 6358 25072 6392 25106
rect 6426 25072 6460 25106
rect 6494 25072 6528 25106
rect 6562 25072 6596 25106
rect 6630 25072 6664 25106
rect 6698 25072 6732 25106
rect 6766 25072 6800 25106
rect 6834 25072 6868 25106
rect 6902 25072 6936 25106
rect 6970 25072 7004 25106
rect 7038 25072 7072 25106
rect 7106 25072 7140 25106
rect 7174 25072 7208 25106
rect 7242 25072 7276 25106
rect 7310 25072 7344 25106
rect 7378 25072 7412 25106
rect 7446 25072 7480 25106
rect 7514 25072 7548 25106
rect 7582 25072 7616 25106
rect 7650 25072 7684 25106
rect 7718 25072 7752 25106
rect 7786 25072 7820 25106
rect 7854 25072 7888 25106
rect 7922 25072 7956 25106
rect 7990 25072 8024 25106
rect 8058 25072 8092 25106
rect 8126 25072 8160 25106
rect 8194 25072 8228 25106
rect 8262 25072 8296 25106
rect 8330 25072 8364 25106
rect 8398 25072 8432 25106
rect 8466 25072 8500 25106
rect 8534 25072 8568 25106
rect 8602 25072 8636 25106
rect 8670 25072 8704 25106
rect 8738 25072 8772 25106
rect 8806 25072 8840 25106
rect 8874 25072 8908 25106
rect 8942 25072 8976 25106
rect 9010 25072 9044 25106
rect 9078 25072 9112 25106
rect 9146 25072 9180 25106
rect 9214 25072 9248 25106
rect 9282 25072 9316 25106
rect 9350 25072 9384 25106
rect 9418 25072 9452 25106
rect 9486 25072 9520 25106
rect 9554 25072 9588 25106
rect 9622 25072 9656 25106
rect 9690 25072 9724 25106
rect 9758 25072 9792 25106
rect 9826 25072 9860 25106
rect 9894 25072 9928 25106
rect 9962 25072 9996 25106
rect 10030 25072 10064 25106
rect 10098 25072 10132 25106
rect 10166 25072 10200 25106
rect 10234 25072 10268 25106
rect 10302 25072 10336 25106
rect 10370 25072 10404 25106
rect 10438 25072 10472 25106
rect 10506 25072 10540 25106
rect 10574 25072 10608 25106
rect 10642 25072 10676 25106
rect 10710 25072 10744 25106
rect 10778 25072 10812 25106
rect 10846 25072 10880 25106
rect 10914 25072 10948 25106
rect 10982 25072 11016 25106
rect 11050 25072 11084 25106
rect 11118 25072 11152 25106
rect 11186 25072 11220 25106
rect 11254 25072 11288 25106
rect 11322 25072 11356 25106
rect 11390 25072 11424 25106
rect 11458 25072 11492 25106
rect 11526 25072 11560 25106
rect 11594 25072 11628 25106
rect 11662 25072 11696 25106
rect 11730 25072 11764 25106
rect 11798 25072 11832 25106
rect 11866 25072 11900 25106
rect 11934 25072 11968 25106
rect 12002 25072 12036 25106
rect 12070 25072 12104 25106
rect 12138 25072 12172 25106
rect 12206 25072 12240 25106
rect 12274 25072 12308 25106
rect 12342 25072 12376 25106
rect 12410 25072 12444 25106
rect 12478 25072 12512 25106
rect 12546 25072 12580 25106
rect 12614 25072 12648 25106
rect 12682 25072 12716 25106
rect 12750 25072 12784 25106
rect 12818 25072 12852 25106
rect 12886 25072 12920 25106
rect 12954 25072 12988 25106
rect 13022 25072 13056 25106
rect 13090 25072 13124 25106
rect 13158 25072 13192 25106
rect 13226 25072 13260 25106
rect 13294 25072 13328 25106
rect 13362 25072 13396 25106
rect 13430 25072 13464 25106
rect 13498 25072 13532 25106
rect 13566 25072 13600 25106
rect 13634 25072 13668 25106
rect 13702 25072 13736 25106
rect 13770 25072 13804 25106
rect 13838 25072 13872 25106
rect 13906 25072 13940 25106
rect 13974 25072 14008 25106
rect 14042 25072 14076 25106
rect 14110 25072 14144 25106
rect 14178 25072 14212 25106
rect 14246 25072 14280 25106
rect 14314 25072 14348 25106
rect 14382 25072 14416 25106
rect 14450 25072 14484 25106
rect 14518 25072 14552 25106
rect 14586 25072 14620 25106
rect 14654 25072 14688 25106
rect 14722 25072 14756 25106
rect 14790 25072 14824 25106
rect 14858 25072 14882 25106
rect 53 25034 14882 25072
rect 53 25000 124 25034
rect 158 25000 193 25034
rect 227 25000 262 25034
rect 296 25000 331 25034
rect 365 25000 400 25034
rect 434 25000 469 25034
rect 503 25000 538 25034
rect 572 25000 607 25034
rect 641 25000 676 25034
rect 710 25000 745 25034
rect 779 25000 814 25034
rect 848 25000 883 25034
rect 917 25000 952 25034
rect 986 25000 1020 25034
rect 1054 25000 1088 25034
rect 1122 25000 1156 25034
rect 1190 25000 1224 25034
rect 1258 25000 1292 25034
rect 1326 25000 1360 25034
rect 1394 25000 1428 25034
rect 1462 25000 1496 25034
rect 1530 25000 1564 25034
rect 1598 25000 1632 25034
rect 1666 25000 1700 25034
rect 1734 25000 1768 25034
rect 1802 25000 1836 25034
rect 1870 25000 1904 25034
rect 1938 25000 1972 25034
rect 2006 25000 2040 25034
rect 2074 25000 2108 25034
rect 2142 25000 2176 25034
rect 2210 25000 2244 25034
rect 2278 25000 2312 25034
rect 2346 25000 2380 25034
rect 2414 25000 2448 25034
rect 2482 25000 2516 25034
rect 2550 25000 2584 25034
rect 2618 25000 2652 25034
rect 2686 25000 2720 25034
rect 2754 25000 2788 25034
rect 2822 25000 2856 25034
rect 2890 25000 2924 25034
rect 2958 25000 2992 25034
rect 3026 25000 3060 25034
rect 3094 25000 3128 25034
rect 3162 25000 3196 25034
rect 3230 25000 3264 25034
rect 3298 25000 3332 25034
rect 3366 25000 3400 25034
rect 3434 25000 3468 25034
rect 3502 25000 3536 25034
rect 3570 25000 3604 25034
rect 3638 25000 3672 25034
rect 3706 25000 3740 25034
rect 3774 25000 3808 25034
rect 3842 25000 3876 25034
rect 3910 25000 3944 25034
rect 3978 25000 4012 25034
rect 4046 25000 4080 25034
rect 4114 25000 4148 25034
rect 4182 25000 4216 25034
rect 4250 25000 4284 25034
rect 4318 25000 4352 25034
rect 4386 25000 4420 25034
rect 4454 25000 4488 25034
rect 4522 25000 4556 25034
rect 4590 25000 4624 25034
rect 4658 25000 4692 25034
rect 4726 25000 4760 25034
rect 4794 25000 4828 25034
rect 4862 25000 4896 25034
rect 4930 25000 4964 25034
rect 4998 25000 5032 25034
rect 5066 25000 5100 25034
rect 5134 25000 5168 25034
rect 5202 25000 5236 25034
rect 5270 25000 5304 25034
rect 5338 25000 5372 25034
rect 5406 25000 5440 25034
rect 5474 25000 5508 25034
rect 5542 25000 5576 25034
rect 5610 25000 5644 25034
rect 5678 25000 5712 25034
rect 5746 25000 5780 25034
rect 5814 25000 5848 25034
rect 5882 25000 5916 25034
rect 5950 25000 5984 25034
rect 6018 25000 6052 25034
rect 6086 25000 6120 25034
rect 6154 25000 6188 25034
rect 6222 25000 6256 25034
rect 6290 25000 6324 25034
rect 6358 25000 6392 25034
rect 6426 25000 6460 25034
rect 6494 25000 6528 25034
rect 6562 25000 6596 25034
rect 6630 25000 6664 25034
rect 6698 25000 6732 25034
rect 6766 25000 6800 25034
rect 6834 25000 6868 25034
rect 6902 25000 6936 25034
rect 6970 25000 7004 25034
rect 7038 25000 7072 25034
rect 7106 25000 7140 25034
rect 7174 25000 7208 25034
rect 7242 25000 7276 25034
rect 7310 25000 7344 25034
rect 7378 25000 7412 25034
rect 7446 25000 7480 25034
rect 7514 25000 7548 25034
rect 7582 25000 7616 25034
rect 7650 25000 7684 25034
rect 7718 25000 7752 25034
rect 7786 25000 7820 25034
rect 7854 25000 7888 25034
rect 7922 25000 7956 25034
rect 7990 25000 8024 25034
rect 8058 25000 8092 25034
rect 8126 25000 8160 25034
rect 8194 25000 8228 25034
rect 8262 25000 8296 25034
rect 8330 25000 8364 25034
rect 8398 25000 8432 25034
rect 8466 25000 8500 25034
rect 8534 25000 8568 25034
rect 8602 25000 8636 25034
rect 8670 25000 8704 25034
rect 8738 25000 8772 25034
rect 8806 25000 8840 25034
rect 8874 25000 8908 25034
rect 8942 25000 8976 25034
rect 9010 25000 9044 25034
rect 9078 25000 9112 25034
rect 9146 25000 9180 25034
rect 9214 25000 9248 25034
rect 9282 25000 9316 25034
rect 9350 25000 9384 25034
rect 9418 25000 9452 25034
rect 9486 25000 9520 25034
rect 9554 25000 9588 25034
rect 9622 25000 9656 25034
rect 9690 25000 9724 25034
rect 9758 25000 9792 25034
rect 9826 25000 9860 25034
rect 9894 25000 9928 25034
rect 9962 25000 9996 25034
rect 10030 25000 10064 25034
rect 10098 25000 10132 25034
rect 10166 25000 10200 25034
rect 10234 25000 10268 25034
rect 10302 25000 10336 25034
rect 10370 25000 10404 25034
rect 10438 25000 10472 25034
rect 10506 25000 10540 25034
rect 10574 25000 10608 25034
rect 10642 25000 10676 25034
rect 10710 25000 10744 25034
rect 10778 25000 10812 25034
rect 10846 25000 10880 25034
rect 10914 25000 10948 25034
rect 10982 25000 11016 25034
rect 11050 25000 11084 25034
rect 11118 25000 11152 25034
rect 11186 25000 11220 25034
rect 11254 25000 11288 25034
rect 11322 25000 11356 25034
rect 11390 25000 11424 25034
rect 11458 25000 11492 25034
rect 11526 25000 11560 25034
rect 11594 25000 11628 25034
rect 11662 25000 11696 25034
rect 11730 25000 11764 25034
rect 11798 25000 11832 25034
rect 11866 25000 11900 25034
rect 11934 25000 11968 25034
rect 12002 25000 12036 25034
rect 12070 25000 12104 25034
rect 12138 25000 12172 25034
rect 12206 25000 12240 25034
rect 12274 25000 12308 25034
rect 12342 25000 12376 25034
rect 12410 25000 12444 25034
rect 12478 25000 12512 25034
rect 12546 25000 12580 25034
rect 12614 25000 12648 25034
rect 12682 25000 12716 25034
rect 12750 25000 12784 25034
rect 12818 25000 12852 25034
rect 12886 25000 12920 25034
rect 12954 25000 12988 25034
rect 13022 25000 13056 25034
rect 13090 25000 13124 25034
rect 13158 25000 13192 25034
rect 13226 25000 13260 25034
rect 13294 25000 13328 25034
rect 13362 25000 13396 25034
rect 13430 25000 13464 25034
rect 13498 25000 13532 25034
rect 13566 25000 13600 25034
rect 13634 25000 13668 25034
rect 13702 25000 13736 25034
rect 13770 25000 13804 25034
rect 13838 25000 13872 25034
rect 13906 25000 13940 25034
rect 13974 25000 14008 25034
rect 14042 25000 14076 25034
rect 14110 25000 14144 25034
rect 14178 25000 14212 25034
rect 14246 25000 14280 25034
rect 14314 25000 14348 25034
rect 14382 25000 14416 25034
rect 14450 25000 14484 25034
rect 14518 25000 14552 25034
rect 14586 25000 14620 25034
rect 14654 25000 14688 25034
rect 14722 25000 14756 25034
rect 14790 25000 14824 25034
rect 14858 25000 14882 25034
rect 53 24962 14882 25000
rect 53 24928 124 24962
rect 158 24928 193 24962
rect 227 24928 262 24962
rect 296 24928 331 24962
rect 365 24928 400 24962
rect 434 24928 469 24962
rect 503 24928 538 24962
rect 572 24928 607 24962
rect 641 24928 676 24962
rect 710 24928 745 24962
rect 779 24928 814 24962
rect 848 24928 883 24962
rect 917 24928 952 24962
rect 986 24928 1020 24962
rect 1054 24928 1088 24962
rect 1122 24928 1156 24962
rect 1190 24928 1224 24962
rect 1258 24928 1292 24962
rect 1326 24928 1360 24962
rect 1394 24928 1428 24962
rect 1462 24928 1496 24962
rect 1530 24928 1564 24962
rect 1598 24928 1632 24962
rect 1666 24928 1700 24962
rect 1734 24928 1768 24962
rect 1802 24928 1836 24962
rect 1870 24928 1904 24962
rect 1938 24928 1972 24962
rect 2006 24928 2040 24962
rect 2074 24928 2108 24962
rect 2142 24928 2176 24962
rect 2210 24928 2244 24962
rect 2278 24928 2312 24962
rect 2346 24928 2380 24962
rect 2414 24928 2448 24962
rect 2482 24928 2516 24962
rect 2550 24928 2584 24962
rect 2618 24928 2652 24962
rect 2686 24928 2720 24962
rect 2754 24928 2788 24962
rect 2822 24928 2856 24962
rect 2890 24928 2924 24962
rect 2958 24928 2992 24962
rect 3026 24928 3060 24962
rect 3094 24928 3128 24962
rect 3162 24928 3196 24962
rect 3230 24928 3264 24962
rect 3298 24928 3332 24962
rect 3366 24928 3400 24962
rect 3434 24928 3468 24962
rect 3502 24928 3536 24962
rect 3570 24928 3604 24962
rect 3638 24928 3672 24962
rect 3706 24928 3740 24962
rect 3774 24928 3808 24962
rect 3842 24928 3876 24962
rect 3910 24928 3944 24962
rect 3978 24928 4012 24962
rect 4046 24928 4080 24962
rect 4114 24928 4148 24962
rect 4182 24928 4216 24962
rect 4250 24928 4284 24962
rect 4318 24928 4352 24962
rect 4386 24928 4420 24962
rect 4454 24928 4488 24962
rect 4522 24928 4556 24962
rect 4590 24928 4624 24962
rect 4658 24928 4692 24962
rect 4726 24928 4760 24962
rect 4794 24928 4828 24962
rect 4862 24928 4896 24962
rect 4930 24928 4964 24962
rect 4998 24928 5032 24962
rect 5066 24928 5100 24962
rect 5134 24928 5168 24962
rect 5202 24928 5236 24962
rect 5270 24928 5304 24962
rect 5338 24928 5372 24962
rect 5406 24928 5440 24962
rect 5474 24928 5508 24962
rect 5542 24928 5576 24962
rect 5610 24928 5644 24962
rect 5678 24928 5712 24962
rect 5746 24928 5780 24962
rect 5814 24928 5848 24962
rect 5882 24928 5916 24962
rect 5950 24928 5984 24962
rect 6018 24928 6052 24962
rect 6086 24928 6120 24962
rect 6154 24928 6188 24962
rect 6222 24928 6256 24962
rect 6290 24928 6324 24962
rect 6358 24928 6392 24962
rect 6426 24928 6460 24962
rect 6494 24928 6528 24962
rect 6562 24928 6596 24962
rect 6630 24928 6664 24962
rect 6698 24928 6732 24962
rect 6766 24928 6800 24962
rect 6834 24928 6868 24962
rect 6902 24928 6936 24962
rect 6970 24928 7004 24962
rect 7038 24928 7072 24962
rect 7106 24928 7140 24962
rect 7174 24928 7208 24962
rect 7242 24928 7276 24962
rect 7310 24928 7344 24962
rect 7378 24928 7412 24962
rect 7446 24928 7480 24962
rect 7514 24928 7548 24962
rect 7582 24928 7616 24962
rect 7650 24928 7684 24962
rect 7718 24928 7752 24962
rect 7786 24928 7820 24962
rect 7854 24928 7888 24962
rect 7922 24928 7956 24962
rect 7990 24928 8024 24962
rect 8058 24928 8092 24962
rect 8126 24928 8160 24962
rect 8194 24928 8228 24962
rect 8262 24928 8296 24962
rect 8330 24928 8364 24962
rect 8398 24928 8432 24962
rect 8466 24928 8500 24962
rect 8534 24928 8568 24962
rect 8602 24928 8636 24962
rect 8670 24928 8704 24962
rect 8738 24928 8772 24962
rect 8806 24928 8840 24962
rect 8874 24928 8908 24962
rect 8942 24928 8976 24962
rect 9010 24928 9044 24962
rect 9078 24928 9112 24962
rect 9146 24928 9180 24962
rect 9214 24928 9248 24962
rect 9282 24928 9316 24962
rect 9350 24928 9384 24962
rect 9418 24928 9452 24962
rect 9486 24928 9520 24962
rect 9554 24928 9588 24962
rect 9622 24928 9656 24962
rect 9690 24928 9724 24962
rect 9758 24928 9792 24962
rect 9826 24928 9860 24962
rect 9894 24928 9928 24962
rect 9962 24928 9996 24962
rect 10030 24928 10064 24962
rect 10098 24928 10132 24962
rect 10166 24928 10200 24962
rect 10234 24928 10268 24962
rect 10302 24928 10336 24962
rect 10370 24928 10404 24962
rect 10438 24928 10472 24962
rect 10506 24928 10540 24962
rect 10574 24928 10608 24962
rect 10642 24928 10676 24962
rect 10710 24928 10744 24962
rect 10778 24928 10812 24962
rect 10846 24928 10880 24962
rect 10914 24928 10948 24962
rect 10982 24928 11016 24962
rect 11050 24928 11084 24962
rect 11118 24928 11152 24962
rect 11186 24928 11220 24962
rect 11254 24928 11288 24962
rect 11322 24928 11356 24962
rect 11390 24928 11424 24962
rect 11458 24928 11492 24962
rect 11526 24928 11560 24962
rect 11594 24928 11628 24962
rect 11662 24928 11696 24962
rect 11730 24928 11764 24962
rect 11798 24928 11832 24962
rect 11866 24928 11900 24962
rect 11934 24928 11968 24962
rect 12002 24928 12036 24962
rect 12070 24928 12104 24962
rect 12138 24928 12172 24962
rect 12206 24928 12240 24962
rect 12274 24928 12308 24962
rect 12342 24928 12376 24962
rect 12410 24928 12444 24962
rect 12478 24928 12512 24962
rect 12546 24928 12580 24962
rect 12614 24928 12648 24962
rect 12682 24928 12716 24962
rect 12750 24928 12784 24962
rect 12818 24928 12852 24962
rect 12886 24928 12920 24962
rect 12954 24928 12988 24962
rect 13022 24928 13056 24962
rect 13090 24928 13124 24962
rect 13158 24928 13192 24962
rect 13226 24928 13260 24962
rect 13294 24928 13328 24962
rect 13362 24928 13396 24962
rect 13430 24928 13464 24962
rect 13498 24928 13532 24962
rect 13566 24928 13600 24962
rect 13634 24928 13668 24962
rect 13702 24928 13736 24962
rect 13770 24928 13804 24962
rect 13838 24928 13872 24962
rect 13906 24928 13940 24962
rect 13974 24928 14008 24962
rect 14042 24928 14076 24962
rect 14110 24928 14144 24962
rect 14178 24928 14212 24962
rect 14246 24928 14280 24962
rect 14314 24928 14348 24962
rect 14382 24928 14416 24962
rect 14450 24928 14484 24962
rect 14518 24928 14552 24962
rect 14586 24928 14620 24962
rect 14654 24928 14688 24962
rect 14722 24928 14756 24962
rect 14790 24928 14824 24962
rect 14858 24928 14882 24962
rect 53 24890 14882 24928
rect 53 24856 124 24890
rect 158 24856 193 24890
rect 227 24856 262 24890
rect 296 24856 331 24890
rect 365 24856 400 24890
rect 434 24856 469 24890
rect 503 24856 538 24890
rect 572 24856 607 24890
rect 641 24856 676 24890
rect 710 24856 745 24890
rect 779 24856 814 24890
rect 848 24856 883 24890
rect 917 24856 952 24890
rect 986 24856 1020 24890
rect 1054 24856 1088 24890
rect 1122 24856 1156 24890
rect 1190 24856 1224 24890
rect 1258 24856 1292 24890
rect 1326 24856 1360 24890
rect 1394 24856 1428 24890
rect 1462 24856 1496 24890
rect 1530 24856 1564 24890
rect 1598 24856 1632 24890
rect 1666 24856 1700 24890
rect 1734 24856 1768 24890
rect 1802 24856 1836 24890
rect 1870 24856 1904 24890
rect 1938 24856 1972 24890
rect 2006 24856 2040 24890
rect 2074 24856 2108 24890
rect 2142 24856 2176 24890
rect 2210 24856 2244 24890
rect 2278 24856 2312 24890
rect 2346 24856 2380 24890
rect 2414 24856 2448 24890
rect 2482 24856 2516 24890
rect 2550 24856 2584 24890
rect 2618 24856 2652 24890
rect 2686 24856 2720 24890
rect 2754 24856 2788 24890
rect 2822 24856 2856 24890
rect 2890 24856 2924 24890
rect 2958 24856 2992 24890
rect 3026 24856 3060 24890
rect 3094 24856 3128 24890
rect 3162 24856 3196 24890
rect 3230 24856 3264 24890
rect 3298 24856 3332 24890
rect 3366 24856 3400 24890
rect 3434 24856 3468 24890
rect 3502 24856 3536 24890
rect 3570 24856 3604 24890
rect 3638 24856 3672 24890
rect 3706 24856 3740 24890
rect 3774 24856 3808 24890
rect 3842 24856 3876 24890
rect 3910 24856 3944 24890
rect 3978 24856 4012 24890
rect 4046 24856 4080 24890
rect 4114 24856 4148 24890
rect 4182 24856 4216 24890
rect 4250 24856 4284 24890
rect 4318 24856 4352 24890
rect 4386 24856 4420 24890
rect 4454 24856 4488 24890
rect 4522 24856 4556 24890
rect 4590 24856 4624 24890
rect 4658 24856 4692 24890
rect 4726 24856 4760 24890
rect 4794 24856 4828 24890
rect 4862 24856 4896 24890
rect 4930 24856 4964 24890
rect 4998 24856 5032 24890
rect 5066 24856 5100 24890
rect 5134 24856 5168 24890
rect 5202 24856 5236 24890
rect 5270 24856 5304 24890
rect 5338 24856 5372 24890
rect 5406 24856 5440 24890
rect 5474 24856 5508 24890
rect 5542 24856 5576 24890
rect 5610 24856 5644 24890
rect 5678 24856 5712 24890
rect 5746 24856 5780 24890
rect 5814 24856 5848 24890
rect 5882 24856 5916 24890
rect 5950 24856 5984 24890
rect 6018 24856 6052 24890
rect 6086 24856 6120 24890
rect 6154 24856 6188 24890
rect 6222 24856 6256 24890
rect 6290 24856 6324 24890
rect 6358 24856 6392 24890
rect 6426 24856 6460 24890
rect 6494 24856 6528 24890
rect 6562 24856 6596 24890
rect 6630 24856 6664 24890
rect 6698 24856 6732 24890
rect 6766 24856 6800 24890
rect 6834 24856 6868 24890
rect 6902 24856 6936 24890
rect 6970 24856 7004 24890
rect 7038 24856 7072 24890
rect 7106 24856 7140 24890
rect 7174 24856 7208 24890
rect 7242 24856 7276 24890
rect 7310 24856 7344 24890
rect 7378 24856 7412 24890
rect 7446 24856 7480 24890
rect 7514 24856 7548 24890
rect 7582 24856 7616 24890
rect 7650 24856 7684 24890
rect 7718 24856 7752 24890
rect 7786 24856 7820 24890
rect 7854 24856 7888 24890
rect 7922 24856 7956 24890
rect 7990 24856 8024 24890
rect 8058 24856 8092 24890
rect 8126 24856 8160 24890
rect 8194 24856 8228 24890
rect 8262 24856 8296 24890
rect 8330 24856 8364 24890
rect 8398 24856 8432 24890
rect 8466 24856 8500 24890
rect 8534 24856 8568 24890
rect 8602 24856 8636 24890
rect 8670 24856 8704 24890
rect 8738 24856 8772 24890
rect 8806 24856 8840 24890
rect 8874 24856 8908 24890
rect 8942 24856 8976 24890
rect 9010 24856 9044 24890
rect 9078 24856 9112 24890
rect 9146 24856 9180 24890
rect 9214 24856 9248 24890
rect 9282 24856 9316 24890
rect 9350 24856 9384 24890
rect 9418 24856 9452 24890
rect 9486 24856 9520 24890
rect 9554 24856 9588 24890
rect 9622 24856 9656 24890
rect 9690 24856 9724 24890
rect 9758 24856 9792 24890
rect 9826 24856 9860 24890
rect 9894 24856 9928 24890
rect 9962 24856 9996 24890
rect 10030 24856 10064 24890
rect 10098 24856 10132 24890
rect 10166 24856 10200 24890
rect 10234 24856 10268 24890
rect 10302 24856 10336 24890
rect 10370 24856 10404 24890
rect 10438 24856 10472 24890
rect 10506 24856 10540 24890
rect 10574 24856 10608 24890
rect 10642 24856 10676 24890
rect 10710 24856 10744 24890
rect 10778 24856 10812 24890
rect 10846 24856 10880 24890
rect 10914 24856 10948 24890
rect 10982 24856 11016 24890
rect 11050 24856 11084 24890
rect 11118 24856 11152 24890
rect 11186 24856 11220 24890
rect 11254 24856 11288 24890
rect 11322 24856 11356 24890
rect 11390 24856 11424 24890
rect 11458 24856 11492 24890
rect 11526 24856 11560 24890
rect 11594 24856 11628 24890
rect 11662 24856 11696 24890
rect 11730 24856 11764 24890
rect 11798 24856 11832 24890
rect 11866 24856 11900 24890
rect 11934 24856 11968 24890
rect 12002 24856 12036 24890
rect 12070 24856 12104 24890
rect 12138 24856 12172 24890
rect 12206 24856 12240 24890
rect 12274 24856 12308 24890
rect 12342 24856 12376 24890
rect 12410 24856 12444 24890
rect 12478 24856 12512 24890
rect 12546 24856 12580 24890
rect 12614 24856 12648 24890
rect 12682 24856 12716 24890
rect 12750 24856 12784 24890
rect 12818 24856 12852 24890
rect 12886 24856 12920 24890
rect 12954 24856 12988 24890
rect 13022 24856 13056 24890
rect 13090 24856 13124 24890
rect 13158 24856 13192 24890
rect 13226 24856 13260 24890
rect 13294 24856 13328 24890
rect 13362 24856 13396 24890
rect 13430 24856 13464 24890
rect 13498 24856 13532 24890
rect 13566 24856 13600 24890
rect 13634 24856 13668 24890
rect 13702 24856 13736 24890
rect 13770 24856 13804 24890
rect 13838 24856 13872 24890
rect 13906 24856 13940 24890
rect 13974 24856 14008 24890
rect 14042 24856 14076 24890
rect 14110 24856 14144 24890
rect 14178 24856 14212 24890
rect 14246 24856 14280 24890
rect 14314 24856 14348 24890
rect 14382 24856 14416 24890
rect 14450 24856 14484 24890
rect 14518 24856 14552 24890
rect 14586 24856 14620 24890
rect 14654 24856 14688 24890
rect 14722 24856 14756 24890
rect 14790 24856 14824 24890
rect 14858 24856 14882 24890
rect 53 24818 14882 24856
rect 53 24784 124 24818
rect 158 24784 193 24818
rect 227 24784 262 24818
rect 296 24784 331 24818
rect 365 24784 400 24818
rect 434 24784 469 24818
rect 503 24784 538 24818
rect 572 24784 607 24818
rect 641 24784 676 24818
rect 710 24784 745 24818
rect 779 24784 814 24818
rect 848 24784 883 24818
rect 917 24784 952 24818
rect 986 24784 1020 24818
rect 1054 24784 1088 24818
rect 1122 24784 1156 24818
rect 1190 24784 1224 24818
rect 1258 24784 1292 24818
rect 1326 24784 1360 24818
rect 1394 24784 1428 24818
rect 1462 24784 1496 24818
rect 1530 24784 1564 24818
rect 1598 24784 1632 24818
rect 1666 24784 1700 24818
rect 1734 24784 1768 24818
rect 1802 24784 1836 24818
rect 1870 24784 1904 24818
rect 1938 24784 1972 24818
rect 2006 24784 2040 24818
rect 2074 24784 2108 24818
rect 2142 24784 2176 24818
rect 2210 24784 2244 24818
rect 2278 24784 2312 24818
rect 2346 24784 2380 24818
rect 2414 24784 2448 24818
rect 2482 24784 2516 24818
rect 2550 24784 2584 24818
rect 2618 24784 2652 24818
rect 2686 24784 2720 24818
rect 2754 24784 2788 24818
rect 2822 24784 2856 24818
rect 2890 24784 2924 24818
rect 2958 24784 2992 24818
rect 3026 24784 3060 24818
rect 3094 24784 3128 24818
rect 3162 24784 3196 24818
rect 3230 24784 3264 24818
rect 3298 24784 3332 24818
rect 3366 24784 3400 24818
rect 3434 24784 3468 24818
rect 3502 24784 3536 24818
rect 3570 24784 3604 24818
rect 3638 24784 3672 24818
rect 3706 24784 3740 24818
rect 3774 24784 3808 24818
rect 3842 24784 3876 24818
rect 3910 24784 3944 24818
rect 3978 24784 4012 24818
rect 4046 24784 4080 24818
rect 4114 24784 4148 24818
rect 4182 24784 4216 24818
rect 4250 24784 4284 24818
rect 4318 24784 4352 24818
rect 4386 24784 4420 24818
rect 4454 24784 4488 24818
rect 4522 24784 4556 24818
rect 4590 24784 4624 24818
rect 4658 24784 4692 24818
rect 4726 24784 4760 24818
rect 4794 24784 4828 24818
rect 4862 24784 4896 24818
rect 4930 24784 4964 24818
rect 4998 24784 5032 24818
rect 5066 24784 5100 24818
rect 5134 24784 5168 24818
rect 5202 24784 5236 24818
rect 5270 24784 5304 24818
rect 5338 24784 5372 24818
rect 5406 24784 5440 24818
rect 5474 24784 5508 24818
rect 5542 24784 5576 24818
rect 5610 24784 5644 24818
rect 5678 24784 5712 24818
rect 5746 24784 5780 24818
rect 5814 24784 5848 24818
rect 5882 24784 5916 24818
rect 5950 24784 5984 24818
rect 6018 24784 6052 24818
rect 6086 24784 6120 24818
rect 6154 24784 6188 24818
rect 6222 24784 6256 24818
rect 6290 24784 6324 24818
rect 6358 24784 6392 24818
rect 6426 24784 6460 24818
rect 6494 24784 6528 24818
rect 6562 24784 6596 24818
rect 6630 24784 6664 24818
rect 6698 24784 6732 24818
rect 6766 24784 6800 24818
rect 6834 24784 6868 24818
rect 6902 24784 6936 24818
rect 6970 24784 7004 24818
rect 7038 24784 7072 24818
rect 7106 24784 7140 24818
rect 7174 24784 7208 24818
rect 7242 24784 7276 24818
rect 7310 24784 7344 24818
rect 7378 24784 7412 24818
rect 7446 24784 7480 24818
rect 7514 24784 7548 24818
rect 7582 24784 7616 24818
rect 7650 24784 7684 24818
rect 7718 24784 7752 24818
rect 7786 24784 7820 24818
rect 7854 24784 7888 24818
rect 7922 24784 7956 24818
rect 7990 24784 8024 24818
rect 8058 24784 8092 24818
rect 8126 24784 8160 24818
rect 8194 24784 8228 24818
rect 8262 24784 8296 24818
rect 8330 24784 8364 24818
rect 8398 24784 8432 24818
rect 8466 24784 8500 24818
rect 8534 24784 8568 24818
rect 8602 24784 8636 24818
rect 8670 24784 8704 24818
rect 8738 24784 8772 24818
rect 8806 24784 8840 24818
rect 8874 24784 8908 24818
rect 8942 24784 8976 24818
rect 9010 24784 9044 24818
rect 9078 24784 9112 24818
rect 9146 24784 9180 24818
rect 9214 24784 9248 24818
rect 9282 24784 9316 24818
rect 9350 24784 9384 24818
rect 9418 24784 9452 24818
rect 9486 24784 9520 24818
rect 9554 24784 9588 24818
rect 9622 24784 9656 24818
rect 9690 24784 9724 24818
rect 9758 24784 9792 24818
rect 9826 24784 9860 24818
rect 9894 24784 9928 24818
rect 9962 24784 9996 24818
rect 10030 24784 10064 24818
rect 10098 24784 10132 24818
rect 10166 24784 10200 24818
rect 10234 24784 10268 24818
rect 10302 24784 10336 24818
rect 10370 24784 10404 24818
rect 10438 24784 10472 24818
rect 10506 24784 10540 24818
rect 10574 24784 10608 24818
rect 10642 24784 10676 24818
rect 10710 24784 10744 24818
rect 10778 24784 10812 24818
rect 10846 24784 10880 24818
rect 10914 24784 10948 24818
rect 10982 24784 11016 24818
rect 11050 24784 11084 24818
rect 11118 24784 11152 24818
rect 11186 24784 11220 24818
rect 11254 24784 11288 24818
rect 11322 24784 11356 24818
rect 11390 24784 11424 24818
rect 11458 24784 11492 24818
rect 11526 24784 11560 24818
rect 11594 24784 11628 24818
rect 11662 24784 11696 24818
rect 11730 24784 11764 24818
rect 11798 24784 11832 24818
rect 11866 24784 11900 24818
rect 11934 24784 11968 24818
rect 12002 24784 12036 24818
rect 12070 24784 12104 24818
rect 12138 24784 12172 24818
rect 12206 24784 12240 24818
rect 12274 24784 12308 24818
rect 12342 24784 12376 24818
rect 12410 24784 12444 24818
rect 12478 24784 12512 24818
rect 12546 24784 12580 24818
rect 12614 24784 12648 24818
rect 12682 24784 12716 24818
rect 12750 24784 12784 24818
rect 12818 24784 12852 24818
rect 12886 24784 12920 24818
rect 12954 24784 12988 24818
rect 13022 24784 13056 24818
rect 13090 24784 13124 24818
rect 13158 24784 13192 24818
rect 13226 24784 13260 24818
rect 13294 24784 13328 24818
rect 13362 24784 13396 24818
rect 13430 24784 13464 24818
rect 13498 24784 13532 24818
rect 13566 24784 13600 24818
rect 13634 24784 13668 24818
rect 13702 24784 13736 24818
rect 13770 24784 13804 24818
rect 13838 24784 13872 24818
rect 13906 24784 13940 24818
rect 13974 24784 14008 24818
rect 14042 24784 14076 24818
rect 14110 24784 14144 24818
rect 14178 24784 14212 24818
rect 14246 24784 14280 24818
rect 14314 24784 14348 24818
rect 14382 24784 14416 24818
rect 14450 24784 14484 24818
rect 14518 24784 14552 24818
rect 14586 24784 14620 24818
rect 14654 24784 14688 24818
rect 14722 24784 14756 24818
rect 14790 24784 14824 24818
rect 14858 24784 14882 24818
rect 53 24746 14882 24784
rect 53 24712 124 24746
rect 158 24712 193 24746
rect 227 24712 262 24746
rect 296 24712 331 24746
rect 365 24712 400 24746
rect 434 24712 469 24746
rect 503 24712 538 24746
rect 572 24712 607 24746
rect 641 24712 676 24746
rect 710 24712 745 24746
rect 779 24712 814 24746
rect 848 24712 883 24746
rect 917 24712 952 24746
rect 986 24712 1020 24746
rect 1054 24712 1088 24746
rect 1122 24712 1156 24746
rect 1190 24712 1224 24746
rect 1258 24712 1292 24746
rect 1326 24712 1360 24746
rect 1394 24712 1428 24746
rect 1462 24712 1496 24746
rect 1530 24712 1564 24746
rect 1598 24712 1632 24746
rect 1666 24712 1700 24746
rect 1734 24712 1768 24746
rect 1802 24712 1836 24746
rect 1870 24712 1904 24746
rect 1938 24712 1972 24746
rect 2006 24712 2040 24746
rect 2074 24712 2108 24746
rect 2142 24712 2176 24746
rect 2210 24712 2244 24746
rect 2278 24712 2312 24746
rect 2346 24712 2380 24746
rect 2414 24712 2448 24746
rect 2482 24712 2516 24746
rect 2550 24712 2584 24746
rect 2618 24712 2652 24746
rect 2686 24712 2720 24746
rect 2754 24712 2788 24746
rect 2822 24712 2856 24746
rect 2890 24712 2924 24746
rect 2958 24712 2992 24746
rect 3026 24712 3060 24746
rect 3094 24712 3128 24746
rect 3162 24712 3196 24746
rect 3230 24712 3264 24746
rect 3298 24712 3332 24746
rect 3366 24712 3400 24746
rect 3434 24712 3468 24746
rect 3502 24712 3536 24746
rect 3570 24712 3604 24746
rect 3638 24712 3672 24746
rect 3706 24712 3740 24746
rect 3774 24712 3808 24746
rect 3842 24712 3876 24746
rect 3910 24712 3944 24746
rect 3978 24712 4012 24746
rect 4046 24712 4080 24746
rect 4114 24712 4148 24746
rect 4182 24712 4216 24746
rect 4250 24712 4284 24746
rect 4318 24712 4352 24746
rect 4386 24712 4420 24746
rect 4454 24712 4488 24746
rect 4522 24712 4556 24746
rect 4590 24712 4624 24746
rect 4658 24712 4692 24746
rect 4726 24712 4760 24746
rect 4794 24712 4828 24746
rect 4862 24712 4896 24746
rect 4930 24712 4964 24746
rect 4998 24712 5032 24746
rect 5066 24712 5100 24746
rect 5134 24712 5168 24746
rect 5202 24712 5236 24746
rect 5270 24712 5304 24746
rect 5338 24712 5372 24746
rect 5406 24712 5440 24746
rect 5474 24712 5508 24746
rect 5542 24712 5576 24746
rect 5610 24712 5644 24746
rect 5678 24712 5712 24746
rect 5746 24712 5780 24746
rect 5814 24712 5848 24746
rect 5882 24712 5916 24746
rect 5950 24712 5984 24746
rect 6018 24712 6052 24746
rect 6086 24712 6120 24746
rect 6154 24712 6188 24746
rect 6222 24712 6256 24746
rect 6290 24712 6324 24746
rect 6358 24712 6392 24746
rect 6426 24712 6460 24746
rect 6494 24712 6528 24746
rect 6562 24712 6596 24746
rect 6630 24712 6664 24746
rect 6698 24712 6732 24746
rect 6766 24712 6800 24746
rect 6834 24712 6868 24746
rect 6902 24712 6936 24746
rect 6970 24712 7004 24746
rect 7038 24712 7072 24746
rect 7106 24712 7140 24746
rect 7174 24712 7208 24746
rect 7242 24712 7276 24746
rect 7310 24712 7344 24746
rect 7378 24712 7412 24746
rect 7446 24712 7480 24746
rect 7514 24712 7548 24746
rect 7582 24712 7616 24746
rect 7650 24712 7684 24746
rect 7718 24712 7752 24746
rect 7786 24712 7820 24746
rect 7854 24712 7888 24746
rect 7922 24712 7956 24746
rect 7990 24712 8024 24746
rect 8058 24712 8092 24746
rect 8126 24712 8160 24746
rect 8194 24712 8228 24746
rect 8262 24712 8296 24746
rect 8330 24712 8364 24746
rect 8398 24712 8432 24746
rect 8466 24712 8500 24746
rect 8534 24712 8568 24746
rect 8602 24712 8636 24746
rect 8670 24712 8704 24746
rect 8738 24712 8772 24746
rect 8806 24712 8840 24746
rect 8874 24712 8908 24746
rect 8942 24712 8976 24746
rect 9010 24712 9044 24746
rect 9078 24712 9112 24746
rect 9146 24712 9180 24746
rect 9214 24712 9248 24746
rect 9282 24712 9316 24746
rect 9350 24712 9384 24746
rect 9418 24712 9452 24746
rect 9486 24712 9520 24746
rect 9554 24712 9588 24746
rect 9622 24712 9656 24746
rect 9690 24712 9724 24746
rect 9758 24712 9792 24746
rect 9826 24712 9860 24746
rect 9894 24712 9928 24746
rect 9962 24712 9996 24746
rect 10030 24712 10064 24746
rect 10098 24712 10132 24746
rect 10166 24712 10200 24746
rect 10234 24712 10268 24746
rect 10302 24712 10336 24746
rect 10370 24712 10404 24746
rect 10438 24712 10472 24746
rect 10506 24712 10540 24746
rect 10574 24712 10608 24746
rect 10642 24712 10676 24746
rect 10710 24712 10744 24746
rect 10778 24712 10812 24746
rect 10846 24712 10880 24746
rect 10914 24712 10948 24746
rect 10982 24712 11016 24746
rect 11050 24712 11084 24746
rect 11118 24712 11152 24746
rect 11186 24712 11220 24746
rect 11254 24712 11288 24746
rect 11322 24712 11356 24746
rect 11390 24712 11424 24746
rect 11458 24712 11492 24746
rect 11526 24712 11560 24746
rect 11594 24712 11628 24746
rect 11662 24712 11696 24746
rect 11730 24712 11764 24746
rect 11798 24712 11832 24746
rect 11866 24712 11900 24746
rect 11934 24712 11968 24746
rect 12002 24712 12036 24746
rect 12070 24712 12104 24746
rect 12138 24712 12172 24746
rect 12206 24712 12240 24746
rect 12274 24712 12308 24746
rect 12342 24712 12376 24746
rect 12410 24712 12444 24746
rect 12478 24712 12512 24746
rect 12546 24712 12580 24746
rect 12614 24712 12648 24746
rect 12682 24712 12716 24746
rect 12750 24712 12784 24746
rect 12818 24712 12852 24746
rect 12886 24712 12920 24746
rect 12954 24712 12988 24746
rect 13022 24712 13056 24746
rect 13090 24712 13124 24746
rect 13158 24712 13192 24746
rect 13226 24712 13260 24746
rect 13294 24712 13328 24746
rect 13362 24712 13396 24746
rect 13430 24712 13464 24746
rect 13498 24712 13532 24746
rect 13566 24712 13600 24746
rect 13634 24712 13668 24746
rect 13702 24712 13736 24746
rect 13770 24712 13804 24746
rect 13838 24712 13872 24746
rect 13906 24712 13940 24746
rect 13974 24712 14008 24746
rect 14042 24712 14076 24746
rect 14110 24712 14144 24746
rect 14178 24712 14212 24746
rect 14246 24712 14280 24746
rect 14314 24712 14348 24746
rect 14382 24712 14416 24746
rect 14450 24712 14484 24746
rect 14518 24712 14552 24746
rect 14586 24712 14620 24746
rect 14654 24712 14688 24746
rect 14722 24712 14756 24746
rect 14790 24712 14824 24746
rect 14858 24712 14882 24746
rect 53 24648 14882 24712
rect 53 24527 14874 24648
rect 53 24463 304 24527
rect 14765 24463 14874 24527
rect 53 19894 261 24463
rect 53 19859 14874 19894
rect 53 19825 77 19859
rect 111 19825 146 19859
rect 180 19825 215 19859
rect 249 19825 284 19859
rect 318 19825 353 19859
rect 387 19825 422 19859
rect 456 19825 491 19859
rect 525 19825 560 19859
rect 594 19825 629 19859
rect 663 19825 698 19859
rect 732 19825 767 19859
rect 801 19825 836 19859
rect 870 19825 905 19859
rect 939 19825 974 19859
rect 1008 19825 1043 19859
rect 1077 19825 1112 19859
rect 1146 19825 1181 19859
rect 1215 19825 1250 19859
rect 1284 19825 1319 19859
rect 1353 19825 1388 19859
rect 1422 19825 1457 19859
rect 1491 19825 1526 19859
rect 1560 19825 1595 19859
rect 1629 19825 1664 19859
rect 1698 19825 1733 19859
rect 1767 19825 1802 19859
rect 1836 19825 1871 19859
rect 1905 19825 1940 19859
rect 1974 19825 2009 19859
rect 2043 19825 2078 19859
rect 2112 19825 2147 19859
rect 2181 19825 2216 19859
rect 2250 19825 2285 19859
rect 2319 19825 2354 19859
rect 2388 19825 2423 19859
rect 2457 19825 2492 19859
rect 2526 19825 2561 19859
rect 2595 19825 2630 19859
rect 2664 19825 2699 19859
rect 2733 19825 2768 19859
rect 2802 19825 2837 19859
rect 2871 19825 2906 19859
rect 2940 19825 2975 19859
rect 3009 19825 3044 19859
rect 3078 19825 3113 19859
rect 3147 19825 3182 19859
rect 53 19791 3182 19825
rect 53 19757 77 19791
rect 111 19757 146 19791
rect 180 19757 215 19791
rect 249 19757 284 19791
rect 318 19757 353 19791
rect 387 19757 422 19791
rect 456 19757 491 19791
rect 525 19757 560 19791
rect 594 19757 629 19791
rect 663 19757 698 19791
rect 732 19757 767 19791
rect 801 19757 836 19791
rect 870 19757 905 19791
rect 939 19757 974 19791
rect 1008 19757 1043 19791
rect 1077 19757 1112 19791
rect 1146 19757 1181 19791
rect 1215 19757 1250 19791
rect 1284 19757 1319 19791
rect 1353 19757 1388 19791
rect 1422 19757 1457 19791
rect 1491 19757 1526 19791
rect 1560 19757 1595 19791
rect 1629 19757 1664 19791
rect 1698 19757 1733 19791
rect 1767 19757 1802 19791
rect 1836 19757 1871 19791
rect 1905 19757 1940 19791
rect 1974 19757 2009 19791
rect 2043 19757 2078 19791
rect 2112 19757 2147 19791
rect 2181 19757 2216 19791
rect 2250 19757 2285 19791
rect 2319 19757 2354 19791
rect 2388 19757 2423 19791
rect 2457 19757 2492 19791
rect 2526 19757 2561 19791
rect 2595 19757 2630 19791
rect 2664 19757 2699 19791
rect 2733 19757 2768 19791
rect 2802 19757 2837 19791
rect 2871 19757 2906 19791
rect 2940 19757 2975 19791
rect 3009 19757 3044 19791
rect 3078 19757 3113 19791
rect 3147 19757 3182 19791
rect 53 19723 3182 19757
rect 53 19689 77 19723
rect 111 19689 146 19723
rect 180 19689 215 19723
rect 249 19689 284 19723
rect 318 19689 353 19723
rect 387 19689 422 19723
rect 456 19689 491 19723
rect 525 19689 560 19723
rect 594 19689 629 19723
rect 663 19689 698 19723
rect 732 19689 767 19723
rect 801 19689 836 19723
rect 870 19689 905 19723
rect 939 19689 974 19723
rect 1008 19689 1043 19723
rect 1077 19689 1112 19723
rect 1146 19689 1181 19723
rect 1215 19689 1250 19723
rect 1284 19689 1319 19723
rect 1353 19689 1388 19723
rect 1422 19689 1457 19723
rect 1491 19689 1526 19723
rect 1560 19689 1595 19723
rect 1629 19689 1664 19723
rect 1698 19689 1733 19723
rect 1767 19689 1802 19723
rect 1836 19689 1871 19723
rect 1905 19689 1940 19723
rect 1974 19689 2009 19723
rect 2043 19689 2078 19723
rect 2112 19689 2147 19723
rect 2181 19689 2216 19723
rect 2250 19689 2285 19723
rect 2319 19689 2354 19723
rect 2388 19689 2423 19723
rect 2457 19689 2492 19723
rect 2526 19689 2561 19723
rect 2595 19689 2630 19723
rect 2664 19689 2699 19723
rect 2733 19689 2768 19723
rect 2802 19689 2837 19723
rect 2871 19689 2906 19723
rect 2940 19689 2975 19723
rect 3009 19689 3044 19723
rect 3078 19689 3113 19723
rect 3147 19689 3182 19723
rect 53 19655 3182 19689
rect 53 19621 77 19655
rect 111 19621 146 19655
rect 180 19621 215 19655
rect 249 19621 284 19655
rect 318 19621 353 19655
rect 387 19621 422 19655
rect 456 19621 491 19655
rect 525 19621 560 19655
rect 594 19621 629 19655
rect 663 19621 698 19655
rect 732 19621 767 19655
rect 801 19621 836 19655
rect 870 19621 905 19655
rect 939 19621 974 19655
rect 1008 19621 1043 19655
rect 1077 19621 1112 19655
rect 1146 19621 1181 19655
rect 1215 19621 1250 19655
rect 1284 19621 1319 19655
rect 1353 19621 1388 19655
rect 1422 19621 1457 19655
rect 1491 19621 1526 19655
rect 1560 19621 1595 19655
rect 1629 19621 1664 19655
rect 1698 19621 1733 19655
rect 1767 19621 1802 19655
rect 1836 19621 1871 19655
rect 1905 19621 1940 19655
rect 1974 19621 2009 19655
rect 2043 19621 2078 19655
rect 2112 19621 2147 19655
rect 2181 19621 2216 19655
rect 2250 19621 2285 19655
rect 2319 19621 2354 19655
rect 2388 19621 2423 19655
rect 2457 19621 2492 19655
rect 2526 19621 2561 19655
rect 2595 19621 2630 19655
rect 2664 19621 2699 19655
rect 2733 19621 2768 19655
rect 2802 19621 2837 19655
rect 2871 19621 2906 19655
rect 2940 19621 2975 19655
rect 3009 19621 3044 19655
rect 3078 19621 3113 19655
rect 3147 19621 3182 19655
rect 14436 19831 14874 19859
rect 14436 19797 14484 19831
rect 14518 19797 14567 19831
rect 14601 19797 14650 19831
rect 14684 19797 14733 19831
rect 14767 19797 14816 19831
rect 14850 19797 14874 19831
rect 14436 19761 14874 19797
rect 14436 19727 14484 19761
rect 14518 19727 14567 19761
rect 14601 19727 14650 19761
rect 14684 19727 14733 19761
rect 14767 19727 14816 19761
rect 14850 19727 14874 19761
rect 14436 19691 14874 19727
rect 14436 19657 14484 19691
rect 14518 19657 14567 19691
rect 14601 19657 14650 19691
rect 14684 19657 14733 19691
rect 14767 19657 14816 19691
rect 14850 19657 14874 19691
rect 14436 19621 14874 19657
rect 53 19587 14484 19621
rect 14518 19587 14567 19621
rect 14601 19587 14650 19621
rect 14684 19587 14733 19621
rect 14767 19587 14816 19621
rect 14850 19587 14874 19621
rect 53 19585 14874 19587
rect 53 19551 77 19585
rect 111 19551 146 19585
rect 180 19551 215 19585
rect 249 19551 284 19585
rect 318 19551 353 19585
rect 387 19551 422 19585
rect 456 19551 491 19585
rect 525 19551 560 19585
rect 594 19551 629 19585
rect 663 19551 698 19585
rect 732 19551 767 19585
rect 801 19551 836 19585
rect 870 19551 905 19585
rect 939 19551 974 19585
rect 1008 19551 1043 19585
rect 1077 19551 1112 19585
rect 1146 19551 1181 19585
rect 1215 19551 1250 19585
rect 1284 19551 1319 19585
rect 1353 19551 1388 19585
rect 1422 19551 1457 19585
rect 1491 19551 1526 19585
rect 1560 19551 1595 19585
rect 1629 19551 1664 19585
rect 1698 19551 1733 19585
rect 1767 19551 1802 19585
rect 1836 19551 1871 19585
rect 1905 19551 1940 19585
rect 1974 19551 2009 19585
rect 2043 19551 2078 19585
rect 2112 19551 2147 19585
rect 2181 19551 2216 19585
rect 2250 19551 2285 19585
rect 2319 19551 2354 19585
rect 2388 19551 2423 19585
rect 2457 19551 2492 19585
rect 2526 19551 2561 19585
rect 2595 19551 2630 19585
rect 2664 19551 2699 19585
rect 2733 19551 2768 19585
rect 2802 19551 2837 19585
rect 2871 19551 2906 19585
rect 2940 19551 2975 19585
rect 3009 19551 3044 19585
rect 3078 19551 3113 19585
rect 3147 19551 3182 19585
rect 3216 19551 3251 19585
rect 3285 19551 3320 19585
rect 3354 19551 3389 19585
rect 3423 19551 3458 19585
rect 3492 19551 3527 19585
rect 3561 19551 3596 19585
rect 3630 19551 3665 19585
rect 3699 19551 3733 19585
rect 3767 19551 3801 19585
rect 3835 19551 3869 19585
rect 3903 19551 3937 19585
rect 3971 19551 4005 19585
rect 4039 19551 4073 19585
rect 4107 19551 4141 19585
rect 4175 19551 4209 19585
rect 4243 19551 4277 19585
rect 4311 19551 4345 19585
rect 4379 19551 4413 19585
rect 4447 19551 4481 19585
rect 4515 19551 4549 19585
rect 4583 19551 4617 19585
rect 4651 19551 4685 19585
rect 4719 19551 4753 19585
rect 4787 19551 4821 19585
rect 4855 19551 4889 19585
rect 4923 19551 4957 19585
rect 4991 19551 5025 19585
rect 5059 19551 5093 19585
rect 5127 19551 5161 19585
rect 5195 19551 5229 19585
rect 5263 19551 5297 19585
rect 5331 19551 5365 19585
rect 5399 19551 5433 19585
rect 5467 19551 5501 19585
rect 5535 19551 5569 19585
rect 5603 19551 5637 19585
rect 5671 19551 5705 19585
rect 5739 19551 5773 19585
rect 5807 19551 5841 19585
rect 5875 19551 5909 19585
rect 5943 19551 5977 19585
rect 6011 19551 6045 19585
rect 6079 19551 6113 19585
rect 6147 19551 6181 19585
rect 6215 19551 6249 19585
rect 6283 19551 6317 19585
rect 6351 19551 6385 19585
rect 6419 19551 6453 19585
rect 6487 19551 6521 19585
rect 6555 19551 6589 19585
rect 6623 19551 6657 19585
rect 6691 19551 6725 19585
rect 6759 19551 6793 19585
rect 6827 19551 6861 19585
rect 6895 19551 6929 19585
rect 6963 19551 6997 19585
rect 7031 19551 7065 19585
rect 7099 19551 7133 19585
rect 7167 19551 7201 19585
rect 7235 19551 7269 19585
rect 7303 19551 7337 19585
rect 7371 19551 7405 19585
rect 7439 19551 7473 19585
rect 7507 19551 7541 19585
rect 7575 19551 7609 19585
rect 7643 19551 7677 19585
rect 7711 19551 7745 19585
rect 7779 19551 7813 19585
rect 7847 19551 7881 19585
rect 7915 19551 7949 19585
rect 7983 19551 8017 19585
rect 8051 19551 8085 19585
rect 8119 19551 8153 19585
rect 8187 19551 8221 19585
rect 8255 19551 8289 19585
rect 8323 19551 8357 19585
rect 8391 19551 8425 19585
rect 8459 19551 8493 19585
rect 8527 19551 8561 19585
rect 8595 19551 8629 19585
rect 8663 19551 8697 19585
rect 8731 19551 8765 19585
rect 8799 19551 8833 19585
rect 8867 19551 8901 19585
rect 8935 19551 8969 19585
rect 9003 19551 9037 19585
rect 9071 19551 9105 19585
rect 9139 19551 9173 19585
rect 9207 19551 9241 19585
rect 9275 19551 9309 19585
rect 9343 19551 9377 19585
rect 9411 19551 9445 19585
rect 9479 19551 9513 19585
rect 9547 19551 9581 19585
rect 9615 19551 9649 19585
rect 9683 19551 9717 19585
rect 9751 19551 9785 19585
rect 9819 19551 9853 19585
rect 9887 19551 9921 19585
rect 9955 19551 9989 19585
rect 10023 19551 10057 19585
rect 10091 19551 10125 19585
rect 10159 19551 10193 19585
rect 10227 19551 10261 19585
rect 10295 19551 10329 19585
rect 10363 19551 10397 19585
rect 10431 19551 10465 19585
rect 10499 19551 10533 19585
rect 10567 19551 10601 19585
rect 10635 19551 10669 19585
rect 10703 19551 10737 19585
rect 10771 19551 10805 19585
rect 10839 19551 10873 19585
rect 10907 19551 10941 19585
rect 10975 19551 11009 19585
rect 11043 19551 11077 19585
rect 11111 19551 11145 19585
rect 11179 19551 11213 19585
rect 11247 19551 11281 19585
rect 11315 19551 11349 19585
rect 11383 19551 11417 19585
rect 11451 19551 11485 19585
rect 11519 19551 11553 19585
rect 11587 19551 11621 19585
rect 11655 19551 11689 19585
rect 11723 19557 14874 19585
rect 11723 19551 11771 19557
rect 53 19523 11771 19551
rect 11805 19523 11841 19557
rect 11875 19523 11911 19557
rect 11945 19523 11981 19557
rect 12015 19523 12051 19557
rect 12085 19523 12121 19557
rect 12155 19523 12191 19557
rect 12225 19523 12261 19557
rect 12295 19523 12331 19557
rect 12365 19523 12401 19557
rect 12435 19523 12470 19557
rect 12504 19523 12539 19557
rect 12573 19523 12608 19557
rect 12642 19523 12677 19557
rect 12711 19523 12746 19557
rect 12780 19523 12815 19557
rect 12849 19523 12884 19557
rect 12918 19523 12953 19557
rect 12987 19523 13022 19557
rect 13056 19523 13091 19557
rect 13125 19523 13160 19557
rect 13194 19523 13229 19557
rect 13263 19523 13298 19557
rect 13332 19523 13367 19557
rect 13401 19523 13436 19557
rect 13470 19523 13505 19557
rect 13539 19523 13574 19557
rect 13608 19523 13643 19557
rect 13677 19523 13712 19557
rect 13746 19523 13781 19557
rect 13815 19523 13850 19557
rect 13884 19523 13919 19557
rect 13953 19523 13988 19557
rect 14022 19523 14057 19557
rect 14091 19523 14126 19557
rect 14160 19523 14195 19557
rect 14229 19523 14264 19557
rect 14298 19523 14333 19557
rect 14367 19523 14402 19557
rect 14436 19551 14874 19557
rect 14436 19523 14484 19551
rect 53 19517 14484 19523
rect 14518 19517 14567 19551
rect 14601 19517 14650 19551
rect 14684 19517 14733 19551
rect 14767 19517 14816 19551
rect 14850 19517 14874 19551
rect 53 19513 14874 19517
rect 53 19479 77 19513
rect 111 19479 146 19513
rect 180 19479 215 19513
rect 249 19479 284 19513
rect 318 19479 353 19513
rect 387 19479 422 19513
rect 456 19479 491 19513
rect 525 19479 560 19513
rect 594 19479 629 19513
rect 663 19479 698 19513
rect 732 19479 767 19513
rect 801 19479 836 19513
rect 870 19479 905 19513
rect 939 19479 974 19513
rect 1008 19479 1043 19513
rect 1077 19479 1112 19513
rect 1146 19479 1181 19513
rect 1215 19479 1250 19513
rect 1284 19479 1319 19513
rect 1353 19479 1388 19513
rect 1422 19479 1457 19513
rect 1491 19479 1526 19513
rect 1560 19479 1595 19513
rect 1629 19479 1664 19513
rect 1698 19479 1733 19513
rect 1767 19479 1802 19513
rect 1836 19479 1871 19513
rect 1905 19479 1940 19513
rect 1974 19479 2009 19513
rect 2043 19479 2078 19513
rect 2112 19479 2147 19513
rect 2181 19479 2216 19513
rect 2250 19479 2285 19513
rect 2319 19479 2354 19513
rect 2388 19479 2423 19513
rect 2457 19479 2492 19513
rect 2526 19479 2561 19513
rect 2595 19479 2630 19513
rect 2664 19479 2699 19513
rect 2733 19479 2768 19513
rect 2802 19479 2837 19513
rect 2871 19479 2906 19513
rect 2940 19479 2975 19513
rect 3009 19479 3044 19513
rect 3078 19479 3113 19513
rect 3147 19479 3182 19513
rect 3216 19479 3251 19513
rect 3285 19479 3320 19513
rect 3354 19479 3389 19513
rect 3423 19479 3458 19513
rect 3492 19479 3527 19513
rect 3561 19479 3596 19513
rect 3630 19479 3665 19513
rect 3699 19479 3733 19513
rect 3767 19479 3801 19513
rect 3835 19479 3869 19513
rect 3903 19479 3937 19513
rect 3971 19479 4005 19513
rect 4039 19479 4073 19513
rect 4107 19479 4141 19513
rect 4175 19479 4209 19513
rect 4243 19479 4277 19513
rect 4311 19479 4345 19513
rect 4379 19479 4413 19513
rect 4447 19479 4481 19513
rect 4515 19479 4549 19513
rect 4583 19479 4617 19513
rect 4651 19479 4685 19513
rect 4719 19479 4753 19513
rect 4787 19479 4821 19513
rect 4855 19479 4889 19513
rect 4923 19479 4957 19513
rect 4991 19479 5025 19513
rect 5059 19479 5093 19513
rect 5127 19479 5161 19513
rect 5195 19479 5229 19513
rect 5263 19479 5297 19513
rect 5331 19479 5365 19513
rect 5399 19479 5433 19513
rect 5467 19479 5501 19513
rect 5535 19479 5569 19513
rect 5603 19479 5637 19513
rect 5671 19479 5705 19513
rect 5739 19479 5773 19513
rect 5807 19479 5841 19513
rect 5875 19479 5909 19513
rect 5943 19479 5977 19513
rect 6011 19479 6045 19513
rect 6079 19479 6113 19513
rect 6147 19479 6181 19513
rect 6215 19479 6249 19513
rect 6283 19479 6317 19513
rect 6351 19479 6385 19513
rect 6419 19479 6453 19513
rect 6487 19479 6521 19513
rect 6555 19479 6589 19513
rect 6623 19479 6657 19513
rect 6691 19479 6725 19513
rect 6759 19479 6793 19513
rect 6827 19479 6861 19513
rect 6895 19479 6929 19513
rect 6963 19479 6997 19513
rect 7031 19479 7065 19513
rect 7099 19479 7133 19513
rect 7167 19479 7201 19513
rect 7235 19479 7269 19513
rect 7303 19479 7337 19513
rect 7371 19479 7405 19513
rect 7439 19479 7473 19513
rect 7507 19479 7541 19513
rect 7575 19479 7609 19513
rect 7643 19479 7677 19513
rect 7711 19479 7745 19513
rect 7779 19479 7813 19513
rect 7847 19479 7881 19513
rect 7915 19479 7949 19513
rect 7983 19479 8017 19513
rect 8051 19479 8085 19513
rect 8119 19479 8153 19513
rect 8187 19479 8221 19513
rect 8255 19479 8289 19513
rect 8323 19479 8357 19513
rect 8391 19479 8425 19513
rect 8459 19479 8493 19513
rect 8527 19479 8561 19513
rect 8595 19479 8629 19513
rect 8663 19479 8697 19513
rect 8731 19479 8765 19513
rect 8799 19479 8833 19513
rect 8867 19479 8901 19513
rect 8935 19479 8969 19513
rect 9003 19479 9037 19513
rect 9071 19479 9105 19513
rect 9139 19479 9173 19513
rect 9207 19479 9241 19513
rect 9275 19479 9309 19513
rect 9343 19479 9377 19513
rect 9411 19479 9445 19513
rect 9479 19479 9513 19513
rect 9547 19479 9581 19513
rect 9615 19479 9649 19513
rect 9683 19479 9717 19513
rect 9751 19479 9785 19513
rect 9819 19479 9853 19513
rect 9887 19479 9921 19513
rect 9955 19479 9989 19513
rect 10023 19479 10057 19513
rect 10091 19479 10125 19513
rect 10159 19479 10193 19513
rect 10227 19479 10261 19513
rect 10295 19479 10329 19513
rect 10363 19479 10397 19513
rect 10431 19479 10465 19513
rect 10499 19479 10533 19513
rect 10567 19479 10601 19513
rect 10635 19479 10669 19513
rect 10703 19479 10737 19513
rect 10771 19479 10805 19513
rect 10839 19479 10873 19513
rect 10907 19479 10941 19513
rect 10975 19479 11009 19513
rect 11043 19479 11077 19513
rect 11111 19479 11145 19513
rect 11179 19479 11213 19513
rect 11247 19479 11281 19513
rect 11315 19479 11349 19513
rect 11383 19479 11417 19513
rect 11451 19479 11485 19513
rect 11519 19479 11553 19513
rect 11587 19479 11621 19513
rect 11655 19479 11689 19513
rect 11723 19481 14874 19513
rect 11723 19479 14484 19481
rect 53 19477 14484 19479
rect 53 19443 11771 19477
rect 11805 19443 11841 19477
rect 11875 19443 11911 19477
rect 11945 19443 11981 19477
rect 12015 19443 12051 19477
rect 12085 19443 12121 19477
rect 12155 19443 12191 19477
rect 12225 19443 12261 19477
rect 12295 19443 12331 19477
rect 12365 19443 12401 19477
rect 12435 19443 12470 19477
rect 12504 19443 12539 19477
rect 12573 19443 12608 19477
rect 12642 19443 12677 19477
rect 12711 19443 12746 19477
rect 12780 19443 12815 19477
rect 12849 19443 12884 19477
rect 12918 19443 12953 19477
rect 12987 19443 13022 19477
rect 13056 19443 13091 19477
rect 13125 19443 13160 19477
rect 13194 19443 13229 19477
rect 13263 19443 13298 19477
rect 13332 19443 13367 19477
rect 13401 19443 13436 19477
rect 13470 19443 13505 19477
rect 13539 19443 13574 19477
rect 13608 19443 13643 19477
rect 13677 19443 13712 19477
rect 13746 19443 13781 19477
rect 13815 19443 13850 19477
rect 13884 19443 13919 19477
rect 13953 19443 13988 19477
rect 14022 19443 14057 19477
rect 14091 19443 14126 19477
rect 14160 19443 14195 19477
rect 14229 19443 14264 19477
rect 14298 19443 14333 19477
rect 14367 19443 14402 19477
rect 14436 19447 14484 19477
rect 14518 19447 14567 19481
rect 14601 19447 14650 19481
rect 14684 19447 14733 19481
rect 14767 19447 14816 19481
rect 14850 19447 14874 19481
rect 14436 19443 14874 19447
rect 53 19441 14874 19443
rect 53 19407 77 19441
rect 111 19407 146 19441
rect 180 19407 215 19441
rect 249 19407 284 19441
rect 318 19407 353 19441
rect 387 19407 422 19441
rect 456 19407 491 19441
rect 525 19407 560 19441
rect 594 19407 629 19441
rect 663 19407 698 19441
rect 732 19407 767 19441
rect 801 19407 836 19441
rect 870 19407 905 19441
rect 939 19407 974 19441
rect 1008 19407 1043 19441
rect 1077 19407 1112 19441
rect 1146 19407 1181 19441
rect 1215 19407 1250 19441
rect 1284 19407 1319 19441
rect 1353 19407 1388 19441
rect 1422 19407 1457 19441
rect 1491 19407 1526 19441
rect 1560 19407 1595 19441
rect 1629 19407 1664 19441
rect 1698 19407 1733 19441
rect 1767 19407 1802 19441
rect 1836 19407 1871 19441
rect 1905 19407 1940 19441
rect 1974 19407 2009 19441
rect 2043 19407 2078 19441
rect 2112 19407 2147 19441
rect 2181 19407 2216 19441
rect 2250 19407 2285 19441
rect 2319 19407 2354 19441
rect 2388 19407 2423 19441
rect 2457 19407 2492 19441
rect 2526 19407 2561 19441
rect 2595 19407 2630 19441
rect 2664 19407 2699 19441
rect 2733 19407 2768 19441
rect 2802 19407 2837 19441
rect 2871 19407 2906 19441
rect 2940 19407 2975 19441
rect 3009 19407 3044 19441
rect 3078 19407 3113 19441
rect 3147 19407 3182 19441
rect 3216 19407 3251 19441
rect 3285 19407 3320 19441
rect 3354 19407 3389 19441
rect 3423 19407 3458 19441
rect 3492 19407 3527 19441
rect 3561 19407 3596 19441
rect 3630 19407 3665 19441
rect 3699 19407 3733 19441
rect 3767 19407 3801 19441
rect 3835 19407 3869 19441
rect 3903 19407 3937 19441
rect 3971 19407 4005 19441
rect 4039 19407 4073 19441
rect 4107 19407 4141 19441
rect 4175 19407 4209 19441
rect 4243 19407 4277 19441
rect 4311 19407 4345 19441
rect 4379 19407 4413 19441
rect 4447 19407 4481 19441
rect 4515 19407 4549 19441
rect 4583 19407 4617 19441
rect 4651 19407 4685 19441
rect 4719 19407 4753 19441
rect 4787 19407 4821 19441
rect 4855 19407 4889 19441
rect 4923 19407 4957 19441
rect 4991 19407 5025 19441
rect 5059 19407 5093 19441
rect 5127 19407 5161 19441
rect 5195 19407 5229 19441
rect 5263 19407 5297 19441
rect 5331 19407 5365 19441
rect 5399 19407 5433 19441
rect 5467 19407 5501 19441
rect 5535 19407 5569 19441
rect 5603 19407 5637 19441
rect 5671 19407 5705 19441
rect 5739 19407 5773 19441
rect 5807 19407 5841 19441
rect 5875 19407 5909 19441
rect 5943 19407 5977 19441
rect 6011 19407 6045 19441
rect 6079 19407 6113 19441
rect 6147 19407 6181 19441
rect 6215 19407 6249 19441
rect 6283 19407 6317 19441
rect 6351 19407 6385 19441
rect 6419 19407 6453 19441
rect 6487 19407 6521 19441
rect 6555 19407 6589 19441
rect 6623 19407 6657 19441
rect 6691 19407 6725 19441
rect 6759 19407 6793 19441
rect 6827 19407 6861 19441
rect 6895 19407 6929 19441
rect 6963 19407 6997 19441
rect 7031 19407 7065 19441
rect 7099 19407 7133 19441
rect 7167 19407 7201 19441
rect 7235 19407 7269 19441
rect 7303 19407 7337 19441
rect 7371 19407 7405 19441
rect 7439 19407 7473 19441
rect 7507 19407 7541 19441
rect 7575 19407 7609 19441
rect 7643 19407 7677 19441
rect 7711 19407 7745 19441
rect 7779 19407 7813 19441
rect 7847 19407 7881 19441
rect 7915 19407 7949 19441
rect 7983 19407 8017 19441
rect 8051 19407 8085 19441
rect 8119 19407 8153 19441
rect 8187 19407 8221 19441
rect 8255 19407 8289 19441
rect 8323 19407 8357 19441
rect 8391 19407 8425 19441
rect 8459 19407 8493 19441
rect 8527 19407 8561 19441
rect 8595 19407 8629 19441
rect 8663 19407 8697 19441
rect 8731 19407 8765 19441
rect 8799 19407 8833 19441
rect 8867 19407 8901 19441
rect 8935 19407 8969 19441
rect 9003 19407 9037 19441
rect 9071 19407 9105 19441
rect 9139 19407 9173 19441
rect 9207 19407 9241 19441
rect 9275 19407 9309 19441
rect 9343 19407 9377 19441
rect 9411 19407 9445 19441
rect 9479 19407 9513 19441
rect 9547 19407 9581 19441
rect 9615 19407 9649 19441
rect 9683 19407 9717 19441
rect 9751 19407 9785 19441
rect 9819 19407 9853 19441
rect 9887 19407 9921 19441
rect 9955 19407 9989 19441
rect 10023 19407 10057 19441
rect 10091 19407 10125 19441
rect 10159 19407 10193 19441
rect 10227 19407 10261 19441
rect 10295 19407 10329 19441
rect 10363 19407 10397 19441
rect 10431 19407 10465 19441
rect 10499 19407 10533 19441
rect 10567 19407 10601 19441
rect 10635 19407 10669 19441
rect 10703 19407 10737 19441
rect 10771 19407 10805 19441
rect 10839 19407 10873 19441
rect 10907 19407 10941 19441
rect 10975 19407 11009 19441
rect 11043 19407 11077 19441
rect 11111 19407 11145 19441
rect 11179 19407 11213 19441
rect 11247 19407 11281 19441
rect 11315 19407 11349 19441
rect 11383 19407 11417 19441
rect 11451 19407 11485 19441
rect 11519 19407 11553 19441
rect 11587 19407 11621 19441
rect 11655 19407 11689 19441
rect 11723 19411 14874 19441
rect 11723 19407 14484 19411
rect 53 19397 14484 19407
rect 53 19369 11771 19397
rect 53 19335 77 19369
rect 111 19335 146 19369
rect 180 19335 215 19369
rect 249 19335 284 19369
rect 318 19335 353 19369
rect 387 19335 422 19369
rect 456 19335 491 19369
rect 525 19335 560 19369
rect 594 19335 629 19369
rect 663 19335 698 19369
rect 732 19335 767 19369
rect 801 19335 836 19369
rect 870 19335 905 19369
rect 939 19335 974 19369
rect 1008 19335 1043 19369
rect 1077 19335 1112 19369
rect 1146 19335 1181 19369
rect 1215 19335 1250 19369
rect 1284 19335 1319 19369
rect 1353 19335 1388 19369
rect 1422 19335 1457 19369
rect 1491 19335 1526 19369
rect 1560 19335 1595 19369
rect 1629 19335 1664 19369
rect 1698 19335 1733 19369
rect 1767 19335 1802 19369
rect 1836 19335 1871 19369
rect 1905 19335 1940 19369
rect 1974 19335 2009 19369
rect 2043 19335 2078 19369
rect 2112 19335 2147 19369
rect 2181 19335 2216 19369
rect 2250 19335 2285 19369
rect 2319 19335 2354 19369
rect 2388 19335 2423 19369
rect 2457 19335 2492 19369
rect 2526 19335 2561 19369
rect 2595 19335 2630 19369
rect 2664 19335 2699 19369
rect 2733 19335 2768 19369
rect 2802 19335 2837 19369
rect 2871 19335 2906 19369
rect 2940 19335 2975 19369
rect 3009 19335 3044 19369
rect 3078 19335 3113 19369
rect 3147 19335 3182 19369
rect 3216 19335 3251 19369
rect 3285 19335 3320 19369
rect 3354 19335 3389 19369
rect 3423 19335 3458 19369
rect 3492 19335 3527 19369
rect 3561 19335 3596 19369
rect 3630 19335 3665 19369
rect 3699 19335 3733 19369
rect 3767 19335 3801 19369
rect 3835 19335 3869 19369
rect 3903 19335 3937 19369
rect 3971 19335 4005 19369
rect 4039 19335 4073 19369
rect 4107 19335 4141 19369
rect 4175 19335 4209 19369
rect 4243 19335 4277 19369
rect 4311 19335 4345 19369
rect 4379 19335 4413 19369
rect 4447 19335 4481 19369
rect 4515 19335 4549 19369
rect 4583 19335 4617 19369
rect 4651 19335 4685 19369
rect 4719 19335 4753 19369
rect 4787 19335 4821 19369
rect 4855 19335 4889 19369
rect 4923 19335 4957 19369
rect 4991 19335 5025 19369
rect 5059 19335 5093 19369
rect 5127 19335 5161 19369
rect 5195 19335 5229 19369
rect 5263 19335 5297 19369
rect 5331 19335 5365 19369
rect 5399 19335 5433 19369
rect 5467 19335 5501 19369
rect 5535 19335 5569 19369
rect 5603 19335 5637 19369
rect 5671 19335 5705 19369
rect 5739 19335 5773 19369
rect 5807 19335 5841 19369
rect 5875 19335 5909 19369
rect 5943 19335 5977 19369
rect 6011 19335 6045 19369
rect 6079 19335 6113 19369
rect 6147 19335 6181 19369
rect 6215 19335 6249 19369
rect 6283 19335 6317 19369
rect 6351 19335 6385 19369
rect 6419 19335 6453 19369
rect 6487 19335 6521 19369
rect 6555 19335 6589 19369
rect 6623 19335 6657 19369
rect 6691 19335 6725 19369
rect 6759 19335 6793 19369
rect 6827 19335 6861 19369
rect 6895 19335 6929 19369
rect 6963 19335 6997 19369
rect 7031 19335 7065 19369
rect 7099 19335 7133 19369
rect 7167 19335 7201 19369
rect 7235 19335 7269 19369
rect 7303 19335 7337 19369
rect 7371 19335 7405 19369
rect 7439 19335 7473 19369
rect 7507 19335 7541 19369
rect 7575 19335 7609 19369
rect 7643 19335 7677 19369
rect 7711 19335 7745 19369
rect 7779 19335 7813 19369
rect 7847 19335 7881 19369
rect 7915 19335 7949 19369
rect 7983 19335 8017 19369
rect 8051 19335 8085 19369
rect 8119 19335 8153 19369
rect 8187 19335 8221 19369
rect 8255 19335 8289 19369
rect 8323 19335 8357 19369
rect 8391 19335 8425 19369
rect 8459 19335 8493 19369
rect 8527 19335 8561 19369
rect 8595 19335 8629 19369
rect 8663 19335 8697 19369
rect 8731 19335 8765 19369
rect 8799 19335 8833 19369
rect 8867 19335 8901 19369
rect 8935 19335 8969 19369
rect 9003 19335 9037 19369
rect 9071 19335 9105 19369
rect 9139 19335 9173 19369
rect 9207 19335 9241 19369
rect 9275 19335 9309 19369
rect 9343 19335 9377 19369
rect 9411 19335 9445 19369
rect 9479 19335 9513 19369
rect 9547 19335 9581 19369
rect 9615 19335 9649 19369
rect 9683 19335 9717 19369
rect 9751 19335 9785 19369
rect 9819 19335 9853 19369
rect 9887 19335 9921 19369
rect 9955 19335 9989 19369
rect 10023 19335 10057 19369
rect 10091 19335 10125 19369
rect 10159 19335 10193 19369
rect 10227 19335 10261 19369
rect 10295 19335 10329 19369
rect 10363 19335 10397 19369
rect 10431 19335 10465 19369
rect 10499 19335 10533 19369
rect 10567 19335 10601 19369
rect 10635 19335 10669 19369
rect 10703 19335 10737 19369
rect 10771 19335 10805 19369
rect 10839 19335 10873 19369
rect 10907 19335 10941 19369
rect 10975 19335 11009 19369
rect 11043 19335 11077 19369
rect 11111 19335 11145 19369
rect 11179 19335 11213 19369
rect 11247 19335 11281 19369
rect 11315 19335 11349 19369
rect 11383 19335 11417 19369
rect 11451 19335 11485 19369
rect 11519 19335 11553 19369
rect 11587 19335 11621 19369
rect 11655 19335 11689 19369
rect 11723 19363 11771 19369
rect 11805 19363 11841 19397
rect 11875 19363 11911 19397
rect 11945 19363 11981 19397
rect 12015 19363 12051 19397
rect 12085 19363 12121 19397
rect 12155 19363 12191 19397
rect 12225 19363 12261 19397
rect 12295 19363 12331 19397
rect 12365 19363 12401 19397
rect 12435 19363 12470 19397
rect 12504 19363 12539 19397
rect 12573 19363 12608 19397
rect 12642 19363 12677 19397
rect 12711 19363 12746 19397
rect 12780 19363 12815 19397
rect 12849 19363 12884 19397
rect 12918 19363 12953 19397
rect 12987 19363 13022 19397
rect 13056 19363 13091 19397
rect 13125 19363 13160 19397
rect 13194 19363 13229 19397
rect 13263 19363 13298 19397
rect 13332 19363 13367 19397
rect 13401 19363 13436 19397
rect 13470 19363 13505 19397
rect 13539 19363 13574 19397
rect 13608 19363 13643 19397
rect 13677 19363 13712 19397
rect 13746 19363 13781 19397
rect 13815 19363 13850 19397
rect 13884 19363 13919 19397
rect 13953 19363 13988 19397
rect 14022 19363 14057 19397
rect 14091 19363 14126 19397
rect 14160 19363 14195 19397
rect 14229 19363 14264 19397
rect 14298 19363 14333 19397
rect 14367 19363 14402 19397
rect 14436 19377 14484 19397
rect 14518 19377 14567 19411
rect 14601 19377 14650 19411
rect 14684 19377 14733 19411
rect 14767 19377 14816 19411
rect 14850 19377 14874 19411
rect 14436 19363 14874 19377
rect 11723 19341 14874 19363
rect 11723 19335 14484 19341
rect 53 19330 14484 19335
rect 53 19297 11747 19330
rect 53 19263 77 19297
rect 111 19263 146 19297
rect 180 19263 215 19297
rect 249 19263 284 19297
rect 318 19263 353 19297
rect 387 19263 422 19297
rect 456 19263 491 19297
rect 525 19263 560 19297
rect 594 19263 629 19297
rect 663 19263 698 19297
rect 732 19263 767 19297
rect 801 19263 836 19297
rect 870 19263 905 19297
rect 939 19263 974 19297
rect 1008 19263 1043 19297
rect 1077 19263 1112 19297
rect 1146 19263 1181 19297
rect 1215 19263 1250 19297
rect 1284 19263 1319 19297
rect 1353 19263 1388 19297
rect 1422 19263 1457 19297
rect 1491 19263 1526 19297
rect 1560 19263 1595 19297
rect 1629 19263 1664 19297
rect 1698 19263 1733 19297
rect 1767 19263 1802 19297
rect 1836 19263 1871 19297
rect 1905 19263 1940 19297
rect 1974 19263 2009 19297
rect 2043 19263 2078 19297
rect 2112 19263 2147 19297
rect 2181 19263 2216 19297
rect 2250 19263 2285 19297
rect 2319 19263 2354 19297
rect 2388 19263 2423 19297
rect 2457 19263 2492 19297
rect 2526 19263 2561 19297
rect 2595 19263 2630 19297
rect 2664 19263 2699 19297
rect 2733 19263 2768 19297
rect 2802 19263 2837 19297
rect 2871 19263 2906 19297
rect 2940 19263 2975 19297
rect 3009 19263 3044 19297
rect 3078 19263 3113 19297
rect 3147 19263 3182 19297
rect 3216 19263 3251 19297
rect 3285 19263 3320 19297
rect 3354 19263 3389 19297
rect 3423 19263 3458 19297
rect 3492 19263 3527 19297
rect 3561 19263 3596 19297
rect 3630 19263 3665 19297
rect 3699 19263 3733 19297
rect 3767 19263 3801 19297
rect 3835 19263 3869 19297
rect 3903 19263 3937 19297
rect 3971 19263 4005 19297
rect 4039 19263 4073 19297
rect 4107 19263 4141 19297
rect 4175 19263 4209 19297
rect 4243 19263 4277 19297
rect 4311 19263 4345 19297
rect 4379 19263 4413 19297
rect 4447 19263 4481 19297
rect 4515 19263 4549 19297
rect 4583 19263 4617 19297
rect 4651 19263 4685 19297
rect 4719 19263 4753 19297
rect 4787 19263 4821 19297
rect 4855 19263 4889 19297
rect 4923 19263 4957 19297
rect 4991 19263 5025 19297
rect 5059 19263 5093 19297
rect 5127 19263 5161 19297
rect 5195 19263 5229 19297
rect 5263 19263 5297 19297
rect 5331 19263 5365 19297
rect 5399 19263 5433 19297
rect 5467 19263 5501 19297
rect 5535 19263 5569 19297
rect 5603 19263 5637 19297
rect 5671 19263 5705 19297
rect 5739 19263 5773 19297
rect 5807 19263 5841 19297
rect 5875 19263 5909 19297
rect 5943 19263 5977 19297
rect 6011 19263 6045 19297
rect 6079 19263 6113 19297
rect 6147 19263 6181 19297
rect 6215 19263 6249 19297
rect 6283 19263 6317 19297
rect 6351 19263 6385 19297
rect 6419 19263 6453 19297
rect 6487 19263 6521 19297
rect 6555 19263 6589 19297
rect 6623 19263 6657 19297
rect 6691 19263 6725 19297
rect 6759 19263 6793 19297
rect 6827 19263 6861 19297
rect 6895 19263 6929 19297
rect 6963 19263 6997 19297
rect 7031 19263 7065 19297
rect 7099 19263 7133 19297
rect 7167 19263 7201 19297
rect 7235 19263 7269 19297
rect 7303 19263 7337 19297
rect 7371 19263 7405 19297
rect 7439 19263 7473 19297
rect 7507 19263 7541 19297
rect 7575 19263 7609 19297
rect 7643 19263 7677 19297
rect 7711 19263 7745 19297
rect 7779 19263 7813 19297
rect 7847 19263 7881 19297
rect 7915 19263 7949 19297
rect 7983 19263 8017 19297
rect 8051 19263 8085 19297
rect 8119 19263 8153 19297
rect 8187 19263 8221 19297
rect 8255 19263 8289 19297
rect 8323 19263 8357 19297
rect 8391 19263 8425 19297
rect 8459 19263 8493 19297
rect 8527 19263 8561 19297
rect 8595 19263 8629 19297
rect 8663 19263 8697 19297
rect 8731 19263 8765 19297
rect 8799 19263 8833 19297
rect 8867 19263 8901 19297
rect 8935 19263 8969 19297
rect 9003 19263 9037 19297
rect 9071 19263 9105 19297
rect 9139 19263 9173 19297
rect 9207 19263 9241 19297
rect 9275 19263 9309 19297
rect 9343 19263 9377 19297
rect 9411 19263 9445 19297
rect 9479 19263 9513 19297
rect 9547 19263 9581 19297
rect 9615 19263 9649 19297
rect 9683 19263 9717 19297
rect 9751 19263 9785 19297
rect 9819 19263 9853 19297
rect 9887 19263 9921 19297
rect 9955 19263 9989 19297
rect 10023 19263 10057 19297
rect 10091 19263 10125 19297
rect 10159 19263 10193 19297
rect 10227 19263 10261 19297
rect 10295 19263 10329 19297
rect 10363 19263 10397 19297
rect 10431 19263 10465 19297
rect 10499 19263 10533 19297
rect 10567 19263 10601 19297
rect 10635 19263 10669 19297
rect 10703 19263 10737 19297
rect 10771 19263 10805 19297
rect 10839 19263 10873 19297
rect 10907 19263 10941 19297
rect 10975 19263 11009 19297
rect 11043 19263 11077 19297
rect 11111 19263 11145 19297
rect 11179 19263 11213 19297
rect 11247 19263 11281 19297
rect 11315 19263 11349 19297
rect 11383 19263 11417 19297
rect 11451 19263 11485 19297
rect 11519 19263 11553 19297
rect 11587 19263 11621 19297
rect 11655 19263 11689 19297
rect 11723 19263 11747 19297
rect 53 19225 11747 19263
rect 53 19191 77 19225
rect 111 19191 146 19225
rect 180 19191 215 19225
rect 249 19191 284 19225
rect 318 19191 353 19225
rect 387 19191 422 19225
rect 456 19191 491 19225
rect 525 19191 560 19225
rect 594 19191 629 19225
rect 663 19191 698 19225
rect 732 19191 767 19225
rect 801 19191 836 19225
rect 870 19191 905 19225
rect 939 19191 974 19225
rect 1008 19191 1043 19225
rect 1077 19191 1112 19225
rect 1146 19191 1181 19225
rect 1215 19191 1250 19225
rect 1284 19191 1319 19225
rect 1353 19191 1388 19225
rect 1422 19191 1457 19225
rect 1491 19191 1526 19225
rect 1560 19191 1595 19225
rect 1629 19191 1664 19225
rect 1698 19191 1733 19225
rect 1767 19191 1802 19225
rect 1836 19191 1871 19225
rect 1905 19191 1940 19225
rect 1974 19191 2009 19225
rect 2043 19191 2078 19225
rect 2112 19191 2147 19225
rect 2181 19191 2216 19225
rect 2250 19191 2285 19225
rect 2319 19191 2354 19225
rect 2388 19191 2423 19225
rect 2457 19191 2492 19225
rect 2526 19191 2561 19225
rect 2595 19191 2630 19225
rect 2664 19191 2699 19225
rect 2733 19191 2768 19225
rect 2802 19191 2837 19225
rect 2871 19191 2906 19225
rect 2940 19191 2975 19225
rect 3009 19191 3044 19225
rect 3078 19191 3113 19225
rect 3147 19191 3182 19225
rect 3216 19191 3251 19225
rect 3285 19191 3320 19225
rect 3354 19191 3389 19225
rect 3423 19191 3458 19225
rect 3492 19191 3527 19225
rect 3561 19191 3596 19225
rect 3630 19191 3665 19225
rect 3699 19191 3733 19225
rect 3767 19191 3801 19225
rect 3835 19191 3869 19225
rect 3903 19191 3937 19225
rect 3971 19191 4005 19225
rect 4039 19191 4073 19225
rect 4107 19191 4141 19225
rect 4175 19191 4209 19225
rect 4243 19191 4277 19225
rect 4311 19191 4345 19225
rect 4379 19191 4413 19225
rect 4447 19191 4481 19225
rect 4515 19191 4549 19225
rect 4583 19191 4617 19225
rect 4651 19191 4685 19225
rect 4719 19191 4753 19225
rect 4787 19191 4821 19225
rect 4855 19191 4889 19225
rect 4923 19191 4957 19225
rect 4991 19191 5025 19225
rect 5059 19191 5093 19225
rect 5127 19191 5161 19225
rect 5195 19191 5229 19225
rect 5263 19191 5297 19225
rect 5331 19191 5365 19225
rect 5399 19191 5433 19225
rect 5467 19191 5501 19225
rect 5535 19191 5569 19225
rect 5603 19191 5637 19225
rect 5671 19191 5705 19225
rect 5739 19191 5773 19225
rect 5807 19191 5841 19225
rect 5875 19191 5909 19225
rect 5943 19191 5977 19225
rect 6011 19191 6045 19225
rect 6079 19191 6113 19225
rect 6147 19191 6181 19225
rect 6215 19191 6249 19225
rect 6283 19191 6317 19225
rect 6351 19191 6385 19225
rect 6419 19191 6453 19225
rect 6487 19191 6521 19225
rect 6555 19191 6589 19225
rect 6623 19191 6657 19225
rect 6691 19191 6725 19225
rect 6759 19191 6793 19225
rect 6827 19191 6861 19225
rect 6895 19191 6929 19225
rect 6963 19191 6997 19225
rect 7031 19191 7065 19225
rect 7099 19191 7133 19225
rect 7167 19191 7201 19225
rect 7235 19191 7269 19225
rect 7303 19191 7337 19225
rect 7371 19191 7405 19225
rect 7439 19191 7473 19225
rect 7507 19191 7541 19225
rect 7575 19191 7609 19225
rect 7643 19191 7677 19225
rect 7711 19191 7745 19225
rect 7779 19191 7813 19225
rect 7847 19191 7881 19225
rect 7915 19191 7949 19225
rect 7983 19191 8017 19225
rect 8051 19191 8085 19225
rect 8119 19191 8153 19225
rect 8187 19191 8221 19225
rect 8255 19191 8289 19225
rect 8323 19191 8357 19225
rect 8391 19191 8425 19225
rect 8459 19191 8493 19225
rect 8527 19191 8561 19225
rect 8595 19191 8629 19225
rect 8663 19191 8697 19225
rect 8731 19191 8765 19225
rect 8799 19191 8833 19225
rect 8867 19191 8901 19225
rect 8935 19191 8969 19225
rect 9003 19191 9037 19225
rect 9071 19191 9105 19225
rect 9139 19191 9173 19225
rect 9207 19191 9241 19225
rect 9275 19191 9309 19225
rect 9343 19191 9377 19225
rect 9411 19191 9445 19225
rect 9479 19191 9513 19225
rect 9547 19191 9581 19225
rect 9615 19191 9649 19225
rect 9683 19191 9717 19225
rect 9751 19191 9785 19225
rect 9819 19191 9853 19225
rect 9887 19191 9921 19225
rect 9955 19191 9989 19225
rect 10023 19191 10057 19225
rect 10091 19191 10125 19225
rect 10159 19191 10193 19225
rect 10227 19191 10261 19225
rect 10295 19191 10329 19225
rect 10363 19191 10397 19225
rect 10431 19191 10465 19225
rect 10499 19191 10533 19225
rect 10567 19191 10601 19225
rect 10635 19191 10669 19225
rect 10703 19191 10737 19225
rect 10771 19191 10805 19225
rect 10839 19191 10873 19225
rect 10907 19191 10941 19225
rect 10975 19191 11009 19225
rect 11043 19191 11077 19225
rect 11111 19191 11145 19225
rect 11179 19191 11213 19225
rect 11247 19191 11281 19225
rect 11315 19191 11349 19225
rect 11383 19191 11417 19225
rect 11451 19191 11485 19225
rect 11519 19191 11553 19225
rect 11587 19191 11621 19225
rect 11655 19191 11689 19225
rect 11723 19191 11747 19225
rect 53 19153 11747 19191
rect 53 19119 77 19153
rect 111 19119 146 19153
rect 180 19119 215 19153
rect 249 19119 284 19153
rect 318 19119 353 19153
rect 387 19119 422 19153
rect 456 19119 491 19153
rect 525 19119 560 19153
rect 594 19119 629 19153
rect 663 19119 698 19153
rect 732 19119 767 19153
rect 801 19119 836 19153
rect 870 19119 905 19153
rect 939 19119 974 19153
rect 1008 19119 1043 19153
rect 1077 19119 1112 19153
rect 1146 19119 1181 19153
rect 1215 19119 1250 19153
rect 1284 19119 1319 19153
rect 1353 19119 1388 19153
rect 1422 19119 1457 19153
rect 1491 19119 1526 19153
rect 1560 19119 1595 19153
rect 1629 19119 1664 19153
rect 1698 19119 1733 19153
rect 1767 19119 1802 19153
rect 1836 19119 1871 19153
rect 1905 19119 1940 19153
rect 1974 19119 2009 19153
rect 2043 19119 2078 19153
rect 2112 19119 2147 19153
rect 2181 19119 2216 19153
rect 2250 19119 2285 19153
rect 2319 19119 2354 19153
rect 2388 19119 2423 19153
rect 2457 19119 2492 19153
rect 2526 19119 2561 19153
rect 2595 19119 2630 19153
rect 2664 19119 2699 19153
rect 2733 19119 2768 19153
rect 2802 19119 2837 19153
rect 2871 19119 2906 19153
rect 2940 19119 2975 19153
rect 3009 19119 3044 19153
rect 3078 19119 3113 19153
rect 3147 19119 3182 19153
rect 3216 19119 3251 19153
rect 3285 19119 3320 19153
rect 3354 19119 3389 19153
rect 3423 19119 3458 19153
rect 3492 19119 3527 19153
rect 3561 19119 3596 19153
rect 3630 19119 3665 19153
rect 3699 19119 3733 19153
rect 3767 19119 3801 19153
rect 3835 19119 3869 19153
rect 3903 19119 3937 19153
rect 3971 19119 4005 19153
rect 4039 19119 4073 19153
rect 4107 19119 4141 19153
rect 4175 19119 4209 19153
rect 4243 19119 4277 19153
rect 4311 19119 4345 19153
rect 4379 19119 4413 19153
rect 4447 19119 4481 19153
rect 4515 19119 4549 19153
rect 4583 19119 4617 19153
rect 4651 19119 4685 19153
rect 4719 19119 4753 19153
rect 4787 19119 4821 19153
rect 4855 19119 4889 19153
rect 4923 19119 4957 19153
rect 4991 19119 5025 19153
rect 5059 19119 5093 19153
rect 5127 19119 5161 19153
rect 5195 19119 5229 19153
rect 5263 19119 5297 19153
rect 5331 19119 5365 19153
rect 5399 19119 5433 19153
rect 5467 19119 5501 19153
rect 5535 19119 5569 19153
rect 5603 19119 5637 19153
rect 5671 19119 5705 19153
rect 5739 19119 5773 19153
rect 5807 19119 5841 19153
rect 5875 19119 5909 19153
rect 5943 19119 5977 19153
rect 6011 19119 6045 19153
rect 6079 19119 6113 19153
rect 6147 19119 6181 19153
rect 6215 19119 6249 19153
rect 6283 19119 6317 19153
rect 6351 19119 6385 19153
rect 6419 19119 6453 19153
rect 6487 19119 6521 19153
rect 6555 19119 6589 19153
rect 6623 19119 6657 19153
rect 6691 19119 6725 19153
rect 6759 19119 6793 19153
rect 6827 19119 6861 19153
rect 6895 19119 6929 19153
rect 6963 19119 6997 19153
rect 7031 19119 7065 19153
rect 7099 19119 7133 19153
rect 7167 19119 7201 19153
rect 7235 19119 7269 19153
rect 7303 19119 7337 19153
rect 7371 19119 7405 19153
rect 7439 19119 7473 19153
rect 7507 19119 7541 19153
rect 7575 19119 7609 19153
rect 7643 19119 7677 19153
rect 7711 19119 7745 19153
rect 7779 19119 7813 19153
rect 7847 19119 7881 19153
rect 7915 19119 7949 19153
rect 7983 19119 8017 19153
rect 8051 19119 8085 19153
rect 8119 19119 8153 19153
rect 8187 19119 8221 19153
rect 8255 19119 8289 19153
rect 8323 19119 8357 19153
rect 8391 19119 8425 19153
rect 8459 19119 8493 19153
rect 8527 19119 8561 19153
rect 8595 19119 8629 19153
rect 8663 19119 8697 19153
rect 8731 19119 8765 19153
rect 8799 19119 8833 19153
rect 8867 19119 8901 19153
rect 8935 19119 8969 19153
rect 9003 19119 9037 19153
rect 9071 19119 9105 19153
rect 9139 19119 9173 19153
rect 9207 19119 9241 19153
rect 9275 19119 9309 19153
rect 9343 19119 9377 19153
rect 9411 19119 9445 19153
rect 9479 19119 9513 19153
rect 9547 19119 9581 19153
rect 9615 19119 9649 19153
rect 9683 19119 9717 19153
rect 9751 19119 9785 19153
rect 9819 19119 9853 19153
rect 9887 19119 9921 19153
rect 9955 19119 9989 19153
rect 10023 19119 10057 19153
rect 10091 19119 10125 19153
rect 10159 19119 10193 19153
rect 10227 19119 10261 19153
rect 10295 19119 10329 19153
rect 10363 19119 10397 19153
rect 10431 19119 10465 19153
rect 10499 19119 10533 19153
rect 10567 19119 10601 19153
rect 10635 19119 10669 19153
rect 10703 19119 10737 19153
rect 10771 19119 10805 19153
rect 10839 19119 10873 19153
rect 10907 19119 10941 19153
rect 10975 19119 11009 19153
rect 11043 19119 11077 19153
rect 11111 19119 11145 19153
rect 11179 19119 11213 19153
rect 11247 19119 11281 19153
rect 11315 19119 11349 19153
rect 11383 19119 11417 19153
rect 11451 19119 11485 19153
rect 11519 19119 11553 19153
rect 11587 19119 11621 19153
rect 11655 19119 11689 19153
rect 11723 19119 11747 19153
rect 53 19081 11747 19119
rect 53 19047 77 19081
rect 111 19047 146 19081
rect 180 19047 215 19081
rect 249 19047 284 19081
rect 318 19047 353 19081
rect 387 19047 422 19081
rect 456 19047 491 19081
rect 525 19047 560 19081
rect 594 19047 629 19081
rect 663 19047 698 19081
rect 732 19047 767 19081
rect 801 19047 836 19081
rect 870 19047 905 19081
rect 939 19047 974 19081
rect 1008 19047 1043 19081
rect 1077 19047 1112 19081
rect 1146 19047 1181 19081
rect 1215 19047 1250 19081
rect 1284 19047 1319 19081
rect 1353 19047 1388 19081
rect 1422 19047 1457 19081
rect 1491 19047 1526 19081
rect 1560 19047 1595 19081
rect 1629 19047 1664 19081
rect 1698 19047 1733 19081
rect 1767 19047 1802 19081
rect 1836 19047 1871 19081
rect 1905 19047 1940 19081
rect 1974 19047 2009 19081
rect 2043 19047 2078 19081
rect 2112 19047 2147 19081
rect 2181 19047 2216 19081
rect 2250 19047 2285 19081
rect 2319 19047 2354 19081
rect 2388 19047 2423 19081
rect 2457 19047 2492 19081
rect 2526 19047 2561 19081
rect 2595 19047 2630 19081
rect 2664 19047 2699 19081
rect 2733 19047 2768 19081
rect 2802 19047 2837 19081
rect 2871 19047 2906 19081
rect 2940 19047 2975 19081
rect 3009 19047 3044 19081
rect 3078 19047 3113 19081
rect 3147 19047 3182 19081
rect 3216 19047 3251 19081
rect 3285 19047 3320 19081
rect 3354 19047 3389 19081
rect 3423 19047 3458 19081
rect 3492 19047 3527 19081
rect 3561 19047 3596 19081
rect 3630 19047 3665 19081
rect 3699 19047 3733 19081
rect 3767 19047 3801 19081
rect 3835 19047 3869 19081
rect 3903 19047 3937 19081
rect 3971 19047 4005 19081
rect 4039 19047 4073 19081
rect 4107 19047 4141 19081
rect 4175 19047 4209 19081
rect 4243 19047 4277 19081
rect 4311 19047 4345 19081
rect 4379 19047 4413 19081
rect 4447 19047 4481 19081
rect 4515 19047 4549 19081
rect 4583 19047 4617 19081
rect 4651 19047 4685 19081
rect 4719 19047 4753 19081
rect 4787 19047 4821 19081
rect 4855 19047 4889 19081
rect 4923 19047 4957 19081
rect 4991 19047 5025 19081
rect 5059 19047 5093 19081
rect 5127 19047 5161 19081
rect 5195 19047 5229 19081
rect 5263 19047 5297 19081
rect 5331 19047 5365 19081
rect 5399 19047 5433 19081
rect 5467 19047 5501 19081
rect 5535 19047 5569 19081
rect 5603 19047 5637 19081
rect 5671 19047 5705 19081
rect 5739 19047 5773 19081
rect 5807 19047 5841 19081
rect 5875 19047 5909 19081
rect 5943 19047 5977 19081
rect 6011 19047 6045 19081
rect 6079 19047 6113 19081
rect 6147 19047 6181 19081
rect 6215 19047 6249 19081
rect 6283 19047 6317 19081
rect 6351 19047 6385 19081
rect 6419 19047 6453 19081
rect 6487 19047 6521 19081
rect 6555 19047 6589 19081
rect 6623 19047 6657 19081
rect 6691 19047 6725 19081
rect 6759 19047 6793 19081
rect 6827 19047 6861 19081
rect 6895 19047 6929 19081
rect 6963 19047 6997 19081
rect 7031 19047 7065 19081
rect 7099 19047 7133 19081
rect 7167 19047 7201 19081
rect 7235 19047 7269 19081
rect 7303 19047 7337 19081
rect 7371 19047 7405 19081
rect 7439 19047 7473 19081
rect 7507 19047 7541 19081
rect 7575 19047 7609 19081
rect 7643 19047 7677 19081
rect 7711 19047 7745 19081
rect 7779 19047 7813 19081
rect 7847 19047 7881 19081
rect 7915 19047 7949 19081
rect 7983 19047 8017 19081
rect 8051 19047 8085 19081
rect 8119 19047 8153 19081
rect 8187 19047 8221 19081
rect 8255 19047 8289 19081
rect 8323 19047 8357 19081
rect 8391 19047 8425 19081
rect 8459 19047 8493 19081
rect 8527 19047 8561 19081
rect 8595 19047 8629 19081
rect 8663 19047 8697 19081
rect 8731 19047 8765 19081
rect 8799 19047 8833 19081
rect 8867 19047 8901 19081
rect 8935 19047 8969 19081
rect 9003 19047 9037 19081
rect 9071 19047 9105 19081
rect 9139 19047 9173 19081
rect 9207 19047 9241 19081
rect 9275 19047 9309 19081
rect 9343 19047 9377 19081
rect 9411 19047 9445 19081
rect 9479 19047 9513 19081
rect 9547 19047 9581 19081
rect 9615 19047 9649 19081
rect 9683 19047 9717 19081
rect 9751 19047 9785 19081
rect 9819 19047 9853 19081
rect 9887 19047 9921 19081
rect 9955 19047 9989 19081
rect 10023 19047 10057 19081
rect 10091 19047 10125 19081
rect 10159 19047 10193 19081
rect 10227 19047 10261 19081
rect 10295 19047 10329 19081
rect 10363 19047 10397 19081
rect 10431 19047 10465 19081
rect 10499 19047 10533 19081
rect 10567 19047 10601 19081
rect 10635 19047 10669 19081
rect 10703 19047 10737 19081
rect 10771 19047 10805 19081
rect 10839 19047 10873 19081
rect 10907 19047 10941 19081
rect 10975 19047 11009 19081
rect 11043 19047 11077 19081
rect 11111 19047 11145 19081
rect 11179 19047 11213 19081
rect 11247 19047 11281 19081
rect 11315 19047 11349 19081
rect 11383 19047 11417 19081
rect 11451 19047 11485 19081
rect 11519 19047 11553 19081
rect 11587 19047 11621 19081
rect 11655 19047 11689 19081
rect 11723 19047 11747 19081
rect 53 19009 11747 19047
rect 53 18975 77 19009
rect 111 18975 146 19009
rect 180 18975 215 19009
rect 249 18975 284 19009
rect 318 18975 353 19009
rect 387 18975 422 19009
rect 456 18975 491 19009
rect 525 18975 560 19009
rect 594 18975 629 19009
rect 663 18975 698 19009
rect 732 18975 767 19009
rect 801 18975 836 19009
rect 870 18975 905 19009
rect 939 18975 974 19009
rect 1008 18975 1043 19009
rect 1077 18975 1112 19009
rect 1146 18975 1181 19009
rect 1215 18975 1250 19009
rect 1284 18975 1319 19009
rect 1353 18975 1388 19009
rect 1422 18975 1457 19009
rect 1491 18975 1526 19009
rect 1560 18975 1595 19009
rect 1629 18975 1664 19009
rect 1698 18975 1733 19009
rect 1767 18975 1802 19009
rect 1836 18975 1871 19009
rect 1905 18975 1940 19009
rect 1974 18975 2009 19009
rect 2043 18975 2078 19009
rect 2112 18975 2147 19009
rect 2181 18975 2216 19009
rect 2250 18975 2285 19009
rect 2319 18975 2354 19009
rect 2388 18975 2423 19009
rect 2457 18975 2492 19009
rect 2526 18975 2561 19009
rect 2595 18975 2630 19009
rect 2664 18975 2699 19009
rect 2733 18975 2768 19009
rect 2802 18975 2837 19009
rect 2871 18975 2906 19009
rect 2940 18975 2975 19009
rect 3009 18975 3044 19009
rect 3078 18975 3113 19009
rect 3147 18975 3182 19009
rect 3216 18975 3251 19009
rect 3285 18975 3320 19009
rect 3354 18975 3389 19009
rect 3423 18975 3458 19009
rect 3492 18975 3527 19009
rect 3561 18975 3596 19009
rect 3630 18975 3665 19009
rect 3699 18975 3733 19009
rect 3767 18975 3801 19009
rect 3835 18975 3869 19009
rect 3903 18975 3937 19009
rect 3971 18975 4005 19009
rect 4039 18975 4073 19009
rect 4107 18975 4141 19009
rect 4175 18975 4209 19009
rect 4243 18975 4277 19009
rect 4311 18975 4345 19009
rect 4379 18975 4413 19009
rect 4447 18975 4481 19009
rect 4515 18975 4549 19009
rect 4583 18975 4617 19009
rect 4651 18975 4685 19009
rect 4719 18975 4753 19009
rect 4787 18975 4821 19009
rect 4855 18975 4889 19009
rect 4923 18975 4957 19009
rect 4991 18975 5025 19009
rect 5059 18975 5093 19009
rect 5127 18975 5161 19009
rect 5195 18975 5229 19009
rect 5263 18975 5297 19009
rect 5331 18975 5365 19009
rect 5399 18975 5433 19009
rect 5467 18975 5501 19009
rect 5535 18975 5569 19009
rect 5603 18975 5637 19009
rect 5671 18975 5705 19009
rect 5739 18975 5773 19009
rect 5807 18975 5841 19009
rect 5875 18975 5909 19009
rect 5943 18975 5977 19009
rect 6011 18975 6045 19009
rect 6079 18975 6113 19009
rect 6147 18975 6181 19009
rect 6215 18975 6249 19009
rect 6283 18975 6317 19009
rect 6351 18975 6385 19009
rect 6419 18975 6453 19009
rect 6487 18975 6521 19009
rect 6555 18975 6589 19009
rect 6623 18975 6657 19009
rect 6691 18975 6725 19009
rect 6759 18975 6793 19009
rect 6827 18975 6861 19009
rect 6895 18975 6929 19009
rect 6963 18975 6997 19009
rect 7031 18975 7065 19009
rect 7099 18975 7133 19009
rect 7167 18975 7201 19009
rect 7235 18975 7269 19009
rect 7303 18975 7337 19009
rect 7371 18975 7405 19009
rect 7439 18975 7473 19009
rect 7507 18975 7541 19009
rect 7575 18975 7609 19009
rect 7643 18975 7677 19009
rect 7711 18975 7745 19009
rect 7779 18975 7813 19009
rect 7847 18975 7881 19009
rect 7915 18975 7949 19009
rect 7983 18975 8017 19009
rect 8051 18975 8085 19009
rect 8119 18975 8153 19009
rect 8187 18975 8221 19009
rect 8255 18975 8289 19009
rect 8323 18975 8357 19009
rect 8391 18975 8425 19009
rect 8459 18975 8493 19009
rect 8527 18975 8561 19009
rect 8595 18975 8629 19009
rect 8663 18975 8697 19009
rect 8731 18975 8765 19009
rect 8799 18975 8833 19009
rect 8867 18975 8901 19009
rect 8935 18975 8969 19009
rect 9003 18975 9037 19009
rect 9071 18975 9105 19009
rect 9139 18975 9173 19009
rect 9207 18975 9241 19009
rect 9275 18975 9309 19009
rect 9343 18975 9377 19009
rect 9411 18975 9445 19009
rect 9479 18975 9513 19009
rect 9547 18975 9581 19009
rect 9615 18975 9649 19009
rect 9683 18975 9717 19009
rect 9751 18975 9785 19009
rect 9819 18975 9853 19009
rect 9887 18975 9921 19009
rect 9955 18975 9989 19009
rect 10023 18975 10057 19009
rect 10091 18975 10125 19009
rect 10159 18975 10193 19009
rect 10227 18975 10261 19009
rect 10295 18975 10329 19009
rect 10363 18975 10397 19009
rect 10431 18975 10465 19009
rect 10499 18975 10533 19009
rect 10567 18975 10601 19009
rect 10635 18975 10669 19009
rect 10703 18975 10737 19009
rect 10771 18975 10805 19009
rect 10839 18975 10873 19009
rect 10907 18975 10941 19009
rect 10975 18975 11009 19009
rect 11043 18975 11077 19009
rect 11111 18975 11145 19009
rect 11179 18975 11213 19009
rect 11247 18975 11281 19009
rect 11315 18975 11349 19009
rect 11383 18975 11417 19009
rect 11451 18975 11485 19009
rect 11519 18975 11553 19009
rect 11587 18975 11621 19009
rect 11655 18975 11689 19009
rect 11723 18975 11747 19009
rect 53 18915 11747 18975
rect 14460 19307 14484 19330
rect 14518 19307 14567 19341
rect 14601 19307 14650 19341
rect 14684 19307 14733 19341
rect 14767 19307 14816 19341
rect 14850 19307 14874 19341
rect 14460 19271 14874 19307
rect 14460 19237 14484 19271
rect 14518 19237 14567 19271
rect 14601 19237 14650 19271
rect 14684 19237 14733 19271
rect 14767 19237 14816 19271
rect 14850 19237 14874 19271
rect 14460 19201 14874 19237
rect 14460 19167 14484 19201
rect 14518 19167 14567 19201
rect 14601 19167 14650 19201
rect 14684 19167 14733 19201
rect 14767 19167 14816 19201
rect 14850 19167 14874 19201
rect 14460 19131 14874 19167
rect 14460 19097 14484 19131
rect 14518 19097 14567 19131
rect 14601 19097 14650 19131
rect 14684 19097 14733 19131
rect 14767 19097 14816 19131
rect 14850 19097 14874 19131
rect 14460 19061 14874 19097
rect 14460 19027 14484 19061
rect 14518 19027 14567 19061
rect 14601 19027 14650 19061
rect 14684 19027 14733 19061
rect 14767 19027 14816 19061
rect 14850 19027 14874 19061
rect 14460 18915 14874 19027
rect 53 18881 77 18915
rect 111 18881 146 18915
rect 180 18881 215 18915
rect 249 18881 284 18915
rect 318 18881 353 18915
rect 387 18881 422 18915
rect 456 18881 491 18915
rect 525 18881 560 18915
rect 594 18881 629 18915
rect 663 18881 698 18915
rect 732 18881 767 18915
rect 801 18881 836 18915
rect 870 18881 905 18915
rect 939 18881 974 18915
rect 1008 18881 1043 18915
rect 1077 18881 1112 18915
rect 1146 18881 1181 18915
rect 1215 18881 1250 18915
rect 1284 18881 1319 18915
rect 1353 18881 1388 18915
rect 1422 18881 1457 18915
rect 1491 18881 1526 18915
rect 1560 18881 1595 18915
rect 1629 18881 1664 18915
rect 1698 18881 1733 18915
rect 1767 18881 1802 18915
rect 1836 18881 1871 18915
rect 1905 18881 1940 18915
rect 1974 18881 2009 18915
rect 2043 18881 2078 18915
rect 2112 18881 2147 18915
rect 2181 18881 2216 18915
rect 2250 18881 2285 18915
rect 2319 18881 2354 18915
rect 2388 18881 2423 18915
rect 2457 18881 2492 18915
rect 2526 18881 2561 18915
rect 2595 18881 2630 18915
rect 2664 18881 2699 18915
rect 2733 18881 2768 18915
rect 2802 18881 2837 18915
rect 2871 18881 2906 18915
rect 2940 18881 2975 18915
rect 3009 18881 3044 18915
rect 3078 18881 3113 18915
rect 3147 18881 3182 18915
rect 3216 18881 3251 18915
rect 3285 18881 3320 18915
rect 3354 18881 3389 18915
rect 3423 18881 3458 18915
rect 3492 18881 3527 18915
rect 3561 18881 3596 18915
rect 53 18847 3596 18881
rect 53 18813 77 18847
rect 111 18813 146 18847
rect 180 18813 215 18847
rect 249 18813 284 18847
rect 318 18813 353 18847
rect 387 18813 422 18847
rect 456 18813 491 18847
rect 525 18813 560 18847
rect 594 18813 629 18847
rect 663 18813 698 18847
rect 732 18813 767 18847
rect 801 18813 836 18847
rect 870 18813 905 18847
rect 939 18813 974 18847
rect 1008 18813 1043 18847
rect 1077 18813 1112 18847
rect 1146 18813 1181 18847
rect 1215 18813 1250 18847
rect 1284 18813 1319 18847
rect 1353 18813 1388 18847
rect 1422 18813 1457 18847
rect 1491 18813 1526 18847
rect 1560 18813 1595 18847
rect 1629 18813 1664 18847
rect 1698 18813 1733 18847
rect 1767 18813 1802 18847
rect 1836 18813 1871 18847
rect 1905 18813 1940 18847
rect 1974 18813 2009 18847
rect 2043 18813 2078 18847
rect 2112 18813 2147 18847
rect 2181 18813 2216 18847
rect 2250 18813 2285 18847
rect 2319 18813 2354 18847
rect 2388 18813 2423 18847
rect 2457 18813 2492 18847
rect 2526 18813 2561 18847
rect 2595 18813 2630 18847
rect 2664 18813 2699 18847
rect 2733 18813 2768 18847
rect 2802 18813 2837 18847
rect 2871 18813 2906 18847
rect 2940 18813 2975 18847
rect 3009 18813 3044 18847
rect 3078 18813 3113 18847
rect 3147 18813 3182 18847
rect 3216 18813 3251 18847
rect 3285 18813 3320 18847
rect 3354 18813 3389 18847
rect 3423 18813 3458 18847
rect 3492 18813 3527 18847
rect 3561 18813 3596 18847
rect 53 18779 3596 18813
rect 53 18745 77 18779
rect 111 18745 146 18779
rect 180 18745 215 18779
rect 249 18745 284 18779
rect 318 18745 353 18779
rect 387 18745 422 18779
rect 456 18745 491 18779
rect 525 18745 560 18779
rect 594 18745 629 18779
rect 663 18745 698 18779
rect 732 18745 767 18779
rect 801 18745 836 18779
rect 870 18745 905 18779
rect 939 18745 974 18779
rect 1008 18745 1043 18779
rect 1077 18745 1112 18779
rect 1146 18745 1181 18779
rect 1215 18745 1250 18779
rect 1284 18745 1319 18779
rect 1353 18745 1388 18779
rect 1422 18745 1457 18779
rect 1491 18745 1526 18779
rect 1560 18745 1595 18779
rect 1629 18745 1664 18779
rect 1698 18745 1733 18779
rect 1767 18745 1802 18779
rect 1836 18745 1871 18779
rect 1905 18745 1940 18779
rect 1974 18745 2009 18779
rect 2043 18745 2078 18779
rect 2112 18745 2147 18779
rect 2181 18745 2216 18779
rect 2250 18745 2285 18779
rect 2319 18745 2354 18779
rect 2388 18745 2423 18779
rect 2457 18745 2492 18779
rect 2526 18745 2561 18779
rect 2595 18745 2630 18779
rect 2664 18745 2699 18779
rect 2733 18745 2768 18779
rect 2802 18745 2837 18779
rect 2871 18745 2906 18779
rect 2940 18745 2975 18779
rect 3009 18745 3044 18779
rect 3078 18745 3113 18779
rect 3147 18745 3182 18779
rect 3216 18745 3251 18779
rect 3285 18745 3320 18779
rect 3354 18745 3389 18779
rect 3423 18745 3458 18779
rect 3492 18745 3527 18779
rect 3561 18745 3596 18779
rect 53 18711 3596 18745
rect 53 18677 77 18711
rect 111 18677 146 18711
rect 180 18677 215 18711
rect 249 18677 284 18711
rect 318 18677 353 18711
rect 387 18677 422 18711
rect 456 18677 491 18711
rect 525 18677 560 18711
rect 594 18677 629 18711
rect 663 18677 698 18711
rect 732 18677 767 18711
rect 801 18677 836 18711
rect 870 18677 905 18711
rect 939 18677 974 18711
rect 1008 18677 1043 18711
rect 1077 18677 1112 18711
rect 1146 18677 1181 18711
rect 1215 18677 1250 18711
rect 1284 18677 1319 18711
rect 1353 18677 1388 18711
rect 1422 18677 1457 18711
rect 1491 18677 1526 18711
rect 1560 18677 1595 18711
rect 1629 18677 1664 18711
rect 1698 18677 1733 18711
rect 1767 18677 1802 18711
rect 1836 18677 1871 18711
rect 1905 18677 1940 18711
rect 1974 18677 2009 18711
rect 2043 18677 2078 18711
rect 2112 18677 2147 18711
rect 2181 18677 2216 18711
rect 2250 18677 2285 18711
rect 2319 18677 2354 18711
rect 2388 18677 2423 18711
rect 2457 18677 2492 18711
rect 2526 18677 2561 18711
rect 2595 18677 2630 18711
rect 2664 18677 2699 18711
rect 2733 18677 2768 18711
rect 2802 18677 2837 18711
rect 2871 18677 2906 18711
rect 2940 18677 2975 18711
rect 3009 18677 3044 18711
rect 3078 18677 3113 18711
rect 3147 18677 3182 18711
rect 3216 18677 3251 18711
rect 3285 18677 3320 18711
rect 3354 18677 3389 18711
rect 3423 18677 3458 18711
rect 3492 18677 3527 18711
rect 3561 18677 3596 18711
rect 14850 18677 14874 18915
rect 53 18621 14874 18677
rect 197 18589 14772 18621
rect 197 18555 221 18589
rect 255 18555 290 18589
rect 324 18555 359 18589
rect 393 18555 427 18589
rect 461 18555 495 18589
rect 529 18555 563 18589
rect 597 18555 631 18589
rect 665 18555 699 18589
rect 733 18555 767 18589
rect 801 18555 835 18589
rect 869 18555 903 18589
rect 937 18555 971 18589
rect 1005 18555 1039 18589
rect 1073 18555 1107 18589
rect 1141 18555 1175 18589
rect 1209 18555 1243 18589
rect 1277 18555 1311 18589
rect 1345 18555 1379 18589
rect 1413 18555 1447 18589
rect 1481 18555 1515 18589
rect 1549 18555 1583 18589
rect 1617 18555 1651 18589
rect 1685 18555 1719 18589
rect 1753 18555 1787 18589
rect 1821 18555 1855 18589
rect 1889 18555 1923 18589
rect 1957 18555 1991 18589
rect 2025 18555 2059 18589
rect 2093 18555 2127 18589
rect 2161 18555 2195 18589
rect 2229 18555 2263 18589
rect 2297 18555 2331 18589
rect 2365 18555 2399 18589
rect 2433 18555 2467 18589
rect 2501 18555 2535 18589
rect 2569 18555 2603 18589
rect 2637 18555 2671 18589
rect 2705 18555 2739 18589
rect 2773 18555 2807 18589
rect 2841 18555 2875 18589
rect 2909 18555 2943 18589
rect 2977 18555 3011 18589
rect 3045 18555 3079 18589
rect 3113 18555 3147 18589
rect 3181 18555 3215 18589
rect 3249 18555 3283 18589
rect 3317 18555 3351 18589
rect 3385 18555 3419 18589
rect 3453 18555 3487 18589
rect 3521 18555 3555 18589
rect 3589 18555 3623 18589
rect 3657 18555 3691 18589
rect 3725 18555 3759 18589
rect 3793 18555 3827 18589
rect 3861 18555 3895 18589
rect 3929 18555 3963 18589
rect 3997 18555 4031 18589
rect 4065 18555 4099 18589
rect 4133 18555 4167 18589
rect 4201 18555 4235 18589
rect 4269 18555 4303 18589
rect 4337 18555 4371 18589
rect 4405 18555 4439 18589
rect 4473 18555 4507 18589
rect 4541 18555 4575 18589
rect 4609 18555 4643 18589
rect 4677 18555 4711 18589
rect 4745 18555 4779 18589
rect 4813 18555 4847 18589
rect 4881 18555 4915 18589
rect 4949 18555 4983 18589
rect 5017 18555 5051 18589
rect 5085 18555 5119 18589
rect 5153 18555 5187 18589
rect 5221 18555 5255 18589
rect 5289 18555 5323 18589
rect 5357 18555 5391 18589
rect 5425 18555 5459 18589
rect 5493 18555 5527 18589
rect 5561 18555 5595 18589
rect 5629 18555 5663 18589
rect 5697 18555 5731 18589
rect 5765 18555 5799 18589
rect 5833 18555 5867 18589
rect 5901 18555 5935 18589
rect 5969 18555 6003 18589
rect 6037 18555 6071 18589
rect 6105 18555 6139 18589
rect 6173 18555 6207 18589
rect 6241 18555 6275 18589
rect 6309 18555 6343 18589
rect 6377 18555 6411 18589
rect 6445 18555 6479 18589
rect 6513 18555 6547 18589
rect 6581 18555 6615 18589
rect 6649 18555 6683 18589
rect 6717 18555 6751 18589
rect 6785 18555 6819 18589
rect 6853 18555 6887 18589
rect 6921 18555 6955 18589
rect 6989 18555 7023 18589
rect 7057 18555 7091 18589
rect 7125 18555 7159 18589
rect 7193 18555 7227 18589
rect 7261 18555 7295 18589
rect 7329 18555 7363 18589
rect 7397 18555 7431 18589
rect 7465 18555 7499 18589
rect 7533 18555 7567 18589
rect 7601 18555 7635 18589
rect 7669 18555 7703 18589
rect 7737 18555 7771 18589
rect 7805 18555 7839 18589
rect 7873 18555 7907 18589
rect 7941 18555 7975 18589
rect 8009 18555 8043 18589
rect 8077 18555 8111 18589
rect 8145 18555 8179 18589
rect 8213 18555 8247 18589
rect 8281 18555 8315 18589
rect 8349 18555 8383 18589
rect 8417 18555 8451 18589
rect 8485 18555 8519 18589
rect 8553 18555 8587 18589
rect 8621 18555 8655 18589
rect 8689 18555 8723 18589
rect 8757 18555 8791 18589
rect 8825 18555 8859 18589
rect 8893 18555 8927 18589
rect 8961 18555 8995 18589
rect 9029 18555 9063 18589
rect 9097 18555 9131 18589
rect 9165 18555 9199 18589
rect 9233 18555 9267 18589
rect 9301 18555 9335 18589
rect 9369 18555 9403 18589
rect 9437 18555 9471 18589
rect 9505 18555 9539 18589
rect 9573 18555 9607 18589
rect 9641 18555 9675 18589
rect 9709 18555 9743 18589
rect 9777 18555 9811 18589
rect 9845 18555 9879 18589
rect 9913 18555 9947 18589
rect 9981 18555 10015 18589
rect 10049 18555 10083 18589
rect 10117 18555 10151 18589
rect 10185 18555 10219 18589
rect 10253 18555 10287 18589
rect 10321 18555 10355 18589
rect 10389 18555 10423 18589
rect 10457 18555 10491 18589
rect 10525 18555 10559 18589
rect 10593 18555 10627 18589
rect 10661 18555 10695 18589
rect 10729 18555 10763 18589
rect 10797 18555 10831 18589
rect 10865 18555 10899 18589
rect 10933 18555 10967 18589
rect 11001 18555 11035 18589
rect 11069 18555 11103 18589
rect 11137 18555 11171 18589
rect 11205 18555 11239 18589
rect 11273 18555 11307 18589
rect 11341 18555 11375 18589
rect 11409 18555 11443 18589
rect 11477 18555 11511 18589
rect 11545 18555 11579 18589
rect 11613 18555 11647 18589
rect 11681 18555 11715 18589
rect 11749 18555 11783 18589
rect 11817 18555 11851 18589
rect 11885 18555 11919 18589
rect 11953 18555 11987 18589
rect 12021 18555 12055 18589
rect 12089 18555 12123 18589
rect 12157 18555 12191 18589
rect 12225 18555 12259 18589
rect 12293 18555 12327 18589
rect 12361 18555 12395 18589
rect 12429 18555 12463 18589
rect 12497 18555 12531 18589
rect 12565 18555 12599 18589
rect 12633 18555 12667 18589
rect 12701 18555 12735 18589
rect 12769 18555 12803 18589
rect 12837 18555 12871 18589
rect 12905 18555 12939 18589
rect 12973 18555 13007 18589
rect 13041 18555 13075 18589
rect 13109 18555 13143 18589
rect 13177 18555 13211 18589
rect 13245 18555 13279 18589
rect 13313 18555 13347 18589
rect 13381 18555 13415 18589
rect 13449 18555 13483 18589
rect 13517 18555 13551 18589
rect 13585 18555 13619 18589
rect 13653 18555 13687 18589
rect 13721 18555 13755 18589
rect 13789 18555 13823 18589
rect 13857 18555 13891 18589
rect 13925 18555 13959 18589
rect 13993 18555 14027 18589
rect 14061 18555 14095 18589
rect 14129 18555 14163 18589
rect 14197 18555 14231 18589
rect 14265 18555 14299 18589
rect 14333 18555 14367 18589
rect 14401 18555 14435 18589
rect 14469 18555 14503 18589
rect 14537 18555 14571 18589
rect 14605 18555 14639 18589
rect 14673 18555 14707 18589
rect 14741 18555 14772 18589
rect 197 18519 14772 18555
rect 197 18485 221 18519
rect 255 18485 290 18519
rect 324 18485 359 18519
rect 393 18485 427 18519
rect 461 18485 495 18519
rect 529 18485 563 18519
rect 597 18485 631 18519
rect 665 18485 699 18519
rect 733 18485 767 18519
rect 801 18485 835 18519
rect 869 18485 903 18519
rect 937 18485 971 18519
rect 1005 18485 1039 18519
rect 1073 18485 1107 18519
rect 1141 18485 1175 18519
rect 1209 18485 1243 18519
rect 1277 18485 1311 18519
rect 1345 18485 1379 18519
rect 1413 18485 1447 18519
rect 1481 18485 1515 18519
rect 1549 18485 1583 18519
rect 1617 18485 1651 18519
rect 1685 18485 1719 18519
rect 1753 18485 1787 18519
rect 1821 18485 1855 18519
rect 1889 18485 1923 18519
rect 1957 18485 1991 18519
rect 2025 18485 2059 18519
rect 2093 18485 2127 18519
rect 2161 18485 2195 18519
rect 2229 18485 2263 18519
rect 2297 18485 2331 18519
rect 2365 18485 2399 18519
rect 2433 18485 2467 18519
rect 2501 18485 2535 18519
rect 2569 18485 2603 18519
rect 2637 18485 2671 18519
rect 2705 18485 2739 18519
rect 2773 18485 2807 18519
rect 2841 18485 2875 18519
rect 2909 18485 2943 18519
rect 2977 18485 3011 18519
rect 3045 18485 3079 18519
rect 3113 18485 3147 18519
rect 3181 18485 3215 18519
rect 3249 18485 3283 18519
rect 3317 18485 3351 18519
rect 3385 18485 3419 18519
rect 3453 18485 3487 18519
rect 3521 18485 3555 18519
rect 3589 18485 3623 18519
rect 3657 18485 3691 18519
rect 3725 18485 3759 18519
rect 3793 18485 3827 18519
rect 3861 18485 3895 18519
rect 3929 18485 3963 18519
rect 3997 18485 4031 18519
rect 4065 18485 4099 18519
rect 4133 18485 4167 18519
rect 4201 18485 4235 18519
rect 4269 18485 4303 18519
rect 4337 18485 4371 18519
rect 4405 18485 4439 18519
rect 4473 18485 4507 18519
rect 4541 18485 4575 18519
rect 4609 18485 4643 18519
rect 4677 18485 4711 18519
rect 4745 18485 4779 18519
rect 4813 18485 4847 18519
rect 4881 18485 4915 18519
rect 4949 18485 4983 18519
rect 5017 18485 5051 18519
rect 5085 18485 5119 18519
rect 5153 18485 5187 18519
rect 5221 18485 5255 18519
rect 5289 18485 5323 18519
rect 5357 18485 5391 18519
rect 5425 18485 5459 18519
rect 5493 18485 5527 18519
rect 5561 18485 5595 18519
rect 5629 18485 5663 18519
rect 5697 18485 5731 18519
rect 5765 18485 5799 18519
rect 5833 18485 5867 18519
rect 5901 18485 5935 18519
rect 5969 18485 6003 18519
rect 6037 18485 6071 18519
rect 6105 18485 6139 18519
rect 6173 18485 6207 18519
rect 6241 18485 6275 18519
rect 6309 18485 6343 18519
rect 6377 18485 6411 18519
rect 6445 18485 6479 18519
rect 6513 18485 6547 18519
rect 6581 18485 6615 18519
rect 6649 18485 6683 18519
rect 6717 18485 6751 18519
rect 6785 18485 6819 18519
rect 6853 18485 6887 18519
rect 6921 18485 6955 18519
rect 6989 18485 7023 18519
rect 7057 18485 7091 18519
rect 7125 18485 7159 18519
rect 7193 18485 7227 18519
rect 7261 18485 7295 18519
rect 7329 18485 7363 18519
rect 7397 18485 7431 18519
rect 7465 18485 7499 18519
rect 7533 18485 7567 18519
rect 7601 18485 7635 18519
rect 7669 18485 7703 18519
rect 7737 18485 7771 18519
rect 7805 18485 7839 18519
rect 7873 18485 7907 18519
rect 7941 18485 7975 18519
rect 8009 18485 8043 18519
rect 8077 18485 8111 18519
rect 8145 18485 8179 18519
rect 8213 18485 8247 18519
rect 8281 18485 8315 18519
rect 8349 18485 8383 18519
rect 8417 18485 8451 18519
rect 8485 18485 8519 18519
rect 8553 18485 8587 18519
rect 8621 18485 8655 18519
rect 8689 18485 8723 18519
rect 8757 18485 8791 18519
rect 8825 18485 8859 18519
rect 8893 18485 8927 18519
rect 8961 18485 8995 18519
rect 9029 18485 9063 18519
rect 9097 18485 9131 18519
rect 9165 18485 9199 18519
rect 9233 18485 9267 18519
rect 9301 18485 9335 18519
rect 9369 18485 9403 18519
rect 9437 18485 9471 18519
rect 9505 18485 9539 18519
rect 9573 18485 9607 18519
rect 9641 18485 9675 18519
rect 9709 18485 9743 18519
rect 9777 18485 9811 18519
rect 9845 18485 9879 18519
rect 9913 18485 9947 18519
rect 9981 18485 10015 18519
rect 10049 18485 10083 18519
rect 10117 18485 10151 18519
rect 10185 18485 10219 18519
rect 10253 18485 10287 18519
rect 10321 18485 10355 18519
rect 10389 18485 10423 18519
rect 10457 18485 10491 18519
rect 10525 18485 10559 18519
rect 10593 18485 10627 18519
rect 10661 18485 10695 18519
rect 10729 18485 10763 18519
rect 10797 18485 10831 18519
rect 10865 18485 10899 18519
rect 10933 18485 10967 18519
rect 11001 18485 11035 18519
rect 11069 18485 11103 18519
rect 11137 18485 11171 18519
rect 11205 18485 11239 18519
rect 11273 18485 11307 18519
rect 11341 18485 11375 18519
rect 11409 18485 11443 18519
rect 11477 18485 11511 18519
rect 11545 18485 11579 18519
rect 11613 18485 11647 18519
rect 11681 18485 11715 18519
rect 11749 18485 11783 18519
rect 11817 18485 11851 18519
rect 11885 18485 11919 18519
rect 11953 18485 11987 18519
rect 12021 18485 12055 18519
rect 12089 18485 12123 18519
rect 12157 18485 12191 18519
rect 12225 18485 12259 18519
rect 12293 18485 12327 18519
rect 12361 18485 12395 18519
rect 12429 18485 12463 18519
rect 12497 18485 12531 18519
rect 12565 18485 12599 18519
rect 12633 18485 12667 18519
rect 12701 18485 12735 18519
rect 12769 18485 12803 18519
rect 12837 18485 12871 18519
rect 12905 18485 12939 18519
rect 12973 18485 13007 18519
rect 13041 18485 13075 18519
rect 13109 18485 13143 18519
rect 13177 18485 13211 18519
rect 13245 18485 13279 18519
rect 13313 18485 13347 18519
rect 13381 18485 13415 18519
rect 13449 18485 13483 18519
rect 13517 18485 13551 18519
rect 13585 18485 13619 18519
rect 13653 18485 13687 18519
rect 13721 18485 13755 18519
rect 13789 18485 13823 18519
rect 13857 18485 13891 18519
rect 13925 18485 13959 18519
rect 13993 18485 14027 18519
rect 14061 18485 14095 18519
rect 14129 18485 14163 18519
rect 14197 18485 14231 18519
rect 14265 18485 14299 18519
rect 14333 18485 14367 18519
rect 14401 18485 14435 18519
rect 14469 18485 14503 18519
rect 14537 18485 14571 18519
rect 14605 18485 14639 18519
rect 14673 18485 14707 18519
rect 14741 18485 14772 18519
rect 197 18449 14772 18485
rect 197 18415 221 18449
rect 255 18415 290 18449
rect 324 18415 359 18449
rect 393 18415 427 18449
rect 461 18415 495 18449
rect 529 18415 563 18449
rect 597 18415 631 18449
rect 665 18415 699 18449
rect 733 18415 767 18449
rect 801 18415 835 18449
rect 869 18415 903 18449
rect 937 18415 971 18449
rect 1005 18415 1039 18449
rect 1073 18415 1107 18449
rect 1141 18415 1175 18449
rect 1209 18415 1243 18449
rect 1277 18415 1311 18449
rect 1345 18415 1379 18449
rect 1413 18415 1447 18449
rect 1481 18415 1515 18449
rect 1549 18415 1583 18449
rect 1617 18415 1651 18449
rect 1685 18415 1719 18449
rect 1753 18415 1787 18449
rect 1821 18415 1855 18449
rect 1889 18415 1923 18449
rect 1957 18415 1991 18449
rect 2025 18415 2059 18449
rect 2093 18415 2127 18449
rect 2161 18415 2195 18449
rect 2229 18415 2263 18449
rect 2297 18415 2331 18449
rect 2365 18415 2399 18449
rect 2433 18415 2467 18449
rect 2501 18415 2535 18449
rect 2569 18415 2603 18449
rect 2637 18415 2671 18449
rect 2705 18415 2739 18449
rect 2773 18415 2807 18449
rect 2841 18415 2875 18449
rect 2909 18415 2943 18449
rect 2977 18415 3011 18449
rect 3045 18415 3079 18449
rect 3113 18415 3147 18449
rect 3181 18415 3215 18449
rect 3249 18415 3283 18449
rect 3317 18415 3351 18449
rect 3385 18415 3419 18449
rect 3453 18415 3487 18449
rect 3521 18415 3555 18449
rect 3589 18415 3623 18449
rect 3657 18415 3691 18449
rect 3725 18415 3759 18449
rect 3793 18415 3827 18449
rect 3861 18415 3895 18449
rect 3929 18415 3963 18449
rect 3997 18415 4031 18449
rect 4065 18415 4099 18449
rect 4133 18415 4167 18449
rect 4201 18415 4235 18449
rect 4269 18415 4303 18449
rect 4337 18415 4371 18449
rect 4405 18415 4439 18449
rect 4473 18415 4507 18449
rect 4541 18415 4575 18449
rect 4609 18415 4643 18449
rect 4677 18415 4711 18449
rect 4745 18415 4779 18449
rect 4813 18415 4847 18449
rect 4881 18415 4915 18449
rect 4949 18415 4983 18449
rect 5017 18415 5051 18449
rect 5085 18415 5119 18449
rect 5153 18415 5187 18449
rect 5221 18415 5255 18449
rect 5289 18415 5323 18449
rect 5357 18415 5391 18449
rect 5425 18415 5459 18449
rect 5493 18415 5527 18449
rect 5561 18415 5595 18449
rect 5629 18415 5663 18449
rect 5697 18415 5731 18449
rect 5765 18415 5799 18449
rect 5833 18415 5867 18449
rect 5901 18415 5935 18449
rect 5969 18415 6003 18449
rect 6037 18415 6071 18449
rect 6105 18415 6139 18449
rect 6173 18415 6207 18449
rect 6241 18415 6275 18449
rect 6309 18415 6343 18449
rect 6377 18415 6411 18449
rect 6445 18415 6479 18449
rect 6513 18415 6547 18449
rect 6581 18415 6615 18449
rect 6649 18415 6683 18449
rect 6717 18415 6751 18449
rect 6785 18415 6819 18449
rect 6853 18415 6887 18449
rect 6921 18415 6955 18449
rect 6989 18415 7023 18449
rect 7057 18415 7091 18449
rect 7125 18415 7159 18449
rect 7193 18415 7227 18449
rect 7261 18415 7295 18449
rect 7329 18415 7363 18449
rect 7397 18415 7431 18449
rect 7465 18415 7499 18449
rect 7533 18415 7567 18449
rect 7601 18415 7635 18449
rect 7669 18415 7703 18449
rect 7737 18415 7771 18449
rect 7805 18415 7839 18449
rect 7873 18415 7907 18449
rect 7941 18415 7975 18449
rect 8009 18415 8043 18449
rect 8077 18415 8111 18449
rect 8145 18415 8179 18449
rect 8213 18415 8247 18449
rect 8281 18415 8315 18449
rect 8349 18415 8383 18449
rect 8417 18415 8451 18449
rect 8485 18415 8519 18449
rect 8553 18415 8587 18449
rect 8621 18415 8655 18449
rect 8689 18415 8723 18449
rect 8757 18415 8791 18449
rect 8825 18415 8859 18449
rect 8893 18415 8927 18449
rect 8961 18415 8995 18449
rect 9029 18415 9063 18449
rect 9097 18415 9131 18449
rect 9165 18415 9199 18449
rect 9233 18415 9267 18449
rect 9301 18415 9335 18449
rect 9369 18415 9403 18449
rect 9437 18415 9471 18449
rect 9505 18415 9539 18449
rect 9573 18415 9607 18449
rect 9641 18415 9675 18449
rect 9709 18415 9743 18449
rect 9777 18415 9811 18449
rect 9845 18415 9879 18449
rect 9913 18415 9947 18449
rect 9981 18415 10015 18449
rect 10049 18415 10083 18449
rect 10117 18415 10151 18449
rect 10185 18415 10219 18449
rect 10253 18415 10287 18449
rect 10321 18415 10355 18449
rect 10389 18415 10423 18449
rect 10457 18415 10491 18449
rect 10525 18415 10559 18449
rect 10593 18415 10627 18449
rect 10661 18415 10695 18449
rect 10729 18415 10763 18449
rect 10797 18415 10831 18449
rect 10865 18415 10899 18449
rect 10933 18415 10967 18449
rect 11001 18415 11035 18449
rect 11069 18415 11103 18449
rect 11137 18415 11171 18449
rect 11205 18415 11239 18449
rect 11273 18415 11307 18449
rect 11341 18415 11375 18449
rect 11409 18415 11443 18449
rect 11477 18415 11511 18449
rect 11545 18415 11579 18449
rect 11613 18415 11647 18449
rect 11681 18415 11715 18449
rect 11749 18415 11783 18449
rect 11817 18415 11851 18449
rect 11885 18415 11919 18449
rect 11953 18415 11987 18449
rect 12021 18415 12055 18449
rect 12089 18415 12123 18449
rect 12157 18415 12191 18449
rect 12225 18415 12259 18449
rect 12293 18415 12327 18449
rect 12361 18415 12395 18449
rect 12429 18415 12463 18449
rect 12497 18415 12531 18449
rect 12565 18415 12599 18449
rect 12633 18415 12667 18449
rect 12701 18415 12735 18449
rect 12769 18415 12803 18449
rect 12837 18415 12871 18449
rect 12905 18415 12939 18449
rect 12973 18415 13007 18449
rect 13041 18415 13075 18449
rect 13109 18415 13143 18449
rect 13177 18415 13211 18449
rect 13245 18415 13279 18449
rect 13313 18415 13347 18449
rect 13381 18415 13415 18449
rect 13449 18415 13483 18449
rect 13517 18415 13551 18449
rect 13585 18415 13619 18449
rect 13653 18415 13687 18449
rect 13721 18415 13755 18449
rect 13789 18415 13823 18449
rect 13857 18415 13891 18449
rect 13925 18415 13959 18449
rect 13993 18415 14027 18449
rect 14061 18415 14095 18449
rect 14129 18415 14163 18449
rect 14197 18415 14231 18449
rect 14265 18415 14299 18449
rect 14333 18415 14367 18449
rect 14401 18415 14435 18449
rect 14469 18415 14503 18449
rect 14537 18415 14571 18449
rect 14605 18415 14639 18449
rect 14673 18415 14707 18449
rect 14741 18415 14772 18449
rect 197 18379 14772 18415
rect 197 18345 221 18379
rect 255 18345 290 18379
rect 324 18345 359 18379
rect 393 18345 427 18379
rect 461 18345 495 18379
rect 529 18345 563 18379
rect 597 18345 631 18379
rect 665 18345 699 18379
rect 733 18345 767 18379
rect 801 18345 835 18379
rect 869 18345 903 18379
rect 937 18345 971 18379
rect 1005 18345 1039 18379
rect 1073 18345 1107 18379
rect 1141 18345 1175 18379
rect 1209 18345 1243 18379
rect 1277 18345 1311 18379
rect 1345 18345 1379 18379
rect 1413 18345 1447 18379
rect 1481 18345 1515 18379
rect 1549 18345 1583 18379
rect 1617 18345 1651 18379
rect 1685 18345 1719 18379
rect 1753 18345 1787 18379
rect 1821 18345 1855 18379
rect 1889 18345 1923 18379
rect 1957 18345 1991 18379
rect 2025 18345 2059 18379
rect 2093 18345 2127 18379
rect 2161 18345 2195 18379
rect 2229 18345 2263 18379
rect 2297 18345 2331 18379
rect 2365 18345 2399 18379
rect 2433 18345 2467 18379
rect 2501 18345 2535 18379
rect 2569 18345 2603 18379
rect 2637 18345 2671 18379
rect 2705 18345 2739 18379
rect 2773 18345 2807 18379
rect 2841 18345 2875 18379
rect 2909 18345 2943 18379
rect 2977 18345 3011 18379
rect 3045 18345 3079 18379
rect 3113 18345 3147 18379
rect 3181 18345 3215 18379
rect 3249 18345 3283 18379
rect 3317 18345 3351 18379
rect 3385 18345 3419 18379
rect 3453 18345 3487 18379
rect 3521 18345 3555 18379
rect 3589 18345 3623 18379
rect 3657 18345 3691 18379
rect 3725 18345 3759 18379
rect 3793 18345 3827 18379
rect 3861 18345 3895 18379
rect 3929 18345 3963 18379
rect 3997 18345 4031 18379
rect 4065 18345 4099 18379
rect 4133 18345 4167 18379
rect 4201 18345 4235 18379
rect 4269 18345 4303 18379
rect 4337 18345 4371 18379
rect 4405 18345 4439 18379
rect 4473 18345 4507 18379
rect 4541 18345 4575 18379
rect 4609 18345 4643 18379
rect 4677 18345 4711 18379
rect 4745 18345 4779 18379
rect 4813 18345 4847 18379
rect 4881 18345 4915 18379
rect 4949 18345 4983 18379
rect 5017 18345 5051 18379
rect 5085 18345 5119 18379
rect 5153 18345 5187 18379
rect 5221 18345 5255 18379
rect 5289 18345 5323 18379
rect 5357 18345 5391 18379
rect 5425 18345 5459 18379
rect 5493 18345 5527 18379
rect 5561 18345 5595 18379
rect 5629 18345 5663 18379
rect 5697 18345 5731 18379
rect 5765 18345 5799 18379
rect 5833 18345 5867 18379
rect 5901 18345 5935 18379
rect 5969 18345 6003 18379
rect 6037 18345 6071 18379
rect 6105 18345 6139 18379
rect 6173 18345 6207 18379
rect 6241 18345 6275 18379
rect 6309 18345 6343 18379
rect 6377 18345 6411 18379
rect 6445 18345 6479 18379
rect 6513 18345 6547 18379
rect 6581 18345 6615 18379
rect 6649 18345 6683 18379
rect 6717 18345 6751 18379
rect 6785 18345 6819 18379
rect 6853 18345 6887 18379
rect 6921 18345 6955 18379
rect 6989 18345 7023 18379
rect 7057 18345 7091 18379
rect 7125 18345 7159 18379
rect 7193 18345 7227 18379
rect 7261 18345 7295 18379
rect 7329 18345 7363 18379
rect 7397 18345 7431 18379
rect 7465 18345 7499 18379
rect 7533 18345 7567 18379
rect 7601 18345 7635 18379
rect 7669 18345 7703 18379
rect 7737 18345 7771 18379
rect 7805 18345 7839 18379
rect 7873 18345 7907 18379
rect 7941 18345 7975 18379
rect 8009 18345 8043 18379
rect 8077 18345 8111 18379
rect 8145 18345 8179 18379
rect 8213 18345 8247 18379
rect 8281 18345 8315 18379
rect 8349 18345 8383 18379
rect 8417 18345 8451 18379
rect 8485 18345 8519 18379
rect 8553 18345 8587 18379
rect 8621 18345 8655 18379
rect 8689 18345 8723 18379
rect 8757 18345 8791 18379
rect 8825 18345 8859 18379
rect 8893 18345 8927 18379
rect 8961 18345 8995 18379
rect 9029 18345 9063 18379
rect 9097 18345 9131 18379
rect 9165 18345 9199 18379
rect 9233 18345 9267 18379
rect 9301 18345 9335 18379
rect 9369 18345 9403 18379
rect 9437 18345 9471 18379
rect 9505 18345 9539 18379
rect 9573 18345 9607 18379
rect 9641 18345 9675 18379
rect 9709 18345 9743 18379
rect 9777 18345 9811 18379
rect 9845 18345 9879 18379
rect 9913 18345 9947 18379
rect 9981 18345 10015 18379
rect 10049 18345 10083 18379
rect 10117 18345 10151 18379
rect 10185 18345 10219 18379
rect 10253 18345 10287 18379
rect 10321 18345 10355 18379
rect 10389 18345 10423 18379
rect 10457 18345 10491 18379
rect 10525 18345 10559 18379
rect 10593 18345 10627 18379
rect 10661 18345 10695 18379
rect 10729 18345 10763 18379
rect 10797 18345 10831 18379
rect 10865 18345 10899 18379
rect 10933 18345 10967 18379
rect 11001 18345 11035 18379
rect 11069 18345 11103 18379
rect 11137 18345 11171 18379
rect 11205 18345 11239 18379
rect 11273 18345 11307 18379
rect 11341 18345 11375 18379
rect 11409 18345 11443 18379
rect 11477 18345 11511 18379
rect 11545 18345 11579 18379
rect 11613 18345 11647 18379
rect 11681 18345 11715 18379
rect 11749 18345 11783 18379
rect 11817 18345 11851 18379
rect 11885 18345 11919 18379
rect 11953 18345 11987 18379
rect 12021 18345 12055 18379
rect 12089 18345 12123 18379
rect 12157 18345 12191 18379
rect 12225 18345 12259 18379
rect 12293 18345 12327 18379
rect 12361 18345 12395 18379
rect 12429 18345 12463 18379
rect 12497 18345 12531 18379
rect 12565 18345 12599 18379
rect 12633 18345 12667 18379
rect 12701 18345 12735 18379
rect 12769 18345 12803 18379
rect 12837 18345 12871 18379
rect 12905 18345 12939 18379
rect 12973 18345 13007 18379
rect 13041 18345 13075 18379
rect 13109 18345 13143 18379
rect 13177 18345 13211 18379
rect 13245 18345 13279 18379
rect 13313 18345 13347 18379
rect 13381 18345 13415 18379
rect 13449 18345 13483 18379
rect 13517 18345 13551 18379
rect 13585 18345 13619 18379
rect 13653 18345 13687 18379
rect 13721 18345 13755 18379
rect 13789 18345 13823 18379
rect 13857 18345 13891 18379
rect 13925 18345 13959 18379
rect 13993 18345 14027 18379
rect 14061 18345 14095 18379
rect 14129 18345 14163 18379
rect 14197 18345 14231 18379
rect 14265 18345 14299 18379
rect 14333 18345 14367 18379
rect 14401 18345 14435 18379
rect 14469 18345 14503 18379
rect 14537 18345 14571 18379
rect 14605 18345 14639 18379
rect 14673 18345 14707 18379
rect 14741 18345 14772 18379
rect 197 18309 14772 18345
rect 197 18275 221 18309
rect 255 18275 290 18309
rect 324 18275 359 18309
rect 393 18275 427 18309
rect 461 18275 495 18309
rect 529 18275 563 18309
rect 597 18275 631 18309
rect 665 18275 699 18309
rect 733 18275 767 18309
rect 801 18275 835 18309
rect 869 18275 903 18309
rect 937 18275 971 18309
rect 1005 18275 1039 18309
rect 1073 18275 1107 18309
rect 1141 18275 1175 18309
rect 1209 18275 1243 18309
rect 1277 18275 1311 18309
rect 1345 18275 1379 18309
rect 1413 18275 1447 18309
rect 1481 18275 1515 18309
rect 1549 18275 1583 18309
rect 1617 18275 1651 18309
rect 1685 18275 1719 18309
rect 1753 18275 1787 18309
rect 1821 18275 1855 18309
rect 1889 18275 1923 18309
rect 1957 18275 1991 18309
rect 2025 18275 2059 18309
rect 2093 18275 2127 18309
rect 2161 18275 2195 18309
rect 2229 18275 2263 18309
rect 2297 18275 2331 18309
rect 2365 18275 2399 18309
rect 2433 18275 2467 18309
rect 2501 18275 2535 18309
rect 2569 18275 2603 18309
rect 2637 18275 2671 18309
rect 2705 18275 2739 18309
rect 2773 18275 2807 18309
rect 2841 18275 2875 18309
rect 2909 18275 2943 18309
rect 2977 18275 3011 18309
rect 3045 18275 3079 18309
rect 3113 18275 3147 18309
rect 3181 18275 3215 18309
rect 3249 18275 3283 18309
rect 3317 18275 3351 18309
rect 3385 18275 3419 18309
rect 3453 18275 3487 18309
rect 3521 18275 3555 18309
rect 3589 18275 3623 18309
rect 3657 18275 3691 18309
rect 3725 18275 3759 18309
rect 3793 18275 3827 18309
rect 3861 18275 3895 18309
rect 3929 18275 3963 18309
rect 3997 18275 4031 18309
rect 4065 18275 4099 18309
rect 4133 18275 4167 18309
rect 4201 18275 4235 18309
rect 4269 18275 4303 18309
rect 4337 18275 4371 18309
rect 4405 18275 4439 18309
rect 4473 18275 4507 18309
rect 4541 18275 4575 18309
rect 4609 18275 4643 18309
rect 4677 18275 4711 18309
rect 4745 18275 4779 18309
rect 4813 18275 4847 18309
rect 4881 18275 4915 18309
rect 4949 18275 4983 18309
rect 5017 18275 5051 18309
rect 5085 18275 5119 18309
rect 5153 18275 5187 18309
rect 5221 18275 5255 18309
rect 5289 18275 5323 18309
rect 5357 18275 5391 18309
rect 5425 18275 5459 18309
rect 5493 18275 5527 18309
rect 5561 18275 5595 18309
rect 5629 18275 5663 18309
rect 5697 18275 5731 18309
rect 5765 18275 5799 18309
rect 5833 18275 5867 18309
rect 5901 18275 5935 18309
rect 5969 18275 6003 18309
rect 6037 18275 6071 18309
rect 6105 18275 6139 18309
rect 6173 18275 6207 18309
rect 6241 18275 6275 18309
rect 6309 18275 6343 18309
rect 6377 18275 6411 18309
rect 6445 18275 6479 18309
rect 6513 18275 6547 18309
rect 6581 18275 6615 18309
rect 6649 18275 6683 18309
rect 6717 18275 6751 18309
rect 6785 18275 6819 18309
rect 6853 18275 6887 18309
rect 6921 18275 6955 18309
rect 6989 18275 7023 18309
rect 7057 18275 7091 18309
rect 7125 18275 7159 18309
rect 7193 18275 7227 18309
rect 7261 18275 7295 18309
rect 7329 18275 7363 18309
rect 7397 18275 7431 18309
rect 7465 18275 7499 18309
rect 7533 18275 7567 18309
rect 7601 18275 7635 18309
rect 7669 18275 7703 18309
rect 7737 18275 7771 18309
rect 7805 18275 7839 18309
rect 7873 18275 7907 18309
rect 7941 18275 7975 18309
rect 8009 18275 8043 18309
rect 8077 18275 8111 18309
rect 8145 18275 8179 18309
rect 8213 18275 8247 18309
rect 8281 18275 8315 18309
rect 8349 18275 8383 18309
rect 8417 18275 8451 18309
rect 8485 18275 8519 18309
rect 8553 18275 8587 18309
rect 8621 18275 8655 18309
rect 8689 18275 8723 18309
rect 8757 18275 8791 18309
rect 8825 18275 8859 18309
rect 8893 18275 8927 18309
rect 8961 18275 8995 18309
rect 9029 18275 9063 18309
rect 9097 18275 9131 18309
rect 9165 18275 9199 18309
rect 9233 18275 9267 18309
rect 9301 18275 9335 18309
rect 9369 18275 9403 18309
rect 9437 18275 9471 18309
rect 9505 18275 9539 18309
rect 9573 18275 9607 18309
rect 9641 18275 9675 18309
rect 9709 18275 9743 18309
rect 9777 18275 9811 18309
rect 9845 18275 9879 18309
rect 9913 18275 9947 18309
rect 9981 18275 10015 18309
rect 10049 18275 10083 18309
rect 10117 18275 10151 18309
rect 10185 18275 10219 18309
rect 10253 18275 10287 18309
rect 10321 18275 10355 18309
rect 10389 18275 10423 18309
rect 10457 18275 10491 18309
rect 10525 18275 10559 18309
rect 10593 18275 10627 18309
rect 10661 18275 10695 18309
rect 10729 18275 10763 18309
rect 10797 18275 10831 18309
rect 10865 18275 10899 18309
rect 10933 18275 10967 18309
rect 11001 18275 11035 18309
rect 11069 18275 11103 18309
rect 11137 18275 11171 18309
rect 11205 18275 11239 18309
rect 11273 18275 11307 18309
rect 11341 18275 11375 18309
rect 11409 18275 11443 18309
rect 11477 18275 11511 18309
rect 11545 18275 11579 18309
rect 11613 18275 11647 18309
rect 11681 18275 11715 18309
rect 11749 18275 11783 18309
rect 11817 18275 11851 18309
rect 11885 18275 11919 18309
rect 11953 18275 11987 18309
rect 12021 18275 12055 18309
rect 12089 18275 12123 18309
rect 12157 18275 12191 18309
rect 12225 18275 12259 18309
rect 12293 18275 12327 18309
rect 12361 18275 12395 18309
rect 12429 18275 12463 18309
rect 12497 18275 12531 18309
rect 12565 18275 12599 18309
rect 12633 18275 12667 18309
rect 12701 18275 12735 18309
rect 12769 18275 12803 18309
rect 12837 18275 12871 18309
rect 12905 18275 12939 18309
rect 12973 18275 13007 18309
rect 13041 18275 13075 18309
rect 13109 18275 13143 18309
rect 13177 18275 13211 18309
rect 13245 18275 13279 18309
rect 13313 18275 13347 18309
rect 13381 18275 13415 18309
rect 13449 18275 13483 18309
rect 13517 18275 13551 18309
rect 13585 18275 13619 18309
rect 13653 18275 13687 18309
rect 13721 18275 13755 18309
rect 13789 18275 13823 18309
rect 13857 18275 13891 18309
rect 13925 18275 13959 18309
rect 13993 18275 14027 18309
rect 14061 18275 14095 18309
rect 14129 18275 14163 18309
rect 14197 18275 14231 18309
rect 14265 18275 14299 18309
rect 14333 18275 14367 18309
rect 14401 18275 14435 18309
rect 14469 18275 14503 18309
rect 14537 18275 14571 18309
rect 14605 18275 14639 18309
rect 14673 18275 14707 18309
rect 14741 18275 14772 18309
rect 197 18239 14772 18275
rect 197 18205 221 18239
rect 255 18205 290 18239
rect 324 18205 359 18239
rect 393 18205 427 18239
rect 461 18205 495 18239
rect 529 18205 563 18239
rect 597 18205 631 18239
rect 665 18205 699 18239
rect 733 18205 767 18239
rect 801 18205 835 18239
rect 869 18205 903 18239
rect 937 18205 971 18239
rect 1005 18205 1039 18239
rect 1073 18205 1107 18239
rect 1141 18205 1175 18239
rect 1209 18205 1243 18239
rect 1277 18205 1311 18239
rect 1345 18205 1379 18239
rect 1413 18205 1447 18239
rect 1481 18205 1515 18239
rect 1549 18205 1583 18239
rect 1617 18205 1651 18239
rect 1685 18205 1719 18239
rect 1753 18205 1787 18239
rect 1821 18205 1855 18239
rect 1889 18205 1923 18239
rect 1957 18205 1991 18239
rect 2025 18205 2059 18239
rect 2093 18205 2127 18239
rect 2161 18205 2195 18239
rect 2229 18205 2263 18239
rect 2297 18205 2331 18239
rect 2365 18205 2399 18239
rect 2433 18205 2467 18239
rect 2501 18205 2535 18239
rect 2569 18205 2603 18239
rect 2637 18205 2671 18239
rect 2705 18205 2739 18239
rect 2773 18205 2807 18239
rect 2841 18205 2875 18239
rect 2909 18205 2943 18239
rect 2977 18205 3011 18239
rect 3045 18205 3079 18239
rect 3113 18205 3147 18239
rect 3181 18205 3215 18239
rect 3249 18205 3283 18239
rect 3317 18205 3351 18239
rect 3385 18205 3419 18239
rect 3453 18205 3487 18239
rect 3521 18205 3555 18239
rect 3589 18205 3623 18239
rect 3657 18205 3691 18239
rect 3725 18205 3759 18239
rect 3793 18205 3827 18239
rect 3861 18205 3895 18239
rect 3929 18205 3963 18239
rect 3997 18205 4031 18239
rect 4065 18205 4099 18239
rect 4133 18205 4167 18239
rect 4201 18205 4235 18239
rect 4269 18205 4303 18239
rect 4337 18205 4371 18239
rect 4405 18205 4439 18239
rect 4473 18205 4507 18239
rect 4541 18205 4575 18239
rect 4609 18205 4643 18239
rect 4677 18205 4711 18239
rect 4745 18205 4779 18239
rect 4813 18205 4847 18239
rect 4881 18205 4915 18239
rect 4949 18205 4983 18239
rect 5017 18205 5051 18239
rect 5085 18205 5119 18239
rect 5153 18205 5187 18239
rect 5221 18205 5255 18239
rect 5289 18205 5323 18239
rect 5357 18205 5391 18239
rect 5425 18205 5459 18239
rect 5493 18205 5527 18239
rect 5561 18205 5595 18239
rect 5629 18205 5663 18239
rect 5697 18205 5731 18239
rect 5765 18205 5799 18239
rect 5833 18205 5867 18239
rect 5901 18205 5935 18239
rect 5969 18205 6003 18239
rect 6037 18205 6071 18239
rect 6105 18205 6139 18239
rect 6173 18205 6207 18239
rect 6241 18205 6275 18239
rect 6309 18205 6343 18239
rect 6377 18205 6411 18239
rect 6445 18205 6479 18239
rect 6513 18205 6547 18239
rect 6581 18205 6615 18239
rect 6649 18205 6683 18239
rect 6717 18205 6751 18239
rect 6785 18205 6819 18239
rect 6853 18205 6887 18239
rect 6921 18205 6955 18239
rect 6989 18205 7023 18239
rect 7057 18205 7091 18239
rect 7125 18205 7159 18239
rect 7193 18205 7227 18239
rect 7261 18205 7295 18239
rect 7329 18205 7363 18239
rect 7397 18205 7431 18239
rect 7465 18205 7499 18239
rect 7533 18205 7567 18239
rect 7601 18205 7635 18239
rect 7669 18205 7703 18239
rect 7737 18205 7771 18239
rect 7805 18205 7839 18239
rect 7873 18205 7907 18239
rect 7941 18205 7975 18239
rect 8009 18205 8043 18239
rect 8077 18205 8111 18239
rect 8145 18205 8179 18239
rect 8213 18205 8247 18239
rect 8281 18205 8315 18239
rect 8349 18205 8383 18239
rect 8417 18205 8451 18239
rect 8485 18205 8519 18239
rect 8553 18205 8587 18239
rect 8621 18205 8655 18239
rect 8689 18205 8723 18239
rect 8757 18205 8791 18239
rect 8825 18205 8859 18239
rect 8893 18205 8927 18239
rect 8961 18205 8995 18239
rect 9029 18205 9063 18239
rect 9097 18205 9131 18239
rect 9165 18205 9199 18239
rect 9233 18205 9267 18239
rect 9301 18205 9335 18239
rect 9369 18205 9403 18239
rect 9437 18205 9471 18239
rect 9505 18205 9539 18239
rect 9573 18205 9607 18239
rect 9641 18205 9675 18239
rect 9709 18205 9743 18239
rect 9777 18205 9811 18239
rect 9845 18205 9879 18239
rect 9913 18205 9947 18239
rect 9981 18205 10015 18239
rect 10049 18205 10083 18239
rect 10117 18205 10151 18239
rect 10185 18205 10219 18239
rect 10253 18205 10287 18239
rect 10321 18205 10355 18239
rect 10389 18205 10423 18239
rect 10457 18205 10491 18239
rect 10525 18205 10559 18239
rect 10593 18205 10627 18239
rect 10661 18205 10695 18239
rect 10729 18205 10763 18239
rect 10797 18205 10831 18239
rect 10865 18205 10899 18239
rect 10933 18205 10967 18239
rect 11001 18205 11035 18239
rect 11069 18205 11103 18239
rect 11137 18205 11171 18239
rect 11205 18205 11239 18239
rect 11273 18205 11307 18239
rect 11341 18205 11375 18239
rect 11409 18205 11443 18239
rect 11477 18205 11511 18239
rect 11545 18205 11579 18239
rect 11613 18205 11647 18239
rect 11681 18205 11715 18239
rect 11749 18205 11783 18239
rect 11817 18205 11851 18239
rect 11885 18205 11919 18239
rect 11953 18205 11987 18239
rect 12021 18205 12055 18239
rect 12089 18205 12123 18239
rect 12157 18205 12191 18239
rect 12225 18205 12259 18239
rect 12293 18205 12327 18239
rect 12361 18205 12395 18239
rect 12429 18205 12463 18239
rect 12497 18205 12531 18239
rect 12565 18205 12599 18239
rect 12633 18205 12667 18239
rect 12701 18205 12735 18239
rect 12769 18205 12803 18239
rect 12837 18205 12871 18239
rect 12905 18205 12939 18239
rect 12973 18205 13007 18239
rect 13041 18205 13075 18239
rect 13109 18205 13143 18239
rect 13177 18205 13211 18239
rect 13245 18205 13279 18239
rect 13313 18205 13347 18239
rect 13381 18205 13415 18239
rect 13449 18205 13483 18239
rect 13517 18205 13551 18239
rect 13585 18205 13619 18239
rect 13653 18205 13687 18239
rect 13721 18205 13755 18239
rect 13789 18205 13823 18239
rect 13857 18205 13891 18239
rect 13925 18205 13959 18239
rect 13993 18205 14027 18239
rect 14061 18205 14095 18239
rect 14129 18205 14163 18239
rect 14197 18205 14231 18239
rect 14265 18205 14299 18239
rect 14333 18205 14367 18239
rect 14401 18205 14435 18239
rect 14469 18205 14503 18239
rect 14537 18205 14571 18239
rect 14605 18205 14639 18239
rect 14673 18205 14707 18239
rect 14741 18205 14772 18239
rect 197 18169 14772 18205
rect 197 18135 221 18169
rect 255 18135 290 18169
rect 324 18135 359 18169
rect 393 18135 427 18169
rect 461 18135 495 18169
rect 529 18135 563 18169
rect 597 18135 631 18169
rect 665 18135 699 18169
rect 733 18135 767 18169
rect 801 18135 835 18169
rect 869 18135 903 18169
rect 937 18135 971 18169
rect 1005 18135 1039 18169
rect 1073 18135 1107 18169
rect 1141 18135 1175 18169
rect 1209 18135 1243 18169
rect 1277 18135 1311 18169
rect 1345 18135 1379 18169
rect 1413 18135 1447 18169
rect 1481 18135 1515 18169
rect 1549 18135 1583 18169
rect 1617 18135 1651 18169
rect 1685 18135 1719 18169
rect 1753 18135 1787 18169
rect 1821 18135 1855 18169
rect 1889 18135 1923 18169
rect 1957 18135 1991 18169
rect 2025 18135 2059 18169
rect 2093 18135 2127 18169
rect 2161 18135 2195 18169
rect 2229 18135 2263 18169
rect 2297 18135 2331 18169
rect 2365 18135 2399 18169
rect 2433 18135 2467 18169
rect 2501 18135 2535 18169
rect 2569 18135 2603 18169
rect 2637 18135 2671 18169
rect 2705 18135 2739 18169
rect 2773 18135 2807 18169
rect 2841 18135 2875 18169
rect 2909 18135 2943 18169
rect 2977 18135 3011 18169
rect 3045 18135 3079 18169
rect 3113 18135 3147 18169
rect 3181 18135 3215 18169
rect 3249 18135 3283 18169
rect 3317 18135 3351 18169
rect 3385 18135 3419 18169
rect 3453 18135 3487 18169
rect 3521 18135 3555 18169
rect 3589 18135 3623 18169
rect 3657 18135 3691 18169
rect 3725 18135 3759 18169
rect 3793 18135 3827 18169
rect 3861 18135 3895 18169
rect 3929 18135 3963 18169
rect 3997 18135 4031 18169
rect 4065 18135 4099 18169
rect 4133 18135 4167 18169
rect 4201 18135 4235 18169
rect 4269 18135 4303 18169
rect 4337 18135 4371 18169
rect 4405 18135 4439 18169
rect 4473 18135 4507 18169
rect 4541 18135 4575 18169
rect 4609 18135 4643 18169
rect 4677 18135 4711 18169
rect 4745 18135 4779 18169
rect 4813 18135 4847 18169
rect 4881 18135 4915 18169
rect 4949 18135 4983 18169
rect 5017 18135 5051 18169
rect 5085 18135 5119 18169
rect 5153 18135 5187 18169
rect 5221 18135 5255 18169
rect 5289 18135 5323 18169
rect 5357 18135 5391 18169
rect 5425 18135 5459 18169
rect 5493 18135 5527 18169
rect 5561 18135 5595 18169
rect 5629 18135 5663 18169
rect 5697 18135 5731 18169
rect 5765 18135 5799 18169
rect 5833 18135 5867 18169
rect 5901 18135 5935 18169
rect 5969 18135 6003 18169
rect 6037 18135 6071 18169
rect 6105 18135 6139 18169
rect 6173 18135 6207 18169
rect 6241 18135 6275 18169
rect 6309 18135 6343 18169
rect 6377 18135 6411 18169
rect 6445 18135 6479 18169
rect 6513 18135 6547 18169
rect 6581 18135 6615 18169
rect 6649 18135 6683 18169
rect 6717 18135 6751 18169
rect 6785 18135 6819 18169
rect 6853 18135 6887 18169
rect 6921 18135 6955 18169
rect 6989 18135 7023 18169
rect 7057 18135 7091 18169
rect 7125 18135 7159 18169
rect 7193 18135 7227 18169
rect 7261 18135 7295 18169
rect 7329 18135 7363 18169
rect 7397 18135 7431 18169
rect 7465 18135 7499 18169
rect 7533 18135 7567 18169
rect 7601 18135 7635 18169
rect 7669 18135 7703 18169
rect 7737 18135 7771 18169
rect 7805 18135 7839 18169
rect 7873 18135 7907 18169
rect 7941 18135 7975 18169
rect 8009 18135 8043 18169
rect 8077 18135 8111 18169
rect 8145 18135 8179 18169
rect 8213 18135 8247 18169
rect 8281 18135 8315 18169
rect 8349 18135 8383 18169
rect 8417 18135 8451 18169
rect 8485 18135 8519 18169
rect 8553 18135 8587 18169
rect 8621 18135 8655 18169
rect 8689 18135 8723 18169
rect 8757 18135 8791 18169
rect 8825 18135 8859 18169
rect 8893 18135 8927 18169
rect 8961 18135 8995 18169
rect 9029 18135 9063 18169
rect 9097 18135 9131 18169
rect 9165 18135 9199 18169
rect 9233 18135 9267 18169
rect 9301 18135 9335 18169
rect 9369 18135 9403 18169
rect 9437 18135 9471 18169
rect 9505 18135 9539 18169
rect 9573 18135 9607 18169
rect 9641 18135 9675 18169
rect 9709 18135 9743 18169
rect 9777 18135 9811 18169
rect 9845 18135 9879 18169
rect 9913 18135 9947 18169
rect 9981 18135 10015 18169
rect 10049 18135 10083 18169
rect 10117 18135 10151 18169
rect 10185 18135 10219 18169
rect 10253 18135 10287 18169
rect 10321 18135 10355 18169
rect 10389 18135 10423 18169
rect 10457 18135 10491 18169
rect 10525 18135 10559 18169
rect 10593 18135 10627 18169
rect 10661 18135 10695 18169
rect 10729 18135 10763 18169
rect 10797 18135 10831 18169
rect 10865 18135 10899 18169
rect 10933 18135 10967 18169
rect 11001 18135 11035 18169
rect 11069 18135 11103 18169
rect 11137 18135 11171 18169
rect 11205 18135 11239 18169
rect 11273 18135 11307 18169
rect 11341 18135 11375 18169
rect 11409 18135 11443 18169
rect 11477 18135 11511 18169
rect 11545 18135 11579 18169
rect 11613 18135 11647 18169
rect 11681 18135 11715 18169
rect 11749 18135 11783 18169
rect 11817 18135 11851 18169
rect 11885 18135 11919 18169
rect 11953 18135 11987 18169
rect 12021 18135 12055 18169
rect 12089 18135 12123 18169
rect 12157 18135 12191 18169
rect 12225 18135 12259 18169
rect 12293 18135 12327 18169
rect 12361 18135 12395 18169
rect 12429 18135 12463 18169
rect 12497 18135 12531 18169
rect 12565 18135 12599 18169
rect 12633 18135 12667 18169
rect 12701 18135 12735 18169
rect 12769 18135 12803 18169
rect 12837 18135 12871 18169
rect 12905 18135 12939 18169
rect 12973 18135 13007 18169
rect 13041 18135 13075 18169
rect 13109 18135 13143 18169
rect 13177 18135 13211 18169
rect 13245 18135 13279 18169
rect 13313 18135 13347 18169
rect 13381 18135 13415 18169
rect 13449 18135 13483 18169
rect 13517 18135 13551 18169
rect 13585 18135 13619 18169
rect 13653 18135 13687 18169
rect 13721 18135 13755 18169
rect 13789 18135 13823 18169
rect 13857 18135 13891 18169
rect 13925 18135 13959 18169
rect 13993 18135 14027 18169
rect 14061 18135 14095 18169
rect 14129 18135 14163 18169
rect 14197 18135 14231 18169
rect 14265 18135 14299 18169
rect 14333 18135 14367 18169
rect 14401 18135 14435 18169
rect 14469 18135 14503 18169
rect 14537 18135 14571 18169
rect 14605 18135 14639 18169
rect 14673 18135 14707 18169
rect 14741 18135 14772 18169
rect 197 18099 14772 18135
rect 197 18065 221 18099
rect 255 18065 290 18099
rect 324 18065 359 18099
rect 393 18065 427 18099
rect 461 18065 495 18099
rect 529 18065 563 18099
rect 597 18065 631 18099
rect 665 18065 699 18099
rect 733 18065 767 18099
rect 801 18065 835 18099
rect 869 18065 903 18099
rect 937 18065 971 18099
rect 1005 18065 1039 18099
rect 1073 18065 1107 18099
rect 1141 18065 1175 18099
rect 1209 18065 1243 18099
rect 1277 18065 1311 18099
rect 1345 18065 1379 18099
rect 1413 18065 1447 18099
rect 1481 18065 1515 18099
rect 1549 18065 1583 18099
rect 1617 18065 1651 18099
rect 1685 18065 1719 18099
rect 1753 18065 1787 18099
rect 1821 18065 1855 18099
rect 1889 18065 1923 18099
rect 1957 18065 1991 18099
rect 2025 18065 2059 18099
rect 2093 18065 2127 18099
rect 2161 18065 2195 18099
rect 2229 18065 2263 18099
rect 2297 18065 2331 18099
rect 2365 18065 2399 18099
rect 2433 18065 2467 18099
rect 2501 18065 2535 18099
rect 2569 18065 2603 18099
rect 2637 18065 2671 18099
rect 2705 18065 2739 18099
rect 2773 18065 2807 18099
rect 2841 18065 2875 18099
rect 2909 18065 2943 18099
rect 2977 18065 3011 18099
rect 3045 18065 3079 18099
rect 3113 18065 3147 18099
rect 3181 18065 3215 18099
rect 3249 18065 3283 18099
rect 3317 18065 3351 18099
rect 3385 18065 3419 18099
rect 3453 18065 3487 18099
rect 3521 18065 3555 18099
rect 3589 18065 3623 18099
rect 3657 18065 3691 18099
rect 3725 18065 3759 18099
rect 3793 18065 3827 18099
rect 3861 18065 3895 18099
rect 3929 18065 3963 18099
rect 3997 18065 4031 18099
rect 4065 18065 4099 18099
rect 4133 18065 4167 18099
rect 4201 18065 4235 18099
rect 4269 18065 4303 18099
rect 4337 18065 4371 18099
rect 4405 18065 4439 18099
rect 4473 18065 4507 18099
rect 4541 18065 4575 18099
rect 4609 18065 4643 18099
rect 4677 18065 4711 18099
rect 4745 18065 4779 18099
rect 4813 18065 4847 18099
rect 4881 18065 4915 18099
rect 4949 18065 4983 18099
rect 5017 18065 5051 18099
rect 5085 18065 5119 18099
rect 5153 18065 5187 18099
rect 5221 18065 5255 18099
rect 5289 18065 5323 18099
rect 5357 18065 5391 18099
rect 5425 18065 5459 18099
rect 5493 18065 5527 18099
rect 5561 18065 5595 18099
rect 5629 18065 5663 18099
rect 5697 18065 5731 18099
rect 5765 18065 5799 18099
rect 5833 18065 5867 18099
rect 5901 18065 5935 18099
rect 5969 18065 6003 18099
rect 6037 18065 6071 18099
rect 6105 18065 6139 18099
rect 6173 18065 6207 18099
rect 6241 18065 6275 18099
rect 6309 18065 6343 18099
rect 6377 18065 6411 18099
rect 6445 18065 6479 18099
rect 6513 18065 6547 18099
rect 6581 18065 6615 18099
rect 6649 18065 6683 18099
rect 6717 18065 6751 18099
rect 6785 18065 6819 18099
rect 6853 18065 6887 18099
rect 6921 18065 6955 18099
rect 6989 18065 7023 18099
rect 7057 18065 7091 18099
rect 7125 18065 7159 18099
rect 7193 18065 7227 18099
rect 7261 18065 7295 18099
rect 7329 18065 7363 18099
rect 7397 18065 7431 18099
rect 7465 18065 7499 18099
rect 7533 18065 7567 18099
rect 7601 18065 7635 18099
rect 7669 18065 7703 18099
rect 7737 18065 7771 18099
rect 7805 18065 7839 18099
rect 7873 18065 7907 18099
rect 7941 18065 7975 18099
rect 8009 18065 8043 18099
rect 8077 18065 8111 18099
rect 8145 18065 8179 18099
rect 8213 18065 8247 18099
rect 8281 18065 8315 18099
rect 8349 18065 8383 18099
rect 8417 18065 8451 18099
rect 8485 18065 8519 18099
rect 8553 18065 8587 18099
rect 8621 18065 8655 18099
rect 8689 18065 8723 18099
rect 8757 18065 8791 18099
rect 8825 18065 8859 18099
rect 8893 18065 8927 18099
rect 8961 18065 8995 18099
rect 9029 18065 9063 18099
rect 9097 18065 9131 18099
rect 9165 18065 9199 18099
rect 9233 18065 9267 18099
rect 9301 18065 9335 18099
rect 9369 18065 9403 18099
rect 9437 18065 9471 18099
rect 9505 18065 9539 18099
rect 9573 18065 9607 18099
rect 9641 18065 9675 18099
rect 9709 18065 9743 18099
rect 9777 18065 9811 18099
rect 9845 18065 9879 18099
rect 9913 18065 9947 18099
rect 9981 18065 10015 18099
rect 10049 18065 10083 18099
rect 10117 18065 10151 18099
rect 10185 18065 10219 18099
rect 10253 18065 10287 18099
rect 10321 18065 10355 18099
rect 10389 18065 10423 18099
rect 10457 18065 10491 18099
rect 10525 18065 10559 18099
rect 10593 18065 10627 18099
rect 10661 18065 10695 18099
rect 10729 18065 10763 18099
rect 10797 18065 10831 18099
rect 10865 18065 10899 18099
rect 10933 18065 10967 18099
rect 11001 18065 11035 18099
rect 11069 18065 11103 18099
rect 11137 18065 11171 18099
rect 11205 18065 11239 18099
rect 11273 18065 11307 18099
rect 11341 18065 11375 18099
rect 11409 18065 11443 18099
rect 11477 18065 11511 18099
rect 11545 18065 11579 18099
rect 11613 18065 11647 18099
rect 11681 18065 11715 18099
rect 11749 18065 11783 18099
rect 11817 18065 11851 18099
rect 11885 18065 11919 18099
rect 11953 18065 11987 18099
rect 12021 18065 12055 18099
rect 12089 18065 12123 18099
rect 12157 18065 12191 18099
rect 12225 18065 12259 18099
rect 12293 18065 12327 18099
rect 12361 18065 12395 18099
rect 12429 18065 12463 18099
rect 12497 18065 12531 18099
rect 12565 18065 12599 18099
rect 12633 18065 12667 18099
rect 12701 18065 12735 18099
rect 12769 18065 12803 18099
rect 12837 18065 12871 18099
rect 12905 18065 12939 18099
rect 12973 18065 13007 18099
rect 13041 18065 13075 18099
rect 13109 18065 13143 18099
rect 13177 18065 13211 18099
rect 13245 18065 13279 18099
rect 13313 18065 13347 18099
rect 13381 18065 13415 18099
rect 13449 18065 13483 18099
rect 13517 18065 13551 18099
rect 13585 18065 13619 18099
rect 13653 18065 13687 18099
rect 13721 18065 13755 18099
rect 13789 18065 13823 18099
rect 13857 18065 13891 18099
rect 13925 18065 13959 18099
rect 13993 18065 14027 18099
rect 14061 18065 14095 18099
rect 14129 18065 14163 18099
rect 14197 18065 14231 18099
rect 14265 18065 14299 18099
rect 14333 18065 14367 18099
rect 14401 18065 14435 18099
rect 14469 18065 14503 18099
rect 14537 18065 14571 18099
rect 14605 18065 14639 18099
rect 14673 18065 14707 18099
rect 14741 18065 14772 18099
rect 197 18029 14772 18065
rect 197 17995 221 18029
rect 255 17995 290 18029
rect 324 17995 359 18029
rect 393 17995 427 18029
rect 461 17995 495 18029
rect 529 17995 563 18029
rect 597 17995 631 18029
rect 665 17995 699 18029
rect 733 17995 767 18029
rect 801 17995 835 18029
rect 869 17995 903 18029
rect 937 17995 971 18029
rect 1005 17995 1039 18029
rect 1073 17995 1107 18029
rect 1141 17995 1175 18029
rect 1209 17995 1243 18029
rect 1277 17995 1311 18029
rect 1345 17995 1379 18029
rect 1413 17995 1447 18029
rect 1481 17995 1515 18029
rect 1549 17995 1583 18029
rect 1617 17995 1651 18029
rect 1685 17995 1719 18029
rect 1753 17995 1787 18029
rect 1821 17995 1855 18029
rect 1889 17995 1923 18029
rect 1957 17995 1991 18029
rect 2025 17995 2059 18029
rect 2093 17995 2127 18029
rect 2161 17995 2195 18029
rect 2229 17995 2263 18029
rect 2297 17995 2331 18029
rect 2365 17995 2399 18029
rect 2433 17995 2467 18029
rect 2501 17995 2535 18029
rect 2569 17995 2603 18029
rect 2637 17995 2671 18029
rect 2705 17995 2739 18029
rect 2773 17995 2807 18029
rect 2841 17995 2875 18029
rect 2909 17995 2943 18029
rect 2977 17995 3011 18029
rect 3045 17995 3079 18029
rect 3113 17995 3147 18029
rect 3181 17995 3215 18029
rect 3249 17995 3283 18029
rect 3317 17995 3351 18029
rect 3385 17995 3419 18029
rect 3453 17995 3487 18029
rect 3521 17995 3555 18029
rect 3589 17995 3623 18029
rect 3657 17995 3691 18029
rect 3725 17995 3759 18029
rect 3793 17995 3827 18029
rect 3861 17995 3895 18029
rect 3929 17995 3963 18029
rect 3997 17995 4031 18029
rect 4065 17995 4099 18029
rect 4133 17995 4167 18029
rect 4201 17995 4235 18029
rect 4269 17995 4303 18029
rect 4337 17995 4371 18029
rect 4405 17995 4439 18029
rect 4473 17995 4507 18029
rect 4541 17995 4575 18029
rect 4609 17995 4643 18029
rect 4677 17995 4711 18029
rect 4745 17995 4779 18029
rect 4813 17995 4847 18029
rect 4881 17995 4915 18029
rect 4949 17995 4983 18029
rect 5017 17995 5051 18029
rect 5085 17995 5119 18029
rect 5153 17995 5187 18029
rect 5221 17995 5255 18029
rect 5289 17995 5323 18029
rect 5357 17995 5391 18029
rect 5425 17995 5459 18029
rect 5493 17995 5527 18029
rect 5561 17995 5595 18029
rect 5629 17995 5663 18029
rect 5697 17995 5731 18029
rect 5765 17995 5799 18029
rect 5833 17995 5867 18029
rect 5901 17995 5935 18029
rect 5969 17995 6003 18029
rect 6037 17995 6071 18029
rect 6105 17995 6139 18029
rect 6173 17995 6207 18029
rect 6241 17995 6275 18029
rect 6309 17995 6343 18029
rect 6377 17995 6411 18029
rect 6445 17995 6479 18029
rect 6513 17995 6547 18029
rect 6581 17995 6615 18029
rect 6649 17995 6683 18029
rect 6717 17995 6751 18029
rect 6785 17995 6819 18029
rect 6853 17995 6887 18029
rect 6921 17995 6955 18029
rect 6989 17995 7023 18029
rect 7057 17995 7091 18029
rect 7125 17995 7159 18029
rect 7193 17995 7227 18029
rect 7261 17995 7295 18029
rect 7329 17995 7363 18029
rect 7397 17995 7431 18029
rect 7465 17995 7499 18029
rect 7533 17995 7567 18029
rect 7601 17995 7635 18029
rect 7669 17995 7703 18029
rect 7737 17995 7771 18029
rect 7805 17995 7839 18029
rect 7873 17995 7907 18029
rect 7941 17995 7975 18029
rect 8009 17995 8043 18029
rect 8077 17995 8111 18029
rect 8145 17995 8179 18029
rect 8213 17995 8247 18029
rect 8281 17995 8315 18029
rect 8349 17995 8383 18029
rect 8417 17995 8451 18029
rect 8485 17995 8519 18029
rect 8553 17995 8587 18029
rect 8621 17995 8655 18029
rect 8689 17995 8723 18029
rect 8757 17995 8791 18029
rect 8825 17995 8859 18029
rect 8893 17995 8927 18029
rect 8961 17995 8995 18029
rect 9029 17995 9063 18029
rect 9097 17995 9131 18029
rect 9165 17995 9199 18029
rect 9233 17995 9267 18029
rect 9301 17995 9335 18029
rect 9369 17995 9403 18029
rect 9437 17995 9471 18029
rect 9505 17995 9539 18029
rect 9573 17995 9607 18029
rect 9641 17995 9675 18029
rect 9709 17995 9743 18029
rect 9777 17995 9811 18029
rect 9845 17995 9879 18029
rect 9913 17995 9947 18029
rect 9981 17995 10015 18029
rect 10049 17995 10083 18029
rect 10117 17995 10151 18029
rect 10185 17995 10219 18029
rect 10253 17995 10287 18029
rect 10321 17995 10355 18029
rect 10389 17995 10423 18029
rect 10457 17995 10491 18029
rect 10525 17995 10559 18029
rect 10593 17995 10627 18029
rect 10661 17995 10695 18029
rect 10729 17995 10763 18029
rect 10797 17995 10831 18029
rect 10865 17995 10899 18029
rect 10933 17995 10967 18029
rect 11001 17995 11035 18029
rect 11069 17995 11103 18029
rect 11137 17995 11171 18029
rect 11205 17995 11239 18029
rect 11273 17995 11307 18029
rect 11341 17995 11375 18029
rect 11409 17995 11443 18029
rect 11477 17995 11511 18029
rect 11545 17995 11579 18029
rect 11613 17995 11647 18029
rect 11681 17995 11715 18029
rect 11749 17995 11783 18029
rect 11817 17995 11851 18029
rect 11885 17995 11919 18029
rect 11953 17995 11987 18029
rect 12021 17995 12055 18029
rect 12089 17995 12123 18029
rect 12157 17995 12191 18029
rect 12225 17995 12259 18029
rect 12293 17995 12327 18029
rect 12361 17995 12395 18029
rect 12429 17995 12463 18029
rect 12497 17995 12531 18029
rect 12565 17995 12599 18029
rect 12633 17995 12667 18029
rect 12701 17995 12735 18029
rect 12769 17995 12803 18029
rect 12837 17995 12871 18029
rect 12905 17995 12939 18029
rect 12973 17995 13007 18029
rect 13041 17995 13075 18029
rect 13109 17995 13143 18029
rect 13177 17995 13211 18029
rect 13245 17995 13279 18029
rect 13313 17995 13347 18029
rect 13381 17995 13415 18029
rect 13449 17995 13483 18029
rect 13517 17995 13551 18029
rect 13585 17995 13619 18029
rect 13653 17995 13687 18029
rect 13721 17995 13755 18029
rect 13789 17995 13823 18029
rect 13857 17995 13891 18029
rect 13925 17995 13959 18029
rect 13993 17995 14027 18029
rect 14061 17995 14095 18029
rect 14129 17995 14163 18029
rect 14197 17995 14231 18029
rect 14265 17995 14299 18029
rect 14333 17995 14367 18029
rect 14401 17995 14435 18029
rect 14469 17995 14503 18029
rect 14537 17995 14571 18029
rect 14605 17995 14639 18029
rect 14673 17995 14707 18029
rect 14741 17995 14772 18029
rect 197 17959 14772 17995
rect 197 17925 221 17959
rect 255 17925 290 17959
rect 324 17925 359 17959
rect 393 17925 427 17959
rect 461 17925 495 17959
rect 529 17925 563 17959
rect 597 17925 631 17959
rect 665 17925 699 17959
rect 733 17925 767 17959
rect 801 17925 835 17959
rect 869 17925 903 17959
rect 937 17925 971 17959
rect 1005 17925 1039 17959
rect 1073 17925 1107 17959
rect 1141 17925 1175 17959
rect 1209 17925 1243 17959
rect 1277 17925 1311 17959
rect 1345 17925 1379 17959
rect 1413 17925 1447 17959
rect 1481 17925 1515 17959
rect 1549 17925 1583 17959
rect 1617 17925 1651 17959
rect 1685 17925 1719 17959
rect 1753 17925 1787 17959
rect 1821 17925 1855 17959
rect 1889 17925 1923 17959
rect 1957 17925 1991 17959
rect 2025 17925 2059 17959
rect 2093 17925 2127 17959
rect 2161 17925 2195 17959
rect 2229 17925 2263 17959
rect 2297 17925 2331 17959
rect 2365 17925 2399 17959
rect 2433 17925 2467 17959
rect 2501 17925 2535 17959
rect 2569 17925 2603 17959
rect 2637 17925 2671 17959
rect 2705 17925 2739 17959
rect 2773 17925 2807 17959
rect 2841 17925 2875 17959
rect 2909 17925 2943 17959
rect 2977 17925 3011 17959
rect 3045 17925 3079 17959
rect 3113 17925 3147 17959
rect 3181 17925 3215 17959
rect 3249 17925 3283 17959
rect 3317 17925 3351 17959
rect 3385 17925 3419 17959
rect 3453 17925 3487 17959
rect 3521 17925 3555 17959
rect 3589 17925 3623 17959
rect 3657 17925 3691 17959
rect 3725 17925 3759 17959
rect 3793 17925 3827 17959
rect 3861 17925 3895 17959
rect 3929 17925 3963 17959
rect 3997 17925 4031 17959
rect 4065 17925 4099 17959
rect 4133 17925 4167 17959
rect 4201 17925 4235 17959
rect 4269 17925 4303 17959
rect 4337 17925 4371 17959
rect 4405 17925 4439 17959
rect 4473 17925 4507 17959
rect 4541 17925 4575 17959
rect 4609 17925 4643 17959
rect 4677 17925 4711 17959
rect 4745 17925 4779 17959
rect 4813 17925 4847 17959
rect 4881 17925 4915 17959
rect 4949 17925 4983 17959
rect 5017 17925 5051 17959
rect 5085 17925 5119 17959
rect 5153 17925 5187 17959
rect 5221 17925 5255 17959
rect 5289 17925 5323 17959
rect 5357 17925 5391 17959
rect 5425 17925 5459 17959
rect 5493 17925 5527 17959
rect 5561 17925 5595 17959
rect 5629 17925 5663 17959
rect 5697 17925 5731 17959
rect 5765 17925 5799 17959
rect 5833 17925 5867 17959
rect 5901 17925 5935 17959
rect 5969 17925 6003 17959
rect 6037 17925 6071 17959
rect 6105 17925 6139 17959
rect 6173 17925 6207 17959
rect 6241 17925 6275 17959
rect 6309 17925 6343 17959
rect 6377 17925 6411 17959
rect 6445 17925 6479 17959
rect 6513 17925 6547 17959
rect 6581 17925 6615 17959
rect 6649 17925 6683 17959
rect 6717 17925 6751 17959
rect 6785 17925 6819 17959
rect 6853 17925 6887 17959
rect 6921 17925 6955 17959
rect 6989 17925 7023 17959
rect 7057 17925 7091 17959
rect 7125 17925 7159 17959
rect 7193 17925 7227 17959
rect 7261 17925 7295 17959
rect 7329 17925 7363 17959
rect 7397 17925 7431 17959
rect 7465 17925 7499 17959
rect 7533 17925 7567 17959
rect 7601 17925 7635 17959
rect 7669 17925 7703 17959
rect 7737 17925 7771 17959
rect 7805 17925 7839 17959
rect 7873 17925 7907 17959
rect 7941 17925 7975 17959
rect 8009 17925 8043 17959
rect 8077 17925 8111 17959
rect 8145 17925 8179 17959
rect 8213 17925 8247 17959
rect 8281 17925 8315 17959
rect 8349 17925 8383 17959
rect 8417 17925 8451 17959
rect 8485 17925 8519 17959
rect 8553 17925 8587 17959
rect 8621 17925 8655 17959
rect 8689 17925 8723 17959
rect 8757 17925 8791 17959
rect 8825 17925 8859 17959
rect 8893 17925 8927 17959
rect 8961 17925 8995 17959
rect 9029 17925 9063 17959
rect 9097 17925 9131 17959
rect 9165 17925 9199 17959
rect 9233 17925 9267 17959
rect 9301 17925 9335 17959
rect 9369 17925 9403 17959
rect 9437 17925 9471 17959
rect 9505 17925 9539 17959
rect 9573 17925 9607 17959
rect 9641 17925 9675 17959
rect 9709 17925 9743 17959
rect 9777 17925 9811 17959
rect 9845 17925 9879 17959
rect 9913 17925 9947 17959
rect 9981 17925 10015 17959
rect 10049 17925 10083 17959
rect 10117 17925 10151 17959
rect 10185 17925 10219 17959
rect 10253 17925 10287 17959
rect 10321 17925 10355 17959
rect 10389 17925 10423 17959
rect 10457 17925 10491 17959
rect 10525 17925 10559 17959
rect 10593 17925 10627 17959
rect 10661 17925 10695 17959
rect 10729 17925 10763 17959
rect 10797 17925 10831 17959
rect 10865 17925 10899 17959
rect 10933 17925 10967 17959
rect 11001 17925 11035 17959
rect 11069 17925 11103 17959
rect 11137 17925 11171 17959
rect 11205 17925 11239 17959
rect 11273 17925 11307 17959
rect 11341 17925 11375 17959
rect 11409 17925 11443 17959
rect 11477 17925 11511 17959
rect 11545 17925 11579 17959
rect 11613 17925 11647 17959
rect 11681 17925 11715 17959
rect 11749 17925 11783 17959
rect 11817 17925 11851 17959
rect 11885 17925 11919 17959
rect 11953 17925 11987 17959
rect 12021 17925 12055 17959
rect 12089 17925 12123 17959
rect 12157 17925 12191 17959
rect 12225 17925 12259 17959
rect 12293 17925 12327 17959
rect 12361 17925 12395 17959
rect 12429 17925 12463 17959
rect 12497 17925 12531 17959
rect 12565 17925 12599 17959
rect 12633 17925 12667 17959
rect 12701 17925 12735 17959
rect 12769 17925 12803 17959
rect 12837 17925 12871 17959
rect 12905 17925 12939 17959
rect 12973 17925 13007 17959
rect 13041 17925 13075 17959
rect 13109 17925 13143 17959
rect 13177 17925 13211 17959
rect 13245 17925 13279 17959
rect 13313 17925 13347 17959
rect 13381 17925 13415 17959
rect 13449 17925 13483 17959
rect 13517 17925 13551 17959
rect 13585 17925 13619 17959
rect 13653 17925 13687 17959
rect 13721 17925 13755 17959
rect 13789 17925 13823 17959
rect 13857 17925 13891 17959
rect 13925 17925 13959 17959
rect 13993 17925 14027 17959
rect 14061 17925 14095 17959
rect 14129 17925 14163 17959
rect 14197 17925 14231 17959
rect 14265 17925 14299 17959
rect 14333 17925 14367 17959
rect 14401 17925 14435 17959
rect 14469 17925 14503 17959
rect 14537 17925 14571 17959
rect 14605 17925 14639 17959
rect 14673 17925 14707 17959
rect 14741 17925 14772 17959
rect 197 17889 14772 17925
rect 197 17855 221 17889
rect 255 17855 290 17889
rect 324 17855 359 17889
rect 393 17855 427 17889
rect 461 17855 495 17889
rect 529 17855 563 17889
rect 597 17855 631 17889
rect 665 17855 699 17889
rect 733 17855 767 17889
rect 801 17855 835 17889
rect 869 17855 903 17889
rect 937 17855 971 17889
rect 1005 17855 1039 17889
rect 1073 17855 1107 17889
rect 1141 17855 1175 17889
rect 1209 17855 1243 17889
rect 1277 17855 1311 17889
rect 1345 17855 1379 17889
rect 1413 17855 1447 17889
rect 1481 17855 1515 17889
rect 1549 17855 1583 17889
rect 1617 17855 1651 17889
rect 1685 17855 1719 17889
rect 1753 17855 1787 17889
rect 1821 17855 1855 17889
rect 1889 17855 1923 17889
rect 1957 17855 1991 17889
rect 2025 17855 2059 17889
rect 2093 17855 2127 17889
rect 2161 17855 2195 17889
rect 2229 17855 2263 17889
rect 2297 17855 2331 17889
rect 2365 17855 2399 17889
rect 2433 17855 2467 17889
rect 2501 17855 2535 17889
rect 2569 17855 2603 17889
rect 2637 17855 2671 17889
rect 2705 17855 2739 17889
rect 2773 17855 2807 17889
rect 2841 17855 2875 17889
rect 2909 17855 2943 17889
rect 2977 17855 3011 17889
rect 3045 17855 3079 17889
rect 3113 17855 3147 17889
rect 3181 17855 3215 17889
rect 3249 17855 3283 17889
rect 3317 17855 3351 17889
rect 3385 17855 3419 17889
rect 3453 17855 3487 17889
rect 3521 17855 3555 17889
rect 3589 17855 3623 17889
rect 3657 17855 3691 17889
rect 3725 17855 3759 17889
rect 3793 17855 3827 17889
rect 3861 17855 3895 17889
rect 3929 17855 3963 17889
rect 3997 17855 4031 17889
rect 4065 17855 4099 17889
rect 4133 17855 4167 17889
rect 4201 17855 4235 17889
rect 4269 17855 4303 17889
rect 4337 17855 4371 17889
rect 4405 17855 4439 17889
rect 4473 17855 4507 17889
rect 4541 17855 4575 17889
rect 4609 17855 4643 17889
rect 4677 17855 4711 17889
rect 4745 17855 4779 17889
rect 4813 17855 4847 17889
rect 4881 17855 4915 17889
rect 4949 17855 4983 17889
rect 5017 17855 5051 17889
rect 5085 17855 5119 17889
rect 5153 17855 5187 17889
rect 5221 17855 5255 17889
rect 5289 17855 5323 17889
rect 5357 17855 5391 17889
rect 5425 17855 5459 17889
rect 5493 17855 5527 17889
rect 5561 17855 5595 17889
rect 5629 17855 5663 17889
rect 5697 17855 5731 17889
rect 5765 17855 5799 17889
rect 5833 17855 5867 17889
rect 5901 17855 5935 17889
rect 5969 17855 6003 17889
rect 6037 17855 6071 17889
rect 6105 17855 6139 17889
rect 6173 17855 6207 17889
rect 6241 17855 6275 17889
rect 6309 17855 6343 17889
rect 6377 17855 6411 17889
rect 6445 17855 6479 17889
rect 6513 17855 6547 17889
rect 6581 17855 6615 17889
rect 6649 17855 6683 17889
rect 6717 17855 6751 17889
rect 6785 17855 6819 17889
rect 6853 17855 6887 17889
rect 6921 17855 6955 17889
rect 6989 17855 7023 17889
rect 7057 17855 7091 17889
rect 7125 17855 7159 17889
rect 7193 17855 7227 17889
rect 7261 17855 7295 17889
rect 7329 17855 7363 17889
rect 7397 17855 7431 17889
rect 7465 17855 7499 17889
rect 7533 17855 7567 17889
rect 7601 17855 7635 17889
rect 7669 17855 7703 17889
rect 7737 17855 7771 17889
rect 7805 17855 7839 17889
rect 7873 17855 7907 17889
rect 7941 17855 7975 17889
rect 8009 17855 8043 17889
rect 8077 17855 8111 17889
rect 8145 17855 8179 17889
rect 8213 17855 8247 17889
rect 8281 17855 8315 17889
rect 8349 17855 8383 17889
rect 8417 17855 8451 17889
rect 8485 17855 8519 17889
rect 8553 17855 8587 17889
rect 8621 17855 8655 17889
rect 8689 17855 8723 17889
rect 8757 17855 8791 17889
rect 8825 17855 8859 17889
rect 8893 17855 8927 17889
rect 8961 17855 8995 17889
rect 9029 17855 9063 17889
rect 9097 17855 9131 17889
rect 9165 17855 9199 17889
rect 9233 17855 9267 17889
rect 9301 17855 9335 17889
rect 9369 17855 9403 17889
rect 9437 17855 9471 17889
rect 9505 17855 9539 17889
rect 9573 17855 9607 17889
rect 9641 17855 9675 17889
rect 9709 17855 9743 17889
rect 9777 17855 9811 17889
rect 9845 17855 9879 17889
rect 9913 17855 9947 17889
rect 9981 17855 10015 17889
rect 10049 17855 10083 17889
rect 10117 17855 10151 17889
rect 10185 17855 10219 17889
rect 10253 17855 10287 17889
rect 10321 17855 10355 17889
rect 10389 17855 10423 17889
rect 10457 17855 10491 17889
rect 10525 17855 10559 17889
rect 10593 17855 10627 17889
rect 10661 17855 10695 17889
rect 10729 17855 10763 17889
rect 10797 17855 10831 17889
rect 10865 17855 10899 17889
rect 10933 17855 10967 17889
rect 11001 17855 11035 17889
rect 11069 17855 11103 17889
rect 11137 17855 11171 17889
rect 11205 17855 11239 17889
rect 11273 17855 11307 17889
rect 11341 17855 11375 17889
rect 11409 17855 11443 17889
rect 11477 17855 11511 17889
rect 11545 17855 11579 17889
rect 11613 17855 11647 17889
rect 11681 17855 11715 17889
rect 11749 17855 11783 17889
rect 11817 17855 11851 17889
rect 11885 17855 11919 17889
rect 11953 17855 11987 17889
rect 12021 17855 12055 17889
rect 12089 17855 12123 17889
rect 12157 17855 12191 17889
rect 12225 17855 12259 17889
rect 12293 17855 12327 17889
rect 12361 17855 12395 17889
rect 12429 17855 12463 17889
rect 12497 17855 12531 17889
rect 12565 17855 12599 17889
rect 12633 17855 12667 17889
rect 12701 17855 12735 17889
rect 12769 17855 12803 17889
rect 12837 17855 12871 17889
rect 12905 17855 12939 17889
rect 12973 17855 13007 17889
rect 13041 17855 13075 17889
rect 13109 17855 13143 17889
rect 13177 17855 13211 17889
rect 13245 17855 13279 17889
rect 13313 17855 13347 17889
rect 13381 17855 13415 17889
rect 13449 17855 13483 17889
rect 13517 17855 13551 17889
rect 13585 17855 13619 17889
rect 13653 17855 13687 17889
rect 13721 17855 13755 17889
rect 13789 17855 13823 17889
rect 13857 17855 13891 17889
rect 13925 17855 13959 17889
rect 13993 17855 14027 17889
rect 14061 17855 14095 17889
rect 14129 17855 14163 17889
rect 14197 17855 14231 17889
rect 14265 17855 14299 17889
rect 14333 17855 14367 17889
rect 14401 17855 14435 17889
rect 14469 17855 14503 17889
rect 14537 17855 14571 17889
rect 14605 17855 14639 17889
rect 14673 17855 14707 17889
rect 14741 17855 14772 17889
<< mvnsubdiff >>
rect 49 27376 14952 27410
rect 49 27342 83 27376
rect 117 27342 152 27376
rect 186 27342 221 27376
rect 255 27342 290 27376
rect 324 27342 359 27376
rect 393 27342 428 27376
rect 462 27342 497 27376
rect 531 27342 566 27376
rect 600 27342 635 27376
rect 669 27342 704 27376
rect 738 27342 773 27376
rect 807 27342 842 27376
rect 876 27342 911 27376
rect 945 27342 980 27376
rect 1014 27342 1049 27376
rect 1083 27342 1118 27376
rect 1152 27342 1187 27376
rect 1221 27342 1256 27376
rect 1290 27342 1325 27376
rect 1359 27342 1394 27376
rect 1428 27342 1463 27376
rect 1497 27342 1532 27376
rect 1566 27342 1601 27376
rect 1635 27342 1670 27376
rect 1704 27342 1739 27376
rect 1773 27342 1808 27376
rect 1842 27342 1877 27376
rect 1911 27342 1946 27376
rect 1980 27342 2014 27376
rect 2048 27342 2082 27376
rect 2116 27342 2150 27376
rect 2184 27342 2218 27376
rect 2252 27342 2286 27376
rect 2320 27342 2354 27376
rect 2388 27342 2422 27376
rect 2456 27342 2490 27376
rect 2524 27342 2558 27376
rect 2592 27342 2626 27376
rect 2660 27342 2694 27376
rect 2728 27342 2762 27376
rect 2796 27372 14952 27376
rect 2796 27342 2848 27372
rect 49 27338 2848 27342
rect 2882 27338 2916 27372
rect 2950 27338 2984 27372
rect 3018 27338 3052 27372
rect 3086 27338 3120 27372
rect 3154 27338 3188 27372
rect 3222 27338 3256 27372
rect 3290 27338 3324 27372
rect 3358 27338 3392 27372
rect 3426 27338 3460 27372
rect 3494 27338 3528 27372
rect 3562 27338 3596 27372
rect 3630 27338 3664 27372
rect 3698 27338 3732 27372
rect 3766 27338 3800 27372
rect 3834 27338 3868 27372
rect 3902 27338 3936 27372
rect 3970 27338 4004 27372
rect 4038 27338 4072 27372
rect 4106 27338 4140 27372
rect 4174 27338 4208 27372
rect 4242 27338 4276 27372
rect 4310 27338 4344 27372
rect 4378 27338 4412 27372
rect 4446 27338 4480 27372
rect 4514 27338 4548 27372
rect 4582 27338 4616 27372
rect 4650 27338 4684 27372
rect 4718 27338 4752 27372
rect 4786 27338 4820 27372
rect 4854 27338 4888 27372
rect 4922 27338 4956 27372
rect 4990 27338 5024 27372
rect 5058 27338 5092 27372
rect 5126 27338 5160 27372
rect 5194 27338 5228 27372
rect 5262 27338 5296 27372
rect 5330 27338 5364 27372
rect 5398 27338 5432 27372
rect 5466 27338 5500 27372
rect 5534 27338 5568 27372
rect 5602 27338 5636 27372
rect 5670 27338 5704 27372
rect 5738 27338 5772 27372
rect 5806 27338 5840 27372
rect 5874 27338 5908 27372
rect 5942 27338 5976 27372
rect 6010 27338 6044 27372
rect 6078 27338 6112 27372
rect 6146 27338 6180 27372
rect 6214 27338 6248 27372
rect 6282 27338 6316 27372
rect 6350 27338 6384 27372
rect 6418 27338 6452 27372
rect 6486 27338 6520 27372
rect 6554 27338 6588 27372
rect 6622 27338 6656 27372
rect 6690 27338 6724 27372
rect 6758 27338 6792 27372
rect 6826 27338 6860 27372
rect 6894 27338 6928 27372
rect 6962 27338 6996 27372
rect 7030 27338 7064 27372
rect 7098 27338 7132 27372
rect 7166 27338 7200 27372
rect 7234 27338 7268 27372
rect 7302 27338 7336 27372
rect 7370 27338 7404 27372
rect 7438 27338 7472 27372
rect 7506 27338 7540 27372
rect 7574 27338 7608 27372
rect 7642 27338 7676 27372
rect 7710 27338 7744 27372
rect 7778 27338 7812 27372
rect 7846 27338 7880 27372
rect 7914 27338 7948 27372
rect 7982 27338 8016 27372
rect 8050 27338 8084 27372
rect 8118 27338 8152 27372
rect 8186 27338 8220 27372
rect 8254 27338 8288 27372
rect 8322 27338 8356 27372
rect 8390 27338 8424 27372
rect 8458 27338 8492 27372
rect 8526 27338 8560 27372
rect 8594 27338 8628 27372
rect 8662 27338 8696 27372
rect 8730 27338 8764 27372
rect 8798 27338 8832 27372
rect 8866 27338 8900 27372
rect 8934 27338 8968 27372
rect 9002 27338 9036 27372
rect 9070 27338 9104 27372
rect 9138 27338 9172 27372
rect 9206 27338 9240 27372
rect 9274 27338 9308 27372
rect 9342 27338 9376 27372
rect 9410 27338 9444 27372
rect 9478 27338 9512 27372
rect 9546 27338 9580 27372
rect 9614 27338 9648 27372
rect 9682 27338 9716 27372
rect 9750 27338 9784 27372
rect 9818 27338 9852 27372
rect 9886 27338 9920 27372
rect 9954 27338 9988 27372
rect 10022 27338 10056 27372
rect 10090 27338 10124 27372
rect 10158 27338 10192 27372
rect 10226 27338 10260 27372
rect 10294 27338 10328 27372
rect 10362 27338 10396 27372
rect 10430 27338 10464 27372
rect 10498 27338 10532 27372
rect 10566 27338 10600 27372
rect 10634 27338 10668 27372
rect 10702 27338 10736 27372
rect 10770 27338 10804 27372
rect 10838 27338 10872 27372
rect 10906 27338 10940 27372
rect 10974 27338 11008 27372
rect 11042 27338 11076 27372
rect 11110 27338 11144 27372
rect 11178 27338 11212 27372
rect 11246 27338 11280 27372
rect 11314 27338 11348 27372
rect 11382 27338 11416 27372
rect 11450 27338 11484 27372
rect 11518 27338 11552 27372
rect 11586 27338 11620 27372
rect 11654 27338 11688 27372
rect 11722 27338 11756 27372
rect 11790 27338 11824 27372
rect 11858 27338 11892 27372
rect 11926 27338 11960 27372
rect 11994 27338 12028 27372
rect 12062 27338 12096 27372
rect 12130 27338 12164 27372
rect 12198 27338 12232 27372
rect 12266 27338 12300 27372
rect 12334 27338 12368 27372
rect 12402 27338 12436 27372
rect 12470 27338 12504 27372
rect 12538 27338 12572 27372
rect 12606 27338 12640 27372
rect 12674 27338 12708 27372
rect 12742 27338 12776 27372
rect 12810 27338 12844 27372
rect 12878 27338 12912 27372
rect 12946 27338 12980 27372
rect 13014 27338 13048 27372
rect 13082 27338 13116 27372
rect 13150 27338 13184 27372
rect 13218 27338 13252 27372
rect 13286 27338 13320 27372
rect 13354 27338 13388 27372
rect 13422 27338 13456 27372
rect 13490 27338 13524 27372
rect 13558 27338 13592 27372
rect 13626 27338 13660 27372
rect 13694 27338 13728 27372
rect 13762 27338 13796 27372
rect 13830 27338 13864 27372
rect 13898 27338 13932 27372
rect 13966 27338 14000 27372
rect 14034 27338 14068 27372
rect 14102 27338 14136 27372
rect 14170 27338 14204 27372
rect 14238 27338 14272 27372
rect 14306 27338 14340 27372
rect 14374 27338 14408 27372
rect 14442 27338 14476 27372
rect 14510 27338 14544 27372
rect 14578 27338 14612 27372
rect 14646 27338 14680 27372
rect 14714 27338 14748 27372
rect 14782 27338 14816 27372
rect 14850 27338 14884 27372
rect 14918 27338 14952 27372
rect 49 27302 14952 27338
rect 49 27268 83 27302
rect 117 27268 152 27302
rect 186 27268 221 27302
rect 255 27268 290 27302
rect 324 27268 359 27302
rect 393 27268 428 27302
rect 462 27268 497 27302
rect 531 27268 566 27302
rect 600 27268 635 27302
rect 669 27268 704 27302
rect 738 27268 773 27302
rect 807 27268 842 27302
rect 876 27268 911 27302
rect 945 27268 980 27302
rect 1014 27268 1049 27302
rect 1083 27268 1118 27302
rect 1152 27268 1187 27302
rect 1221 27268 1256 27302
rect 1290 27268 1325 27302
rect 1359 27268 1394 27302
rect 1428 27268 1463 27302
rect 1497 27268 1532 27302
rect 1566 27268 1601 27302
rect 1635 27268 1670 27302
rect 1704 27268 1739 27302
rect 1773 27268 1808 27302
rect 1842 27268 1877 27302
rect 1911 27268 1946 27302
rect 1980 27268 2014 27302
rect 2048 27268 2082 27302
rect 2116 27268 2150 27302
rect 2184 27268 2218 27302
rect 2252 27268 2286 27302
rect 2320 27268 2354 27302
rect 2388 27268 2422 27302
rect 2456 27268 2490 27302
rect 2524 27268 2558 27302
rect 2592 27268 2626 27302
rect 2660 27268 2694 27302
rect 2728 27268 2762 27302
rect 2796 27268 2848 27302
rect 2882 27268 2916 27302
rect 2950 27268 2984 27302
rect 3018 27268 3052 27302
rect 3086 27268 3120 27302
rect 3154 27268 3188 27302
rect 3222 27268 3256 27302
rect 3290 27268 3324 27302
rect 3358 27268 3392 27302
rect 3426 27268 3460 27302
rect 3494 27268 3528 27302
rect 3562 27268 3596 27302
rect 3630 27268 3664 27302
rect 3698 27268 3732 27302
rect 3766 27268 3800 27302
rect 3834 27268 3868 27302
rect 3902 27268 3936 27302
rect 3970 27268 4004 27302
rect 4038 27268 4072 27302
rect 4106 27268 4140 27302
rect 4174 27268 4208 27302
rect 4242 27268 4276 27302
rect 4310 27268 4344 27302
rect 4378 27268 4412 27302
rect 4446 27268 4480 27302
rect 4514 27268 4548 27302
rect 4582 27268 4616 27302
rect 4650 27268 4684 27302
rect 4718 27268 4752 27302
rect 4786 27268 4820 27302
rect 4854 27268 4888 27302
rect 4922 27268 4956 27302
rect 4990 27268 5024 27302
rect 5058 27268 5092 27302
rect 5126 27268 5160 27302
rect 5194 27268 5228 27302
rect 5262 27268 5296 27302
rect 5330 27268 5364 27302
rect 5398 27268 5432 27302
rect 5466 27268 5500 27302
rect 5534 27268 5568 27302
rect 5602 27268 5636 27302
rect 5670 27268 5704 27302
rect 5738 27268 5772 27302
rect 5806 27268 5840 27302
rect 5874 27268 5908 27302
rect 5942 27268 5976 27302
rect 6010 27268 6044 27302
rect 6078 27268 6112 27302
rect 6146 27268 6180 27302
rect 6214 27268 6248 27302
rect 6282 27268 6316 27302
rect 6350 27268 6384 27302
rect 6418 27268 6452 27302
rect 6486 27268 6520 27302
rect 6554 27268 6588 27302
rect 6622 27268 6656 27302
rect 6690 27268 6724 27302
rect 6758 27268 6792 27302
rect 6826 27268 6860 27302
rect 6894 27268 6928 27302
rect 6962 27268 6996 27302
rect 7030 27268 7064 27302
rect 7098 27268 7132 27302
rect 7166 27268 7200 27302
rect 7234 27268 7268 27302
rect 7302 27268 7336 27302
rect 7370 27268 7404 27302
rect 7438 27268 7472 27302
rect 7506 27268 7540 27302
rect 7574 27268 7608 27302
rect 7642 27268 7676 27302
rect 7710 27268 7744 27302
rect 7778 27268 7812 27302
rect 7846 27268 7880 27302
rect 7914 27268 7948 27302
rect 7982 27268 8016 27302
rect 8050 27268 8084 27302
rect 8118 27268 8152 27302
rect 8186 27268 8220 27302
rect 8254 27268 8288 27302
rect 8322 27268 8356 27302
rect 8390 27268 8424 27302
rect 8458 27268 8492 27302
rect 8526 27268 8560 27302
rect 8594 27268 8628 27302
rect 8662 27268 8696 27302
rect 8730 27268 8764 27302
rect 8798 27268 8832 27302
rect 8866 27268 8900 27302
rect 8934 27268 8968 27302
rect 9002 27268 9036 27302
rect 9070 27268 9104 27302
rect 9138 27268 9172 27302
rect 9206 27268 9240 27302
rect 9274 27268 9308 27302
rect 9342 27268 9376 27302
rect 9410 27268 9444 27302
rect 9478 27268 9512 27302
rect 9546 27268 9580 27302
rect 9614 27268 9648 27302
rect 9682 27268 9716 27302
rect 9750 27268 9784 27302
rect 9818 27268 9852 27302
rect 9886 27268 9920 27302
rect 9954 27268 9988 27302
rect 10022 27268 10056 27302
rect 10090 27268 10124 27302
rect 10158 27268 10192 27302
rect 10226 27268 10260 27302
rect 10294 27268 10328 27302
rect 10362 27268 10396 27302
rect 10430 27268 10464 27302
rect 10498 27268 10532 27302
rect 10566 27268 10600 27302
rect 10634 27268 10668 27302
rect 10702 27268 10736 27302
rect 10770 27268 10804 27302
rect 10838 27268 10872 27302
rect 10906 27268 10940 27302
rect 10974 27268 11008 27302
rect 11042 27268 11076 27302
rect 11110 27268 11144 27302
rect 11178 27268 11212 27302
rect 11246 27268 11280 27302
rect 11314 27268 11348 27302
rect 11382 27268 11416 27302
rect 11450 27268 11484 27302
rect 11518 27268 11552 27302
rect 11586 27268 11620 27302
rect 11654 27268 11688 27302
rect 11722 27268 11756 27302
rect 11790 27268 11824 27302
rect 11858 27268 11892 27302
rect 11926 27268 11960 27302
rect 11994 27268 12028 27302
rect 12062 27268 12096 27302
rect 12130 27268 12164 27302
rect 12198 27268 12232 27302
rect 12266 27268 12300 27302
rect 12334 27268 12368 27302
rect 12402 27268 12436 27302
rect 12470 27268 12504 27302
rect 12538 27268 12572 27302
rect 12606 27268 12640 27302
rect 12674 27268 12708 27302
rect 12742 27268 12776 27302
rect 12810 27268 12844 27302
rect 12878 27268 12912 27302
rect 12946 27268 12980 27302
rect 13014 27268 13048 27302
rect 13082 27268 13116 27302
rect 13150 27268 13184 27302
rect 13218 27268 13252 27302
rect 13286 27268 13320 27302
rect 13354 27268 13388 27302
rect 13422 27268 13456 27302
rect 13490 27268 13524 27302
rect 13558 27268 13592 27302
rect 13626 27268 13660 27302
rect 13694 27268 13728 27302
rect 13762 27268 13796 27302
rect 13830 27268 13864 27302
rect 13898 27268 13932 27302
rect 13966 27268 14000 27302
rect 14034 27268 14068 27302
rect 14102 27268 14136 27302
rect 14170 27268 14204 27302
rect 14238 27268 14272 27302
rect 14306 27268 14340 27302
rect 14374 27268 14408 27302
rect 14442 27268 14476 27302
rect 14510 27268 14544 27302
rect 14578 27268 14612 27302
rect 14646 27268 14680 27302
rect 14714 27268 14748 27302
rect 14782 27268 14816 27302
rect 14850 27268 14884 27302
rect 14918 27268 14952 27302
rect 49 27232 14952 27268
rect 49 27228 2848 27232
rect 49 27194 83 27228
rect 117 27194 152 27228
rect 186 27194 221 27228
rect 255 27194 290 27228
rect 324 27194 359 27228
rect 393 27194 428 27228
rect 462 27194 497 27228
rect 531 27194 566 27228
rect 600 27194 635 27228
rect 669 27194 704 27228
rect 738 27194 773 27228
rect 807 27194 842 27228
rect 876 27194 911 27228
rect 945 27194 980 27228
rect 1014 27194 1049 27228
rect 1083 27194 1118 27228
rect 1152 27194 1187 27228
rect 1221 27194 1256 27228
rect 1290 27194 1325 27228
rect 1359 27194 1394 27228
rect 1428 27194 1463 27228
rect 1497 27194 1532 27228
rect 1566 27194 1601 27228
rect 1635 27194 1670 27228
rect 1704 27194 1739 27228
rect 1773 27194 1808 27228
rect 1842 27194 1877 27228
rect 1911 27194 1946 27228
rect 1980 27194 2014 27228
rect 2048 27194 2082 27228
rect 2116 27194 2150 27228
rect 2184 27194 2218 27228
rect 2252 27194 2286 27228
rect 2320 27194 2354 27228
rect 2388 27194 2422 27228
rect 2456 27194 2490 27228
rect 2524 27194 2558 27228
rect 2592 27194 2626 27228
rect 2660 27194 2694 27228
rect 2728 27194 2762 27228
rect 2796 27198 2848 27228
rect 2882 27198 2916 27232
rect 2950 27198 2984 27232
rect 3018 27198 3052 27232
rect 3086 27198 3120 27232
rect 3154 27198 3188 27232
rect 3222 27198 3256 27232
rect 3290 27198 3324 27232
rect 3358 27198 3392 27232
rect 3426 27198 3460 27232
rect 3494 27198 3528 27232
rect 3562 27198 3596 27232
rect 3630 27198 3664 27232
rect 3698 27198 3732 27232
rect 3766 27198 3800 27232
rect 3834 27198 3868 27232
rect 3902 27198 3936 27232
rect 3970 27198 4004 27232
rect 4038 27198 4072 27232
rect 4106 27198 4140 27232
rect 4174 27198 4208 27232
rect 4242 27198 4276 27232
rect 4310 27198 4344 27232
rect 4378 27198 4412 27232
rect 4446 27198 4480 27232
rect 4514 27198 4548 27232
rect 4582 27198 4616 27232
rect 4650 27198 4684 27232
rect 4718 27198 4752 27232
rect 4786 27198 4820 27232
rect 4854 27198 4888 27232
rect 4922 27198 4956 27232
rect 4990 27198 5024 27232
rect 5058 27198 5092 27232
rect 5126 27198 5160 27232
rect 5194 27198 5228 27232
rect 5262 27198 5296 27232
rect 5330 27198 5364 27232
rect 5398 27198 5432 27232
rect 5466 27198 5500 27232
rect 5534 27198 5568 27232
rect 5602 27198 5636 27232
rect 5670 27198 5704 27232
rect 5738 27198 5772 27232
rect 5806 27198 5840 27232
rect 5874 27198 5908 27232
rect 5942 27198 5976 27232
rect 6010 27198 6044 27232
rect 6078 27198 6112 27232
rect 6146 27198 6180 27232
rect 6214 27198 6248 27232
rect 6282 27198 6316 27232
rect 6350 27198 6384 27232
rect 6418 27198 6452 27232
rect 6486 27198 6520 27232
rect 6554 27198 6588 27232
rect 6622 27198 6656 27232
rect 6690 27198 6724 27232
rect 6758 27198 6792 27232
rect 6826 27198 6860 27232
rect 6894 27198 6928 27232
rect 6962 27198 6996 27232
rect 7030 27198 7064 27232
rect 7098 27198 7132 27232
rect 7166 27198 7200 27232
rect 7234 27198 7268 27232
rect 7302 27198 7336 27232
rect 7370 27198 7404 27232
rect 7438 27198 7472 27232
rect 7506 27198 7540 27232
rect 7574 27198 7608 27232
rect 7642 27198 7676 27232
rect 7710 27198 7744 27232
rect 7778 27198 7812 27232
rect 7846 27198 7880 27232
rect 7914 27198 7948 27232
rect 7982 27198 8016 27232
rect 8050 27198 8084 27232
rect 8118 27198 8152 27232
rect 8186 27198 8220 27232
rect 8254 27198 8288 27232
rect 8322 27198 8356 27232
rect 8390 27198 8424 27232
rect 8458 27198 8492 27232
rect 8526 27198 8560 27232
rect 8594 27198 8628 27232
rect 8662 27198 8696 27232
rect 8730 27198 8764 27232
rect 8798 27198 8832 27232
rect 8866 27198 8900 27232
rect 8934 27198 8968 27232
rect 9002 27198 9036 27232
rect 9070 27198 9104 27232
rect 9138 27198 9172 27232
rect 9206 27198 9240 27232
rect 9274 27198 9308 27232
rect 9342 27198 9376 27232
rect 9410 27198 9444 27232
rect 9478 27198 9512 27232
rect 9546 27198 9580 27232
rect 9614 27198 9648 27232
rect 9682 27198 9716 27232
rect 9750 27198 9784 27232
rect 9818 27198 9852 27232
rect 9886 27198 9920 27232
rect 9954 27198 9988 27232
rect 10022 27198 10056 27232
rect 10090 27198 10124 27232
rect 10158 27198 10192 27232
rect 10226 27198 10260 27232
rect 10294 27198 10328 27232
rect 10362 27198 10396 27232
rect 10430 27198 10464 27232
rect 10498 27198 10532 27232
rect 10566 27198 10600 27232
rect 10634 27198 10668 27232
rect 10702 27198 10736 27232
rect 10770 27198 10804 27232
rect 10838 27198 10872 27232
rect 10906 27198 10940 27232
rect 10974 27198 11008 27232
rect 11042 27198 11076 27232
rect 11110 27198 11144 27232
rect 11178 27198 11212 27232
rect 11246 27198 11280 27232
rect 11314 27198 11348 27232
rect 11382 27198 11416 27232
rect 11450 27198 11484 27232
rect 11518 27198 11552 27232
rect 11586 27198 11620 27232
rect 11654 27198 11688 27232
rect 11722 27198 11756 27232
rect 11790 27198 11824 27232
rect 11858 27198 11892 27232
rect 11926 27198 11960 27232
rect 11994 27198 12028 27232
rect 12062 27198 12096 27232
rect 12130 27198 12164 27232
rect 12198 27198 12232 27232
rect 12266 27198 12300 27232
rect 12334 27198 12368 27232
rect 12402 27198 12436 27232
rect 12470 27198 12504 27232
rect 12538 27198 12572 27232
rect 12606 27198 12640 27232
rect 12674 27198 12708 27232
rect 12742 27198 12776 27232
rect 12810 27198 12844 27232
rect 12878 27198 12912 27232
rect 12946 27198 12980 27232
rect 13014 27198 13048 27232
rect 13082 27198 13116 27232
rect 13150 27198 13184 27232
rect 13218 27198 13252 27232
rect 13286 27198 13320 27232
rect 13354 27198 13388 27232
rect 13422 27198 13456 27232
rect 13490 27198 13524 27232
rect 13558 27198 13592 27232
rect 13626 27198 13660 27232
rect 13694 27198 13728 27232
rect 13762 27198 13796 27232
rect 13830 27198 13864 27232
rect 13898 27198 13932 27232
rect 13966 27198 14000 27232
rect 14034 27198 14068 27232
rect 14102 27198 14136 27232
rect 14170 27198 14204 27232
rect 14238 27198 14272 27232
rect 14306 27198 14340 27232
rect 14374 27198 14408 27232
rect 14442 27198 14476 27232
rect 14510 27198 14544 27232
rect 14578 27198 14612 27232
rect 14646 27198 14680 27232
rect 14714 27198 14748 27232
rect 14782 27198 14816 27232
rect 14850 27198 14884 27232
rect 14918 27198 14952 27232
rect 2796 27194 14952 27198
rect 49 27162 14952 27194
rect 49 27154 2848 27162
rect 49 27120 83 27154
rect 117 27120 152 27154
rect 186 27120 221 27154
rect 255 27120 290 27154
rect 324 27120 359 27154
rect 393 27120 428 27154
rect 462 27120 497 27154
rect 531 27120 566 27154
rect 600 27120 635 27154
rect 669 27120 704 27154
rect 738 27120 773 27154
rect 807 27120 842 27154
rect 876 27120 911 27154
rect 945 27120 980 27154
rect 1014 27120 1049 27154
rect 1083 27120 1118 27154
rect 1152 27120 1187 27154
rect 1221 27120 1256 27154
rect 1290 27120 1325 27154
rect 1359 27120 1394 27154
rect 1428 27120 1463 27154
rect 1497 27120 1532 27154
rect 1566 27120 1601 27154
rect 1635 27120 1670 27154
rect 1704 27120 1739 27154
rect 1773 27120 1808 27154
rect 1842 27120 1877 27154
rect 1911 27120 1946 27154
rect 1980 27120 2014 27154
rect 2048 27120 2082 27154
rect 2116 27120 2150 27154
rect 2184 27120 2218 27154
rect 2252 27120 2286 27154
rect 2320 27120 2354 27154
rect 2388 27120 2422 27154
rect 2456 27120 2490 27154
rect 2524 27120 2558 27154
rect 2592 27120 2626 27154
rect 2660 27120 2694 27154
rect 2728 27120 2762 27154
rect 2796 27128 2848 27154
rect 2882 27128 2916 27162
rect 2950 27128 2984 27162
rect 3018 27128 3052 27162
rect 3086 27128 3120 27162
rect 3154 27128 3188 27162
rect 3222 27128 3256 27162
rect 3290 27128 3324 27162
rect 3358 27128 3392 27162
rect 3426 27128 3460 27162
rect 3494 27128 3528 27162
rect 3562 27128 3596 27162
rect 3630 27128 3664 27162
rect 3698 27128 3732 27162
rect 3766 27128 3800 27162
rect 3834 27128 3868 27162
rect 3902 27128 3936 27162
rect 3970 27128 4004 27162
rect 4038 27128 4072 27162
rect 4106 27128 4140 27162
rect 4174 27128 4208 27162
rect 4242 27128 4276 27162
rect 4310 27128 4344 27162
rect 4378 27128 4412 27162
rect 4446 27128 4480 27162
rect 4514 27128 4548 27162
rect 4582 27128 4616 27162
rect 4650 27128 4684 27162
rect 4718 27128 4752 27162
rect 4786 27128 4820 27162
rect 4854 27128 4888 27162
rect 4922 27128 4956 27162
rect 4990 27128 5024 27162
rect 5058 27128 5092 27162
rect 5126 27128 5160 27162
rect 5194 27128 5228 27162
rect 5262 27128 5296 27162
rect 5330 27128 5364 27162
rect 5398 27128 5432 27162
rect 5466 27128 5500 27162
rect 5534 27128 5568 27162
rect 5602 27128 5636 27162
rect 5670 27128 5704 27162
rect 5738 27128 5772 27162
rect 5806 27128 5840 27162
rect 5874 27128 5908 27162
rect 5942 27128 5976 27162
rect 6010 27128 6044 27162
rect 6078 27128 6112 27162
rect 6146 27128 6180 27162
rect 6214 27128 6248 27162
rect 6282 27128 6316 27162
rect 6350 27128 6384 27162
rect 6418 27128 6452 27162
rect 6486 27128 6520 27162
rect 6554 27128 6588 27162
rect 6622 27128 6656 27162
rect 6690 27128 6724 27162
rect 6758 27128 6792 27162
rect 6826 27128 6860 27162
rect 6894 27128 6928 27162
rect 6962 27128 6996 27162
rect 7030 27128 7064 27162
rect 7098 27128 7132 27162
rect 7166 27128 7200 27162
rect 7234 27128 7268 27162
rect 7302 27128 7336 27162
rect 7370 27128 7404 27162
rect 7438 27128 7472 27162
rect 7506 27128 7540 27162
rect 7574 27128 7608 27162
rect 7642 27128 7676 27162
rect 7710 27128 7744 27162
rect 7778 27128 7812 27162
rect 7846 27128 7880 27162
rect 7914 27128 7948 27162
rect 7982 27128 8016 27162
rect 8050 27128 8084 27162
rect 8118 27128 8152 27162
rect 8186 27128 8220 27162
rect 8254 27128 8288 27162
rect 8322 27128 8356 27162
rect 8390 27128 8424 27162
rect 8458 27128 8492 27162
rect 8526 27128 8560 27162
rect 8594 27128 8628 27162
rect 8662 27128 8696 27162
rect 8730 27128 8764 27162
rect 8798 27128 8832 27162
rect 8866 27128 8900 27162
rect 8934 27128 8968 27162
rect 9002 27128 9036 27162
rect 9070 27128 9104 27162
rect 9138 27128 9172 27162
rect 9206 27128 9240 27162
rect 9274 27128 9308 27162
rect 9342 27128 9376 27162
rect 9410 27128 9444 27162
rect 9478 27128 9512 27162
rect 9546 27128 9580 27162
rect 9614 27128 9648 27162
rect 9682 27128 9716 27162
rect 9750 27128 9784 27162
rect 9818 27128 9852 27162
rect 9886 27128 9920 27162
rect 9954 27128 9988 27162
rect 10022 27128 10056 27162
rect 10090 27128 10124 27162
rect 10158 27128 10192 27162
rect 10226 27128 10260 27162
rect 10294 27128 10328 27162
rect 10362 27128 10396 27162
rect 10430 27128 10464 27162
rect 10498 27128 10532 27162
rect 10566 27128 10600 27162
rect 10634 27128 10668 27162
rect 10702 27128 10736 27162
rect 10770 27128 10804 27162
rect 10838 27128 10872 27162
rect 10906 27128 10940 27162
rect 10974 27128 11008 27162
rect 11042 27128 11076 27162
rect 11110 27128 11144 27162
rect 11178 27128 11212 27162
rect 11246 27128 11280 27162
rect 11314 27128 11348 27162
rect 11382 27128 11416 27162
rect 11450 27128 11484 27162
rect 11518 27128 11552 27162
rect 11586 27128 11620 27162
rect 11654 27128 11688 27162
rect 11722 27128 11756 27162
rect 11790 27128 11824 27162
rect 11858 27128 11892 27162
rect 11926 27128 11960 27162
rect 11994 27128 12028 27162
rect 12062 27128 12096 27162
rect 12130 27128 12164 27162
rect 12198 27128 12232 27162
rect 12266 27128 12300 27162
rect 12334 27128 12368 27162
rect 12402 27128 12436 27162
rect 12470 27128 12504 27162
rect 12538 27128 12572 27162
rect 12606 27128 12640 27162
rect 12674 27128 12708 27162
rect 12742 27128 12776 27162
rect 12810 27128 12844 27162
rect 12878 27128 12912 27162
rect 12946 27128 12980 27162
rect 13014 27128 13048 27162
rect 13082 27128 13116 27162
rect 13150 27128 13184 27162
rect 13218 27128 13252 27162
rect 13286 27128 13320 27162
rect 13354 27128 13388 27162
rect 13422 27128 13456 27162
rect 13490 27128 13524 27162
rect 13558 27128 13592 27162
rect 13626 27128 13660 27162
rect 13694 27128 13728 27162
rect 13762 27128 13796 27162
rect 13830 27128 13864 27162
rect 13898 27128 13932 27162
rect 13966 27128 14000 27162
rect 14034 27128 14068 27162
rect 14102 27128 14136 27162
rect 14170 27128 14204 27162
rect 14238 27128 14272 27162
rect 14306 27128 14340 27162
rect 14374 27128 14408 27162
rect 14442 27128 14476 27162
rect 14510 27128 14544 27162
rect 14578 27128 14612 27162
rect 14646 27128 14680 27162
rect 14714 27128 14748 27162
rect 14782 27128 14816 27162
rect 14850 27128 14884 27162
rect 14918 27128 14952 27162
rect 2796 27120 14952 27128
rect 49 27092 14952 27120
rect 49 27086 2848 27092
rect 49 26794 151 27086
rect 2814 27058 2848 27086
rect 2882 27058 2916 27092
rect 2950 27058 2984 27092
rect 3018 27058 3052 27092
rect 3086 27058 3120 27092
rect 3154 27058 3188 27092
rect 3222 27058 3256 27092
rect 3290 27058 3324 27092
rect 3358 27058 3392 27092
rect 3426 27058 3460 27092
rect 3494 27058 3528 27092
rect 3562 27058 3596 27092
rect 3630 27058 3664 27092
rect 3698 27058 3732 27092
rect 3766 27058 3800 27092
rect 3834 27058 3868 27092
rect 3902 27058 3936 27092
rect 3970 27058 4004 27092
rect 4038 27058 4072 27092
rect 4106 27058 4140 27092
rect 4174 27058 4208 27092
rect 4242 27058 4276 27092
rect 4310 27058 4344 27092
rect 4378 27058 4412 27092
rect 4446 27058 4480 27092
rect 4514 27058 4548 27092
rect 4582 27058 4616 27092
rect 4650 27058 4684 27092
rect 4718 27058 4752 27092
rect 4786 27058 4820 27092
rect 4854 27058 4888 27092
rect 4922 27058 4956 27092
rect 4990 27058 5024 27092
rect 5058 27058 5092 27092
rect 5126 27058 5160 27092
rect 5194 27058 5228 27092
rect 5262 27058 5296 27092
rect 5330 27058 5364 27092
rect 5398 27058 5432 27092
rect 5466 27058 5500 27092
rect 5534 27058 5568 27092
rect 5602 27058 5636 27092
rect 5670 27058 5704 27092
rect 5738 27058 5772 27092
rect 5806 27058 5840 27092
rect 5874 27058 5908 27092
rect 5942 27058 5976 27092
rect 6010 27058 6044 27092
rect 6078 27058 6112 27092
rect 6146 27058 6180 27092
rect 6214 27058 6248 27092
rect 6282 27058 6316 27092
rect 6350 27058 6384 27092
rect 6418 27058 6452 27092
rect 6486 27058 6520 27092
rect 6554 27058 6588 27092
rect 6622 27058 6656 27092
rect 6690 27058 6724 27092
rect 6758 27058 6792 27092
rect 6826 27058 6860 27092
rect 6894 27058 6928 27092
rect 6962 27058 6996 27092
rect 7030 27058 7064 27092
rect 7098 27058 7132 27092
rect 7166 27058 7200 27092
rect 7234 27058 7268 27092
rect 7302 27058 7336 27092
rect 7370 27058 7404 27092
rect 7438 27058 7472 27092
rect 7506 27058 7540 27092
rect 7574 27058 7608 27092
rect 7642 27058 7676 27092
rect 7710 27058 7744 27092
rect 7778 27058 7812 27092
rect 7846 27058 7880 27092
rect 7914 27058 7948 27092
rect 7982 27058 8016 27092
rect 8050 27058 8084 27092
rect 8118 27058 8152 27092
rect 8186 27058 8220 27092
rect 8254 27058 8288 27092
rect 8322 27058 8356 27092
rect 8390 27058 8424 27092
rect 8458 27058 8492 27092
rect 8526 27058 8560 27092
rect 8594 27058 8628 27092
rect 8662 27058 8696 27092
rect 8730 27058 8764 27092
rect 8798 27058 8832 27092
rect 8866 27058 8900 27092
rect 8934 27058 8968 27092
rect 9002 27058 9036 27092
rect 9070 27058 9104 27092
rect 9138 27058 9172 27092
rect 9206 27058 9240 27092
rect 9274 27058 9308 27092
rect 9342 27058 9376 27092
rect 9410 27058 9444 27092
rect 9478 27058 9512 27092
rect 9546 27058 9580 27092
rect 9614 27058 9648 27092
rect 9682 27058 9716 27092
rect 9750 27058 9784 27092
rect 9818 27058 9852 27092
rect 9886 27058 9920 27092
rect 9954 27058 9988 27092
rect 10022 27058 10056 27092
rect 10090 27058 10124 27092
rect 10158 27058 10192 27092
rect 10226 27058 10260 27092
rect 10294 27058 10328 27092
rect 10362 27058 10396 27092
rect 10430 27058 10464 27092
rect 10498 27058 10532 27092
rect 10566 27058 10600 27092
rect 10634 27058 10668 27092
rect 10702 27058 10736 27092
rect 10770 27058 10804 27092
rect 10838 27058 10872 27092
rect 10906 27058 10940 27092
rect 10974 27058 11008 27092
rect 11042 27058 11076 27092
rect 11110 27058 11144 27092
rect 11178 27058 11212 27092
rect 11246 27058 11280 27092
rect 11314 27058 11348 27092
rect 11382 27058 11416 27092
rect 11450 27058 11484 27092
rect 11518 27058 11552 27092
rect 11586 27058 11620 27092
rect 11654 27058 11688 27092
rect 11722 27058 11756 27092
rect 11790 27058 11824 27092
rect 11858 27058 11892 27092
rect 11926 27058 11960 27092
rect 11994 27058 12028 27092
rect 12062 27058 12096 27092
rect 12130 27058 12164 27092
rect 12198 27058 12232 27092
rect 12266 27058 12300 27092
rect 12334 27058 12368 27092
rect 12402 27058 12436 27092
rect 12470 27058 12504 27092
rect 12538 27058 12572 27092
rect 12606 27058 12640 27092
rect 12674 27058 12708 27092
rect 12742 27058 12776 27092
rect 12810 27058 12844 27092
rect 12878 27058 12912 27092
rect 12946 27058 12980 27092
rect 13014 27058 13048 27092
rect 13082 27058 13116 27092
rect 13150 27058 13184 27092
rect 13218 27058 13252 27092
rect 13286 27058 13320 27092
rect 13354 27058 13388 27092
rect 13422 27058 13456 27092
rect 13490 27058 13524 27092
rect 13558 27058 13592 27092
rect 13626 27058 13660 27092
rect 13694 27058 13728 27092
rect 13762 27058 13796 27092
rect 13830 27058 13864 27092
rect 13898 27058 13932 27092
rect 13966 27058 14000 27092
rect 14034 27058 14068 27092
rect 14102 27058 14136 27092
rect 14170 27058 14204 27092
rect 14238 27058 14272 27092
rect 14306 27058 14340 27092
rect 14374 27058 14408 27092
rect 14442 27058 14476 27092
rect 14510 27058 14544 27092
rect 14578 27058 14612 27092
rect 14646 27058 14680 27092
rect 14714 27058 14748 27092
rect 14782 27058 14816 27092
rect 14850 27058 14884 27092
rect 14918 27058 14952 27092
rect 2814 27022 14952 27058
rect 2814 26988 2848 27022
rect 2882 26988 2916 27022
rect 2950 26988 2984 27022
rect 3018 26988 3052 27022
rect 3086 26988 3120 27022
rect 3154 26988 3188 27022
rect 3222 26988 3256 27022
rect 3290 26988 3324 27022
rect 3358 26988 3392 27022
rect 3426 26988 3460 27022
rect 3494 26988 3528 27022
rect 3562 26988 3596 27022
rect 3630 26988 3664 27022
rect 3698 26988 3732 27022
rect 3766 26988 3800 27022
rect 3834 26988 3868 27022
rect 3902 26988 3936 27022
rect 3970 26988 4004 27022
rect 4038 26988 4072 27022
rect 4106 26988 4140 27022
rect 4174 26988 4208 27022
rect 4242 26988 4276 27022
rect 4310 26988 4344 27022
rect 4378 26988 4412 27022
rect 4446 26988 4480 27022
rect 4514 26988 4548 27022
rect 4582 26988 4616 27022
rect 4650 26988 4684 27022
rect 4718 26988 4752 27022
rect 4786 26988 4820 27022
rect 4854 26988 4888 27022
rect 4922 26988 4956 27022
rect 4990 26988 5024 27022
rect 5058 26988 5092 27022
rect 5126 26988 5160 27022
rect 5194 26988 5228 27022
rect 5262 26988 5296 27022
rect 5330 26988 5364 27022
rect 5398 26988 5432 27022
rect 5466 26988 5500 27022
rect 5534 26988 5568 27022
rect 5602 26988 5636 27022
rect 5670 26988 5704 27022
rect 5738 26988 5772 27022
rect 5806 26988 5840 27022
rect 5874 26988 5908 27022
rect 5942 26988 5976 27022
rect 6010 26988 6044 27022
rect 6078 26988 6112 27022
rect 6146 26988 6180 27022
rect 6214 26988 6248 27022
rect 6282 26988 6316 27022
rect 6350 26988 6384 27022
rect 6418 26988 6452 27022
rect 6486 26988 6520 27022
rect 6554 26988 6588 27022
rect 6622 26988 6656 27022
rect 6690 26988 6724 27022
rect 6758 26988 6792 27022
rect 6826 26988 6860 27022
rect 6894 26988 6928 27022
rect 6962 26988 6996 27022
rect 7030 26988 7064 27022
rect 7098 26988 7132 27022
rect 7166 26988 7200 27022
rect 7234 26988 7268 27022
rect 7302 26988 7336 27022
rect 7370 26988 7404 27022
rect 7438 26988 7472 27022
rect 7506 26988 7540 27022
rect 7574 26988 7608 27022
rect 7642 26988 7676 27022
rect 7710 26988 7744 27022
rect 7778 26988 7812 27022
rect 7846 26988 7880 27022
rect 7914 26988 7948 27022
rect 7982 26988 8016 27022
rect 8050 26988 8084 27022
rect 8118 26988 8152 27022
rect 8186 26988 8220 27022
rect 8254 26988 8288 27022
rect 8322 26988 8356 27022
rect 8390 26988 8424 27022
rect 8458 26988 8492 27022
rect 8526 26988 8560 27022
rect 8594 26988 8628 27022
rect 8662 26988 8696 27022
rect 8730 26988 8764 27022
rect 8798 26988 8832 27022
rect 8866 26988 8900 27022
rect 8934 26988 8968 27022
rect 9002 26988 9036 27022
rect 9070 26988 9104 27022
rect 9138 26988 9172 27022
rect 9206 26988 9240 27022
rect 9274 26988 9308 27022
rect 9342 26988 9376 27022
rect 9410 26988 9444 27022
rect 9478 26988 9512 27022
rect 9546 26988 9580 27022
rect 9614 26988 9648 27022
rect 9682 26988 9716 27022
rect 9750 26988 9784 27022
rect 9818 26988 9852 27022
rect 9886 26988 9920 27022
rect 9954 26988 9988 27022
rect 10022 26988 10056 27022
rect 10090 26988 10124 27022
rect 10158 26988 10192 27022
rect 10226 26988 10260 27022
rect 10294 26988 10328 27022
rect 10362 26988 10396 27022
rect 10430 26988 10464 27022
rect 10498 26988 10532 27022
rect 10566 26988 10600 27022
rect 10634 26988 10668 27022
rect 10702 26988 10736 27022
rect 10770 26988 10804 27022
rect 10838 26988 10872 27022
rect 10906 26988 10940 27022
rect 10974 26988 11008 27022
rect 11042 26988 11076 27022
rect 11110 26988 11144 27022
rect 11178 26988 11212 27022
rect 11246 26988 11280 27022
rect 11314 26988 11348 27022
rect 11382 26988 11416 27022
rect 11450 26988 11484 27022
rect 11518 26988 11552 27022
rect 11586 26988 11620 27022
rect 11654 26988 11688 27022
rect 11722 26988 11756 27022
rect 11790 26988 11824 27022
rect 11858 26988 11892 27022
rect 11926 26988 11960 27022
rect 11994 26988 12028 27022
rect 12062 26988 12096 27022
rect 12130 26988 12164 27022
rect 12198 26988 12232 27022
rect 12266 26988 12300 27022
rect 12334 26988 12368 27022
rect 12402 26988 12436 27022
rect 12470 26988 12504 27022
rect 12538 26988 12572 27022
rect 12606 26988 12640 27022
rect 12674 26988 12708 27022
rect 12742 26988 12776 27022
rect 12810 26988 12844 27022
rect 12878 26988 12912 27022
rect 12946 26988 12980 27022
rect 13014 26988 13048 27022
rect 13082 26988 13116 27022
rect 13150 26988 13184 27022
rect 13218 26988 13252 27022
rect 13286 26988 13320 27022
rect 13354 26988 13388 27022
rect 13422 26988 13456 27022
rect 13490 26988 13524 27022
rect 13558 26988 13592 27022
rect 13626 26988 13660 27022
rect 13694 26988 13728 27022
rect 13762 26988 13796 27022
rect 13830 26988 13864 27022
rect 13898 26988 13932 27022
rect 13966 26988 14000 27022
rect 14034 26988 14068 27022
rect 14102 26988 14136 27022
rect 14170 26988 14204 27022
rect 14238 26988 14272 27022
rect 14306 26988 14340 27022
rect 14374 26988 14408 27022
rect 14442 26988 14476 27022
rect 14510 26988 14544 27022
rect 14578 26988 14612 27022
rect 14646 26988 14680 27022
rect 14714 26988 14748 27022
rect 14782 26988 14816 27022
rect 14850 26988 14884 27022
rect 14918 26988 14952 27022
rect 2814 26952 14952 26988
rect 2814 26918 2848 26952
rect 2882 26918 2916 26952
rect 2950 26918 2984 26952
rect 3018 26918 3052 26952
rect 3086 26918 3120 26952
rect 3154 26918 3188 26952
rect 3222 26918 3256 26952
rect 3290 26918 3324 26952
rect 3358 26918 3392 26952
rect 3426 26918 3460 26952
rect 3494 26918 3528 26952
rect 3562 26918 3596 26952
rect 3630 26918 3664 26952
rect 3698 26918 3732 26952
rect 3766 26918 3800 26952
rect 3834 26918 3868 26952
rect 3902 26918 3936 26952
rect 3970 26918 4004 26952
rect 4038 26918 4072 26952
rect 4106 26918 4140 26952
rect 4174 26918 4208 26952
rect 4242 26918 4276 26952
rect 4310 26918 4344 26952
rect 4378 26918 4412 26952
rect 4446 26918 4480 26952
rect 4514 26918 4548 26952
rect 4582 26918 4616 26952
rect 4650 26918 4684 26952
rect 4718 26918 4752 26952
rect 4786 26918 4820 26952
rect 4854 26918 4888 26952
rect 4922 26918 4956 26952
rect 4990 26918 5024 26952
rect 5058 26918 5092 26952
rect 5126 26918 5160 26952
rect 5194 26918 5228 26952
rect 5262 26918 5296 26952
rect 5330 26918 5364 26952
rect 5398 26918 5432 26952
rect 5466 26918 5500 26952
rect 5534 26918 5568 26952
rect 5602 26918 5636 26952
rect 5670 26918 5704 26952
rect 5738 26918 5772 26952
rect 5806 26918 5840 26952
rect 5874 26918 5908 26952
rect 5942 26918 5976 26952
rect 6010 26918 6044 26952
rect 6078 26918 6112 26952
rect 6146 26918 6180 26952
rect 6214 26918 6248 26952
rect 6282 26918 6316 26952
rect 6350 26918 6384 26952
rect 6418 26918 6452 26952
rect 6486 26918 6520 26952
rect 6554 26918 6588 26952
rect 6622 26918 6656 26952
rect 6690 26918 6724 26952
rect 6758 26918 6792 26952
rect 6826 26918 6860 26952
rect 6894 26918 6928 26952
rect 6962 26918 6996 26952
rect 7030 26918 7064 26952
rect 7098 26918 7132 26952
rect 7166 26918 7200 26952
rect 7234 26918 7268 26952
rect 7302 26918 7336 26952
rect 7370 26918 7404 26952
rect 7438 26918 7472 26952
rect 7506 26918 7540 26952
rect 7574 26918 7608 26952
rect 7642 26918 7676 26952
rect 7710 26918 7744 26952
rect 7778 26918 7812 26952
rect 7846 26918 7880 26952
rect 7914 26918 7948 26952
rect 7982 26918 8016 26952
rect 8050 26918 8084 26952
rect 8118 26918 8152 26952
rect 8186 26918 8220 26952
rect 8254 26918 8288 26952
rect 8322 26918 8356 26952
rect 8390 26918 8424 26952
rect 8458 26918 8492 26952
rect 8526 26918 8560 26952
rect 8594 26918 8628 26952
rect 8662 26918 8696 26952
rect 8730 26918 8764 26952
rect 8798 26918 8832 26952
rect 8866 26918 8900 26952
rect 8934 26918 8968 26952
rect 9002 26918 9036 26952
rect 9070 26918 9104 26952
rect 9138 26918 9172 26952
rect 9206 26918 9240 26952
rect 9274 26918 9308 26952
rect 9342 26918 9376 26952
rect 9410 26918 9444 26952
rect 9478 26918 9512 26952
rect 9546 26918 9580 26952
rect 9614 26918 9648 26952
rect 9682 26918 9716 26952
rect 9750 26918 9784 26952
rect 9818 26918 9852 26952
rect 9886 26918 9920 26952
rect 9954 26918 9988 26952
rect 10022 26918 10056 26952
rect 10090 26918 10124 26952
rect 10158 26918 10192 26952
rect 10226 26918 10260 26952
rect 10294 26918 10328 26952
rect 10362 26918 10396 26952
rect 10430 26918 10464 26952
rect 10498 26918 10532 26952
rect 10566 26918 10600 26952
rect 10634 26918 10668 26952
rect 10702 26918 10736 26952
rect 10770 26918 10804 26952
rect 10838 26918 10872 26952
rect 10906 26918 10940 26952
rect 10974 26918 11008 26952
rect 11042 26918 11076 26952
rect 11110 26918 11144 26952
rect 11178 26918 11212 26952
rect 11246 26918 11280 26952
rect 11314 26918 11348 26952
rect 11382 26918 11416 26952
rect 11450 26918 11484 26952
rect 11518 26918 11552 26952
rect 11586 26918 11620 26952
rect 11654 26918 11688 26952
rect 11722 26918 11756 26952
rect 11790 26918 11824 26952
rect 11858 26918 11892 26952
rect 11926 26918 11960 26952
rect 11994 26918 12028 26952
rect 12062 26918 12096 26952
rect 12130 26918 12164 26952
rect 12198 26918 12232 26952
rect 12266 26918 12300 26952
rect 12334 26918 12368 26952
rect 12402 26918 12436 26952
rect 12470 26918 12504 26952
rect 12538 26918 12572 26952
rect 12606 26918 12640 26952
rect 12674 26918 12708 26952
rect 12742 26918 12776 26952
rect 12810 26918 12844 26952
rect 12878 26918 12912 26952
rect 12946 26918 12980 26952
rect 13014 26918 13048 26952
rect 13082 26918 13116 26952
rect 13150 26918 13184 26952
rect 13218 26918 13252 26952
rect 13286 26918 13320 26952
rect 13354 26918 13388 26952
rect 13422 26918 13456 26952
rect 13490 26918 13524 26952
rect 13558 26918 13592 26952
rect 13626 26918 13660 26952
rect 13694 26918 13728 26952
rect 13762 26918 13796 26952
rect 13830 26918 13864 26952
rect 13898 26918 13932 26952
rect 13966 26918 14000 26952
rect 14034 26918 14068 26952
rect 14102 26918 14136 26952
rect 14170 26918 14204 26952
rect 14238 26918 14272 26952
rect 14306 26918 14340 26952
rect 14374 26918 14408 26952
rect 14442 26918 14476 26952
rect 14510 26918 14544 26952
rect 14578 26918 14612 26952
rect 14646 26918 14680 26952
rect 14714 26918 14748 26952
rect 14782 26918 14816 26952
rect 14850 26918 14884 26952
rect 14918 26918 14952 26952
rect 2814 26882 14952 26918
rect 2814 26848 2848 26882
rect 2882 26848 2916 26882
rect 2950 26848 2984 26882
rect 3018 26848 3052 26882
rect 3086 26848 3120 26882
rect 3154 26848 3188 26882
rect 3222 26848 3256 26882
rect 3290 26848 3324 26882
rect 3358 26848 3392 26882
rect 3426 26848 3460 26882
rect 3494 26848 3528 26882
rect 3562 26848 3596 26882
rect 3630 26848 3664 26882
rect 3698 26848 3732 26882
rect 3766 26848 3800 26882
rect 3834 26848 3868 26882
rect 3902 26848 3936 26882
rect 3970 26848 4004 26882
rect 4038 26848 4072 26882
rect 4106 26848 4140 26882
rect 4174 26848 4208 26882
rect 4242 26848 4276 26882
rect 4310 26848 4344 26882
rect 4378 26848 4412 26882
rect 4446 26848 4480 26882
rect 4514 26848 4548 26882
rect 4582 26848 4616 26882
rect 4650 26848 4684 26882
rect 4718 26848 4752 26882
rect 4786 26848 4820 26882
rect 4854 26848 4888 26882
rect 4922 26848 4956 26882
rect 4990 26848 5024 26882
rect 5058 26848 5092 26882
rect 5126 26848 5160 26882
rect 5194 26848 5228 26882
rect 5262 26848 5296 26882
rect 5330 26848 5364 26882
rect 5398 26848 5432 26882
rect 5466 26848 5500 26882
rect 5534 26848 5568 26882
rect 5602 26848 5636 26882
rect 5670 26848 5704 26882
rect 5738 26848 5772 26882
rect 5806 26848 5840 26882
rect 5874 26848 5908 26882
rect 5942 26848 5976 26882
rect 6010 26848 6044 26882
rect 6078 26848 6112 26882
rect 6146 26848 6180 26882
rect 6214 26848 6248 26882
rect 6282 26848 6316 26882
rect 6350 26848 6384 26882
rect 6418 26848 6452 26882
rect 6486 26848 6520 26882
rect 6554 26848 6588 26882
rect 6622 26848 6656 26882
rect 6690 26848 6724 26882
rect 6758 26848 6792 26882
rect 6826 26848 6860 26882
rect 6894 26848 6928 26882
rect 6962 26848 6996 26882
rect 7030 26848 7064 26882
rect 7098 26848 7132 26882
rect 7166 26848 7200 26882
rect 7234 26848 7268 26882
rect 7302 26848 7336 26882
rect 7370 26848 7404 26882
rect 7438 26848 7472 26882
rect 7506 26848 7540 26882
rect 7574 26848 7608 26882
rect 7642 26848 7676 26882
rect 7710 26848 7744 26882
rect 7778 26848 7812 26882
rect 7846 26848 7880 26882
rect 7914 26848 7948 26882
rect 7982 26848 8016 26882
rect 8050 26848 8084 26882
rect 8118 26848 8152 26882
rect 8186 26848 8220 26882
rect 8254 26848 8288 26882
rect 8322 26848 8356 26882
rect 8390 26848 8424 26882
rect 8458 26848 8492 26882
rect 8526 26848 8560 26882
rect 8594 26848 8628 26882
rect 8662 26848 8696 26882
rect 8730 26848 8764 26882
rect 8798 26848 8832 26882
rect 8866 26848 8900 26882
rect 8934 26848 8968 26882
rect 9002 26848 9036 26882
rect 9070 26848 9104 26882
rect 9138 26848 9172 26882
rect 9206 26848 9240 26882
rect 9274 26848 9308 26882
rect 9342 26848 9376 26882
rect 9410 26848 9444 26882
rect 9478 26848 9512 26882
rect 9546 26848 9580 26882
rect 9614 26848 9648 26882
rect 9682 26848 9716 26882
rect 9750 26848 9784 26882
rect 9818 26848 9852 26882
rect 9886 26848 9920 26882
rect 9954 26848 9988 26882
rect 10022 26848 10056 26882
rect 10090 26848 10124 26882
rect 10158 26848 10192 26882
rect 10226 26848 10260 26882
rect 10294 26848 10328 26882
rect 10362 26848 10396 26882
rect 10430 26848 10464 26882
rect 10498 26848 10532 26882
rect 10566 26848 10600 26882
rect 10634 26848 10668 26882
rect 10702 26848 10736 26882
rect 10770 26848 10804 26882
rect 10838 26848 10872 26882
rect 10906 26848 10940 26882
rect 10974 26848 11008 26882
rect 11042 26848 11076 26882
rect 11110 26848 11144 26882
rect 11178 26848 11212 26882
rect 11246 26848 11280 26882
rect 11314 26848 11348 26882
rect 11382 26848 11416 26882
rect 11450 26848 11484 26882
rect 11518 26848 11552 26882
rect 11586 26848 11620 26882
rect 11654 26848 11688 26882
rect 11722 26848 11756 26882
rect 11790 26848 11824 26882
rect 11858 26848 11892 26882
rect 11926 26848 11960 26882
rect 11994 26848 12028 26882
rect 12062 26848 12096 26882
rect 12130 26848 12164 26882
rect 12198 26848 12232 26882
rect 12266 26848 12300 26882
rect 12334 26848 12368 26882
rect 12402 26848 12436 26882
rect 12470 26848 12504 26882
rect 12538 26848 12572 26882
rect 12606 26848 12640 26882
rect 12674 26848 12708 26882
rect 12742 26848 12776 26882
rect 12810 26848 12844 26882
rect 12878 26848 12912 26882
rect 12946 26848 12980 26882
rect 13014 26848 13048 26882
rect 13082 26848 13116 26882
rect 13150 26848 13184 26882
rect 13218 26848 13252 26882
rect 13286 26848 13320 26882
rect 13354 26848 13388 26882
rect 13422 26848 13456 26882
rect 13490 26848 13524 26882
rect 13558 26848 13592 26882
rect 13626 26848 13660 26882
rect 13694 26848 13728 26882
rect 13762 26848 13796 26882
rect 13830 26848 13864 26882
rect 13898 26848 13932 26882
rect 13966 26848 14000 26882
rect 14034 26848 14068 26882
rect 14102 26848 14136 26882
rect 14170 26848 14204 26882
rect 14238 26848 14272 26882
rect 14306 26848 14340 26882
rect 14374 26848 14408 26882
rect 14442 26848 14476 26882
rect 14510 26848 14544 26882
rect 14578 26848 14612 26882
rect 14646 26848 14680 26882
rect 14714 26848 14748 26882
rect 14782 26848 14816 26882
rect 14850 26848 14884 26882
rect 14918 26848 14952 26882
rect 2814 26812 14952 26848
rect 2814 26794 2848 26812
rect 49 26778 2848 26794
rect 2882 26778 2916 26812
rect 2950 26778 2984 26812
rect 3018 26778 3052 26812
rect 3086 26778 3120 26812
rect 3154 26778 3188 26812
rect 3222 26778 3256 26812
rect 3290 26778 3324 26812
rect 3358 26778 3392 26812
rect 3426 26778 3460 26812
rect 3494 26778 3528 26812
rect 3562 26778 3596 26812
rect 3630 26778 3664 26812
rect 3698 26778 3732 26812
rect 3766 26778 3800 26812
rect 3834 26778 3868 26812
rect 3902 26778 3936 26812
rect 3970 26778 4004 26812
rect 4038 26778 4072 26812
rect 4106 26778 4140 26812
rect 4174 26778 4208 26812
rect 4242 26778 4276 26812
rect 4310 26778 4344 26812
rect 4378 26778 4412 26812
rect 4446 26778 4480 26812
rect 4514 26778 4548 26812
rect 4582 26778 4616 26812
rect 4650 26778 4684 26812
rect 4718 26778 4752 26812
rect 4786 26778 4820 26812
rect 4854 26778 4888 26812
rect 4922 26778 4956 26812
rect 4990 26778 5024 26812
rect 5058 26778 5092 26812
rect 5126 26778 5160 26812
rect 5194 26778 5228 26812
rect 5262 26778 5296 26812
rect 5330 26778 5364 26812
rect 5398 26778 5432 26812
rect 5466 26778 5500 26812
rect 5534 26778 5568 26812
rect 5602 26778 5636 26812
rect 5670 26778 5704 26812
rect 5738 26778 5772 26812
rect 5806 26778 5840 26812
rect 5874 26778 5908 26812
rect 5942 26778 5976 26812
rect 6010 26778 6044 26812
rect 6078 26778 6112 26812
rect 6146 26778 6180 26812
rect 6214 26778 6248 26812
rect 6282 26778 6316 26812
rect 6350 26778 6384 26812
rect 6418 26778 6452 26812
rect 6486 26778 6520 26812
rect 6554 26778 6588 26812
rect 6622 26778 6656 26812
rect 6690 26778 6724 26812
rect 6758 26778 6792 26812
rect 6826 26778 6860 26812
rect 6894 26778 6928 26812
rect 6962 26778 6996 26812
rect 7030 26778 7064 26812
rect 7098 26778 7132 26812
rect 7166 26778 7200 26812
rect 7234 26778 7268 26812
rect 7302 26778 7336 26812
rect 7370 26778 7404 26812
rect 7438 26778 7472 26812
rect 7506 26778 7540 26812
rect 7574 26778 7608 26812
rect 7642 26778 7676 26812
rect 7710 26778 7744 26812
rect 7778 26778 7812 26812
rect 7846 26778 7880 26812
rect 7914 26778 7948 26812
rect 7982 26778 8016 26812
rect 8050 26778 8084 26812
rect 8118 26778 8152 26812
rect 8186 26778 8220 26812
rect 8254 26778 8288 26812
rect 8322 26778 8356 26812
rect 8390 26778 8424 26812
rect 8458 26778 8492 26812
rect 8526 26778 8560 26812
rect 8594 26778 8628 26812
rect 8662 26778 8696 26812
rect 8730 26778 8764 26812
rect 8798 26778 8832 26812
rect 8866 26778 8900 26812
rect 8934 26778 8968 26812
rect 9002 26778 9036 26812
rect 9070 26778 9104 26812
rect 9138 26778 9172 26812
rect 9206 26778 9240 26812
rect 9274 26778 9308 26812
rect 9342 26778 9376 26812
rect 9410 26778 9444 26812
rect 9478 26778 9512 26812
rect 9546 26778 9580 26812
rect 9614 26778 9648 26812
rect 9682 26778 9716 26812
rect 9750 26778 9784 26812
rect 9818 26778 9852 26812
rect 9886 26778 9920 26812
rect 9954 26778 9988 26812
rect 10022 26778 10056 26812
rect 10090 26778 10124 26812
rect 10158 26778 10192 26812
rect 10226 26778 10260 26812
rect 10294 26778 10328 26812
rect 10362 26778 10396 26812
rect 10430 26778 10464 26812
rect 10498 26778 10532 26812
rect 10566 26778 10600 26812
rect 10634 26778 10668 26812
rect 10702 26778 10736 26812
rect 10770 26778 10804 26812
rect 10838 26778 10872 26812
rect 10906 26778 10940 26812
rect 10974 26778 11008 26812
rect 11042 26778 11076 26812
rect 11110 26778 11144 26812
rect 11178 26778 11212 26812
rect 11246 26778 11280 26812
rect 11314 26778 11348 26812
rect 11382 26778 11416 26812
rect 11450 26778 11484 26812
rect 11518 26778 11552 26812
rect 11586 26778 11620 26812
rect 11654 26778 11688 26812
rect 11722 26778 11756 26812
rect 11790 26778 11824 26812
rect 11858 26778 11892 26812
rect 11926 26778 11960 26812
rect 11994 26778 12028 26812
rect 12062 26778 12096 26812
rect 12130 26778 12164 26812
rect 12198 26778 12232 26812
rect 12266 26778 12300 26812
rect 12334 26778 12368 26812
rect 12402 26778 12436 26812
rect 12470 26778 12504 26812
rect 12538 26778 12572 26812
rect 12606 26778 12640 26812
rect 12674 26778 12708 26812
rect 12742 26778 12776 26812
rect 12810 26778 12844 26812
rect 12878 26778 12912 26812
rect 12946 26778 12980 26812
rect 13014 26778 13048 26812
rect 13082 26778 13116 26812
rect 13150 26778 13184 26812
rect 13218 26778 13252 26812
rect 13286 26778 13320 26812
rect 13354 26778 13388 26812
rect 13422 26778 13456 26812
rect 13490 26778 13524 26812
rect 13558 26778 13592 26812
rect 13626 26778 13660 26812
rect 13694 26778 13728 26812
rect 13762 26778 13796 26812
rect 13830 26778 13864 26812
rect 13898 26778 13932 26812
rect 13966 26778 14000 26812
rect 14034 26778 14068 26812
rect 14102 26778 14136 26812
rect 14170 26778 14204 26812
rect 14238 26778 14272 26812
rect 14306 26778 14340 26812
rect 14374 26778 14408 26812
rect 14442 26778 14476 26812
rect 14510 26778 14544 26812
rect 14578 26778 14612 26812
rect 14646 26778 14680 26812
rect 14714 26778 14748 26812
rect 14782 26778 14816 26812
rect 14850 26778 14884 26812
rect 14918 26778 14952 26812
rect 49 26757 14952 26778
rect 49 26723 83 26757
rect 117 26723 152 26757
rect 186 26723 221 26757
rect 255 26723 290 26757
rect 324 26723 359 26757
rect 393 26723 428 26757
rect 462 26723 497 26757
rect 531 26723 566 26757
rect 600 26723 635 26757
rect 669 26723 704 26757
rect 738 26723 773 26757
rect 807 26723 842 26757
rect 876 26723 911 26757
rect 945 26723 980 26757
rect 1014 26723 1049 26757
rect 1083 26723 1118 26757
rect 1152 26723 1187 26757
rect 1221 26723 1256 26757
rect 1290 26723 1325 26757
rect 1359 26723 1394 26757
rect 1428 26723 1463 26757
rect 1497 26723 1532 26757
rect 1566 26723 1601 26757
rect 1635 26723 1670 26757
rect 1704 26723 1739 26757
rect 1773 26723 1808 26757
rect 1842 26723 1877 26757
rect 1911 26723 1946 26757
rect 1980 26723 2014 26757
rect 2048 26723 2082 26757
rect 2116 26723 2150 26757
rect 2184 26723 2218 26757
rect 2252 26723 2286 26757
rect 2320 26723 2354 26757
rect 2388 26723 2422 26757
rect 2456 26723 2490 26757
rect 2524 26723 2558 26757
rect 2592 26723 2626 26757
rect 2660 26723 2694 26757
rect 2728 26723 2762 26757
rect 2796 26742 14952 26757
rect 2796 26723 2848 26742
rect 49 26708 2848 26723
rect 2882 26708 2916 26742
rect 2950 26708 2984 26742
rect 3018 26708 3052 26742
rect 3086 26708 3120 26742
rect 3154 26708 3188 26742
rect 3222 26708 3256 26742
rect 3290 26708 3324 26742
rect 3358 26708 3392 26742
rect 3426 26708 3460 26742
rect 3494 26708 3528 26742
rect 3562 26708 3596 26742
rect 3630 26708 3664 26742
rect 3698 26708 3732 26742
rect 3766 26708 3800 26742
rect 3834 26708 3868 26742
rect 3902 26708 3936 26742
rect 3970 26708 4004 26742
rect 4038 26708 4072 26742
rect 4106 26708 4140 26742
rect 4174 26708 4208 26742
rect 4242 26708 4276 26742
rect 4310 26708 4344 26742
rect 4378 26708 4412 26742
rect 4446 26708 4480 26742
rect 4514 26708 4548 26742
rect 4582 26708 4616 26742
rect 4650 26708 4684 26742
rect 4718 26708 4752 26742
rect 4786 26708 4820 26742
rect 4854 26708 4888 26742
rect 4922 26708 4956 26742
rect 4990 26708 5024 26742
rect 5058 26708 5092 26742
rect 5126 26708 5160 26742
rect 5194 26708 5228 26742
rect 5262 26708 5296 26742
rect 5330 26708 5364 26742
rect 5398 26708 5432 26742
rect 5466 26708 5500 26742
rect 5534 26708 5568 26742
rect 5602 26708 5636 26742
rect 5670 26708 5704 26742
rect 5738 26708 5772 26742
rect 5806 26708 5840 26742
rect 5874 26708 5908 26742
rect 5942 26708 5976 26742
rect 6010 26708 6044 26742
rect 6078 26708 6112 26742
rect 6146 26708 6180 26742
rect 6214 26708 6248 26742
rect 6282 26708 6316 26742
rect 6350 26708 6384 26742
rect 6418 26708 6452 26742
rect 6486 26708 6520 26742
rect 6554 26708 6588 26742
rect 6622 26708 6656 26742
rect 6690 26708 6724 26742
rect 6758 26708 6792 26742
rect 6826 26708 6860 26742
rect 6894 26708 6928 26742
rect 6962 26708 6996 26742
rect 7030 26708 7064 26742
rect 7098 26708 7132 26742
rect 7166 26708 7200 26742
rect 7234 26708 7268 26742
rect 7302 26708 7336 26742
rect 7370 26708 7404 26742
rect 7438 26708 7472 26742
rect 7506 26708 7540 26742
rect 7574 26708 7608 26742
rect 7642 26708 7676 26742
rect 7710 26708 7744 26742
rect 7778 26708 7812 26742
rect 7846 26708 7880 26742
rect 7914 26708 7948 26742
rect 7982 26708 8016 26742
rect 8050 26708 8084 26742
rect 8118 26708 8152 26742
rect 8186 26708 8220 26742
rect 8254 26708 8288 26742
rect 8322 26708 8356 26742
rect 8390 26708 8424 26742
rect 8458 26708 8492 26742
rect 8526 26708 8560 26742
rect 8594 26708 8628 26742
rect 8662 26708 8696 26742
rect 8730 26708 8764 26742
rect 8798 26708 8832 26742
rect 8866 26708 8900 26742
rect 8934 26708 8968 26742
rect 9002 26708 9036 26742
rect 9070 26708 9104 26742
rect 9138 26708 9172 26742
rect 9206 26708 9240 26742
rect 9274 26708 9308 26742
rect 9342 26708 9376 26742
rect 9410 26708 9444 26742
rect 9478 26708 9512 26742
rect 9546 26708 9580 26742
rect 9614 26708 9648 26742
rect 9682 26708 9716 26742
rect 9750 26708 9784 26742
rect 9818 26708 9852 26742
rect 9886 26708 9920 26742
rect 9954 26708 9988 26742
rect 10022 26708 10056 26742
rect 10090 26708 10124 26742
rect 10158 26708 10192 26742
rect 10226 26708 10260 26742
rect 10294 26708 10328 26742
rect 10362 26708 10396 26742
rect 10430 26708 10464 26742
rect 10498 26708 10532 26742
rect 10566 26708 10600 26742
rect 10634 26708 10668 26742
rect 10702 26708 10736 26742
rect 10770 26708 10804 26742
rect 10838 26708 10872 26742
rect 10906 26708 10940 26742
rect 10974 26708 11008 26742
rect 11042 26708 11076 26742
rect 11110 26708 11144 26742
rect 11178 26708 11212 26742
rect 11246 26708 11280 26742
rect 11314 26708 11348 26742
rect 11382 26708 11416 26742
rect 11450 26708 11484 26742
rect 11518 26708 11552 26742
rect 11586 26708 11620 26742
rect 11654 26708 11688 26742
rect 11722 26708 11756 26742
rect 11790 26708 11824 26742
rect 11858 26708 11892 26742
rect 11926 26708 11960 26742
rect 11994 26708 12028 26742
rect 12062 26708 12096 26742
rect 12130 26708 12164 26742
rect 12198 26708 12232 26742
rect 12266 26708 12300 26742
rect 12334 26708 12368 26742
rect 12402 26708 12436 26742
rect 12470 26708 12504 26742
rect 12538 26708 12572 26742
rect 12606 26708 12640 26742
rect 12674 26708 12708 26742
rect 12742 26708 12776 26742
rect 12810 26708 12844 26742
rect 12878 26708 12912 26742
rect 12946 26708 12980 26742
rect 13014 26708 13048 26742
rect 13082 26708 13116 26742
rect 13150 26708 13184 26742
rect 13218 26708 13252 26742
rect 13286 26708 13320 26742
rect 13354 26708 13388 26742
rect 13422 26708 13456 26742
rect 13490 26708 13524 26742
rect 13558 26708 13592 26742
rect 13626 26708 13660 26742
rect 13694 26708 13728 26742
rect 13762 26708 13796 26742
rect 13830 26708 13864 26742
rect 13898 26708 13932 26742
rect 13966 26708 14000 26742
rect 14034 26708 14068 26742
rect 14102 26708 14136 26742
rect 14170 26708 14204 26742
rect 14238 26708 14272 26742
rect 14306 26708 14340 26742
rect 14374 26708 14408 26742
rect 14442 26708 14476 26742
rect 14510 26708 14544 26742
rect 14578 26708 14612 26742
rect 14646 26708 14680 26742
rect 14714 26708 14748 26742
rect 14782 26708 14816 26742
rect 14850 26708 14884 26742
rect 14918 26708 14952 26742
rect 49 26683 14952 26708
rect 49 26649 83 26683
rect 117 26649 152 26683
rect 186 26649 221 26683
rect 255 26649 290 26683
rect 324 26649 359 26683
rect 393 26649 428 26683
rect 462 26649 497 26683
rect 531 26649 566 26683
rect 600 26649 635 26683
rect 669 26649 704 26683
rect 738 26649 773 26683
rect 807 26649 842 26683
rect 876 26649 911 26683
rect 945 26649 980 26683
rect 1014 26649 1049 26683
rect 1083 26649 1118 26683
rect 1152 26649 1187 26683
rect 1221 26649 1256 26683
rect 1290 26649 1325 26683
rect 1359 26649 1394 26683
rect 1428 26649 1463 26683
rect 1497 26649 1532 26683
rect 1566 26649 1601 26683
rect 1635 26649 1670 26683
rect 1704 26649 1739 26683
rect 1773 26649 1808 26683
rect 1842 26649 1877 26683
rect 1911 26649 1946 26683
rect 1980 26649 2014 26683
rect 2048 26649 2082 26683
rect 2116 26649 2150 26683
rect 2184 26649 2218 26683
rect 2252 26649 2286 26683
rect 2320 26649 2354 26683
rect 2388 26649 2422 26683
rect 2456 26649 2490 26683
rect 2524 26649 2558 26683
rect 2592 26649 2626 26683
rect 2660 26649 2694 26683
rect 2728 26649 2762 26683
rect 2796 26672 14952 26683
rect 2796 26649 2848 26672
rect 49 26638 2848 26649
rect 2882 26638 2916 26672
rect 2950 26638 2984 26672
rect 3018 26638 3052 26672
rect 3086 26638 3120 26672
rect 3154 26638 3188 26672
rect 3222 26638 3256 26672
rect 3290 26638 3324 26672
rect 3358 26638 3392 26672
rect 3426 26638 3460 26672
rect 3494 26638 3528 26672
rect 3562 26638 3596 26672
rect 3630 26638 3664 26672
rect 3698 26638 3732 26672
rect 3766 26638 3800 26672
rect 3834 26638 3868 26672
rect 3902 26638 3936 26672
rect 3970 26638 4004 26672
rect 4038 26638 4072 26672
rect 4106 26638 4140 26672
rect 4174 26638 4208 26672
rect 4242 26638 4276 26672
rect 4310 26638 4344 26672
rect 4378 26638 4412 26672
rect 4446 26638 4480 26672
rect 4514 26638 4548 26672
rect 4582 26638 4616 26672
rect 4650 26638 4684 26672
rect 4718 26638 4752 26672
rect 4786 26638 4820 26672
rect 4854 26638 4888 26672
rect 4922 26638 4956 26672
rect 4990 26638 5024 26672
rect 5058 26638 5092 26672
rect 5126 26638 5160 26672
rect 5194 26638 5228 26672
rect 5262 26638 5296 26672
rect 5330 26638 5364 26672
rect 5398 26638 5432 26672
rect 5466 26638 5500 26672
rect 5534 26638 5568 26672
rect 5602 26638 5636 26672
rect 5670 26638 5704 26672
rect 5738 26638 5772 26672
rect 5806 26638 5840 26672
rect 5874 26638 5908 26672
rect 5942 26638 5976 26672
rect 6010 26638 6044 26672
rect 6078 26638 6112 26672
rect 6146 26638 6180 26672
rect 6214 26638 6248 26672
rect 6282 26638 6316 26672
rect 6350 26638 6384 26672
rect 6418 26638 6452 26672
rect 6486 26638 6520 26672
rect 6554 26638 6588 26672
rect 6622 26638 6656 26672
rect 6690 26638 6724 26672
rect 6758 26638 6792 26672
rect 6826 26638 6860 26672
rect 6894 26638 6928 26672
rect 6962 26638 6996 26672
rect 7030 26638 7064 26672
rect 7098 26638 7132 26672
rect 7166 26638 7200 26672
rect 7234 26638 7268 26672
rect 7302 26638 7336 26672
rect 7370 26638 7404 26672
rect 7438 26638 7472 26672
rect 7506 26638 7540 26672
rect 7574 26638 7608 26672
rect 7642 26638 7676 26672
rect 7710 26638 7744 26672
rect 7778 26638 7812 26672
rect 7846 26638 7880 26672
rect 7914 26638 7948 26672
rect 7982 26638 8016 26672
rect 8050 26638 8084 26672
rect 8118 26638 8152 26672
rect 8186 26638 8220 26672
rect 8254 26638 8288 26672
rect 8322 26638 8356 26672
rect 8390 26638 8424 26672
rect 8458 26638 8492 26672
rect 8526 26638 8560 26672
rect 8594 26638 8628 26672
rect 8662 26638 8696 26672
rect 8730 26638 8764 26672
rect 8798 26638 8832 26672
rect 8866 26638 8900 26672
rect 8934 26638 8968 26672
rect 9002 26638 9036 26672
rect 9070 26638 9104 26672
rect 9138 26638 9172 26672
rect 9206 26638 9240 26672
rect 9274 26638 9308 26672
rect 9342 26638 9376 26672
rect 9410 26638 9444 26672
rect 9478 26638 9512 26672
rect 9546 26638 9580 26672
rect 9614 26638 9648 26672
rect 9682 26638 9716 26672
rect 9750 26638 9784 26672
rect 9818 26638 9852 26672
rect 9886 26638 9920 26672
rect 9954 26638 9988 26672
rect 10022 26638 10056 26672
rect 10090 26638 10124 26672
rect 10158 26638 10192 26672
rect 10226 26638 10260 26672
rect 10294 26638 10328 26672
rect 10362 26638 10396 26672
rect 10430 26638 10464 26672
rect 10498 26638 10532 26672
rect 10566 26638 10600 26672
rect 10634 26638 10668 26672
rect 10702 26638 10736 26672
rect 10770 26638 10804 26672
rect 10838 26638 10872 26672
rect 10906 26638 10940 26672
rect 10974 26638 11008 26672
rect 11042 26638 11076 26672
rect 11110 26638 11144 26672
rect 11178 26638 11212 26672
rect 11246 26638 11280 26672
rect 11314 26638 11348 26672
rect 11382 26638 11416 26672
rect 11450 26638 11484 26672
rect 11518 26638 11552 26672
rect 11586 26638 11620 26672
rect 11654 26638 11688 26672
rect 11722 26638 11756 26672
rect 11790 26638 11824 26672
rect 11858 26638 11892 26672
rect 11926 26638 11960 26672
rect 11994 26638 12028 26672
rect 12062 26638 12096 26672
rect 12130 26638 12164 26672
rect 12198 26638 12232 26672
rect 12266 26638 12300 26672
rect 12334 26638 12368 26672
rect 12402 26638 12436 26672
rect 12470 26638 12504 26672
rect 12538 26638 12572 26672
rect 12606 26638 12640 26672
rect 12674 26638 12708 26672
rect 12742 26638 12776 26672
rect 12810 26638 12844 26672
rect 12878 26638 12912 26672
rect 12946 26638 12980 26672
rect 13014 26638 13048 26672
rect 13082 26638 13116 26672
rect 13150 26638 13184 26672
rect 13218 26638 13252 26672
rect 13286 26638 13320 26672
rect 13354 26638 13388 26672
rect 13422 26638 13456 26672
rect 13490 26638 13524 26672
rect 13558 26638 13592 26672
rect 13626 26638 13660 26672
rect 13694 26638 13728 26672
rect 13762 26638 13796 26672
rect 13830 26638 13864 26672
rect 13898 26638 13932 26672
rect 13966 26638 14000 26672
rect 14034 26638 14068 26672
rect 14102 26638 14136 26672
rect 14170 26638 14204 26672
rect 14238 26638 14272 26672
rect 14306 26638 14340 26672
rect 14374 26638 14408 26672
rect 14442 26638 14476 26672
rect 14510 26638 14544 26672
rect 14578 26638 14612 26672
rect 14646 26638 14680 26672
rect 14714 26638 14748 26672
rect 14782 26638 14816 26672
rect 14850 26638 14884 26672
rect 14918 26638 14952 26672
rect 49 26609 14952 26638
rect 49 26575 83 26609
rect 117 26575 152 26609
rect 186 26575 221 26609
rect 255 26575 290 26609
rect 324 26575 359 26609
rect 393 26575 428 26609
rect 462 26575 497 26609
rect 531 26575 566 26609
rect 600 26575 635 26609
rect 669 26575 704 26609
rect 738 26575 773 26609
rect 807 26575 842 26609
rect 876 26575 911 26609
rect 945 26575 980 26609
rect 1014 26575 1049 26609
rect 1083 26575 1118 26609
rect 1152 26575 1187 26609
rect 1221 26575 1256 26609
rect 1290 26575 1325 26609
rect 1359 26575 1394 26609
rect 1428 26575 1463 26609
rect 1497 26575 1532 26609
rect 1566 26575 1601 26609
rect 1635 26575 1670 26609
rect 1704 26575 1739 26609
rect 1773 26575 1808 26609
rect 1842 26575 1877 26609
rect 1911 26575 1946 26609
rect 1980 26575 2014 26609
rect 2048 26575 2082 26609
rect 2116 26575 2150 26609
rect 2184 26575 2218 26609
rect 2252 26575 2286 26609
rect 2320 26575 2354 26609
rect 2388 26575 2422 26609
rect 2456 26575 2490 26609
rect 2524 26575 2558 26609
rect 2592 26575 2626 26609
rect 2660 26575 2694 26609
rect 2728 26575 2762 26609
rect 2796 26602 14952 26609
rect 2796 26575 2848 26602
rect 49 26568 2848 26575
rect 2882 26568 2916 26602
rect 2950 26568 2984 26602
rect 3018 26568 3052 26602
rect 3086 26568 3120 26602
rect 3154 26568 3188 26602
rect 3222 26568 3256 26602
rect 3290 26568 3324 26602
rect 3358 26568 3392 26602
rect 3426 26568 3460 26602
rect 3494 26568 3528 26602
rect 3562 26568 3596 26602
rect 3630 26568 3664 26602
rect 3698 26568 3732 26602
rect 3766 26568 3800 26602
rect 3834 26568 3868 26602
rect 3902 26568 3936 26602
rect 3970 26568 4004 26602
rect 4038 26568 4072 26602
rect 4106 26568 4140 26602
rect 4174 26568 4208 26602
rect 4242 26568 4276 26602
rect 4310 26568 4344 26602
rect 4378 26568 4412 26602
rect 4446 26568 4480 26602
rect 4514 26568 4548 26602
rect 4582 26568 4616 26602
rect 4650 26568 4684 26602
rect 4718 26568 4752 26602
rect 4786 26568 4820 26602
rect 4854 26568 4888 26602
rect 4922 26568 4956 26602
rect 4990 26568 5024 26602
rect 5058 26568 5092 26602
rect 5126 26568 5160 26602
rect 5194 26568 5228 26602
rect 5262 26568 5296 26602
rect 5330 26568 5364 26602
rect 5398 26568 5432 26602
rect 5466 26568 5500 26602
rect 5534 26568 5568 26602
rect 5602 26568 5636 26602
rect 5670 26568 5704 26602
rect 5738 26568 5772 26602
rect 5806 26568 5840 26602
rect 5874 26568 5908 26602
rect 5942 26568 5976 26602
rect 6010 26568 6044 26602
rect 6078 26568 6112 26602
rect 6146 26568 6180 26602
rect 6214 26568 6248 26602
rect 6282 26568 6316 26602
rect 6350 26568 6384 26602
rect 6418 26568 6452 26602
rect 6486 26568 6520 26602
rect 6554 26568 6588 26602
rect 6622 26568 6656 26602
rect 6690 26568 6724 26602
rect 6758 26568 6792 26602
rect 6826 26568 6860 26602
rect 6894 26568 6928 26602
rect 6962 26568 6996 26602
rect 7030 26568 7064 26602
rect 7098 26568 7132 26602
rect 7166 26568 7200 26602
rect 7234 26568 7268 26602
rect 7302 26568 7336 26602
rect 7370 26568 7404 26602
rect 7438 26568 7472 26602
rect 7506 26568 7540 26602
rect 7574 26568 7608 26602
rect 7642 26568 7676 26602
rect 7710 26568 7744 26602
rect 7778 26568 7812 26602
rect 7846 26568 7880 26602
rect 7914 26568 7948 26602
rect 7982 26568 8016 26602
rect 8050 26568 8084 26602
rect 8118 26568 8152 26602
rect 8186 26568 8220 26602
rect 8254 26568 8288 26602
rect 8322 26568 8356 26602
rect 8390 26568 8424 26602
rect 8458 26568 8492 26602
rect 8526 26568 8560 26602
rect 8594 26568 8628 26602
rect 8662 26568 8696 26602
rect 8730 26568 8764 26602
rect 8798 26568 8832 26602
rect 8866 26568 8900 26602
rect 8934 26568 8968 26602
rect 9002 26568 9036 26602
rect 9070 26568 9104 26602
rect 9138 26568 9172 26602
rect 9206 26568 9240 26602
rect 9274 26568 9308 26602
rect 9342 26568 9376 26602
rect 9410 26568 9444 26602
rect 9478 26568 9512 26602
rect 9546 26568 9580 26602
rect 9614 26568 9648 26602
rect 9682 26568 9716 26602
rect 9750 26568 9784 26602
rect 9818 26568 9852 26602
rect 9886 26568 9920 26602
rect 9954 26568 9988 26602
rect 10022 26568 10056 26602
rect 10090 26568 10124 26602
rect 10158 26568 10192 26602
rect 10226 26568 10260 26602
rect 10294 26568 10328 26602
rect 10362 26568 10396 26602
rect 10430 26568 10464 26602
rect 10498 26568 10532 26602
rect 10566 26568 10600 26602
rect 10634 26568 10668 26602
rect 10702 26568 10736 26602
rect 10770 26568 10804 26602
rect 10838 26568 10872 26602
rect 10906 26568 10940 26602
rect 10974 26568 11008 26602
rect 11042 26568 11076 26602
rect 11110 26568 11144 26602
rect 11178 26568 11212 26602
rect 11246 26568 11280 26602
rect 11314 26568 11348 26602
rect 11382 26568 11416 26602
rect 11450 26568 11484 26602
rect 11518 26568 11552 26602
rect 11586 26568 11620 26602
rect 11654 26568 11688 26602
rect 11722 26568 11756 26602
rect 11790 26568 11824 26602
rect 11858 26568 11892 26602
rect 11926 26568 11960 26602
rect 11994 26568 12028 26602
rect 12062 26568 12096 26602
rect 12130 26568 12164 26602
rect 12198 26568 12232 26602
rect 12266 26568 12300 26602
rect 12334 26568 12368 26602
rect 12402 26568 12436 26602
rect 12470 26568 12504 26602
rect 12538 26568 12572 26602
rect 12606 26568 12640 26602
rect 12674 26568 12708 26602
rect 12742 26568 12776 26602
rect 12810 26568 12844 26602
rect 12878 26568 12912 26602
rect 12946 26568 12980 26602
rect 13014 26568 13048 26602
rect 13082 26568 13116 26602
rect 13150 26568 13184 26602
rect 13218 26568 13252 26602
rect 13286 26568 13320 26602
rect 13354 26568 13388 26602
rect 13422 26568 13456 26602
rect 13490 26568 13524 26602
rect 13558 26568 13592 26602
rect 13626 26568 13660 26602
rect 13694 26568 13728 26602
rect 13762 26568 13796 26602
rect 13830 26568 13864 26602
rect 13898 26568 13932 26602
rect 13966 26568 14000 26602
rect 14034 26568 14068 26602
rect 14102 26568 14136 26602
rect 14170 26568 14204 26602
rect 14238 26568 14272 26602
rect 14306 26568 14340 26602
rect 14374 26568 14408 26602
rect 14442 26568 14476 26602
rect 14510 26568 14544 26602
rect 14578 26568 14612 26602
rect 14646 26568 14680 26602
rect 14714 26568 14748 26602
rect 14782 26568 14816 26602
rect 14850 26568 14884 26602
rect 14918 26568 14952 26602
rect 49 26535 14952 26568
rect 49 26501 83 26535
rect 117 26501 152 26535
rect 186 26501 221 26535
rect 255 26501 290 26535
rect 324 26501 359 26535
rect 393 26501 428 26535
rect 462 26501 497 26535
rect 531 26501 566 26535
rect 600 26501 635 26535
rect 669 26501 704 26535
rect 738 26501 773 26535
rect 807 26501 842 26535
rect 876 26501 911 26535
rect 945 26501 980 26535
rect 1014 26501 1049 26535
rect 1083 26501 1118 26535
rect 1152 26501 1187 26535
rect 1221 26501 1256 26535
rect 1290 26501 1325 26535
rect 1359 26501 1394 26535
rect 1428 26501 1463 26535
rect 1497 26501 1532 26535
rect 1566 26501 1601 26535
rect 1635 26501 1670 26535
rect 1704 26501 1739 26535
rect 1773 26501 1808 26535
rect 1842 26501 1877 26535
rect 1911 26501 1946 26535
rect 1980 26501 2014 26535
rect 2048 26501 2082 26535
rect 2116 26501 2150 26535
rect 2184 26501 2218 26535
rect 2252 26501 2286 26535
rect 2320 26501 2354 26535
rect 2388 26501 2422 26535
rect 2456 26501 2490 26535
rect 2524 26501 2558 26535
rect 2592 26501 2626 26535
rect 2660 26501 2694 26535
rect 2728 26501 2762 26535
rect 2796 26532 14952 26535
rect 2796 26501 2848 26532
rect 49 26498 2848 26501
rect 2882 26498 2916 26532
rect 2950 26498 2984 26532
rect 3018 26498 3052 26532
rect 3086 26498 3120 26532
rect 3154 26498 3188 26532
rect 3222 26498 3256 26532
rect 3290 26498 3324 26532
rect 3358 26498 3392 26532
rect 3426 26498 3460 26532
rect 3494 26498 3528 26532
rect 3562 26498 3596 26532
rect 3630 26498 3664 26532
rect 3698 26498 3732 26532
rect 3766 26498 3800 26532
rect 3834 26498 3868 26532
rect 3902 26498 3936 26532
rect 3970 26498 4004 26532
rect 4038 26498 4072 26532
rect 4106 26498 4140 26532
rect 4174 26498 4208 26532
rect 4242 26498 4276 26532
rect 4310 26498 4344 26532
rect 4378 26498 4412 26532
rect 4446 26498 4480 26532
rect 4514 26498 4548 26532
rect 4582 26498 4616 26532
rect 4650 26498 4684 26532
rect 4718 26498 4752 26532
rect 4786 26498 4820 26532
rect 4854 26498 4888 26532
rect 4922 26498 4956 26532
rect 4990 26498 5024 26532
rect 5058 26498 5092 26532
rect 5126 26498 5160 26532
rect 5194 26498 5228 26532
rect 5262 26498 5296 26532
rect 5330 26498 5364 26532
rect 5398 26498 5432 26532
rect 5466 26498 5500 26532
rect 5534 26498 5568 26532
rect 5602 26498 5636 26532
rect 5670 26498 5704 26532
rect 5738 26498 5772 26532
rect 5806 26498 5840 26532
rect 5874 26498 5908 26532
rect 5942 26498 5976 26532
rect 6010 26498 6044 26532
rect 6078 26498 6112 26532
rect 6146 26498 6180 26532
rect 6214 26498 6248 26532
rect 6282 26498 6316 26532
rect 6350 26498 6384 26532
rect 6418 26498 6452 26532
rect 6486 26498 6520 26532
rect 6554 26498 6588 26532
rect 6622 26498 6656 26532
rect 6690 26498 6724 26532
rect 6758 26498 6792 26532
rect 6826 26498 6860 26532
rect 6894 26498 6928 26532
rect 6962 26498 6996 26532
rect 7030 26498 7064 26532
rect 7098 26498 7132 26532
rect 7166 26498 7200 26532
rect 7234 26498 7268 26532
rect 7302 26498 7336 26532
rect 7370 26498 7404 26532
rect 7438 26498 7472 26532
rect 7506 26498 7540 26532
rect 7574 26498 7608 26532
rect 7642 26498 7676 26532
rect 7710 26498 7744 26532
rect 7778 26498 7812 26532
rect 7846 26498 7880 26532
rect 7914 26498 7948 26532
rect 7982 26498 8016 26532
rect 8050 26498 8084 26532
rect 8118 26498 8152 26532
rect 8186 26498 8220 26532
rect 8254 26498 8288 26532
rect 8322 26498 8356 26532
rect 8390 26498 8424 26532
rect 8458 26498 8492 26532
rect 8526 26498 8560 26532
rect 8594 26498 8628 26532
rect 8662 26498 8696 26532
rect 8730 26498 8764 26532
rect 8798 26498 8832 26532
rect 8866 26498 8900 26532
rect 8934 26498 8968 26532
rect 9002 26498 9036 26532
rect 9070 26498 9104 26532
rect 9138 26498 9172 26532
rect 9206 26498 9240 26532
rect 9274 26498 9308 26532
rect 9342 26498 9376 26532
rect 9410 26498 9444 26532
rect 9478 26498 9512 26532
rect 9546 26498 9580 26532
rect 9614 26498 9648 26532
rect 9682 26498 9716 26532
rect 9750 26498 9784 26532
rect 9818 26498 9852 26532
rect 9886 26498 9920 26532
rect 9954 26498 9988 26532
rect 10022 26498 10056 26532
rect 10090 26498 10124 26532
rect 10158 26498 10192 26532
rect 10226 26498 10260 26532
rect 10294 26498 10328 26532
rect 10362 26498 10396 26532
rect 10430 26498 10464 26532
rect 10498 26498 10532 26532
rect 10566 26498 10600 26532
rect 10634 26498 10668 26532
rect 10702 26498 10736 26532
rect 10770 26498 10804 26532
rect 10838 26498 10872 26532
rect 10906 26498 10940 26532
rect 10974 26498 11008 26532
rect 11042 26498 11076 26532
rect 11110 26498 11144 26532
rect 11178 26498 11212 26532
rect 11246 26498 11280 26532
rect 11314 26498 11348 26532
rect 11382 26498 11416 26532
rect 11450 26498 11484 26532
rect 11518 26498 11552 26532
rect 11586 26498 11620 26532
rect 11654 26498 11688 26532
rect 11722 26498 11756 26532
rect 11790 26498 11824 26532
rect 11858 26498 11892 26532
rect 11926 26498 11960 26532
rect 11994 26498 12028 26532
rect 12062 26498 12096 26532
rect 12130 26498 12164 26532
rect 12198 26498 12232 26532
rect 12266 26498 12300 26532
rect 12334 26498 12368 26532
rect 12402 26498 12436 26532
rect 12470 26498 12504 26532
rect 12538 26498 12572 26532
rect 12606 26498 12640 26532
rect 12674 26498 12708 26532
rect 12742 26498 12776 26532
rect 12810 26498 12844 26532
rect 12878 26498 12912 26532
rect 12946 26498 12980 26532
rect 13014 26498 13048 26532
rect 13082 26498 13116 26532
rect 13150 26498 13184 26532
rect 13218 26498 13252 26532
rect 13286 26498 13320 26532
rect 13354 26498 13388 26532
rect 13422 26498 13456 26532
rect 13490 26498 13524 26532
rect 13558 26498 13592 26532
rect 13626 26498 13660 26532
rect 13694 26498 13728 26532
rect 13762 26498 13796 26532
rect 13830 26498 13864 26532
rect 13898 26498 13932 26532
rect 13966 26498 14000 26532
rect 14034 26498 14068 26532
rect 14102 26498 14136 26532
rect 14170 26498 14204 26532
rect 14238 26498 14272 26532
rect 14306 26498 14340 26532
rect 14374 26498 14408 26532
rect 14442 26498 14476 26532
rect 14510 26498 14544 26532
rect 14578 26498 14612 26532
rect 14646 26498 14680 26532
rect 14714 26498 14748 26532
rect 14782 26498 14816 26532
rect 14850 26498 14884 26532
rect 14918 26498 14952 26532
rect 49 26462 14952 26498
rect 49 26461 2848 26462
rect 49 26427 83 26461
rect 117 26427 152 26461
rect 186 26427 221 26461
rect 255 26427 290 26461
rect 324 26427 359 26461
rect 393 26427 428 26461
rect 462 26427 497 26461
rect 531 26427 566 26461
rect 600 26427 635 26461
rect 669 26427 704 26461
rect 738 26427 773 26461
rect 807 26427 842 26461
rect 876 26427 911 26461
rect 945 26427 980 26461
rect 1014 26427 1049 26461
rect 1083 26427 1118 26461
rect 1152 26427 1187 26461
rect 1221 26427 1256 26461
rect 1290 26427 1325 26461
rect 1359 26427 1394 26461
rect 1428 26427 1463 26461
rect 1497 26427 1532 26461
rect 1566 26427 1601 26461
rect 1635 26427 1670 26461
rect 1704 26427 1739 26461
rect 1773 26427 1808 26461
rect 1842 26427 1877 26461
rect 1911 26427 1946 26461
rect 1980 26427 2014 26461
rect 2048 26427 2082 26461
rect 2116 26427 2150 26461
rect 2184 26427 2218 26461
rect 2252 26427 2286 26461
rect 2320 26427 2354 26461
rect 2388 26427 2422 26461
rect 2456 26427 2490 26461
rect 2524 26427 2558 26461
rect 2592 26427 2626 26461
rect 2660 26427 2694 26461
rect 2728 26427 2762 26461
rect 2796 26428 2848 26461
rect 2882 26428 2916 26462
rect 2950 26428 2984 26462
rect 3018 26428 3052 26462
rect 3086 26428 3120 26462
rect 3154 26428 3188 26462
rect 3222 26428 3256 26462
rect 3290 26428 3324 26462
rect 3358 26428 3392 26462
rect 3426 26428 3460 26462
rect 3494 26428 3528 26462
rect 3562 26428 3596 26462
rect 3630 26428 3664 26462
rect 3698 26428 3732 26462
rect 3766 26428 3800 26462
rect 3834 26428 3868 26462
rect 3902 26428 3936 26462
rect 3970 26428 4004 26462
rect 4038 26428 4072 26462
rect 4106 26428 4140 26462
rect 4174 26428 4208 26462
rect 4242 26428 4276 26462
rect 4310 26428 4344 26462
rect 4378 26428 4412 26462
rect 4446 26428 4480 26462
rect 4514 26428 4548 26462
rect 4582 26428 4616 26462
rect 4650 26428 4684 26462
rect 4718 26428 4752 26462
rect 4786 26428 4820 26462
rect 4854 26428 4888 26462
rect 4922 26428 4956 26462
rect 4990 26428 5024 26462
rect 5058 26428 5092 26462
rect 5126 26428 5160 26462
rect 5194 26428 5228 26462
rect 5262 26428 5296 26462
rect 5330 26428 5364 26462
rect 5398 26428 5432 26462
rect 5466 26428 5500 26462
rect 5534 26428 5568 26462
rect 5602 26428 5636 26462
rect 5670 26428 5704 26462
rect 5738 26428 5772 26462
rect 5806 26428 5840 26462
rect 5874 26428 5908 26462
rect 5942 26428 5976 26462
rect 6010 26428 6044 26462
rect 6078 26428 6112 26462
rect 6146 26428 6180 26462
rect 6214 26428 6248 26462
rect 6282 26428 6316 26462
rect 6350 26428 6384 26462
rect 6418 26428 6452 26462
rect 6486 26428 6520 26462
rect 6554 26428 6588 26462
rect 6622 26428 6656 26462
rect 6690 26428 6724 26462
rect 6758 26428 6792 26462
rect 6826 26428 6860 26462
rect 6894 26428 6928 26462
rect 6962 26428 6996 26462
rect 7030 26428 7064 26462
rect 7098 26428 7132 26462
rect 7166 26428 7200 26462
rect 7234 26428 7268 26462
rect 7302 26428 7336 26462
rect 7370 26428 7404 26462
rect 7438 26428 7472 26462
rect 7506 26428 7540 26462
rect 7574 26428 7608 26462
rect 7642 26428 7676 26462
rect 7710 26428 7744 26462
rect 7778 26428 7812 26462
rect 7846 26428 7880 26462
rect 7914 26428 7948 26462
rect 7982 26428 8016 26462
rect 8050 26428 8084 26462
rect 8118 26428 8152 26462
rect 8186 26428 8220 26462
rect 8254 26428 8288 26462
rect 8322 26428 8356 26462
rect 8390 26428 8424 26462
rect 8458 26428 8492 26462
rect 8526 26428 8560 26462
rect 8594 26428 8628 26462
rect 8662 26428 8696 26462
rect 8730 26428 8764 26462
rect 8798 26428 8832 26462
rect 8866 26428 8900 26462
rect 8934 26428 8968 26462
rect 9002 26428 9036 26462
rect 9070 26428 9104 26462
rect 9138 26428 9172 26462
rect 9206 26428 9240 26462
rect 9274 26428 9308 26462
rect 9342 26428 9376 26462
rect 9410 26428 9444 26462
rect 9478 26428 9512 26462
rect 9546 26428 9580 26462
rect 9614 26428 9648 26462
rect 9682 26428 9716 26462
rect 9750 26428 9784 26462
rect 9818 26428 9852 26462
rect 9886 26428 9920 26462
rect 9954 26428 9988 26462
rect 10022 26428 10056 26462
rect 10090 26428 10124 26462
rect 10158 26428 10192 26462
rect 10226 26428 10260 26462
rect 10294 26428 10328 26462
rect 10362 26428 10396 26462
rect 10430 26428 10464 26462
rect 10498 26428 10532 26462
rect 10566 26428 10600 26462
rect 10634 26428 10668 26462
rect 10702 26428 10736 26462
rect 10770 26428 10804 26462
rect 10838 26428 10872 26462
rect 10906 26428 10940 26462
rect 10974 26428 11008 26462
rect 11042 26428 11076 26462
rect 11110 26428 11144 26462
rect 11178 26428 11212 26462
rect 11246 26428 11280 26462
rect 11314 26428 11348 26462
rect 11382 26428 11416 26462
rect 11450 26428 11484 26462
rect 11518 26428 11552 26462
rect 11586 26428 11620 26462
rect 11654 26428 11688 26462
rect 11722 26428 11756 26462
rect 11790 26428 11824 26462
rect 11858 26428 11892 26462
rect 11926 26428 11960 26462
rect 11994 26428 12028 26462
rect 12062 26428 12096 26462
rect 12130 26428 12164 26462
rect 12198 26428 12232 26462
rect 12266 26428 12300 26462
rect 12334 26428 12368 26462
rect 12402 26428 12436 26462
rect 12470 26428 12504 26462
rect 12538 26428 12572 26462
rect 12606 26428 12640 26462
rect 12674 26428 12708 26462
rect 12742 26428 12776 26462
rect 12810 26428 12844 26462
rect 12878 26428 12912 26462
rect 12946 26428 12980 26462
rect 13014 26428 13048 26462
rect 13082 26428 13116 26462
rect 13150 26428 13184 26462
rect 13218 26428 13252 26462
rect 13286 26428 13320 26462
rect 13354 26428 13388 26462
rect 13422 26428 13456 26462
rect 13490 26428 13524 26462
rect 13558 26428 13592 26462
rect 13626 26428 13660 26462
rect 13694 26428 13728 26462
rect 13762 26428 13796 26462
rect 13830 26428 13864 26462
rect 13898 26428 13932 26462
rect 13966 26428 14000 26462
rect 14034 26428 14068 26462
rect 14102 26428 14136 26462
rect 14170 26428 14204 26462
rect 14238 26428 14272 26462
rect 14306 26428 14340 26462
rect 14374 26428 14408 26462
rect 14442 26428 14476 26462
rect 14510 26428 14544 26462
rect 14578 26428 14612 26462
rect 14646 26428 14680 26462
rect 14714 26428 14748 26462
rect 14782 26428 14816 26462
rect 14850 26428 14884 26462
rect 14918 26428 14952 26462
rect 2796 26427 14952 26428
rect 49 26351 14952 26427
rect 49 26317 83 26351
rect 117 26317 152 26351
rect 186 26317 221 26351
rect 255 26317 290 26351
rect 324 26317 359 26351
rect 393 26317 428 26351
rect 462 26317 497 26351
rect 531 26317 566 26351
rect 600 26317 635 26351
rect 669 26317 704 26351
rect 738 26317 773 26351
rect 807 26317 842 26351
rect 876 26317 911 26351
rect 945 26317 980 26351
rect 1014 26317 1049 26351
rect 1083 26317 1118 26351
rect 1152 26317 1187 26351
rect 1221 26317 1256 26351
rect 1290 26317 1325 26351
rect 1359 26317 1394 26351
rect 1428 26317 1463 26351
rect 1497 26317 1532 26351
rect 1566 26317 1601 26351
rect 1635 26317 1670 26351
rect 1704 26317 1739 26351
rect 1773 26317 1808 26351
rect 1842 26317 1877 26351
rect 1911 26317 1946 26351
rect 1980 26317 2015 26351
rect 2049 26317 2084 26351
rect 2118 26317 2153 26351
rect 2187 26317 2222 26351
rect 2256 26317 2291 26351
rect 2325 26317 2360 26351
rect 2394 26317 2429 26351
rect 2463 26317 2498 26351
rect 2532 26317 2567 26351
rect 2601 26317 2636 26351
rect 2670 26317 2705 26351
rect 2739 26317 2774 26351
rect 2808 26317 2843 26351
rect 2877 26317 2912 26351
rect 2946 26317 2981 26351
rect 3015 26317 3050 26351
rect 3084 26317 3119 26351
rect 3153 26317 3188 26351
rect 3222 26317 3256 26351
rect 3290 26317 3324 26351
rect 3358 26317 3392 26351
rect 3426 26317 3460 26351
rect 3494 26317 3528 26351
rect 3562 26317 3596 26351
rect 3630 26317 3664 26351
rect 3698 26317 3732 26351
rect 3766 26317 3800 26351
rect 3834 26317 3868 26351
rect 3902 26317 3936 26351
rect 3970 26317 4004 26351
rect 4038 26317 4072 26351
rect 4106 26317 4140 26351
rect 4174 26317 4208 26351
rect 4242 26317 4276 26351
rect 4310 26317 4344 26351
rect 4378 26317 4412 26351
rect 4446 26317 4480 26351
rect 4514 26317 4548 26351
rect 4582 26317 4616 26351
rect 4650 26317 4684 26351
rect 4718 26317 4752 26351
rect 4786 26317 4820 26351
rect 4854 26317 4888 26351
rect 4922 26317 4956 26351
rect 4990 26317 5024 26351
rect 5058 26317 5092 26351
rect 5126 26317 5160 26351
rect 5194 26317 5228 26351
rect 5262 26317 5296 26351
rect 5330 26317 5364 26351
rect 5398 26317 5432 26351
rect 5466 26317 5500 26351
rect 5534 26317 5568 26351
rect 5602 26317 5636 26351
rect 5670 26317 5704 26351
rect 5738 26317 5772 26351
rect 5806 26317 5840 26351
rect 5874 26317 5908 26351
rect 5942 26317 5976 26351
rect 6010 26317 6044 26351
rect 6078 26317 6112 26351
rect 6146 26317 6180 26351
rect 6214 26317 6248 26351
rect 6282 26317 6316 26351
rect 6350 26317 6384 26351
rect 6418 26317 6452 26351
rect 6486 26317 6520 26351
rect 6554 26317 6588 26351
rect 6622 26317 6656 26351
rect 6690 26317 6724 26351
rect 6758 26317 6792 26351
rect 6826 26317 6860 26351
rect 6894 26317 6928 26351
rect 6962 26317 6996 26351
rect 7030 26317 7064 26351
rect 7098 26317 7132 26351
rect 7166 26317 7200 26351
rect 7234 26317 7268 26351
rect 7302 26317 7336 26351
rect 7370 26317 7404 26351
rect 7438 26317 7472 26351
rect 7506 26317 7540 26351
rect 7574 26317 7608 26351
rect 7642 26317 7676 26351
rect 7710 26317 7744 26351
rect 7778 26317 7812 26351
rect 7846 26317 7880 26351
rect 7914 26317 7948 26351
rect 7982 26317 8016 26351
rect 8050 26317 8084 26351
rect 8118 26317 8152 26351
rect 8186 26317 8220 26351
rect 8254 26317 8288 26351
rect 8322 26317 8356 26351
rect 8390 26317 8424 26351
rect 8458 26317 8492 26351
rect 8526 26317 8560 26351
rect 8594 26317 8628 26351
rect 8662 26317 8696 26351
rect 8730 26317 8764 26351
rect 8798 26317 8832 26351
rect 8866 26317 8900 26351
rect 8934 26317 8968 26351
rect 9002 26317 9036 26351
rect 9070 26317 9104 26351
rect 9138 26317 9172 26351
rect 9206 26317 9240 26351
rect 9274 26317 9308 26351
rect 9342 26317 9376 26351
rect 9410 26317 9444 26351
rect 9478 26317 9512 26351
rect 9546 26317 9580 26351
rect 9614 26317 9648 26351
rect 9682 26317 9716 26351
rect 9750 26317 9784 26351
rect 9818 26317 9852 26351
rect 9886 26317 9920 26351
rect 9954 26317 9988 26351
rect 10022 26317 10056 26351
rect 10090 26317 10124 26351
rect 10158 26317 10192 26351
rect 10226 26317 10260 26351
rect 10294 26317 10328 26351
rect 10362 26317 10396 26351
rect 10430 26317 10464 26351
rect 10498 26317 10532 26351
rect 10566 26317 10600 26351
rect 10634 26317 10668 26351
rect 10702 26317 10736 26351
rect 10770 26317 10804 26351
rect 10838 26317 10872 26351
rect 10906 26317 10940 26351
rect 10974 26317 11008 26351
rect 11042 26317 11076 26351
rect 11110 26317 11144 26351
rect 11178 26317 11212 26351
rect 11246 26317 11280 26351
rect 11314 26317 11348 26351
rect 11382 26317 11416 26351
rect 11450 26317 11484 26351
rect 11518 26317 11552 26351
rect 11586 26317 11620 26351
rect 11654 26317 11688 26351
rect 11722 26317 11756 26351
rect 11790 26317 11824 26351
rect 11858 26317 11892 26351
rect 11926 26317 11960 26351
rect 11994 26317 12028 26351
rect 12062 26317 12096 26351
rect 12130 26317 12164 26351
rect 12198 26317 12232 26351
rect 12266 26317 12300 26351
rect 12334 26317 12368 26351
rect 12402 26317 12436 26351
rect 12470 26317 12504 26351
rect 12538 26317 12572 26351
rect 12606 26317 12640 26351
rect 12674 26317 12708 26351
rect 12742 26317 12776 26351
rect 12810 26317 12844 26351
rect 12878 26317 12912 26351
rect 12946 26317 12980 26351
rect 13014 26317 13048 26351
rect 13082 26317 13116 26351
rect 13150 26317 13184 26351
rect 13218 26317 13252 26351
rect 13286 26317 13320 26351
rect 13354 26317 13388 26351
rect 13422 26317 13456 26351
rect 13490 26317 13524 26351
rect 13558 26317 13592 26351
rect 13626 26317 13660 26351
rect 13694 26317 13728 26351
rect 13762 26317 13796 26351
rect 13830 26317 13864 26351
rect 13898 26317 13932 26351
rect 13966 26317 14000 26351
rect 14034 26317 14068 26351
rect 14102 26317 14136 26351
rect 14170 26317 14204 26351
rect 14238 26317 14272 26351
rect 14306 26317 14340 26351
rect 14374 26317 14408 26351
rect 14442 26317 14476 26351
rect 14510 26317 14544 26351
rect 14578 26317 14612 26351
rect 14646 26317 14680 26351
rect 14714 26317 14748 26351
rect 14782 26317 14816 26351
rect 14850 26317 14884 26351
rect 14918 26317 14952 26351
rect 49 26244 14952 26317
rect 49 26210 69 26244
rect 103 26210 138 26244
rect 172 26210 207 26244
rect 241 26210 276 26244
rect 310 26210 345 26244
rect 379 26210 414 26244
rect 448 26210 483 26244
rect 517 26210 552 26244
rect 586 26210 621 26244
rect 655 26210 690 26244
rect 724 26210 759 26244
rect 793 26210 828 26244
rect 862 26210 897 26244
rect 931 26210 966 26244
rect 1000 26210 1035 26244
rect 1069 26210 1104 26244
rect 1138 26210 1173 26244
rect 1207 26210 1242 26244
rect 1276 26210 1311 26244
rect 1345 26210 1380 26244
rect 1414 26210 1449 26244
rect 1483 26210 1518 26244
rect 1552 26210 1587 26244
rect 1621 26210 1656 26244
rect 1690 26210 1725 26244
rect 1759 26210 1794 26244
rect 1828 26210 1863 26244
rect 1897 26210 1932 26244
rect 1966 26210 2001 26244
rect 2035 26210 2070 26244
rect 2104 26210 2139 26244
rect 2173 26210 2208 26244
rect 2242 26210 2277 26244
rect 2311 26210 2346 26244
rect 2380 26210 2415 26244
rect 2449 26210 2484 26244
rect 2518 26210 2553 26244
rect 2587 26210 2622 26244
rect 2656 26210 2691 26244
rect 2725 26210 2760 26244
rect 2794 26210 2829 26244
rect 2863 26210 2898 26244
rect 2932 26210 2967 26244
rect 3001 26210 3036 26244
rect 3070 26210 3105 26244
rect 3139 26210 3174 26244
rect 3208 26210 3243 26244
rect 3277 26210 3312 26244
rect 3346 26210 3381 26244
rect 3415 26210 3450 26244
rect 3484 26210 3519 26244
rect 3553 26210 3588 26244
rect 3622 26210 3657 26244
rect 3691 26210 3726 26244
rect 3760 26210 3795 26244
rect 3829 26210 3864 26244
rect 3898 26210 3933 26244
rect 3967 26210 4002 26244
rect 4036 26210 4071 26244
rect 4105 26210 4140 26244
rect 4174 26210 4208 26244
rect 4242 26210 4276 26244
rect 4310 26210 4344 26244
rect 4378 26210 4412 26244
rect 4446 26210 4480 26244
rect 4514 26210 4548 26244
rect 4582 26210 4616 26244
rect 4650 26210 4684 26244
rect 4718 26210 4752 26244
rect 4786 26210 4820 26244
rect 4854 26210 4888 26244
rect 4922 26210 4956 26244
rect 4990 26210 5024 26244
rect 5058 26210 5092 26244
rect 5126 26210 5160 26244
rect 5194 26210 5228 26244
rect 5262 26210 5296 26244
rect 5330 26210 5364 26244
rect 5398 26210 5432 26244
rect 5466 26210 5500 26244
rect 5534 26210 5568 26244
rect 5602 26210 5636 26244
rect 5670 26210 5704 26244
rect 5738 26210 5772 26244
rect 5806 26210 5840 26244
rect 5874 26210 5908 26244
rect 5942 26210 5976 26244
rect 6010 26210 6044 26244
rect 6078 26210 6112 26244
rect 6146 26210 6180 26244
rect 6214 26210 6248 26244
rect 6282 26210 6316 26244
rect 6350 26210 6384 26244
rect 6418 26210 6452 26244
rect 6486 26210 6520 26244
rect 6554 26210 6588 26244
rect 6622 26210 6656 26244
rect 6690 26210 6724 26244
rect 6758 26210 6792 26244
rect 6826 26210 6860 26244
rect 6894 26210 6928 26244
rect 6962 26210 6996 26244
rect 7030 26210 7064 26244
rect 7098 26210 7132 26244
rect 7166 26210 7200 26244
rect 7234 26210 7268 26244
rect 7302 26210 7336 26244
rect 7370 26210 7404 26244
rect 7438 26210 7472 26244
rect 7506 26210 7540 26244
rect 7574 26210 7608 26244
rect 7642 26210 7676 26244
rect 7710 26210 7744 26244
rect 7778 26210 7812 26244
rect 7846 26210 7880 26244
rect 7914 26210 7948 26244
rect 7982 26210 8016 26244
rect 8050 26210 8084 26244
rect 8118 26210 8152 26244
rect 8186 26210 8220 26244
rect 8254 26210 8288 26244
rect 8322 26210 8356 26244
rect 8390 26210 8424 26244
rect 8458 26210 8492 26244
rect 8526 26210 8560 26244
rect 8594 26210 8628 26244
rect 8662 26210 8696 26244
rect 8730 26210 8764 26244
rect 8798 26210 8832 26244
rect 8866 26210 8900 26244
rect 8934 26210 8968 26244
rect 9002 26210 9036 26244
rect 9070 26210 9104 26244
rect 9138 26210 9172 26244
rect 9206 26210 9240 26244
rect 9274 26210 9308 26244
rect 9342 26210 9376 26244
rect 9410 26210 9444 26244
rect 9478 26210 9512 26244
rect 9546 26210 9580 26244
rect 9614 26210 9648 26244
rect 9682 26210 9716 26244
rect 9750 26210 9784 26244
rect 9818 26210 9852 26244
rect 9886 26210 9920 26244
rect 9954 26210 9988 26244
rect 10022 26210 10056 26244
rect 10090 26210 10124 26244
rect 10158 26210 10192 26244
rect 10226 26210 10260 26244
rect 10294 26210 10328 26244
rect 10362 26210 10396 26244
rect 10430 26210 10464 26244
rect 10498 26210 10532 26244
rect 10566 26210 10600 26244
rect 10634 26210 10668 26244
rect 10702 26210 10736 26244
rect 10770 26210 10804 26244
rect 10838 26210 10872 26244
rect 10906 26210 10940 26244
rect 10974 26210 11008 26244
rect 11042 26210 11076 26244
rect 11110 26210 11144 26244
rect 11178 26210 11212 26244
rect 11246 26210 11280 26244
rect 11314 26210 11348 26244
rect 11382 26210 11416 26244
rect 11450 26210 11484 26244
rect 11518 26210 11552 26244
rect 11586 26210 11620 26244
rect 11654 26210 11688 26244
rect 11722 26210 11756 26244
rect 11790 26210 11824 26244
rect 11858 26210 11892 26244
rect 11926 26210 11960 26244
rect 11994 26210 12028 26244
rect 12062 26210 12096 26244
rect 12130 26210 12164 26244
rect 12198 26210 12232 26244
rect 12266 26210 12300 26244
rect 12334 26210 12368 26244
rect 12402 26210 12436 26244
rect 12470 26210 12504 26244
rect 12538 26210 12572 26244
rect 12606 26210 12640 26244
rect 12674 26210 12708 26244
rect 12742 26210 12776 26244
rect 12810 26210 12844 26244
rect 12878 26210 12912 26244
rect 12946 26210 12980 26244
rect 13014 26210 13048 26244
rect 13082 26210 13116 26244
rect 13150 26210 13184 26244
rect 13218 26210 13252 26244
rect 13286 26210 13320 26244
rect 13354 26210 13388 26244
rect 13422 26210 13456 26244
rect 13490 26210 13524 26244
rect 13558 26210 13592 26244
rect 13626 26210 13660 26244
rect 13694 26210 13728 26244
rect 13762 26210 13796 26244
rect 13830 26210 13864 26244
rect 13898 26210 13932 26244
rect 13966 26210 14000 26244
rect 14034 26210 14068 26244
rect 14102 26210 14136 26244
rect 14170 26210 14204 26244
rect 14238 26210 14272 26244
rect 14306 26210 14340 26244
rect 14374 26210 14408 26244
rect 14442 26210 14476 26244
rect 14510 26210 14544 26244
rect 14578 26210 14612 26244
rect 14646 26210 14680 26244
rect 14714 26210 14748 26244
rect 14782 26210 14816 26244
rect 14850 26210 14884 26244
rect 14918 26210 14952 26244
rect 49 26172 14952 26210
rect 49 26138 69 26172
rect 103 26138 138 26172
rect 172 26138 207 26172
rect 241 26138 276 26172
rect 310 26138 345 26172
rect 379 26138 414 26172
rect 448 26138 483 26172
rect 517 26138 552 26172
rect 586 26138 621 26172
rect 655 26138 690 26172
rect 724 26138 759 26172
rect 793 26138 828 26172
rect 862 26138 897 26172
rect 931 26138 966 26172
rect 1000 26138 1035 26172
rect 1069 26138 1104 26172
rect 1138 26138 1173 26172
rect 1207 26138 1242 26172
rect 1276 26138 1311 26172
rect 1345 26138 1380 26172
rect 1414 26138 1449 26172
rect 1483 26138 1518 26172
rect 1552 26138 1587 26172
rect 1621 26138 1656 26172
rect 1690 26138 1725 26172
rect 1759 26138 1794 26172
rect 1828 26138 1863 26172
rect 1897 26138 1932 26172
rect 1966 26138 2001 26172
rect 2035 26138 2070 26172
rect 2104 26138 2139 26172
rect 2173 26138 2208 26172
rect 2242 26138 2277 26172
rect 2311 26138 2346 26172
rect 2380 26138 2415 26172
rect 2449 26138 2484 26172
rect 2518 26138 2553 26172
rect 2587 26138 2622 26172
rect 2656 26138 2691 26172
rect 2725 26138 2760 26172
rect 2794 26138 2829 26172
rect 2863 26138 2898 26172
rect 2932 26138 2967 26172
rect 3001 26138 3036 26172
rect 3070 26138 3105 26172
rect 3139 26138 3174 26172
rect 3208 26138 3243 26172
rect 3277 26138 3312 26172
rect 3346 26138 3381 26172
rect 3415 26138 3450 26172
rect 3484 26138 3519 26172
rect 3553 26138 3588 26172
rect 3622 26138 3657 26172
rect 3691 26138 3726 26172
rect 3760 26138 3795 26172
rect 3829 26138 3864 26172
rect 3898 26138 3933 26172
rect 3967 26138 4002 26172
rect 4036 26138 4071 26172
rect 4105 26138 4140 26172
rect 4174 26138 4208 26172
rect 4242 26138 4276 26172
rect 4310 26138 4344 26172
rect 4378 26138 4412 26172
rect 4446 26138 4480 26172
rect 4514 26138 4548 26172
rect 4582 26138 4616 26172
rect 4650 26138 4684 26172
rect 4718 26138 4752 26172
rect 4786 26138 4820 26172
rect 4854 26138 4888 26172
rect 4922 26138 4956 26172
rect 4990 26138 5024 26172
rect 5058 26138 5092 26172
rect 5126 26138 5160 26172
rect 5194 26138 5228 26172
rect 5262 26138 5296 26172
rect 5330 26138 5364 26172
rect 5398 26138 5432 26172
rect 5466 26138 5500 26172
rect 5534 26138 5568 26172
rect 5602 26138 5636 26172
rect 5670 26138 5704 26172
rect 5738 26138 5772 26172
rect 5806 26138 5840 26172
rect 5874 26138 5908 26172
rect 5942 26138 5976 26172
rect 6010 26138 6044 26172
rect 6078 26138 6112 26172
rect 6146 26138 6180 26172
rect 6214 26138 6248 26172
rect 6282 26138 6316 26172
rect 6350 26138 6384 26172
rect 6418 26138 6452 26172
rect 6486 26138 6520 26172
rect 6554 26138 6588 26172
rect 6622 26138 6656 26172
rect 6690 26138 6724 26172
rect 6758 26138 6792 26172
rect 6826 26138 6860 26172
rect 6894 26138 6928 26172
rect 6962 26138 6996 26172
rect 7030 26138 7064 26172
rect 7098 26138 7132 26172
rect 7166 26138 7200 26172
rect 7234 26138 7268 26172
rect 7302 26138 7336 26172
rect 7370 26138 7404 26172
rect 7438 26138 7472 26172
rect 7506 26138 7540 26172
rect 7574 26138 7608 26172
rect 7642 26138 7676 26172
rect 7710 26138 7744 26172
rect 7778 26138 7812 26172
rect 7846 26138 7880 26172
rect 7914 26138 7948 26172
rect 7982 26138 8016 26172
rect 8050 26138 8084 26172
rect 8118 26138 8152 26172
rect 8186 26138 8220 26172
rect 8254 26138 8288 26172
rect 8322 26138 8356 26172
rect 8390 26138 8424 26172
rect 8458 26138 8492 26172
rect 8526 26138 8560 26172
rect 8594 26138 8628 26172
rect 8662 26138 8696 26172
rect 8730 26138 8764 26172
rect 8798 26138 8832 26172
rect 8866 26138 8900 26172
rect 8934 26138 8968 26172
rect 9002 26138 9036 26172
rect 9070 26138 9104 26172
rect 9138 26138 9172 26172
rect 9206 26138 9240 26172
rect 9274 26138 9308 26172
rect 9342 26138 9376 26172
rect 9410 26138 9444 26172
rect 9478 26138 9512 26172
rect 9546 26138 9580 26172
rect 9614 26138 9648 26172
rect 9682 26138 9716 26172
rect 9750 26138 9784 26172
rect 9818 26138 9852 26172
rect 9886 26138 9920 26172
rect 9954 26138 9988 26172
rect 10022 26138 10056 26172
rect 10090 26138 10124 26172
rect 10158 26138 10192 26172
rect 10226 26138 10260 26172
rect 10294 26138 10328 26172
rect 10362 26138 10396 26172
rect 10430 26138 10464 26172
rect 10498 26138 10532 26172
rect 10566 26138 10600 26172
rect 10634 26138 10668 26172
rect 10702 26138 10736 26172
rect 10770 26138 10804 26172
rect 10838 26138 10872 26172
rect 10906 26138 10940 26172
rect 10974 26138 11008 26172
rect 11042 26138 11076 26172
rect 11110 26138 11144 26172
rect 11178 26138 11212 26172
rect 11246 26138 11280 26172
rect 11314 26138 11348 26172
rect 11382 26138 11416 26172
rect 11450 26138 11484 26172
rect 11518 26138 11552 26172
rect 11586 26138 11620 26172
rect 11654 26138 11688 26172
rect 11722 26138 11756 26172
rect 11790 26138 11824 26172
rect 11858 26138 11892 26172
rect 11926 26138 11960 26172
rect 11994 26138 12028 26172
rect 12062 26138 12096 26172
rect 12130 26138 12164 26172
rect 12198 26138 12232 26172
rect 12266 26138 12300 26172
rect 12334 26138 12368 26172
rect 12402 26138 12436 26172
rect 12470 26138 12504 26172
rect 12538 26138 12572 26172
rect 12606 26138 12640 26172
rect 12674 26138 12708 26172
rect 12742 26138 12776 26172
rect 12810 26138 12844 26172
rect 12878 26138 12912 26172
rect 12946 26138 12980 26172
rect 13014 26138 13048 26172
rect 13082 26138 13116 26172
rect 13150 26138 13184 26172
rect 13218 26138 13252 26172
rect 13286 26138 13320 26172
rect 13354 26138 13388 26172
rect 13422 26138 13456 26172
rect 13490 26138 13524 26172
rect 13558 26138 13592 26172
rect 13626 26138 13660 26172
rect 13694 26138 13728 26172
rect 13762 26138 13796 26172
rect 13830 26138 13864 26172
rect 13898 26138 13932 26172
rect 13966 26138 14000 26172
rect 14034 26138 14068 26172
rect 14102 26138 14136 26172
rect 14170 26138 14204 26172
rect 14238 26138 14272 26172
rect 14306 26138 14340 26172
rect 14374 26138 14408 26172
rect 14442 26138 14476 26172
rect 14510 26138 14544 26172
rect 14578 26138 14612 26172
rect 14646 26138 14680 26172
rect 14714 26138 14748 26172
rect 14782 26138 14816 26172
rect 14850 26138 14884 26172
rect 14918 26138 14952 26172
rect 49 26100 14952 26138
rect 49 26066 69 26100
rect 103 26066 138 26100
rect 172 26066 207 26100
rect 241 26066 276 26100
rect 310 26066 345 26100
rect 379 26066 414 26100
rect 448 26066 483 26100
rect 517 26066 552 26100
rect 586 26066 621 26100
rect 655 26066 690 26100
rect 724 26066 759 26100
rect 793 26066 828 26100
rect 862 26066 897 26100
rect 931 26066 966 26100
rect 1000 26066 1035 26100
rect 1069 26066 1104 26100
rect 1138 26066 1173 26100
rect 1207 26066 1242 26100
rect 1276 26066 1311 26100
rect 1345 26066 1380 26100
rect 1414 26066 1449 26100
rect 1483 26066 1518 26100
rect 1552 26066 1587 26100
rect 1621 26066 1656 26100
rect 1690 26066 1725 26100
rect 1759 26066 1794 26100
rect 1828 26066 1863 26100
rect 1897 26066 1932 26100
rect 1966 26066 2001 26100
rect 2035 26066 2070 26100
rect 2104 26066 2139 26100
rect 2173 26066 2208 26100
rect 2242 26066 2277 26100
rect 2311 26066 2346 26100
rect 2380 26066 2415 26100
rect 2449 26066 2484 26100
rect 2518 26066 2553 26100
rect 2587 26066 2622 26100
rect 2656 26066 2691 26100
rect 2725 26066 2760 26100
rect 2794 26066 2829 26100
rect 2863 26066 2898 26100
rect 2932 26066 2967 26100
rect 3001 26066 3036 26100
rect 3070 26066 3105 26100
rect 3139 26066 3174 26100
rect 3208 26066 3243 26100
rect 3277 26066 3312 26100
rect 3346 26066 3381 26100
rect 3415 26066 3450 26100
rect 3484 26066 3519 26100
rect 3553 26066 3588 26100
rect 3622 26066 3657 26100
rect 3691 26066 3726 26100
rect 3760 26066 3795 26100
rect 3829 26066 3864 26100
rect 3898 26066 3933 26100
rect 3967 26066 4002 26100
rect 4036 26066 4071 26100
rect 4105 26066 4140 26100
rect 4174 26066 4208 26100
rect 4242 26066 4276 26100
rect 4310 26066 4344 26100
rect 4378 26066 4412 26100
rect 4446 26066 4480 26100
rect 4514 26066 4548 26100
rect 4582 26066 4616 26100
rect 4650 26066 4684 26100
rect 4718 26066 4752 26100
rect 4786 26066 4820 26100
rect 4854 26066 4888 26100
rect 4922 26066 4956 26100
rect 4990 26066 5024 26100
rect 5058 26066 5092 26100
rect 5126 26066 5160 26100
rect 5194 26066 5228 26100
rect 5262 26066 5296 26100
rect 5330 26066 5364 26100
rect 5398 26066 5432 26100
rect 5466 26066 5500 26100
rect 5534 26066 5568 26100
rect 5602 26066 5636 26100
rect 5670 26066 5704 26100
rect 5738 26066 5772 26100
rect 5806 26066 5840 26100
rect 5874 26066 5908 26100
rect 5942 26066 5976 26100
rect 6010 26066 6044 26100
rect 6078 26066 6112 26100
rect 6146 26066 6180 26100
rect 6214 26066 6248 26100
rect 6282 26066 6316 26100
rect 6350 26066 6384 26100
rect 6418 26066 6452 26100
rect 6486 26066 6520 26100
rect 6554 26066 6588 26100
rect 6622 26066 6656 26100
rect 6690 26066 6724 26100
rect 6758 26066 6792 26100
rect 6826 26066 6860 26100
rect 6894 26066 6928 26100
rect 6962 26066 6996 26100
rect 7030 26066 7064 26100
rect 7098 26066 7132 26100
rect 7166 26066 7200 26100
rect 7234 26066 7268 26100
rect 7302 26066 7336 26100
rect 7370 26066 7404 26100
rect 7438 26066 7472 26100
rect 7506 26066 7540 26100
rect 7574 26066 7608 26100
rect 7642 26066 7676 26100
rect 7710 26066 7744 26100
rect 7778 26066 7812 26100
rect 7846 26066 7880 26100
rect 7914 26066 7948 26100
rect 7982 26066 8016 26100
rect 8050 26066 8084 26100
rect 8118 26066 8152 26100
rect 8186 26066 8220 26100
rect 8254 26066 8288 26100
rect 8322 26066 8356 26100
rect 8390 26066 8424 26100
rect 8458 26066 8492 26100
rect 8526 26066 8560 26100
rect 8594 26066 8628 26100
rect 8662 26066 8696 26100
rect 8730 26066 8764 26100
rect 8798 26066 8832 26100
rect 8866 26066 8900 26100
rect 8934 26066 8968 26100
rect 9002 26066 9036 26100
rect 9070 26066 9104 26100
rect 9138 26066 9172 26100
rect 9206 26066 9240 26100
rect 9274 26066 9308 26100
rect 9342 26066 9376 26100
rect 9410 26066 9444 26100
rect 9478 26066 9512 26100
rect 9546 26066 9580 26100
rect 9614 26066 9648 26100
rect 9682 26066 9716 26100
rect 9750 26066 9784 26100
rect 9818 26066 9852 26100
rect 9886 26066 9920 26100
rect 9954 26066 9988 26100
rect 10022 26066 10056 26100
rect 10090 26066 10124 26100
rect 10158 26066 10192 26100
rect 10226 26066 10260 26100
rect 10294 26066 10328 26100
rect 10362 26066 10396 26100
rect 10430 26066 10464 26100
rect 10498 26066 10532 26100
rect 10566 26066 10600 26100
rect 10634 26066 10668 26100
rect 10702 26066 10736 26100
rect 10770 26066 10804 26100
rect 10838 26066 10872 26100
rect 10906 26066 10940 26100
rect 10974 26066 11008 26100
rect 11042 26066 11076 26100
rect 11110 26066 11144 26100
rect 11178 26066 11212 26100
rect 11246 26066 11280 26100
rect 11314 26066 11348 26100
rect 11382 26066 11416 26100
rect 11450 26066 11484 26100
rect 11518 26066 11552 26100
rect 11586 26066 11620 26100
rect 11654 26066 11688 26100
rect 11722 26066 11756 26100
rect 11790 26066 11824 26100
rect 11858 26066 11892 26100
rect 11926 26066 11960 26100
rect 11994 26066 12028 26100
rect 12062 26066 12096 26100
rect 12130 26066 12164 26100
rect 12198 26066 12232 26100
rect 12266 26066 12300 26100
rect 12334 26066 12368 26100
rect 12402 26066 12436 26100
rect 12470 26066 12504 26100
rect 12538 26066 12572 26100
rect 12606 26066 12640 26100
rect 12674 26066 12708 26100
rect 12742 26066 12776 26100
rect 12810 26066 12844 26100
rect 12878 26066 12912 26100
rect 12946 26066 12980 26100
rect 13014 26066 13048 26100
rect 13082 26066 13116 26100
rect 13150 26066 13184 26100
rect 13218 26066 13252 26100
rect 13286 26066 13320 26100
rect 13354 26066 13388 26100
rect 13422 26066 13456 26100
rect 13490 26066 13524 26100
rect 13558 26066 13592 26100
rect 13626 26066 13660 26100
rect 13694 26066 13728 26100
rect 13762 26066 13796 26100
rect 13830 26066 13864 26100
rect 13898 26066 13932 26100
rect 13966 26066 14000 26100
rect 14034 26066 14068 26100
rect 14102 26066 14136 26100
rect 14170 26066 14204 26100
rect 14238 26066 14272 26100
rect 14306 26066 14340 26100
rect 14374 26066 14408 26100
rect 14442 26066 14476 26100
rect 14510 26066 14544 26100
rect 14578 26066 14612 26100
rect 14646 26066 14680 26100
rect 14714 26066 14748 26100
rect 14782 26066 14816 26100
rect 14850 26066 14884 26100
rect 14918 26066 14952 26100
rect 49 26028 14952 26066
rect 49 25994 69 26028
rect 103 25994 138 26028
rect 172 25994 207 26028
rect 241 25994 276 26028
rect 310 25994 345 26028
rect 379 25994 414 26028
rect 448 25994 483 26028
rect 517 25994 552 26028
rect 586 25994 621 26028
rect 655 25994 690 26028
rect 724 25994 759 26028
rect 793 25994 828 26028
rect 862 25994 897 26028
rect 931 25994 966 26028
rect 1000 25994 1035 26028
rect 1069 25994 1104 26028
rect 1138 25994 1173 26028
rect 1207 25994 1242 26028
rect 1276 25994 1311 26028
rect 1345 25994 1380 26028
rect 1414 25994 1449 26028
rect 1483 25994 1518 26028
rect 1552 25994 1587 26028
rect 1621 25994 1656 26028
rect 1690 25994 1725 26028
rect 1759 25994 1794 26028
rect 1828 25994 1863 26028
rect 1897 25994 1932 26028
rect 1966 25994 2001 26028
rect 2035 25994 2070 26028
rect 2104 25994 2139 26028
rect 2173 25994 2208 26028
rect 2242 25994 2277 26028
rect 2311 25994 2346 26028
rect 2380 25994 2415 26028
rect 2449 25994 2484 26028
rect 2518 25994 2553 26028
rect 2587 25994 2622 26028
rect 2656 25994 2691 26028
rect 2725 25994 2760 26028
rect 2794 25994 2829 26028
rect 2863 25994 2898 26028
rect 2932 25994 2967 26028
rect 3001 25994 3036 26028
rect 3070 25994 3105 26028
rect 3139 25994 3174 26028
rect 3208 25994 3243 26028
rect 3277 25994 3312 26028
rect 3346 25994 3381 26028
rect 3415 25994 3450 26028
rect 3484 25994 3519 26028
rect 3553 25994 3588 26028
rect 3622 25994 3657 26028
rect 3691 25994 3726 26028
rect 3760 25994 3795 26028
rect 3829 25994 3864 26028
rect 3898 25994 3933 26028
rect 3967 25994 4002 26028
rect 4036 25994 4071 26028
rect 4105 25994 4140 26028
rect 4174 25994 4208 26028
rect 4242 25994 4276 26028
rect 4310 25994 4344 26028
rect 4378 25994 4412 26028
rect 4446 25994 4480 26028
rect 4514 25994 4548 26028
rect 4582 25994 4616 26028
rect 4650 25994 4684 26028
rect 4718 25994 4752 26028
rect 4786 25994 4820 26028
rect 4854 25994 4888 26028
rect 4922 25994 4956 26028
rect 4990 25994 5024 26028
rect 5058 25994 5092 26028
rect 5126 25994 5160 26028
rect 5194 25994 5228 26028
rect 5262 25994 5296 26028
rect 5330 25994 5364 26028
rect 5398 25994 5432 26028
rect 5466 25994 5500 26028
rect 5534 25994 5568 26028
rect 5602 25994 5636 26028
rect 5670 25994 5704 26028
rect 5738 25994 5772 26028
rect 5806 25994 5840 26028
rect 5874 25994 5908 26028
rect 5942 25994 5976 26028
rect 6010 25994 6044 26028
rect 6078 25994 6112 26028
rect 6146 25994 6180 26028
rect 6214 25994 6248 26028
rect 6282 25994 6316 26028
rect 6350 25994 6384 26028
rect 6418 25994 6452 26028
rect 6486 25994 6520 26028
rect 6554 25994 6588 26028
rect 6622 25994 6656 26028
rect 6690 25994 6724 26028
rect 6758 25994 6792 26028
rect 6826 25994 6860 26028
rect 6894 25994 6928 26028
rect 6962 25994 6996 26028
rect 7030 25994 7064 26028
rect 7098 25994 7132 26028
rect 7166 25994 7200 26028
rect 7234 25994 7268 26028
rect 7302 25994 7336 26028
rect 7370 25994 7404 26028
rect 7438 25994 7472 26028
rect 7506 25994 7540 26028
rect 7574 25994 7608 26028
rect 7642 25994 7676 26028
rect 7710 25994 7744 26028
rect 7778 25994 7812 26028
rect 7846 25994 7880 26028
rect 7914 25994 7948 26028
rect 7982 25994 8016 26028
rect 8050 25994 8084 26028
rect 8118 25994 8152 26028
rect 8186 25994 8220 26028
rect 8254 25994 8288 26028
rect 8322 25994 8356 26028
rect 8390 25994 8424 26028
rect 8458 25994 8492 26028
rect 8526 25994 8560 26028
rect 8594 25994 8628 26028
rect 8662 25994 8696 26028
rect 8730 25994 8764 26028
rect 8798 25994 8832 26028
rect 8866 25994 8900 26028
rect 8934 25994 8968 26028
rect 9002 25994 9036 26028
rect 9070 25994 9104 26028
rect 9138 25994 9172 26028
rect 9206 25994 9240 26028
rect 9274 25994 9308 26028
rect 9342 25994 9376 26028
rect 9410 25994 9444 26028
rect 9478 25994 9512 26028
rect 9546 25994 9580 26028
rect 9614 25994 9648 26028
rect 9682 25994 9716 26028
rect 9750 25994 9784 26028
rect 9818 25994 9852 26028
rect 9886 25994 9920 26028
rect 9954 25994 9988 26028
rect 10022 25994 10056 26028
rect 10090 25994 10124 26028
rect 10158 25994 10192 26028
rect 10226 25994 10260 26028
rect 10294 25994 10328 26028
rect 10362 25994 10396 26028
rect 10430 25994 10464 26028
rect 10498 25994 10532 26028
rect 10566 25994 10600 26028
rect 10634 25994 10668 26028
rect 10702 25994 10736 26028
rect 10770 25994 10804 26028
rect 10838 25994 10872 26028
rect 10906 25994 10940 26028
rect 10974 25994 11008 26028
rect 11042 25994 11076 26028
rect 11110 25994 11144 26028
rect 11178 25994 11212 26028
rect 11246 25994 11280 26028
rect 11314 25994 11348 26028
rect 11382 25994 11416 26028
rect 11450 25994 11484 26028
rect 11518 25994 11552 26028
rect 11586 25994 11620 26028
rect 11654 25994 11688 26028
rect 11722 25994 11756 26028
rect 11790 25994 11824 26028
rect 11858 25994 11892 26028
rect 11926 25994 11960 26028
rect 11994 25994 12028 26028
rect 12062 25994 12096 26028
rect 12130 25994 12164 26028
rect 12198 25994 12232 26028
rect 12266 25994 12300 26028
rect 12334 25994 12368 26028
rect 12402 25994 12436 26028
rect 12470 25994 12504 26028
rect 12538 25994 12572 26028
rect 12606 25994 12640 26028
rect 12674 25994 12708 26028
rect 12742 25994 12776 26028
rect 12810 25994 12844 26028
rect 12878 25994 12912 26028
rect 12946 25994 12980 26028
rect 13014 25994 13048 26028
rect 13082 25994 13116 26028
rect 13150 25994 13184 26028
rect 13218 25994 13252 26028
rect 13286 25994 13320 26028
rect 13354 25994 13388 26028
rect 13422 25994 13456 26028
rect 13490 25994 13524 26028
rect 13558 25994 13592 26028
rect 13626 25994 13660 26028
rect 13694 25994 13728 26028
rect 13762 25994 13796 26028
rect 13830 25994 13864 26028
rect 13898 25994 13932 26028
rect 13966 25994 14000 26028
rect 14034 25994 14068 26028
rect 14102 25994 14136 26028
rect 14170 25994 14204 26028
rect 14238 25994 14272 26028
rect 14306 25994 14340 26028
rect 14374 25994 14408 26028
rect 14442 25994 14476 26028
rect 14510 25994 14544 26028
rect 14578 25994 14612 26028
rect 14646 25994 14680 26028
rect 14714 25994 14748 26028
rect 14782 25994 14816 26028
rect 14850 25994 14884 26028
rect 14918 25994 14952 26028
rect 49 25956 14952 25994
rect 49 25922 69 25956
rect 103 25922 138 25956
rect 172 25922 207 25956
rect 241 25922 276 25956
rect 310 25922 345 25956
rect 379 25922 414 25956
rect 448 25922 483 25956
rect 517 25922 552 25956
rect 586 25922 621 25956
rect 655 25922 690 25956
rect 724 25922 759 25956
rect 793 25922 828 25956
rect 862 25922 897 25956
rect 931 25922 966 25956
rect 1000 25922 1035 25956
rect 1069 25922 1104 25956
rect 1138 25922 1173 25956
rect 1207 25922 1242 25956
rect 1276 25922 1311 25956
rect 1345 25922 1380 25956
rect 1414 25922 1449 25956
rect 1483 25922 1518 25956
rect 1552 25922 1587 25956
rect 1621 25922 1656 25956
rect 1690 25922 1725 25956
rect 1759 25922 1794 25956
rect 1828 25922 1863 25956
rect 1897 25922 1932 25956
rect 1966 25922 2001 25956
rect 2035 25922 2070 25956
rect 2104 25922 2139 25956
rect 2173 25922 2208 25956
rect 2242 25922 2277 25956
rect 2311 25922 2346 25956
rect 2380 25922 2415 25956
rect 2449 25922 2484 25956
rect 2518 25922 2553 25956
rect 2587 25922 2622 25956
rect 2656 25922 2691 25956
rect 2725 25922 2760 25956
rect 2794 25922 2829 25956
rect 2863 25922 2898 25956
rect 2932 25922 2967 25956
rect 3001 25922 3036 25956
rect 3070 25922 3105 25956
rect 3139 25922 3174 25956
rect 3208 25922 3243 25956
rect 3277 25922 3312 25956
rect 3346 25922 3381 25956
rect 3415 25922 3450 25956
rect 3484 25922 3519 25956
rect 3553 25922 3588 25956
rect 3622 25922 3657 25956
rect 3691 25922 3726 25956
rect 3760 25922 3795 25956
rect 3829 25922 3864 25956
rect 3898 25922 3933 25956
rect 3967 25922 4002 25956
rect 4036 25922 4071 25956
rect 4105 25922 4140 25956
rect 4174 25922 4208 25956
rect 4242 25922 4276 25956
rect 4310 25922 4344 25956
rect 4378 25922 4412 25956
rect 4446 25922 4480 25956
rect 4514 25922 4548 25956
rect 4582 25922 4616 25956
rect 4650 25922 4684 25956
rect 4718 25922 4752 25956
rect 4786 25922 4820 25956
rect 4854 25922 4888 25956
rect 4922 25922 4956 25956
rect 4990 25922 5024 25956
rect 5058 25922 5092 25956
rect 5126 25922 5160 25956
rect 5194 25922 5228 25956
rect 5262 25922 5296 25956
rect 5330 25922 5364 25956
rect 5398 25922 5432 25956
rect 5466 25922 5500 25956
rect 5534 25922 5568 25956
rect 5602 25922 5636 25956
rect 5670 25922 5704 25956
rect 5738 25922 5772 25956
rect 5806 25922 5840 25956
rect 5874 25922 5908 25956
rect 5942 25922 5976 25956
rect 6010 25922 6044 25956
rect 6078 25922 6112 25956
rect 6146 25922 6180 25956
rect 6214 25922 6248 25956
rect 6282 25922 6316 25956
rect 6350 25922 6384 25956
rect 6418 25922 6452 25956
rect 6486 25922 6520 25956
rect 6554 25922 6588 25956
rect 6622 25922 6656 25956
rect 6690 25922 6724 25956
rect 6758 25922 6792 25956
rect 6826 25922 6860 25956
rect 6894 25922 6928 25956
rect 6962 25922 6996 25956
rect 7030 25922 7064 25956
rect 7098 25922 7132 25956
rect 7166 25922 7200 25956
rect 7234 25922 7268 25956
rect 7302 25922 7336 25956
rect 7370 25922 7404 25956
rect 7438 25922 7472 25956
rect 7506 25922 7540 25956
rect 7574 25922 7608 25956
rect 7642 25922 7676 25956
rect 7710 25922 7744 25956
rect 7778 25922 7812 25956
rect 7846 25922 7880 25956
rect 7914 25922 7948 25956
rect 7982 25922 8016 25956
rect 8050 25922 8084 25956
rect 8118 25922 8152 25956
rect 8186 25922 8220 25956
rect 8254 25922 8288 25956
rect 8322 25922 8356 25956
rect 8390 25922 8424 25956
rect 8458 25922 8492 25956
rect 8526 25922 8560 25956
rect 8594 25922 8628 25956
rect 8662 25922 8696 25956
rect 8730 25922 8764 25956
rect 8798 25922 8832 25956
rect 8866 25922 8900 25956
rect 8934 25922 8968 25956
rect 9002 25922 9036 25956
rect 9070 25922 9104 25956
rect 9138 25922 9172 25956
rect 9206 25922 9240 25956
rect 9274 25922 9308 25956
rect 9342 25922 9376 25956
rect 9410 25922 9444 25956
rect 9478 25922 9512 25956
rect 9546 25922 9580 25956
rect 9614 25922 9648 25956
rect 9682 25922 9716 25956
rect 9750 25922 9784 25956
rect 9818 25922 9852 25956
rect 9886 25922 9920 25956
rect 9954 25922 9988 25956
rect 10022 25922 10056 25956
rect 10090 25922 10124 25956
rect 10158 25922 10192 25956
rect 10226 25922 10260 25956
rect 10294 25922 10328 25956
rect 10362 25922 10396 25956
rect 10430 25922 10464 25956
rect 10498 25922 10532 25956
rect 10566 25922 10600 25956
rect 10634 25922 10668 25956
rect 10702 25922 10736 25956
rect 10770 25922 10804 25956
rect 10838 25922 10872 25956
rect 10906 25922 10940 25956
rect 10974 25922 11008 25956
rect 11042 25922 11076 25956
rect 11110 25922 11144 25956
rect 11178 25922 11212 25956
rect 11246 25922 11280 25956
rect 11314 25922 11348 25956
rect 11382 25922 11416 25956
rect 11450 25922 11484 25956
rect 11518 25922 11552 25956
rect 11586 25922 11620 25956
rect 11654 25922 11688 25956
rect 11722 25922 11756 25956
rect 11790 25922 11824 25956
rect 11858 25922 11892 25956
rect 11926 25922 11960 25956
rect 11994 25922 12028 25956
rect 12062 25922 12096 25956
rect 12130 25922 12164 25956
rect 12198 25922 12232 25956
rect 12266 25922 12300 25956
rect 12334 25922 12368 25956
rect 12402 25922 12436 25956
rect 12470 25922 12504 25956
rect 12538 25922 12572 25956
rect 12606 25922 12640 25956
rect 12674 25922 12708 25956
rect 12742 25922 12776 25956
rect 12810 25922 12844 25956
rect 12878 25922 12912 25956
rect 12946 25922 12980 25956
rect 13014 25922 13048 25956
rect 13082 25922 13116 25956
rect 13150 25922 13184 25956
rect 13218 25922 13252 25956
rect 13286 25922 13320 25956
rect 13354 25922 13388 25956
rect 13422 25922 13456 25956
rect 13490 25922 13524 25956
rect 13558 25922 13592 25956
rect 13626 25922 13660 25956
rect 13694 25922 13728 25956
rect 13762 25922 13796 25956
rect 13830 25922 13864 25956
rect 13898 25922 13932 25956
rect 13966 25922 14000 25956
rect 14034 25922 14068 25956
rect 14102 25922 14136 25956
rect 14170 25922 14204 25956
rect 14238 25922 14272 25956
rect 14306 25922 14340 25956
rect 14374 25922 14408 25956
rect 14442 25922 14476 25956
rect 14510 25922 14544 25956
rect 14578 25922 14612 25956
rect 14646 25922 14680 25956
rect 14714 25922 14748 25956
rect 14782 25922 14816 25956
rect 14850 25922 14884 25956
rect 14918 25922 14952 25956
rect 49 25884 14952 25922
rect 49 25850 69 25884
rect 103 25850 138 25884
rect 172 25850 207 25884
rect 241 25850 276 25884
rect 310 25850 345 25884
rect 379 25850 414 25884
rect 448 25850 483 25884
rect 517 25850 552 25884
rect 586 25850 621 25884
rect 655 25850 690 25884
rect 724 25850 759 25884
rect 793 25850 828 25884
rect 862 25850 897 25884
rect 931 25850 966 25884
rect 1000 25850 1035 25884
rect 1069 25850 1104 25884
rect 1138 25850 1173 25884
rect 1207 25850 1242 25884
rect 1276 25850 1311 25884
rect 1345 25850 1380 25884
rect 1414 25850 1449 25884
rect 1483 25850 1518 25884
rect 1552 25850 1587 25884
rect 1621 25850 1656 25884
rect 1690 25850 1725 25884
rect 1759 25850 1794 25884
rect 1828 25850 1863 25884
rect 1897 25850 1932 25884
rect 1966 25850 2001 25884
rect 2035 25850 2070 25884
rect 2104 25850 2139 25884
rect 2173 25850 2208 25884
rect 2242 25850 2277 25884
rect 2311 25850 2346 25884
rect 2380 25850 2415 25884
rect 2449 25850 2484 25884
rect 2518 25850 2553 25884
rect 2587 25850 2622 25884
rect 2656 25850 2691 25884
rect 2725 25850 2760 25884
rect 2794 25850 2829 25884
rect 2863 25850 2898 25884
rect 2932 25850 2967 25884
rect 3001 25850 3036 25884
rect 3070 25850 3105 25884
rect 3139 25850 3174 25884
rect 3208 25850 3243 25884
rect 3277 25850 3312 25884
rect 3346 25850 3381 25884
rect 3415 25850 3450 25884
rect 3484 25850 3519 25884
rect 3553 25850 3588 25884
rect 3622 25850 3657 25884
rect 3691 25850 3726 25884
rect 3760 25850 3795 25884
rect 3829 25850 3864 25884
rect 3898 25850 3933 25884
rect 3967 25850 4002 25884
rect 4036 25850 4071 25884
rect 4105 25850 4140 25884
rect 4174 25850 4208 25884
rect 4242 25850 4276 25884
rect 4310 25850 4344 25884
rect 4378 25850 4412 25884
rect 4446 25850 4480 25884
rect 4514 25850 4548 25884
rect 4582 25850 4616 25884
rect 4650 25850 4684 25884
rect 4718 25850 4752 25884
rect 4786 25850 4820 25884
rect 4854 25850 4888 25884
rect 4922 25850 4956 25884
rect 4990 25850 5024 25884
rect 5058 25850 5092 25884
rect 5126 25850 5160 25884
rect 5194 25850 5228 25884
rect 5262 25850 5296 25884
rect 5330 25850 5364 25884
rect 5398 25850 5432 25884
rect 5466 25850 5500 25884
rect 5534 25850 5568 25884
rect 5602 25850 5636 25884
rect 5670 25850 5704 25884
rect 5738 25850 5772 25884
rect 5806 25850 5840 25884
rect 5874 25850 5908 25884
rect 5942 25850 5976 25884
rect 6010 25850 6044 25884
rect 6078 25850 6112 25884
rect 6146 25850 6180 25884
rect 6214 25850 6248 25884
rect 6282 25850 6316 25884
rect 6350 25850 6384 25884
rect 6418 25850 6452 25884
rect 6486 25850 6520 25884
rect 6554 25850 6588 25884
rect 6622 25850 6656 25884
rect 6690 25850 6724 25884
rect 6758 25850 6792 25884
rect 6826 25850 6860 25884
rect 6894 25850 6928 25884
rect 6962 25850 6996 25884
rect 7030 25850 7064 25884
rect 7098 25850 7132 25884
rect 7166 25850 7200 25884
rect 7234 25850 7268 25884
rect 7302 25850 7336 25884
rect 7370 25850 7404 25884
rect 7438 25850 7472 25884
rect 7506 25850 7540 25884
rect 7574 25850 7608 25884
rect 7642 25850 7676 25884
rect 7710 25850 7744 25884
rect 7778 25850 7812 25884
rect 7846 25850 7880 25884
rect 7914 25850 7948 25884
rect 7982 25850 8016 25884
rect 8050 25850 8084 25884
rect 8118 25850 8152 25884
rect 8186 25850 8220 25884
rect 8254 25850 8288 25884
rect 8322 25850 8356 25884
rect 8390 25850 8424 25884
rect 8458 25850 8492 25884
rect 8526 25850 8560 25884
rect 8594 25850 8628 25884
rect 8662 25850 8696 25884
rect 8730 25850 8764 25884
rect 8798 25850 8832 25884
rect 8866 25850 8900 25884
rect 8934 25850 8968 25884
rect 9002 25850 9036 25884
rect 9070 25850 9104 25884
rect 9138 25850 9172 25884
rect 9206 25850 9240 25884
rect 9274 25850 9308 25884
rect 9342 25850 9376 25884
rect 9410 25850 9444 25884
rect 9478 25850 9512 25884
rect 9546 25850 9580 25884
rect 9614 25850 9648 25884
rect 9682 25850 9716 25884
rect 9750 25850 9784 25884
rect 9818 25850 9852 25884
rect 9886 25850 9920 25884
rect 9954 25850 9988 25884
rect 10022 25850 10056 25884
rect 10090 25850 10124 25884
rect 10158 25850 10192 25884
rect 10226 25850 10260 25884
rect 10294 25850 10328 25884
rect 10362 25850 10396 25884
rect 10430 25850 10464 25884
rect 10498 25850 10532 25884
rect 10566 25850 10600 25884
rect 10634 25850 10668 25884
rect 10702 25850 10736 25884
rect 10770 25850 10804 25884
rect 10838 25850 10872 25884
rect 10906 25850 10940 25884
rect 10974 25850 11008 25884
rect 11042 25850 11076 25884
rect 11110 25850 11144 25884
rect 11178 25850 11212 25884
rect 11246 25850 11280 25884
rect 11314 25850 11348 25884
rect 11382 25850 11416 25884
rect 11450 25850 11484 25884
rect 11518 25850 11552 25884
rect 11586 25850 11620 25884
rect 11654 25850 11688 25884
rect 11722 25850 11756 25884
rect 11790 25850 11824 25884
rect 11858 25850 11892 25884
rect 11926 25850 11960 25884
rect 11994 25850 12028 25884
rect 12062 25850 12096 25884
rect 12130 25850 12164 25884
rect 12198 25850 12232 25884
rect 12266 25850 12300 25884
rect 12334 25850 12368 25884
rect 12402 25850 12436 25884
rect 12470 25850 12504 25884
rect 12538 25850 12572 25884
rect 12606 25850 12640 25884
rect 12674 25850 12708 25884
rect 12742 25850 12776 25884
rect 12810 25850 12844 25884
rect 12878 25850 12912 25884
rect 12946 25850 12980 25884
rect 13014 25850 13048 25884
rect 13082 25850 13116 25884
rect 13150 25850 13184 25884
rect 13218 25850 13252 25884
rect 13286 25850 13320 25884
rect 13354 25850 13388 25884
rect 13422 25850 13456 25884
rect 13490 25850 13524 25884
rect 13558 25850 13592 25884
rect 13626 25850 13660 25884
rect 13694 25850 13728 25884
rect 13762 25850 13796 25884
rect 13830 25850 13864 25884
rect 13898 25850 13932 25884
rect 13966 25850 14000 25884
rect 14034 25850 14068 25884
rect 14102 25850 14136 25884
rect 14170 25850 14204 25884
rect 14238 25850 14272 25884
rect 14306 25850 14340 25884
rect 14374 25850 14408 25884
rect 14442 25850 14476 25884
rect 14510 25850 14544 25884
rect 14578 25850 14612 25884
rect 14646 25850 14680 25884
rect 14714 25850 14748 25884
rect 14782 25850 14816 25884
rect 14850 25850 14884 25884
rect 14918 25850 14952 25884
rect 49 25812 14952 25850
rect 49 25778 69 25812
rect 103 25778 138 25812
rect 172 25778 207 25812
rect 241 25778 276 25812
rect 310 25778 345 25812
rect 379 25778 414 25812
rect 448 25778 483 25812
rect 517 25778 552 25812
rect 586 25778 621 25812
rect 655 25778 690 25812
rect 724 25778 759 25812
rect 793 25778 828 25812
rect 862 25778 897 25812
rect 931 25778 966 25812
rect 1000 25778 1035 25812
rect 1069 25778 1104 25812
rect 1138 25778 1173 25812
rect 1207 25778 1242 25812
rect 1276 25778 1311 25812
rect 1345 25778 1380 25812
rect 1414 25778 1449 25812
rect 1483 25778 1518 25812
rect 1552 25778 1587 25812
rect 1621 25778 1656 25812
rect 1690 25778 1725 25812
rect 1759 25778 1794 25812
rect 1828 25778 1863 25812
rect 1897 25778 1932 25812
rect 1966 25778 2001 25812
rect 2035 25778 2070 25812
rect 2104 25778 2139 25812
rect 2173 25778 2208 25812
rect 2242 25778 2277 25812
rect 2311 25778 2346 25812
rect 2380 25778 2415 25812
rect 2449 25778 2484 25812
rect 2518 25778 2553 25812
rect 2587 25778 2622 25812
rect 2656 25778 2691 25812
rect 2725 25778 2760 25812
rect 2794 25778 2829 25812
rect 2863 25778 2898 25812
rect 2932 25778 2967 25812
rect 3001 25778 3036 25812
rect 3070 25778 3105 25812
rect 3139 25778 3174 25812
rect 3208 25778 3243 25812
rect 3277 25778 3312 25812
rect 3346 25778 3381 25812
rect 3415 25778 3450 25812
rect 3484 25778 3519 25812
rect 3553 25778 3588 25812
rect 3622 25778 3657 25812
rect 3691 25778 3726 25812
rect 3760 25778 3795 25812
rect 3829 25778 3864 25812
rect 3898 25778 3933 25812
rect 3967 25778 4002 25812
rect 4036 25778 4071 25812
rect 4105 25778 4140 25812
rect 4174 25778 4208 25812
rect 4242 25778 4276 25812
rect 4310 25778 4344 25812
rect 4378 25778 4412 25812
rect 4446 25778 4480 25812
rect 4514 25778 4548 25812
rect 4582 25778 4616 25812
rect 4650 25778 4684 25812
rect 4718 25778 4752 25812
rect 4786 25778 4820 25812
rect 4854 25778 4888 25812
rect 4922 25778 4956 25812
rect 4990 25778 5024 25812
rect 5058 25778 5092 25812
rect 5126 25778 5160 25812
rect 5194 25778 5228 25812
rect 5262 25778 5296 25812
rect 5330 25778 5364 25812
rect 5398 25778 5432 25812
rect 5466 25778 5500 25812
rect 5534 25778 5568 25812
rect 5602 25778 5636 25812
rect 5670 25778 5704 25812
rect 5738 25778 5772 25812
rect 5806 25778 5840 25812
rect 5874 25778 5908 25812
rect 5942 25778 5976 25812
rect 6010 25778 6044 25812
rect 6078 25778 6112 25812
rect 6146 25778 6180 25812
rect 6214 25778 6248 25812
rect 6282 25778 6316 25812
rect 6350 25778 6384 25812
rect 6418 25778 6452 25812
rect 6486 25778 6520 25812
rect 6554 25778 6588 25812
rect 6622 25778 6656 25812
rect 6690 25778 6724 25812
rect 6758 25778 6792 25812
rect 6826 25778 6860 25812
rect 6894 25778 6928 25812
rect 6962 25778 6996 25812
rect 7030 25778 7064 25812
rect 7098 25778 7132 25812
rect 7166 25778 7200 25812
rect 7234 25778 7268 25812
rect 7302 25778 7336 25812
rect 7370 25778 7404 25812
rect 7438 25778 7472 25812
rect 7506 25778 7540 25812
rect 7574 25778 7608 25812
rect 7642 25778 7676 25812
rect 7710 25778 7744 25812
rect 7778 25778 7812 25812
rect 7846 25778 7880 25812
rect 7914 25778 7948 25812
rect 7982 25778 8016 25812
rect 8050 25778 8084 25812
rect 8118 25778 8152 25812
rect 8186 25778 8220 25812
rect 8254 25778 8288 25812
rect 8322 25778 8356 25812
rect 8390 25778 8424 25812
rect 8458 25778 8492 25812
rect 8526 25778 8560 25812
rect 8594 25778 8628 25812
rect 8662 25778 8696 25812
rect 8730 25778 8764 25812
rect 8798 25778 8832 25812
rect 8866 25778 8900 25812
rect 8934 25778 8968 25812
rect 9002 25778 9036 25812
rect 9070 25778 9104 25812
rect 9138 25778 9172 25812
rect 9206 25778 9240 25812
rect 9274 25778 9308 25812
rect 9342 25778 9376 25812
rect 9410 25778 9444 25812
rect 9478 25778 9512 25812
rect 9546 25778 9580 25812
rect 9614 25778 9648 25812
rect 9682 25778 9716 25812
rect 9750 25778 9784 25812
rect 9818 25778 9852 25812
rect 9886 25778 9920 25812
rect 9954 25778 9988 25812
rect 10022 25778 10056 25812
rect 10090 25778 10124 25812
rect 10158 25778 10192 25812
rect 10226 25778 10260 25812
rect 10294 25778 10328 25812
rect 10362 25778 10396 25812
rect 10430 25778 10464 25812
rect 10498 25778 10532 25812
rect 10566 25778 10600 25812
rect 10634 25778 10668 25812
rect 10702 25778 10736 25812
rect 10770 25778 10804 25812
rect 10838 25778 10872 25812
rect 10906 25778 10940 25812
rect 10974 25778 11008 25812
rect 11042 25778 11076 25812
rect 11110 25778 11144 25812
rect 11178 25778 11212 25812
rect 11246 25778 11280 25812
rect 11314 25778 11348 25812
rect 11382 25778 11416 25812
rect 11450 25778 11484 25812
rect 11518 25778 11552 25812
rect 11586 25778 11620 25812
rect 11654 25778 11688 25812
rect 11722 25778 11756 25812
rect 11790 25778 11824 25812
rect 11858 25778 11892 25812
rect 11926 25778 11960 25812
rect 11994 25778 12028 25812
rect 12062 25778 12096 25812
rect 12130 25778 12164 25812
rect 12198 25778 12232 25812
rect 12266 25778 12300 25812
rect 12334 25778 12368 25812
rect 12402 25778 12436 25812
rect 12470 25778 12504 25812
rect 12538 25778 12572 25812
rect 12606 25778 12640 25812
rect 12674 25778 12708 25812
rect 12742 25778 12776 25812
rect 12810 25778 12844 25812
rect 12878 25778 12912 25812
rect 12946 25778 12980 25812
rect 13014 25778 13048 25812
rect 13082 25778 13116 25812
rect 13150 25778 13184 25812
rect 13218 25778 13252 25812
rect 13286 25778 13320 25812
rect 13354 25778 13388 25812
rect 13422 25778 13456 25812
rect 13490 25778 13524 25812
rect 13558 25778 13592 25812
rect 13626 25778 13660 25812
rect 13694 25778 13728 25812
rect 13762 25778 13796 25812
rect 13830 25778 13864 25812
rect 13898 25778 13932 25812
rect 13966 25778 14000 25812
rect 14034 25778 14068 25812
rect 14102 25778 14136 25812
rect 14170 25778 14204 25812
rect 14238 25778 14272 25812
rect 14306 25778 14340 25812
rect 14374 25778 14408 25812
rect 14442 25778 14476 25812
rect 14510 25778 14544 25812
rect 14578 25778 14612 25812
rect 14646 25778 14680 25812
rect 14714 25778 14748 25812
rect 14782 25778 14816 25812
rect 14850 25778 14884 25812
rect 14918 25778 14952 25812
rect 49 25740 14952 25778
rect 49 25706 69 25740
rect 103 25706 138 25740
rect 172 25706 207 25740
rect 241 25706 276 25740
rect 310 25706 345 25740
rect 379 25706 414 25740
rect 448 25706 483 25740
rect 517 25706 552 25740
rect 586 25706 621 25740
rect 655 25706 690 25740
rect 724 25706 759 25740
rect 793 25706 828 25740
rect 862 25706 897 25740
rect 931 25706 966 25740
rect 1000 25706 1035 25740
rect 1069 25706 1104 25740
rect 1138 25706 1173 25740
rect 1207 25706 1242 25740
rect 1276 25706 1311 25740
rect 1345 25706 1380 25740
rect 1414 25706 1449 25740
rect 1483 25706 1518 25740
rect 1552 25706 1587 25740
rect 1621 25706 1656 25740
rect 1690 25706 1725 25740
rect 1759 25706 1794 25740
rect 1828 25706 1863 25740
rect 1897 25706 1932 25740
rect 1966 25706 2001 25740
rect 2035 25706 2070 25740
rect 2104 25706 2139 25740
rect 2173 25706 2208 25740
rect 2242 25706 2277 25740
rect 2311 25706 2346 25740
rect 2380 25706 2415 25740
rect 2449 25706 2484 25740
rect 2518 25706 2553 25740
rect 2587 25706 2622 25740
rect 2656 25706 2691 25740
rect 2725 25706 2760 25740
rect 2794 25706 2829 25740
rect 2863 25706 2898 25740
rect 2932 25706 2967 25740
rect 3001 25706 3036 25740
rect 3070 25706 3105 25740
rect 3139 25706 3174 25740
rect 3208 25706 3243 25740
rect 3277 25706 3312 25740
rect 3346 25706 3381 25740
rect 3415 25706 3450 25740
rect 3484 25706 3519 25740
rect 3553 25706 3588 25740
rect 3622 25706 3657 25740
rect 3691 25706 3726 25740
rect 3760 25706 3795 25740
rect 3829 25706 3864 25740
rect 3898 25706 3933 25740
rect 3967 25706 4002 25740
rect 4036 25706 4071 25740
rect 4105 25706 4140 25740
rect 4174 25706 4208 25740
rect 4242 25706 4276 25740
rect 4310 25706 4344 25740
rect 4378 25706 4412 25740
rect 4446 25706 4480 25740
rect 4514 25706 4548 25740
rect 4582 25706 4616 25740
rect 4650 25706 4684 25740
rect 4718 25706 4752 25740
rect 4786 25706 4820 25740
rect 4854 25706 4888 25740
rect 4922 25706 4956 25740
rect 4990 25706 5024 25740
rect 5058 25706 5092 25740
rect 5126 25706 5160 25740
rect 5194 25706 5228 25740
rect 5262 25706 5296 25740
rect 5330 25706 5364 25740
rect 5398 25706 5432 25740
rect 5466 25706 5500 25740
rect 5534 25706 5568 25740
rect 5602 25706 5636 25740
rect 5670 25706 5704 25740
rect 5738 25706 5772 25740
rect 5806 25706 5840 25740
rect 5874 25706 5908 25740
rect 5942 25706 5976 25740
rect 6010 25706 6044 25740
rect 6078 25706 6112 25740
rect 6146 25706 6180 25740
rect 6214 25706 6248 25740
rect 6282 25706 6316 25740
rect 6350 25706 6384 25740
rect 6418 25706 6452 25740
rect 6486 25706 6520 25740
rect 6554 25706 6588 25740
rect 6622 25706 6656 25740
rect 6690 25706 6724 25740
rect 6758 25706 6792 25740
rect 6826 25706 6860 25740
rect 6894 25706 6928 25740
rect 6962 25706 6996 25740
rect 7030 25706 7064 25740
rect 7098 25706 7132 25740
rect 7166 25706 7200 25740
rect 7234 25706 7268 25740
rect 7302 25706 7336 25740
rect 7370 25706 7404 25740
rect 7438 25706 7472 25740
rect 7506 25706 7540 25740
rect 7574 25706 7608 25740
rect 7642 25706 7676 25740
rect 7710 25706 7744 25740
rect 7778 25706 7812 25740
rect 7846 25706 7880 25740
rect 7914 25706 7948 25740
rect 7982 25706 8016 25740
rect 8050 25706 8084 25740
rect 8118 25706 8152 25740
rect 8186 25706 8220 25740
rect 8254 25706 8288 25740
rect 8322 25706 8356 25740
rect 8390 25706 8424 25740
rect 8458 25706 8492 25740
rect 8526 25706 8560 25740
rect 8594 25706 8628 25740
rect 8662 25706 8696 25740
rect 8730 25706 8764 25740
rect 8798 25706 8832 25740
rect 8866 25706 8900 25740
rect 8934 25706 8968 25740
rect 9002 25706 9036 25740
rect 9070 25706 9104 25740
rect 9138 25706 9172 25740
rect 9206 25706 9240 25740
rect 9274 25706 9308 25740
rect 9342 25706 9376 25740
rect 9410 25706 9444 25740
rect 9478 25706 9512 25740
rect 9546 25706 9580 25740
rect 9614 25706 9648 25740
rect 9682 25706 9716 25740
rect 9750 25706 9784 25740
rect 9818 25706 9852 25740
rect 9886 25706 9920 25740
rect 9954 25706 9988 25740
rect 10022 25706 10056 25740
rect 10090 25706 10124 25740
rect 10158 25706 10192 25740
rect 10226 25706 10260 25740
rect 10294 25706 10328 25740
rect 10362 25706 10396 25740
rect 10430 25706 10464 25740
rect 10498 25706 10532 25740
rect 10566 25706 10600 25740
rect 10634 25706 10668 25740
rect 10702 25706 10736 25740
rect 10770 25706 10804 25740
rect 10838 25706 10872 25740
rect 10906 25706 10940 25740
rect 10974 25706 11008 25740
rect 11042 25706 11076 25740
rect 11110 25706 11144 25740
rect 11178 25706 11212 25740
rect 11246 25706 11280 25740
rect 11314 25706 11348 25740
rect 11382 25706 11416 25740
rect 11450 25706 11484 25740
rect 11518 25706 11552 25740
rect 11586 25706 11620 25740
rect 11654 25706 11688 25740
rect 11722 25706 11756 25740
rect 11790 25706 11824 25740
rect 11858 25706 11892 25740
rect 11926 25706 11960 25740
rect 11994 25706 12028 25740
rect 12062 25706 12096 25740
rect 12130 25706 12164 25740
rect 12198 25706 12232 25740
rect 12266 25706 12300 25740
rect 12334 25706 12368 25740
rect 12402 25706 12436 25740
rect 12470 25706 12504 25740
rect 12538 25706 12572 25740
rect 12606 25706 12640 25740
rect 12674 25706 12708 25740
rect 12742 25706 12776 25740
rect 12810 25706 12844 25740
rect 12878 25706 12912 25740
rect 12946 25706 12980 25740
rect 13014 25706 13048 25740
rect 13082 25706 13116 25740
rect 13150 25706 13184 25740
rect 13218 25706 13252 25740
rect 13286 25706 13320 25740
rect 13354 25706 13388 25740
rect 13422 25706 13456 25740
rect 13490 25706 13524 25740
rect 13558 25706 13592 25740
rect 13626 25706 13660 25740
rect 13694 25706 13728 25740
rect 13762 25706 13796 25740
rect 13830 25706 13864 25740
rect 13898 25706 13932 25740
rect 13966 25706 14000 25740
rect 14034 25706 14068 25740
rect 14102 25706 14136 25740
rect 14170 25706 14204 25740
rect 14238 25706 14272 25740
rect 14306 25706 14340 25740
rect 14374 25706 14408 25740
rect 14442 25706 14476 25740
rect 14510 25706 14544 25740
rect 14578 25706 14612 25740
rect 14646 25706 14680 25740
rect 14714 25706 14748 25740
rect 14782 25706 14816 25740
rect 14850 25706 14884 25740
rect 14918 25706 14952 25740
rect 49 25668 14952 25706
rect 49 25634 69 25668
rect 103 25634 138 25668
rect 172 25634 207 25668
rect 241 25634 276 25668
rect 310 25634 345 25668
rect 379 25634 414 25668
rect 448 25634 483 25668
rect 517 25634 552 25668
rect 586 25634 621 25668
rect 655 25634 690 25668
rect 724 25634 759 25668
rect 793 25634 828 25668
rect 862 25634 897 25668
rect 931 25634 966 25668
rect 1000 25634 1035 25668
rect 1069 25634 1104 25668
rect 1138 25634 1173 25668
rect 1207 25634 1242 25668
rect 1276 25634 1311 25668
rect 1345 25634 1380 25668
rect 1414 25634 1449 25668
rect 1483 25634 1518 25668
rect 1552 25634 1587 25668
rect 1621 25634 1656 25668
rect 1690 25634 1725 25668
rect 1759 25634 1794 25668
rect 1828 25634 1863 25668
rect 1897 25634 1932 25668
rect 1966 25634 2001 25668
rect 2035 25634 2070 25668
rect 2104 25634 2139 25668
rect 2173 25634 2208 25668
rect 2242 25634 2277 25668
rect 2311 25634 2346 25668
rect 2380 25634 2415 25668
rect 2449 25634 2484 25668
rect 2518 25634 2553 25668
rect 2587 25634 2622 25668
rect 2656 25634 2691 25668
rect 2725 25634 2760 25668
rect 2794 25634 2829 25668
rect 2863 25634 2898 25668
rect 2932 25634 2967 25668
rect 3001 25634 3036 25668
rect 3070 25634 3105 25668
rect 3139 25634 3174 25668
rect 3208 25634 3243 25668
rect 3277 25634 3312 25668
rect 3346 25634 3381 25668
rect 3415 25634 3450 25668
rect 3484 25634 3519 25668
rect 3553 25634 3588 25668
rect 3622 25634 3657 25668
rect 3691 25634 3726 25668
rect 3760 25634 3795 25668
rect 3829 25634 3864 25668
rect 3898 25634 3933 25668
rect 3967 25634 4002 25668
rect 4036 25634 4071 25668
rect 4105 25634 4140 25668
rect 4174 25634 4208 25668
rect 4242 25634 4276 25668
rect 4310 25634 4344 25668
rect 4378 25634 4412 25668
rect 4446 25634 4480 25668
rect 4514 25634 4548 25668
rect 4582 25634 4616 25668
rect 4650 25634 4684 25668
rect 4718 25634 4752 25668
rect 4786 25634 4820 25668
rect 4854 25634 4888 25668
rect 4922 25634 4956 25668
rect 4990 25634 5024 25668
rect 5058 25634 5092 25668
rect 5126 25634 5160 25668
rect 5194 25634 5228 25668
rect 5262 25634 5296 25668
rect 5330 25634 5364 25668
rect 5398 25634 5432 25668
rect 5466 25634 5500 25668
rect 5534 25634 5568 25668
rect 5602 25634 5636 25668
rect 5670 25634 5704 25668
rect 5738 25634 5772 25668
rect 5806 25634 5840 25668
rect 5874 25634 5908 25668
rect 5942 25634 5976 25668
rect 6010 25634 6044 25668
rect 6078 25634 6112 25668
rect 6146 25634 6180 25668
rect 6214 25634 6248 25668
rect 6282 25634 6316 25668
rect 6350 25634 6384 25668
rect 6418 25634 6452 25668
rect 6486 25634 6520 25668
rect 6554 25634 6588 25668
rect 6622 25634 6656 25668
rect 6690 25634 6724 25668
rect 6758 25634 6792 25668
rect 6826 25634 6860 25668
rect 6894 25634 6928 25668
rect 6962 25634 6996 25668
rect 7030 25634 7064 25668
rect 7098 25634 7132 25668
rect 7166 25634 7200 25668
rect 7234 25634 7268 25668
rect 7302 25634 7336 25668
rect 7370 25634 7404 25668
rect 7438 25634 7472 25668
rect 7506 25634 7540 25668
rect 7574 25634 7608 25668
rect 7642 25634 7676 25668
rect 7710 25634 7744 25668
rect 7778 25634 7812 25668
rect 7846 25634 7880 25668
rect 7914 25634 7948 25668
rect 7982 25634 8016 25668
rect 8050 25634 8084 25668
rect 8118 25634 8152 25668
rect 8186 25634 8220 25668
rect 8254 25634 8288 25668
rect 8322 25634 8356 25668
rect 8390 25634 8424 25668
rect 8458 25634 8492 25668
rect 8526 25634 8560 25668
rect 8594 25634 8628 25668
rect 8662 25634 8696 25668
rect 8730 25634 8764 25668
rect 8798 25634 8832 25668
rect 8866 25634 8900 25668
rect 8934 25634 8968 25668
rect 9002 25634 9036 25668
rect 9070 25634 9104 25668
rect 9138 25634 9172 25668
rect 9206 25634 9240 25668
rect 9274 25634 9308 25668
rect 9342 25634 9376 25668
rect 9410 25634 9444 25668
rect 9478 25634 9512 25668
rect 9546 25634 9580 25668
rect 9614 25634 9648 25668
rect 9682 25634 9716 25668
rect 9750 25634 9784 25668
rect 9818 25634 9852 25668
rect 9886 25634 9920 25668
rect 9954 25634 9988 25668
rect 10022 25634 10056 25668
rect 10090 25634 10124 25668
rect 10158 25634 10192 25668
rect 10226 25634 10260 25668
rect 10294 25634 10328 25668
rect 10362 25634 10396 25668
rect 10430 25634 10464 25668
rect 10498 25634 10532 25668
rect 10566 25634 10600 25668
rect 10634 25634 10668 25668
rect 10702 25634 10736 25668
rect 10770 25634 10804 25668
rect 10838 25634 10872 25668
rect 10906 25634 10940 25668
rect 10974 25634 11008 25668
rect 11042 25634 11076 25668
rect 11110 25634 11144 25668
rect 11178 25634 11212 25668
rect 11246 25634 11280 25668
rect 11314 25634 11348 25668
rect 11382 25634 11416 25668
rect 11450 25634 11484 25668
rect 11518 25634 11552 25668
rect 11586 25634 11620 25668
rect 11654 25634 11688 25668
rect 11722 25634 11756 25668
rect 11790 25634 11824 25668
rect 11858 25634 11892 25668
rect 11926 25634 11960 25668
rect 11994 25634 12028 25668
rect 12062 25634 12096 25668
rect 12130 25634 12164 25668
rect 12198 25634 12232 25668
rect 12266 25634 12300 25668
rect 12334 25634 12368 25668
rect 12402 25634 12436 25668
rect 12470 25634 12504 25668
rect 12538 25634 12572 25668
rect 12606 25634 12640 25668
rect 12674 25634 12708 25668
rect 12742 25634 12776 25668
rect 12810 25634 12844 25668
rect 12878 25634 12912 25668
rect 12946 25634 12980 25668
rect 13014 25634 13048 25668
rect 13082 25634 13116 25668
rect 13150 25634 13184 25668
rect 13218 25634 13252 25668
rect 13286 25634 13320 25668
rect 13354 25634 13388 25668
rect 13422 25634 13456 25668
rect 13490 25634 13524 25668
rect 13558 25634 13592 25668
rect 13626 25634 13660 25668
rect 13694 25634 13728 25668
rect 13762 25634 13796 25668
rect 13830 25634 13864 25668
rect 13898 25634 13932 25668
rect 13966 25634 14000 25668
rect 14034 25634 14068 25668
rect 14102 25634 14136 25668
rect 14170 25634 14204 25668
rect 14238 25634 14272 25668
rect 14306 25634 14340 25668
rect 14374 25634 14408 25668
rect 14442 25634 14476 25668
rect 14510 25634 14544 25668
rect 14578 25634 14612 25668
rect 14646 25634 14680 25668
rect 14714 25634 14748 25668
rect 14782 25634 14816 25668
rect 14850 25634 14884 25668
rect 14918 25634 14952 25668
rect 49 25599 14952 25634
<< mvpsubdiffcont >>
rect 121 28249 155 28283
rect 190 28249 224 28283
rect 259 28249 293 28283
rect 328 28249 362 28283
rect 397 28249 431 28283
rect 466 28249 500 28283
rect 535 28249 569 28283
rect 604 28249 638 28283
rect 673 28249 707 28283
rect 742 28249 776 28283
rect 811 28249 845 28283
rect 880 28249 914 28283
rect 949 28249 983 28283
rect 1018 28249 1052 28283
rect 1087 28249 1121 28283
rect 121 28181 155 28215
rect 190 28181 224 28215
rect 259 28181 293 28215
rect 328 28181 362 28215
rect 397 28181 431 28215
rect 466 28181 500 28215
rect 535 28181 569 28215
rect 604 28181 638 28215
rect 673 28181 707 28215
rect 742 28181 776 28215
rect 811 28181 845 28215
rect 880 28181 914 28215
rect 949 28181 983 28215
rect 1018 28181 1052 28215
rect 1087 28181 1121 28215
rect 121 28113 155 28147
rect 190 28113 224 28147
rect 259 28113 293 28147
rect 328 28113 362 28147
rect 397 28113 431 28147
rect 466 28113 500 28147
rect 535 28113 569 28147
rect 604 28113 638 28147
rect 673 28113 707 28147
rect 742 28113 776 28147
rect 811 28113 845 28147
rect 880 28113 914 28147
rect 949 28113 983 28147
rect 1018 28113 1052 28147
rect 1087 28113 1121 28147
rect 121 28045 155 28079
rect 190 28045 224 28079
rect 259 28045 293 28079
rect 328 28045 362 28079
rect 397 28045 431 28079
rect 466 28045 500 28079
rect 535 28045 569 28079
rect 604 28045 638 28079
rect 673 28045 707 28079
rect 742 28045 776 28079
rect 811 28045 845 28079
rect 880 28045 914 28079
rect 949 28045 983 28079
rect 1018 28045 1052 28079
rect 1087 28045 1121 28079
rect 121 27977 155 28011
rect 190 27977 224 28011
rect 259 27977 293 28011
rect 328 27977 362 28011
rect 397 27977 431 28011
rect 466 27977 500 28011
rect 535 27977 569 28011
rect 604 27977 638 28011
rect 673 27977 707 28011
rect 742 27977 776 28011
rect 811 27977 845 28011
rect 880 27977 914 28011
rect 949 27977 983 28011
rect 1018 27977 1052 28011
rect 1087 27977 1121 28011
rect 121 27909 155 27943
rect 190 27909 224 27943
rect 259 27909 293 27943
rect 328 27909 362 27943
rect 397 27909 431 27943
rect 466 27909 500 27943
rect 535 27909 569 27943
rect 604 27909 638 27943
rect 673 27909 707 27943
rect 742 27909 776 27943
rect 811 27909 845 27943
rect 880 27909 914 27943
rect 949 27909 983 27943
rect 1018 27909 1052 27943
rect 1087 27909 1121 27943
rect 121 27841 155 27875
rect 190 27841 224 27875
rect 259 27841 293 27875
rect 328 27841 362 27875
rect 397 27841 431 27875
rect 466 27841 500 27875
rect 535 27841 569 27875
rect 604 27841 638 27875
rect 673 27841 707 27875
rect 742 27841 776 27875
rect 811 27841 845 27875
rect 880 27841 914 27875
rect 949 27841 983 27875
rect 1018 27841 1052 27875
rect 1087 27841 1121 27875
rect 121 27773 155 27807
rect 190 27773 224 27807
rect 259 27773 293 27807
rect 328 27773 362 27807
rect 397 27773 431 27807
rect 466 27773 500 27807
rect 535 27773 569 27807
rect 604 27773 638 27807
rect 673 27773 707 27807
rect 742 27773 776 27807
rect 811 27773 845 27807
rect 880 27773 914 27807
rect 949 27773 983 27807
rect 1018 27773 1052 27807
rect 1087 27773 1121 27807
rect 121 27705 155 27739
rect 190 27705 224 27739
rect 259 27705 293 27739
rect 328 27705 362 27739
rect 397 27705 431 27739
rect 466 27705 500 27739
rect 535 27705 569 27739
rect 604 27705 638 27739
rect 673 27705 707 27739
rect 742 27705 776 27739
rect 811 27705 845 27739
rect 880 27705 914 27739
rect 949 27705 983 27739
rect 1018 27705 1052 27739
rect 1087 27705 1121 27739
rect 121 27637 155 27671
rect 190 27637 224 27671
rect 259 27637 293 27671
rect 328 27637 362 27671
rect 397 27637 431 27671
rect 466 27637 500 27671
rect 535 27637 569 27671
rect 604 27637 638 27671
rect 673 27637 707 27671
rect 742 27637 776 27671
rect 811 27637 845 27671
rect 880 27637 914 27671
rect 949 27637 983 27671
rect 1018 27637 1052 27671
rect 1087 27637 1121 27671
rect 121 27569 155 27603
rect 190 27569 224 27603
rect 259 27569 293 27603
rect 328 27569 362 27603
rect 397 27569 431 27603
rect 466 27569 500 27603
rect 535 27569 569 27603
rect 604 27569 638 27603
rect 673 27569 707 27603
rect 742 27569 776 27603
rect 811 27569 845 27603
rect 880 27569 914 27603
rect 949 27569 983 27603
rect 1018 27569 1052 27603
rect 1087 27569 1121 27603
rect 1156 27569 14858 28283
rect 77 25410 111 25444
rect 146 25410 180 25444
rect 215 25410 249 25444
rect 284 25410 318 25444
rect 353 25410 387 25444
rect 422 25410 456 25444
rect 491 25410 525 25444
rect 560 25410 594 25444
rect 629 25410 663 25444
rect 698 25410 732 25444
rect 766 25410 800 25444
rect 834 25410 868 25444
rect 902 25410 936 25444
rect 970 25410 1004 25444
rect 1038 25410 1072 25444
rect 1106 25410 1140 25444
rect 1174 25410 1208 25444
rect 1242 25410 1276 25444
rect 1310 25410 1344 25444
rect 1378 25410 1412 25444
rect 1446 25410 1480 25444
rect 1514 25410 1548 25444
rect 1582 25410 1616 25444
rect 1650 25410 1684 25444
rect 1718 25410 1752 25444
rect 1786 25410 1820 25444
rect 1854 25410 1888 25444
rect 1922 25410 1956 25444
rect 1990 25410 2024 25444
rect 2058 25410 2092 25444
rect 2126 25410 2160 25444
rect 2194 25410 2228 25444
rect 2262 25410 2296 25444
rect 2330 25410 2364 25444
rect 2398 25410 2432 25444
rect 2466 25410 2500 25444
rect 2534 25410 2568 25444
rect 2602 25410 2636 25444
rect 2670 25410 2704 25444
rect 2738 25410 2772 25444
rect 2806 25410 2840 25444
rect 2874 25410 2908 25444
rect 2942 25410 2976 25444
rect 3010 25410 3044 25444
rect 3078 25410 3112 25444
rect 3146 25410 3180 25444
rect 3214 25410 3248 25444
rect 3282 25410 3316 25444
rect 3350 25410 3384 25444
rect 3418 25410 3452 25444
rect 3486 25410 3520 25444
rect 3554 25410 3588 25444
rect 3622 25410 3656 25444
rect 3690 25410 3724 25444
rect 3758 25410 3792 25444
rect 3826 25410 3860 25444
rect 3894 25410 3928 25444
rect 3962 25410 3996 25444
rect 4030 25410 4064 25444
rect 4098 25410 4132 25444
rect 4166 25410 4200 25444
rect 4234 25410 4268 25444
rect 4302 25410 4336 25444
rect 4370 25410 4404 25444
rect 4438 25410 4472 25444
rect 4506 25410 4540 25444
rect 4574 25410 4608 25444
rect 4642 25410 4676 25444
rect 4710 25410 4744 25444
rect 4778 25410 4812 25444
rect 4846 25410 4880 25444
rect 4914 25410 4948 25444
rect 4982 25410 5016 25444
rect 5050 25410 5084 25444
rect 5118 25410 5152 25444
rect 5186 25410 5220 25444
rect 5254 25410 5288 25444
rect 5322 25410 5356 25444
rect 5390 25410 5424 25444
rect 5458 25410 5492 25444
rect 5526 25410 5560 25444
rect 5594 25410 5628 25444
rect 5662 25410 5696 25444
rect 5730 25410 5764 25444
rect 5798 25410 5832 25444
rect 5866 25410 5900 25444
rect 5934 25410 5968 25444
rect 6002 25410 6036 25444
rect 6070 25410 6104 25444
rect 6138 25410 6172 25444
rect 6206 25410 6240 25444
rect 6274 25410 6308 25444
rect 6342 25410 6376 25444
rect 6410 25410 6444 25444
rect 6478 25410 6512 25444
rect 6546 25410 6580 25444
rect 6614 25410 6648 25444
rect 6682 25410 6716 25444
rect 6750 25410 6784 25444
rect 6818 25410 6852 25444
rect 6886 25410 6920 25444
rect 6954 25410 6988 25444
rect 7022 25410 7056 25444
rect 7090 25410 7124 25444
rect 7158 25410 7192 25444
rect 7226 25410 7260 25444
rect 7294 25410 7328 25444
rect 7362 25410 7396 25444
rect 7430 25410 7464 25444
rect 7498 25410 7532 25444
rect 7566 25410 7600 25444
rect 7634 25410 7668 25444
rect 7702 25410 7736 25444
rect 7770 25410 7804 25444
rect 7838 25410 7872 25444
rect 7906 25410 7940 25444
rect 7974 25410 8008 25444
rect 8042 25410 8076 25444
rect 8110 25410 8144 25444
rect 8178 25410 8212 25444
rect 8246 25410 8280 25444
rect 77 25324 111 25358
rect 146 25324 180 25358
rect 215 25324 249 25358
rect 284 25324 318 25358
rect 353 25324 387 25358
rect 422 25324 456 25358
rect 491 25324 525 25358
rect 560 25324 594 25358
rect 629 25324 663 25358
rect 698 25324 732 25358
rect 766 25324 800 25358
rect 834 25324 868 25358
rect 902 25324 936 25358
rect 970 25324 1004 25358
rect 1038 25324 1072 25358
rect 1106 25324 1140 25358
rect 1174 25324 1208 25358
rect 1242 25324 1276 25358
rect 1310 25324 1344 25358
rect 1378 25324 1412 25358
rect 1446 25324 1480 25358
rect 1514 25324 1548 25358
rect 1582 25324 1616 25358
rect 1650 25324 1684 25358
rect 1718 25324 1752 25358
rect 1786 25324 1820 25358
rect 1854 25324 1888 25358
rect 1922 25324 1956 25358
rect 1990 25324 2024 25358
rect 2058 25324 2092 25358
rect 2126 25324 2160 25358
rect 2194 25324 2228 25358
rect 2262 25324 2296 25358
rect 2330 25324 2364 25358
rect 2398 25324 2432 25358
rect 2466 25324 2500 25358
rect 2534 25324 2568 25358
rect 2602 25324 2636 25358
rect 2670 25324 2704 25358
rect 2738 25324 2772 25358
rect 2806 25324 2840 25358
rect 2874 25324 2908 25358
rect 2942 25324 2976 25358
rect 3010 25324 3044 25358
rect 3078 25324 3112 25358
rect 3146 25324 3180 25358
rect 3214 25324 3248 25358
rect 3282 25324 3316 25358
rect 3350 25324 3384 25358
rect 3418 25324 3452 25358
rect 3486 25324 3520 25358
rect 3554 25324 3588 25358
rect 3622 25324 3656 25358
rect 3690 25324 3724 25358
rect 3758 25324 3792 25358
rect 3826 25324 3860 25358
rect 3894 25324 3928 25358
rect 3962 25324 3996 25358
rect 4030 25324 4064 25358
rect 4098 25324 4132 25358
rect 4166 25324 4200 25358
rect 4234 25324 4268 25358
rect 4302 25324 4336 25358
rect 4370 25324 4404 25358
rect 4438 25324 4472 25358
rect 4506 25324 4540 25358
rect 4574 25324 4608 25358
rect 4642 25324 4676 25358
rect 4710 25324 4744 25358
rect 4778 25324 4812 25358
rect 4846 25324 4880 25358
rect 4914 25324 4948 25358
rect 4982 25324 5016 25358
rect 5050 25324 5084 25358
rect 5118 25324 5152 25358
rect 5186 25324 5220 25358
rect 5254 25324 5288 25358
rect 5322 25324 5356 25358
rect 5390 25324 5424 25358
rect 5458 25324 5492 25358
rect 5526 25324 5560 25358
rect 5594 25324 5628 25358
rect 5662 25324 5696 25358
rect 5730 25324 5764 25358
rect 5798 25324 5832 25358
rect 5866 25324 5900 25358
rect 5934 25324 5968 25358
rect 6002 25324 6036 25358
rect 6070 25324 6104 25358
rect 6138 25324 6172 25358
rect 6206 25324 6240 25358
rect 6274 25324 6308 25358
rect 6342 25324 6376 25358
rect 6410 25324 6444 25358
rect 6478 25324 6512 25358
rect 6546 25324 6580 25358
rect 6614 25324 6648 25358
rect 6682 25324 6716 25358
rect 6750 25324 6784 25358
rect 6818 25324 6852 25358
rect 6886 25324 6920 25358
rect 6954 25324 6988 25358
rect 7022 25324 7056 25358
rect 7090 25324 7124 25358
rect 7158 25324 7192 25358
rect 7226 25324 7260 25358
rect 7294 25324 7328 25358
rect 7362 25324 7396 25358
rect 7430 25324 7464 25358
rect 7498 25324 7532 25358
rect 7566 25324 7600 25358
rect 7634 25324 7668 25358
rect 7702 25324 7736 25358
rect 7770 25324 7804 25358
rect 7838 25324 7872 25358
rect 7906 25324 7940 25358
rect 7974 25324 8008 25358
rect 8042 25324 8076 25358
rect 8110 25324 8144 25358
rect 8178 25324 8212 25358
rect 8246 25324 8280 25358
rect 77 25238 111 25272
rect 146 25238 180 25272
rect 215 25238 249 25272
rect 284 25238 318 25272
rect 353 25238 387 25272
rect 422 25238 456 25272
rect 491 25238 525 25272
rect 560 25238 594 25272
rect 629 25238 663 25272
rect 698 25238 732 25272
rect 766 25238 800 25272
rect 834 25238 868 25272
rect 902 25238 936 25272
rect 970 25238 1004 25272
rect 1038 25238 1072 25272
rect 1106 25238 1140 25272
rect 1174 25238 1208 25272
rect 1242 25238 1276 25272
rect 1310 25238 1344 25272
rect 1378 25238 1412 25272
rect 1446 25238 1480 25272
rect 1514 25238 1548 25272
rect 1582 25238 1616 25272
rect 1650 25238 1684 25272
rect 1718 25238 1752 25272
rect 1786 25238 1820 25272
rect 1854 25238 1888 25272
rect 1922 25238 1956 25272
rect 1990 25238 2024 25272
rect 2058 25238 2092 25272
rect 2126 25238 2160 25272
rect 2194 25238 2228 25272
rect 2262 25238 2296 25272
rect 2330 25238 2364 25272
rect 2398 25238 2432 25272
rect 2466 25238 2500 25272
rect 2534 25238 2568 25272
rect 2602 25238 2636 25272
rect 2670 25238 2704 25272
rect 2738 25238 2772 25272
rect 2806 25238 2840 25272
rect 2874 25238 2908 25272
rect 2942 25238 2976 25272
rect 3010 25238 3044 25272
rect 3078 25238 3112 25272
rect 3146 25238 3180 25272
rect 3214 25238 3248 25272
rect 3282 25238 3316 25272
rect 3350 25238 3384 25272
rect 3418 25238 3452 25272
rect 3486 25238 3520 25272
rect 3554 25238 3588 25272
rect 3622 25238 3656 25272
rect 3690 25238 3724 25272
rect 3758 25238 3792 25272
rect 3826 25238 3860 25272
rect 3894 25238 3928 25272
rect 3962 25238 3996 25272
rect 4030 25238 4064 25272
rect 4098 25238 4132 25272
rect 4166 25238 4200 25272
rect 4234 25238 4268 25272
rect 4302 25238 4336 25272
rect 4370 25238 4404 25272
rect 4438 25238 4472 25272
rect 4506 25238 4540 25272
rect 4574 25238 4608 25272
rect 4642 25238 4676 25272
rect 4710 25238 4744 25272
rect 4778 25238 4812 25272
rect 4846 25238 4880 25272
rect 4914 25238 4948 25272
rect 4982 25238 5016 25272
rect 5050 25238 5084 25272
rect 5118 25238 5152 25272
rect 5186 25238 5220 25272
rect 5254 25238 5288 25272
rect 5322 25238 5356 25272
rect 5390 25238 5424 25272
rect 5458 25238 5492 25272
rect 5526 25238 5560 25272
rect 5594 25238 5628 25272
rect 5662 25238 5696 25272
rect 5730 25238 5764 25272
rect 5798 25238 5832 25272
rect 5866 25238 5900 25272
rect 5934 25238 5968 25272
rect 6002 25238 6036 25272
rect 6070 25238 6104 25272
rect 6138 25238 6172 25272
rect 6206 25238 6240 25272
rect 6274 25238 6308 25272
rect 6342 25238 6376 25272
rect 6410 25238 6444 25272
rect 6478 25238 6512 25272
rect 6546 25238 6580 25272
rect 6614 25238 6648 25272
rect 6682 25238 6716 25272
rect 6750 25238 6784 25272
rect 6818 25238 6852 25272
rect 6886 25238 6920 25272
rect 6954 25238 6988 25272
rect 7022 25238 7056 25272
rect 7090 25238 7124 25272
rect 7158 25238 7192 25272
rect 7226 25238 7260 25272
rect 7294 25238 7328 25272
rect 7362 25238 7396 25272
rect 7430 25238 7464 25272
rect 7498 25238 7532 25272
rect 7566 25238 7600 25272
rect 7634 25238 7668 25272
rect 7702 25238 7736 25272
rect 7770 25238 7804 25272
rect 7838 25238 7872 25272
rect 7906 25238 7940 25272
rect 7974 25238 8008 25272
rect 8042 25238 8076 25272
rect 8110 25238 8144 25272
rect 8178 25238 8212 25272
rect 8246 25238 8280 25272
rect 12432 25410 12466 25444
rect 12501 25410 12535 25444
rect 12570 25410 12604 25444
rect 12639 25410 12673 25444
rect 12708 25410 12742 25444
rect 12777 25410 12811 25444
rect 12846 25410 12880 25444
rect 12915 25410 12949 25444
rect 12984 25410 13018 25444
rect 13053 25410 13087 25444
rect 13122 25410 13156 25444
rect 13191 25410 13225 25444
rect 13260 25410 13294 25444
rect 13328 25410 13362 25444
rect 13396 25410 13430 25444
rect 13464 25410 13498 25444
rect 13532 25410 13566 25444
rect 13600 25410 13634 25444
rect 13668 25410 13702 25444
rect 13736 25410 13770 25444
rect 13804 25410 13838 25444
rect 13872 25410 13906 25444
rect 13940 25410 13974 25444
rect 14008 25410 14042 25444
rect 14076 25410 14110 25444
rect 14144 25410 14178 25444
rect 14212 25410 14246 25444
rect 14280 25410 14314 25444
rect 14348 25410 14382 25444
rect 14416 25410 14450 25444
rect 14484 25410 14518 25444
rect 14552 25410 14586 25444
rect 14620 25410 14654 25444
rect 14688 25410 14722 25444
rect 14756 25410 14790 25444
rect 14824 25410 14858 25444
rect 12432 25324 12466 25358
rect 12501 25324 12535 25358
rect 12570 25324 12604 25358
rect 12639 25324 12673 25358
rect 12708 25324 12742 25358
rect 12777 25324 12811 25358
rect 12846 25324 12880 25358
rect 12915 25324 12949 25358
rect 12984 25324 13018 25358
rect 13053 25324 13087 25358
rect 13122 25324 13156 25358
rect 13191 25324 13225 25358
rect 13260 25324 13294 25358
rect 13328 25324 13362 25358
rect 13396 25324 13430 25358
rect 13464 25324 13498 25358
rect 13532 25324 13566 25358
rect 13600 25324 13634 25358
rect 13668 25324 13702 25358
rect 13736 25324 13770 25358
rect 13804 25324 13838 25358
rect 13872 25324 13906 25358
rect 13940 25324 13974 25358
rect 14008 25324 14042 25358
rect 14076 25324 14110 25358
rect 14144 25324 14178 25358
rect 14212 25324 14246 25358
rect 14280 25324 14314 25358
rect 14348 25324 14382 25358
rect 14416 25324 14450 25358
rect 14484 25324 14518 25358
rect 14552 25324 14586 25358
rect 14620 25324 14654 25358
rect 14688 25324 14722 25358
rect 14756 25324 14790 25358
rect 14824 25324 14858 25358
rect 12432 25238 12466 25272
rect 12501 25238 12535 25272
rect 12570 25238 12604 25272
rect 12639 25238 12673 25272
rect 12708 25238 12742 25272
rect 12777 25238 12811 25272
rect 12846 25238 12880 25272
rect 12915 25238 12949 25272
rect 12984 25238 13018 25272
rect 13053 25238 13087 25272
rect 13122 25238 13156 25272
rect 13191 25238 13225 25272
rect 13260 25238 13294 25272
rect 13328 25238 13362 25272
rect 13396 25238 13430 25272
rect 13464 25238 13498 25272
rect 13532 25238 13566 25272
rect 13600 25238 13634 25272
rect 13668 25238 13702 25272
rect 13736 25238 13770 25272
rect 13804 25238 13838 25272
rect 13872 25238 13906 25272
rect 13940 25238 13974 25272
rect 14008 25238 14042 25272
rect 14076 25238 14110 25272
rect 14144 25238 14178 25272
rect 14212 25238 14246 25272
rect 14280 25238 14314 25272
rect 14348 25238 14382 25272
rect 14416 25238 14450 25272
rect 14484 25238 14518 25272
rect 14552 25238 14586 25272
rect 14620 25238 14654 25272
rect 14688 25238 14722 25272
rect 14756 25238 14790 25272
rect 14824 25238 14858 25272
rect 124 25144 158 25178
rect 193 25144 227 25178
rect 262 25144 296 25178
rect 331 25144 365 25178
rect 400 25144 434 25178
rect 469 25144 503 25178
rect 538 25144 572 25178
rect 607 25144 641 25178
rect 676 25144 710 25178
rect 745 25144 779 25178
rect 814 25144 848 25178
rect 883 25144 917 25178
rect 952 25144 986 25178
rect 1020 25144 1054 25178
rect 1088 25144 1122 25178
rect 1156 25144 1190 25178
rect 1224 25144 1258 25178
rect 1292 25144 1326 25178
rect 1360 25144 1394 25178
rect 1428 25144 1462 25178
rect 1496 25144 1530 25178
rect 1564 25144 1598 25178
rect 1632 25144 1666 25178
rect 1700 25144 1734 25178
rect 1768 25144 1802 25178
rect 1836 25144 1870 25178
rect 1904 25144 1938 25178
rect 1972 25144 2006 25178
rect 2040 25144 2074 25178
rect 2108 25144 2142 25178
rect 2176 25144 2210 25178
rect 2244 25144 2278 25178
rect 2312 25144 2346 25178
rect 2380 25144 2414 25178
rect 2448 25144 2482 25178
rect 2516 25144 2550 25178
rect 2584 25144 2618 25178
rect 2652 25144 2686 25178
rect 2720 25144 2754 25178
rect 2788 25144 2822 25178
rect 2856 25144 2890 25178
rect 2924 25144 2958 25178
rect 2992 25144 3026 25178
rect 3060 25144 3094 25178
rect 3128 25144 3162 25178
rect 3196 25144 3230 25178
rect 3264 25144 3298 25178
rect 3332 25144 3366 25178
rect 3400 25144 3434 25178
rect 3468 25144 3502 25178
rect 3536 25144 3570 25178
rect 3604 25144 3638 25178
rect 3672 25144 3706 25178
rect 3740 25144 3774 25178
rect 3808 25144 3842 25178
rect 3876 25144 3910 25178
rect 3944 25144 3978 25178
rect 4012 25144 4046 25178
rect 4080 25144 4114 25178
rect 4148 25144 4182 25178
rect 4216 25144 4250 25178
rect 4284 25144 4318 25178
rect 4352 25144 4386 25178
rect 4420 25144 4454 25178
rect 4488 25144 4522 25178
rect 4556 25144 4590 25178
rect 4624 25144 4658 25178
rect 4692 25144 4726 25178
rect 4760 25144 4794 25178
rect 4828 25144 4862 25178
rect 4896 25144 4930 25178
rect 4964 25144 4998 25178
rect 5032 25144 5066 25178
rect 5100 25144 5134 25178
rect 5168 25144 5202 25178
rect 5236 25144 5270 25178
rect 5304 25144 5338 25178
rect 5372 25144 5406 25178
rect 5440 25144 5474 25178
rect 5508 25144 5542 25178
rect 5576 25144 5610 25178
rect 5644 25144 5678 25178
rect 5712 25144 5746 25178
rect 5780 25144 5814 25178
rect 5848 25144 5882 25178
rect 5916 25144 5950 25178
rect 5984 25144 6018 25178
rect 6052 25144 6086 25178
rect 6120 25144 6154 25178
rect 6188 25144 6222 25178
rect 6256 25144 6290 25178
rect 6324 25144 6358 25178
rect 6392 25144 6426 25178
rect 6460 25144 6494 25178
rect 6528 25144 6562 25178
rect 6596 25144 6630 25178
rect 6664 25144 6698 25178
rect 6732 25144 6766 25178
rect 6800 25144 6834 25178
rect 6868 25144 6902 25178
rect 6936 25144 6970 25178
rect 7004 25144 7038 25178
rect 7072 25144 7106 25178
rect 7140 25144 7174 25178
rect 7208 25144 7242 25178
rect 7276 25144 7310 25178
rect 7344 25144 7378 25178
rect 7412 25144 7446 25178
rect 7480 25144 7514 25178
rect 7548 25144 7582 25178
rect 7616 25144 7650 25178
rect 7684 25144 7718 25178
rect 7752 25144 7786 25178
rect 7820 25144 7854 25178
rect 7888 25144 7922 25178
rect 7956 25144 7990 25178
rect 8024 25144 8058 25178
rect 8092 25144 8126 25178
rect 8160 25144 8194 25178
rect 8228 25144 8262 25178
rect 8296 25144 8330 25178
rect 8364 25144 8398 25178
rect 8432 25144 8466 25178
rect 8500 25144 8534 25178
rect 8568 25144 8602 25178
rect 8636 25144 8670 25178
rect 8704 25144 8738 25178
rect 8772 25144 8806 25178
rect 8840 25144 8874 25178
rect 8908 25144 8942 25178
rect 8976 25144 9010 25178
rect 9044 25144 9078 25178
rect 9112 25144 9146 25178
rect 9180 25144 9214 25178
rect 9248 25144 9282 25178
rect 9316 25144 9350 25178
rect 9384 25144 9418 25178
rect 9452 25144 9486 25178
rect 9520 25144 9554 25178
rect 9588 25144 9622 25178
rect 9656 25144 9690 25178
rect 9724 25144 9758 25178
rect 9792 25144 9826 25178
rect 9860 25144 9894 25178
rect 9928 25144 9962 25178
rect 9996 25144 10030 25178
rect 10064 25144 10098 25178
rect 10132 25144 10166 25178
rect 10200 25144 10234 25178
rect 10268 25144 10302 25178
rect 10336 25144 10370 25178
rect 10404 25144 10438 25178
rect 10472 25144 10506 25178
rect 10540 25144 10574 25178
rect 10608 25144 10642 25178
rect 10676 25144 10710 25178
rect 10744 25144 10778 25178
rect 10812 25144 10846 25178
rect 10880 25144 10914 25178
rect 10948 25144 10982 25178
rect 11016 25144 11050 25178
rect 11084 25144 11118 25178
rect 11152 25144 11186 25178
rect 11220 25144 11254 25178
rect 11288 25144 11322 25178
rect 11356 25144 11390 25178
rect 11424 25144 11458 25178
rect 11492 25144 11526 25178
rect 11560 25144 11594 25178
rect 11628 25144 11662 25178
rect 11696 25144 11730 25178
rect 11764 25144 11798 25178
rect 11832 25144 11866 25178
rect 11900 25144 11934 25178
rect 11968 25144 12002 25178
rect 12036 25144 12070 25178
rect 12104 25144 12138 25178
rect 12172 25144 12206 25178
rect 12240 25144 12274 25178
rect 12308 25144 12342 25178
rect 12376 25144 12410 25178
rect 12444 25144 12478 25178
rect 12512 25144 12546 25178
rect 12580 25144 12614 25178
rect 12648 25144 12682 25178
rect 12716 25144 12750 25178
rect 12784 25144 12818 25178
rect 12852 25144 12886 25178
rect 12920 25144 12954 25178
rect 12988 25144 13022 25178
rect 13056 25144 13090 25178
rect 13124 25144 13158 25178
rect 13192 25144 13226 25178
rect 13260 25144 13294 25178
rect 13328 25144 13362 25178
rect 13396 25144 13430 25178
rect 13464 25144 13498 25178
rect 13532 25144 13566 25178
rect 13600 25144 13634 25178
rect 13668 25144 13702 25178
rect 13736 25144 13770 25178
rect 13804 25144 13838 25178
rect 13872 25144 13906 25178
rect 13940 25144 13974 25178
rect 14008 25144 14042 25178
rect 14076 25144 14110 25178
rect 14144 25144 14178 25178
rect 14212 25144 14246 25178
rect 14280 25144 14314 25178
rect 14348 25144 14382 25178
rect 14416 25144 14450 25178
rect 14484 25144 14518 25178
rect 14552 25144 14586 25178
rect 14620 25144 14654 25178
rect 14688 25144 14722 25178
rect 14756 25144 14790 25178
rect 14824 25144 14858 25178
rect 124 25072 158 25106
rect 193 25072 227 25106
rect 262 25072 296 25106
rect 331 25072 365 25106
rect 400 25072 434 25106
rect 469 25072 503 25106
rect 538 25072 572 25106
rect 607 25072 641 25106
rect 676 25072 710 25106
rect 745 25072 779 25106
rect 814 25072 848 25106
rect 883 25072 917 25106
rect 952 25072 986 25106
rect 1020 25072 1054 25106
rect 1088 25072 1122 25106
rect 1156 25072 1190 25106
rect 1224 25072 1258 25106
rect 1292 25072 1326 25106
rect 1360 25072 1394 25106
rect 1428 25072 1462 25106
rect 1496 25072 1530 25106
rect 1564 25072 1598 25106
rect 1632 25072 1666 25106
rect 1700 25072 1734 25106
rect 1768 25072 1802 25106
rect 1836 25072 1870 25106
rect 1904 25072 1938 25106
rect 1972 25072 2006 25106
rect 2040 25072 2074 25106
rect 2108 25072 2142 25106
rect 2176 25072 2210 25106
rect 2244 25072 2278 25106
rect 2312 25072 2346 25106
rect 2380 25072 2414 25106
rect 2448 25072 2482 25106
rect 2516 25072 2550 25106
rect 2584 25072 2618 25106
rect 2652 25072 2686 25106
rect 2720 25072 2754 25106
rect 2788 25072 2822 25106
rect 2856 25072 2890 25106
rect 2924 25072 2958 25106
rect 2992 25072 3026 25106
rect 3060 25072 3094 25106
rect 3128 25072 3162 25106
rect 3196 25072 3230 25106
rect 3264 25072 3298 25106
rect 3332 25072 3366 25106
rect 3400 25072 3434 25106
rect 3468 25072 3502 25106
rect 3536 25072 3570 25106
rect 3604 25072 3638 25106
rect 3672 25072 3706 25106
rect 3740 25072 3774 25106
rect 3808 25072 3842 25106
rect 3876 25072 3910 25106
rect 3944 25072 3978 25106
rect 4012 25072 4046 25106
rect 4080 25072 4114 25106
rect 4148 25072 4182 25106
rect 4216 25072 4250 25106
rect 4284 25072 4318 25106
rect 4352 25072 4386 25106
rect 4420 25072 4454 25106
rect 4488 25072 4522 25106
rect 4556 25072 4590 25106
rect 4624 25072 4658 25106
rect 4692 25072 4726 25106
rect 4760 25072 4794 25106
rect 4828 25072 4862 25106
rect 4896 25072 4930 25106
rect 4964 25072 4998 25106
rect 5032 25072 5066 25106
rect 5100 25072 5134 25106
rect 5168 25072 5202 25106
rect 5236 25072 5270 25106
rect 5304 25072 5338 25106
rect 5372 25072 5406 25106
rect 5440 25072 5474 25106
rect 5508 25072 5542 25106
rect 5576 25072 5610 25106
rect 5644 25072 5678 25106
rect 5712 25072 5746 25106
rect 5780 25072 5814 25106
rect 5848 25072 5882 25106
rect 5916 25072 5950 25106
rect 5984 25072 6018 25106
rect 6052 25072 6086 25106
rect 6120 25072 6154 25106
rect 6188 25072 6222 25106
rect 6256 25072 6290 25106
rect 6324 25072 6358 25106
rect 6392 25072 6426 25106
rect 6460 25072 6494 25106
rect 6528 25072 6562 25106
rect 6596 25072 6630 25106
rect 6664 25072 6698 25106
rect 6732 25072 6766 25106
rect 6800 25072 6834 25106
rect 6868 25072 6902 25106
rect 6936 25072 6970 25106
rect 7004 25072 7038 25106
rect 7072 25072 7106 25106
rect 7140 25072 7174 25106
rect 7208 25072 7242 25106
rect 7276 25072 7310 25106
rect 7344 25072 7378 25106
rect 7412 25072 7446 25106
rect 7480 25072 7514 25106
rect 7548 25072 7582 25106
rect 7616 25072 7650 25106
rect 7684 25072 7718 25106
rect 7752 25072 7786 25106
rect 7820 25072 7854 25106
rect 7888 25072 7922 25106
rect 7956 25072 7990 25106
rect 8024 25072 8058 25106
rect 8092 25072 8126 25106
rect 8160 25072 8194 25106
rect 8228 25072 8262 25106
rect 8296 25072 8330 25106
rect 8364 25072 8398 25106
rect 8432 25072 8466 25106
rect 8500 25072 8534 25106
rect 8568 25072 8602 25106
rect 8636 25072 8670 25106
rect 8704 25072 8738 25106
rect 8772 25072 8806 25106
rect 8840 25072 8874 25106
rect 8908 25072 8942 25106
rect 8976 25072 9010 25106
rect 9044 25072 9078 25106
rect 9112 25072 9146 25106
rect 9180 25072 9214 25106
rect 9248 25072 9282 25106
rect 9316 25072 9350 25106
rect 9384 25072 9418 25106
rect 9452 25072 9486 25106
rect 9520 25072 9554 25106
rect 9588 25072 9622 25106
rect 9656 25072 9690 25106
rect 9724 25072 9758 25106
rect 9792 25072 9826 25106
rect 9860 25072 9894 25106
rect 9928 25072 9962 25106
rect 9996 25072 10030 25106
rect 10064 25072 10098 25106
rect 10132 25072 10166 25106
rect 10200 25072 10234 25106
rect 10268 25072 10302 25106
rect 10336 25072 10370 25106
rect 10404 25072 10438 25106
rect 10472 25072 10506 25106
rect 10540 25072 10574 25106
rect 10608 25072 10642 25106
rect 10676 25072 10710 25106
rect 10744 25072 10778 25106
rect 10812 25072 10846 25106
rect 10880 25072 10914 25106
rect 10948 25072 10982 25106
rect 11016 25072 11050 25106
rect 11084 25072 11118 25106
rect 11152 25072 11186 25106
rect 11220 25072 11254 25106
rect 11288 25072 11322 25106
rect 11356 25072 11390 25106
rect 11424 25072 11458 25106
rect 11492 25072 11526 25106
rect 11560 25072 11594 25106
rect 11628 25072 11662 25106
rect 11696 25072 11730 25106
rect 11764 25072 11798 25106
rect 11832 25072 11866 25106
rect 11900 25072 11934 25106
rect 11968 25072 12002 25106
rect 12036 25072 12070 25106
rect 12104 25072 12138 25106
rect 12172 25072 12206 25106
rect 12240 25072 12274 25106
rect 12308 25072 12342 25106
rect 12376 25072 12410 25106
rect 12444 25072 12478 25106
rect 12512 25072 12546 25106
rect 12580 25072 12614 25106
rect 12648 25072 12682 25106
rect 12716 25072 12750 25106
rect 12784 25072 12818 25106
rect 12852 25072 12886 25106
rect 12920 25072 12954 25106
rect 12988 25072 13022 25106
rect 13056 25072 13090 25106
rect 13124 25072 13158 25106
rect 13192 25072 13226 25106
rect 13260 25072 13294 25106
rect 13328 25072 13362 25106
rect 13396 25072 13430 25106
rect 13464 25072 13498 25106
rect 13532 25072 13566 25106
rect 13600 25072 13634 25106
rect 13668 25072 13702 25106
rect 13736 25072 13770 25106
rect 13804 25072 13838 25106
rect 13872 25072 13906 25106
rect 13940 25072 13974 25106
rect 14008 25072 14042 25106
rect 14076 25072 14110 25106
rect 14144 25072 14178 25106
rect 14212 25072 14246 25106
rect 14280 25072 14314 25106
rect 14348 25072 14382 25106
rect 14416 25072 14450 25106
rect 14484 25072 14518 25106
rect 14552 25072 14586 25106
rect 14620 25072 14654 25106
rect 14688 25072 14722 25106
rect 14756 25072 14790 25106
rect 14824 25072 14858 25106
rect 124 25000 158 25034
rect 193 25000 227 25034
rect 262 25000 296 25034
rect 331 25000 365 25034
rect 400 25000 434 25034
rect 469 25000 503 25034
rect 538 25000 572 25034
rect 607 25000 641 25034
rect 676 25000 710 25034
rect 745 25000 779 25034
rect 814 25000 848 25034
rect 883 25000 917 25034
rect 952 25000 986 25034
rect 1020 25000 1054 25034
rect 1088 25000 1122 25034
rect 1156 25000 1190 25034
rect 1224 25000 1258 25034
rect 1292 25000 1326 25034
rect 1360 25000 1394 25034
rect 1428 25000 1462 25034
rect 1496 25000 1530 25034
rect 1564 25000 1598 25034
rect 1632 25000 1666 25034
rect 1700 25000 1734 25034
rect 1768 25000 1802 25034
rect 1836 25000 1870 25034
rect 1904 25000 1938 25034
rect 1972 25000 2006 25034
rect 2040 25000 2074 25034
rect 2108 25000 2142 25034
rect 2176 25000 2210 25034
rect 2244 25000 2278 25034
rect 2312 25000 2346 25034
rect 2380 25000 2414 25034
rect 2448 25000 2482 25034
rect 2516 25000 2550 25034
rect 2584 25000 2618 25034
rect 2652 25000 2686 25034
rect 2720 25000 2754 25034
rect 2788 25000 2822 25034
rect 2856 25000 2890 25034
rect 2924 25000 2958 25034
rect 2992 25000 3026 25034
rect 3060 25000 3094 25034
rect 3128 25000 3162 25034
rect 3196 25000 3230 25034
rect 3264 25000 3298 25034
rect 3332 25000 3366 25034
rect 3400 25000 3434 25034
rect 3468 25000 3502 25034
rect 3536 25000 3570 25034
rect 3604 25000 3638 25034
rect 3672 25000 3706 25034
rect 3740 25000 3774 25034
rect 3808 25000 3842 25034
rect 3876 25000 3910 25034
rect 3944 25000 3978 25034
rect 4012 25000 4046 25034
rect 4080 25000 4114 25034
rect 4148 25000 4182 25034
rect 4216 25000 4250 25034
rect 4284 25000 4318 25034
rect 4352 25000 4386 25034
rect 4420 25000 4454 25034
rect 4488 25000 4522 25034
rect 4556 25000 4590 25034
rect 4624 25000 4658 25034
rect 4692 25000 4726 25034
rect 4760 25000 4794 25034
rect 4828 25000 4862 25034
rect 4896 25000 4930 25034
rect 4964 25000 4998 25034
rect 5032 25000 5066 25034
rect 5100 25000 5134 25034
rect 5168 25000 5202 25034
rect 5236 25000 5270 25034
rect 5304 25000 5338 25034
rect 5372 25000 5406 25034
rect 5440 25000 5474 25034
rect 5508 25000 5542 25034
rect 5576 25000 5610 25034
rect 5644 25000 5678 25034
rect 5712 25000 5746 25034
rect 5780 25000 5814 25034
rect 5848 25000 5882 25034
rect 5916 25000 5950 25034
rect 5984 25000 6018 25034
rect 6052 25000 6086 25034
rect 6120 25000 6154 25034
rect 6188 25000 6222 25034
rect 6256 25000 6290 25034
rect 6324 25000 6358 25034
rect 6392 25000 6426 25034
rect 6460 25000 6494 25034
rect 6528 25000 6562 25034
rect 6596 25000 6630 25034
rect 6664 25000 6698 25034
rect 6732 25000 6766 25034
rect 6800 25000 6834 25034
rect 6868 25000 6902 25034
rect 6936 25000 6970 25034
rect 7004 25000 7038 25034
rect 7072 25000 7106 25034
rect 7140 25000 7174 25034
rect 7208 25000 7242 25034
rect 7276 25000 7310 25034
rect 7344 25000 7378 25034
rect 7412 25000 7446 25034
rect 7480 25000 7514 25034
rect 7548 25000 7582 25034
rect 7616 25000 7650 25034
rect 7684 25000 7718 25034
rect 7752 25000 7786 25034
rect 7820 25000 7854 25034
rect 7888 25000 7922 25034
rect 7956 25000 7990 25034
rect 8024 25000 8058 25034
rect 8092 25000 8126 25034
rect 8160 25000 8194 25034
rect 8228 25000 8262 25034
rect 8296 25000 8330 25034
rect 8364 25000 8398 25034
rect 8432 25000 8466 25034
rect 8500 25000 8534 25034
rect 8568 25000 8602 25034
rect 8636 25000 8670 25034
rect 8704 25000 8738 25034
rect 8772 25000 8806 25034
rect 8840 25000 8874 25034
rect 8908 25000 8942 25034
rect 8976 25000 9010 25034
rect 9044 25000 9078 25034
rect 9112 25000 9146 25034
rect 9180 25000 9214 25034
rect 9248 25000 9282 25034
rect 9316 25000 9350 25034
rect 9384 25000 9418 25034
rect 9452 25000 9486 25034
rect 9520 25000 9554 25034
rect 9588 25000 9622 25034
rect 9656 25000 9690 25034
rect 9724 25000 9758 25034
rect 9792 25000 9826 25034
rect 9860 25000 9894 25034
rect 9928 25000 9962 25034
rect 9996 25000 10030 25034
rect 10064 25000 10098 25034
rect 10132 25000 10166 25034
rect 10200 25000 10234 25034
rect 10268 25000 10302 25034
rect 10336 25000 10370 25034
rect 10404 25000 10438 25034
rect 10472 25000 10506 25034
rect 10540 25000 10574 25034
rect 10608 25000 10642 25034
rect 10676 25000 10710 25034
rect 10744 25000 10778 25034
rect 10812 25000 10846 25034
rect 10880 25000 10914 25034
rect 10948 25000 10982 25034
rect 11016 25000 11050 25034
rect 11084 25000 11118 25034
rect 11152 25000 11186 25034
rect 11220 25000 11254 25034
rect 11288 25000 11322 25034
rect 11356 25000 11390 25034
rect 11424 25000 11458 25034
rect 11492 25000 11526 25034
rect 11560 25000 11594 25034
rect 11628 25000 11662 25034
rect 11696 25000 11730 25034
rect 11764 25000 11798 25034
rect 11832 25000 11866 25034
rect 11900 25000 11934 25034
rect 11968 25000 12002 25034
rect 12036 25000 12070 25034
rect 12104 25000 12138 25034
rect 12172 25000 12206 25034
rect 12240 25000 12274 25034
rect 12308 25000 12342 25034
rect 12376 25000 12410 25034
rect 12444 25000 12478 25034
rect 12512 25000 12546 25034
rect 12580 25000 12614 25034
rect 12648 25000 12682 25034
rect 12716 25000 12750 25034
rect 12784 25000 12818 25034
rect 12852 25000 12886 25034
rect 12920 25000 12954 25034
rect 12988 25000 13022 25034
rect 13056 25000 13090 25034
rect 13124 25000 13158 25034
rect 13192 25000 13226 25034
rect 13260 25000 13294 25034
rect 13328 25000 13362 25034
rect 13396 25000 13430 25034
rect 13464 25000 13498 25034
rect 13532 25000 13566 25034
rect 13600 25000 13634 25034
rect 13668 25000 13702 25034
rect 13736 25000 13770 25034
rect 13804 25000 13838 25034
rect 13872 25000 13906 25034
rect 13940 25000 13974 25034
rect 14008 25000 14042 25034
rect 14076 25000 14110 25034
rect 14144 25000 14178 25034
rect 14212 25000 14246 25034
rect 14280 25000 14314 25034
rect 14348 25000 14382 25034
rect 14416 25000 14450 25034
rect 14484 25000 14518 25034
rect 14552 25000 14586 25034
rect 14620 25000 14654 25034
rect 14688 25000 14722 25034
rect 14756 25000 14790 25034
rect 14824 25000 14858 25034
rect 124 24928 158 24962
rect 193 24928 227 24962
rect 262 24928 296 24962
rect 331 24928 365 24962
rect 400 24928 434 24962
rect 469 24928 503 24962
rect 538 24928 572 24962
rect 607 24928 641 24962
rect 676 24928 710 24962
rect 745 24928 779 24962
rect 814 24928 848 24962
rect 883 24928 917 24962
rect 952 24928 986 24962
rect 1020 24928 1054 24962
rect 1088 24928 1122 24962
rect 1156 24928 1190 24962
rect 1224 24928 1258 24962
rect 1292 24928 1326 24962
rect 1360 24928 1394 24962
rect 1428 24928 1462 24962
rect 1496 24928 1530 24962
rect 1564 24928 1598 24962
rect 1632 24928 1666 24962
rect 1700 24928 1734 24962
rect 1768 24928 1802 24962
rect 1836 24928 1870 24962
rect 1904 24928 1938 24962
rect 1972 24928 2006 24962
rect 2040 24928 2074 24962
rect 2108 24928 2142 24962
rect 2176 24928 2210 24962
rect 2244 24928 2278 24962
rect 2312 24928 2346 24962
rect 2380 24928 2414 24962
rect 2448 24928 2482 24962
rect 2516 24928 2550 24962
rect 2584 24928 2618 24962
rect 2652 24928 2686 24962
rect 2720 24928 2754 24962
rect 2788 24928 2822 24962
rect 2856 24928 2890 24962
rect 2924 24928 2958 24962
rect 2992 24928 3026 24962
rect 3060 24928 3094 24962
rect 3128 24928 3162 24962
rect 3196 24928 3230 24962
rect 3264 24928 3298 24962
rect 3332 24928 3366 24962
rect 3400 24928 3434 24962
rect 3468 24928 3502 24962
rect 3536 24928 3570 24962
rect 3604 24928 3638 24962
rect 3672 24928 3706 24962
rect 3740 24928 3774 24962
rect 3808 24928 3842 24962
rect 3876 24928 3910 24962
rect 3944 24928 3978 24962
rect 4012 24928 4046 24962
rect 4080 24928 4114 24962
rect 4148 24928 4182 24962
rect 4216 24928 4250 24962
rect 4284 24928 4318 24962
rect 4352 24928 4386 24962
rect 4420 24928 4454 24962
rect 4488 24928 4522 24962
rect 4556 24928 4590 24962
rect 4624 24928 4658 24962
rect 4692 24928 4726 24962
rect 4760 24928 4794 24962
rect 4828 24928 4862 24962
rect 4896 24928 4930 24962
rect 4964 24928 4998 24962
rect 5032 24928 5066 24962
rect 5100 24928 5134 24962
rect 5168 24928 5202 24962
rect 5236 24928 5270 24962
rect 5304 24928 5338 24962
rect 5372 24928 5406 24962
rect 5440 24928 5474 24962
rect 5508 24928 5542 24962
rect 5576 24928 5610 24962
rect 5644 24928 5678 24962
rect 5712 24928 5746 24962
rect 5780 24928 5814 24962
rect 5848 24928 5882 24962
rect 5916 24928 5950 24962
rect 5984 24928 6018 24962
rect 6052 24928 6086 24962
rect 6120 24928 6154 24962
rect 6188 24928 6222 24962
rect 6256 24928 6290 24962
rect 6324 24928 6358 24962
rect 6392 24928 6426 24962
rect 6460 24928 6494 24962
rect 6528 24928 6562 24962
rect 6596 24928 6630 24962
rect 6664 24928 6698 24962
rect 6732 24928 6766 24962
rect 6800 24928 6834 24962
rect 6868 24928 6902 24962
rect 6936 24928 6970 24962
rect 7004 24928 7038 24962
rect 7072 24928 7106 24962
rect 7140 24928 7174 24962
rect 7208 24928 7242 24962
rect 7276 24928 7310 24962
rect 7344 24928 7378 24962
rect 7412 24928 7446 24962
rect 7480 24928 7514 24962
rect 7548 24928 7582 24962
rect 7616 24928 7650 24962
rect 7684 24928 7718 24962
rect 7752 24928 7786 24962
rect 7820 24928 7854 24962
rect 7888 24928 7922 24962
rect 7956 24928 7990 24962
rect 8024 24928 8058 24962
rect 8092 24928 8126 24962
rect 8160 24928 8194 24962
rect 8228 24928 8262 24962
rect 8296 24928 8330 24962
rect 8364 24928 8398 24962
rect 8432 24928 8466 24962
rect 8500 24928 8534 24962
rect 8568 24928 8602 24962
rect 8636 24928 8670 24962
rect 8704 24928 8738 24962
rect 8772 24928 8806 24962
rect 8840 24928 8874 24962
rect 8908 24928 8942 24962
rect 8976 24928 9010 24962
rect 9044 24928 9078 24962
rect 9112 24928 9146 24962
rect 9180 24928 9214 24962
rect 9248 24928 9282 24962
rect 9316 24928 9350 24962
rect 9384 24928 9418 24962
rect 9452 24928 9486 24962
rect 9520 24928 9554 24962
rect 9588 24928 9622 24962
rect 9656 24928 9690 24962
rect 9724 24928 9758 24962
rect 9792 24928 9826 24962
rect 9860 24928 9894 24962
rect 9928 24928 9962 24962
rect 9996 24928 10030 24962
rect 10064 24928 10098 24962
rect 10132 24928 10166 24962
rect 10200 24928 10234 24962
rect 10268 24928 10302 24962
rect 10336 24928 10370 24962
rect 10404 24928 10438 24962
rect 10472 24928 10506 24962
rect 10540 24928 10574 24962
rect 10608 24928 10642 24962
rect 10676 24928 10710 24962
rect 10744 24928 10778 24962
rect 10812 24928 10846 24962
rect 10880 24928 10914 24962
rect 10948 24928 10982 24962
rect 11016 24928 11050 24962
rect 11084 24928 11118 24962
rect 11152 24928 11186 24962
rect 11220 24928 11254 24962
rect 11288 24928 11322 24962
rect 11356 24928 11390 24962
rect 11424 24928 11458 24962
rect 11492 24928 11526 24962
rect 11560 24928 11594 24962
rect 11628 24928 11662 24962
rect 11696 24928 11730 24962
rect 11764 24928 11798 24962
rect 11832 24928 11866 24962
rect 11900 24928 11934 24962
rect 11968 24928 12002 24962
rect 12036 24928 12070 24962
rect 12104 24928 12138 24962
rect 12172 24928 12206 24962
rect 12240 24928 12274 24962
rect 12308 24928 12342 24962
rect 12376 24928 12410 24962
rect 12444 24928 12478 24962
rect 12512 24928 12546 24962
rect 12580 24928 12614 24962
rect 12648 24928 12682 24962
rect 12716 24928 12750 24962
rect 12784 24928 12818 24962
rect 12852 24928 12886 24962
rect 12920 24928 12954 24962
rect 12988 24928 13022 24962
rect 13056 24928 13090 24962
rect 13124 24928 13158 24962
rect 13192 24928 13226 24962
rect 13260 24928 13294 24962
rect 13328 24928 13362 24962
rect 13396 24928 13430 24962
rect 13464 24928 13498 24962
rect 13532 24928 13566 24962
rect 13600 24928 13634 24962
rect 13668 24928 13702 24962
rect 13736 24928 13770 24962
rect 13804 24928 13838 24962
rect 13872 24928 13906 24962
rect 13940 24928 13974 24962
rect 14008 24928 14042 24962
rect 14076 24928 14110 24962
rect 14144 24928 14178 24962
rect 14212 24928 14246 24962
rect 14280 24928 14314 24962
rect 14348 24928 14382 24962
rect 14416 24928 14450 24962
rect 14484 24928 14518 24962
rect 14552 24928 14586 24962
rect 14620 24928 14654 24962
rect 14688 24928 14722 24962
rect 14756 24928 14790 24962
rect 14824 24928 14858 24962
rect 124 24856 158 24890
rect 193 24856 227 24890
rect 262 24856 296 24890
rect 331 24856 365 24890
rect 400 24856 434 24890
rect 469 24856 503 24890
rect 538 24856 572 24890
rect 607 24856 641 24890
rect 676 24856 710 24890
rect 745 24856 779 24890
rect 814 24856 848 24890
rect 883 24856 917 24890
rect 952 24856 986 24890
rect 1020 24856 1054 24890
rect 1088 24856 1122 24890
rect 1156 24856 1190 24890
rect 1224 24856 1258 24890
rect 1292 24856 1326 24890
rect 1360 24856 1394 24890
rect 1428 24856 1462 24890
rect 1496 24856 1530 24890
rect 1564 24856 1598 24890
rect 1632 24856 1666 24890
rect 1700 24856 1734 24890
rect 1768 24856 1802 24890
rect 1836 24856 1870 24890
rect 1904 24856 1938 24890
rect 1972 24856 2006 24890
rect 2040 24856 2074 24890
rect 2108 24856 2142 24890
rect 2176 24856 2210 24890
rect 2244 24856 2278 24890
rect 2312 24856 2346 24890
rect 2380 24856 2414 24890
rect 2448 24856 2482 24890
rect 2516 24856 2550 24890
rect 2584 24856 2618 24890
rect 2652 24856 2686 24890
rect 2720 24856 2754 24890
rect 2788 24856 2822 24890
rect 2856 24856 2890 24890
rect 2924 24856 2958 24890
rect 2992 24856 3026 24890
rect 3060 24856 3094 24890
rect 3128 24856 3162 24890
rect 3196 24856 3230 24890
rect 3264 24856 3298 24890
rect 3332 24856 3366 24890
rect 3400 24856 3434 24890
rect 3468 24856 3502 24890
rect 3536 24856 3570 24890
rect 3604 24856 3638 24890
rect 3672 24856 3706 24890
rect 3740 24856 3774 24890
rect 3808 24856 3842 24890
rect 3876 24856 3910 24890
rect 3944 24856 3978 24890
rect 4012 24856 4046 24890
rect 4080 24856 4114 24890
rect 4148 24856 4182 24890
rect 4216 24856 4250 24890
rect 4284 24856 4318 24890
rect 4352 24856 4386 24890
rect 4420 24856 4454 24890
rect 4488 24856 4522 24890
rect 4556 24856 4590 24890
rect 4624 24856 4658 24890
rect 4692 24856 4726 24890
rect 4760 24856 4794 24890
rect 4828 24856 4862 24890
rect 4896 24856 4930 24890
rect 4964 24856 4998 24890
rect 5032 24856 5066 24890
rect 5100 24856 5134 24890
rect 5168 24856 5202 24890
rect 5236 24856 5270 24890
rect 5304 24856 5338 24890
rect 5372 24856 5406 24890
rect 5440 24856 5474 24890
rect 5508 24856 5542 24890
rect 5576 24856 5610 24890
rect 5644 24856 5678 24890
rect 5712 24856 5746 24890
rect 5780 24856 5814 24890
rect 5848 24856 5882 24890
rect 5916 24856 5950 24890
rect 5984 24856 6018 24890
rect 6052 24856 6086 24890
rect 6120 24856 6154 24890
rect 6188 24856 6222 24890
rect 6256 24856 6290 24890
rect 6324 24856 6358 24890
rect 6392 24856 6426 24890
rect 6460 24856 6494 24890
rect 6528 24856 6562 24890
rect 6596 24856 6630 24890
rect 6664 24856 6698 24890
rect 6732 24856 6766 24890
rect 6800 24856 6834 24890
rect 6868 24856 6902 24890
rect 6936 24856 6970 24890
rect 7004 24856 7038 24890
rect 7072 24856 7106 24890
rect 7140 24856 7174 24890
rect 7208 24856 7242 24890
rect 7276 24856 7310 24890
rect 7344 24856 7378 24890
rect 7412 24856 7446 24890
rect 7480 24856 7514 24890
rect 7548 24856 7582 24890
rect 7616 24856 7650 24890
rect 7684 24856 7718 24890
rect 7752 24856 7786 24890
rect 7820 24856 7854 24890
rect 7888 24856 7922 24890
rect 7956 24856 7990 24890
rect 8024 24856 8058 24890
rect 8092 24856 8126 24890
rect 8160 24856 8194 24890
rect 8228 24856 8262 24890
rect 8296 24856 8330 24890
rect 8364 24856 8398 24890
rect 8432 24856 8466 24890
rect 8500 24856 8534 24890
rect 8568 24856 8602 24890
rect 8636 24856 8670 24890
rect 8704 24856 8738 24890
rect 8772 24856 8806 24890
rect 8840 24856 8874 24890
rect 8908 24856 8942 24890
rect 8976 24856 9010 24890
rect 9044 24856 9078 24890
rect 9112 24856 9146 24890
rect 9180 24856 9214 24890
rect 9248 24856 9282 24890
rect 9316 24856 9350 24890
rect 9384 24856 9418 24890
rect 9452 24856 9486 24890
rect 9520 24856 9554 24890
rect 9588 24856 9622 24890
rect 9656 24856 9690 24890
rect 9724 24856 9758 24890
rect 9792 24856 9826 24890
rect 9860 24856 9894 24890
rect 9928 24856 9962 24890
rect 9996 24856 10030 24890
rect 10064 24856 10098 24890
rect 10132 24856 10166 24890
rect 10200 24856 10234 24890
rect 10268 24856 10302 24890
rect 10336 24856 10370 24890
rect 10404 24856 10438 24890
rect 10472 24856 10506 24890
rect 10540 24856 10574 24890
rect 10608 24856 10642 24890
rect 10676 24856 10710 24890
rect 10744 24856 10778 24890
rect 10812 24856 10846 24890
rect 10880 24856 10914 24890
rect 10948 24856 10982 24890
rect 11016 24856 11050 24890
rect 11084 24856 11118 24890
rect 11152 24856 11186 24890
rect 11220 24856 11254 24890
rect 11288 24856 11322 24890
rect 11356 24856 11390 24890
rect 11424 24856 11458 24890
rect 11492 24856 11526 24890
rect 11560 24856 11594 24890
rect 11628 24856 11662 24890
rect 11696 24856 11730 24890
rect 11764 24856 11798 24890
rect 11832 24856 11866 24890
rect 11900 24856 11934 24890
rect 11968 24856 12002 24890
rect 12036 24856 12070 24890
rect 12104 24856 12138 24890
rect 12172 24856 12206 24890
rect 12240 24856 12274 24890
rect 12308 24856 12342 24890
rect 12376 24856 12410 24890
rect 12444 24856 12478 24890
rect 12512 24856 12546 24890
rect 12580 24856 12614 24890
rect 12648 24856 12682 24890
rect 12716 24856 12750 24890
rect 12784 24856 12818 24890
rect 12852 24856 12886 24890
rect 12920 24856 12954 24890
rect 12988 24856 13022 24890
rect 13056 24856 13090 24890
rect 13124 24856 13158 24890
rect 13192 24856 13226 24890
rect 13260 24856 13294 24890
rect 13328 24856 13362 24890
rect 13396 24856 13430 24890
rect 13464 24856 13498 24890
rect 13532 24856 13566 24890
rect 13600 24856 13634 24890
rect 13668 24856 13702 24890
rect 13736 24856 13770 24890
rect 13804 24856 13838 24890
rect 13872 24856 13906 24890
rect 13940 24856 13974 24890
rect 14008 24856 14042 24890
rect 14076 24856 14110 24890
rect 14144 24856 14178 24890
rect 14212 24856 14246 24890
rect 14280 24856 14314 24890
rect 14348 24856 14382 24890
rect 14416 24856 14450 24890
rect 14484 24856 14518 24890
rect 14552 24856 14586 24890
rect 14620 24856 14654 24890
rect 14688 24856 14722 24890
rect 14756 24856 14790 24890
rect 14824 24856 14858 24890
rect 124 24784 158 24818
rect 193 24784 227 24818
rect 262 24784 296 24818
rect 331 24784 365 24818
rect 400 24784 434 24818
rect 469 24784 503 24818
rect 538 24784 572 24818
rect 607 24784 641 24818
rect 676 24784 710 24818
rect 745 24784 779 24818
rect 814 24784 848 24818
rect 883 24784 917 24818
rect 952 24784 986 24818
rect 1020 24784 1054 24818
rect 1088 24784 1122 24818
rect 1156 24784 1190 24818
rect 1224 24784 1258 24818
rect 1292 24784 1326 24818
rect 1360 24784 1394 24818
rect 1428 24784 1462 24818
rect 1496 24784 1530 24818
rect 1564 24784 1598 24818
rect 1632 24784 1666 24818
rect 1700 24784 1734 24818
rect 1768 24784 1802 24818
rect 1836 24784 1870 24818
rect 1904 24784 1938 24818
rect 1972 24784 2006 24818
rect 2040 24784 2074 24818
rect 2108 24784 2142 24818
rect 2176 24784 2210 24818
rect 2244 24784 2278 24818
rect 2312 24784 2346 24818
rect 2380 24784 2414 24818
rect 2448 24784 2482 24818
rect 2516 24784 2550 24818
rect 2584 24784 2618 24818
rect 2652 24784 2686 24818
rect 2720 24784 2754 24818
rect 2788 24784 2822 24818
rect 2856 24784 2890 24818
rect 2924 24784 2958 24818
rect 2992 24784 3026 24818
rect 3060 24784 3094 24818
rect 3128 24784 3162 24818
rect 3196 24784 3230 24818
rect 3264 24784 3298 24818
rect 3332 24784 3366 24818
rect 3400 24784 3434 24818
rect 3468 24784 3502 24818
rect 3536 24784 3570 24818
rect 3604 24784 3638 24818
rect 3672 24784 3706 24818
rect 3740 24784 3774 24818
rect 3808 24784 3842 24818
rect 3876 24784 3910 24818
rect 3944 24784 3978 24818
rect 4012 24784 4046 24818
rect 4080 24784 4114 24818
rect 4148 24784 4182 24818
rect 4216 24784 4250 24818
rect 4284 24784 4318 24818
rect 4352 24784 4386 24818
rect 4420 24784 4454 24818
rect 4488 24784 4522 24818
rect 4556 24784 4590 24818
rect 4624 24784 4658 24818
rect 4692 24784 4726 24818
rect 4760 24784 4794 24818
rect 4828 24784 4862 24818
rect 4896 24784 4930 24818
rect 4964 24784 4998 24818
rect 5032 24784 5066 24818
rect 5100 24784 5134 24818
rect 5168 24784 5202 24818
rect 5236 24784 5270 24818
rect 5304 24784 5338 24818
rect 5372 24784 5406 24818
rect 5440 24784 5474 24818
rect 5508 24784 5542 24818
rect 5576 24784 5610 24818
rect 5644 24784 5678 24818
rect 5712 24784 5746 24818
rect 5780 24784 5814 24818
rect 5848 24784 5882 24818
rect 5916 24784 5950 24818
rect 5984 24784 6018 24818
rect 6052 24784 6086 24818
rect 6120 24784 6154 24818
rect 6188 24784 6222 24818
rect 6256 24784 6290 24818
rect 6324 24784 6358 24818
rect 6392 24784 6426 24818
rect 6460 24784 6494 24818
rect 6528 24784 6562 24818
rect 6596 24784 6630 24818
rect 6664 24784 6698 24818
rect 6732 24784 6766 24818
rect 6800 24784 6834 24818
rect 6868 24784 6902 24818
rect 6936 24784 6970 24818
rect 7004 24784 7038 24818
rect 7072 24784 7106 24818
rect 7140 24784 7174 24818
rect 7208 24784 7242 24818
rect 7276 24784 7310 24818
rect 7344 24784 7378 24818
rect 7412 24784 7446 24818
rect 7480 24784 7514 24818
rect 7548 24784 7582 24818
rect 7616 24784 7650 24818
rect 7684 24784 7718 24818
rect 7752 24784 7786 24818
rect 7820 24784 7854 24818
rect 7888 24784 7922 24818
rect 7956 24784 7990 24818
rect 8024 24784 8058 24818
rect 8092 24784 8126 24818
rect 8160 24784 8194 24818
rect 8228 24784 8262 24818
rect 8296 24784 8330 24818
rect 8364 24784 8398 24818
rect 8432 24784 8466 24818
rect 8500 24784 8534 24818
rect 8568 24784 8602 24818
rect 8636 24784 8670 24818
rect 8704 24784 8738 24818
rect 8772 24784 8806 24818
rect 8840 24784 8874 24818
rect 8908 24784 8942 24818
rect 8976 24784 9010 24818
rect 9044 24784 9078 24818
rect 9112 24784 9146 24818
rect 9180 24784 9214 24818
rect 9248 24784 9282 24818
rect 9316 24784 9350 24818
rect 9384 24784 9418 24818
rect 9452 24784 9486 24818
rect 9520 24784 9554 24818
rect 9588 24784 9622 24818
rect 9656 24784 9690 24818
rect 9724 24784 9758 24818
rect 9792 24784 9826 24818
rect 9860 24784 9894 24818
rect 9928 24784 9962 24818
rect 9996 24784 10030 24818
rect 10064 24784 10098 24818
rect 10132 24784 10166 24818
rect 10200 24784 10234 24818
rect 10268 24784 10302 24818
rect 10336 24784 10370 24818
rect 10404 24784 10438 24818
rect 10472 24784 10506 24818
rect 10540 24784 10574 24818
rect 10608 24784 10642 24818
rect 10676 24784 10710 24818
rect 10744 24784 10778 24818
rect 10812 24784 10846 24818
rect 10880 24784 10914 24818
rect 10948 24784 10982 24818
rect 11016 24784 11050 24818
rect 11084 24784 11118 24818
rect 11152 24784 11186 24818
rect 11220 24784 11254 24818
rect 11288 24784 11322 24818
rect 11356 24784 11390 24818
rect 11424 24784 11458 24818
rect 11492 24784 11526 24818
rect 11560 24784 11594 24818
rect 11628 24784 11662 24818
rect 11696 24784 11730 24818
rect 11764 24784 11798 24818
rect 11832 24784 11866 24818
rect 11900 24784 11934 24818
rect 11968 24784 12002 24818
rect 12036 24784 12070 24818
rect 12104 24784 12138 24818
rect 12172 24784 12206 24818
rect 12240 24784 12274 24818
rect 12308 24784 12342 24818
rect 12376 24784 12410 24818
rect 12444 24784 12478 24818
rect 12512 24784 12546 24818
rect 12580 24784 12614 24818
rect 12648 24784 12682 24818
rect 12716 24784 12750 24818
rect 12784 24784 12818 24818
rect 12852 24784 12886 24818
rect 12920 24784 12954 24818
rect 12988 24784 13022 24818
rect 13056 24784 13090 24818
rect 13124 24784 13158 24818
rect 13192 24784 13226 24818
rect 13260 24784 13294 24818
rect 13328 24784 13362 24818
rect 13396 24784 13430 24818
rect 13464 24784 13498 24818
rect 13532 24784 13566 24818
rect 13600 24784 13634 24818
rect 13668 24784 13702 24818
rect 13736 24784 13770 24818
rect 13804 24784 13838 24818
rect 13872 24784 13906 24818
rect 13940 24784 13974 24818
rect 14008 24784 14042 24818
rect 14076 24784 14110 24818
rect 14144 24784 14178 24818
rect 14212 24784 14246 24818
rect 14280 24784 14314 24818
rect 14348 24784 14382 24818
rect 14416 24784 14450 24818
rect 14484 24784 14518 24818
rect 14552 24784 14586 24818
rect 14620 24784 14654 24818
rect 14688 24784 14722 24818
rect 14756 24784 14790 24818
rect 14824 24784 14858 24818
rect 124 24712 158 24746
rect 193 24712 227 24746
rect 262 24712 296 24746
rect 331 24712 365 24746
rect 400 24712 434 24746
rect 469 24712 503 24746
rect 538 24712 572 24746
rect 607 24712 641 24746
rect 676 24712 710 24746
rect 745 24712 779 24746
rect 814 24712 848 24746
rect 883 24712 917 24746
rect 952 24712 986 24746
rect 1020 24712 1054 24746
rect 1088 24712 1122 24746
rect 1156 24712 1190 24746
rect 1224 24712 1258 24746
rect 1292 24712 1326 24746
rect 1360 24712 1394 24746
rect 1428 24712 1462 24746
rect 1496 24712 1530 24746
rect 1564 24712 1598 24746
rect 1632 24712 1666 24746
rect 1700 24712 1734 24746
rect 1768 24712 1802 24746
rect 1836 24712 1870 24746
rect 1904 24712 1938 24746
rect 1972 24712 2006 24746
rect 2040 24712 2074 24746
rect 2108 24712 2142 24746
rect 2176 24712 2210 24746
rect 2244 24712 2278 24746
rect 2312 24712 2346 24746
rect 2380 24712 2414 24746
rect 2448 24712 2482 24746
rect 2516 24712 2550 24746
rect 2584 24712 2618 24746
rect 2652 24712 2686 24746
rect 2720 24712 2754 24746
rect 2788 24712 2822 24746
rect 2856 24712 2890 24746
rect 2924 24712 2958 24746
rect 2992 24712 3026 24746
rect 3060 24712 3094 24746
rect 3128 24712 3162 24746
rect 3196 24712 3230 24746
rect 3264 24712 3298 24746
rect 3332 24712 3366 24746
rect 3400 24712 3434 24746
rect 3468 24712 3502 24746
rect 3536 24712 3570 24746
rect 3604 24712 3638 24746
rect 3672 24712 3706 24746
rect 3740 24712 3774 24746
rect 3808 24712 3842 24746
rect 3876 24712 3910 24746
rect 3944 24712 3978 24746
rect 4012 24712 4046 24746
rect 4080 24712 4114 24746
rect 4148 24712 4182 24746
rect 4216 24712 4250 24746
rect 4284 24712 4318 24746
rect 4352 24712 4386 24746
rect 4420 24712 4454 24746
rect 4488 24712 4522 24746
rect 4556 24712 4590 24746
rect 4624 24712 4658 24746
rect 4692 24712 4726 24746
rect 4760 24712 4794 24746
rect 4828 24712 4862 24746
rect 4896 24712 4930 24746
rect 4964 24712 4998 24746
rect 5032 24712 5066 24746
rect 5100 24712 5134 24746
rect 5168 24712 5202 24746
rect 5236 24712 5270 24746
rect 5304 24712 5338 24746
rect 5372 24712 5406 24746
rect 5440 24712 5474 24746
rect 5508 24712 5542 24746
rect 5576 24712 5610 24746
rect 5644 24712 5678 24746
rect 5712 24712 5746 24746
rect 5780 24712 5814 24746
rect 5848 24712 5882 24746
rect 5916 24712 5950 24746
rect 5984 24712 6018 24746
rect 6052 24712 6086 24746
rect 6120 24712 6154 24746
rect 6188 24712 6222 24746
rect 6256 24712 6290 24746
rect 6324 24712 6358 24746
rect 6392 24712 6426 24746
rect 6460 24712 6494 24746
rect 6528 24712 6562 24746
rect 6596 24712 6630 24746
rect 6664 24712 6698 24746
rect 6732 24712 6766 24746
rect 6800 24712 6834 24746
rect 6868 24712 6902 24746
rect 6936 24712 6970 24746
rect 7004 24712 7038 24746
rect 7072 24712 7106 24746
rect 7140 24712 7174 24746
rect 7208 24712 7242 24746
rect 7276 24712 7310 24746
rect 7344 24712 7378 24746
rect 7412 24712 7446 24746
rect 7480 24712 7514 24746
rect 7548 24712 7582 24746
rect 7616 24712 7650 24746
rect 7684 24712 7718 24746
rect 7752 24712 7786 24746
rect 7820 24712 7854 24746
rect 7888 24712 7922 24746
rect 7956 24712 7990 24746
rect 8024 24712 8058 24746
rect 8092 24712 8126 24746
rect 8160 24712 8194 24746
rect 8228 24712 8262 24746
rect 8296 24712 8330 24746
rect 8364 24712 8398 24746
rect 8432 24712 8466 24746
rect 8500 24712 8534 24746
rect 8568 24712 8602 24746
rect 8636 24712 8670 24746
rect 8704 24712 8738 24746
rect 8772 24712 8806 24746
rect 8840 24712 8874 24746
rect 8908 24712 8942 24746
rect 8976 24712 9010 24746
rect 9044 24712 9078 24746
rect 9112 24712 9146 24746
rect 9180 24712 9214 24746
rect 9248 24712 9282 24746
rect 9316 24712 9350 24746
rect 9384 24712 9418 24746
rect 9452 24712 9486 24746
rect 9520 24712 9554 24746
rect 9588 24712 9622 24746
rect 9656 24712 9690 24746
rect 9724 24712 9758 24746
rect 9792 24712 9826 24746
rect 9860 24712 9894 24746
rect 9928 24712 9962 24746
rect 9996 24712 10030 24746
rect 10064 24712 10098 24746
rect 10132 24712 10166 24746
rect 10200 24712 10234 24746
rect 10268 24712 10302 24746
rect 10336 24712 10370 24746
rect 10404 24712 10438 24746
rect 10472 24712 10506 24746
rect 10540 24712 10574 24746
rect 10608 24712 10642 24746
rect 10676 24712 10710 24746
rect 10744 24712 10778 24746
rect 10812 24712 10846 24746
rect 10880 24712 10914 24746
rect 10948 24712 10982 24746
rect 11016 24712 11050 24746
rect 11084 24712 11118 24746
rect 11152 24712 11186 24746
rect 11220 24712 11254 24746
rect 11288 24712 11322 24746
rect 11356 24712 11390 24746
rect 11424 24712 11458 24746
rect 11492 24712 11526 24746
rect 11560 24712 11594 24746
rect 11628 24712 11662 24746
rect 11696 24712 11730 24746
rect 11764 24712 11798 24746
rect 11832 24712 11866 24746
rect 11900 24712 11934 24746
rect 11968 24712 12002 24746
rect 12036 24712 12070 24746
rect 12104 24712 12138 24746
rect 12172 24712 12206 24746
rect 12240 24712 12274 24746
rect 12308 24712 12342 24746
rect 12376 24712 12410 24746
rect 12444 24712 12478 24746
rect 12512 24712 12546 24746
rect 12580 24712 12614 24746
rect 12648 24712 12682 24746
rect 12716 24712 12750 24746
rect 12784 24712 12818 24746
rect 12852 24712 12886 24746
rect 12920 24712 12954 24746
rect 12988 24712 13022 24746
rect 13056 24712 13090 24746
rect 13124 24712 13158 24746
rect 13192 24712 13226 24746
rect 13260 24712 13294 24746
rect 13328 24712 13362 24746
rect 13396 24712 13430 24746
rect 13464 24712 13498 24746
rect 13532 24712 13566 24746
rect 13600 24712 13634 24746
rect 13668 24712 13702 24746
rect 13736 24712 13770 24746
rect 13804 24712 13838 24746
rect 13872 24712 13906 24746
rect 13940 24712 13974 24746
rect 14008 24712 14042 24746
rect 14076 24712 14110 24746
rect 14144 24712 14178 24746
rect 14212 24712 14246 24746
rect 14280 24712 14314 24746
rect 14348 24712 14382 24746
rect 14416 24712 14450 24746
rect 14484 24712 14518 24746
rect 14552 24712 14586 24746
rect 14620 24712 14654 24746
rect 14688 24712 14722 24746
rect 14756 24712 14790 24746
rect 14824 24712 14858 24746
rect 77 19825 111 19859
rect 146 19825 180 19859
rect 215 19825 249 19859
rect 284 19825 318 19859
rect 353 19825 387 19859
rect 422 19825 456 19859
rect 491 19825 525 19859
rect 560 19825 594 19859
rect 629 19825 663 19859
rect 698 19825 732 19859
rect 767 19825 801 19859
rect 836 19825 870 19859
rect 905 19825 939 19859
rect 974 19825 1008 19859
rect 1043 19825 1077 19859
rect 1112 19825 1146 19859
rect 1181 19825 1215 19859
rect 1250 19825 1284 19859
rect 1319 19825 1353 19859
rect 1388 19825 1422 19859
rect 1457 19825 1491 19859
rect 1526 19825 1560 19859
rect 1595 19825 1629 19859
rect 1664 19825 1698 19859
rect 1733 19825 1767 19859
rect 1802 19825 1836 19859
rect 1871 19825 1905 19859
rect 1940 19825 1974 19859
rect 2009 19825 2043 19859
rect 2078 19825 2112 19859
rect 2147 19825 2181 19859
rect 2216 19825 2250 19859
rect 2285 19825 2319 19859
rect 2354 19825 2388 19859
rect 2423 19825 2457 19859
rect 2492 19825 2526 19859
rect 2561 19825 2595 19859
rect 2630 19825 2664 19859
rect 2699 19825 2733 19859
rect 2768 19825 2802 19859
rect 2837 19825 2871 19859
rect 2906 19825 2940 19859
rect 2975 19825 3009 19859
rect 3044 19825 3078 19859
rect 3113 19825 3147 19859
rect 77 19757 111 19791
rect 146 19757 180 19791
rect 215 19757 249 19791
rect 284 19757 318 19791
rect 353 19757 387 19791
rect 422 19757 456 19791
rect 491 19757 525 19791
rect 560 19757 594 19791
rect 629 19757 663 19791
rect 698 19757 732 19791
rect 767 19757 801 19791
rect 836 19757 870 19791
rect 905 19757 939 19791
rect 974 19757 1008 19791
rect 1043 19757 1077 19791
rect 1112 19757 1146 19791
rect 1181 19757 1215 19791
rect 1250 19757 1284 19791
rect 1319 19757 1353 19791
rect 1388 19757 1422 19791
rect 1457 19757 1491 19791
rect 1526 19757 1560 19791
rect 1595 19757 1629 19791
rect 1664 19757 1698 19791
rect 1733 19757 1767 19791
rect 1802 19757 1836 19791
rect 1871 19757 1905 19791
rect 1940 19757 1974 19791
rect 2009 19757 2043 19791
rect 2078 19757 2112 19791
rect 2147 19757 2181 19791
rect 2216 19757 2250 19791
rect 2285 19757 2319 19791
rect 2354 19757 2388 19791
rect 2423 19757 2457 19791
rect 2492 19757 2526 19791
rect 2561 19757 2595 19791
rect 2630 19757 2664 19791
rect 2699 19757 2733 19791
rect 2768 19757 2802 19791
rect 2837 19757 2871 19791
rect 2906 19757 2940 19791
rect 2975 19757 3009 19791
rect 3044 19757 3078 19791
rect 3113 19757 3147 19791
rect 77 19689 111 19723
rect 146 19689 180 19723
rect 215 19689 249 19723
rect 284 19689 318 19723
rect 353 19689 387 19723
rect 422 19689 456 19723
rect 491 19689 525 19723
rect 560 19689 594 19723
rect 629 19689 663 19723
rect 698 19689 732 19723
rect 767 19689 801 19723
rect 836 19689 870 19723
rect 905 19689 939 19723
rect 974 19689 1008 19723
rect 1043 19689 1077 19723
rect 1112 19689 1146 19723
rect 1181 19689 1215 19723
rect 1250 19689 1284 19723
rect 1319 19689 1353 19723
rect 1388 19689 1422 19723
rect 1457 19689 1491 19723
rect 1526 19689 1560 19723
rect 1595 19689 1629 19723
rect 1664 19689 1698 19723
rect 1733 19689 1767 19723
rect 1802 19689 1836 19723
rect 1871 19689 1905 19723
rect 1940 19689 1974 19723
rect 2009 19689 2043 19723
rect 2078 19689 2112 19723
rect 2147 19689 2181 19723
rect 2216 19689 2250 19723
rect 2285 19689 2319 19723
rect 2354 19689 2388 19723
rect 2423 19689 2457 19723
rect 2492 19689 2526 19723
rect 2561 19689 2595 19723
rect 2630 19689 2664 19723
rect 2699 19689 2733 19723
rect 2768 19689 2802 19723
rect 2837 19689 2871 19723
rect 2906 19689 2940 19723
rect 2975 19689 3009 19723
rect 3044 19689 3078 19723
rect 3113 19689 3147 19723
rect 77 19621 111 19655
rect 146 19621 180 19655
rect 215 19621 249 19655
rect 284 19621 318 19655
rect 353 19621 387 19655
rect 422 19621 456 19655
rect 491 19621 525 19655
rect 560 19621 594 19655
rect 629 19621 663 19655
rect 698 19621 732 19655
rect 767 19621 801 19655
rect 836 19621 870 19655
rect 905 19621 939 19655
rect 974 19621 1008 19655
rect 1043 19621 1077 19655
rect 1112 19621 1146 19655
rect 1181 19621 1215 19655
rect 1250 19621 1284 19655
rect 1319 19621 1353 19655
rect 1388 19621 1422 19655
rect 1457 19621 1491 19655
rect 1526 19621 1560 19655
rect 1595 19621 1629 19655
rect 1664 19621 1698 19655
rect 1733 19621 1767 19655
rect 1802 19621 1836 19655
rect 1871 19621 1905 19655
rect 1940 19621 1974 19655
rect 2009 19621 2043 19655
rect 2078 19621 2112 19655
rect 2147 19621 2181 19655
rect 2216 19621 2250 19655
rect 2285 19621 2319 19655
rect 2354 19621 2388 19655
rect 2423 19621 2457 19655
rect 2492 19621 2526 19655
rect 2561 19621 2595 19655
rect 2630 19621 2664 19655
rect 2699 19621 2733 19655
rect 2768 19621 2802 19655
rect 2837 19621 2871 19655
rect 2906 19621 2940 19655
rect 2975 19621 3009 19655
rect 3044 19621 3078 19655
rect 3113 19621 3147 19655
rect 3182 19621 14436 19859
rect 14484 19797 14518 19831
rect 14567 19797 14601 19831
rect 14650 19797 14684 19831
rect 14733 19797 14767 19831
rect 14816 19797 14850 19831
rect 14484 19727 14518 19761
rect 14567 19727 14601 19761
rect 14650 19727 14684 19761
rect 14733 19727 14767 19761
rect 14816 19727 14850 19761
rect 14484 19657 14518 19691
rect 14567 19657 14601 19691
rect 14650 19657 14684 19691
rect 14733 19657 14767 19691
rect 14816 19657 14850 19691
rect 14484 19587 14518 19621
rect 14567 19587 14601 19621
rect 14650 19587 14684 19621
rect 14733 19587 14767 19621
rect 14816 19587 14850 19621
rect 77 19551 111 19585
rect 146 19551 180 19585
rect 215 19551 249 19585
rect 284 19551 318 19585
rect 353 19551 387 19585
rect 422 19551 456 19585
rect 491 19551 525 19585
rect 560 19551 594 19585
rect 629 19551 663 19585
rect 698 19551 732 19585
rect 767 19551 801 19585
rect 836 19551 870 19585
rect 905 19551 939 19585
rect 974 19551 1008 19585
rect 1043 19551 1077 19585
rect 1112 19551 1146 19585
rect 1181 19551 1215 19585
rect 1250 19551 1284 19585
rect 1319 19551 1353 19585
rect 1388 19551 1422 19585
rect 1457 19551 1491 19585
rect 1526 19551 1560 19585
rect 1595 19551 1629 19585
rect 1664 19551 1698 19585
rect 1733 19551 1767 19585
rect 1802 19551 1836 19585
rect 1871 19551 1905 19585
rect 1940 19551 1974 19585
rect 2009 19551 2043 19585
rect 2078 19551 2112 19585
rect 2147 19551 2181 19585
rect 2216 19551 2250 19585
rect 2285 19551 2319 19585
rect 2354 19551 2388 19585
rect 2423 19551 2457 19585
rect 2492 19551 2526 19585
rect 2561 19551 2595 19585
rect 2630 19551 2664 19585
rect 2699 19551 2733 19585
rect 2768 19551 2802 19585
rect 2837 19551 2871 19585
rect 2906 19551 2940 19585
rect 2975 19551 3009 19585
rect 3044 19551 3078 19585
rect 3113 19551 3147 19585
rect 3182 19551 3216 19585
rect 3251 19551 3285 19585
rect 3320 19551 3354 19585
rect 3389 19551 3423 19585
rect 3458 19551 3492 19585
rect 3527 19551 3561 19585
rect 3596 19551 3630 19585
rect 3665 19551 3699 19585
rect 3733 19551 3767 19585
rect 3801 19551 3835 19585
rect 3869 19551 3903 19585
rect 3937 19551 3971 19585
rect 4005 19551 4039 19585
rect 4073 19551 4107 19585
rect 4141 19551 4175 19585
rect 4209 19551 4243 19585
rect 4277 19551 4311 19585
rect 4345 19551 4379 19585
rect 4413 19551 4447 19585
rect 4481 19551 4515 19585
rect 4549 19551 4583 19585
rect 4617 19551 4651 19585
rect 4685 19551 4719 19585
rect 4753 19551 4787 19585
rect 4821 19551 4855 19585
rect 4889 19551 4923 19585
rect 4957 19551 4991 19585
rect 5025 19551 5059 19585
rect 5093 19551 5127 19585
rect 5161 19551 5195 19585
rect 5229 19551 5263 19585
rect 5297 19551 5331 19585
rect 5365 19551 5399 19585
rect 5433 19551 5467 19585
rect 5501 19551 5535 19585
rect 5569 19551 5603 19585
rect 5637 19551 5671 19585
rect 5705 19551 5739 19585
rect 5773 19551 5807 19585
rect 5841 19551 5875 19585
rect 5909 19551 5943 19585
rect 5977 19551 6011 19585
rect 6045 19551 6079 19585
rect 6113 19551 6147 19585
rect 6181 19551 6215 19585
rect 6249 19551 6283 19585
rect 6317 19551 6351 19585
rect 6385 19551 6419 19585
rect 6453 19551 6487 19585
rect 6521 19551 6555 19585
rect 6589 19551 6623 19585
rect 6657 19551 6691 19585
rect 6725 19551 6759 19585
rect 6793 19551 6827 19585
rect 6861 19551 6895 19585
rect 6929 19551 6963 19585
rect 6997 19551 7031 19585
rect 7065 19551 7099 19585
rect 7133 19551 7167 19585
rect 7201 19551 7235 19585
rect 7269 19551 7303 19585
rect 7337 19551 7371 19585
rect 7405 19551 7439 19585
rect 7473 19551 7507 19585
rect 7541 19551 7575 19585
rect 7609 19551 7643 19585
rect 7677 19551 7711 19585
rect 7745 19551 7779 19585
rect 7813 19551 7847 19585
rect 7881 19551 7915 19585
rect 7949 19551 7983 19585
rect 8017 19551 8051 19585
rect 8085 19551 8119 19585
rect 8153 19551 8187 19585
rect 8221 19551 8255 19585
rect 8289 19551 8323 19585
rect 8357 19551 8391 19585
rect 8425 19551 8459 19585
rect 8493 19551 8527 19585
rect 8561 19551 8595 19585
rect 8629 19551 8663 19585
rect 8697 19551 8731 19585
rect 8765 19551 8799 19585
rect 8833 19551 8867 19585
rect 8901 19551 8935 19585
rect 8969 19551 9003 19585
rect 9037 19551 9071 19585
rect 9105 19551 9139 19585
rect 9173 19551 9207 19585
rect 9241 19551 9275 19585
rect 9309 19551 9343 19585
rect 9377 19551 9411 19585
rect 9445 19551 9479 19585
rect 9513 19551 9547 19585
rect 9581 19551 9615 19585
rect 9649 19551 9683 19585
rect 9717 19551 9751 19585
rect 9785 19551 9819 19585
rect 9853 19551 9887 19585
rect 9921 19551 9955 19585
rect 9989 19551 10023 19585
rect 10057 19551 10091 19585
rect 10125 19551 10159 19585
rect 10193 19551 10227 19585
rect 10261 19551 10295 19585
rect 10329 19551 10363 19585
rect 10397 19551 10431 19585
rect 10465 19551 10499 19585
rect 10533 19551 10567 19585
rect 10601 19551 10635 19585
rect 10669 19551 10703 19585
rect 10737 19551 10771 19585
rect 10805 19551 10839 19585
rect 10873 19551 10907 19585
rect 10941 19551 10975 19585
rect 11009 19551 11043 19585
rect 11077 19551 11111 19585
rect 11145 19551 11179 19585
rect 11213 19551 11247 19585
rect 11281 19551 11315 19585
rect 11349 19551 11383 19585
rect 11417 19551 11451 19585
rect 11485 19551 11519 19585
rect 11553 19551 11587 19585
rect 11621 19551 11655 19585
rect 11689 19551 11723 19585
rect 11771 19523 11805 19557
rect 11841 19523 11875 19557
rect 11911 19523 11945 19557
rect 11981 19523 12015 19557
rect 12051 19523 12085 19557
rect 12121 19523 12155 19557
rect 12191 19523 12225 19557
rect 12261 19523 12295 19557
rect 12331 19523 12365 19557
rect 12401 19523 12435 19557
rect 12470 19523 12504 19557
rect 12539 19523 12573 19557
rect 12608 19523 12642 19557
rect 12677 19523 12711 19557
rect 12746 19523 12780 19557
rect 12815 19523 12849 19557
rect 12884 19523 12918 19557
rect 12953 19523 12987 19557
rect 13022 19523 13056 19557
rect 13091 19523 13125 19557
rect 13160 19523 13194 19557
rect 13229 19523 13263 19557
rect 13298 19523 13332 19557
rect 13367 19523 13401 19557
rect 13436 19523 13470 19557
rect 13505 19523 13539 19557
rect 13574 19523 13608 19557
rect 13643 19523 13677 19557
rect 13712 19523 13746 19557
rect 13781 19523 13815 19557
rect 13850 19523 13884 19557
rect 13919 19523 13953 19557
rect 13988 19523 14022 19557
rect 14057 19523 14091 19557
rect 14126 19523 14160 19557
rect 14195 19523 14229 19557
rect 14264 19523 14298 19557
rect 14333 19523 14367 19557
rect 14402 19523 14436 19557
rect 14484 19517 14518 19551
rect 14567 19517 14601 19551
rect 14650 19517 14684 19551
rect 14733 19517 14767 19551
rect 14816 19517 14850 19551
rect 77 19479 111 19513
rect 146 19479 180 19513
rect 215 19479 249 19513
rect 284 19479 318 19513
rect 353 19479 387 19513
rect 422 19479 456 19513
rect 491 19479 525 19513
rect 560 19479 594 19513
rect 629 19479 663 19513
rect 698 19479 732 19513
rect 767 19479 801 19513
rect 836 19479 870 19513
rect 905 19479 939 19513
rect 974 19479 1008 19513
rect 1043 19479 1077 19513
rect 1112 19479 1146 19513
rect 1181 19479 1215 19513
rect 1250 19479 1284 19513
rect 1319 19479 1353 19513
rect 1388 19479 1422 19513
rect 1457 19479 1491 19513
rect 1526 19479 1560 19513
rect 1595 19479 1629 19513
rect 1664 19479 1698 19513
rect 1733 19479 1767 19513
rect 1802 19479 1836 19513
rect 1871 19479 1905 19513
rect 1940 19479 1974 19513
rect 2009 19479 2043 19513
rect 2078 19479 2112 19513
rect 2147 19479 2181 19513
rect 2216 19479 2250 19513
rect 2285 19479 2319 19513
rect 2354 19479 2388 19513
rect 2423 19479 2457 19513
rect 2492 19479 2526 19513
rect 2561 19479 2595 19513
rect 2630 19479 2664 19513
rect 2699 19479 2733 19513
rect 2768 19479 2802 19513
rect 2837 19479 2871 19513
rect 2906 19479 2940 19513
rect 2975 19479 3009 19513
rect 3044 19479 3078 19513
rect 3113 19479 3147 19513
rect 3182 19479 3216 19513
rect 3251 19479 3285 19513
rect 3320 19479 3354 19513
rect 3389 19479 3423 19513
rect 3458 19479 3492 19513
rect 3527 19479 3561 19513
rect 3596 19479 3630 19513
rect 3665 19479 3699 19513
rect 3733 19479 3767 19513
rect 3801 19479 3835 19513
rect 3869 19479 3903 19513
rect 3937 19479 3971 19513
rect 4005 19479 4039 19513
rect 4073 19479 4107 19513
rect 4141 19479 4175 19513
rect 4209 19479 4243 19513
rect 4277 19479 4311 19513
rect 4345 19479 4379 19513
rect 4413 19479 4447 19513
rect 4481 19479 4515 19513
rect 4549 19479 4583 19513
rect 4617 19479 4651 19513
rect 4685 19479 4719 19513
rect 4753 19479 4787 19513
rect 4821 19479 4855 19513
rect 4889 19479 4923 19513
rect 4957 19479 4991 19513
rect 5025 19479 5059 19513
rect 5093 19479 5127 19513
rect 5161 19479 5195 19513
rect 5229 19479 5263 19513
rect 5297 19479 5331 19513
rect 5365 19479 5399 19513
rect 5433 19479 5467 19513
rect 5501 19479 5535 19513
rect 5569 19479 5603 19513
rect 5637 19479 5671 19513
rect 5705 19479 5739 19513
rect 5773 19479 5807 19513
rect 5841 19479 5875 19513
rect 5909 19479 5943 19513
rect 5977 19479 6011 19513
rect 6045 19479 6079 19513
rect 6113 19479 6147 19513
rect 6181 19479 6215 19513
rect 6249 19479 6283 19513
rect 6317 19479 6351 19513
rect 6385 19479 6419 19513
rect 6453 19479 6487 19513
rect 6521 19479 6555 19513
rect 6589 19479 6623 19513
rect 6657 19479 6691 19513
rect 6725 19479 6759 19513
rect 6793 19479 6827 19513
rect 6861 19479 6895 19513
rect 6929 19479 6963 19513
rect 6997 19479 7031 19513
rect 7065 19479 7099 19513
rect 7133 19479 7167 19513
rect 7201 19479 7235 19513
rect 7269 19479 7303 19513
rect 7337 19479 7371 19513
rect 7405 19479 7439 19513
rect 7473 19479 7507 19513
rect 7541 19479 7575 19513
rect 7609 19479 7643 19513
rect 7677 19479 7711 19513
rect 7745 19479 7779 19513
rect 7813 19479 7847 19513
rect 7881 19479 7915 19513
rect 7949 19479 7983 19513
rect 8017 19479 8051 19513
rect 8085 19479 8119 19513
rect 8153 19479 8187 19513
rect 8221 19479 8255 19513
rect 8289 19479 8323 19513
rect 8357 19479 8391 19513
rect 8425 19479 8459 19513
rect 8493 19479 8527 19513
rect 8561 19479 8595 19513
rect 8629 19479 8663 19513
rect 8697 19479 8731 19513
rect 8765 19479 8799 19513
rect 8833 19479 8867 19513
rect 8901 19479 8935 19513
rect 8969 19479 9003 19513
rect 9037 19479 9071 19513
rect 9105 19479 9139 19513
rect 9173 19479 9207 19513
rect 9241 19479 9275 19513
rect 9309 19479 9343 19513
rect 9377 19479 9411 19513
rect 9445 19479 9479 19513
rect 9513 19479 9547 19513
rect 9581 19479 9615 19513
rect 9649 19479 9683 19513
rect 9717 19479 9751 19513
rect 9785 19479 9819 19513
rect 9853 19479 9887 19513
rect 9921 19479 9955 19513
rect 9989 19479 10023 19513
rect 10057 19479 10091 19513
rect 10125 19479 10159 19513
rect 10193 19479 10227 19513
rect 10261 19479 10295 19513
rect 10329 19479 10363 19513
rect 10397 19479 10431 19513
rect 10465 19479 10499 19513
rect 10533 19479 10567 19513
rect 10601 19479 10635 19513
rect 10669 19479 10703 19513
rect 10737 19479 10771 19513
rect 10805 19479 10839 19513
rect 10873 19479 10907 19513
rect 10941 19479 10975 19513
rect 11009 19479 11043 19513
rect 11077 19479 11111 19513
rect 11145 19479 11179 19513
rect 11213 19479 11247 19513
rect 11281 19479 11315 19513
rect 11349 19479 11383 19513
rect 11417 19479 11451 19513
rect 11485 19479 11519 19513
rect 11553 19479 11587 19513
rect 11621 19479 11655 19513
rect 11689 19479 11723 19513
rect 11771 19443 11805 19477
rect 11841 19443 11875 19477
rect 11911 19443 11945 19477
rect 11981 19443 12015 19477
rect 12051 19443 12085 19477
rect 12121 19443 12155 19477
rect 12191 19443 12225 19477
rect 12261 19443 12295 19477
rect 12331 19443 12365 19477
rect 12401 19443 12435 19477
rect 12470 19443 12504 19477
rect 12539 19443 12573 19477
rect 12608 19443 12642 19477
rect 12677 19443 12711 19477
rect 12746 19443 12780 19477
rect 12815 19443 12849 19477
rect 12884 19443 12918 19477
rect 12953 19443 12987 19477
rect 13022 19443 13056 19477
rect 13091 19443 13125 19477
rect 13160 19443 13194 19477
rect 13229 19443 13263 19477
rect 13298 19443 13332 19477
rect 13367 19443 13401 19477
rect 13436 19443 13470 19477
rect 13505 19443 13539 19477
rect 13574 19443 13608 19477
rect 13643 19443 13677 19477
rect 13712 19443 13746 19477
rect 13781 19443 13815 19477
rect 13850 19443 13884 19477
rect 13919 19443 13953 19477
rect 13988 19443 14022 19477
rect 14057 19443 14091 19477
rect 14126 19443 14160 19477
rect 14195 19443 14229 19477
rect 14264 19443 14298 19477
rect 14333 19443 14367 19477
rect 14402 19443 14436 19477
rect 14484 19447 14518 19481
rect 14567 19447 14601 19481
rect 14650 19447 14684 19481
rect 14733 19447 14767 19481
rect 14816 19447 14850 19481
rect 77 19407 111 19441
rect 146 19407 180 19441
rect 215 19407 249 19441
rect 284 19407 318 19441
rect 353 19407 387 19441
rect 422 19407 456 19441
rect 491 19407 525 19441
rect 560 19407 594 19441
rect 629 19407 663 19441
rect 698 19407 732 19441
rect 767 19407 801 19441
rect 836 19407 870 19441
rect 905 19407 939 19441
rect 974 19407 1008 19441
rect 1043 19407 1077 19441
rect 1112 19407 1146 19441
rect 1181 19407 1215 19441
rect 1250 19407 1284 19441
rect 1319 19407 1353 19441
rect 1388 19407 1422 19441
rect 1457 19407 1491 19441
rect 1526 19407 1560 19441
rect 1595 19407 1629 19441
rect 1664 19407 1698 19441
rect 1733 19407 1767 19441
rect 1802 19407 1836 19441
rect 1871 19407 1905 19441
rect 1940 19407 1974 19441
rect 2009 19407 2043 19441
rect 2078 19407 2112 19441
rect 2147 19407 2181 19441
rect 2216 19407 2250 19441
rect 2285 19407 2319 19441
rect 2354 19407 2388 19441
rect 2423 19407 2457 19441
rect 2492 19407 2526 19441
rect 2561 19407 2595 19441
rect 2630 19407 2664 19441
rect 2699 19407 2733 19441
rect 2768 19407 2802 19441
rect 2837 19407 2871 19441
rect 2906 19407 2940 19441
rect 2975 19407 3009 19441
rect 3044 19407 3078 19441
rect 3113 19407 3147 19441
rect 3182 19407 3216 19441
rect 3251 19407 3285 19441
rect 3320 19407 3354 19441
rect 3389 19407 3423 19441
rect 3458 19407 3492 19441
rect 3527 19407 3561 19441
rect 3596 19407 3630 19441
rect 3665 19407 3699 19441
rect 3733 19407 3767 19441
rect 3801 19407 3835 19441
rect 3869 19407 3903 19441
rect 3937 19407 3971 19441
rect 4005 19407 4039 19441
rect 4073 19407 4107 19441
rect 4141 19407 4175 19441
rect 4209 19407 4243 19441
rect 4277 19407 4311 19441
rect 4345 19407 4379 19441
rect 4413 19407 4447 19441
rect 4481 19407 4515 19441
rect 4549 19407 4583 19441
rect 4617 19407 4651 19441
rect 4685 19407 4719 19441
rect 4753 19407 4787 19441
rect 4821 19407 4855 19441
rect 4889 19407 4923 19441
rect 4957 19407 4991 19441
rect 5025 19407 5059 19441
rect 5093 19407 5127 19441
rect 5161 19407 5195 19441
rect 5229 19407 5263 19441
rect 5297 19407 5331 19441
rect 5365 19407 5399 19441
rect 5433 19407 5467 19441
rect 5501 19407 5535 19441
rect 5569 19407 5603 19441
rect 5637 19407 5671 19441
rect 5705 19407 5739 19441
rect 5773 19407 5807 19441
rect 5841 19407 5875 19441
rect 5909 19407 5943 19441
rect 5977 19407 6011 19441
rect 6045 19407 6079 19441
rect 6113 19407 6147 19441
rect 6181 19407 6215 19441
rect 6249 19407 6283 19441
rect 6317 19407 6351 19441
rect 6385 19407 6419 19441
rect 6453 19407 6487 19441
rect 6521 19407 6555 19441
rect 6589 19407 6623 19441
rect 6657 19407 6691 19441
rect 6725 19407 6759 19441
rect 6793 19407 6827 19441
rect 6861 19407 6895 19441
rect 6929 19407 6963 19441
rect 6997 19407 7031 19441
rect 7065 19407 7099 19441
rect 7133 19407 7167 19441
rect 7201 19407 7235 19441
rect 7269 19407 7303 19441
rect 7337 19407 7371 19441
rect 7405 19407 7439 19441
rect 7473 19407 7507 19441
rect 7541 19407 7575 19441
rect 7609 19407 7643 19441
rect 7677 19407 7711 19441
rect 7745 19407 7779 19441
rect 7813 19407 7847 19441
rect 7881 19407 7915 19441
rect 7949 19407 7983 19441
rect 8017 19407 8051 19441
rect 8085 19407 8119 19441
rect 8153 19407 8187 19441
rect 8221 19407 8255 19441
rect 8289 19407 8323 19441
rect 8357 19407 8391 19441
rect 8425 19407 8459 19441
rect 8493 19407 8527 19441
rect 8561 19407 8595 19441
rect 8629 19407 8663 19441
rect 8697 19407 8731 19441
rect 8765 19407 8799 19441
rect 8833 19407 8867 19441
rect 8901 19407 8935 19441
rect 8969 19407 9003 19441
rect 9037 19407 9071 19441
rect 9105 19407 9139 19441
rect 9173 19407 9207 19441
rect 9241 19407 9275 19441
rect 9309 19407 9343 19441
rect 9377 19407 9411 19441
rect 9445 19407 9479 19441
rect 9513 19407 9547 19441
rect 9581 19407 9615 19441
rect 9649 19407 9683 19441
rect 9717 19407 9751 19441
rect 9785 19407 9819 19441
rect 9853 19407 9887 19441
rect 9921 19407 9955 19441
rect 9989 19407 10023 19441
rect 10057 19407 10091 19441
rect 10125 19407 10159 19441
rect 10193 19407 10227 19441
rect 10261 19407 10295 19441
rect 10329 19407 10363 19441
rect 10397 19407 10431 19441
rect 10465 19407 10499 19441
rect 10533 19407 10567 19441
rect 10601 19407 10635 19441
rect 10669 19407 10703 19441
rect 10737 19407 10771 19441
rect 10805 19407 10839 19441
rect 10873 19407 10907 19441
rect 10941 19407 10975 19441
rect 11009 19407 11043 19441
rect 11077 19407 11111 19441
rect 11145 19407 11179 19441
rect 11213 19407 11247 19441
rect 11281 19407 11315 19441
rect 11349 19407 11383 19441
rect 11417 19407 11451 19441
rect 11485 19407 11519 19441
rect 11553 19407 11587 19441
rect 11621 19407 11655 19441
rect 11689 19407 11723 19441
rect 77 19335 111 19369
rect 146 19335 180 19369
rect 215 19335 249 19369
rect 284 19335 318 19369
rect 353 19335 387 19369
rect 422 19335 456 19369
rect 491 19335 525 19369
rect 560 19335 594 19369
rect 629 19335 663 19369
rect 698 19335 732 19369
rect 767 19335 801 19369
rect 836 19335 870 19369
rect 905 19335 939 19369
rect 974 19335 1008 19369
rect 1043 19335 1077 19369
rect 1112 19335 1146 19369
rect 1181 19335 1215 19369
rect 1250 19335 1284 19369
rect 1319 19335 1353 19369
rect 1388 19335 1422 19369
rect 1457 19335 1491 19369
rect 1526 19335 1560 19369
rect 1595 19335 1629 19369
rect 1664 19335 1698 19369
rect 1733 19335 1767 19369
rect 1802 19335 1836 19369
rect 1871 19335 1905 19369
rect 1940 19335 1974 19369
rect 2009 19335 2043 19369
rect 2078 19335 2112 19369
rect 2147 19335 2181 19369
rect 2216 19335 2250 19369
rect 2285 19335 2319 19369
rect 2354 19335 2388 19369
rect 2423 19335 2457 19369
rect 2492 19335 2526 19369
rect 2561 19335 2595 19369
rect 2630 19335 2664 19369
rect 2699 19335 2733 19369
rect 2768 19335 2802 19369
rect 2837 19335 2871 19369
rect 2906 19335 2940 19369
rect 2975 19335 3009 19369
rect 3044 19335 3078 19369
rect 3113 19335 3147 19369
rect 3182 19335 3216 19369
rect 3251 19335 3285 19369
rect 3320 19335 3354 19369
rect 3389 19335 3423 19369
rect 3458 19335 3492 19369
rect 3527 19335 3561 19369
rect 3596 19335 3630 19369
rect 3665 19335 3699 19369
rect 3733 19335 3767 19369
rect 3801 19335 3835 19369
rect 3869 19335 3903 19369
rect 3937 19335 3971 19369
rect 4005 19335 4039 19369
rect 4073 19335 4107 19369
rect 4141 19335 4175 19369
rect 4209 19335 4243 19369
rect 4277 19335 4311 19369
rect 4345 19335 4379 19369
rect 4413 19335 4447 19369
rect 4481 19335 4515 19369
rect 4549 19335 4583 19369
rect 4617 19335 4651 19369
rect 4685 19335 4719 19369
rect 4753 19335 4787 19369
rect 4821 19335 4855 19369
rect 4889 19335 4923 19369
rect 4957 19335 4991 19369
rect 5025 19335 5059 19369
rect 5093 19335 5127 19369
rect 5161 19335 5195 19369
rect 5229 19335 5263 19369
rect 5297 19335 5331 19369
rect 5365 19335 5399 19369
rect 5433 19335 5467 19369
rect 5501 19335 5535 19369
rect 5569 19335 5603 19369
rect 5637 19335 5671 19369
rect 5705 19335 5739 19369
rect 5773 19335 5807 19369
rect 5841 19335 5875 19369
rect 5909 19335 5943 19369
rect 5977 19335 6011 19369
rect 6045 19335 6079 19369
rect 6113 19335 6147 19369
rect 6181 19335 6215 19369
rect 6249 19335 6283 19369
rect 6317 19335 6351 19369
rect 6385 19335 6419 19369
rect 6453 19335 6487 19369
rect 6521 19335 6555 19369
rect 6589 19335 6623 19369
rect 6657 19335 6691 19369
rect 6725 19335 6759 19369
rect 6793 19335 6827 19369
rect 6861 19335 6895 19369
rect 6929 19335 6963 19369
rect 6997 19335 7031 19369
rect 7065 19335 7099 19369
rect 7133 19335 7167 19369
rect 7201 19335 7235 19369
rect 7269 19335 7303 19369
rect 7337 19335 7371 19369
rect 7405 19335 7439 19369
rect 7473 19335 7507 19369
rect 7541 19335 7575 19369
rect 7609 19335 7643 19369
rect 7677 19335 7711 19369
rect 7745 19335 7779 19369
rect 7813 19335 7847 19369
rect 7881 19335 7915 19369
rect 7949 19335 7983 19369
rect 8017 19335 8051 19369
rect 8085 19335 8119 19369
rect 8153 19335 8187 19369
rect 8221 19335 8255 19369
rect 8289 19335 8323 19369
rect 8357 19335 8391 19369
rect 8425 19335 8459 19369
rect 8493 19335 8527 19369
rect 8561 19335 8595 19369
rect 8629 19335 8663 19369
rect 8697 19335 8731 19369
rect 8765 19335 8799 19369
rect 8833 19335 8867 19369
rect 8901 19335 8935 19369
rect 8969 19335 9003 19369
rect 9037 19335 9071 19369
rect 9105 19335 9139 19369
rect 9173 19335 9207 19369
rect 9241 19335 9275 19369
rect 9309 19335 9343 19369
rect 9377 19335 9411 19369
rect 9445 19335 9479 19369
rect 9513 19335 9547 19369
rect 9581 19335 9615 19369
rect 9649 19335 9683 19369
rect 9717 19335 9751 19369
rect 9785 19335 9819 19369
rect 9853 19335 9887 19369
rect 9921 19335 9955 19369
rect 9989 19335 10023 19369
rect 10057 19335 10091 19369
rect 10125 19335 10159 19369
rect 10193 19335 10227 19369
rect 10261 19335 10295 19369
rect 10329 19335 10363 19369
rect 10397 19335 10431 19369
rect 10465 19335 10499 19369
rect 10533 19335 10567 19369
rect 10601 19335 10635 19369
rect 10669 19335 10703 19369
rect 10737 19335 10771 19369
rect 10805 19335 10839 19369
rect 10873 19335 10907 19369
rect 10941 19335 10975 19369
rect 11009 19335 11043 19369
rect 11077 19335 11111 19369
rect 11145 19335 11179 19369
rect 11213 19335 11247 19369
rect 11281 19335 11315 19369
rect 11349 19335 11383 19369
rect 11417 19335 11451 19369
rect 11485 19335 11519 19369
rect 11553 19335 11587 19369
rect 11621 19335 11655 19369
rect 11689 19335 11723 19369
rect 11771 19363 11805 19397
rect 11841 19363 11875 19397
rect 11911 19363 11945 19397
rect 11981 19363 12015 19397
rect 12051 19363 12085 19397
rect 12121 19363 12155 19397
rect 12191 19363 12225 19397
rect 12261 19363 12295 19397
rect 12331 19363 12365 19397
rect 12401 19363 12435 19397
rect 12470 19363 12504 19397
rect 12539 19363 12573 19397
rect 12608 19363 12642 19397
rect 12677 19363 12711 19397
rect 12746 19363 12780 19397
rect 12815 19363 12849 19397
rect 12884 19363 12918 19397
rect 12953 19363 12987 19397
rect 13022 19363 13056 19397
rect 13091 19363 13125 19397
rect 13160 19363 13194 19397
rect 13229 19363 13263 19397
rect 13298 19363 13332 19397
rect 13367 19363 13401 19397
rect 13436 19363 13470 19397
rect 13505 19363 13539 19397
rect 13574 19363 13608 19397
rect 13643 19363 13677 19397
rect 13712 19363 13746 19397
rect 13781 19363 13815 19397
rect 13850 19363 13884 19397
rect 13919 19363 13953 19397
rect 13988 19363 14022 19397
rect 14057 19363 14091 19397
rect 14126 19363 14160 19397
rect 14195 19363 14229 19397
rect 14264 19363 14298 19397
rect 14333 19363 14367 19397
rect 14402 19363 14436 19397
rect 14484 19377 14518 19411
rect 14567 19377 14601 19411
rect 14650 19377 14684 19411
rect 14733 19377 14767 19411
rect 14816 19377 14850 19411
rect 77 19263 111 19297
rect 146 19263 180 19297
rect 215 19263 249 19297
rect 284 19263 318 19297
rect 353 19263 387 19297
rect 422 19263 456 19297
rect 491 19263 525 19297
rect 560 19263 594 19297
rect 629 19263 663 19297
rect 698 19263 732 19297
rect 767 19263 801 19297
rect 836 19263 870 19297
rect 905 19263 939 19297
rect 974 19263 1008 19297
rect 1043 19263 1077 19297
rect 1112 19263 1146 19297
rect 1181 19263 1215 19297
rect 1250 19263 1284 19297
rect 1319 19263 1353 19297
rect 1388 19263 1422 19297
rect 1457 19263 1491 19297
rect 1526 19263 1560 19297
rect 1595 19263 1629 19297
rect 1664 19263 1698 19297
rect 1733 19263 1767 19297
rect 1802 19263 1836 19297
rect 1871 19263 1905 19297
rect 1940 19263 1974 19297
rect 2009 19263 2043 19297
rect 2078 19263 2112 19297
rect 2147 19263 2181 19297
rect 2216 19263 2250 19297
rect 2285 19263 2319 19297
rect 2354 19263 2388 19297
rect 2423 19263 2457 19297
rect 2492 19263 2526 19297
rect 2561 19263 2595 19297
rect 2630 19263 2664 19297
rect 2699 19263 2733 19297
rect 2768 19263 2802 19297
rect 2837 19263 2871 19297
rect 2906 19263 2940 19297
rect 2975 19263 3009 19297
rect 3044 19263 3078 19297
rect 3113 19263 3147 19297
rect 3182 19263 3216 19297
rect 3251 19263 3285 19297
rect 3320 19263 3354 19297
rect 3389 19263 3423 19297
rect 3458 19263 3492 19297
rect 3527 19263 3561 19297
rect 3596 19263 3630 19297
rect 3665 19263 3699 19297
rect 3733 19263 3767 19297
rect 3801 19263 3835 19297
rect 3869 19263 3903 19297
rect 3937 19263 3971 19297
rect 4005 19263 4039 19297
rect 4073 19263 4107 19297
rect 4141 19263 4175 19297
rect 4209 19263 4243 19297
rect 4277 19263 4311 19297
rect 4345 19263 4379 19297
rect 4413 19263 4447 19297
rect 4481 19263 4515 19297
rect 4549 19263 4583 19297
rect 4617 19263 4651 19297
rect 4685 19263 4719 19297
rect 4753 19263 4787 19297
rect 4821 19263 4855 19297
rect 4889 19263 4923 19297
rect 4957 19263 4991 19297
rect 5025 19263 5059 19297
rect 5093 19263 5127 19297
rect 5161 19263 5195 19297
rect 5229 19263 5263 19297
rect 5297 19263 5331 19297
rect 5365 19263 5399 19297
rect 5433 19263 5467 19297
rect 5501 19263 5535 19297
rect 5569 19263 5603 19297
rect 5637 19263 5671 19297
rect 5705 19263 5739 19297
rect 5773 19263 5807 19297
rect 5841 19263 5875 19297
rect 5909 19263 5943 19297
rect 5977 19263 6011 19297
rect 6045 19263 6079 19297
rect 6113 19263 6147 19297
rect 6181 19263 6215 19297
rect 6249 19263 6283 19297
rect 6317 19263 6351 19297
rect 6385 19263 6419 19297
rect 6453 19263 6487 19297
rect 6521 19263 6555 19297
rect 6589 19263 6623 19297
rect 6657 19263 6691 19297
rect 6725 19263 6759 19297
rect 6793 19263 6827 19297
rect 6861 19263 6895 19297
rect 6929 19263 6963 19297
rect 6997 19263 7031 19297
rect 7065 19263 7099 19297
rect 7133 19263 7167 19297
rect 7201 19263 7235 19297
rect 7269 19263 7303 19297
rect 7337 19263 7371 19297
rect 7405 19263 7439 19297
rect 7473 19263 7507 19297
rect 7541 19263 7575 19297
rect 7609 19263 7643 19297
rect 7677 19263 7711 19297
rect 7745 19263 7779 19297
rect 7813 19263 7847 19297
rect 7881 19263 7915 19297
rect 7949 19263 7983 19297
rect 8017 19263 8051 19297
rect 8085 19263 8119 19297
rect 8153 19263 8187 19297
rect 8221 19263 8255 19297
rect 8289 19263 8323 19297
rect 8357 19263 8391 19297
rect 8425 19263 8459 19297
rect 8493 19263 8527 19297
rect 8561 19263 8595 19297
rect 8629 19263 8663 19297
rect 8697 19263 8731 19297
rect 8765 19263 8799 19297
rect 8833 19263 8867 19297
rect 8901 19263 8935 19297
rect 8969 19263 9003 19297
rect 9037 19263 9071 19297
rect 9105 19263 9139 19297
rect 9173 19263 9207 19297
rect 9241 19263 9275 19297
rect 9309 19263 9343 19297
rect 9377 19263 9411 19297
rect 9445 19263 9479 19297
rect 9513 19263 9547 19297
rect 9581 19263 9615 19297
rect 9649 19263 9683 19297
rect 9717 19263 9751 19297
rect 9785 19263 9819 19297
rect 9853 19263 9887 19297
rect 9921 19263 9955 19297
rect 9989 19263 10023 19297
rect 10057 19263 10091 19297
rect 10125 19263 10159 19297
rect 10193 19263 10227 19297
rect 10261 19263 10295 19297
rect 10329 19263 10363 19297
rect 10397 19263 10431 19297
rect 10465 19263 10499 19297
rect 10533 19263 10567 19297
rect 10601 19263 10635 19297
rect 10669 19263 10703 19297
rect 10737 19263 10771 19297
rect 10805 19263 10839 19297
rect 10873 19263 10907 19297
rect 10941 19263 10975 19297
rect 11009 19263 11043 19297
rect 11077 19263 11111 19297
rect 11145 19263 11179 19297
rect 11213 19263 11247 19297
rect 11281 19263 11315 19297
rect 11349 19263 11383 19297
rect 11417 19263 11451 19297
rect 11485 19263 11519 19297
rect 11553 19263 11587 19297
rect 11621 19263 11655 19297
rect 11689 19263 11723 19297
rect 77 19191 111 19225
rect 146 19191 180 19225
rect 215 19191 249 19225
rect 284 19191 318 19225
rect 353 19191 387 19225
rect 422 19191 456 19225
rect 491 19191 525 19225
rect 560 19191 594 19225
rect 629 19191 663 19225
rect 698 19191 732 19225
rect 767 19191 801 19225
rect 836 19191 870 19225
rect 905 19191 939 19225
rect 974 19191 1008 19225
rect 1043 19191 1077 19225
rect 1112 19191 1146 19225
rect 1181 19191 1215 19225
rect 1250 19191 1284 19225
rect 1319 19191 1353 19225
rect 1388 19191 1422 19225
rect 1457 19191 1491 19225
rect 1526 19191 1560 19225
rect 1595 19191 1629 19225
rect 1664 19191 1698 19225
rect 1733 19191 1767 19225
rect 1802 19191 1836 19225
rect 1871 19191 1905 19225
rect 1940 19191 1974 19225
rect 2009 19191 2043 19225
rect 2078 19191 2112 19225
rect 2147 19191 2181 19225
rect 2216 19191 2250 19225
rect 2285 19191 2319 19225
rect 2354 19191 2388 19225
rect 2423 19191 2457 19225
rect 2492 19191 2526 19225
rect 2561 19191 2595 19225
rect 2630 19191 2664 19225
rect 2699 19191 2733 19225
rect 2768 19191 2802 19225
rect 2837 19191 2871 19225
rect 2906 19191 2940 19225
rect 2975 19191 3009 19225
rect 3044 19191 3078 19225
rect 3113 19191 3147 19225
rect 3182 19191 3216 19225
rect 3251 19191 3285 19225
rect 3320 19191 3354 19225
rect 3389 19191 3423 19225
rect 3458 19191 3492 19225
rect 3527 19191 3561 19225
rect 3596 19191 3630 19225
rect 3665 19191 3699 19225
rect 3733 19191 3767 19225
rect 3801 19191 3835 19225
rect 3869 19191 3903 19225
rect 3937 19191 3971 19225
rect 4005 19191 4039 19225
rect 4073 19191 4107 19225
rect 4141 19191 4175 19225
rect 4209 19191 4243 19225
rect 4277 19191 4311 19225
rect 4345 19191 4379 19225
rect 4413 19191 4447 19225
rect 4481 19191 4515 19225
rect 4549 19191 4583 19225
rect 4617 19191 4651 19225
rect 4685 19191 4719 19225
rect 4753 19191 4787 19225
rect 4821 19191 4855 19225
rect 4889 19191 4923 19225
rect 4957 19191 4991 19225
rect 5025 19191 5059 19225
rect 5093 19191 5127 19225
rect 5161 19191 5195 19225
rect 5229 19191 5263 19225
rect 5297 19191 5331 19225
rect 5365 19191 5399 19225
rect 5433 19191 5467 19225
rect 5501 19191 5535 19225
rect 5569 19191 5603 19225
rect 5637 19191 5671 19225
rect 5705 19191 5739 19225
rect 5773 19191 5807 19225
rect 5841 19191 5875 19225
rect 5909 19191 5943 19225
rect 5977 19191 6011 19225
rect 6045 19191 6079 19225
rect 6113 19191 6147 19225
rect 6181 19191 6215 19225
rect 6249 19191 6283 19225
rect 6317 19191 6351 19225
rect 6385 19191 6419 19225
rect 6453 19191 6487 19225
rect 6521 19191 6555 19225
rect 6589 19191 6623 19225
rect 6657 19191 6691 19225
rect 6725 19191 6759 19225
rect 6793 19191 6827 19225
rect 6861 19191 6895 19225
rect 6929 19191 6963 19225
rect 6997 19191 7031 19225
rect 7065 19191 7099 19225
rect 7133 19191 7167 19225
rect 7201 19191 7235 19225
rect 7269 19191 7303 19225
rect 7337 19191 7371 19225
rect 7405 19191 7439 19225
rect 7473 19191 7507 19225
rect 7541 19191 7575 19225
rect 7609 19191 7643 19225
rect 7677 19191 7711 19225
rect 7745 19191 7779 19225
rect 7813 19191 7847 19225
rect 7881 19191 7915 19225
rect 7949 19191 7983 19225
rect 8017 19191 8051 19225
rect 8085 19191 8119 19225
rect 8153 19191 8187 19225
rect 8221 19191 8255 19225
rect 8289 19191 8323 19225
rect 8357 19191 8391 19225
rect 8425 19191 8459 19225
rect 8493 19191 8527 19225
rect 8561 19191 8595 19225
rect 8629 19191 8663 19225
rect 8697 19191 8731 19225
rect 8765 19191 8799 19225
rect 8833 19191 8867 19225
rect 8901 19191 8935 19225
rect 8969 19191 9003 19225
rect 9037 19191 9071 19225
rect 9105 19191 9139 19225
rect 9173 19191 9207 19225
rect 9241 19191 9275 19225
rect 9309 19191 9343 19225
rect 9377 19191 9411 19225
rect 9445 19191 9479 19225
rect 9513 19191 9547 19225
rect 9581 19191 9615 19225
rect 9649 19191 9683 19225
rect 9717 19191 9751 19225
rect 9785 19191 9819 19225
rect 9853 19191 9887 19225
rect 9921 19191 9955 19225
rect 9989 19191 10023 19225
rect 10057 19191 10091 19225
rect 10125 19191 10159 19225
rect 10193 19191 10227 19225
rect 10261 19191 10295 19225
rect 10329 19191 10363 19225
rect 10397 19191 10431 19225
rect 10465 19191 10499 19225
rect 10533 19191 10567 19225
rect 10601 19191 10635 19225
rect 10669 19191 10703 19225
rect 10737 19191 10771 19225
rect 10805 19191 10839 19225
rect 10873 19191 10907 19225
rect 10941 19191 10975 19225
rect 11009 19191 11043 19225
rect 11077 19191 11111 19225
rect 11145 19191 11179 19225
rect 11213 19191 11247 19225
rect 11281 19191 11315 19225
rect 11349 19191 11383 19225
rect 11417 19191 11451 19225
rect 11485 19191 11519 19225
rect 11553 19191 11587 19225
rect 11621 19191 11655 19225
rect 11689 19191 11723 19225
rect 77 19119 111 19153
rect 146 19119 180 19153
rect 215 19119 249 19153
rect 284 19119 318 19153
rect 353 19119 387 19153
rect 422 19119 456 19153
rect 491 19119 525 19153
rect 560 19119 594 19153
rect 629 19119 663 19153
rect 698 19119 732 19153
rect 767 19119 801 19153
rect 836 19119 870 19153
rect 905 19119 939 19153
rect 974 19119 1008 19153
rect 1043 19119 1077 19153
rect 1112 19119 1146 19153
rect 1181 19119 1215 19153
rect 1250 19119 1284 19153
rect 1319 19119 1353 19153
rect 1388 19119 1422 19153
rect 1457 19119 1491 19153
rect 1526 19119 1560 19153
rect 1595 19119 1629 19153
rect 1664 19119 1698 19153
rect 1733 19119 1767 19153
rect 1802 19119 1836 19153
rect 1871 19119 1905 19153
rect 1940 19119 1974 19153
rect 2009 19119 2043 19153
rect 2078 19119 2112 19153
rect 2147 19119 2181 19153
rect 2216 19119 2250 19153
rect 2285 19119 2319 19153
rect 2354 19119 2388 19153
rect 2423 19119 2457 19153
rect 2492 19119 2526 19153
rect 2561 19119 2595 19153
rect 2630 19119 2664 19153
rect 2699 19119 2733 19153
rect 2768 19119 2802 19153
rect 2837 19119 2871 19153
rect 2906 19119 2940 19153
rect 2975 19119 3009 19153
rect 3044 19119 3078 19153
rect 3113 19119 3147 19153
rect 3182 19119 3216 19153
rect 3251 19119 3285 19153
rect 3320 19119 3354 19153
rect 3389 19119 3423 19153
rect 3458 19119 3492 19153
rect 3527 19119 3561 19153
rect 3596 19119 3630 19153
rect 3665 19119 3699 19153
rect 3733 19119 3767 19153
rect 3801 19119 3835 19153
rect 3869 19119 3903 19153
rect 3937 19119 3971 19153
rect 4005 19119 4039 19153
rect 4073 19119 4107 19153
rect 4141 19119 4175 19153
rect 4209 19119 4243 19153
rect 4277 19119 4311 19153
rect 4345 19119 4379 19153
rect 4413 19119 4447 19153
rect 4481 19119 4515 19153
rect 4549 19119 4583 19153
rect 4617 19119 4651 19153
rect 4685 19119 4719 19153
rect 4753 19119 4787 19153
rect 4821 19119 4855 19153
rect 4889 19119 4923 19153
rect 4957 19119 4991 19153
rect 5025 19119 5059 19153
rect 5093 19119 5127 19153
rect 5161 19119 5195 19153
rect 5229 19119 5263 19153
rect 5297 19119 5331 19153
rect 5365 19119 5399 19153
rect 5433 19119 5467 19153
rect 5501 19119 5535 19153
rect 5569 19119 5603 19153
rect 5637 19119 5671 19153
rect 5705 19119 5739 19153
rect 5773 19119 5807 19153
rect 5841 19119 5875 19153
rect 5909 19119 5943 19153
rect 5977 19119 6011 19153
rect 6045 19119 6079 19153
rect 6113 19119 6147 19153
rect 6181 19119 6215 19153
rect 6249 19119 6283 19153
rect 6317 19119 6351 19153
rect 6385 19119 6419 19153
rect 6453 19119 6487 19153
rect 6521 19119 6555 19153
rect 6589 19119 6623 19153
rect 6657 19119 6691 19153
rect 6725 19119 6759 19153
rect 6793 19119 6827 19153
rect 6861 19119 6895 19153
rect 6929 19119 6963 19153
rect 6997 19119 7031 19153
rect 7065 19119 7099 19153
rect 7133 19119 7167 19153
rect 7201 19119 7235 19153
rect 7269 19119 7303 19153
rect 7337 19119 7371 19153
rect 7405 19119 7439 19153
rect 7473 19119 7507 19153
rect 7541 19119 7575 19153
rect 7609 19119 7643 19153
rect 7677 19119 7711 19153
rect 7745 19119 7779 19153
rect 7813 19119 7847 19153
rect 7881 19119 7915 19153
rect 7949 19119 7983 19153
rect 8017 19119 8051 19153
rect 8085 19119 8119 19153
rect 8153 19119 8187 19153
rect 8221 19119 8255 19153
rect 8289 19119 8323 19153
rect 8357 19119 8391 19153
rect 8425 19119 8459 19153
rect 8493 19119 8527 19153
rect 8561 19119 8595 19153
rect 8629 19119 8663 19153
rect 8697 19119 8731 19153
rect 8765 19119 8799 19153
rect 8833 19119 8867 19153
rect 8901 19119 8935 19153
rect 8969 19119 9003 19153
rect 9037 19119 9071 19153
rect 9105 19119 9139 19153
rect 9173 19119 9207 19153
rect 9241 19119 9275 19153
rect 9309 19119 9343 19153
rect 9377 19119 9411 19153
rect 9445 19119 9479 19153
rect 9513 19119 9547 19153
rect 9581 19119 9615 19153
rect 9649 19119 9683 19153
rect 9717 19119 9751 19153
rect 9785 19119 9819 19153
rect 9853 19119 9887 19153
rect 9921 19119 9955 19153
rect 9989 19119 10023 19153
rect 10057 19119 10091 19153
rect 10125 19119 10159 19153
rect 10193 19119 10227 19153
rect 10261 19119 10295 19153
rect 10329 19119 10363 19153
rect 10397 19119 10431 19153
rect 10465 19119 10499 19153
rect 10533 19119 10567 19153
rect 10601 19119 10635 19153
rect 10669 19119 10703 19153
rect 10737 19119 10771 19153
rect 10805 19119 10839 19153
rect 10873 19119 10907 19153
rect 10941 19119 10975 19153
rect 11009 19119 11043 19153
rect 11077 19119 11111 19153
rect 11145 19119 11179 19153
rect 11213 19119 11247 19153
rect 11281 19119 11315 19153
rect 11349 19119 11383 19153
rect 11417 19119 11451 19153
rect 11485 19119 11519 19153
rect 11553 19119 11587 19153
rect 11621 19119 11655 19153
rect 11689 19119 11723 19153
rect 77 19047 111 19081
rect 146 19047 180 19081
rect 215 19047 249 19081
rect 284 19047 318 19081
rect 353 19047 387 19081
rect 422 19047 456 19081
rect 491 19047 525 19081
rect 560 19047 594 19081
rect 629 19047 663 19081
rect 698 19047 732 19081
rect 767 19047 801 19081
rect 836 19047 870 19081
rect 905 19047 939 19081
rect 974 19047 1008 19081
rect 1043 19047 1077 19081
rect 1112 19047 1146 19081
rect 1181 19047 1215 19081
rect 1250 19047 1284 19081
rect 1319 19047 1353 19081
rect 1388 19047 1422 19081
rect 1457 19047 1491 19081
rect 1526 19047 1560 19081
rect 1595 19047 1629 19081
rect 1664 19047 1698 19081
rect 1733 19047 1767 19081
rect 1802 19047 1836 19081
rect 1871 19047 1905 19081
rect 1940 19047 1974 19081
rect 2009 19047 2043 19081
rect 2078 19047 2112 19081
rect 2147 19047 2181 19081
rect 2216 19047 2250 19081
rect 2285 19047 2319 19081
rect 2354 19047 2388 19081
rect 2423 19047 2457 19081
rect 2492 19047 2526 19081
rect 2561 19047 2595 19081
rect 2630 19047 2664 19081
rect 2699 19047 2733 19081
rect 2768 19047 2802 19081
rect 2837 19047 2871 19081
rect 2906 19047 2940 19081
rect 2975 19047 3009 19081
rect 3044 19047 3078 19081
rect 3113 19047 3147 19081
rect 3182 19047 3216 19081
rect 3251 19047 3285 19081
rect 3320 19047 3354 19081
rect 3389 19047 3423 19081
rect 3458 19047 3492 19081
rect 3527 19047 3561 19081
rect 3596 19047 3630 19081
rect 3665 19047 3699 19081
rect 3733 19047 3767 19081
rect 3801 19047 3835 19081
rect 3869 19047 3903 19081
rect 3937 19047 3971 19081
rect 4005 19047 4039 19081
rect 4073 19047 4107 19081
rect 4141 19047 4175 19081
rect 4209 19047 4243 19081
rect 4277 19047 4311 19081
rect 4345 19047 4379 19081
rect 4413 19047 4447 19081
rect 4481 19047 4515 19081
rect 4549 19047 4583 19081
rect 4617 19047 4651 19081
rect 4685 19047 4719 19081
rect 4753 19047 4787 19081
rect 4821 19047 4855 19081
rect 4889 19047 4923 19081
rect 4957 19047 4991 19081
rect 5025 19047 5059 19081
rect 5093 19047 5127 19081
rect 5161 19047 5195 19081
rect 5229 19047 5263 19081
rect 5297 19047 5331 19081
rect 5365 19047 5399 19081
rect 5433 19047 5467 19081
rect 5501 19047 5535 19081
rect 5569 19047 5603 19081
rect 5637 19047 5671 19081
rect 5705 19047 5739 19081
rect 5773 19047 5807 19081
rect 5841 19047 5875 19081
rect 5909 19047 5943 19081
rect 5977 19047 6011 19081
rect 6045 19047 6079 19081
rect 6113 19047 6147 19081
rect 6181 19047 6215 19081
rect 6249 19047 6283 19081
rect 6317 19047 6351 19081
rect 6385 19047 6419 19081
rect 6453 19047 6487 19081
rect 6521 19047 6555 19081
rect 6589 19047 6623 19081
rect 6657 19047 6691 19081
rect 6725 19047 6759 19081
rect 6793 19047 6827 19081
rect 6861 19047 6895 19081
rect 6929 19047 6963 19081
rect 6997 19047 7031 19081
rect 7065 19047 7099 19081
rect 7133 19047 7167 19081
rect 7201 19047 7235 19081
rect 7269 19047 7303 19081
rect 7337 19047 7371 19081
rect 7405 19047 7439 19081
rect 7473 19047 7507 19081
rect 7541 19047 7575 19081
rect 7609 19047 7643 19081
rect 7677 19047 7711 19081
rect 7745 19047 7779 19081
rect 7813 19047 7847 19081
rect 7881 19047 7915 19081
rect 7949 19047 7983 19081
rect 8017 19047 8051 19081
rect 8085 19047 8119 19081
rect 8153 19047 8187 19081
rect 8221 19047 8255 19081
rect 8289 19047 8323 19081
rect 8357 19047 8391 19081
rect 8425 19047 8459 19081
rect 8493 19047 8527 19081
rect 8561 19047 8595 19081
rect 8629 19047 8663 19081
rect 8697 19047 8731 19081
rect 8765 19047 8799 19081
rect 8833 19047 8867 19081
rect 8901 19047 8935 19081
rect 8969 19047 9003 19081
rect 9037 19047 9071 19081
rect 9105 19047 9139 19081
rect 9173 19047 9207 19081
rect 9241 19047 9275 19081
rect 9309 19047 9343 19081
rect 9377 19047 9411 19081
rect 9445 19047 9479 19081
rect 9513 19047 9547 19081
rect 9581 19047 9615 19081
rect 9649 19047 9683 19081
rect 9717 19047 9751 19081
rect 9785 19047 9819 19081
rect 9853 19047 9887 19081
rect 9921 19047 9955 19081
rect 9989 19047 10023 19081
rect 10057 19047 10091 19081
rect 10125 19047 10159 19081
rect 10193 19047 10227 19081
rect 10261 19047 10295 19081
rect 10329 19047 10363 19081
rect 10397 19047 10431 19081
rect 10465 19047 10499 19081
rect 10533 19047 10567 19081
rect 10601 19047 10635 19081
rect 10669 19047 10703 19081
rect 10737 19047 10771 19081
rect 10805 19047 10839 19081
rect 10873 19047 10907 19081
rect 10941 19047 10975 19081
rect 11009 19047 11043 19081
rect 11077 19047 11111 19081
rect 11145 19047 11179 19081
rect 11213 19047 11247 19081
rect 11281 19047 11315 19081
rect 11349 19047 11383 19081
rect 11417 19047 11451 19081
rect 11485 19047 11519 19081
rect 11553 19047 11587 19081
rect 11621 19047 11655 19081
rect 11689 19047 11723 19081
rect 77 18975 111 19009
rect 146 18975 180 19009
rect 215 18975 249 19009
rect 284 18975 318 19009
rect 353 18975 387 19009
rect 422 18975 456 19009
rect 491 18975 525 19009
rect 560 18975 594 19009
rect 629 18975 663 19009
rect 698 18975 732 19009
rect 767 18975 801 19009
rect 836 18975 870 19009
rect 905 18975 939 19009
rect 974 18975 1008 19009
rect 1043 18975 1077 19009
rect 1112 18975 1146 19009
rect 1181 18975 1215 19009
rect 1250 18975 1284 19009
rect 1319 18975 1353 19009
rect 1388 18975 1422 19009
rect 1457 18975 1491 19009
rect 1526 18975 1560 19009
rect 1595 18975 1629 19009
rect 1664 18975 1698 19009
rect 1733 18975 1767 19009
rect 1802 18975 1836 19009
rect 1871 18975 1905 19009
rect 1940 18975 1974 19009
rect 2009 18975 2043 19009
rect 2078 18975 2112 19009
rect 2147 18975 2181 19009
rect 2216 18975 2250 19009
rect 2285 18975 2319 19009
rect 2354 18975 2388 19009
rect 2423 18975 2457 19009
rect 2492 18975 2526 19009
rect 2561 18975 2595 19009
rect 2630 18975 2664 19009
rect 2699 18975 2733 19009
rect 2768 18975 2802 19009
rect 2837 18975 2871 19009
rect 2906 18975 2940 19009
rect 2975 18975 3009 19009
rect 3044 18975 3078 19009
rect 3113 18975 3147 19009
rect 3182 18975 3216 19009
rect 3251 18975 3285 19009
rect 3320 18975 3354 19009
rect 3389 18975 3423 19009
rect 3458 18975 3492 19009
rect 3527 18975 3561 19009
rect 3596 18975 3630 19009
rect 3665 18975 3699 19009
rect 3733 18975 3767 19009
rect 3801 18975 3835 19009
rect 3869 18975 3903 19009
rect 3937 18975 3971 19009
rect 4005 18975 4039 19009
rect 4073 18975 4107 19009
rect 4141 18975 4175 19009
rect 4209 18975 4243 19009
rect 4277 18975 4311 19009
rect 4345 18975 4379 19009
rect 4413 18975 4447 19009
rect 4481 18975 4515 19009
rect 4549 18975 4583 19009
rect 4617 18975 4651 19009
rect 4685 18975 4719 19009
rect 4753 18975 4787 19009
rect 4821 18975 4855 19009
rect 4889 18975 4923 19009
rect 4957 18975 4991 19009
rect 5025 18975 5059 19009
rect 5093 18975 5127 19009
rect 5161 18975 5195 19009
rect 5229 18975 5263 19009
rect 5297 18975 5331 19009
rect 5365 18975 5399 19009
rect 5433 18975 5467 19009
rect 5501 18975 5535 19009
rect 5569 18975 5603 19009
rect 5637 18975 5671 19009
rect 5705 18975 5739 19009
rect 5773 18975 5807 19009
rect 5841 18975 5875 19009
rect 5909 18975 5943 19009
rect 5977 18975 6011 19009
rect 6045 18975 6079 19009
rect 6113 18975 6147 19009
rect 6181 18975 6215 19009
rect 6249 18975 6283 19009
rect 6317 18975 6351 19009
rect 6385 18975 6419 19009
rect 6453 18975 6487 19009
rect 6521 18975 6555 19009
rect 6589 18975 6623 19009
rect 6657 18975 6691 19009
rect 6725 18975 6759 19009
rect 6793 18975 6827 19009
rect 6861 18975 6895 19009
rect 6929 18975 6963 19009
rect 6997 18975 7031 19009
rect 7065 18975 7099 19009
rect 7133 18975 7167 19009
rect 7201 18975 7235 19009
rect 7269 18975 7303 19009
rect 7337 18975 7371 19009
rect 7405 18975 7439 19009
rect 7473 18975 7507 19009
rect 7541 18975 7575 19009
rect 7609 18975 7643 19009
rect 7677 18975 7711 19009
rect 7745 18975 7779 19009
rect 7813 18975 7847 19009
rect 7881 18975 7915 19009
rect 7949 18975 7983 19009
rect 8017 18975 8051 19009
rect 8085 18975 8119 19009
rect 8153 18975 8187 19009
rect 8221 18975 8255 19009
rect 8289 18975 8323 19009
rect 8357 18975 8391 19009
rect 8425 18975 8459 19009
rect 8493 18975 8527 19009
rect 8561 18975 8595 19009
rect 8629 18975 8663 19009
rect 8697 18975 8731 19009
rect 8765 18975 8799 19009
rect 8833 18975 8867 19009
rect 8901 18975 8935 19009
rect 8969 18975 9003 19009
rect 9037 18975 9071 19009
rect 9105 18975 9139 19009
rect 9173 18975 9207 19009
rect 9241 18975 9275 19009
rect 9309 18975 9343 19009
rect 9377 18975 9411 19009
rect 9445 18975 9479 19009
rect 9513 18975 9547 19009
rect 9581 18975 9615 19009
rect 9649 18975 9683 19009
rect 9717 18975 9751 19009
rect 9785 18975 9819 19009
rect 9853 18975 9887 19009
rect 9921 18975 9955 19009
rect 9989 18975 10023 19009
rect 10057 18975 10091 19009
rect 10125 18975 10159 19009
rect 10193 18975 10227 19009
rect 10261 18975 10295 19009
rect 10329 18975 10363 19009
rect 10397 18975 10431 19009
rect 10465 18975 10499 19009
rect 10533 18975 10567 19009
rect 10601 18975 10635 19009
rect 10669 18975 10703 19009
rect 10737 18975 10771 19009
rect 10805 18975 10839 19009
rect 10873 18975 10907 19009
rect 10941 18975 10975 19009
rect 11009 18975 11043 19009
rect 11077 18975 11111 19009
rect 11145 18975 11179 19009
rect 11213 18975 11247 19009
rect 11281 18975 11315 19009
rect 11349 18975 11383 19009
rect 11417 18975 11451 19009
rect 11485 18975 11519 19009
rect 11553 18975 11587 19009
rect 11621 18975 11655 19009
rect 11689 18975 11723 19009
rect 14484 19307 14518 19341
rect 14567 19307 14601 19341
rect 14650 19307 14684 19341
rect 14733 19307 14767 19341
rect 14816 19307 14850 19341
rect 14484 19237 14518 19271
rect 14567 19237 14601 19271
rect 14650 19237 14684 19271
rect 14733 19237 14767 19271
rect 14816 19237 14850 19271
rect 14484 19167 14518 19201
rect 14567 19167 14601 19201
rect 14650 19167 14684 19201
rect 14733 19167 14767 19201
rect 14816 19167 14850 19201
rect 14484 19097 14518 19131
rect 14567 19097 14601 19131
rect 14650 19097 14684 19131
rect 14733 19097 14767 19131
rect 14816 19097 14850 19131
rect 14484 19027 14518 19061
rect 14567 19027 14601 19061
rect 14650 19027 14684 19061
rect 14733 19027 14767 19061
rect 14816 19027 14850 19061
rect 77 18881 111 18915
rect 146 18881 180 18915
rect 215 18881 249 18915
rect 284 18881 318 18915
rect 353 18881 387 18915
rect 422 18881 456 18915
rect 491 18881 525 18915
rect 560 18881 594 18915
rect 629 18881 663 18915
rect 698 18881 732 18915
rect 767 18881 801 18915
rect 836 18881 870 18915
rect 905 18881 939 18915
rect 974 18881 1008 18915
rect 1043 18881 1077 18915
rect 1112 18881 1146 18915
rect 1181 18881 1215 18915
rect 1250 18881 1284 18915
rect 1319 18881 1353 18915
rect 1388 18881 1422 18915
rect 1457 18881 1491 18915
rect 1526 18881 1560 18915
rect 1595 18881 1629 18915
rect 1664 18881 1698 18915
rect 1733 18881 1767 18915
rect 1802 18881 1836 18915
rect 1871 18881 1905 18915
rect 1940 18881 1974 18915
rect 2009 18881 2043 18915
rect 2078 18881 2112 18915
rect 2147 18881 2181 18915
rect 2216 18881 2250 18915
rect 2285 18881 2319 18915
rect 2354 18881 2388 18915
rect 2423 18881 2457 18915
rect 2492 18881 2526 18915
rect 2561 18881 2595 18915
rect 2630 18881 2664 18915
rect 2699 18881 2733 18915
rect 2768 18881 2802 18915
rect 2837 18881 2871 18915
rect 2906 18881 2940 18915
rect 2975 18881 3009 18915
rect 3044 18881 3078 18915
rect 3113 18881 3147 18915
rect 3182 18881 3216 18915
rect 3251 18881 3285 18915
rect 3320 18881 3354 18915
rect 3389 18881 3423 18915
rect 3458 18881 3492 18915
rect 3527 18881 3561 18915
rect 77 18813 111 18847
rect 146 18813 180 18847
rect 215 18813 249 18847
rect 284 18813 318 18847
rect 353 18813 387 18847
rect 422 18813 456 18847
rect 491 18813 525 18847
rect 560 18813 594 18847
rect 629 18813 663 18847
rect 698 18813 732 18847
rect 767 18813 801 18847
rect 836 18813 870 18847
rect 905 18813 939 18847
rect 974 18813 1008 18847
rect 1043 18813 1077 18847
rect 1112 18813 1146 18847
rect 1181 18813 1215 18847
rect 1250 18813 1284 18847
rect 1319 18813 1353 18847
rect 1388 18813 1422 18847
rect 1457 18813 1491 18847
rect 1526 18813 1560 18847
rect 1595 18813 1629 18847
rect 1664 18813 1698 18847
rect 1733 18813 1767 18847
rect 1802 18813 1836 18847
rect 1871 18813 1905 18847
rect 1940 18813 1974 18847
rect 2009 18813 2043 18847
rect 2078 18813 2112 18847
rect 2147 18813 2181 18847
rect 2216 18813 2250 18847
rect 2285 18813 2319 18847
rect 2354 18813 2388 18847
rect 2423 18813 2457 18847
rect 2492 18813 2526 18847
rect 2561 18813 2595 18847
rect 2630 18813 2664 18847
rect 2699 18813 2733 18847
rect 2768 18813 2802 18847
rect 2837 18813 2871 18847
rect 2906 18813 2940 18847
rect 2975 18813 3009 18847
rect 3044 18813 3078 18847
rect 3113 18813 3147 18847
rect 3182 18813 3216 18847
rect 3251 18813 3285 18847
rect 3320 18813 3354 18847
rect 3389 18813 3423 18847
rect 3458 18813 3492 18847
rect 3527 18813 3561 18847
rect 77 18745 111 18779
rect 146 18745 180 18779
rect 215 18745 249 18779
rect 284 18745 318 18779
rect 353 18745 387 18779
rect 422 18745 456 18779
rect 491 18745 525 18779
rect 560 18745 594 18779
rect 629 18745 663 18779
rect 698 18745 732 18779
rect 767 18745 801 18779
rect 836 18745 870 18779
rect 905 18745 939 18779
rect 974 18745 1008 18779
rect 1043 18745 1077 18779
rect 1112 18745 1146 18779
rect 1181 18745 1215 18779
rect 1250 18745 1284 18779
rect 1319 18745 1353 18779
rect 1388 18745 1422 18779
rect 1457 18745 1491 18779
rect 1526 18745 1560 18779
rect 1595 18745 1629 18779
rect 1664 18745 1698 18779
rect 1733 18745 1767 18779
rect 1802 18745 1836 18779
rect 1871 18745 1905 18779
rect 1940 18745 1974 18779
rect 2009 18745 2043 18779
rect 2078 18745 2112 18779
rect 2147 18745 2181 18779
rect 2216 18745 2250 18779
rect 2285 18745 2319 18779
rect 2354 18745 2388 18779
rect 2423 18745 2457 18779
rect 2492 18745 2526 18779
rect 2561 18745 2595 18779
rect 2630 18745 2664 18779
rect 2699 18745 2733 18779
rect 2768 18745 2802 18779
rect 2837 18745 2871 18779
rect 2906 18745 2940 18779
rect 2975 18745 3009 18779
rect 3044 18745 3078 18779
rect 3113 18745 3147 18779
rect 3182 18745 3216 18779
rect 3251 18745 3285 18779
rect 3320 18745 3354 18779
rect 3389 18745 3423 18779
rect 3458 18745 3492 18779
rect 3527 18745 3561 18779
rect 77 18677 111 18711
rect 146 18677 180 18711
rect 215 18677 249 18711
rect 284 18677 318 18711
rect 353 18677 387 18711
rect 422 18677 456 18711
rect 491 18677 525 18711
rect 560 18677 594 18711
rect 629 18677 663 18711
rect 698 18677 732 18711
rect 767 18677 801 18711
rect 836 18677 870 18711
rect 905 18677 939 18711
rect 974 18677 1008 18711
rect 1043 18677 1077 18711
rect 1112 18677 1146 18711
rect 1181 18677 1215 18711
rect 1250 18677 1284 18711
rect 1319 18677 1353 18711
rect 1388 18677 1422 18711
rect 1457 18677 1491 18711
rect 1526 18677 1560 18711
rect 1595 18677 1629 18711
rect 1664 18677 1698 18711
rect 1733 18677 1767 18711
rect 1802 18677 1836 18711
rect 1871 18677 1905 18711
rect 1940 18677 1974 18711
rect 2009 18677 2043 18711
rect 2078 18677 2112 18711
rect 2147 18677 2181 18711
rect 2216 18677 2250 18711
rect 2285 18677 2319 18711
rect 2354 18677 2388 18711
rect 2423 18677 2457 18711
rect 2492 18677 2526 18711
rect 2561 18677 2595 18711
rect 2630 18677 2664 18711
rect 2699 18677 2733 18711
rect 2768 18677 2802 18711
rect 2837 18677 2871 18711
rect 2906 18677 2940 18711
rect 2975 18677 3009 18711
rect 3044 18677 3078 18711
rect 3113 18677 3147 18711
rect 3182 18677 3216 18711
rect 3251 18677 3285 18711
rect 3320 18677 3354 18711
rect 3389 18677 3423 18711
rect 3458 18677 3492 18711
rect 3527 18677 3561 18711
rect 3596 18677 14850 18915
rect 221 18555 255 18589
rect 290 18555 324 18589
rect 359 18555 393 18589
rect 427 18555 461 18589
rect 495 18555 529 18589
rect 563 18555 597 18589
rect 631 18555 665 18589
rect 699 18555 733 18589
rect 767 18555 801 18589
rect 835 18555 869 18589
rect 903 18555 937 18589
rect 971 18555 1005 18589
rect 1039 18555 1073 18589
rect 1107 18555 1141 18589
rect 1175 18555 1209 18589
rect 1243 18555 1277 18589
rect 1311 18555 1345 18589
rect 1379 18555 1413 18589
rect 1447 18555 1481 18589
rect 1515 18555 1549 18589
rect 1583 18555 1617 18589
rect 1651 18555 1685 18589
rect 1719 18555 1753 18589
rect 1787 18555 1821 18589
rect 1855 18555 1889 18589
rect 1923 18555 1957 18589
rect 1991 18555 2025 18589
rect 2059 18555 2093 18589
rect 2127 18555 2161 18589
rect 2195 18555 2229 18589
rect 2263 18555 2297 18589
rect 2331 18555 2365 18589
rect 2399 18555 2433 18589
rect 2467 18555 2501 18589
rect 2535 18555 2569 18589
rect 2603 18555 2637 18589
rect 2671 18555 2705 18589
rect 2739 18555 2773 18589
rect 2807 18555 2841 18589
rect 2875 18555 2909 18589
rect 2943 18555 2977 18589
rect 3011 18555 3045 18589
rect 3079 18555 3113 18589
rect 3147 18555 3181 18589
rect 3215 18555 3249 18589
rect 3283 18555 3317 18589
rect 3351 18555 3385 18589
rect 3419 18555 3453 18589
rect 3487 18555 3521 18589
rect 3555 18555 3589 18589
rect 3623 18555 3657 18589
rect 3691 18555 3725 18589
rect 3759 18555 3793 18589
rect 3827 18555 3861 18589
rect 3895 18555 3929 18589
rect 3963 18555 3997 18589
rect 4031 18555 4065 18589
rect 4099 18555 4133 18589
rect 4167 18555 4201 18589
rect 4235 18555 4269 18589
rect 4303 18555 4337 18589
rect 4371 18555 4405 18589
rect 4439 18555 4473 18589
rect 4507 18555 4541 18589
rect 4575 18555 4609 18589
rect 4643 18555 4677 18589
rect 4711 18555 4745 18589
rect 4779 18555 4813 18589
rect 4847 18555 4881 18589
rect 4915 18555 4949 18589
rect 4983 18555 5017 18589
rect 5051 18555 5085 18589
rect 5119 18555 5153 18589
rect 5187 18555 5221 18589
rect 5255 18555 5289 18589
rect 5323 18555 5357 18589
rect 5391 18555 5425 18589
rect 5459 18555 5493 18589
rect 5527 18555 5561 18589
rect 5595 18555 5629 18589
rect 5663 18555 5697 18589
rect 5731 18555 5765 18589
rect 5799 18555 5833 18589
rect 5867 18555 5901 18589
rect 5935 18555 5969 18589
rect 6003 18555 6037 18589
rect 6071 18555 6105 18589
rect 6139 18555 6173 18589
rect 6207 18555 6241 18589
rect 6275 18555 6309 18589
rect 6343 18555 6377 18589
rect 6411 18555 6445 18589
rect 6479 18555 6513 18589
rect 6547 18555 6581 18589
rect 6615 18555 6649 18589
rect 6683 18555 6717 18589
rect 6751 18555 6785 18589
rect 6819 18555 6853 18589
rect 6887 18555 6921 18589
rect 6955 18555 6989 18589
rect 7023 18555 7057 18589
rect 7091 18555 7125 18589
rect 7159 18555 7193 18589
rect 7227 18555 7261 18589
rect 7295 18555 7329 18589
rect 7363 18555 7397 18589
rect 7431 18555 7465 18589
rect 7499 18555 7533 18589
rect 7567 18555 7601 18589
rect 7635 18555 7669 18589
rect 7703 18555 7737 18589
rect 7771 18555 7805 18589
rect 7839 18555 7873 18589
rect 7907 18555 7941 18589
rect 7975 18555 8009 18589
rect 8043 18555 8077 18589
rect 8111 18555 8145 18589
rect 8179 18555 8213 18589
rect 8247 18555 8281 18589
rect 8315 18555 8349 18589
rect 8383 18555 8417 18589
rect 8451 18555 8485 18589
rect 8519 18555 8553 18589
rect 8587 18555 8621 18589
rect 8655 18555 8689 18589
rect 8723 18555 8757 18589
rect 8791 18555 8825 18589
rect 8859 18555 8893 18589
rect 8927 18555 8961 18589
rect 8995 18555 9029 18589
rect 9063 18555 9097 18589
rect 9131 18555 9165 18589
rect 9199 18555 9233 18589
rect 9267 18555 9301 18589
rect 9335 18555 9369 18589
rect 9403 18555 9437 18589
rect 9471 18555 9505 18589
rect 9539 18555 9573 18589
rect 9607 18555 9641 18589
rect 9675 18555 9709 18589
rect 9743 18555 9777 18589
rect 9811 18555 9845 18589
rect 9879 18555 9913 18589
rect 9947 18555 9981 18589
rect 10015 18555 10049 18589
rect 10083 18555 10117 18589
rect 10151 18555 10185 18589
rect 10219 18555 10253 18589
rect 10287 18555 10321 18589
rect 10355 18555 10389 18589
rect 10423 18555 10457 18589
rect 10491 18555 10525 18589
rect 10559 18555 10593 18589
rect 10627 18555 10661 18589
rect 10695 18555 10729 18589
rect 10763 18555 10797 18589
rect 10831 18555 10865 18589
rect 10899 18555 10933 18589
rect 10967 18555 11001 18589
rect 11035 18555 11069 18589
rect 11103 18555 11137 18589
rect 11171 18555 11205 18589
rect 11239 18555 11273 18589
rect 11307 18555 11341 18589
rect 11375 18555 11409 18589
rect 11443 18555 11477 18589
rect 11511 18555 11545 18589
rect 11579 18555 11613 18589
rect 11647 18555 11681 18589
rect 11715 18555 11749 18589
rect 11783 18555 11817 18589
rect 11851 18555 11885 18589
rect 11919 18555 11953 18589
rect 11987 18555 12021 18589
rect 12055 18555 12089 18589
rect 12123 18555 12157 18589
rect 12191 18555 12225 18589
rect 12259 18555 12293 18589
rect 12327 18555 12361 18589
rect 12395 18555 12429 18589
rect 12463 18555 12497 18589
rect 12531 18555 12565 18589
rect 12599 18555 12633 18589
rect 12667 18555 12701 18589
rect 12735 18555 12769 18589
rect 12803 18555 12837 18589
rect 12871 18555 12905 18589
rect 12939 18555 12973 18589
rect 13007 18555 13041 18589
rect 13075 18555 13109 18589
rect 13143 18555 13177 18589
rect 13211 18555 13245 18589
rect 13279 18555 13313 18589
rect 13347 18555 13381 18589
rect 13415 18555 13449 18589
rect 13483 18555 13517 18589
rect 13551 18555 13585 18589
rect 13619 18555 13653 18589
rect 13687 18555 13721 18589
rect 13755 18555 13789 18589
rect 13823 18555 13857 18589
rect 13891 18555 13925 18589
rect 13959 18555 13993 18589
rect 14027 18555 14061 18589
rect 14095 18555 14129 18589
rect 14163 18555 14197 18589
rect 14231 18555 14265 18589
rect 14299 18555 14333 18589
rect 14367 18555 14401 18589
rect 14435 18555 14469 18589
rect 14503 18555 14537 18589
rect 14571 18555 14605 18589
rect 14639 18555 14673 18589
rect 14707 18555 14741 18589
rect 221 18485 255 18519
rect 290 18485 324 18519
rect 359 18485 393 18519
rect 427 18485 461 18519
rect 495 18485 529 18519
rect 563 18485 597 18519
rect 631 18485 665 18519
rect 699 18485 733 18519
rect 767 18485 801 18519
rect 835 18485 869 18519
rect 903 18485 937 18519
rect 971 18485 1005 18519
rect 1039 18485 1073 18519
rect 1107 18485 1141 18519
rect 1175 18485 1209 18519
rect 1243 18485 1277 18519
rect 1311 18485 1345 18519
rect 1379 18485 1413 18519
rect 1447 18485 1481 18519
rect 1515 18485 1549 18519
rect 1583 18485 1617 18519
rect 1651 18485 1685 18519
rect 1719 18485 1753 18519
rect 1787 18485 1821 18519
rect 1855 18485 1889 18519
rect 1923 18485 1957 18519
rect 1991 18485 2025 18519
rect 2059 18485 2093 18519
rect 2127 18485 2161 18519
rect 2195 18485 2229 18519
rect 2263 18485 2297 18519
rect 2331 18485 2365 18519
rect 2399 18485 2433 18519
rect 2467 18485 2501 18519
rect 2535 18485 2569 18519
rect 2603 18485 2637 18519
rect 2671 18485 2705 18519
rect 2739 18485 2773 18519
rect 2807 18485 2841 18519
rect 2875 18485 2909 18519
rect 2943 18485 2977 18519
rect 3011 18485 3045 18519
rect 3079 18485 3113 18519
rect 3147 18485 3181 18519
rect 3215 18485 3249 18519
rect 3283 18485 3317 18519
rect 3351 18485 3385 18519
rect 3419 18485 3453 18519
rect 3487 18485 3521 18519
rect 3555 18485 3589 18519
rect 3623 18485 3657 18519
rect 3691 18485 3725 18519
rect 3759 18485 3793 18519
rect 3827 18485 3861 18519
rect 3895 18485 3929 18519
rect 3963 18485 3997 18519
rect 4031 18485 4065 18519
rect 4099 18485 4133 18519
rect 4167 18485 4201 18519
rect 4235 18485 4269 18519
rect 4303 18485 4337 18519
rect 4371 18485 4405 18519
rect 4439 18485 4473 18519
rect 4507 18485 4541 18519
rect 4575 18485 4609 18519
rect 4643 18485 4677 18519
rect 4711 18485 4745 18519
rect 4779 18485 4813 18519
rect 4847 18485 4881 18519
rect 4915 18485 4949 18519
rect 4983 18485 5017 18519
rect 5051 18485 5085 18519
rect 5119 18485 5153 18519
rect 5187 18485 5221 18519
rect 5255 18485 5289 18519
rect 5323 18485 5357 18519
rect 5391 18485 5425 18519
rect 5459 18485 5493 18519
rect 5527 18485 5561 18519
rect 5595 18485 5629 18519
rect 5663 18485 5697 18519
rect 5731 18485 5765 18519
rect 5799 18485 5833 18519
rect 5867 18485 5901 18519
rect 5935 18485 5969 18519
rect 6003 18485 6037 18519
rect 6071 18485 6105 18519
rect 6139 18485 6173 18519
rect 6207 18485 6241 18519
rect 6275 18485 6309 18519
rect 6343 18485 6377 18519
rect 6411 18485 6445 18519
rect 6479 18485 6513 18519
rect 6547 18485 6581 18519
rect 6615 18485 6649 18519
rect 6683 18485 6717 18519
rect 6751 18485 6785 18519
rect 6819 18485 6853 18519
rect 6887 18485 6921 18519
rect 6955 18485 6989 18519
rect 7023 18485 7057 18519
rect 7091 18485 7125 18519
rect 7159 18485 7193 18519
rect 7227 18485 7261 18519
rect 7295 18485 7329 18519
rect 7363 18485 7397 18519
rect 7431 18485 7465 18519
rect 7499 18485 7533 18519
rect 7567 18485 7601 18519
rect 7635 18485 7669 18519
rect 7703 18485 7737 18519
rect 7771 18485 7805 18519
rect 7839 18485 7873 18519
rect 7907 18485 7941 18519
rect 7975 18485 8009 18519
rect 8043 18485 8077 18519
rect 8111 18485 8145 18519
rect 8179 18485 8213 18519
rect 8247 18485 8281 18519
rect 8315 18485 8349 18519
rect 8383 18485 8417 18519
rect 8451 18485 8485 18519
rect 8519 18485 8553 18519
rect 8587 18485 8621 18519
rect 8655 18485 8689 18519
rect 8723 18485 8757 18519
rect 8791 18485 8825 18519
rect 8859 18485 8893 18519
rect 8927 18485 8961 18519
rect 8995 18485 9029 18519
rect 9063 18485 9097 18519
rect 9131 18485 9165 18519
rect 9199 18485 9233 18519
rect 9267 18485 9301 18519
rect 9335 18485 9369 18519
rect 9403 18485 9437 18519
rect 9471 18485 9505 18519
rect 9539 18485 9573 18519
rect 9607 18485 9641 18519
rect 9675 18485 9709 18519
rect 9743 18485 9777 18519
rect 9811 18485 9845 18519
rect 9879 18485 9913 18519
rect 9947 18485 9981 18519
rect 10015 18485 10049 18519
rect 10083 18485 10117 18519
rect 10151 18485 10185 18519
rect 10219 18485 10253 18519
rect 10287 18485 10321 18519
rect 10355 18485 10389 18519
rect 10423 18485 10457 18519
rect 10491 18485 10525 18519
rect 10559 18485 10593 18519
rect 10627 18485 10661 18519
rect 10695 18485 10729 18519
rect 10763 18485 10797 18519
rect 10831 18485 10865 18519
rect 10899 18485 10933 18519
rect 10967 18485 11001 18519
rect 11035 18485 11069 18519
rect 11103 18485 11137 18519
rect 11171 18485 11205 18519
rect 11239 18485 11273 18519
rect 11307 18485 11341 18519
rect 11375 18485 11409 18519
rect 11443 18485 11477 18519
rect 11511 18485 11545 18519
rect 11579 18485 11613 18519
rect 11647 18485 11681 18519
rect 11715 18485 11749 18519
rect 11783 18485 11817 18519
rect 11851 18485 11885 18519
rect 11919 18485 11953 18519
rect 11987 18485 12021 18519
rect 12055 18485 12089 18519
rect 12123 18485 12157 18519
rect 12191 18485 12225 18519
rect 12259 18485 12293 18519
rect 12327 18485 12361 18519
rect 12395 18485 12429 18519
rect 12463 18485 12497 18519
rect 12531 18485 12565 18519
rect 12599 18485 12633 18519
rect 12667 18485 12701 18519
rect 12735 18485 12769 18519
rect 12803 18485 12837 18519
rect 12871 18485 12905 18519
rect 12939 18485 12973 18519
rect 13007 18485 13041 18519
rect 13075 18485 13109 18519
rect 13143 18485 13177 18519
rect 13211 18485 13245 18519
rect 13279 18485 13313 18519
rect 13347 18485 13381 18519
rect 13415 18485 13449 18519
rect 13483 18485 13517 18519
rect 13551 18485 13585 18519
rect 13619 18485 13653 18519
rect 13687 18485 13721 18519
rect 13755 18485 13789 18519
rect 13823 18485 13857 18519
rect 13891 18485 13925 18519
rect 13959 18485 13993 18519
rect 14027 18485 14061 18519
rect 14095 18485 14129 18519
rect 14163 18485 14197 18519
rect 14231 18485 14265 18519
rect 14299 18485 14333 18519
rect 14367 18485 14401 18519
rect 14435 18485 14469 18519
rect 14503 18485 14537 18519
rect 14571 18485 14605 18519
rect 14639 18485 14673 18519
rect 14707 18485 14741 18519
rect 221 18415 255 18449
rect 290 18415 324 18449
rect 359 18415 393 18449
rect 427 18415 461 18449
rect 495 18415 529 18449
rect 563 18415 597 18449
rect 631 18415 665 18449
rect 699 18415 733 18449
rect 767 18415 801 18449
rect 835 18415 869 18449
rect 903 18415 937 18449
rect 971 18415 1005 18449
rect 1039 18415 1073 18449
rect 1107 18415 1141 18449
rect 1175 18415 1209 18449
rect 1243 18415 1277 18449
rect 1311 18415 1345 18449
rect 1379 18415 1413 18449
rect 1447 18415 1481 18449
rect 1515 18415 1549 18449
rect 1583 18415 1617 18449
rect 1651 18415 1685 18449
rect 1719 18415 1753 18449
rect 1787 18415 1821 18449
rect 1855 18415 1889 18449
rect 1923 18415 1957 18449
rect 1991 18415 2025 18449
rect 2059 18415 2093 18449
rect 2127 18415 2161 18449
rect 2195 18415 2229 18449
rect 2263 18415 2297 18449
rect 2331 18415 2365 18449
rect 2399 18415 2433 18449
rect 2467 18415 2501 18449
rect 2535 18415 2569 18449
rect 2603 18415 2637 18449
rect 2671 18415 2705 18449
rect 2739 18415 2773 18449
rect 2807 18415 2841 18449
rect 2875 18415 2909 18449
rect 2943 18415 2977 18449
rect 3011 18415 3045 18449
rect 3079 18415 3113 18449
rect 3147 18415 3181 18449
rect 3215 18415 3249 18449
rect 3283 18415 3317 18449
rect 3351 18415 3385 18449
rect 3419 18415 3453 18449
rect 3487 18415 3521 18449
rect 3555 18415 3589 18449
rect 3623 18415 3657 18449
rect 3691 18415 3725 18449
rect 3759 18415 3793 18449
rect 3827 18415 3861 18449
rect 3895 18415 3929 18449
rect 3963 18415 3997 18449
rect 4031 18415 4065 18449
rect 4099 18415 4133 18449
rect 4167 18415 4201 18449
rect 4235 18415 4269 18449
rect 4303 18415 4337 18449
rect 4371 18415 4405 18449
rect 4439 18415 4473 18449
rect 4507 18415 4541 18449
rect 4575 18415 4609 18449
rect 4643 18415 4677 18449
rect 4711 18415 4745 18449
rect 4779 18415 4813 18449
rect 4847 18415 4881 18449
rect 4915 18415 4949 18449
rect 4983 18415 5017 18449
rect 5051 18415 5085 18449
rect 5119 18415 5153 18449
rect 5187 18415 5221 18449
rect 5255 18415 5289 18449
rect 5323 18415 5357 18449
rect 5391 18415 5425 18449
rect 5459 18415 5493 18449
rect 5527 18415 5561 18449
rect 5595 18415 5629 18449
rect 5663 18415 5697 18449
rect 5731 18415 5765 18449
rect 5799 18415 5833 18449
rect 5867 18415 5901 18449
rect 5935 18415 5969 18449
rect 6003 18415 6037 18449
rect 6071 18415 6105 18449
rect 6139 18415 6173 18449
rect 6207 18415 6241 18449
rect 6275 18415 6309 18449
rect 6343 18415 6377 18449
rect 6411 18415 6445 18449
rect 6479 18415 6513 18449
rect 6547 18415 6581 18449
rect 6615 18415 6649 18449
rect 6683 18415 6717 18449
rect 6751 18415 6785 18449
rect 6819 18415 6853 18449
rect 6887 18415 6921 18449
rect 6955 18415 6989 18449
rect 7023 18415 7057 18449
rect 7091 18415 7125 18449
rect 7159 18415 7193 18449
rect 7227 18415 7261 18449
rect 7295 18415 7329 18449
rect 7363 18415 7397 18449
rect 7431 18415 7465 18449
rect 7499 18415 7533 18449
rect 7567 18415 7601 18449
rect 7635 18415 7669 18449
rect 7703 18415 7737 18449
rect 7771 18415 7805 18449
rect 7839 18415 7873 18449
rect 7907 18415 7941 18449
rect 7975 18415 8009 18449
rect 8043 18415 8077 18449
rect 8111 18415 8145 18449
rect 8179 18415 8213 18449
rect 8247 18415 8281 18449
rect 8315 18415 8349 18449
rect 8383 18415 8417 18449
rect 8451 18415 8485 18449
rect 8519 18415 8553 18449
rect 8587 18415 8621 18449
rect 8655 18415 8689 18449
rect 8723 18415 8757 18449
rect 8791 18415 8825 18449
rect 8859 18415 8893 18449
rect 8927 18415 8961 18449
rect 8995 18415 9029 18449
rect 9063 18415 9097 18449
rect 9131 18415 9165 18449
rect 9199 18415 9233 18449
rect 9267 18415 9301 18449
rect 9335 18415 9369 18449
rect 9403 18415 9437 18449
rect 9471 18415 9505 18449
rect 9539 18415 9573 18449
rect 9607 18415 9641 18449
rect 9675 18415 9709 18449
rect 9743 18415 9777 18449
rect 9811 18415 9845 18449
rect 9879 18415 9913 18449
rect 9947 18415 9981 18449
rect 10015 18415 10049 18449
rect 10083 18415 10117 18449
rect 10151 18415 10185 18449
rect 10219 18415 10253 18449
rect 10287 18415 10321 18449
rect 10355 18415 10389 18449
rect 10423 18415 10457 18449
rect 10491 18415 10525 18449
rect 10559 18415 10593 18449
rect 10627 18415 10661 18449
rect 10695 18415 10729 18449
rect 10763 18415 10797 18449
rect 10831 18415 10865 18449
rect 10899 18415 10933 18449
rect 10967 18415 11001 18449
rect 11035 18415 11069 18449
rect 11103 18415 11137 18449
rect 11171 18415 11205 18449
rect 11239 18415 11273 18449
rect 11307 18415 11341 18449
rect 11375 18415 11409 18449
rect 11443 18415 11477 18449
rect 11511 18415 11545 18449
rect 11579 18415 11613 18449
rect 11647 18415 11681 18449
rect 11715 18415 11749 18449
rect 11783 18415 11817 18449
rect 11851 18415 11885 18449
rect 11919 18415 11953 18449
rect 11987 18415 12021 18449
rect 12055 18415 12089 18449
rect 12123 18415 12157 18449
rect 12191 18415 12225 18449
rect 12259 18415 12293 18449
rect 12327 18415 12361 18449
rect 12395 18415 12429 18449
rect 12463 18415 12497 18449
rect 12531 18415 12565 18449
rect 12599 18415 12633 18449
rect 12667 18415 12701 18449
rect 12735 18415 12769 18449
rect 12803 18415 12837 18449
rect 12871 18415 12905 18449
rect 12939 18415 12973 18449
rect 13007 18415 13041 18449
rect 13075 18415 13109 18449
rect 13143 18415 13177 18449
rect 13211 18415 13245 18449
rect 13279 18415 13313 18449
rect 13347 18415 13381 18449
rect 13415 18415 13449 18449
rect 13483 18415 13517 18449
rect 13551 18415 13585 18449
rect 13619 18415 13653 18449
rect 13687 18415 13721 18449
rect 13755 18415 13789 18449
rect 13823 18415 13857 18449
rect 13891 18415 13925 18449
rect 13959 18415 13993 18449
rect 14027 18415 14061 18449
rect 14095 18415 14129 18449
rect 14163 18415 14197 18449
rect 14231 18415 14265 18449
rect 14299 18415 14333 18449
rect 14367 18415 14401 18449
rect 14435 18415 14469 18449
rect 14503 18415 14537 18449
rect 14571 18415 14605 18449
rect 14639 18415 14673 18449
rect 14707 18415 14741 18449
rect 221 18345 255 18379
rect 290 18345 324 18379
rect 359 18345 393 18379
rect 427 18345 461 18379
rect 495 18345 529 18379
rect 563 18345 597 18379
rect 631 18345 665 18379
rect 699 18345 733 18379
rect 767 18345 801 18379
rect 835 18345 869 18379
rect 903 18345 937 18379
rect 971 18345 1005 18379
rect 1039 18345 1073 18379
rect 1107 18345 1141 18379
rect 1175 18345 1209 18379
rect 1243 18345 1277 18379
rect 1311 18345 1345 18379
rect 1379 18345 1413 18379
rect 1447 18345 1481 18379
rect 1515 18345 1549 18379
rect 1583 18345 1617 18379
rect 1651 18345 1685 18379
rect 1719 18345 1753 18379
rect 1787 18345 1821 18379
rect 1855 18345 1889 18379
rect 1923 18345 1957 18379
rect 1991 18345 2025 18379
rect 2059 18345 2093 18379
rect 2127 18345 2161 18379
rect 2195 18345 2229 18379
rect 2263 18345 2297 18379
rect 2331 18345 2365 18379
rect 2399 18345 2433 18379
rect 2467 18345 2501 18379
rect 2535 18345 2569 18379
rect 2603 18345 2637 18379
rect 2671 18345 2705 18379
rect 2739 18345 2773 18379
rect 2807 18345 2841 18379
rect 2875 18345 2909 18379
rect 2943 18345 2977 18379
rect 3011 18345 3045 18379
rect 3079 18345 3113 18379
rect 3147 18345 3181 18379
rect 3215 18345 3249 18379
rect 3283 18345 3317 18379
rect 3351 18345 3385 18379
rect 3419 18345 3453 18379
rect 3487 18345 3521 18379
rect 3555 18345 3589 18379
rect 3623 18345 3657 18379
rect 3691 18345 3725 18379
rect 3759 18345 3793 18379
rect 3827 18345 3861 18379
rect 3895 18345 3929 18379
rect 3963 18345 3997 18379
rect 4031 18345 4065 18379
rect 4099 18345 4133 18379
rect 4167 18345 4201 18379
rect 4235 18345 4269 18379
rect 4303 18345 4337 18379
rect 4371 18345 4405 18379
rect 4439 18345 4473 18379
rect 4507 18345 4541 18379
rect 4575 18345 4609 18379
rect 4643 18345 4677 18379
rect 4711 18345 4745 18379
rect 4779 18345 4813 18379
rect 4847 18345 4881 18379
rect 4915 18345 4949 18379
rect 4983 18345 5017 18379
rect 5051 18345 5085 18379
rect 5119 18345 5153 18379
rect 5187 18345 5221 18379
rect 5255 18345 5289 18379
rect 5323 18345 5357 18379
rect 5391 18345 5425 18379
rect 5459 18345 5493 18379
rect 5527 18345 5561 18379
rect 5595 18345 5629 18379
rect 5663 18345 5697 18379
rect 5731 18345 5765 18379
rect 5799 18345 5833 18379
rect 5867 18345 5901 18379
rect 5935 18345 5969 18379
rect 6003 18345 6037 18379
rect 6071 18345 6105 18379
rect 6139 18345 6173 18379
rect 6207 18345 6241 18379
rect 6275 18345 6309 18379
rect 6343 18345 6377 18379
rect 6411 18345 6445 18379
rect 6479 18345 6513 18379
rect 6547 18345 6581 18379
rect 6615 18345 6649 18379
rect 6683 18345 6717 18379
rect 6751 18345 6785 18379
rect 6819 18345 6853 18379
rect 6887 18345 6921 18379
rect 6955 18345 6989 18379
rect 7023 18345 7057 18379
rect 7091 18345 7125 18379
rect 7159 18345 7193 18379
rect 7227 18345 7261 18379
rect 7295 18345 7329 18379
rect 7363 18345 7397 18379
rect 7431 18345 7465 18379
rect 7499 18345 7533 18379
rect 7567 18345 7601 18379
rect 7635 18345 7669 18379
rect 7703 18345 7737 18379
rect 7771 18345 7805 18379
rect 7839 18345 7873 18379
rect 7907 18345 7941 18379
rect 7975 18345 8009 18379
rect 8043 18345 8077 18379
rect 8111 18345 8145 18379
rect 8179 18345 8213 18379
rect 8247 18345 8281 18379
rect 8315 18345 8349 18379
rect 8383 18345 8417 18379
rect 8451 18345 8485 18379
rect 8519 18345 8553 18379
rect 8587 18345 8621 18379
rect 8655 18345 8689 18379
rect 8723 18345 8757 18379
rect 8791 18345 8825 18379
rect 8859 18345 8893 18379
rect 8927 18345 8961 18379
rect 8995 18345 9029 18379
rect 9063 18345 9097 18379
rect 9131 18345 9165 18379
rect 9199 18345 9233 18379
rect 9267 18345 9301 18379
rect 9335 18345 9369 18379
rect 9403 18345 9437 18379
rect 9471 18345 9505 18379
rect 9539 18345 9573 18379
rect 9607 18345 9641 18379
rect 9675 18345 9709 18379
rect 9743 18345 9777 18379
rect 9811 18345 9845 18379
rect 9879 18345 9913 18379
rect 9947 18345 9981 18379
rect 10015 18345 10049 18379
rect 10083 18345 10117 18379
rect 10151 18345 10185 18379
rect 10219 18345 10253 18379
rect 10287 18345 10321 18379
rect 10355 18345 10389 18379
rect 10423 18345 10457 18379
rect 10491 18345 10525 18379
rect 10559 18345 10593 18379
rect 10627 18345 10661 18379
rect 10695 18345 10729 18379
rect 10763 18345 10797 18379
rect 10831 18345 10865 18379
rect 10899 18345 10933 18379
rect 10967 18345 11001 18379
rect 11035 18345 11069 18379
rect 11103 18345 11137 18379
rect 11171 18345 11205 18379
rect 11239 18345 11273 18379
rect 11307 18345 11341 18379
rect 11375 18345 11409 18379
rect 11443 18345 11477 18379
rect 11511 18345 11545 18379
rect 11579 18345 11613 18379
rect 11647 18345 11681 18379
rect 11715 18345 11749 18379
rect 11783 18345 11817 18379
rect 11851 18345 11885 18379
rect 11919 18345 11953 18379
rect 11987 18345 12021 18379
rect 12055 18345 12089 18379
rect 12123 18345 12157 18379
rect 12191 18345 12225 18379
rect 12259 18345 12293 18379
rect 12327 18345 12361 18379
rect 12395 18345 12429 18379
rect 12463 18345 12497 18379
rect 12531 18345 12565 18379
rect 12599 18345 12633 18379
rect 12667 18345 12701 18379
rect 12735 18345 12769 18379
rect 12803 18345 12837 18379
rect 12871 18345 12905 18379
rect 12939 18345 12973 18379
rect 13007 18345 13041 18379
rect 13075 18345 13109 18379
rect 13143 18345 13177 18379
rect 13211 18345 13245 18379
rect 13279 18345 13313 18379
rect 13347 18345 13381 18379
rect 13415 18345 13449 18379
rect 13483 18345 13517 18379
rect 13551 18345 13585 18379
rect 13619 18345 13653 18379
rect 13687 18345 13721 18379
rect 13755 18345 13789 18379
rect 13823 18345 13857 18379
rect 13891 18345 13925 18379
rect 13959 18345 13993 18379
rect 14027 18345 14061 18379
rect 14095 18345 14129 18379
rect 14163 18345 14197 18379
rect 14231 18345 14265 18379
rect 14299 18345 14333 18379
rect 14367 18345 14401 18379
rect 14435 18345 14469 18379
rect 14503 18345 14537 18379
rect 14571 18345 14605 18379
rect 14639 18345 14673 18379
rect 14707 18345 14741 18379
rect 221 18275 255 18309
rect 290 18275 324 18309
rect 359 18275 393 18309
rect 427 18275 461 18309
rect 495 18275 529 18309
rect 563 18275 597 18309
rect 631 18275 665 18309
rect 699 18275 733 18309
rect 767 18275 801 18309
rect 835 18275 869 18309
rect 903 18275 937 18309
rect 971 18275 1005 18309
rect 1039 18275 1073 18309
rect 1107 18275 1141 18309
rect 1175 18275 1209 18309
rect 1243 18275 1277 18309
rect 1311 18275 1345 18309
rect 1379 18275 1413 18309
rect 1447 18275 1481 18309
rect 1515 18275 1549 18309
rect 1583 18275 1617 18309
rect 1651 18275 1685 18309
rect 1719 18275 1753 18309
rect 1787 18275 1821 18309
rect 1855 18275 1889 18309
rect 1923 18275 1957 18309
rect 1991 18275 2025 18309
rect 2059 18275 2093 18309
rect 2127 18275 2161 18309
rect 2195 18275 2229 18309
rect 2263 18275 2297 18309
rect 2331 18275 2365 18309
rect 2399 18275 2433 18309
rect 2467 18275 2501 18309
rect 2535 18275 2569 18309
rect 2603 18275 2637 18309
rect 2671 18275 2705 18309
rect 2739 18275 2773 18309
rect 2807 18275 2841 18309
rect 2875 18275 2909 18309
rect 2943 18275 2977 18309
rect 3011 18275 3045 18309
rect 3079 18275 3113 18309
rect 3147 18275 3181 18309
rect 3215 18275 3249 18309
rect 3283 18275 3317 18309
rect 3351 18275 3385 18309
rect 3419 18275 3453 18309
rect 3487 18275 3521 18309
rect 3555 18275 3589 18309
rect 3623 18275 3657 18309
rect 3691 18275 3725 18309
rect 3759 18275 3793 18309
rect 3827 18275 3861 18309
rect 3895 18275 3929 18309
rect 3963 18275 3997 18309
rect 4031 18275 4065 18309
rect 4099 18275 4133 18309
rect 4167 18275 4201 18309
rect 4235 18275 4269 18309
rect 4303 18275 4337 18309
rect 4371 18275 4405 18309
rect 4439 18275 4473 18309
rect 4507 18275 4541 18309
rect 4575 18275 4609 18309
rect 4643 18275 4677 18309
rect 4711 18275 4745 18309
rect 4779 18275 4813 18309
rect 4847 18275 4881 18309
rect 4915 18275 4949 18309
rect 4983 18275 5017 18309
rect 5051 18275 5085 18309
rect 5119 18275 5153 18309
rect 5187 18275 5221 18309
rect 5255 18275 5289 18309
rect 5323 18275 5357 18309
rect 5391 18275 5425 18309
rect 5459 18275 5493 18309
rect 5527 18275 5561 18309
rect 5595 18275 5629 18309
rect 5663 18275 5697 18309
rect 5731 18275 5765 18309
rect 5799 18275 5833 18309
rect 5867 18275 5901 18309
rect 5935 18275 5969 18309
rect 6003 18275 6037 18309
rect 6071 18275 6105 18309
rect 6139 18275 6173 18309
rect 6207 18275 6241 18309
rect 6275 18275 6309 18309
rect 6343 18275 6377 18309
rect 6411 18275 6445 18309
rect 6479 18275 6513 18309
rect 6547 18275 6581 18309
rect 6615 18275 6649 18309
rect 6683 18275 6717 18309
rect 6751 18275 6785 18309
rect 6819 18275 6853 18309
rect 6887 18275 6921 18309
rect 6955 18275 6989 18309
rect 7023 18275 7057 18309
rect 7091 18275 7125 18309
rect 7159 18275 7193 18309
rect 7227 18275 7261 18309
rect 7295 18275 7329 18309
rect 7363 18275 7397 18309
rect 7431 18275 7465 18309
rect 7499 18275 7533 18309
rect 7567 18275 7601 18309
rect 7635 18275 7669 18309
rect 7703 18275 7737 18309
rect 7771 18275 7805 18309
rect 7839 18275 7873 18309
rect 7907 18275 7941 18309
rect 7975 18275 8009 18309
rect 8043 18275 8077 18309
rect 8111 18275 8145 18309
rect 8179 18275 8213 18309
rect 8247 18275 8281 18309
rect 8315 18275 8349 18309
rect 8383 18275 8417 18309
rect 8451 18275 8485 18309
rect 8519 18275 8553 18309
rect 8587 18275 8621 18309
rect 8655 18275 8689 18309
rect 8723 18275 8757 18309
rect 8791 18275 8825 18309
rect 8859 18275 8893 18309
rect 8927 18275 8961 18309
rect 8995 18275 9029 18309
rect 9063 18275 9097 18309
rect 9131 18275 9165 18309
rect 9199 18275 9233 18309
rect 9267 18275 9301 18309
rect 9335 18275 9369 18309
rect 9403 18275 9437 18309
rect 9471 18275 9505 18309
rect 9539 18275 9573 18309
rect 9607 18275 9641 18309
rect 9675 18275 9709 18309
rect 9743 18275 9777 18309
rect 9811 18275 9845 18309
rect 9879 18275 9913 18309
rect 9947 18275 9981 18309
rect 10015 18275 10049 18309
rect 10083 18275 10117 18309
rect 10151 18275 10185 18309
rect 10219 18275 10253 18309
rect 10287 18275 10321 18309
rect 10355 18275 10389 18309
rect 10423 18275 10457 18309
rect 10491 18275 10525 18309
rect 10559 18275 10593 18309
rect 10627 18275 10661 18309
rect 10695 18275 10729 18309
rect 10763 18275 10797 18309
rect 10831 18275 10865 18309
rect 10899 18275 10933 18309
rect 10967 18275 11001 18309
rect 11035 18275 11069 18309
rect 11103 18275 11137 18309
rect 11171 18275 11205 18309
rect 11239 18275 11273 18309
rect 11307 18275 11341 18309
rect 11375 18275 11409 18309
rect 11443 18275 11477 18309
rect 11511 18275 11545 18309
rect 11579 18275 11613 18309
rect 11647 18275 11681 18309
rect 11715 18275 11749 18309
rect 11783 18275 11817 18309
rect 11851 18275 11885 18309
rect 11919 18275 11953 18309
rect 11987 18275 12021 18309
rect 12055 18275 12089 18309
rect 12123 18275 12157 18309
rect 12191 18275 12225 18309
rect 12259 18275 12293 18309
rect 12327 18275 12361 18309
rect 12395 18275 12429 18309
rect 12463 18275 12497 18309
rect 12531 18275 12565 18309
rect 12599 18275 12633 18309
rect 12667 18275 12701 18309
rect 12735 18275 12769 18309
rect 12803 18275 12837 18309
rect 12871 18275 12905 18309
rect 12939 18275 12973 18309
rect 13007 18275 13041 18309
rect 13075 18275 13109 18309
rect 13143 18275 13177 18309
rect 13211 18275 13245 18309
rect 13279 18275 13313 18309
rect 13347 18275 13381 18309
rect 13415 18275 13449 18309
rect 13483 18275 13517 18309
rect 13551 18275 13585 18309
rect 13619 18275 13653 18309
rect 13687 18275 13721 18309
rect 13755 18275 13789 18309
rect 13823 18275 13857 18309
rect 13891 18275 13925 18309
rect 13959 18275 13993 18309
rect 14027 18275 14061 18309
rect 14095 18275 14129 18309
rect 14163 18275 14197 18309
rect 14231 18275 14265 18309
rect 14299 18275 14333 18309
rect 14367 18275 14401 18309
rect 14435 18275 14469 18309
rect 14503 18275 14537 18309
rect 14571 18275 14605 18309
rect 14639 18275 14673 18309
rect 14707 18275 14741 18309
rect 221 18205 255 18239
rect 290 18205 324 18239
rect 359 18205 393 18239
rect 427 18205 461 18239
rect 495 18205 529 18239
rect 563 18205 597 18239
rect 631 18205 665 18239
rect 699 18205 733 18239
rect 767 18205 801 18239
rect 835 18205 869 18239
rect 903 18205 937 18239
rect 971 18205 1005 18239
rect 1039 18205 1073 18239
rect 1107 18205 1141 18239
rect 1175 18205 1209 18239
rect 1243 18205 1277 18239
rect 1311 18205 1345 18239
rect 1379 18205 1413 18239
rect 1447 18205 1481 18239
rect 1515 18205 1549 18239
rect 1583 18205 1617 18239
rect 1651 18205 1685 18239
rect 1719 18205 1753 18239
rect 1787 18205 1821 18239
rect 1855 18205 1889 18239
rect 1923 18205 1957 18239
rect 1991 18205 2025 18239
rect 2059 18205 2093 18239
rect 2127 18205 2161 18239
rect 2195 18205 2229 18239
rect 2263 18205 2297 18239
rect 2331 18205 2365 18239
rect 2399 18205 2433 18239
rect 2467 18205 2501 18239
rect 2535 18205 2569 18239
rect 2603 18205 2637 18239
rect 2671 18205 2705 18239
rect 2739 18205 2773 18239
rect 2807 18205 2841 18239
rect 2875 18205 2909 18239
rect 2943 18205 2977 18239
rect 3011 18205 3045 18239
rect 3079 18205 3113 18239
rect 3147 18205 3181 18239
rect 3215 18205 3249 18239
rect 3283 18205 3317 18239
rect 3351 18205 3385 18239
rect 3419 18205 3453 18239
rect 3487 18205 3521 18239
rect 3555 18205 3589 18239
rect 3623 18205 3657 18239
rect 3691 18205 3725 18239
rect 3759 18205 3793 18239
rect 3827 18205 3861 18239
rect 3895 18205 3929 18239
rect 3963 18205 3997 18239
rect 4031 18205 4065 18239
rect 4099 18205 4133 18239
rect 4167 18205 4201 18239
rect 4235 18205 4269 18239
rect 4303 18205 4337 18239
rect 4371 18205 4405 18239
rect 4439 18205 4473 18239
rect 4507 18205 4541 18239
rect 4575 18205 4609 18239
rect 4643 18205 4677 18239
rect 4711 18205 4745 18239
rect 4779 18205 4813 18239
rect 4847 18205 4881 18239
rect 4915 18205 4949 18239
rect 4983 18205 5017 18239
rect 5051 18205 5085 18239
rect 5119 18205 5153 18239
rect 5187 18205 5221 18239
rect 5255 18205 5289 18239
rect 5323 18205 5357 18239
rect 5391 18205 5425 18239
rect 5459 18205 5493 18239
rect 5527 18205 5561 18239
rect 5595 18205 5629 18239
rect 5663 18205 5697 18239
rect 5731 18205 5765 18239
rect 5799 18205 5833 18239
rect 5867 18205 5901 18239
rect 5935 18205 5969 18239
rect 6003 18205 6037 18239
rect 6071 18205 6105 18239
rect 6139 18205 6173 18239
rect 6207 18205 6241 18239
rect 6275 18205 6309 18239
rect 6343 18205 6377 18239
rect 6411 18205 6445 18239
rect 6479 18205 6513 18239
rect 6547 18205 6581 18239
rect 6615 18205 6649 18239
rect 6683 18205 6717 18239
rect 6751 18205 6785 18239
rect 6819 18205 6853 18239
rect 6887 18205 6921 18239
rect 6955 18205 6989 18239
rect 7023 18205 7057 18239
rect 7091 18205 7125 18239
rect 7159 18205 7193 18239
rect 7227 18205 7261 18239
rect 7295 18205 7329 18239
rect 7363 18205 7397 18239
rect 7431 18205 7465 18239
rect 7499 18205 7533 18239
rect 7567 18205 7601 18239
rect 7635 18205 7669 18239
rect 7703 18205 7737 18239
rect 7771 18205 7805 18239
rect 7839 18205 7873 18239
rect 7907 18205 7941 18239
rect 7975 18205 8009 18239
rect 8043 18205 8077 18239
rect 8111 18205 8145 18239
rect 8179 18205 8213 18239
rect 8247 18205 8281 18239
rect 8315 18205 8349 18239
rect 8383 18205 8417 18239
rect 8451 18205 8485 18239
rect 8519 18205 8553 18239
rect 8587 18205 8621 18239
rect 8655 18205 8689 18239
rect 8723 18205 8757 18239
rect 8791 18205 8825 18239
rect 8859 18205 8893 18239
rect 8927 18205 8961 18239
rect 8995 18205 9029 18239
rect 9063 18205 9097 18239
rect 9131 18205 9165 18239
rect 9199 18205 9233 18239
rect 9267 18205 9301 18239
rect 9335 18205 9369 18239
rect 9403 18205 9437 18239
rect 9471 18205 9505 18239
rect 9539 18205 9573 18239
rect 9607 18205 9641 18239
rect 9675 18205 9709 18239
rect 9743 18205 9777 18239
rect 9811 18205 9845 18239
rect 9879 18205 9913 18239
rect 9947 18205 9981 18239
rect 10015 18205 10049 18239
rect 10083 18205 10117 18239
rect 10151 18205 10185 18239
rect 10219 18205 10253 18239
rect 10287 18205 10321 18239
rect 10355 18205 10389 18239
rect 10423 18205 10457 18239
rect 10491 18205 10525 18239
rect 10559 18205 10593 18239
rect 10627 18205 10661 18239
rect 10695 18205 10729 18239
rect 10763 18205 10797 18239
rect 10831 18205 10865 18239
rect 10899 18205 10933 18239
rect 10967 18205 11001 18239
rect 11035 18205 11069 18239
rect 11103 18205 11137 18239
rect 11171 18205 11205 18239
rect 11239 18205 11273 18239
rect 11307 18205 11341 18239
rect 11375 18205 11409 18239
rect 11443 18205 11477 18239
rect 11511 18205 11545 18239
rect 11579 18205 11613 18239
rect 11647 18205 11681 18239
rect 11715 18205 11749 18239
rect 11783 18205 11817 18239
rect 11851 18205 11885 18239
rect 11919 18205 11953 18239
rect 11987 18205 12021 18239
rect 12055 18205 12089 18239
rect 12123 18205 12157 18239
rect 12191 18205 12225 18239
rect 12259 18205 12293 18239
rect 12327 18205 12361 18239
rect 12395 18205 12429 18239
rect 12463 18205 12497 18239
rect 12531 18205 12565 18239
rect 12599 18205 12633 18239
rect 12667 18205 12701 18239
rect 12735 18205 12769 18239
rect 12803 18205 12837 18239
rect 12871 18205 12905 18239
rect 12939 18205 12973 18239
rect 13007 18205 13041 18239
rect 13075 18205 13109 18239
rect 13143 18205 13177 18239
rect 13211 18205 13245 18239
rect 13279 18205 13313 18239
rect 13347 18205 13381 18239
rect 13415 18205 13449 18239
rect 13483 18205 13517 18239
rect 13551 18205 13585 18239
rect 13619 18205 13653 18239
rect 13687 18205 13721 18239
rect 13755 18205 13789 18239
rect 13823 18205 13857 18239
rect 13891 18205 13925 18239
rect 13959 18205 13993 18239
rect 14027 18205 14061 18239
rect 14095 18205 14129 18239
rect 14163 18205 14197 18239
rect 14231 18205 14265 18239
rect 14299 18205 14333 18239
rect 14367 18205 14401 18239
rect 14435 18205 14469 18239
rect 14503 18205 14537 18239
rect 14571 18205 14605 18239
rect 14639 18205 14673 18239
rect 14707 18205 14741 18239
rect 221 18135 255 18169
rect 290 18135 324 18169
rect 359 18135 393 18169
rect 427 18135 461 18169
rect 495 18135 529 18169
rect 563 18135 597 18169
rect 631 18135 665 18169
rect 699 18135 733 18169
rect 767 18135 801 18169
rect 835 18135 869 18169
rect 903 18135 937 18169
rect 971 18135 1005 18169
rect 1039 18135 1073 18169
rect 1107 18135 1141 18169
rect 1175 18135 1209 18169
rect 1243 18135 1277 18169
rect 1311 18135 1345 18169
rect 1379 18135 1413 18169
rect 1447 18135 1481 18169
rect 1515 18135 1549 18169
rect 1583 18135 1617 18169
rect 1651 18135 1685 18169
rect 1719 18135 1753 18169
rect 1787 18135 1821 18169
rect 1855 18135 1889 18169
rect 1923 18135 1957 18169
rect 1991 18135 2025 18169
rect 2059 18135 2093 18169
rect 2127 18135 2161 18169
rect 2195 18135 2229 18169
rect 2263 18135 2297 18169
rect 2331 18135 2365 18169
rect 2399 18135 2433 18169
rect 2467 18135 2501 18169
rect 2535 18135 2569 18169
rect 2603 18135 2637 18169
rect 2671 18135 2705 18169
rect 2739 18135 2773 18169
rect 2807 18135 2841 18169
rect 2875 18135 2909 18169
rect 2943 18135 2977 18169
rect 3011 18135 3045 18169
rect 3079 18135 3113 18169
rect 3147 18135 3181 18169
rect 3215 18135 3249 18169
rect 3283 18135 3317 18169
rect 3351 18135 3385 18169
rect 3419 18135 3453 18169
rect 3487 18135 3521 18169
rect 3555 18135 3589 18169
rect 3623 18135 3657 18169
rect 3691 18135 3725 18169
rect 3759 18135 3793 18169
rect 3827 18135 3861 18169
rect 3895 18135 3929 18169
rect 3963 18135 3997 18169
rect 4031 18135 4065 18169
rect 4099 18135 4133 18169
rect 4167 18135 4201 18169
rect 4235 18135 4269 18169
rect 4303 18135 4337 18169
rect 4371 18135 4405 18169
rect 4439 18135 4473 18169
rect 4507 18135 4541 18169
rect 4575 18135 4609 18169
rect 4643 18135 4677 18169
rect 4711 18135 4745 18169
rect 4779 18135 4813 18169
rect 4847 18135 4881 18169
rect 4915 18135 4949 18169
rect 4983 18135 5017 18169
rect 5051 18135 5085 18169
rect 5119 18135 5153 18169
rect 5187 18135 5221 18169
rect 5255 18135 5289 18169
rect 5323 18135 5357 18169
rect 5391 18135 5425 18169
rect 5459 18135 5493 18169
rect 5527 18135 5561 18169
rect 5595 18135 5629 18169
rect 5663 18135 5697 18169
rect 5731 18135 5765 18169
rect 5799 18135 5833 18169
rect 5867 18135 5901 18169
rect 5935 18135 5969 18169
rect 6003 18135 6037 18169
rect 6071 18135 6105 18169
rect 6139 18135 6173 18169
rect 6207 18135 6241 18169
rect 6275 18135 6309 18169
rect 6343 18135 6377 18169
rect 6411 18135 6445 18169
rect 6479 18135 6513 18169
rect 6547 18135 6581 18169
rect 6615 18135 6649 18169
rect 6683 18135 6717 18169
rect 6751 18135 6785 18169
rect 6819 18135 6853 18169
rect 6887 18135 6921 18169
rect 6955 18135 6989 18169
rect 7023 18135 7057 18169
rect 7091 18135 7125 18169
rect 7159 18135 7193 18169
rect 7227 18135 7261 18169
rect 7295 18135 7329 18169
rect 7363 18135 7397 18169
rect 7431 18135 7465 18169
rect 7499 18135 7533 18169
rect 7567 18135 7601 18169
rect 7635 18135 7669 18169
rect 7703 18135 7737 18169
rect 7771 18135 7805 18169
rect 7839 18135 7873 18169
rect 7907 18135 7941 18169
rect 7975 18135 8009 18169
rect 8043 18135 8077 18169
rect 8111 18135 8145 18169
rect 8179 18135 8213 18169
rect 8247 18135 8281 18169
rect 8315 18135 8349 18169
rect 8383 18135 8417 18169
rect 8451 18135 8485 18169
rect 8519 18135 8553 18169
rect 8587 18135 8621 18169
rect 8655 18135 8689 18169
rect 8723 18135 8757 18169
rect 8791 18135 8825 18169
rect 8859 18135 8893 18169
rect 8927 18135 8961 18169
rect 8995 18135 9029 18169
rect 9063 18135 9097 18169
rect 9131 18135 9165 18169
rect 9199 18135 9233 18169
rect 9267 18135 9301 18169
rect 9335 18135 9369 18169
rect 9403 18135 9437 18169
rect 9471 18135 9505 18169
rect 9539 18135 9573 18169
rect 9607 18135 9641 18169
rect 9675 18135 9709 18169
rect 9743 18135 9777 18169
rect 9811 18135 9845 18169
rect 9879 18135 9913 18169
rect 9947 18135 9981 18169
rect 10015 18135 10049 18169
rect 10083 18135 10117 18169
rect 10151 18135 10185 18169
rect 10219 18135 10253 18169
rect 10287 18135 10321 18169
rect 10355 18135 10389 18169
rect 10423 18135 10457 18169
rect 10491 18135 10525 18169
rect 10559 18135 10593 18169
rect 10627 18135 10661 18169
rect 10695 18135 10729 18169
rect 10763 18135 10797 18169
rect 10831 18135 10865 18169
rect 10899 18135 10933 18169
rect 10967 18135 11001 18169
rect 11035 18135 11069 18169
rect 11103 18135 11137 18169
rect 11171 18135 11205 18169
rect 11239 18135 11273 18169
rect 11307 18135 11341 18169
rect 11375 18135 11409 18169
rect 11443 18135 11477 18169
rect 11511 18135 11545 18169
rect 11579 18135 11613 18169
rect 11647 18135 11681 18169
rect 11715 18135 11749 18169
rect 11783 18135 11817 18169
rect 11851 18135 11885 18169
rect 11919 18135 11953 18169
rect 11987 18135 12021 18169
rect 12055 18135 12089 18169
rect 12123 18135 12157 18169
rect 12191 18135 12225 18169
rect 12259 18135 12293 18169
rect 12327 18135 12361 18169
rect 12395 18135 12429 18169
rect 12463 18135 12497 18169
rect 12531 18135 12565 18169
rect 12599 18135 12633 18169
rect 12667 18135 12701 18169
rect 12735 18135 12769 18169
rect 12803 18135 12837 18169
rect 12871 18135 12905 18169
rect 12939 18135 12973 18169
rect 13007 18135 13041 18169
rect 13075 18135 13109 18169
rect 13143 18135 13177 18169
rect 13211 18135 13245 18169
rect 13279 18135 13313 18169
rect 13347 18135 13381 18169
rect 13415 18135 13449 18169
rect 13483 18135 13517 18169
rect 13551 18135 13585 18169
rect 13619 18135 13653 18169
rect 13687 18135 13721 18169
rect 13755 18135 13789 18169
rect 13823 18135 13857 18169
rect 13891 18135 13925 18169
rect 13959 18135 13993 18169
rect 14027 18135 14061 18169
rect 14095 18135 14129 18169
rect 14163 18135 14197 18169
rect 14231 18135 14265 18169
rect 14299 18135 14333 18169
rect 14367 18135 14401 18169
rect 14435 18135 14469 18169
rect 14503 18135 14537 18169
rect 14571 18135 14605 18169
rect 14639 18135 14673 18169
rect 14707 18135 14741 18169
rect 221 18065 255 18099
rect 290 18065 324 18099
rect 359 18065 393 18099
rect 427 18065 461 18099
rect 495 18065 529 18099
rect 563 18065 597 18099
rect 631 18065 665 18099
rect 699 18065 733 18099
rect 767 18065 801 18099
rect 835 18065 869 18099
rect 903 18065 937 18099
rect 971 18065 1005 18099
rect 1039 18065 1073 18099
rect 1107 18065 1141 18099
rect 1175 18065 1209 18099
rect 1243 18065 1277 18099
rect 1311 18065 1345 18099
rect 1379 18065 1413 18099
rect 1447 18065 1481 18099
rect 1515 18065 1549 18099
rect 1583 18065 1617 18099
rect 1651 18065 1685 18099
rect 1719 18065 1753 18099
rect 1787 18065 1821 18099
rect 1855 18065 1889 18099
rect 1923 18065 1957 18099
rect 1991 18065 2025 18099
rect 2059 18065 2093 18099
rect 2127 18065 2161 18099
rect 2195 18065 2229 18099
rect 2263 18065 2297 18099
rect 2331 18065 2365 18099
rect 2399 18065 2433 18099
rect 2467 18065 2501 18099
rect 2535 18065 2569 18099
rect 2603 18065 2637 18099
rect 2671 18065 2705 18099
rect 2739 18065 2773 18099
rect 2807 18065 2841 18099
rect 2875 18065 2909 18099
rect 2943 18065 2977 18099
rect 3011 18065 3045 18099
rect 3079 18065 3113 18099
rect 3147 18065 3181 18099
rect 3215 18065 3249 18099
rect 3283 18065 3317 18099
rect 3351 18065 3385 18099
rect 3419 18065 3453 18099
rect 3487 18065 3521 18099
rect 3555 18065 3589 18099
rect 3623 18065 3657 18099
rect 3691 18065 3725 18099
rect 3759 18065 3793 18099
rect 3827 18065 3861 18099
rect 3895 18065 3929 18099
rect 3963 18065 3997 18099
rect 4031 18065 4065 18099
rect 4099 18065 4133 18099
rect 4167 18065 4201 18099
rect 4235 18065 4269 18099
rect 4303 18065 4337 18099
rect 4371 18065 4405 18099
rect 4439 18065 4473 18099
rect 4507 18065 4541 18099
rect 4575 18065 4609 18099
rect 4643 18065 4677 18099
rect 4711 18065 4745 18099
rect 4779 18065 4813 18099
rect 4847 18065 4881 18099
rect 4915 18065 4949 18099
rect 4983 18065 5017 18099
rect 5051 18065 5085 18099
rect 5119 18065 5153 18099
rect 5187 18065 5221 18099
rect 5255 18065 5289 18099
rect 5323 18065 5357 18099
rect 5391 18065 5425 18099
rect 5459 18065 5493 18099
rect 5527 18065 5561 18099
rect 5595 18065 5629 18099
rect 5663 18065 5697 18099
rect 5731 18065 5765 18099
rect 5799 18065 5833 18099
rect 5867 18065 5901 18099
rect 5935 18065 5969 18099
rect 6003 18065 6037 18099
rect 6071 18065 6105 18099
rect 6139 18065 6173 18099
rect 6207 18065 6241 18099
rect 6275 18065 6309 18099
rect 6343 18065 6377 18099
rect 6411 18065 6445 18099
rect 6479 18065 6513 18099
rect 6547 18065 6581 18099
rect 6615 18065 6649 18099
rect 6683 18065 6717 18099
rect 6751 18065 6785 18099
rect 6819 18065 6853 18099
rect 6887 18065 6921 18099
rect 6955 18065 6989 18099
rect 7023 18065 7057 18099
rect 7091 18065 7125 18099
rect 7159 18065 7193 18099
rect 7227 18065 7261 18099
rect 7295 18065 7329 18099
rect 7363 18065 7397 18099
rect 7431 18065 7465 18099
rect 7499 18065 7533 18099
rect 7567 18065 7601 18099
rect 7635 18065 7669 18099
rect 7703 18065 7737 18099
rect 7771 18065 7805 18099
rect 7839 18065 7873 18099
rect 7907 18065 7941 18099
rect 7975 18065 8009 18099
rect 8043 18065 8077 18099
rect 8111 18065 8145 18099
rect 8179 18065 8213 18099
rect 8247 18065 8281 18099
rect 8315 18065 8349 18099
rect 8383 18065 8417 18099
rect 8451 18065 8485 18099
rect 8519 18065 8553 18099
rect 8587 18065 8621 18099
rect 8655 18065 8689 18099
rect 8723 18065 8757 18099
rect 8791 18065 8825 18099
rect 8859 18065 8893 18099
rect 8927 18065 8961 18099
rect 8995 18065 9029 18099
rect 9063 18065 9097 18099
rect 9131 18065 9165 18099
rect 9199 18065 9233 18099
rect 9267 18065 9301 18099
rect 9335 18065 9369 18099
rect 9403 18065 9437 18099
rect 9471 18065 9505 18099
rect 9539 18065 9573 18099
rect 9607 18065 9641 18099
rect 9675 18065 9709 18099
rect 9743 18065 9777 18099
rect 9811 18065 9845 18099
rect 9879 18065 9913 18099
rect 9947 18065 9981 18099
rect 10015 18065 10049 18099
rect 10083 18065 10117 18099
rect 10151 18065 10185 18099
rect 10219 18065 10253 18099
rect 10287 18065 10321 18099
rect 10355 18065 10389 18099
rect 10423 18065 10457 18099
rect 10491 18065 10525 18099
rect 10559 18065 10593 18099
rect 10627 18065 10661 18099
rect 10695 18065 10729 18099
rect 10763 18065 10797 18099
rect 10831 18065 10865 18099
rect 10899 18065 10933 18099
rect 10967 18065 11001 18099
rect 11035 18065 11069 18099
rect 11103 18065 11137 18099
rect 11171 18065 11205 18099
rect 11239 18065 11273 18099
rect 11307 18065 11341 18099
rect 11375 18065 11409 18099
rect 11443 18065 11477 18099
rect 11511 18065 11545 18099
rect 11579 18065 11613 18099
rect 11647 18065 11681 18099
rect 11715 18065 11749 18099
rect 11783 18065 11817 18099
rect 11851 18065 11885 18099
rect 11919 18065 11953 18099
rect 11987 18065 12021 18099
rect 12055 18065 12089 18099
rect 12123 18065 12157 18099
rect 12191 18065 12225 18099
rect 12259 18065 12293 18099
rect 12327 18065 12361 18099
rect 12395 18065 12429 18099
rect 12463 18065 12497 18099
rect 12531 18065 12565 18099
rect 12599 18065 12633 18099
rect 12667 18065 12701 18099
rect 12735 18065 12769 18099
rect 12803 18065 12837 18099
rect 12871 18065 12905 18099
rect 12939 18065 12973 18099
rect 13007 18065 13041 18099
rect 13075 18065 13109 18099
rect 13143 18065 13177 18099
rect 13211 18065 13245 18099
rect 13279 18065 13313 18099
rect 13347 18065 13381 18099
rect 13415 18065 13449 18099
rect 13483 18065 13517 18099
rect 13551 18065 13585 18099
rect 13619 18065 13653 18099
rect 13687 18065 13721 18099
rect 13755 18065 13789 18099
rect 13823 18065 13857 18099
rect 13891 18065 13925 18099
rect 13959 18065 13993 18099
rect 14027 18065 14061 18099
rect 14095 18065 14129 18099
rect 14163 18065 14197 18099
rect 14231 18065 14265 18099
rect 14299 18065 14333 18099
rect 14367 18065 14401 18099
rect 14435 18065 14469 18099
rect 14503 18065 14537 18099
rect 14571 18065 14605 18099
rect 14639 18065 14673 18099
rect 14707 18065 14741 18099
rect 221 17995 255 18029
rect 290 17995 324 18029
rect 359 17995 393 18029
rect 427 17995 461 18029
rect 495 17995 529 18029
rect 563 17995 597 18029
rect 631 17995 665 18029
rect 699 17995 733 18029
rect 767 17995 801 18029
rect 835 17995 869 18029
rect 903 17995 937 18029
rect 971 17995 1005 18029
rect 1039 17995 1073 18029
rect 1107 17995 1141 18029
rect 1175 17995 1209 18029
rect 1243 17995 1277 18029
rect 1311 17995 1345 18029
rect 1379 17995 1413 18029
rect 1447 17995 1481 18029
rect 1515 17995 1549 18029
rect 1583 17995 1617 18029
rect 1651 17995 1685 18029
rect 1719 17995 1753 18029
rect 1787 17995 1821 18029
rect 1855 17995 1889 18029
rect 1923 17995 1957 18029
rect 1991 17995 2025 18029
rect 2059 17995 2093 18029
rect 2127 17995 2161 18029
rect 2195 17995 2229 18029
rect 2263 17995 2297 18029
rect 2331 17995 2365 18029
rect 2399 17995 2433 18029
rect 2467 17995 2501 18029
rect 2535 17995 2569 18029
rect 2603 17995 2637 18029
rect 2671 17995 2705 18029
rect 2739 17995 2773 18029
rect 2807 17995 2841 18029
rect 2875 17995 2909 18029
rect 2943 17995 2977 18029
rect 3011 17995 3045 18029
rect 3079 17995 3113 18029
rect 3147 17995 3181 18029
rect 3215 17995 3249 18029
rect 3283 17995 3317 18029
rect 3351 17995 3385 18029
rect 3419 17995 3453 18029
rect 3487 17995 3521 18029
rect 3555 17995 3589 18029
rect 3623 17995 3657 18029
rect 3691 17995 3725 18029
rect 3759 17995 3793 18029
rect 3827 17995 3861 18029
rect 3895 17995 3929 18029
rect 3963 17995 3997 18029
rect 4031 17995 4065 18029
rect 4099 17995 4133 18029
rect 4167 17995 4201 18029
rect 4235 17995 4269 18029
rect 4303 17995 4337 18029
rect 4371 17995 4405 18029
rect 4439 17995 4473 18029
rect 4507 17995 4541 18029
rect 4575 17995 4609 18029
rect 4643 17995 4677 18029
rect 4711 17995 4745 18029
rect 4779 17995 4813 18029
rect 4847 17995 4881 18029
rect 4915 17995 4949 18029
rect 4983 17995 5017 18029
rect 5051 17995 5085 18029
rect 5119 17995 5153 18029
rect 5187 17995 5221 18029
rect 5255 17995 5289 18029
rect 5323 17995 5357 18029
rect 5391 17995 5425 18029
rect 5459 17995 5493 18029
rect 5527 17995 5561 18029
rect 5595 17995 5629 18029
rect 5663 17995 5697 18029
rect 5731 17995 5765 18029
rect 5799 17995 5833 18029
rect 5867 17995 5901 18029
rect 5935 17995 5969 18029
rect 6003 17995 6037 18029
rect 6071 17995 6105 18029
rect 6139 17995 6173 18029
rect 6207 17995 6241 18029
rect 6275 17995 6309 18029
rect 6343 17995 6377 18029
rect 6411 17995 6445 18029
rect 6479 17995 6513 18029
rect 6547 17995 6581 18029
rect 6615 17995 6649 18029
rect 6683 17995 6717 18029
rect 6751 17995 6785 18029
rect 6819 17995 6853 18029
rect 6887 17995 6921 18029
rect 6955 17995 6989 18029
rect 7023 17995 7057 18029
rect 7091 17995 7125 18029
rect 7159 17995 7193 18029
rect 7227 17995 7261 18029
rect 7295 17995 7329 18029
rect 7363 17995 7397 18029
rect 7431 17995 7465 18029
rect 7499 17995 7533 18029
rect 7567 17995 7601 18029
rect 7635 17995 7669 18029
rect 7703 17995 7737 18029
rect 7771 17995 7805 18029
rect 7839 17995 7873 18029
rect 7907 17995 7941 18029
rect 7975 17995 8009 18029
rect 8043 17995 8077 18029
rect 8111 17995 8145 18029
rect 8179 17995 8213 18029
rect 8247 17995 8281 18029
rect 8315 17995 8349 18029
rect 8383 17995 8417 18029
rect 8451 17995 8485 18029
rect 8519 17995 8553 18029
rect 8587 17995 8621 18029
rect 8655 17995 8689 18029
rect 8723 17995 8757 18029
rect 8791 17995 8825 18029
rect 8859 17995 8893 18029
rect 8927 17995 8961 18029
rect 8995 17995 9029 18029
rect 9063 17995 9097 18029
rect 9131 17995 9165 18029
rect 9199 17995 9233 18029
rect 9267 17995 9301 18029
rect 9335 17995 9369 18029
rect 9403 17995 9437 18029
rect 9471 17995 9505 18029
rect 9539 17995 9573 18029
rect 9607 17995 9641 18029
rect 9675 17995 9709 18029
rect 9743 17995 9777 18029
rect 9811 17995 9845 18029
rect 9879 17995 9913 18029
rect 9947 17995 9981 18029
rect 10015 17995 10049 18029
rect 10083 17995 10117 18029
rect 10151 17995 10185 18029
rect 10219 17995 10253 18029
rect 10287 17995 10321 18029
rect 10355 17995 10389 18029
rect 10423 17995 10457 18029
rect 10491 17995 10525 18029
rect 10559 17995 10593 18029
rect 10627 17995 10661 18029
rect 10695 17995 10729 18029
rect 10763 17995 10797 18029
rect 10831 17995 10865 18029
rect 10899 17995 10933 18029
rect 10967 17995 11001 18029
rect 11035 17995 11069 18029
rect 11103 17995 11137 18029
rect 11171 17995 11205 18029
rect 11239 17995 11273 18029
rect 11307 17995 11341 18029
rect 11375 17995 11409 18029
rect 11443 17995 11477 18029
rect 11511 17995 11545 18029
rect 11579 17995 11613 18029
rect 11647 17995 11681 18029
rect 11715 17995 11749 18029
rect 11783 17995 11817 18029
rect 11851 17995 11885 18029
rect 11919 17995 11953 18029
rect 11987 17995 12021 18029
rect 12055 17995 12089 18029
rect 12123 17995 12157 18029
rect 12191 17995 12225 18029
rect 12259 17995 12293 18029
rect 12327 17995 12361 18029
rect 12395 17995 12429 18029
rect 12463 17995 12497 18029
rect 12531 17995 12565 18029
rect 12599 17995 12633 18029
rect 12667 17995 12701 18029
rect 12735 17995 12769 18029
rect 12803 17995 12837 18029
rect 12871 17995 12905 18029
rect 12939 17995 12973 18029
rect 13007 17995 13041 18029
rect 13075 17995 13109 18029
rect 13143 17995 13177 18029
rect 13211 17995 13245 18029
rect 13279 17995 13313 18029
rect 13347 17995 13381 18029
rect 13415 17995 13449 18029
rect 13483 17995 13517 18029
rect 13551 17995 13585 18029
rect 13619 17995 13653 18029
rect 13687 17995 13721 18029
rect 13755 17995 13789 18029
rect 13823 17995 13857 18029
rect 13891 17995 13925 18029
rect 13959 17995 13993 18029
rect 14027 17995 14061 18029
rect 14095 17995 14129 18029
rect 14163 17995 14197 18029
rect 14231 17995 14265 18029
rect 14299 17995 14333 18029
rect 14367 17995 14401 18029
rect 14435 17995 14469 18029
rect 14503 17995 14537 18029
rect 14571 17995 14605 18029
rect 14639 17995 14673 18029
rect 14707 17995 14741 18029
rect 221 17925 255 17959
rect 290 17925 324 17959
rect 359 17925 393 17959
rect 427 17925 461 17959
rect 495 17925 529 17959
rect 563 17925 597 17959
rect 631 17925 665 17959
rect 699 17925 733 17959
rect 767 17925 801 17959
rect 835 17925 869 17959
rect 903 17925 937 17959
rect 971 17925 1005 17959
rect 1039 17925 1073 17959
rect 1107 17925 1141 17959
rect 1175 17925 1209 17959
rect 1243 17925 1277 17959
rect 1311 17925 1345 17959
rect 1379 17925 1413 17959
rect 1447 17925 1481 17959
rect 1515 17925 1549 17959
rect 1583 17925 1617 17959
rect 1651 17925 1685 17959
rect 1719 17925 1753 17959
rect 1787 17925 1821 17959
rect 1855 17925 1889 17959
rect 1923 17925 1957 17959
rect 1991 17925 2025 17959
rect 2059 17925 2093 17959
rect 2127 17925 2161 17959
rect 2195 17925 2229 17959
rect 2263 17925 2297 17959
rect 2331 17925 2365 17959
rect 2399 17925 2433 17959
rect 2467 17925 2501 17959
rect 2535 17925 2569 17959
rect 2603 17925 2637 17959
rect 2671 17925 2705 17959
rect 2739 17925 2773 17959
rect 2807 17925 2841 17959
rect 2875 17925 2909 17959
rect 2943 17925 2977 17959
rect 3011 17925 3045 17959
rect 3079 17925 3113 17959
rect 3147 17925 3181 17959
rect 3215 17925 3249 17959
rect 3283 17925 3317 17959
rect 3351 17925 3385 17959
rect 3419 17925 3453 17959
rect 3487 17925 3521 17959
rect 3555 17925 3589 17959
rect 3623 17925 3657 17959
rect 3691 17925 3725 17959
rect 3759 17925 3793 17959
rect 3827 17925 3861 17959
rect 3895 17925 3929 17959
rect 3963 17925 3997 17959
rect 4031 17925 4065 17959
rect 4099 17925 4133 17959
rect 4167 17925 4201 17959
rect 4235 17925 4269 17959
rect 4303 17925 4337 17959
rect 4371 17925 4405 17959
rect 4439 17925 4473 17959
rect 4507 17925 4541 17959
rect 4575 17925 4609 17959
rect 4643 17925 4677 17959
rect 4711 17925 4745 17959
rect 4779 17925 4813 17959
rect 4847 17925 4881 17959
rect 4915 17925 4949 17959
rect 4983 17925 5017 17959
rect 5051 17925 5085 17959
rect 5119 17925 5153 17959
rect 5187 17925 5221 17959
rect 5255 17925 5289 17959
rect 5323 17925 5357 17959
rect 5391 17925 5425 17959
rect 5459 17925 5493 17959
rect 5527 17925 5561 17959
rect 5595 17925 5629 17959
rect 5663 17925 5697 17959
rect 5731 17925 5765 17959
rect 5799 17925 5833 17959
rect 5867 17925 5901 17959
rect 5935 17925 5969 17959
rect 6003 17925 6037 17959
rect 6071 17925 6105 17959
rect 6139 17925 6173 17959
rect 6207 17925 6241 17959
rect 6275 17925 6309 17959
rect 6343 17925 6377 17959
rect 6411 17925 6445 17959
rect 6479 17925 6513 17959
rect 6547 17925 6581 17959
rect 6615 17925 6649 17959
rect 6683 17925 6717 17959
rect 6751 17925 6785 17959
rect 6819 17925 6853 17959
rect 6887 17925 6921 17959
rect 6955 17925 6989 17959
rect 7023 17925 7057 17959
rect 7091 17925 7125 17959
rect 7159 17925 7193 17959
rect 7227 17925 7261 17959
rect 7295 17925 7329 17959
rect 7363 17925 7397 17959
rect 7431 17925 7465 17959
rect 7499 17925 7533 17959
rect 7567 17925 7601 17959
rect 7635 17925 7669 17959
rect 7703 17925 7737 17959
rect 7771 17925 7805 17959
rect 7839 17925 7873 17959
rect 7907 17925 7941 17959
rect 7975 17925 8009 17959
rect 8043 17925 8077 17959
rect 8111 17925 8145 17959
rect 8179 17925 8213 17959
rect 8247 17925 8281 17959
rect 8315 17925 8349 17959
rect 8383 17925 8417 17959
rect 8451 17925 8485 17959
rect 8519 17925 8553 17959
rect 8587 17925 8621 17959
rect 8655 17925 8689 17959
rect 8723 17925 8757 17959
rect 8791 17925 8825 17959
rect 8859 17925 8893 17959
rect 8927 17925 8961 17959
rect 8995 17925 9029 17959
rect 9063 17925 9097 17959
rect 9131 17925 9165 17959
rect 9199 17925 9233 17959
rect 9267 17925 9301 17959
rect 9335 17925 9369 17959
rect 9403 17925 9437 17959
rect 9471 17925 9505 17959
rect 9539 17925 9573 17959
rect 9607 17925 9641 17959
rect 9675 17925 9709 17959
rect 9743 17925 9777 17959
rect 9811 17925 9845 17959
rect 9879 17925 9913 17959
rect 9947 17925 9981 17959
rect 10015 17925 10049 17959
rect 10083 17925 10117 17959
rect 10151 17925 10185 17959
rect 10219 17925 10253 17959
rect 10287 17925 10321 17959
rect 10355 17925 10389 17959
rect 10423 17925 10457 17959
rect 10491 17925 10525 17959
rect 10559 17925 10593 17959
rect 10627 17925 10661 17959
rect 10695 17925 10729 17959
rect 10763 17925 10797 17959
rect 10831 17925 10865 17959
rect 10899 17925 10933 17959
rect 10967 17925 11001 17959
rect 11035 17925 11069 17959
rect 11103 17925 11137 17959
rect 11171 17925 11205 17959
rect 11239 17925 11273 17959
rect 11307 17925 11341 17959
rect 11375 17925 11409 17959
rect 11443 17925 11477 17959
rect 11511 17925 11545 17959
rect 11579 17925 11613 17959
rect 11647 17925 11681 17959
rect 11715 17925 11749 17959
rect 11783 17925 11817 17959
rect 11851 17925 11885 17959
rect 11919 17925 11953 17959
rect 11987 17925 12021 17959
rect 12055 17925 12089 17959
rect 12123 17925 12157 17959
rect 12191 17925 12225 17959
rect 12259 17925 12293 17959
rect 12327 17925 12361 17959
rect 12395 17925 12429 17959
rect 12463 17925 12497 17959
rect 12531 17925 12565 17959
rect 12599 17925 12633 17959
rect 12667 17925 12701 17959
rect 12735 17925 12769 17959
rect 12803 17925 12837 17959
rect 12871 17925 12905 17959
rect 12939 17925 12973 17959
rect 13007 17925 13041 17959
rect 13075 17925 13109 17959
rect 13143 17925 13177 17959
rect 13211 17925 13245 17959
rect 13279 17925 13313 17959
rect 13347 17925 13381 17959
rect 13415 17925 13449 17959
rect 13483 17925 13517 17959
rect 13551 17925 13585 17959
rect 13619 17925 13653 17959
rect 13687 17925 13721 17959
rect 13755 17925 13789 17959
rect 13823 17925 13857 17959
rect 13891 17925 13925 17959
rect 13959 17925 13993 17959
rect 14027 17925 14061 17959
rect 14095 17925 14129 17959
rect 14163 17925 14197 17959
rect 14231 17925 14265 17959
rect 14299 17925 14333 17959
rect 14367 17925 14401 17959
rect 14435 17925 14469 17959
rect 14503 17925 14537 17959
rect 14571 17925 14605 17959
rect 14639 17925 14673 17959
rect 14707 17925 14741 17959
rect 221 17855 255 17889
rect 290 17855 324 17889
rect 359 17855 393 17889
rect 427 17855 461 17889
rect 495 17855 529 17889
rect 563 17855 597 17889
rect 631 17855 665 17889
rect 699 17855 733 17889
rect 767 17855 801 17889
rect 835 17855 869 17889
rect 903 17855 937 17889
rect 971 17855 1005 17889
rect 1039 17855 1073 17889
rect 1107 17855 1141 17889
rect 1175 17855 1209 17889
rect 1243 17855 1277 17889
rect 1311 17855 1345 17889
rect 1379 17855 1413 17889
rect 1447 17855 1481 17889
rect 1515 17855 1549 17889
rect 1583 17855 1617 17889
rect 1651 17855 1685 17889
rect 1719 17855 1753 17889
rect 1787 17855 1821 17889
rect 1855 17855 1889 17889
rect 1923 17855 1957 17889
rect 1991 17855 2025 17889
rect 2059 17855 2093 17889
rect 2127 17855 2161 17889
rect 2195 17855 2229 17889
rect 2263 17855 2297 17889
rect 2331 17855 2365 17889
rect 2399 17855 2433 17889
rect 2467 17855 2501 17889
rect 2535 17855 2569 17889
rect 2603 17855 2637 17889
rect 2671 17855 2705 17889
rect 2739 17855 2773 17889
rect 2807 17855 2841 17889
rect 2875 17855 2909 17889
rect 2943 17855 2977 17889
rect 3011 17855 3045 17889
rect 3079 17855 3113 17889
rect 3147 17855 3181 17889
rect 3215 17855 3249 17889
rect 3283 17855 3317 17889
rect 3351 17855 3385 17889
rect 3419 17855 3453 17889
rect 3487 17855 3521 17889
rect 3555 17855 3589 17889
rect 3623 17855 3657 17889
rect 3691 17855 3725 17889
rect 3759 17855 3793 17889
rect 3827 17855 3861 17889
rect 3895 17855 3929 17889
rect 3963 17855 3997 17889
rect 4031 17855 4065 17889
rect 4099 17855 4133 17889
rect 4167 17855 4201 17889
rect 4235 17855 4269 17889
rect 4303 17855 4337 17889
rect 4371 17855 4405 17889
rect 4439 17855 4473 17889
rect 4507 17855 4541 17889
rect 4575 17855 4609 17889
rect 4643 17855 4677 17889
rect 4711 17855 4745 17889
rect 4779 17855 4813 17889
rect 4847 17855 4881 17889
rect 4915 17855 4949 17889
rect 4983 17855 5017 17889
rect 5051 17855 5085 17889
rect 5119 17855 5153 17889
rect 5187 17855 5221 17889
rect 5255 17855 5289 17889
rect 5323 17855 5357 17889
rect 5391 17855 5425 17889
rect 5459 17855 5493 17889
rect 5527 17855 5561 17889
rect 5595 17855 5629 17889
rect 5663 17855 5697 17889
rect 5731 17855 5765 17889
rect 5799 17855 5833 17889
rect 5867 17855 5901 17889
rect 5935 17855 5969 17889
rect 6003 17855 6037 17889
rect 6071 17855 6105 17889
rect 6139 17855 6173 17889
rect 6207 17855 6241 17889
rect 6275 17855 6309 17889
rect 6343 17855 6377 17889
rect 6411 17855 6445 17889
rect 6479 17855 6513 17889
rect 6547 17855 6581 17889
rect 6615 17855 6649 17889
rect 6683 17855 6717 17889
rect 6751 17855 6785 17889
rect 6819 17855 6853 17889
rect 6887 17855 6921 17889
rect 6955 17855 6989 17889
rect 7023 17855 7057 17889
rect 7091 17855 7125 17889
rect 7159 17855 7193 17889
rect 7227 17855 7261 17889
rect 7295 17855 7329 17889
rect 7363 17855 7397 17889
rect 7431 17855 7465 17889
rect 7499 17855 7533 17889
rect 7567 17855 7601 17889
rect 7635 17855 7669 17889
rect 7703 17855 7737 17889
rect 7771 17855 7805 17889
rect 7839 17855 7873 17889
rect 7907 17855 7941 17889
rect 7975 17855 8009 17889
rect 8043 17855 8077 17889
rect 8111 17855 8145 17889
rect 8179 17855 8213 17889
rect 8247 17855 8281 17889
rect 8315 17855 8349 17889
rect 8383 17855 8417 17889
rect 8451 17855 8485 17889
rect 8519 17855 8553 17889
rect 8587 17855 8621 17889
rect 8655 17855 8689 17889
rect 8723 17855 8757 17889
rect 8791 17855 8825 17889
rect 8859 17855 8893 17889
rect 8927 17855 8961 17889
rect 8995 17855 9029 17889
rect 9063 17855 9097 17889
rect 9131 17855 9165 17889
rect 9199 17855 9233 17889
rect 9267 17855 9301 17889
rect 9335 17855 9369 17889
rect 9403 17855 9437 17889
rect 9471 17855 9505 17889
rect 9539 17855 9573 17889
rect 9607 17855 9641 17889
rect 9675 17855 9709 17889
rect 9743 17855 9777 17889
rect 9811 17855 9845 17889
rect 9879 17855 9913 17889
rect 9947 17855 9981 17889
rect 10015 17855 10049 17889
rect 10083 17855 10117 17889
rect 10151 17855 10185 17889
rect 10219 17855 10253 17889
rect 10287 17855 10321 17889
rect 10355 17855 10389 17889
rect 10423 17855 10457 17889
rect 10491 17855 10525 17889
rect 10559 17855 10593 17889
rect 10627 17855 10661 17889
rect 10695 17855 10729 17889
rect 10763 17855 10797 17889
rect 10831 17855 10865 17889
rect 10899 17855 10933 17889
rect 10967 17855 11001 17889
rect 11035 17855 11069 17889
rect 11103 17855 11137 17889
rect 11171 17855 11205 17889
rect 11239 17855 11273 17889
rect 11307 17855 11341 17889
rect 11375 17855 11409 17889
rect 11443 17855 11477 17889
rect 11511 17855 11545 17889
rect 11579 17855 11613 17889
rect 11647 17855 11681 17889
rect 11715 17855 11749 17889
rect 11783 17855 11817 17889
rect 11851 17855 11885 17889
rect 11919 17855 11953 17889
rect 11987 17855 12021 17889
rect 12055 17855 12089 17889
rect 12123 17855 12157 17889
rect 12191 17855 12225 17889
rect 12259 17855 12293 17889
rect 12327 17855 12361 17889
rect 12395 17855 12429 17889
rect 12463 17855 12497 17889
rect 12531 17855 12565 17889
rect 12599 17855 12633 17889
rect 12667 17855 12701 17889
rect 12735 17855 12769 17889
rect 12803 17855 12837 17889
rect 12871 17855 12905 17889
rect 12939 17855 12973 17889
rect 13007 17855 13041 17889
rect 13075 17855 13109 17889
rect 13143 17855 13177 17889
rect 13211 17855 13245 17889
rect 13279 17855 13313 17889
rect 13347 17855 13381 17889
rect 13415 17855 13449 17889
rect 13483 17855 13517 17889
rect 13551 17855 13585 17889
rect 13619 17855 13653 17889
rect 13687 17855 13721 17889
rect 13755 17855 13789 17889
rect 13823 17855 13857 17889
rect 13891 17855 13925 17889
rect 13959 17855 13993 17889
rect 14027 17855 14061 17889
rect 14095 17855 14129 17889
rect 14163 17855 14197 17889
rect 14231 17855 14265 17889
rect 14299 17855 14333 17889
rect 14367 17855 14401 17889
rect 14435 17855 14469 17889
rect 14503 17855 14537 17889
rect 14571 17855 14605 17889
rect 14639 17855 14673 17889
rect 14707 17855 14741 17889
<< mvnsubdiffcont >>
rect 83 27342 117 27376
rect 152 27342 186 27376
rect 221 27342 255 27376
rect 290 27342 324 27376
rect 359 27342 393 27376
rect 428 27342 462 27376
rect 497 27342 531 27376
rect 566 27342 600 27376
rect 635 27342 669 27376
rect 704 27342 738 27376
rect 773 27342 807 27376
rect 842 27342 876 27376
rect 911 27342 945 27376
rect 980 27342 1014 27376
rect 1049 27342 1083 27376
rect 1118 27342 1152 27376
rect 1187 27342 1221 27376
rect 1256 27342 1290 27376
rect 1325 27342 1359 27376
rect 1394 27342 1428 27376
rect 1463 27342 1497 27376
rect 1532 27342 1566 27376
rect 1601 27342 1635 27376
rect 1670 27342 1704 27376
rect 1739 27342 1773 27376
rect 1808 27342 1842 27376
rect 1877 27342 1911 27376
rect 1946 27342 1980 27376
rect 2014 27342 2048 27376
rect 2082 27342 2116 27376
rect 2150 27342 2184 27376
rect 2218 27342 2252 27376
rect 2286 27342 2320 27376
rect 2354 27342 2388 27376
rect 2422 27342 2456 27376
rect 2490 27342 2524 27376
rect 2558 27342 2592 27376
rect 2626 27342 2660 27376
rect 2694 27342 2728 27376
rect 2762 27342 2796 27376
rect 2848 27338 2882 27372
rect 2916 27338 2950 27372
rect 2984 27338 3018 27372
rect 3052 27338 3086 27372
rect 3120 27338 3154 27372
rect 3188 27338 3222 27372
rect 3256 27338 3290 27372
rect 3324 27338 3358 27372
rect 3392 27338 3426 27372
rect 3460 27338 3494 27372
rect 3528 27338 3562 27372
rect 3596 27338 3630 27372
rect 3664 27338 3698 27372
rect 3732 27338 3766 27372
rect 3800 27338 3834 27372
rect 3868 27338 3902 27372
rect 3936 27338 3970 27372
rect 4004 27338 4038 27372
rect 4072 27338 4106 27372
rect 4140 27338 4174 27372
rect 4208 27338 4242 27372
rect 4276 27338 4310 27372
rect 4344 27338 4378 27372
rect 4412 27338 4446 27372
rect 4480 27338 4514 27372
rect 4548 27338 4582 27372
rect 4616 27338 4650 27372
rect 4684 27338 4718 27372
rect 4752 27338 4786 27372
rect 4820 27338 4854 27372
rect 4888 27338 4922 27372
rect 4956 27338 4990 27372
rect 5024 27338 5058 27372
rect 5092 27338 5126 27372
rect 5160 27338 5194 27372
rect 5228 27338 5262 27372
rect 5296 27338 5330 27372
rect 5364 27338 5398 27372
rect 5432 27338 5466 27372
rect 5500 27338 5534 27372
rect 5568 27338 5602 27372
rect 5636 27338 5670 27372
rect 5704 27338 5738 27372
rect 5772 27338 5806 27372
rect 5840 27338 5874 27372
rect 5908 27338 5942 27372
rect 5976 27338 6010 27372
rect 6044 27338 6078 27372
rect 6112 27338 6146 27372
rect 6180 27338 6214 27372
rect 6248 27338 6282 27372
rect 6316 27338 6350 27372
rect 6384 27338 6418 27372
rect 6452 27338 6486 27372
rect 6520 27338 6554 27372
rect 6588 27338 6622 27372
rect 6656 27338 6690 27372
rect 6724 27338 6758 27372
rect 6792 27338 6826 27372
rect 6860 27338 6894 27372
rect 6928 27338 6962 27372
rect 6996 27338 7030 27372
rect 7064 27338 7098 27372
rect 7132 27338 7166 27372
rect 7200 27338 7234 27372
rect 7268 27338 7302 27372
rect 7336 27338 7370 27372
rect 7404 27338 7438 27372
rect 7472 27338 7506 27372
rect 7540 27338 7574 27372
rect 7608 27338 7642 27372
rect 7676 27338 7710 27372
rect 7744 27338 7778 27372
rect 7812 27338 7846 27372
rect 7880 27338 7914 27372
rect 7948 27338 7982 27372
rect 8016 27338 8050 27372
rect 8084 27338 8118 27372
rect 8152 27338 8186 27372
rect 8220 27338 8254 27372
rect 8288 27338 8322 27372
rect 8356 27338 8390 27372
rect 8424 27338 8458 27372
rect 8492 27338 8526 27372
rect 8560 27338 8594 27372
rect 8628 27338 8662 27372
rect 8696 27338 8730 27372
rect 8764 27338 8798 27372
rect 8832 27338 8866 27372
rect 8900 27338 8934 27372
rect 8968 27338 9002 27372
rect 9036 27338 9070 27372
rect 9104 27338 9138 27372
rect 9172 27338 9206 27372
rect 9240 27338 9274 27372
rect 9308 27338 9342 27372
rect 9376 27338 9410 27372
rect 9444 27338 9478 27372
rect 9512 27338 9546 27372
rect 9580 27338 9614 27372
rect 9648 27338 9682 27372
rect 9716 27338 9750 27372
rect 9784 27338 9818 27372
rect 9852 27338 9886 27372
rect 9920 27338 9954 27372
rect 9988 27338 10022 27372
rect 10056 27338 10090 27372
rect 10124 27338 10158 27372
rect 10192 27338 10226 27372
rect 10260 27338 10294 27372
rect 10328 27338 10362 27372
rect 10396 27338 10430 27372
rect 10464 27338 10498 27372
rect 10532 27338 10566 27372
rect 10600 27338 10634 27372
rect 10668 27338 10702 27372
rect 10736 27338 10770 27372
rect 10804 27338 10838 27372
rect 10872 27338 10906 27372
rect 10940 27338 10974 27372
rect 11008 27338 11042 27372
rect 11076 27338 11110 27372
rect 11144 27338 11178 27372
rect 11212 27338 11246 27372
rect 11280 27338 11314 27372
rect 11348 27338 11382 27372
rect 11416 27338 11450 27372
rect 11484 27338 11518 27372
rect 11552 27338 11586 27372
rect 11620 27338 11654 27372
rect 11688 27338 11722 27372
rect 11756 27338 11790 27372
rect 11824 27338 11858 27372
rect 11892 27338 11926 27372
rect 11960 27338 11994 27372
rect 12028 27338 12062 27372
rect 12096 27338 12130 27372
rect 12164 27338 12198 27372
rect 12232 27338 12266 27372
rect 12300 27338 12334 27372
rect 12368 27338 12402 27372
rect 12436 27338 12470 27372
rect 12504 27338 12538 27372
rect 12572 27338 12606 27372
rect 12640 27338 12674 27372
rect 12708 27338 12742 27372
rect 12776 27338 12810 27372
rect 12844 27338 12878 27372
rect 12912 27338 12946 27372
rect 12980 27338 13014 27372
rect 13048 27338 13082 27372
rect 13116 27338 13150 27372
rect 13184 27338 13218 27372
rect 13252 27338 13286 27372
rect 13320 27338 13354 27372
rect 13388 27338 13422 27372
rect 13456 27338 13490 27372
rect 13524 27338 13558 27372
rect 13592 27338 13626 27372
rect 13660 27338 13694 27372
rect 13728 27338 13762 27372
rect 13796 27338 13830 27372
rect 13864 27338 13898 27372
rect 13932 27338 13966 27372
rect 14000 27338 14034 27372
rect 14068 27338 14102 27372
rect 14136 27338 14170 27372
rect 14204 27338 14238 27372
rect 14272 27338 14306 27372
rect 14340 27338 14374 27372
rect 14408 27338 14442 27372
rect 14476 27338 14510 27372
rect 14544 27338 14578 27372
rect 14612 27338 14646 27372
rect 14680 27338 14714 27372
rect 14748 27338 14782 27372
rect 14816 27338 14850 27372
rect 14884 27338 14918 27372
rect 83 27268 117 27302
rect 152 27268 186 27302
rect 221 27268 255 27302
rect 290 27268 324 27302
rect 359 27268 393 27302
rect 428 27268 462 27302
rect 497 27268 531 27302
rect 566 27268 600 27302
rect 635 27268 669 27302
rect 704 27268 738 27302
rect 773 27268 807 27302
rect 842 27268 876 27302
rect 911 27268 945 27302
rect 980 27268 1014 27302
rect 1049 27268 1083 27302
rect 1118 27268 1152 27302
rect 1187 27268 1221 27302
rect 1256 27268 1290 27302
rect 1325 27268 1359 27302
rect 1394 27268 1428 27302
rect 1463 27268 1497 27302
rect 1532 27268 1566 27302
rect 1601 27268 1635 27302
rect 1670 27268 1704 27302
rect 1739 27268 1773 27302
rect 1808 27268 1842 27302
rect 1877 27268 1911 27302
rect 1946 27268 1980 27302
rect 2014 27268 2048 27302
rect 2082 27268 2116 27302
rect 2150 27268 2184 27302
rect 2218 27268 2252 27302
rect 2286 27268 2320 27302
rect 2354 27268 2388 27302
rect 2422 27268 2456 27302
rect 2490 27268 2524 27302
rect 2558 27268 2592 27302
rect 2626 27268 2660 27302
rect 2694 27268 2728 27302
rect 2762 27268 2796 27302
rect 2848 27268 2882 27302
rect 2916 27268 2950 27302
rect 2984 27268 3018 27302
rect 3052 27268 3086 27302
rect 3120 27268 3154 27302
rect 3188 27268 3222 27302
rect 3256 27268 3290 27302
rect 3324 27268 3358 27302
rect 3392 27268 3426 27302
rect 3460 27268 3494 27302
rect 3528 27268 3562 27302
rect 3596 27268 3630 27302
rect 3664 27268 3698 27302
rect 3732 27268 3766 27302
rect 3800 27268 3834 27302
rect 3868 27268 3902 27302
rect 3936 27268 3970 27302
rect 4004 27268 4038 27302
rect 4072 27268 4106 27302
rect 4140 27268 4174 27302
rect 4208 27268 4242 27302
rect 4276 27268 4310 27302
rect 4344 27268 4378 27302
rect 4412 27268 4446 27302
rect 4480 27268 4514 27302
rect 4548 27268 4582 27302
rect 4616 27268 4650 27302
rect 4684 27268 4718 27302
rect 4752 27268 4786 27302
rect 4820 27268 4854 27302
rect 4888 27268 4922 27302
rect 4956 27268 4990 27302
rect 5024 27268 5058 27302
rect 5092 27268 5126 27302
rect 5160 27268 5194 27302
rect 5228 27268 5262 27302
rect 5296 27268 5330 27302
rect 5364 27268 5398 27302
rect 5432 27268 5466 27302
rect 5500 27268 5534 27302
rect 5568 27268 5602 27302
rect 5636 27268 5670 27302
rect 5704 27268 5738 27302
rect 5772 27268 5806 27302
rect 5840 27268 5874 27302
rect 5908 27268 5942 27302
rect 5976 27268 6010 27302
rect 6044 27268 6078 27302
rect 6112 27268 6146 27302
rect 6180 27268 6214 27302
rect 6248 27268 6282 27302
rect 6316 27268 6350 27302
rect 6384 27268 6418 27302
rect 6452 27268 6486 27302
rect 6520 27268 6554 27302
rect 6588 27268 6622 27302
rect 6656 27268 6690 27302
rect 6724 27268 6758 27302
rect 6792 27268 6826 27302
rect 6860 27268 6894 27302
rect 6928 27268 6962 27302
rect 6996 27268 7030 27302
rect 7064 27268 7098 27302
rect 7132 27268 7166 27302
rect 7200 27268 7234 27302
rect 7268 27268 7302 27302
rect 7336 27268 7370 27302
rect 7404 27268 7438 27302
rect 7472 27268 7506 27302
rect 7540 27268 7574 27302
rect 7608 27268 7642 27302
rect 7676 27268 7710 27302
rect 7744 27268 7778 27302
rect 7812 27268 7846 27302
rect 7880 27268 7914 27302
rect 7948 27268 7982 27302
rect 8016 27268 8050 27302
rect 8084 27268 8118 27302
rect 8152 27268 8186 27302
rect 8220 27268 8254 27302
rect 8288 27268 8322 27302
rect 8356 27268 8390 27302
rect 8424 27268 8458 27302
rect 8492 27268 8526 27302
rect 8560 27268 8594 27302
rect 8628 27268 8662 27302
rect 8696 27268 8730 27302
rect 8764 27268 8798 27302
rect 8832 27268 8866 27302
rect 8900 27268 8934 27302
rect 8968 27268 9002 27302
rect 9036 27268 9070 27302
rect 9104 27268 9138 27302
rect 9172 27268 9206 27302
rect 9240 27268 9274 27302
rect 9308 27268 9342 27302
rect 9376 27268 9410 27302
rect 9444 27268 9478 27302
rect 9512 27268 9546 27302
rect 9580 27268 9614 27302
rect 9648 27268 9682 27302
rect 9716 27268 9750 27302
rect 9784 27268 9818 27302
rect 9852 27268 9886 27302
rect 9920 27268 9954 27302
rect 9988 27268 10022 27302
rect 10056 27268 10090 27302
rect 10124 27268 10158 27302
rect 10192 27268 10226 27302
rect 10260 27268 10294 27302
rect 10328 27268 10362 27302
rect 10396 27268 10430 27302
rect 10464 27268 10498 27302
rect 10532 27268 10566 27302
rect 10600 27268 10634 27302
rect 10668 27268 10702 27302
rect 10736 27268 10770 27302
rect 10804 27268 10838 27302
rect 10872 27268 10906 27302
rect 10940 27268 10974 27302
rect 11008 27268 11042 27302
rect 11076 27268 11110 27302
rect 11144 27268 11178 27302
rect 11212 27268 11246 27302
rect 11280 27268 11314 27302
rect 11348 27268 11382 27302
rect 11416 27268 11450 27302
rect 11484 27268 11518 27302
rect 11552 27268 11586 27302
rect 11620 27268 11654 27302
rect 11688 27268 11722 27302
rect 11756 27268 11790 27302
rect 11824 27268 11858 27302
rect 11892 27268 11926 27302
rect 11960 27268 11994 27302
rect 12028 27268 12062 27302
rect 12096 27268 12130 27302
rect 12164 27268 12198 27302
rect 12232 27268 12266 27302
rect 12300 27268 12334 27302
rect 12368 27268 12402 27302
rect 12436 27268 12470 27302
rect 12504 27268 12538 27302
rect 12572 27268 12606 27302
rect 12640 27268 12674 27302
rect 12708 27268 12742 27302
rect 12776 27268 12810 27302
rect 12844 27268 12878 27302
rect 12912 27268 12946 27302
rect 12980 27268 13014 27302
rect 13048 27268 13082 27302
rect 13116 27268 13150 27302
rect 13184 27268 13218 27302
rect 13252 27268 13286 27302
rect 13320 27268 13354 27302
rect 13388 27268 13422 27302
rect 13456 27268 13490 27302
rect 13524 27268 13558 27302
rect 13592 27268 13626 27302
rect 13660 27268 13694 27302
rect 13728 27268 13762 27302
rect 13796 27268 13830 27302
rect 13864 27268 13898 27302
rect 13932 27268 13966 27302
rect 14000 27268 14034 27302
rect 14068 27268 14102 27302
rect 14136 27268 14170 27302
rect 14204 27268 14238 27302
rect 14272 27268 14306 27302
rect 14340 27268 14374 27302
rect 14408 27268 14442 27302
rect 14476 27268 14510 27302
rect 14544 27268 14578 27302
rect 14612 27268 14646 27302
rect 14680 27268 14714 27302
rect 14748 27268 14782 27302
rect 14816 27268 14850 27302
rect 14884 27268 14918 27302
rect 83 27194 117 27228
rect 152 27194 186 27228
rect 221 27194 255 27228
rect 290 27194 324 27228
rect 359 27194 393 27228
rect 428 27194 462 27228
rect 497 27194 531 27228
rect 566 27194 600 27228
rect 635 27194 669 27228
rect 704 27194 738 27228
rect 773 27194 807 27228
rect 842 27194 876 27228
rect 911 27194 945 27228
rect 980 27194 1014 27228
rect 1049 27194 1083 27228
rect 1118 27194 1152 27228
rect 1187 27194 1221 27228
rect 1256 27194 1290 27228
rect 1325 27194 1359 27228
rect 1394 27194 1428 27228
rect 1463 27194 1497 27228
rect 1532 27194 1566 27228
rect 1601 27194 1635 27228
rect 1670 27194 1704 27228
rect 1739 27194 1773 27228
rect 1808 27194 1842 27228
rect 1877 27194 1911 27228
rect 1946 27194 1980 27228
rect 2014 27194 2048 27228
rect 2082 27194 2116 27228
rect 2150 27194 2184 27228
rect 2218 27194 2252 27228
rect 2286 27194 2320 27228
rect 2354 27194 2388 27228
rect 2422 27194 2456 27228
rect 2490 27194 2524 27228
rect 2558 27194 2592 27228
rect 2626 27194 2660 27228
rect 2694 27194 2728 27228
rect 2762 27194 2796 27228
rect 2848 27198 2882 27232
rect 2916 27198 2950 27232
rect 2984 27198 3018 27232
rect 3052 27198 3086 27232
rect 3120 27198 3154 27232
rect 3188 27198 3222 27232
rect 3256 27198 3290 27232
rect 3324 27198 3358 27232
rect 3392 27198 3426 27232
rect 3460 27198 3494 27232
rect 3528 27198 3562 27232
rect 3596 27198 3630 27232
rect 3664 27198 3698 27232
rect 3732 27198 3766 27232
rect 3800 27198 3834 27232
rect 3868 27198 3902 27232
rect 3936 27198 3970 27232
rect 4004 27198 4038 27232
rect 4072 27198 4106 27232
rect 4140 27198 4174 27232
rect 4208 27198 4242 27232
rect 4276 27198 4310 27232
rect 4344 27198 4378 27232
rect 4412 27198 4446 27232
rect 4480 27198 4514 27232
rect 4548 27198 4582 27232
rect 4616 27198 4650 27232
rect 4684 27198 4718 27232
rect 4752 27198 4786 27232
rect 4820 27198 4854 27232
rect 4888 27198 4922 27232
rect 4956 27198 4990 27232
rect 5024 27198 5058 27232
rect 5092 27198 5126 27232
rect 5160 27198 5194 27232
rect 5228 27198 5262 27232
rect 5296 27198 5330 27232
rect 5364 27198 5398 27232
rect 5432 27198 5466 27232
rect 5500 27198 5534 27232
rect 5568 27198 5602 27232
rect 5636 27198 5670 27232
rect 5704 27198 5738 27232
rect 5772 27198 5806 27232
rect 5840 27198 5874 27232
rect 5908 27198 5942 27232
rect 5976 27198 6010 27232
rect 6044 27198 6078 27232
rect 6112 27198 6146 27232
rect 6180 27198 6214 27232
rect 6248 27198 6282 27232
rect 6316 27198 6350 27232
rect 6384 27198 6418 27232
rect 6452 27198 6486 27232
rect 6520 27198 6554 27232
rect 6588 27198 6622 27232
rect 6656 27198 6690 27232
rect 6724 27198 6758 27232
rect 6792 27198 6826 27232
rect 6860 27198 6894 27232
rect 6928 27198 6962 27232
rect 6996 27198 7030 27232
rect 7064 27198 7098 27232
rect 7132 27198 7166 27232
rect 7200 27198 7234 27232
rect 7268 27198 7302 27232
rect 7336 27198 7370 27232
rect 7404 27198 7438 27232
rect 7472 27198 7506 27232
rect 7540 27198 7574 27232
rect 7608 27198 7642 27232
rect 7676 27198 7710 27232
rect 7744 27198 7778 27232
rect 7812 27198 7846 27232
rect 7880 27198 7914 27232
rect 7948 27198 7982 27232
rect 8016 27198 8050 27232
rect 8084 27198 8118 27232
rect 8152 27198 8186 27232
rect 8220 27198 8254 27232
rect 8288 27198 8322 27232
rect 8356 27198 8390 27232
rect 8424 27198 8458 27232
rect 8492 27198 8526 27232
rect 8560 27198 8594 27232
rect 8628 27198 8662 27232
rect 8696 27198 8730 27232
rect 8764 27198 8798 27232
rect 8832 27198 8866 27232
rect 8900 27198 8934 27232
rect 8968 27198 9002 27232
rect 9036 27198 9070 27232
rect 9104 27198 9138 27232
rect 9172 27198 9206 27232
rect 9240 27198 9274 27232
rect 9308 27198 9342 27232
rect 9376 27198 9410 27232
rect 9444 27198 9478 27232
rect 9512 27198 9546 27232
rect 9580 27198 9614 27232
rect 9648 27198 9682 27232
rect 9716 27198 9750 27232
rect 9784 27198 9818 27232
rect 9852 27198 9886 27232
rect 9920 27198 9954 27232
rect 9988 27198 10022 27232
rect 10056 27198 10090 27232
rect 10124 27198 10158 27232
rect 10192 27198 10226 27232
rect 10260 27198 10294 27232
rect 10328 27198 10362 27232
rect 10396 27198 10430 27232
rect 10464 27198 10498 27232
rect 10532 27198 10566 27232
rect 10600 27198 10634 27232
rect 10668 27198 10702 27232
rect 10736 27198 10770 27232
rect 10804 27198 10838 27232
rect 10872 27198 10906 27232
rect 10940 27198 10974 27232
rect 11008 27198 11042 27232
rect 11076 27198 11110 27232
rect 11144 27198 11178 27232
rect 11212 27198 11246 27232
rect 11280 27198 11314 27232
rect 11348 27198 11382 27232
rect 11416 27198 11450 27232
rect 11484 27198 11518 27232
rect 11552 27198 11586 27232
rect 11620 27198 11654 27232
rect 11688 27198 11722 27232
rect 11756 27198 11790 27232
rect 11824 27198 11858 27232
rect 11892 27198 11926 27232
rect 11960 27198 11994 27232
rect 12028 27198 12062 27232
rect 12096 27198 12130 27232
rect 12164 27198 12198 27232
rect 12232 27198 12266 27232
rect 12300 27198 12334 27232
rect 12368 27198 12402 27232
rect 12436 27198 12470 27232
rect 12504 27198 12538 27232
rect 12572 27198 12606 27232
rect 12640 27198 12674 27232
rect 12708 27198 12742 27232
rect 12776 27198 12810 27232
rect 12844 27198 12878 27232
rect 12912 27198 12946 27232
rect 12980 27198 13014 27232
rect 13048 27198 13082 27232
rect 13116 27198 13150 27232
rect 13184 27198 13218 27232
rect 13252 27198 13286 27232
rect 13320 27198 13354 27232
rect 13388 27198 13422 27232
rect 13456 27198 13490 27232
rect 13524 27198 13558 27232
rect 13592 27198 13626 27232
rect 13660 27198 13694 27232
rect 13728 27198 13762 27232
rect 13796 27198 13830 27232
rect 13864 27198 13898 27232
rect 13932 27198 13966 27232
rect 14000 27198 14034 27232
rect 14068 27198 14102 27232
rect 14136 27198 14170 27232
rect 14204 27198 14238 27232
rect 14272 27198 14306 27232
rect 14340 27198 14374 27232
rect 14408 27198 14442 27232
rect 14476 27198 14510 27232
rect 14544 27198 14578 27232
rect 14612 27198 14646 27232
rect 14680 27198 14714 27232
rect 14748 27198 14782 27232
rect 14816 27198 14850 27232
rect 14884 27198 14918 27232
rect 83 27120 117 27154
rect 152 27120 186 27154
rect 221 27120 255 27154
rect 290 27120 324 27154
rect 359 27120 393 27154
rect 428 27120 462 27154
rect 497 27120 531 27154
rect 566 27120 600 27154
rect 635 27120 669 27154
rect 704 27120 738 27154
rect 773 27120 807 27154
rect 842 27120 876 27154
rect 911 27120 945 27154
rect 980 27120 1014 27154
rect 1049 27120 1083 27154
rect 1118 27120 1152 27154
rect 1187 27120 1221 27154
rect 1256 27120 1290 27154
rect 1325 27120 1359 27154
rect 1394 27120 1428 27154
rect 1463 27120 1497 27154
rect 1532 27120 1566 27154
rect 1601 27120 1635 27154
rect 1670 27120 1704 27154
rect 1739 27120 1773 27154
rect 1808 27120 1842 27154
rect 1877 27120 1911 27154
rect 1946 27120 1980 27154
rect 2014 27120 2048 27154
rect 2082 27120 2116 27154
rect 2150 27120 2184 27154
rect 2218 27120 2252 27154
rect 2286 27120 2320 27154
rect 2354 27120 2388 27154
rect 2422 27120 2456 27154
rect 2490 27120 2524 27154
rect 2558 27120 2592 27154
rect 2626 27120 2660 27154
rect 2694 27120 2728 27154
rect 2762 27120 2796 27154
rect 2848 27128 2882 27162
rect 2916 27128 2950 27162
rect 2984 27128 3018 27162
rect 3052 27128 3086 27162
rect 3120 27128 3154 27162
rect 3188 27128 3222 27162
rect 3256 27128 3290 27162
rect 3324 27128 3358 27162
rect 3392 27128 3426 27162
rect 3460 27128 3494 27162
rect 3528 27128 3562 27162
rect 3596 27128 3630 27162
rect 3664 27128 3698 27162
rect 3732 27128 3766 27162
rect 3800 27128 3834 27162
rect 3868 27128 3902 27162
rect 3936 27128 3970 27162
rect 4004 27128 4038 27162
rect 4072 27128 4106 27162
rect 4140 27128 4174 27162
rect 4208 27128 4242 27162
rect 4276 27128 4310 27162
rect 4344 27128 4378 27162
rect 4412 27128 4446 27162
rect 4480 27128 4514 27162
rect 4548 27128 4582 27162
rect 4616 27128 4650 27162
rect 4684 27128 4718 27162
rect 4752 27128 4786 27162
rect 4820 27128 4854 27162
rect 4888 27128 4922 27162
rect 4956 27128 4990 27162
rect 5024 27128 5058 27162
rect 5092 27128 5126 27162
rect 5160 27128 5194 27162
rect 5228 27128 5262 27162
rect 5296 27128 5330 27162
rect 5364 27128 5398 27162
rect 5432 27128 5466 27162
rect 5500 27128 5534 27162
rect 5568 27128 5602 27162
rect 5636 27128 5670 27162
rect 5704 27128 5738 27162
rect 5772 27128 5806 27162
rect 5840 27128 5874 27162
rect 5908 27128 5942 27162
rect 5976 27128 6010 27162
rect 6044 27128 6078 27162
rect 6112 27128 6146 27162
rect 6180 27128 6214 27162
rect 6248 27128 6282 27162
rect 6316 27128 6350 27162
rect 6384 27128 6418 27162
rect 6452 27128 6486 27162
rect 6520 27128 6554 27162
rect 6588 27128 6622 27162
rect 6656 27128 6690 27162
rect 6724 27128 6758 27162
rect 6792 27128 6826 27162
rect 6860 27128 6894 27162
rect 6928 27128 6962 27162
rect 6996 27128 7030 27162
rect 7064 27128 7098 27162
rect 7132 27128 7166 27162
rect 7200 27128 7234 27162
rect 7268 27128 7302 27162
rect 7336 27128 7370 27162
rect 7404 27128 7438 27162
rect 7472 27128 7506 27162
rect 7540 27128 7574 27162
rect 7608 27128 7642 27162
rect 7676 27128 7710 27162
rect 7744 27128 7778 27162
rect 7812 27128 7846 27162
rect 7880 27128 7914 27162
rect 7948 27128 7982 27162
rect 8016 27128 8050 27162
rect 8084 27128 8118 27162
rect 8152 27128 8186 27162
rect 8220 27128 8254 27162
rect 8288 27128 8322 27162
rect 8356 27128 8390 27162
rect 8424 27128 8458 27162
rect 8492 27128 8526 27162
rect 8560 27128 8594 27162
rect 8628 27128 8662 27162
rect 8696 27128 8730 27162
rect 8764 27128 8798 27162
rect 8832 27128 8866 27162
rect 8900 27128 8934 27162
rect 8968 27128 9002 27162
rect 9036 27128 9070 27162
rect 9104 27128 9138 27162
rect 9172 27128 9206 27162
rect 9240 27128 9274 27162
rect 9308 27128 9342 27162
rect 9376 27128 9410 27162
rect 9444 27128 9478 27162
rect 9512 27128 9546 27162
rect 9580 27128 9614 27162
rect 9648 27128 9682 27162
rect 9716 27128 9750 27162
rect 9784 27128 9818 27162
rect 9852 27128 9886 27162
rect 9920 27128 9954 27162
rect 9988 27128 10022 27162
rect 10056 27128 10090 27162
rect 10124 27128 10158 27162
rect 10192 27128 10226 27162
rect 10260 27128 10294 27162
rect 10328 27128 10362 27162
rect 10396 27128 10430 27162
rect 10464 27128 10498 27162
rect 10532 27128 10566 27162
rect 10600 27128 10634 27162
rect 10668 27128 10702 27162
rect 10736 27128 10770 27162
rect 10804 27128 10838 27162
rect 10872 27128 10906 27162
rect 10940 27128 10974 27162
rect 11008 27128 11042 27162
rect 11076 27128 11110 27162
rect 11144 27128 11178 27162
rect 11212 27128 11246 27162
rect 11280 27128 11314 27162
rect 11348 27128 11382 27162
rect 11416 27128 11450 27162
rect 11484 27128 11518 27162
rect 11552 27128 11586 27162
rect 11620 27128 11654 27162
rect 11688 27128 11722 27162
rect 11756 27128 11790 27162
rect 11824 27128 11858 27162
rect 11892 27128 11926 27162
rect 11960 27128 11994 27162
rect 12028 27128 12062 27162
rect 12096 27128 12130 27162
rect 12164 27128 12198 27162
rect 12232 27128 12266 27162
rect 12300 27128 12334 27162
rect 12368 27128 12402 27162
rect 12436 27128 12470 27162
rect 12504 27128 12538 27162
rect 12572 27128 12606 27162
rect 12640 27128 12674 27162
rect 12708 27128 12742 27162
rect 12776 27128 12810 27162
rect 12844 27128 12878 27162
rect 12912 27128 12946 27162
rect 12980 27128 13014 27162
rect 13048 27128 13082 27162
rect 13116 27128 13150 27162
rect 13184 27128 13218 27162
rect 13252 27128 13286 27162
rect 13320 27128 13354 27162
rect 13388 27128 13422 27162
rect 13456 27128 13490 27162
rect 13524 27128 13558 27162
rect 13592 27128 13626 27162
rect 13660 27128 13694 27162
rect 13728 27128 13762 27162
rect 13796 27128 13830 27162
rect 13864 27128 13898 27162
rect 13932 27128 13966 27162
rect 14000 27128 14034 27162
rect 14068 27128 14102 27162
rect 14136 27128 14170 27162
rect 14204 27128 14238 27162
rect 14272 27128 14306 27162
rect 14340 27128 14374 27162
rect 14408 27128 14442 27162
rect 14476 27128 14510 27162
rect 14544 27128 14578 27162
rect 14612 27128 14646 27162
rect 14680 27128 14714 27162
rect 14748 27128 14782 27162
rect 14816 27128 14850 27162
rect 14884 27128 14918 27162
rect 2848 27058 2882 27092
rect 2916 27058 2950 27092
rect 2984 27058 3018 27092
rect 3052 27058 3086 27092
rect 3120 27058 3154 27092
rect 3188 27058 3222 27092
rect 3256 27058 3290 27092
rect 3324 27058 3358 27092
rect 3392 27058 3426 27092
rect 3460 27058 3494 27092
rect 3528 27058 3562 27092
rect 3596 27058 3630 27092
rect 3664 27058 3698 27092
rect 3732 27058 3766 27092
rect 3800 27058 3834 27092
rect 3868 27058 3902 27092
rect 3936 27058 3970 27092
rect 4004 27058 4038 27092
rect 4072 27058 4106 27092
rect 4140 27058 4174 27092
rect 4208 27058 4242 27092
rect 4276 27058 4310 27092
rect 4344 27058 4378 27092
rect 4412 27058 4446 27092
rect 4480 27058 4514 27092
rect 4548 27058 4582 27092
rect 4616 27058 4650 27092
rect 4684 27058 4718 27092
rect 4752 27058 4786 27092
rect 4820 27058 4854 27092
rect 4888 27058 4922 27092
rect 4956 27058 4990 27092
rect 5024 27058 5058 27092
rect 5092 27058 5126 27092
rect 5160 27058 5194 27092
rect 5228 27058 5262 27092
rect 5296 27058 5330 27092
rect 5364 27058 5398 27092
rect 5432 27058 5466 27092
rect 5500 27058 5534 27092
rect 5568 27058 5602 27092
rect 5636 27058 5670 27092
rect 5704 27058 5738 27092
rect 5772 27058 5806 27092
rect 5840 27058 5874 27092
rect 5908 27058 5942 27092
rect 5976 27058 6010 27092
rect 6044 27058 6078 27092
rect 6112 27058 6146 27092
rect 6180 27058 6214 27092
rect 6248 27058 6282 27092
rect 6316 27058 6350 27092
rect 6384 27058 6418 27092
rect 6452 27058 6486 27092
rect 6520 27058 6554 27092
rect 6588 27058 6622 27092
rect 6656 27058 6690 27092
rect 6724 27058 6758 27092
rect 6792 27058 6826 27092
rect 6860 27058 6894 27092
rect 6928 27058 6962 27092
rect 6996 27058 7030 27092
rect 7064 27058 7098 27092
rect 7132 27058 7166 27092
rect 7200 27058 7234 27092
rect 7268 27058 7302 27092
rect 7336 27058 7370 27092
rect 7404 27058 7438 27092
rect 7472 27058 7506 27092
rect 7540 27058 7574 27092
rect 7608 27058 7642 27092
rect 7676 27058 7710 27092
rect 7744 27058 7778 27092
rect 7812 27058 7846 27092
rect 7880 27058 7914 27092
rect 7948 27058 7982 27092
rect 8016 27058 8050 27092
rect 8084 27058 8118 27092
rect 8152 27058 8186 27092
rect 8220 27058 8254 27092
rect 8288 27058 8322 27092
rect 8356 27058 8390 27092
rect 8424 27058 8458 27092
rect 8492 27058 8526 27092
rect 8560 27058 8594 27092
rect 8628 27058 8662 27092
rect 8696 27058 8730 27092
rect 8764 27058 8798 27092
rect 8832 27058 8866 27092
rect 8900 27058 8934 27092
rect 8968 27058 9002 27092
rect 9036 27058 9070 27092
rect 9104 27058 9138 27092
rect 9172 27058 9206 27092
rect 9240 27058 9274 27092
rect 9308 27058 9342 27092
rect 9376 27058 9410 27092
rect 9444 27058 9478 27092
rect 9512 27058 9546 27092
rect 9580 27058 9614 27092
rect 9648 27058 9682 27092
rect 9716 27058 9750 27092
rect 9784 27058 9818 27092
rect 9852 27058 9886 27092
rect 9920 27058 9954 27092
rect 9988 27058 10022 27092
rect 10056 27058 10090 27092
rect 10124 27058 10158 27092
rect 10192 27058 10226 27092
rect 10260 27058 10294 27092
rect 10328 27058 10362 27092
rect 10396 27058 10430 27092
rect 10464 27058 10498 27092
rect 10532 27058 10566 27092
rect 10600 27058 10634 27092
rect 10668 27058 10702 27092
rect 10736 27058 10770 27092
rect 10804 27058 10838 27092
rect 10872 27058 10906 27092
rect 10940 27058 10974 27092
rect 11008 27058 11042 27092
rect 11076 27058 11110 27092
rect 11144 27058 11178 27092
rect 11212 27058 11246 27092
rect 11280 27058 11314 27092
rect 11348 27058 11382 27092
rect 11416 27058 11450 27092
rect 11484 27058 11518 27092
rect 11552 27058 11586 27092
rect 11620 27058 11654 27092
rect 11688 27058 11722 27092
rect 11756 27058 11790 27092
rect 11824 27058 11858 27092
rect 11892 27058 11926 27092
rect 11960 27058 11994 27092
rect 12028 27058 12062 27092
rect 12096 27058 12130 27092
rect 12164 27058 12198 27092
rect 12232 27058 12266 27092
rect 12300 27058 12334 27092
rect 12368 27058 12402 27092
rect 12436 27058 12470 27092
rect 12504 27058 12538 27092
rect 12572 27058 12606 27092
rect 12640 27058 12674 27092
rect 12708 27058 12742 27092
rect 12776 27058 12810 27092
rect 12844 27058 12878 27092
rect 12912 27058 12946 27092
rect 12980 27058 13014 27092
rect 13048 27058 13082 27092
rect 13116 27058 13150 27092
rect 13184 27058 13218 27092
rect 13252 27058 13286 27092
rect 13320 27058 13354 27092
rect 13388 27058 13422 27092
rect 13456 27058 13490 27092
rect 13524 27058 13558 27092
rect 13592 27058 13626 27092
rect 13660 27058 13694 27092
rect 13728 27058 13762 27092
rect 13796 27058 13830 27092
rect 13864 27058 13898 27092
rect 13932 27058 13966 27092
rect 14000 27058 14034 27092
rect 14068 27058 14102 27092
rect 14136 27058 14170 27092
rect 14204 27058 14238 27092
rect 14272 27058 14306 27092
rect 14340 27058 14374 27092
rect 14408 27058 14442 27092
rect 14476 27058 14510 27092
rect 14544 27058 14578 27092
rect 14612 27058 14646 27092
rect 14680 27058 14714 27092
rect 14748 27058 14782 27092
rect 14816 27058 14850 27092
rect 14884 27058 14918 27092
rect 2848 26988 2882 27022
rect 2916 26988 2950 27022
rect 2984 26988 3018 27022
rect 3052 26988 3086 27022
rect 3120 26988 3154 27022
rect 3188 26988 3222 27022
rect 3256 26988 3290 27022
rect 3324 26988 3358 27022
rect 3392 26988 3426 27022
rect 3460 26988 3494 27022
rect 3528 26988 3562 27022
rect 3596 26988 3630 27022
rect 3664 26988 3698 27022
rect 3732 26988 3766 27022
rect 3800 26988 3834 27022
rect 3868 26988 3902 27022
rect 3936 26988 3970 27022
rect 4004 26988 4038 27022
rect 4072 26988 4106 27022
rect 4140 26988 4174 27022
rect 4208 26988 4242 27022
rect 4276 26988 4310 27022
rect 4344 26988 4378 27022
rect 4412 26988 4446 27022
rect 4480 26988 4514 27022
rect 4548 26988 4582 27022
rect 4616 26988 4650 27022
rect 4684 26988 4718 27022
rect 4752 26988 4786 27022
rect 4820 26988 4854 27022
rect 4888 26988 4922 27022
rect 4956 26988 4990 27022
rect 5024 26988 5058 27022
rect 5092 26988 5126 27022
rect 5160 26988 5194 27022
rect 5228 26988 5262 27022
rect 5296 26988 5330 27022
rect 5364 26988 5398 27022
rect 5432 26988 5466 27022
rect 5500 26988 5534 27022
rect 5568 26988 5602 27022
rect 5636 26988 5670 27022
rect 5704 26988 5738 27022
rect 5772 26988 5806 27022
rect 5840 26988 5874 27022
rect 5908 26988 5942 27022
rect 5976 26988 6010 27022
rect 6044 26988 6078 27022
rect 6112 26988 6146 27022
rect 6180 26988 6214 27022
rect 6248 26988 6282 27022
rect 6316 26988 6350 27022
rect 6384 26988 6418 27022
rect 6452 26988 6486 27022
rect 6520 26988 6554 27022
rect 6588 26988 6622 27022
rect 6656 26988 6690 27022
rect 6724 26988 6758 27022
rect 6792 26988 6826 27022
rect 6860 26988 6894 27022
rect 6928 26988 6962 27022
rect 6996 26988 7030 27022
rect 7064 26988 7098 27022
rect 7132 26988 7166 27022
rect 7200 26988 7234 27022
rect 7268 26988 7302 27022
rect 7336 26988 7370 27022
rect 7404 26988 7438 27022
rect 7472 26988 7506 27022
rect 7540 26988 7574 27022
rect 7608 26988 7642 27022
rect 7676 26988 7710 27022
rect 7744 26988 7778 27022
rect 7812 26988 7846 27022
rect 7880 26988 7914 27022
rect 7948 26988 7982 27022
rect 8016 26988 8050 27022
rect 8084 26988 8118 27022
rect 8152 26988 8186 27022
rect 8220 26988 8254 27022
rect 8288 26988 8322 27022
rect 8356 26988 8390 27022
rect 8424 26988 8458 27022
rect 8492 26988 8526 27022
rect 8560 26988 8594 27022
rect 8628 26988 8662 27022
rect 8696 26988 8730 27022
rect 8764 26988 8798 27022
rect 8832 26988 8866 27022
rect 8900 26988 8934 27022
rect 8968 26988 9002 27022
rect 9036 26988 9070 27022
rect 9104 26988 9138 27022
rect 9172 26988 9206 27022
rect 9240 26988 9274 27022
rect 9308 26988 9342 27022
rect 9376 26988 9410 27022
rect 9444 26988 9478 27022
rect 9512 26988 9546 27022
rect 9580 26988 9614 27022
rect 9648 26988 9682 27022
rect 9716 26988 9750 27022
rect 9784 26988 9818 27022
rect 9852 26988 9886 27022
rect 9920 26988 9954 27022
rect 9988 26988 10022 27022
rect 10056 26988 10090 27022
rect 10124 26988 10158 27022
rect 10192 26988 10226 27022
rect 10260 26988 10294 27022
rect 10328 26988 10362 27022
rect 10396 26988 10430 27022
rect 10464 26988 10498 27022
rect 10532 26988 10566 27022
rect 10600 26988 10634 27022
rect 10668 26988 10702 27022
rect 10736 26988 10770 27022
rect 10804 26988 10838 27022
rect 10872 26988 10906 27022
rect 10940 26988 10974 27022
rect 11008 26988 11042 27022
rect 11076 26988 11110 27022
rect 11144 26988 11178 27022
rect 11212 26988 11246 27022
rect 11280 26988 11314 27022
rect 11348 26988 11382 27022
rect 11416 26988 11450 27022
rect 11484 26988 11518 27022
rect 11552 26988 11586 27022
rect 11620 26988 11654 27022
rect 11688 26988 11722 27022
rect 11756 26988 11790 27022
rect 11824 26988 11858 27022
rect 11892 26988 11926 27022
rect 11960 26988 11994 27022
rect 12028 26988 12062 27022
rect 12096 26988 12130 27022
rect 12164 26988 12198 27022
rect 12232 26988 12266 27022
rect 12300 26988 12334 27022
rect 12368 26988 12402 27022
rect 12436 26988 12470 27022
rect 12504 26988 12538 27022
rect 12572 26988 12606 27022
rect 12640 26988 12674 27022
rect 12708 26988 12742 27022
rect 12776 26988 12810 27022
rect 12844 26988 12878 27022
rect 12912 26988 12946 27022
rect 12980 26988 13014 27022
rect 13048 26988 13082 27022
rect 13116 26988 13150 27022
rect 13184 26988 13218 27022
rect 13252 26988 13286 27022
rect 13320 26988 13354 27022
rect 13388 26988 13422 27022
rect 13456 26988 13490 27022
rect 13524 26988 13558 27022
rect 13592 26988 13626 27022
rect 13660 26988 13694 27022
rect 13728 26988 13762 27022
rect 13796 26988 13830 27022
rect 13864 26988 13898 27022
rect 13932 26988 13966 27022
rect 14000 26988 14034 27022
rect 14068 26988 14102 27022
rect 14136 26988 14170 27022
rect 14204 26988 14238 27022
rect 14272 26988 14306 27022
rect 14340 26988 14374 27022
rect 14408 26988 14442 27022
rect 14476 26988 14510 27022
rect 14544 26988 14578 27022
rect 14612 26988 14646 27022
rect 14680 26988 14714 27022
rect 14748 26988 14782 27022
rect 14816 26988 14850 27022
rect 14884 26988 14918 27022
rect 2848 26918 2882 26952
rect 2916 26918 2950 26952
rect 2984 26918 3018 26952
rect 3052 26918 3086 26952
rect 3120 26918 3154 26952
rect 3188 26918 3222 26952
rect 3256 26918 3290 26952
rect 3324 26918 3358 26952
rect 3392 26918 3426 26952
rect 3460 26918 3494 26952
rect 3528 26918 3562 26952
rect 3596 26918 3630 26952
rect 3664 26918 3698 26952
rect 3732 26918 3766 26952
rect 3800 26918 3834 26952
rect 3868 26918 3902 26952
rect 3936 26918 3970 26952
rect 4004 26918 4038 26952
rect 4072 26918 4106 26952
rect 4140 26918 4174 26952
rect 4208 26918 4242 26952
rect 4276 26918 4310 26952
rect 4344 26918 4378 26952
rect 4412 26918 4446 26952
rect 4480 26918 4514 26952
rect 4548 26918 4582 26952
rect 4616 26918 4650 26952
rect 4684 26918 4718 26952
rect 4752 26918 4786 26952
rect 4820 26918 4854 26952
rect 4888 26918 4922 26952
rect 4956 26918 4990 26952
rect 5024 26918 5058 26952
rect 5092 26918 5126 26952
rect 5160 26918 5194 26952
rect 5228 26918 5262 26952
rect 5296 26918 5330 26952
rect 5364 26918 5398 26952
rect 5432 26918 5466 26952
rect 5500 26918 5534 26952
rect 5568 26918 5602 26952
rect 5636 26918 5670 26952
rect 5704 26918 5738 26952
rect 5772 26918 5806 26952
rect 5840 26918 5874 26952
rect 5908 26918 5942 26952
rect 5976 26918 6010 26952
rect 6044 26918 6078 26952
rect 6112 26918 6146 26952
rect 6180 26918 6214 26952
rect 6248 26918 6282 26952
rect 6316 26918 6350 26952
rect 6384 26918 6418 26952
rect 6452 26918 6486 26952
rect 6520 26918 6554 26952
rect 6588 26918 6622 26952
rect 6656 26918 6690 26952
rect 6724 26918 6758 26952
rect 6792 26918 6826 26952
rect 6860 26918 6894 26952
rect 6928 26918 6962 26952
rect 6996 26918 7030 26952
rect 7064 26918 7098 26952
rect 7132 26918 7166 26952
rect 7200 26918 7234 26952
rect 7268 26918 7302 26952
rect 7336 26918 7370 26952
rect 7404 26918 7438 26952
rect 7472 26918 7506 26952
rect 7540 26918 7574 26952
rect 7608 26918 7642 26952
rect 7676 26918 7710 26952
rect 7744 26918 7778 26952
rect 7812 26918 7846 26952
rect 7880 26918 7914 26952
rect 7948 26918 7982 26952
rect 8016 26918 8050 26952
rect 8084 26918 8118 26952
rect 8152 26918 8186 26952
rect 8220 26918 8254 26952
rect 8288 26918 8322 26952
rect 8356 26918 8390 26952
rect 8424 26918 8458 26952
rect 8492 26918 8526 26952
rect 8560 26918 8594 26952
rect 8628 26918 8662 26952
rect 8696 26918 8730 26952
rect 8764 26918 8798 26952
rect 8832 26918 8866 26952
rect 8900 26918 8934 26952
rect 8968 26918 9002 26952
rect 9036 26918 9070 26952
rect 9104 26918 9138 26952
rect 9172 26918 9206 26952
rect 9240 26918 9274 26952
rect 9308 26918 9342 26952
rect 9376 26918 9410 26952
rect 9444 26918 9478 26952
rect 9512 26918 9546 26952
rect 9580 26918 9614 26952
rect 9648 26918 9682 26952
rect 9716 26918 9750 26952
rect 9784 26918 9818 26952
rect 9852 26918 9886 26952
rect 9920 26918 9954 26952
rect 9988 26918 10022 26952
rect 10056 26918 10090 26952
rect 10124 26918 10158 26952
rect 10192 26918 10226 26952
rect 10260 26918 10294 26952
rect 10328 26918 10362 26952
rect 10396 26918 10430 26952
rect 10464 26918 10498 26952
rect 10532 26918 10566 26952
rect 10600 26918 10634 26952
rect 10668 26918 10702 26952
rect 10736 26918 10770 26952
rect 10804 26918 10838 26952
rect 10872 26918 10906 26952
rect 10940 26918 10974 26952
rect 11008 26918 11042 26952
rect 11076 26918 11110 26952
rect 11144 26918 11178 26952
rect 11212 26918 11246 26952
rect 11280 26918 11314 26952
rect 11348 26918 11382 26952
rect 11416 26918 11450 26952
rect 11484 26918 11518 26952
rect 11552 26918 11586 26952
rect 11620 26918 11654 26952
rect 11688 26918 11722 26952
rect 11756 26918 11790 26952
rect 11824 26918 11858 26952
rect 11892 26918 11926 26952
rect 11960 26918 11994 26952
rect 12028 26918 12062 26952
rect 12096 26918 12130 26952
rect 12164 26918 12198 26952
rect 12232 26918 12266 26952
rect 12300 26918 12334 26952
rect 12368 26918 12402 26952
rect 12436 26918 12470 26952
rect 12504 26918 12538 26952
rect 12572 26918 12606 26952
rect 12640 26918 12674 26952
rect 12708 26918 12742 26952
rect 12776 26918 12810 26952
rect 12844 26918 12878 26952
rect 12912 26918 12946 26952
rect 12980 26918 13014 26952
rect 13048 26918 13082 26952
rect 13116 26918 13150 26952
rect 13184 26918 13218 26952
rect 13252 26918 13286 26952
rect 13320 26918 13354 26952
rect 13388 26918 13422 26952
rect 13456 26918 13490 26952
rect 13524 26918 13558 26952
rect 13592 26918 13626 26952
rect 13660 26918 13694 26952
rect 13728 26918 13762 26952
rect 13796 26918 13830 26952
rect 13864 26918 13898 26952
rect 13932 26918 13966 26952
rect 14000 26918 14034 26952
rect 14068 26918 14102 26952
rect 14136 26918 14170 26952
rect 14204 26918 14238 26952
rect 14272 26918 14306 26952
rect 14340 26918 14374 26952
rect 14408 26918 14442 26952
rect 14476 26918 14510 26952
rect 14544 26918 14578 26952
rect 14612 26918 14646 26952
rect 14680 26918 14714 26952
rect 14748 26918 14782 26952
rect 14816 26918 14850 26952
rect 14884 26918 14918 26952
rect 2848 26848 2882 26882
rect 2916 26848 2950 26882
rect 2984 26848 3018 26882
rect 3052 26848 3086 26882
rect 3120 26848 3154 26882
rect 3188 26848 3222 26882
rect 3256 26848 3290 26882
rect 3324 26848 3358 26882
rect 3392 26848 3426 26882
rect 3460 26848 3494 26882
rect 3528 26848 3562 26882
rect 3596 26848 3630 26882
rect 3664 26848 3698 26882
rect 3732 26848 3766 26882
rect 3800 26848 3834 26882
rect 3868 26848 3902 26882
rect 3936 26848 3970 26882
rect 4004 26848 4038 26882
rect 4072 26848 4106 26882
rect 4140 26848 4174 26882
rect 4208 26848 4242 26882
rect 4276 26848 4310 26882
rect 4344 26848 4378 26882
rect 4412 26848 4446 26882
rect 4480 26848 4514 26882
rect 4548 26848 4582 26882
rect 4616 26848 4650 26882
rect 4684 26848 4718 26882
rect 4752 26848 4786 26882
rect 4820 26848 4854 26882
rect 4888 26848 4922 26882
rect 4956 26848 4990 26882
rect 5024 26848 5058 26882
rect 5092 26848 5126 26882
rect 5160 26848 5194 26882
rect 5228 26848 5262 26882
rect 5296 26848 5330 26882
rect 5364 26848 5398 26882
rect 5432 26848 5466 26882
rect 5500 26848 5534 26882
rect 5568 26848 5602 26882
rect 5636 26848 5670 26882
rect 5704 26848 5738 26882
rect 5772 26848 5806 26882
rect 5840 26848 5874 26882
rect 5908 26848 5942 26882
rect 5976 26848 6010 26882
rect 6044 26848 6078 26882
rect 6112 26848 6146 26882
rect 6180 26848 6214 26882
rect 6248 26848 6282 26882
rect 6316 26848 6350 26882
rect 6384 26848 6418 26882
rect 6452 26848 6486 26882
rect 6520 26848 6554 26882
rect 6588 26848 6622 26882
rect 6656 26848 6690 26882
rect 6724 26848 6758 26882
rect 6792 26848 6826 26882
rect 6860 26848 6894 26882
rect 6928 26848 6962 26882
rect 6996 26848 7030 26882
rect 7064 26848 7098 26882
rect 7132 26848 7166 26882
rect 7200 26848 7234 26882
rect 7268 26848 7302 26882
rect 7336 26848 7370 26882
rect 7404 26848 7438 26882
rect 7472 26848 7506 26882
rect 7540 26848 7574 26882
rect 7608 26848 7642 26882
rect 7676 26848 7710 26882
rect 7744 26848 7778 26882
rect 7812 26848 7846 26882
rect 7880 26848 7914 26882
rect 7948 26848 7982 26882
rect 8016 26848 8050 26882
rect 8084 26848 8118 26882
rect 8152 26848 8186 26882
rect 8220 26848 8254 26882
rect 8288 26848 8322 26882
rect 8356 26848 8390 26882
rect 8424 26848 8458 26882
rect 8492 26848 8526 26882
rect 8560 26848 8594 26882
rect 8628 26848 8662 26882
rect 8696 26848 8730 26882
rect 8764 26848 8798 26882
rect 8832 26848 8866 26882
rect 8900 26848 8934 26882
rect 8968 26848 9002 26882
rect 9036 26848 9070 26882
rect 9104 26848 9138 26882
rect 9172 26848 9206 26882
rect 9240 26848 9274 26882
rect 9308 26848 9342 26882
rect 9376 26848 9410 26882
rect 9444 26848 9478 26882
rect 9512 26848 9546 26882
rect 9580 26848 9614 26882
rect 9648 26848 9682 26882
rect 9716 26848 9750 26882
rect 9784 26848 9818 26882
rect 9852 26848 9886 26882
rect 9920 26848 9954 26882
rect 9988 26848 10022 26882
rect 10056 26848 10090 26882
rect 10124 26848 10158 26882
rect 10192 26848 10226 26882
rect 10260 26848 10294 26882
rect 10328 26848 10362 26882
rect 10396 26848 10430 26882
rect 10464 26848 10498 26882
rect 10532 26848 10566 26882
rect 10600 26848 10634 26882
rect 10668 26848 10702 26882
rect 10736 26848 10770 26882
rect 10804 26848 10838 26882
rect 10872 26848 10906 26882
rect 10940 26848 10974 26882
rect 11008 26848 11042 26882
rect 11076 26848 11110 26882
rect 11144 26848 11178 26882
rect 11212 26848 11246 26882
rect 11280 26848 11314 26882
rect 11348 26848 11382 26882
rect 11416 26848 11450 26882
rect 11484 26848 11518 26882
rect 11552 26848 11586 26882
rect 11620 26848 11654 26882
rect 11688 26848 11722 26882
rect 11756 26848 11790 26882
rect 11824 26848 11858 26882
rect 11892 26848 11926 26882
rect 11960 26848 11994 26882
rect 12028 26848 12062 26882
rect 12096 26848 12130 26882
rect 12164 26848 12198 26882
rect 12232 26848 12266 26882
rect 12300 26848 12334 26882
rect 12368 26848 12402 26882
rect 12436 26848 12470 26882
rect 12504 26848 12538 26882
rect 12572 26848 12606 26882
rect 12640 26848 12674 26882
rect 12708 26848 12742 26882
rect 12776 26848 12810 26882
rect 12844 26848 12878 26882
rect 12912 26848 12946 26882
rect 12980 26848 13014 26882
rect 13048 26848 13082 26882
rect 13116 26848 13150 26882
rect 13184 26848 13218 26882
rect 13252 26848 13286 26882
rect 13320 26848 13354 26882
rect 13388 26848 13422 26882
rect 13456 26848 13490 26882
rect 13524 26848 13558 26882
rect 13592 26848 13626 26882
rect 13660 26848 13694 26882
rect 13728 26848 13762 26882
rect 13796 26848 13830 26882
rect 13864 26848 13898 26882
rect 13932 26848 13966 26882
rect 14000 26848 14034 26882
rect 14068 26848 14102 26882
rect 14136 26848 14170 26882
rect 14204 26848 14238 26882
rect 14272 26848 14306 26882
rect 14340 26848 14374 26882
rect 14408 26848 14442 26882
rect 14476 26848 14510 26882
rect 14544 26848 14578 26882
rect 14612 26848 14646 26882
rect 14680 26848 14714 26882
rect 14748 26848 14782 26882
rect 14816 26848 14850 26882
rect 14884 26848 14918 26882
rect 2848 26778 2882 26812
rect 2916 26778 2950 26812
rect 2984 26778 3018 26812
rect 3052 26778 3086 26812
rect 3120 26778 3154 26812
rect 3188 26778 3222 26812
rect 3256 26778 3290 26812
rect 3324 26778 3358 26812
rect 3392 26778 3426 26812
rect 3460 26778 3494 26812
rect 3528 26778 3562 26812
rect 3596 26778 3630 26812
rect 3664 26778 3698 26812
rect 3732 26778 3766 26812
rect 3800 26778 3834 26812
rect 3868 26778 3902 26812
rect 3936 26778 3970 26812
rect 4004 26778 4038 26812
rect 4072 26778 4106 26812
rect 4140 26778 4174 26812
rect 4208 26778 4242 26812
rect 4276 26778 4310 26812
rect 4344 26778 4378 26812
rect 4412 26778 4446 26812
rect 4480 26778 4514 26812
rect 4548 26778 4582 26812
rect 4616 26778 4650 26812
rect 4684 26778 4718 26812
rect 4752 26778 4786 26812
rect 4820 26778 4854 26812
rect 4888 26778 4922 26812
rect 4956 26778 4990 26812
rect 5024 26778 5058 26812
rect 5092 26778 5126 26812
rect 5160 26778 5194 26812
rect 5228 26778 5262 26812
rect 5296 26778 5330 26812
rect 5364 26778 5398 26812
rect 5432 26778 5466 26812
rect 5500 26778 5534 26812
rect 5568 26778 5602 26812
rect 5636 26778 5670 26812
rect 5704 26778 5738 26812
rect 5772 26778 5806 26812
rect 5840 26778 5874 26812
rect 5908 26778 5942 26812
rect 5976 26778 6010 26812
rect 6044 26778 6078 26812
rect 6112 26778 6146 26812
rect 6180 26778 6214 26812
rect 6248 26778 6282 26812
rect 6316 26778 6350 26812
rect 6384 26778 6418 26812
rect 6452 26778 6486 26812
rect 6520 26778 6554 26812
rect 6588 26778 6622 26812
rect 6656 26778 6690 26812
rect 6724 26778 6758 26812
rect 6792 26778 6826 26812
rect 6860 26778 6894 26812
rect 6928 26778 6962 26812
rect 6996 26778 7030 26812
rect 7064 26778 7098 26812
rect 7132 26778 7166 26812
rect 7200 26778 7234 26812
rect 7268 26778 7302 26812
rect 7336 26778 7370 26812
rect 7404 26778 7438 26812
rect 7472 26778 7506 26812
rect 7540 26778 7574 26812
rect 7608 26778 7642 26812
rect 7676 26778 7710 26812
rect 7744 26778 7778 26812
rect 7812 26778 7846 26812
rect 7880 26778 7914 26812
rect 7948 26778 7982 26812
rect 8016 26778 8050 26812
rect 8084 26778 8118 26812
rect 8152 26778 8186 26812
rect 8220 26778 8254 26812
rect 8288 26778 8322 26812
rect 8356 26778 8390 26812
rect 8424 26778 8458 26812
rect 8492 26778 8526 26812
rect 8560 26778 8594 26812
rect 8628 26778 8662 26812
rect 8696 26778 8730 26812
rect 8764 26778 8798 26812
rect 8832 26778 8866 26812
rect 8900 26778 8934 26812
rect 8968 26778 9002 26812
rect 9036 26778 9070 26812
rect 9104 26778 9138 26812
rect 9172 26778 9206 26812
rect 9240 26778 9274 26812
rect 9308 26778 9342 26812
rect 9376 26778 9410 26812
rect 9444 26778 9478 26812
rect 9512 26778 9546 26812
rect 9580 26778 9614 26812
rect 9648 26778 9682 26812
rect 9716 26778 9750 26812
rect 9784 26778 9818 26812
rect 9852 26778 9886 26812
rect 9920 26778 9954 26812
rect 9988 26778 10022 26812
rect 10056 26778 10090 26812
rect 10124 26778 10158 26812
rect 10192 26778 10226 26812
rect 10260 26778 10294 26812
rect 10328 26778 10362 26812
rect 10396 26778 10430 26812
rect 10464 26778 10498 26812
rect 10532 26778 10566 26812
rect 10600 26778 10634 26812
rect 10668 26778 10702 26812
rect 10736 26778 10770 26812
rect 10804 26778 10838 26812
rect 10872 26778 10906 26812
rect 10940 26778 10974 26812
rect 11008 26778 11042 26812
rect 11076 26778 11110 26812
rect 11144 26778 11178 26812
rect 11212 26778 11246 26812
rect 11280 26778 11314 26812
rect 11348 26778 11382 26812
rect 11416 26778 11450 26812
rect 11484 26778 11518 26812
rect 11552 26778 11586 26812
rect 11620 26778 11654 26812
rect 11688 26778 11722 26812
rect 11756 26778 11790 26812
rect 11824 26778 11858 26812
rect 11892 26778 11926 26812
rect 11960 26778 11994 26812
rect 12028 26778 12062 26812
rect 12096 26778 12130 26812
rect 12164 26778 12198 26812
rect 12232 26778 12266 26812
rect 12300 26778 12334 26812
rect 12368 26778 12402 26812
rect 12436 26778 12470 26812
rect 12504 26778 12538 26812
rect 12572 26778 12606 26812
rect 12640 26778 12674 26812
rect 12708 26778 12742 26812
rect 12776 26778 12810 26812
rect 12844 26778 12878 26812
rect 12912 26778 12946 26812
rect 12980 26778 13014 26812
rect 13048 26778 13082 26812
rect 13116 26778 13150 26812
rect 13184 26778 13218 26812
rect 13252 26778 13286 26812
rect 13320 26778 13354 26812
rect 13388 26778 13422 26812
rect 13456 26778 13490 26812
rect 13524 26778 13558 26812
rect 13592 26778 13626 26812
rect 13660 26778 13694 26812
rect 13728 26778 13762 26812
rect 13796 26778 13830 26812
rect 13864 26778 13898 26812
rect 13932 26778 13966 26812
rect 14000 26778 14034 26812
rect 14068 26778 14102 26812
rect 14136 26778 14170 26812
rect 14204 26778 14238 26812
rect 14272 26778 14306 26812
rect 14340 26778 14374 26812
rect 14408 26778 14442 26812
rect 14476 26778 14510 26812
rect 14544 26778 14578 26812
rect 14612 26778 14646 26812
rect 14680 26778 14714 26812
rect 14748 26778 14782 26812
rect 14816 26778 14850 26812
rect 14884 26778 14918 26812
rect 83 26723 117 26757
rect 152 26723 186 26757
rect 221 26723 255 26757
rect 290 26723 324 26757
rect 359 26723 393 26757
rect 428 26723 462 26757
rect 497 26723 531 26757
rect 566 26723 600 26757
rect 635 26723 669 26757
rect 704 26723 738 26757
rect 773 26723 807 26757
rect 842 26723 876 26757
rect 911 26723 945 26757
rect 980 26723 1014 26757
rect 1049 26723 1083 26757
rect 1118 26723 1152 26757
rect 1187 26723 1221 26757
rect 1256 26723 1290 26757
rect 1325 26723 1359 26757
rect 1394 26723 1428 26757
rect 1463 26723 1497 26757
rect 1532 26723 1566 26757
rect 1601 26723 1635 26757
rect 1670 26723 1704 26757
rect 1739 26723 1773 26757
rect 1808 26723 1842 26757
rect 1877 26723 1911 26757
rect 1946 26723 1980 26757
rect 2014 26723 2048 26757
rect 2082 26723 2116 26757
rect 2150 26723 2184 26757
rect 2218 26723 2252 26757
rect 2286 26723 2320 26757
rect 2354 26723 2388 26757
rect 2422 26723 2456 26757
rect 2490 26723 2524 26757
rect 2558 26723 2592 26757
rect 2626 26723 2660 26757
rect 2694 26723 2728 26757
rect 2762 26723 2796 26757
rect 2848 26708 2882 26742
rect 2916 26708 2950 26742
rect 2984 26708 3018 26742
rect 3052 26708 3086 26742
rect 3120 26708 3154 26742
rect 3188 26708 3222 26742
rect 3256 26708 3290 26742
rect 3324 26708 3358 26742
rect 3392 26708 3426 26742
rect 3460 26708 3494 26742
rect 3528 26708 3562 26742
rect 3596 26708 3630 26742
rect 3664 26708 3698 26742
rect 3732 26708 3766 26742
rect 3800 26708 3834 26742
rect 3868 26708 3902 26742
rect 3936 26708 3970 26742
rect 4004 26708 4038 26742
rect 4072 26708 4106 26742
rect 4140 26708 4174 26742
rect 4208 26708 4242 26742
rect 4276 26708 4310 26742
rect 4344 26708 4378 26742
rect 4412 26708 4446 26742
rect 4480 26708 4514 26742
rect 4548 26708 4582 26742
rect 4616 26708 4650 26742
rect 4684 26708 4718 26742
rect 4752 26708 4786 26742
rect 4820 26708 4854 26742
rect 4888 26708 4922 26742
rect 4956 26708 4990 26742
rect 5024 26708 5058 26742
rect 5092 26708 5126 26742
rect 5160 26708 5194 26742
rect 5228 26708 5262 26742
rect 5296 26708 5330 26742
rect 5364 26708 5398 26742
rect 5432 26708 5466 26742
rect 5500 26708 5534 26742
rect 5568 26708 5602 26742
rect 5636 26708 5670 26742
rect 5704 26708 5738 26742
rect 5772 26708 5806 26742
rect 5840 26708 5874 26742
rect 5908 26708 5942 26742
rect 5976 26708 6010 26742
rect 6044 26708 6078 26742
rect 6112 26708 6146 26742
rect 6180 26708 6214 26742
rect 6248 26708 6282 26742
rect 6316 26708 6350 26742
rect 6384 26708 6418 26742
rect 6452 26708 6486 26742
rect 6520 26708 6554 26742
rect 6588 26708 6622 26742
rect 6656 26708 6690 26742
rect 6724 26708 6758 26742
rect 6792 26708 6826 26742
rect 6860 26708 6894 26742
rect 6928 26708 6962 26742
rect 6996 26708 7030 26742
rect 7064 26708 7098 26742
rect 7132 26708 7166 26742
rect 7200 26708 7234 26742
rect 7268 26708 7302 26742
rect 7336 26708 7370 26742
rect 7404 26708 7438 26742
rect 7472 26708 7506 26742
rect 7540 26708 7574 26742
rect 7608 26708 7642 26742
rect 7676 26708 7710 26742
rect 7744 26708 7778 26742
rect 7812 26708 7846 26742
rect 7880 26708 7914 26742
rect 7948 26708 7982 26742
rect 8016 26708 8050 26742
rect 8084 26708 8118 26742
rect 8152 26708 8186 26742
rect 8220 26708 8254 26742
rect 8288 26708 8322 26742
rect 8356 26708 8390 26742
rect 8424 26708 8458 26742
rect 8492 26708 8526 26742
rect 8560 26708 8594 26742
rect 8628 26708 8662 26742
rect 8696 26708 8730 26742
rect 8764 26708 8798 26742
rect 8832 26708 8866 26742
rect 8900 26708 8934 26742
rect 8968 26708 9002 26742
rect 9036 26708 9070 26742
rect 9104 26708 9138 26742
rect 9172 26708 9206 26742
rect 9240 26708 9274 26742
rect 9308 26708 9342 26742
rect 9376 26708 9410 26742
rect 9444 26708 9478 26742
rect 9512 26708 9546 26742
rect 9580 26708 9614 26742
rect 9648 26708 9682 26742
rect 9716 26708 9750 26742
rect 9784 26708 9818 26742
rect 9852 26708 9886 26742
rect 9920 26708 9954 26742
rect 9988 26708 10022 26742
rect 10056 26708 10090 26742
rect 10124 26708 10158 26742
rect 10192 26708 10226 26742
rect 10260 26708 10294 26742
rect 10328 26708 10362 26742
rect 10396 26708 10430 26742
rect 10464 26708 10498 26742
rect 10532 26708 10566 26742
rect 10600 26708 10634 26742
rect 10668 26708 10702 26742
rect 10736 26708 10770 26742
rect 10804 26708 10838 26742
rect 10872 26708 10906 26742
rect 10940 26708 10974 26742
rect 11008 26708 11042 26742
rect 11076 26708 11110 26742
rect 11144 26708 11178 26742
rect 11212 26708 11246 26742
rect 11280 26708 11314 26742
rect 11348 26708 11382 26742
rect 11416 26708 11450 26742
rect 11484 26708 11518 26742
rect 11552 26708 11586 26742
rect 11620 26708 11654 26742
rect 11688 26708 11722 26742
rect 11756 26708 11790 26742
rect 11824 26708 11858 26742
rect 11892 26708 11926 26742
rect 11960 26708 11994 26742
rect 12028 26708 12062 26742
rect 12096 26708 12130 26742
rect 12164 26708 12198 26742
rect 12232 26708 12266 26742
rect 12300 26708 12334 26742
rect 12368 26708 12402 26742
rect 12436 26708 12470 26742
rect 12504 26708 12538 26742
rect 12572 26708 12606 26742
rect 12640 26708 12674 26742
rect 12708 26708 12742 26742
rect 12776 26708 12810 26742
rect 12844 26708 12878 26742
rect 12912 26708 12946 26742
rect 12980 26708 13014 26742
rect 13048 26708 13082 26742
rect 13116 26708 13150 26742
rect 13184 26708 13218 26742
rect 13252 26708 13286 26742
rect 13320 26708 13354 26742
rect 13388 26708 13422 26742
rect 13456 26708 13490 26742
rect 13524 26708 13558 26742
rect 13592 26708 13626 26742
rect 13660 26708 13694 26742
rect 13728 26708 13762 26742
rect 13796 26708 13830 26742
rect 13864 26708 13898 26742
rect 13932 26708 13966 26742
rect 14000 26708 14034 26742
rect 14068 26708 14102 26742
rect 14136 26708 14170 26742
rect 14204 26708 14238 26742
rect 14272 26708 14306 26742
rect 14340 26708 14374 26742
rect 14408 26708 14442 26742
rect 14476 26708 14510 26742
rect 14544 26708 14578 26742
rect 14612 26708 14646 26742
rect 14680 26708 14714 26742
rect 14748 26708 14782 26742
rect 14816 26708 14850 26742
rect 14884 26708 14918 26742
rect 83 26649 117 26683
rect 152 26649 186 26683
rect 221 26649 255 26683
rect 290 26649 324 26683
rect 359 26649 393 26683
rect 428 26649 462 26683
rect 497 26649 531 26683
rect 566 26649 600 26683
rect 635 26649 669 26683
rect 704 26649 738 26683
rect 773 26649 807 26683
rect 842 26649 876 26683
rect 911 26649 945 26683
rect 980 26649 1014 26683
rect 1049 26649 1083 26683
rect 1118 26649 1152 26683
rect 1187 26649 1221 26683
rect 1256 26649 1290 26683
rect 1325 26649 1359 26683
rect 1394 26649 1428 26683
rect 1463 26649 1497 26683
rect 1532 26649 1566 26683
rect 1601 26649 1635 26683
rect 1670 26649 1704 26683
rect 1739 26649 1773 26683
rect 1808 26649 1842 26683
rect 1877 26649 1911 26683
rect 1946 26649 1980 26683
rect 2014 26649 2048 26683
rect 2082 26649 2116 26683
rect 2150 26649 2184 26683
rect 2218 26649 2252 26683
rect 2286 26649 2320 26683
rect 2354 26649 2388 26683
rect 2422 26649 2456 26683
rect 2490 26649 2524 26683
rect 2558 26649 2592 26683
rect 2626 26649 2660 26683
rect 2694 26649 2728 26683
rect 2762 26649 2796 26683
rect 2848 26638 2882 26672
rect 2916 26638 2950 26672
rect 2984 26638 3018 26672
rect 3052 26638 3086 26672
rect 3120 26638 3154 26672
rect 3188 26638 3222 26672
rect 3256 26638 3290 26672
rect 3324 26638 3358 26672
rect 3392 26638 3426 26672
rect 3460 26638 3494 26672
rect 3528 26638 3562 26672
rect 3596 26638 3630 26672
rect 3664 26638 3698 26672
rect 3732 26638 3766 26672
rect 3800 26638 3834 26672
rect 3868 26638 3902 26672
rect 3936 26638 3970 26672
rect 4004 26638 4038 26672
rect 4072 26638 4106 26672
rect 4140 26638 4174 26672
rect 4208 26638 4242 26672
rect 4276 26638 4310 26672
rect 4344 26638 4378 26672
rect 4412 26638 4446 26672
rect 4480 26638 4514 26672
rect 4548 26638 4582 26672
rect 4616 26638 4650 26672
rect 4684 26638 4718 26672
rect 4752 26638 4786 26672
rect 4820 26638 4854 26672
rect 4888 26638 4922 26672
rect 4956 26638 4990 26672
rect 5024 26638 5058 26672
rect 5092 26638 5126 26672
rect 5160 26638 5194 26672
rect 5228 26638 5262 26672
rect 5296 26638 5330 26672
rect 5364 26638 5398 26672
rect 5432 26638 5466 26672
rect 5500 26638 5534 26672
rect 5568 26638 5602 26672
rect 5636 26638 5670 26672
rect 5704 26638 5738 26672
rect 5772 26638 5806 26672
rect 5840 26638 5874 26672
rect 5908 26638 5942 26672
rect 5976 26638 6010 26672
rect 6044 26638 6078 26672
rect 6112 26638 6146 26672
rect 6180 26638 6214 26672
rect 6248 26638 6282 26672
rect 6316 26638 6350 26672
rect 6384 26638 6418 26672
rect 6452 26638 6486 26672
rect 6520 26638 6554 26672
rect 6588 26638 6622 26672
rect 6656 26638 6690 26672
rect 6724 26638 6758 26672
rect 6792 26638 6826 26672
rect 6860 26638 6894 26672
rect 6928 26638 6962 26672
rect 6996 26638 7030 26672
rect 7064 26638 7098 26672
rect 7132 26638 7166 26672
rect 7200 26638 7234 26672
rect 7268 26638 7302 26672
rect 7336 26638 7370 26672
rect 7404 26638 7438 26672
rect 7472 26638 7506 26672
rect 7540 26638 7574 26672
rect 7608 26638 7642 26672
rect 7676 26638 7710 26672
rect 7744 26638 7778 26672
rect 7812 26638 7846 26672
rect 7880 26638 7914 26672
rect 7948 26638 7982 26672
rect 8016 26638 8050 26672
rect 8084 26638 8118 26672
rect 8152 26638 8186 26672
rect 8220 26638 8254 26672
rect 8288 26638 8322 26672
rect 8356 26638 8390 26672
rect 8424 26638 8458 26672
rect 8492 26638 8526 26672
rect 8560 26638 8594 26672
rect 8628 26638 8662 26672
rect 8696 26638 8730 26672
rect 8764 26638 8798 26672
rect 8832 26638 8866 26672
rect 8900 26638 8934 26672
rect 8968 26638 9002 26672
rect 9036 26638 9070 26672
rect 9104 26638 9138 26672
rect 9172 26638 9206 26672
rect 9240 26638 9274 26672
rect 9308 26638 9342 26672
rect 9376 26638 9410 26672
rect 9444 26638 9478 26672
rect 9512 26638 9546 26672
rect 9580 26638 9614 26672
rect 9648 26638 9682 26672
rect 9716 26638 9750 26672
rect 9784 26638 9818 26672
rect 9852 26638 9886 26672
rect 9920 26638 9954 26672
rect 9988 26638 10022 26672
rect 10056 26638 10090 26672
rect 10124 26638 10158 26672
rect 10192 26638 10226 26672
rect 10260 26638 10294 26672
rect 10328 26638 10362 26672
rect 10396 26638 10430 26672
rect 10464 26638 10498 26672
rect 10532 26638 10566 26672
rect 10600 26638 10634 26672
rect 10668 26638 10702 26672
rect 10736 26638 10770 26672
rect 10804 26638 10838 26672
rect 10872 26638 10906 26672
rect 10940 26638 10974 26672
rect 11008 26638 11042 26672
rect 11076 26638 11110 26672
rect 11144 26638 11178 26672
rect 11212 26638 11246 26672
rect 11280 26638 11314 26672
rect 11348 26638 11382 26672
rect 11416 26638 11450 26672
rect 11484 26638 11518 26672
rect 11552 26638 11586 26672
rect 11620 26638 11654 26672
rect 11688 26638 11722 26672
rect 11756 26638 11790 26672
rect 11824 26638 11858 26672
rect 11892 26638 11926 26672
rect 11960 26638 11994 26672
rect 12028 26638 12062 26672
rect 12096 26638 12130 26672
rect 12164 26638 12198 26672
rect 12232 26638 12266 26672
rect 12300 26638 12334 26672
rect 12368 26638 12402 26672
rect 12436 26638 12470 26672
rect 12504 26638 12538 26672
rect 12572 26638 12606 26672
rect 12640 26638 12674 26672
rect 12708 26638 12742 26672
rect 12776 26638 12810 26672
rect 12844 26638 12878 26672
rect 12912 26638 12946 26672
rect 12980 26638 13014 26672
rect 13048 26638 13082 26672
rect 13116 26638 13150 26672
rect 13184 26638 13218 26672
rect 13252 26638 13286 26672
rect 13320 26638 13354 26672
rect 13388 26638 13422 26672
rect 13456 26638 13490 26672
rect 13524 26638 13558 26672
rect 13592 26638 13626 26672
rect 13660 26638 13694 26672
rect 13728 26638 13762 26672
rect 13796 26638 13830 26672
rect 13864 26638 13898 26672
rect 13932 26638 13966 26672
rect 14000 26638 14034 26672
rect 14068 26638 14102 26672
rect 14136 26638 14170 26672
rect 14204 26638 14238 26672
rect 14272 26638 14306 26672
rect 14340 26638 14374 26672
rect 14408 26638 14442 26672
rect 14476 26638 14510 26672
rect 14544 26638 14578 26672
rect 14612 26638 14646 26672
rect 14680 26638 14714 26672
rect 14748 26638 14782 26672
rect 14816 26638 14850 26672
rect 14884 26638 14918 26672
rect 83 26575 117 26609
rect 152 26575 186 26609
rect 221 26575 255 26609
rect 290 26575 324 26609
rect 359 26575 393 26609
rect 428 26575 462 26609
rect 497 26575 531 26609
rect 566 26575 600 26609
rect 635 26575 669 26609
rect 704 26575 738 26609
rect 773 26575 807 26609
rect 842 26575 876 26609
rect 911 26575 945 26609
rect 980 26575 1014 26609
rect 1049 26575 1083 26609
rect 1118 26575 1152 26609
rect 1187 26575 1221 26609
rect 1256 26575 1290 26609
rect 1325 26575 1359 26609
rect 1394 26575 1428 26609
rect 1463 26575 1497 26609
rect 1532 26575 1566 26609
rect 1601 26575 1635 26609
rect 1670 26575 1704 26609
rect 1739 26575 1773 26609
rect 1808 26575 1842 26609
rect 1877 26575 1911 26609
rect 1946 26575 1980 26609
rect 2014 26575 2048 26609
rect 2082 26575 2116 26609
rect 2150 26575 2184 26609
rect 2218 26575 2252 26609
rect 2286 26575 2320 26609
rect 2354 26575 2388 26609
rect 2422 26575 2456 26609
rect 2490 26575 2524 26609
rect 2558 26575 2592 26609
rect 2626 26575 2660 26609
rect 2694 26575 2728 26609
rect 2762 26575 2796 26609
rect 2848 26568 2882 26602
rect 2916 26568 2950 26602
rect 2984 26568 3018 26602
rect 3052 26568 3086 26602
rect 3120 26568 3154 26602
rect 3188 26568 3222 26602
rect 3256 26568 3290 26602
rect 3324 26568 3358 26602
rect 3392 26568 3426 26602
rect 3460 26568 3494 26602
rect 3528 26568 3562 26602
rect 3596 26568 3630 26602
rect 3664 26568 3698 26602
rect 3732 26568 3766 26602
rect 3800 26568 3834 26602
rect 3868 26568 3902 26602
rect 3936 26568 3970 26602
rect 4004 26568 4038 26602
rect 4072 26568 4106 26602
rect 4140 26568 4174 26602
rect 4208 26568 4242 26602
rect 4276 26568 4310 26602
rect 4344 26568 4378 26602
rect 4412 26568 4446 26602
rect 4480 26568 4514 26602
rect 4548 26568 4582 26602
rect 4616 26568 4650 26602
rect 4684 26568 4718 26602
rect 4752 26568 4786 26602
rect 4820 26568 4854 26602
rect 4888 26568 4922 26602
rect 4956 26568 4990 26602
rect 5024 26568 5058 26602
rect 5092 26568 5126 26602
rect 5160 26568 5194 26602
rect 5228 26568 5262 26602
rect 5296 26568 5330 26602
rect 5364 26568 5398 26602
rect 5432 26568 5466 26602
rect 5500 26568 5534 26602
rect 5568 26568 5602 26602
rect 5636 26568 5670 26602
rect 5704 26568 5738 26602
rect 5772 26568 5806 26602
rect 5840 26568 5874 26602
rect 5908 26568 5942 26602
rect 5976 26568 6010 26602
rect 6044 26568 6078 26602
rect 6112 26568 6146 26602
rect 6180 26568 6214 26602
rect 6248 26568 6282 26602
rect 6316 26568 6350 26602
rect 6384 26568 6418 26602
rect 6452 26568 6486 26602
rect 6520 26568 6554 26602
rect 6588 26568 6622 26602
rect 6656 26568 6690 26602
rect 6724 26568 6758 26602
rect 6792 26568 6826 26602
rect 6860 26568 6894 26602
rect 6928 26568 6962 26602
rect 6996 26568 7030 26602
rect 7064 26568 7098 26602
rect 7132 26568 7166 26602
rect 7200 26568 7234 26602
rect 7268 26568 7302 26602
rect 7336 26568 7370 26602
rect 7404 26568 7438 26602
rect 7472 26568 7506 26602
rect 7540 26568 7574 26602
rect 7608 26568 7642 26602
rect 7676 26568 7710 26602
rect 7744 26568 7778 26602
rect 7812 26568 7846 26602
rect 7880 26568 7914 26602
rect 7948 26568 7982 26602
rect 8016 26568 8050 26602
rect 8084 26568 8118 26602
rect 8152 26568 8186 26602
rect 8220 26568 8254 26602
rect 8288 26568 8322 26602
rect 8356 26568 8390 26602
rect 8424 26568 8458 26602
rect 8492 26568 8526 26602
rect 8560 26568 8594 26602
rect 8628 26568 8662 26602
rect 8696 26568 8730 26602
rect 8764 26568 8798 26602
rect 8832 26568 8866 26602
rect 8900 26568 8934 26602
rect 8968 26568 9002 26602
rect 9036 26568 9070 26602
rect 9104 26568 9138 26602
rect 9172 26568 9206 26602
rect 9240 26568 9274 26602
rect 9308 26568 9342 26602
rect 9376 26568 9410 26602
rect 9444 26568 9478 26602
rect 9512 26568 9546 26602
rect 9580 26568 9614 26602
rect 9648 26568 9682 26602
rect 9716 26568 9750 26602
rect 9784 26568 9818 26602
rect 9852 26568 9886 26602
rect 9920 26568 9954 26602
rect 9988 26568 10022 26602
rect 10056 26568 10090 26602
rect 10124 26568 10158 26602
rect 10192 26568 10226 26602
rect 10260 26568 10294 26602
rect 10328 26568 10362 26602
rect 10396 26568 10430 26602
rect 10464 26568 10498 26602
rect 10532 26568 10566 26602
rect 10600 26568 10634 26602
rect 10668 26568 10702 26602
rect 10736 26568 10770 26602
rect 10804 26568 10838 26602
rect 10872 26568 10906 26602
rect 10940 26568 10974 26602
rect 11008 26568 11042 26602
rect 11076 26568 11110 26602
rect 11144 26568 11178 26602
rect 11212 26568 11246 26602
rect 11280 26568 11314 26602
rect 11348 26568 11382 26602
rect 11416 26568 11450 26602
rect 11484 26568 11518 26602
rect 11552 26568 11586 26602
rect 11620 26568 11654 26602
rect 11688 26568 11722 26602
rect 11756 26568 11790 26602
rect 11824 26568 11858 26602
rect 11892 26568 11926 26602
rect 11960 26568 11994 26602
rect 12028 26568 12062 26602
rect 12096 26568 12130 26602
rect 12164 26568 12198 26602
rect 12232 26568 12266 26602
rect 12300 26568 12334 26602
rect 12368 26568 12402 26602
rect 12436 26568 12470 26602
rect 12504 26568 12538 26602
rect 12572 26568 12606 26602
rect 12640 26568 12674 26602
rect 12708 26568 12742 26602
rect 12776 26568 12810 26602
rect 12844 26568 12878 26602
rect 12912 26568 12946 26602
rect 12980 26568 13014 26602
rect 13048 26568 13082 26602
rect 13116 26568 13150 26602
rect 13184 26568 13218 26602
rect 13252 26568 13286 26602
rect 13320 26568 13354 26602
rect 13388 26568 13422 26602
rect 13456 26568 13490 26602
rect 13524 26568 13558 26602
rect 13592 26568 13626 26602
rect 13660 26568 13694 26602
rect 13728 26568 13762 26602
rect 13796 26568 13830 26602
rect 13864 26568 13898 26602
rect 13932 26568 13966 26602
rect 14000 26568 14034 26602
rect 14068 26568 14102 26602
rect 14136 26568 14170 26602
rect 14204 26568 14238 26602
rect 14272 26568 14306 26602
rect 14340 26568 14374 26602
rect 14408 26568 14442 26602
rect 14476 26568 14510 26602
rect 14544 26568 14578 26602
rect 14612 26568 14646 26602
rect 14680 26568 14714 26602
rect 14748 26568 14782 26602
rect 14816 26568 14850 26602
rect 14884 26568 14918 26602
rect 83 26501 117 26535
rect 152 26501 186 26535
rect 221 26501 255 26535
rect 290 26501 324 26535
rect 359 26501 393 26535
rect 428 26501 462 26535
rect 497 26501 531 26535
rect 566 26501 600 26535
rect 635 26501 669 26535
rect 704 26501 738 26535
rect 773 26501 807 26535
rect 842 26501 876 26535
rect 911 26501 945 26535
rect 980 26501 1014 26535
rect 1049 26501 1083 26535
rect 1118 26501 1152 26535
rect 1187 26501 1221 26535
rect 1256 26501 1290 26535
rect 1325 26501 1359 26535
rect 1394 26501 1428 26535
rect 1463 26501 1497 26535
rect 1532 26501 1566 26535
rect 1601 26501 1635 26535
rect 1670 26501 1704 26535
rect 1739 26501 1773 26535
rect 1808 26501 1842 26535
rect 1877 26501 1911 26535
rect 1946 26501 1980 26535
rect 2014 26501 2048 26535
rect 2082 26501 2116 26535
rect 2150 26501 2184 26535
rect 2218 26501 2252 26535
rect 2286 26501 2320 26535
rect 2354 26501 2388 26535
rect 2422 26501 2456 26535
rect 2490 26501 2524 26535
rect 2558 26501 2592 26535
rect 2626 26501 2660 26535
rect 2694 26501 2728 26535
rect 2762 26501 2796 26535
rect 2848 26498 2882 26532
rect 2916 26498 2950 26532
rect 2984 26498 3018 26532
rect 3052 26498 3086 26532
rect 3120 26498 3154 26532
rect 3188 26498 3222 26532
rect 3256 26498 3290 26532
rect 3324 26498 3358 26532
rect 3392 26498 3426 26532
rect 3460 26498 3494 26532
rect 3528 26498 3562 26532
rect 3596 26498 3630 26532
rect 3664 26498 3698 26532
rect 3732 26498 3766 26532
rect 3800 26498 3834 26532
rect 3868 26498 3902 26532
rect 3936 26498 3970 26532
rect 4004 26498 4038 26532
rect 4072 26498 4106 26532
rect 4140 26498 4174 26532
rect 4208 26498 4242 26532
rect 4276 26498 4310 26532
rect 4344 26498 4378 26532
rect 4412 26498 4446 26532
rect 4480 26498 4514 26532
rect 4548 26498 4582 26532
rect 4616 26498 4650 26532
rect 4684 26498 4718 26532
rect 4752 26498 4786 26532
rect 4820 26498 4854 26532
rect 4888 26498 4922 26532
rect 4956 26498 4990 26532
rect 5024 26498 5058 26532
rect 5092 26498 5126 26532
rect 5160 26498 5194 26532
rect 5228 26498 5262 26532
rect 5296 26498 5330 26532
rect 5364 26498 5398 26532
rect 5432 26498 5466 26532
rect 5500 26498 5534 26532
rect 5568 26498 5602 26532
rect 5636 26498 5670 26532
rect 5704 26498 5738 26532
rect 5772 26498 5806 26532
rect 5840 26498 5874 26532
rect 5908 26498 5942 26532
rect 5976 26498 6010 26532
rect 6044 26498 6078 26532
rect 6112 26498 6146 26532
rect 6180 26498 6214 26532
rect 6248 26498 6282 26532
rect 6316 26498 6350 26532
rect 6384 26498 6418 26532
rect 6452 26498 6486 26532
rect 6520 26498 6554 26532
rect 6588 26498 6622 26532
rect 6656 26498 6690 26532
rect 6724 26498 6758 26532
rect 6792 26498 6826 26532
rect 6860 26498 6894 26532
rect 6928 26498 6962 26532
rect 6996 26498 7030 26532
rect 7064 26498 7098 26532
rect 7132 26498 7166 26532
rect 7200 26498 7234 26532
rect 7268 26498 7302 26532
rect 7336 26498 7370 26532
rect 7404 26498 7438 26532
rect 7472 26498 7506 26532
rect 7540 26498 7574 26532
rect 7608 26498 7642 26532
rect 7676 26498 7710 26532
rect 7744 26498 7778 26532
rect 7812 26498 7846 26532
rect 7880 26498 7914 26532
rect 7948 26498 7982 26532
rect 8016 26498 8050 26532
rect 8084 26498 8118 26532
rect 8152 26498 8186 26532
rect 8220 26498 8254 26532
rect 8288 26498 8322 26532
rect 8356 26498 8390 26532
rect 8424 26498 8458 26532
rect 8492 26498 8526 26532
rect 8560 26498 8594 26532
rect 8628 26498 8662 26532
rect 8696 26498 8730 26532
rect 8764 26498 8798 26532
rect 8832 26498 8866 26532
rect 8900 26498 8934 26532
rect 8968 26498 9002 26532
rect 9036 26498 9070 26532
rect 9104 26498 9138 26532
rect 9172 26498 9206 26532
rect 9240 26498 9274 26532
rect 9308 26498 9342 26532
rect 9376 26498 9410 26532
rect 9444 26498 9478 26532
rect 9512 26498 9546 26532
rect 9580 26498 9614 26532
rect 9648 26498 9682 26532
rect 9716 26498 9750 26532
rect 9784 26498 9818 26532
rect 9852 26498 9886 26532
rect 9920 26498 9954 26532
rect 9988 26498 10022 26532
rect 10056 26498 10090 26532
rect 10124 26498 10158 26532
rect 10192 26498 10226 26532
rect 10260 26498 10294 26532
rect 10328 26498 10362 26532
rect 10396 26498 10430 26532
rect 10464 26498 10498 26532
rect 10532 26498 10566 26532
rect 10600 26498 10634 26532
rect 10668 26498 10702 26532
rect 10736 26498 10770 26532
rect 10804 26498 10838 26532
rect 10872 26498 10906 26532
rect 10940 26498 10974 26532
rect 11008 26498 11042 26532
rect 11076 26498 11110 26532
rect 11144 26498 11178 26532
rect 11212 26498 11246 26532
rect 11280 26498 11314 26532
rect 11348 26498 11382 26532
rect 11416 26498 11450 26532
rect 11484 26498 11518 26532
rect 11552 26498 11586 26532
rect 11620 26498 11654 26532
rect 11688 26498 11722 26532
rect 11756 26498 11790 26532
rect 11824 26498 11858 26532
rect 11892 26498 11926 26532
rect 11960 26498 11994 26532
rect 12028 26498 12062 26532
rect 12096 26498 12130 26532
rect 12164 26498 12198 26532
rect 12232 26498 12266 26532
rect 12300 26498 12334 26532
rect 12368 26498 12402 26532
rect 12436 26498 12470 26532
rect 12504 26498 12538 26532
rect 12572 26498 12606 26532
rect 12640 26498 12674 26532
rect 12708 26498 12742 26532
rect 12776 26498 12810 26532
rect 12844 26498 12878 26532
rect 12912 26498 12946 26532
rect 12980 26498 13014 26532
rect 13048 26498 13082 26532
rect 13116 26498 13150 26532
rect 13184 26498 13218 26532
rect 13252 26498 13286 26532
rect 13320 26498 13354 26532
rect 13388 26498 13422 26532
rect 13456 26498 13490 26532
rect 13524 26498 13558 26532
rect 13592 26498 13626 26532
rect 13660 26498 13694 26532
rect 13728 26498 13762 26532
rect 13796 26498 13830 26532
rect 13864 26498 13898 26532
rect 13932 26498 13966 26532
rect 14000 26498 14034 26532
rect 14068 26498 14102 26532
rect 14136 26498 14170 26532
rect 14204 26498 14238 26532
rect 14272 26498 14306 26532
rect 14340 26498 14374 26532
rect 14408 26498 14442 26532
rect 14476 26498 14510 26532
rect 14544 26498 14578 26532
rect 14612 26498 14646 26532
rect 14680 26498 14714 26532
rect 14748 26498 14782 26532
rect 14816 26498 14850 26532
rect 14884 26498 14918 26532
rect 83 26427 117 26461
rect 152 26427 186 26461
rect 221 26427 255 26461
rect 290 26427 324 26461
rect 359 26427 393 26461
rect 428 26427 462 26461
rect 497 26427 531 26461
rect 566 26427 600 26461
rect 635 26427 669 26461
rect 704 26427 738 26461
rect 773 26427 807 26461
rect 842 26427 876 26461
rect 911 26427 945 26461
rect 980 26427 1014 26461
rect 1049 26427 1083 26461
rect 1118 26427 1152 26461
rect 1187 26427 1221 26461
rect 1256 26427 1290 26461
rect 1325 26427 1359 26461
rect 1394 26427 1428 26461
rect 1463 26427 1497 26461
rect 1532 26427 1566 26461
rect 1601 26427 1635 26461
rect 1670 26427 1704 26461
rect 1739 26427 1773 26461
rect 1808 26427 1842 26461
rect 1877 26427 1911 26461
rect 1946 26427 1980 26461
rect 2014 26427 2048 26461
rect 2082 26427 2116 26461
rect 2150 26427 2184 26461
rect 2218 26427 2252 26461
rect 2286 26427 2320 26461
rect 2354 26427 2388 26461
rect 2422 26427 2456 26461
rect 2490 26427 2524 26461
rect 2558 26427 2592 26461
rect 2626 26427 2660 26461
rect 2694 26427 2728 26461
rect 2762 26427 2796 26461
rect 2848 26428 2882 26462
rect 2916 26428 2950 26462
rect 2984 26428 3018 26462
rect 3052 26428 3086 26462
rect 3120 26428 3154 26462
rect 3188 26428 3222 26462
rect 3256 26428 3290 26462
rect 3324 26428 3358 26462
rect 3392 26428 3426 26462
rect 3460 26428 3494 26462
rect 3528 26428 3562 26462
rect 3596 26428 3630 26462
rect 3664 26428 3698 26462
rect 3732 26428 3766 26462
rect 3800 26428 3834 26462
rect 3868 26428 3902 26462
rect 3936 26428 3970 26462
rect 4004 26428 4038 26462
rect 4072 26428 4106 26462
rect 4140 26428 4174 26462
rect 4208 26428 4242 26462
rect 4276 26428 4310 26462
rect 4344 26428 4378 26462
rect 4412 26428 4446 26462
rect 4480 26428 4514 26462
rect 4548 26428 4582 26462
rect 4616 26428 4650 26462
rect 4684 26428 4718 26462
rect 4752 26428 4786 26462
rect 4820 26428 4854 26462
rect 4888 26428 4922 26462
rect 4956 26428 4990 26462
rect 5024 26428 5058 26462
rect 5092 26428 5126 26462
rect 5160 26428 5194 26462
rect 5228 26428 5262 26462
rect 5296 26428 5330 26462
rect 5364 26428 5398 26462
rect 5432 26428 5466 26462
rect 5500 26428 5534 26462
rect 5568 26428 5602 26462
rect 5636 26428 5670 26462
rect 5704 26428 5738 26462
rect 5772 26428 5806 26462
rect 5840 26428 5874 26462
rect 5908 26428 5942 26462
rect 5976 26428 6010 26462
rect 6044 26428 6078 26462
rect 6112 26428 6146 26462
rect 6180 26428 6214 26462
rect 6248 26428 6282 26462
rect 6316 26428 6350 26462
rect 6384 26428 6418 26462
rect 6452 26428 6486 26462
rect 6520 26428 6554 26462
rect 6588 26428 6622 26462
rect 6656 26428 6690 26462
rect 6724 26428 6758 26462
rect 6792 26428 6826 26462
rect 6860 26428 6894 26462
rect 6928 26428 6962 26462
rect 6996 26428 7030 26462
rect 7064 26428 7098 26462
rect 7132 26428 7166 26462
rect 7200 26428 7234 26462
rect 7268 26428 7302 26462
rect 7336 26428 7370 26462
rect 7404 26428 7438 26462
rect 7472 26428 7506 26462
rect 7540 26428 7574 26462
rect 7608 26428 7642 26462
rect 7676 26428 7710 26462
rect 7744 26428 7778 26462
rect 7812 26428 7846 26462
rect 7880 26428 7914 26462
rect 7948 26428 7982 26462
rect 8016 26428 8050 26462
rect 8084 26428 8118 26462
rect 8152 26428 8186 26462
rect 8220 26428 8254 26462
rect 8288 26428 8322 26462
rect 8356 26428 8390 26462
rect 8424 26428 8458 26462
rect 8492 26428 8526 26462
rect 8560 26428 8594 26462
rect 8628 26428 8662 26462
rect 8696 26428 8730 26462
rect 8764 26428 8798 26462
rect 8832 26428 8866 26462
rect 8900 26428 8934 26462
rect 8968 26428 9002 26462
rect 9036 26428 9070 26462
rect 9104 26428 9138 26462
rect 9172 26428 9206 26462
rect 9240 26428 9274 26462
rect 9308 26428 9342 26462
rect 9376 26428 9410 26462
rect 9444 26428 9478 26462
rect 9512 26428 9546 26462
rect 9580 26428 9614 26462
rect 9648 26428 9682 26462
rect 9716 26428 9750 26462
rect 9784 26428 9818 26462
rect 9852 26428 9886 26462
rect 9920 26428 9954 26462
rect 9988 26428 10022 26462
rect 10056 26428 10090 26462
rect 10124 26428 10158 26462
rect 10192 26428 10226 26462
rect 10260 26428 10294 26462
rect 10328 26428 10362 26462
rect 10396 26428 10430 26462
rect 10464 26428 10498 26462
rect 10532 26428 10566 26462
rect 10600 26428 10634 26462
rect 10668 26428 10702 26462
rect 10736 26428 10770 26462
rect 10804 26428 10838 26462
rect 10872 26428 10906 26462
rect 10940 26428 10974 26462
rect 11008 26428 11042 26462
rect 11076 26428 11110 26462
rect 11144 26428 11178 26462
rect 11212 26428 11246 26462
rect 11280 26428 11314 26462
rect 11348 26428 11382 26462
rect 11416 26428 11450 26462
rect 11484 26428 11518 26462
rect 11552 26428 11586 26462
rect 11620 26428 11654 26462
rect 11688 26428 11722 26462
rect 11756 26428 11790 26462
rect 11824 26428 11858 26462
rect 11892 26428 11926 26462
rect 11960 26428 11994 26462
rect 12028 26428 12062 26462
rect 12096 26428 12130 26462
rect 12164 26428 12198 26462
rect 12232 26428 12266 26462
rect 12300 26428 12334 26462
rect 12368 26428 12402 26462
rect 12436 26428 12470 26462
rect 12504 26428 12538 26462
rect 12572 26428 12606 26462
rect 12640 26428 12674 26462
rect 12708 26428 12742 26462
rect 12776 26428 12810 26462
rect 12844 26428 12878 26462
rect 12912 26428 12946 26462
rect 12980 26428 13014 26462
rect 13048 26428 13082 26462
rect 13116 26428 13150 26462
rect 13184 26428 13218 26462
rect 13252 26428 13286 26462
rect 13320 26428 13354 26462
rect 13388 26428 13422 26462
rect 13456 26428 13490 26462
rect 13524 26428 13558 26462
rect 13592 26428 13626 26462
rect 13660 26428 13694 26462
rect 13728 26428 13762 26462
rect 13796 26428 13830 26462
rect 13864 26428 13898 26462
rect 13932 26428 13966 26462
rect 14000 26428 14034 26462
rect 14068 26428 14102 26462
rect 14136 26428 14170 26462
rect 14204 26428 14238 26462
rect 14272 26428 14306 26462
rect 14340 26428 14374 26462
rect 14408 26428 14442 26462
rect 14476 26428 14510 26462
rect 14544 26428 14578 26462
rect 14612 26428 14646 26462
rect 14680 26428 14714 26462
rect 14748 26428 14782 26462
rect 14816 26428 14850 26462
rect 14884 26428 14918 26462
rect 83 26317 117 26351
rect 152 26317 186 26351
rect 221 26317 255 26351
rect 290 26317 324 26351
rect 359 26317 393 26351
rect 428 26317 462 26351
rect 497 26317 531 26351
rect 566 26317 600 26351
rect 635 26317 669 26351
rect 704 26317 738 26351
rect 773 26317 807 26351
rect 842 26317 876 26351
rect 911 26317 945 26351
rect 980 26317 1014 26351
rect 1049 26317 1083 26351
rect 1118 26317 1152 26351
rect 1187 26317 1221 26351
rect 1256 26317 1290 26351
rect 1325 26317 1359 26351
rect 1394 26317 1428 26351
rect 1463 26317 1497 26351
rect 1532 26317 1566 26351
rect 1601 26317 1635 26351
rect 1670 26317 1704 26351
rect 1739 26317 1773 26351
rect 1808 26317 1842 26351
rect 1877 26317 1911 26351
rect 1946 26317 1980 26351
rect 2015 26317 2049 26351
rect 2084 26317 2118 26351
rect 2153 26317 2187 26351
rect 2222 26317 2256 26351
rect 2291 26317 2325 26351
rect 2360 26317 2394 26351
rect 2429 26317 2463 26351
rect 2498 26317 2532 26351
rect 2567 26317 2601 26351
rect 2636 26317 2670 26351
rect 2705 26317 2739 26351
rect 2774 26317 2808 26351
rect 2843 26317 2877 26351
rect 2912 26317 2946 26351
rect 2981 26317 3015 26351
rect 3050 26317 3084 26351
rect 3119 26317 3153 26351
rect 3188 26317 3222 26351
rect 3256 26317 3290 26351
rect 3324 26317 3358 26351
rect 3392 26317 3426 26351
rect 3460 26317 3494 26351
rect 3528 26317 3562 26351
rect 3596 26317 3630 26351
rect 3664 26317 3698 26351
rect 3732 26317 3766 26351
rect 3800 26317 3834 26351
rect 3868 26317 3902 26351
rect 3936 26317 3970 26351
rect 4004 26317 4038 26351
rect 4072 26317 4106 26351
rect 4140 26317 4174 26351
rect 4208 26317 4242 26351
rect 4276 26317 4310 26351
rect 4344 26317 4378 26351
rect 4412 26317 4446 26351
rect 4480 26317 4514 26351
rect 4548 26317 4582 26351
rect 4616 26317 4650 26351
rect 4684 26317 4718 26351
rect 4752 26317 4786 26351
rect 4820 26317 4854 26351
rect 4888 26317 4922 26351
rect 4956 26317 4990 26351
rect 5024 26317 5058 26351
rect 5092 26317 5126 26351
rect 5160 26317 5194 26351
rect 5228 26317 5262 26351
rect 5296 26317 5330 26351
rect 5364 26317 5398 26351
rect 5432 26317 5466 26351
rect 5500 26317 5534 26351
rect 5568 26317 5602 26351
rect 5636 26317 5670 26351
rect 5704 26317 5738 26351
rect 5772 26317 5806 26351
rect 5840 26317 5874 26351
rect 5908 26317 5942 26351
rect 5976 26317 6010 26351
rect 6044 26317 6078 26351
rect 6112 26317 6146 26351
rect 6180 26317 6214 26351
rect 6248 26317 6282 26351
rect 6316 26317 6350 26351
rect 6384 26317 6418 26351
rect 6452 26317 6486 26351
rect 6520 26317 6554 26351
rect 6588 26317 6622 26351
rect 6656 26317 6690 26351
rect 6724 26317 6758 26351
rect 6792 26317 6826 26351
rect 6860 26317 6894 26351
rect 6928 26317 6962 26351
rect 6996 26317 7030 26351
rect 7064 26317 7098 26351
rect 7132 26317 7166 26351
rect 7200 26317 7234 26351
rect 7268 26317 7302 26351
rect 7336 26317 7370 26351
rect 7404 26317 7438 26351
rect 7472 26317 7506 26351
rect 7540 26317 7574 26351
rect 7608 26317 7642 26351
rect 7676 26317 7710 26351
rect 7744 26317 7778 26351
rect 7812 26317 7846 26351
rect 7880 26317 7914 26351
rect 7948 26317 7982 26351
rect 8016 26317 8050 26351
rect 8084 26317 8118 26351
rect 8152 26317 8186 26351
rect 8220 26317 8254 26351
rect 8288 26317 8322 26351
rect 8356 26317 8390 26351
rect 8424 26317 8458 26351
rect 8492 26317 8526 26351
rect 8560 26317 8594 26351
rect 8628 26317 8662 26351
rect 8696 26317 8730 26351
rect 8764 26317 8798 26351
rect 8832 26317 8866 26351
rect 8900 26317 8934 26351
rect 8968 26317 9002 26351
rect 9036 26317 9070 26351
rect 9104 26317 9138 26351
rect 9172 26317 9206 26351
rect 9240 26317 9274 26351
rect 9308 26317 9342 26351
rect 9376 26317 9410 26351
rect 9444 26317 9478 26351
rect 9512 26317 9546 26351
rect 9580 26317 9614 26351
rect 9648 26317 9682 26351
rect 9716 26317 9750 26351
rect 9784 26317 9818 26351
rect 9852 26317 9886 26351
rect 9920 26317 9954 26351
rect 9988 26317 10022 26351
rect 10056 26317 10090 26351
rect 10124 26317 10158 26351
rect 10192 26317 10226 26351
rect 10260 26317 10294 26351
rect 10328 26317 10362 26351
rect 10396 26317 10430 26351
rect 10464 26317 10498 26351
rect 10532 26317 10566 26351
rect 10600 26317 10634 26351
rect 10668 26317 10702 26351
rect 10736 26317 10770 26351
rect 10804 26317 10838 26351
rect 10872 26317 10906 26351
rect 10940 26317 10974 26351
rect 11008 26317 11042 26351
rect 11076 26317 11110 26351
rect 11144 26317 11178 26351
rect 11212 26317 11246 26351
rect 11280 26317 11314 26351
rect 11348 26317 11382 26351
rect 11416 26317 11450 26351
rect 11484 26317 11518 26351
rect 11552 26317 11586 26351
rect 11620 26317 11654 26351
rect 11688 26317 11722 26351
rect 11756 26317 11790 26351
rect 11824 26317 11858 26351
rect 11892 26317 11926 26351
rect 11960 26317 11994 26351
rect 12028 26317 12062 26351
rect 12096 26317 12130 26351
rect 12164 26317 12198 26351
rect 12232 26317 12266 26351
rect 12300 26317 12334 26351
rect 12368 26317 12402 26351
rect 12436 26317 12470 26351
rect 12504 26317 12538 26351
rect 12572 26317 12606 26351
rect 12640 26317 12674 26351
rect 12708 26317 12742 26351
rect 12776 26317 12810 26351
rect 12844 26317 12878 26351
rect 12912 26317 12946 26351
rect 12980 26317 13014 26351
rect 13048 26317 13082 26351
rect 13116 26317 13150 26351
rect 13184 26317 13218 26351
rect 13252 26317 13286 26351
rect 13320 26317 13354 26351
rect 13388 26317 13422 26351
rect 13456 26317 13490 26351
rect 13524 26317 13558 26351
rect 13592 26317 13626 26351
rect 13660 26317 13694 26351
rect 13728 26317 13762 26351
rect 13796 26317 13830 26351
rect 13864 26317 13898 26351
rect 13932 26317 13966 26351
rect 14000 26317 14034 26351
rect 14068 26317 14102 26351
rect 14136 26317 14170 26351
rect 14204 26317 14238 26351
rect 14272 26317 14306 26351
rect 14340 26317 14374 26351
rect 14408 26317 14442 26351
rect 14476 26317 14510 26351
rect 14544 26317 14578 26351
rect 14612 26317 14646 26351
rect 14680 26317 14714 26351
rect 14748 26317 14782 26351
rect 14816 26317 14850 26351
rect 14884 26317 14918 26351
rect 69 26210 103 26244
rect 138 26210 172 26244
rect 207 26210 241 26244
rect 276 26210 310 26244
rect 345 26210 379 26244
rect 414 26210 448 26244
rect 483 26210 517 26244
rect 552 26210 586 26244
rect 621 26210 655 26244
rect 690 26210 724 26244
rect 759 26210 793 26244
rect 828 26210 862 26244
rect 897 26210 931 26244
rect 966 26210 1000 26244
rect 1035 26210 1069 26244
rect 1104 26210 1138 26244
rect 1173 26210 1207 26244
rect 1242 26210 1276 26244
rect 1311 26210 1345 26244
rect 1380 26210 1414 26244
rect 1449 26210 1483 26244
rect 1518 26210 1552 26244
rect 1587 26210 1621 26244
rect 1656 26210 1690 26244
rect 1725 26210 1759 26244
rect 1794 26210 1828 26244
rect 1863 26210 1897 26244
rect 1932 26210 1966 26244
rect 2001 26210 2035 26244
rect 2070 26210 2104 26244
rect 2139 26210 2173 26244
rect 2208 26210 2242 26244
rect 2277 26210 2311 26244
rect 2346 26210 2380 26244
rect 2415 26210 2449 26244
rect 2484 26210 2518 26244
rect 2553 26210 2587 26244
rect 2622 26210 2656 26244
rect 2691 26210 2725 26244
rect 2760 26210 2794 26244
rect 2829 26210 2863 26244
rect 2898 26210 2932 26244
rect 2967 26210 3001 26244
rect 3036 26210 3070 26244
rect 3105 26210 3139 26244
rect 3174 26210 3208 26244
rect 3243 26210 3277 26244
rect 3312 26210 3346 26244
rect 3381 26210 3415 26244
rect 3450 26210 3484 26244
rect 3519 26210 3553 26244
rect 3588 26210 3622 26244
rect 3657 26210 3691 26244
rect 3726 26210 3760 26244
rect 3795 26210 3829 26244
rect 3864 26210 3898 26244
rect 3933 26210 3967 26244
rect 4002 26210 4036 26244
rect 4071 26210 4105 26244
rect 4140 26210 4174 26244
rect 4208 26210 4242 26244
rect 4276 26210 4310 26244
rect 4344 26210 4378 26244
rect 4412 26210 4446 26244
rect 4480 26210 4514 26244
rect 4548 26210 4582 26244
rect 4616 26210 4650 26244
rect 4684 26210 4718 26244
rect 4752 26210 4786 26244
rect 4820 26210 4854 26244
rect 4888 26210 4922 26244
rect 4956 26210 4990 26244
rect 5024 26210 5058 26244
rect 5092 26210 5126 26244
rect 5160 26210 5194 26244
rect 5228 26210 5262 26244
rect 5296 26210 5330 26244
rect 5364 26210 5398 26244
rect 5432 26210 5466 26244
rect 5500 26210 5534 26244
rect 5568 26210 5602 26244
rect 5636 26210 5670 26244
rect 5704 26210 5738 26244
rect 5772 26210 5806 26244
rect 5840 26210 5874 26244
rect 5908 26210 5942 26244
rect 5976 26210 6010 26244
rect 6044 26210 6078 26244
rect 6112 26210 6146 26244
rect 6180 26210 6214 26244
rect 6248 26210 6282 26244
rect 6316 26210 6350 26244
rect 6384 26210 6418 26244
rect 6452 26210 6486 26244
rect 6520 26210 6554 26244
rect 6588 26210 6622 26244
rect 6656 26210 6690 26244
rect 6724 26210 6758 26244
rect 6792 26210 6826 26244
rect 6860 26210 6894 26244
rect 6928 26210 6962 26244
rect 6996 26210 7030 26244
rect 7064 26210 7098 26244
rect 7132 26210 7166 26244
rect 7200 26210 7234 26244
rect 7268 26210 7302 26244
rect 7336 26210 7370 26244
rect 7404 26210 7438 26244
rect 7472 26210 7506 26244
rect 7540 26210 7574 26244
rect 7608 26210 7642 26244
rect 7676 26210 7710 26244
rect 7744 26210 7778 26244
rect 7812 26210 7846 26244
rect 7880 26210 7914 26244
rect 7948 26210 7982 26244
rect 8016 26210 8050 26244
rect 8084 26210 8118 26244
rect 8152 26210 8186 26244
rect 8220 26210 8254 26244
rect 8288 26210 8322 26244
rect 8356 26210 8390 26244
rect 8424 26210 8458 26244
rect 8492 26210 8526 26244
rect 8560 26210 8594 26244
rect 8628 26210 8662 26244
rect 8696 26210 8730 26244
rect 8764 26210 8798 26244
rect 8832 26210 8866 26244
rect 8900 26210 8934 26244
rect 8968 26210 9002 26244
rect 9036 26210 9070 26244
rect 9104 26210 9138 26244
rect 9172 26210 9206 26244
rect 9240 26210 9274 26244
rect 9308 26210 9342 26244
rect 9376 26210 9410 26244
rect 9444 26210 9478 26244
rect 9512 26210 9546 26244
rect 9580 26210 9614 26244
rect 9648 26210 9682 26244
rect 9716 26210 9750 26244
rect 9784 26210 9818 26244
rect 9852 26210 9886 26244
rect 9920 26210 9954 26244
rect 9988 26210 10022 26244
rect 10056 26210 10090 26244
rect 10124 26210 10158 26244
rect 10192 26210 10226 26244
rect 10260 26210 10294 26244
rect 10328 26210 10362 26244
rect 10396 26210 10430 26244
rect 10464 26210 10498 26244
rect 10532 26210 10566 26244
rect 10600 26210 10634 26244
rect 10668 26210 10702 26244
rect 10736 26210 10770 26244
rect 10804 26210 10838 26244
rect 10872 26210 10906 26244
rect 10940 26210 10974 26244
rect 11008 26210 11042 26244
rect 11076 26210 11110 26244
rect 11144 26210 11178 26244
rect 11212 26210 11246 26244
rect 11280 26210 11314 26244
rect 11348 26210 11382 26244
rect 11416 26210 11450 26244
rect 11484 26210 11518 26244
rect 11552 26210 11586 26244
rect 11620 26210 11654 26244
rect 11688 26210 11722 26244
rect 11756 26210 11790 26244
rect 11824 26210 11858 26244
rect 11892 26210 11926 26244
rect 11960 26210 11994 26244
rect 12028 26210 12062 26244
rect 12096 26210 12130 26244
rect 12164 26210 12198 26244
rect 12232 26210 12266 26244
rect 12300 26210 12334 26244
rect 12368 26210 12402 26244
rect 12436 26210 12470 26244
rect 12504 26210 12538 26244
rect 12572 26210 12606 26244
rect 12640 26210 12674 26244
rect 12708 26210 12742 26244
rect 12776 26210 12810 26244
rect 12844 26210 12878 26244
rect 12912 26210 12946 26244
rect 12980 26210 13014 26244
rect 13048 26210 13082 26244
rect 13116 26210 13150 26244
rect 13184 26210 13218 26244
rect 13252 26210 13286 26244
rect 13320 26210 13354 26244
rect 13388 26210 13422 26244
rect 13456 26210 13490 26244
rect 13524 26210 13558 26244
rect 13592 26210 13626 26244
rect 13660 26210 13694 26244
rect 13728 26210 13762 26244
rect 13796 26210 13830 26244
rect 13864 26210 13898 26244
rect 13932 26210 13966 26244
rect 14000 26210 14034 26244
rect 14068 26210 14102 26244
rect 14136 26210 14170 26244
rect 14204 26210 14238 26244
rect 14272 26210 14306 26244
rect 14340 26210 14374 26244
rect 14408 26210 14442 26244
rect 14476 26210 14510 26244
rect 14544 26210 14578 26244
rect 14612 26210 14646 26244
rect 14680 26210 14714 26244
rect 14748 26210 14782 26244
rect 14816 26210 14850 26244
rect 14884 26210 14918 26244
rect 69 26138 103 26172
rect 138 26138 172 26172
rect 207 26138 241 26172
rect 276 26138 310 26172
rect 345 26138 379 26172
rect 414 26138 448 26172
rect 483 26138 517 26172
rect 552 26138 586 26172
rect 621 26138 655 26172
rect 690 26138 724 26172
rect 759 26138 793 26172
rect 828 26138 862 26172
rect 897 26138 931 26172
rect 966 26138 1000 26172
rect 1035 26138 1069 26172
rect 1104 26138 1138 26172
rect 1173 26138 1207 26172
rect 1242 26138 1276 26172
rect 1311 26138 1345 26172
rect 1380 26138 1414 26172
rect 1449 26138 1483 26172
rect 1518 26138 1552 26172
rect 1587 26138 1621 26172
rect 1656 26138 1690 26172
rect 1725 26138 1759 26172
rect 1794 26138 1828 26172
rect 1863 26138 1897 26172
rect 1932 26138 1966 26172
rect 2001 26138 2035 26172
rect 2070 26138 2104 26172
rect 2139 26138 2173 26172
rect 2208 26138 2242 26172
rect 2277 26138 2311 26172
rect 2346 26138 2380 26172
rect 2415 26138 2449 26172
rect 2484 26138 2518 26172
rect 2553 26138 2587 26172
rect 2622 26138 2656 26172
rect 2691 26138 2725 26172
rect 2760 26138 2794 26172
rect 2829 26138 2863 26172
rect 2898 26138 2932 26172
rect 2967 26138 3001 26172
rect 3036 26138 3070 26172
rect 3105 26138 3139 26172
rect 3174 26138 3208 26172
rect 3243 26138 3277 26172
rect 3312 26138 3346 26172
rect 3381 26138 3415 26172
rect 3450 26138 3484 26172
rect 3519 26138 3553 26172
rect 3588 26138 3622 26172
rect 3657 26138 3691 26172
rect 3726 26138 3760 26172
rect 3795 26138 3829 26172
rect 3864 26138 3898 26172
rect 3933 26138 3967 26172
rect 4002 26138 4036 26172
rect 4071 26138 4105 26172
rect 4140 26138 4174 26172
rect 4208 26138 4242 26172
rect 4276 26138 4310 26172
rect 4344 26138 4378 26172
rect 4412 26138 4446 26172
rect 4480 26138 4514 26172
rect 4548 26138 4582 26172
rect 4616 26138 4650 26172
rect 4684 26138 4718 26172
rect 4752 26138 4786 26172
rect 4820 26138 4854 26172
rect 4888 26138 4922 26172
rect 4956 26138 4990 26172
rect 5024 26138 5058 26172
rect 5092 26138 5126 26172
rect 5160 26138 5194 26172
rect 5228 26138 5262 26172
rect 5296 26138 5330 26172
rect 5364 26138 5398 26172
rect 5432 26138 5466 26172
rect 5500 26138 5534 26172
rect 5568 26138 5602 26172
rect 5636 26138 5670 26172
rect 5704 26138 5738 26172
rect 5772 26138 5806 26172
rect 5840 26138 5874 26172
rect 5908 26138 5942 26172
rect 5976 26138 6010 26172
rect 6044 26138 6078 26172
rect 6112 26138 6146 26172
rect 6180 26138 6214 26172
rect 6248 26138 6282 26172
rect 6316 26138 6350 26172
rect 6384 26138 6418 26172
rect 6452 26138 6486 26172
rect 6520 26138 6554 26172
rect 6588 26138 6622 26172
rect 6656 26138 6690 26172
rect 6724 26138 6758 26172
rect 6792 26138 6826 26172
rect 6860 26138 6894 26172
rect 6928 26138 6962 26172
rect 6996 26138 7030 26172
rect 7064 26138 7098 26172
rect 7132 26138 7166 26172
rect 7200 26138 7234 26172
rect 7268 26138 7302 26172
rect 7336 26138 7370 26172
rect 7404 26138 7438 26172
rect 7472 26138 7506 26172
rect 7540 26138 7574 26172
rect 7608 26138 7642 26172
rect 7676 26138 7710 26172
rect 7744 26138 7778 26172
rect 7812 26138 7846 26172
rect 7880 26138 7914 26172
rect 7948 26138 7982 26172
rect 8016 26138 8050 26172
rect 8084 26138 8118 26172
rect 8152 26138 8186 26172
rect 8220 26138 8254 26172
rect 8288 26138 8322 26172
rect 8356 26138 8390 26172
rect 8424 26138 8458 26172
rect 8492 26138 8526 26172
rect 8560 26138 8594 26172
rect 8628 26138 8662 26172
rect 8696 26138 8730 26172
rect 8764 26138 8798 26172
rect 8832 26138 8866 26172
rect 8900 26138 8934 26172
rect 8968 26138 9002 26172
rect 9036 26138 9070 26172
rect 9104 26138 9138 26172
rect 9172 26138 9206 26172
rect 9240 26138 9274 26172
rect 9308 26138 9342 26172
rect 9376 26138 9410 26172
rect 9444 26138 9478 26172
rect 9512 26138 9546 26172
rect 9580 26138 9614 26172
rect 9648 26138 9682 26172
rect 9716 26138 9750 26172
rect 9784 26138 9818 26172
rect 9852 26138 9886 26172
rect 9920 26138 9954 26172
rect 9988 26138 10022 26172
rect 10056 26138 10090 26172
rect 10124 26138 10158 26172
rect 10192 26138 10226 26172
rect 10260 26138 10294 26172
rect 10328 26138 10362 26172
rect 10396 26138 10430 26172
rect 10464 26138 10498 26172
rect 10532 26138 10566 26172
rect 10600 26138 10634 26172
rect 10668 26138 10702 26172
rect 10736 26138 10770 26172
rect 10804 26138 10838 26172
rect 10872 26138 10906 26172
rect 10940 26138 10974 26172
rect 11008 26138 11042 26172
rect 11076 26138 11110 26172
rect 11144 26138 11178 26172
rect 11212 26138 11246 26172
rect 11280 26138 11314 26172
rect 11348 26138 11382 26172
rect 11416 26138 11450 26172
rect 11484 26138 11518 26172
rect 11552 26138 11586 26172
rect 11620 26138 11654 26172
rect 11688 26138 11722 26172
rect 11756 26138 11790 26172
rect 11824 26138 11858 26172
rect 11892 26138 11926 26172
rect 11960 26138 11994 26172
rect 12028 26138 12062 26172
rect 12096 26138 12130 26172
rect 12164 26138 12198 26172
rect 12232 26138 12266 26172
rect 12300 26138 12334 26172
rect 12368 26138 12402 26172
rect 12436 26138 12470 26172
rect 12504 26138 12538 26172
rect 12572 26138 12606 26172
rect 12640 26138 12674 26172
rect 12708 26138 12742 26172
rect 12776 26138 12810 26172
rect 12844 26138 12878 26172
rect 12912 26138 12946 26172
rect 12980 26138 13014 26172
rect 13048 26138 13082 26172
rect 13116 26138 13150 26172
rect 13184 26138 13218 26172
rect 13252 26138 13286 26172
rect 13320 26138 13354 26172
rect 13388 26138 13422 26172
rect 13456 26138 13490 26172
rect 13524 26138 13558 26172
rect 13592 26138 13626 26172
rect 13660 26138 13694 26172
rect 13728 26138 13762 26172
rect 13796 26138 13830 26172
rect 13864 26138 13898 26172
rect 13932 26138 13966 26172
rect 14000 26138 14034 26172
rect 14068 26138 14102 26172
rect 14136 26138 14170 26172
rect 14204 26138 14238 26172
rect 14272 26138 14306 26172
rect 14340 26138 14374 26172
rect 14408 26138 14442 26172
rect 14476 26138 14510 26172
rect 14544 26138 14578 26172
rect 14612 26138 14646 26172
rect 14680 26138 14714 26172
rect 14748 26138 14782 26172
rect 14816 26138 14850 26172
rect 14884 26138 14918 26172
rect 69 26066 103 26100
rect 138 26066 172 26100
rect 207 26066 241 26100
rect 276 26066 310 26100
rect 345 26066 379 26100
rect 414 26066 448 26100
rect 483 26066 517 26100
rect 552 26066 586 26100
rect 621 26066 655 26100
rect 690 26066 724 26100
rect 759 26066 793 26100
rect 828 26066 862 26100
rect 897 26066 931 26100
rect 966 26066 1000 26100
rect 1035 26066 1069 26100
rect 1104 26066 1138 26100
rect 1173 26066 1207 26100
rect 1242 26066 1276 26100
rect 1311 26066 1345 26100
rect 1380 26066 1414 26100
rect 1449 26066 1483 26100
rect 1518 26066 1552 26100
rect 1587 26066 1621 26100
rect 1656 26066 1690 26100
rect 1725 26066 1759 26100
rect 1794 26066 1828 26100
rect 1863 26066 1897 26100
rect 1932 26066 1966 26100
rect 2001 26066 2035 26100
rect 2070 26066 2104 26100
rect 2139 26066 2173 26100
rect 2208 26066 2242 26100
rect 2277 26066 2311 26100
rect 2346 26066 2380 26100
rect 2415 26066 2449 26100
rect 2484 26066 2518 26100
rect 2553 26066 2587 26100
rect 2622 26066 2656 26100
rect 2691 26066 2725 26100
rect 2760 26066 2794 26100
rect 2829 26066 2863 26100
rect 2898 26066 2932 26100
rect 2967 26066 3001 26100
rect 3036 26066 3070 26100
rect 3105 26066 3139 26100
rect 3174 26066 3208 26100
rect 3243 26066 3277 26100
rect 3312 26066 3346 26100
rect 3381 26066 3415 26100
rect 3450 26066 3484 26100
rect 3519 26066 3553 26100
rect 3588 26066 3622 26100
rect 3657 26066 3691 26100
rect 3726 26066 3760 26100
rect 3795 26066 3829 26100
rect 3864 26066 3898 26100
rect 3933 26066 3967 26100
rect 4002 26066 4036 26100
rect 4071 26066 4105 26100
rect 4140 26066 4174 26100
rect 4208 26066 4242 26100
rect 4276 26066 4310 26100
rect 4344 26066 4378 26100
rect 4412 26066 4446 26100
rect 4480 26066 4514 26100
rect 4548 26066 4582 26100
rect 4616 26066 4650 26100
rect 4684 26066 4718 26100
rect 4752 26066 4786 26100
rect 4820 26066 4854 26100
rect 4888 26066 4922 26100
rect 4956 26066 4990 26100
rect 5024 26066 5058 26100
rect 5092 26066 5126 26100
rect 5160 26066 5194 26100
rect 5228 26066 5262 26100
rect 5296 26066 5330 26100
rect 5364 26066 5398 26100
rect 5432 26066 5466 26100
rect 5500 26066 5534 26100
rect 5568 26066 5602 26100
rect 5636 26066 5670 26100
rect 5704 26066 5738 26100
rect 5772 26066 5806 26100
rect 5840 26066 5874 26100
rect 5908 26066 5942 26100
rect 5976 26066 6010 26100
rect 6044 26066 6078 26100
rect 6112 26066 6146 26100
rect 6180 26066 6214 26100
rect 6248 26066 6282 26100
rect 6316 26066 6350 26100
rect 6384 26066 6418 26100
rect 6452 26066 6486 26100
rect 6520 26066 6554 26100
rect 6588 26066 6622 26100
rect 6656 26066 6690 26100
rect 6724 26066 6758 26100
rect 6792 26066 6826 26100
rect 6860 26066 6894 26100
rect 6928 26066 6962 26100
rect 6996 26066 7030 26100
rect 7064 26066 7098 26100
rect 7132 26066 7166 26100
rect 7200 26066 7234 26100
rect 7268 26066 7302 26100
rect 7336 26066 7370 26100
rect 7404 26066 7438 26100
rect 7472 26066 7506 26100
rect 7540 26066 7574 26100
rect 7608 26066 7642 26100
rect 7676 26066 7710 26100
rect 7744 26066 7778 26100
rect 7812 26066 7846 26100
rect 7880 26066 7914 26100
rect 7948 26066 7982 26100
rect 8016 26066 8050 26100
rect 8084 26066 8118 26100
rect 8152 26066 8186 26100
rect 8220 26066 8254 26100
rect 8288 26066 8322 26100
rect 8356 26066 8390 26100
rect 8424 26066 8458 26100
rect 8492 26066 8526 26100
rect 8560 26066 8594 26100
rect 8628 26066 8662 26100
rect 8696 26066 8730 26100
rect 8764 26066 8798 26100
rect 8832 26066 8866 26100
rect 8900 26066 8934 26100
rect 8968 26066 9002 26100
rect 9036 26066 9070 26100
rect 9104 26066 9138 26100
rect 9172 26066 9206 26100
rect 9240 26066 9274 26100
rect 9308 26066 9342 26100
rect 9376 26066 9410 26100
rect 9444 26066 9478 26100
rect 9512 26066 9546 26100
rect 9580 26066 9614 26100
rect 9648 26066 9682 26100
rect 9716 26066 9750 26100
rect 9784 26066 9818 26100
rect 9852 26066 9886 26100
rect 9920 26066 9954 26100
rect 9988 26066 10022 26100
rect 10056 26066 10090 26100
rect 10124 26066 10158 26100
rect 10192 26066 10226 26100
rect 10260 26066 10294 26100
rect 10328 26066 10362 26100
rect 10396 26066 10430 26100
rect 10464 26066 10498 26100
rect 10532 26066 10566 26100
rect 10600 26066 10634 26100
rect 10668 26066 10702 26100
rect 10736 26066 10770 26100
rect 10804 26066 10838 26100
rect 10872 26066 10906 26100
rect 10940 26066 10974 26100
rect 11008 26066 11042 26100
rect 11076 26066 11110 26100
rect 11144 26066 11178 26100
rect 11212 26066 11246 26100
rect 11280 26066 11314 26100
rect 11348 26066 11382 26100
rect 11416 26066 11450 26100
rect 11484 26066 11518 26100
rect 11552 26066 11586 26100
rect 11620 26066 11654 26100
rect 11688 26066 11722 26100
rect 11756 26066 11790 26100
rect 11824 26066 11858 26100
rect 11892 26066 11926 26100
rect 11960 26066 11994 26100
rect 12028 26066 12062 26100
rect 12096 26066 12130 26100
rect 12164 26066 12198 26100
rect 12232 26066 12266 26100
rect 12300 26066 12334 26100
rect 12368 26066 12402 26100
rect 12436 26066 12470 26100
rect 12504 26066 12538 26100
rect 12572 26066 12606 26100
rect 12640 26066 12674 26100
rect 12708 26066 12742 26100
rect 12776 26066 12810 26100
rect 12844 26066 12878 26100
rect 12912 26066 12946 26100
rect 12980 26066 13014 26100
rect 13048 26066 13082 26100
rect 13116 26066 13150 26100
rect 13184 26066 13218 26100
rect 13252 26066 13286 26100
rect 13320 26066 13354 26100
rect 13388 26066 13422 26100
rect 13456 26066 13490 26100
rect 13524 26066 13558 26100
rect 13592 26066 13626 26100
rect 13660 26066 13694 26100
rect 13728 26066 13762 26100
rect 13796 26066 13830 26100
rect 13864 26066 13898 26100
rect 13932 26066 13966 26100
rect 14000 26066 14034 26100
rect 14068 26066 14102 26100
rect 14136 26066 14170 26100
rect 14204 26066 14238 26100
rect 14272 26066 14306 26100
rect 14340 26066 14374 26100
rect 14408 26066 14442 26100
rect 14476 26066 14510 26100
rect 14544 26066 14578 26100
rect 14612 26066 14646 26100
rect 14680 26066 14714 26100
rect 14748 26066 14782 26100
rect 14816 26066 14850 26100
rect 14884 26066 14918 26100
rect 69 25994 103 26028
rect 138 25994 172 26028
rect 207 25994 241 26028
rect 276 25994 310 26028
rect 345 25994 379 26028
rect 414 25994 448 26028
rect 483 25994 517 26028
rect 552 25994 586 26028
rect 621 25994 655 26028
rect 690 25994 724 26028
rect 759 25994 793 26028
rect 828 25994 862 26028
rect 897 25994 931 26028
rect 966 25994 1000 26028
rect 1035 25994 1069 26028
rect 1104 25994 1138 26028
rect 1173 25994 1207 26028
rect 1242 25994 1276 26028
rect 1311 25994 1345 26028
rect 1380 25994 1414 26028
rect 1449 25994 1483 26028
rect 1518 25994 1552 26028
rect 1587 25994 1621 26028
rect 1656 25994 1690 26028
rect 1725 25994 1759 26028
rect 1794 25994 1828 26028
rect 1863 25994 1897 26028
rect 1932 25994 1966 26028
rect 2001 25994 2035 26028
rect 2070 25994 2104 26028
rect 2139 25994 2173 26028
rect 2208 25994 2242 26028
rect 2277 25994 2311 26028
rect 2346 25994 2380 26028
rect 2415 25994 2449 26028
rect 2484 25994 2518 26028
rect 2553 25994 2587 26028
rect 2622 25994 2656 26028
rect 2691 25994 2725 26028
rect 2760 25994 2794 26028
rect 2829 25994 2863 26028
rect 2898 25994 2932 26028
rect 2967 25994 3001 26028
rect 3036 25994 3070 26028
rect 3105 25994 3139 26028
rect 3174 25994 3208 26028
rect 3243 25994 3277 26028
rect 3312 25994 3346 26028
rect 3381 25994 3415 26028
rect 3450 25994 3484 26028
rect 3519 25994 3553 26028
rect 3588 25994 3622 26028
rect 3657 25994 3691 26028
rect 3726 25994 3760 26028
rect 3795 25994 3829 26028
rect 3864 25994 3898 26028
rect 3933 25994 3967 26028
rect 4002 25994 4036 26028
rect 4071 25994 4105 26028
rect 4140 25994 4174 26028
rect 4208 25994 4242 26028
rect 4276 25994 4310 26028
rect 4344 25994 4378 26028
rect 4412 25994 4446 26028
rect 4480 25994 4514 26028
rect 4548 25994 4582 26028
rect 4616 25994 4650 26028
rect 4684 25994 4718 26028
rect 4752 25994 4786 26028
rect 4820 25994 4854 26028
rect 4888 25994 4922 26028
rect 4956 25994 4990 26028
rect 5024 25994 5058 26028
rect 5092 25994 5126 26028
rect 5160 25994 5194 26028
rect 5228 25994 5262 26028
rect 5296 25994 5330 26028
rect 5364 25994 5398 26028
rect 5432 25994 5466 26028
rect 5500 25994 5534 26028
rect 5568 25994 5602 26028
rect 5636 25994 5670 26028
rect 5704 25994 5738 26028
rect 5772 25994 5806 26028
rect 5840 25994 5874 26028
rect 5908 25994 5942 26028
rect 5976 25994 6010 26028
rect 6044 25994 6078 26028
rect 6112 25994 6146 26028
rect 6180 25994 6214 26028
rect 6248 25994 6282 26028
rect 6316 25994 6350 26028
rect 6384 25994 6418 26028
rect 6452 25994 6486 26028
rect 6520 25994 6554 26028
rect 6588 25994 6622 26028
rect 6656 25994 6690 26028
rect 6724 25994 6758 26028
rect 6792 25994 6826 26028
rect 6860 25994 6894 26028
rect 6928 25994 6962 26028
rect 6996 25994 7030 26028
rect 7064 25994 7098 26028
rect 7132 25994 7166 26028
rect 7200 25994 7234 26028
rect 7268 25994 7302 26028
rect 7336 25994 7370 26028
rect 7404 25994 7438 26028
rect 7472 25994 7506 26028
rect 7540 25994 7574 26028
rect 7608 25994 7642 26028
rect 7676 25994 7710 26028
rect 7744 25994 7778 26028
rect 7812 25994 7846 26028
rect 7880 25994 7914 26028
rect 7948 25994 7982 26028
rect 8016 25994 8050 26028
rect 8084 25994 8118 26028
rect 8152 25994 8186 26028
rect 8220 25994 8254 26028
rect 8288 25994 8322 26028
rect 8356 25994 8390 26028
rect 8424 25994 8458 26028
rect 8492 25994 8526 26028
rect 8560 25994 8594 26028
rect 8628 25994 8662 26028
rect 8696 25994 8730 26028
rect 8764 25994 8798 26028
rect 8832 25994 8866 26028
rect 8900 25994 8934 26028
rect 8968 25994 9002 26028
rect 9036 25994 9070 26028
rect 9104 25994 9138 26028
rect 9172 25994 9206 26028
rect 9240 25994 9274 26028
rect 9308 25994 9342 26028
rect 9376 25994 9410 26028
rect 9444 25994 9478 26028
rect 9512 25994 9546 26028
rect 9580 25994 9614 26028
rect 9648 25994 9682 26028
rect 9716 25994 9750 26028
rect 9784 25994 9818 26028
rect 9852 25994 9886 26028
rect 9920 25994 9954 26028
rect 9988 25994 10022 26028
rect 10056 25994 10090 26028
rect 10124 25994 10158 26028
rect 10192 25994 10226 26028
rect 10260 25994 10294 26028
rect 10328 25994 10362 26028
rect 10396 25994 10430 26028
rect 10464 25994 10498 26028
rect 10532 25994 10566 26028
rect 10600 25994 10634 26028
rect 10668 25994 10702 26028
rect 10736 25994 10770 26028
rect 10804 25994 10838 26028
rect 10872 25994 10906 26028
rect 10940 25994 10974 26028
rect 11008 25994 11042 26028
rect 11076 25994 11110 26028
rect 11144 25994 11178 26028
rect 11212 25994 11246 26028
rect 11280 25994 11314 26028
rect 11348 25994 11382 26028
rect 11416 25994 11450 26028
rect 11484 25994 11518 26028
rect 11552 25994 11586 26028
rect 11620 25994 11654 26028
rect 11688 25994 11722 26028
rect 11756 25994 11790 26028
rect 11824 25994 11858 26028
rect 11892 25994 11926 26028
rect 11960 25994 11994 26028
rect 12028 25994 12062 26028
rect 12096 25994 12130 26028
rect 12164 25994 12198 26028
rect 12232 25994 12266 26028
rect 12300 25994 12334 26028
rect 12368 25994 12402 26028
rect 12436 25994 12470 26028
rect 12504 25994 12538 26028
rect 12572 25994 12606 26028
rect 12640 25994 12674 26028
rect 12708 25994 12742 26028
rect 12776 25994 12810 26028
rect 12844 25994 12878 26028
rect 12912 25994 12946 26028
rect 12980 25994 13014 26028
rect 13048 25994 13082 26028
rect 13116 25994 13150 26028
rect 13184 25994 13218 26028
rect 13252 25994 13286 26028
rect 13320 25994 13354 26028
rect 13388 25994 13422 26028
rect 13456 25994 13490 26028
rect 13524 25994 13558 26028
rect 13592 25994 13626 26028
rect 13660 25994 13694 26028
rect 13728 25994 13762 26028
rect 13796 25994 13830 26028
rect 13864 25994 13898 26028
rect 13932 25994 13966 26028
rect 14000 25994 14034 26028
rect 14068 25994 14102 26028
rect 14136 25994 14170 26028
rect 14204 25994 14238 26028
rect 14272 25994 14306 26028
rect 14340 25994 14374 26028
rect 14408 25994 14442 26028
rect 14476 25994 14510 26028
rect 14544 25994 14578 26028
rect 14612 25994 14646 26028
rect 14680 25994 14714 26028
rect 14748 25994 14782 26028
rect 14816 25994 14850 26028
rect 14884 25994 14918 26028
rect 69 25922 103 25956
rect 138 25922 172 25956
rect 207 25922 241 25956
rect 276 25922 310 25956
rect 345 25922 379 25956
rect 414 25922 448 25956
rect 483 25922 517 25956
rect 552 25922 586 25956
rect 621 25922 655 25956
rect 690 25922 724 25956
rect 759 25922 793 25956
rect 828 25922 862 25956
rect 897 25922 931 25956
rect 966 25922 1000 25956
rect 1035 25922 1069 25956
rect 1104 25922 1138 25956
rect 1173 25922 1207 25956
rect 1242 25922 1276 25956
rect 1311 25922 1345 25956
rect 1380 25922 1414 25956
rect 1449 25922 1483 25956
rect 1518 25922 1552 25956
rect 1587 25922 1621 25956
rect 1656 25922 1690 25956
rect 1725 25922 1759 25956
rect 1794 25922 1828 25956
rect 1863 25922 1897 25956
rect 1932 25922 1966 25956
rect 2001 25922 2035 25956
rect 2070 25922 2104 25956
rect 2139 25922 2173 25956
rect 2208 25922 2242 25956
rect 2277 25922 2311 25956
rect 2346 25922 2380 25956
rect 2415 25922 2449 25956
rect 2484 25922 2518 25956
rect 2553 25922 2587 25956
rect 2622 25922 2656 25956
rect 2691 25922 2725 25956
rect 2760 25922 2794 25956
rect 2829 25922 2863 25956
rect 2898 25922 2932 25956
rect 2967 25922 3001 25956
rect 3036 25922 3070 25956
rect 3105 25922 3139 25956
rect 3174 25922 3208 25956
rect 3243 25922 3277 25956
rect 3312 25922 3346 25956
rect 3381 25922 3415 25956
rect 3450 25922 3484 25956
rect 3519 25922 3553 25956
rect 3588 25922 3622 25956
rect 3657 25922 3691 25956
rect 3726 25922 3760 25956
rect 3795 25922 3829 25956
rect 3864 25922 3898 25956
rect 3933 25922 3967 25956
rect 4002 25922 4036 25956
rect 4071 25922 4105 25956
rect 4140 25922 4174 25956
rect 4208 25922 4242 25956
rect 4276 25922 4310 25956
rect 4344 25922 4378 25956
rect 4412 25922 4446 25956
rect 4480 25922 4514 25956
rect 4548 25922 4582 25956
rect 4616 25922 4650 25956
rect 4684 25922 4718 25956
rect 4752 25922 4786 25956
rect 4820 25922 4854 25956
rect 4888 25922 4922 25956
rect 4956 25922 4990 25956
rect 5024 25922 5058 25956
rect 5092 25922 5126 25956
rect 5160 25922 5194 25956
rect 5228 25922 5262 25956
rect 5296 25922 5330 25956
rect 5364 25922 5398 25956
rect 5432 25922 5466 25956
rect 5500 25922 5534 25956
rect 5568 25922 5602 25956
rect 5636 25922 5670 25956
rect 5704 25922 5738 25956
rect 5772 25922 5806 25956
rect 5840 25922 5874 25956
rect 5908 25922 5942 25956
rect 5976 25922 6010 25956
rect 6044 25922 6078 25956
rect 6112 25922 6146 25956
rect 6180 25922 6214 25956
rect 6248 25922 6282 25956
rect 6316 25922 6350 25956
rect 6384 25922 6418 25956
rect 6452 25922 6486 25956
rect 6520 25922 6554 25956
rect 6588 25922 6622 25956
rect 6656 25922 6690 25956
rect 6724 25922 6758 25956
rect 6792 25922 6826 25956
rect 6860 25922 6894 25956
rect 6928 25922 6962 25956
rect 6996 25922 7030 25956
rect 7064 25922 7098 25956
rect 7132 25922 7166 25956
rect 7200 25922 7234 25956
rect 7268 25922 7302 25956
rect 7336 25922 7370 25956
rect 7404 25922 7438 25956
rect 7472 25922 7506 25956
rect 7540 25922 7574 25956
rect 7608 25922 7642 25956
rect 7676 25922 7710 25956
rect 7744 25922 7778 25956
rect 7812 25922 7846 25956
rect 7880 25922 7914 25956
rect 7948 25922 7982 25956
rect 8016 25922 8050 25956
rect 8084 25922 8118 25956
rect 8152 25922 8186 25956
rect 8220 25922 8254 25956
rect 8288 25922 8322 25956
rect 8356 25922 8390 25956
rect 8424 25922 8458 25956
rect 8492 25922 8526 25956
rect 8560 25922 8594 25956
rect 8628 25922 8662 25956
rect 8696 25922 8730 25956
rect 8764 25922 8798 25956
rect 8832 25922 8866 25956
rect 8900 25922 8934 25956
rect 8968 25922 9002 25956
rect 9036 25922 9070 25956
rect 9104 25922 9138 25956
rect 9172 25922 9206 25956
rect 9240 25922 9274 25956
rect 9308 25922 9342 25956
rect 9376 25922 9410 25956
rect 9444 25922 9478 25956
rect 9512 25922 9546 25956
rect 9580 25922 9614 25956
rect 9648 25922 9682 25956
rect 9716 25922 9750 25956
rect 9784 25922 9818 25956
rect 9852 25922 9886 25956
rect 9920 25922 9954 25956
rect 9988 25922 10022 25956
rect 10056 25922 10090 25956
rect 10124 25922 10158 25956
rect 10192 25922 10226 25956
rect 10260 25922 10294 25956
rect 10328 25922 10362 25956
rect 10396 25922 10430 25956
rect 10464 25922 10498 25956
rect 10532 25922 10566 25956
rect 10600 25922 10634 25956
rect 10668 25922 10702 25956
rect 10736 25922 10770 25956
rect 10804 25922 10838 25956
rect 10872 25922 10906 25956
rect 10940 25922 10974 25956
rect 11008 25922 11042 25956
rect 11076 25922 11110 25956
rect 11144 25922 11178 25956
rect 11212 25922 11246 25956
rect 11280 25922 11314 25956
rect 11348 25922 11382 25956
rect 11416 25922 11450 25956
rect 11484 25922 11518 25956
rect 11552 25922 11586 25956
rect 11620 25922 11654 25956
rect 11688 25922 11722 25956
rect 11756 25922 11790 25956
rect 11824 25922 11858 25956
rect 11892 25922 11926 25956
rect 11960 25922 11994 25956
rect 12028 25922 12062 25956
rect 12096 25922 12130 25956
rect 12164 25922 12198 25956
rect 12232 25922 12266 25956
rect 12300 25922 12334 25956
rect 12368 25922 12402 25956
rect 12436 25922 12470 25956
rect 12504 25922 12538 25956
rect 12572 25922 12606 25956
rect 12640 25922 12674 25956
rect 12708 25922 12742 25956
rect 12776 25922 12810 25956
rect 12844 25922 12878 25956
rect 12912 25922 12946 25956
rect 12980 25922 13014 25956
rect 13048 25922 13082 25956
rect 13116 25922 13150 25956
rect 13184 25922 13218 25956
rect 13252 25922 13286 25956
rect 13320 25922 13354 25956
rect 13388 25922 13422 25956
rect 13456 25922 13490 25956
rect 13524 25922 13558 25956
rect 13592 25922 13626 25956
rect 13660 25922 13694 25956
rect 13728 25922 13762 25956
rect 13796 25922 13830 25956
rect 13864 25922 13898 25956
rect 13932 25922 13966 25956
rect 14000 25922 14034 25956
rect 14068 25922 14102 25956
rect 14136 25922 14170 25956
rect 14204 25922 14238 25956
rect 14272 25922 14306 25956
rect 14340 25922 14374 25956
rect 14408 25922 14442 25956
rect 14476 25922 14510 25956
rect 14544 25922 14578 25956
rect 14612 25922 14646 25956
rect 14680 25922 14714 25956
rect 14748 25922 14782 25956
rect 14816 25922 14850 25956
rect 14884 25922 14918 25956
rect 69 25850 103 25884
rect 138 25850 172 25884
rect 207 25850 241 25884
rect 276 25850 310 25884
rect 345 25850 379 25884
rect 414 25850 448 25884
rect 483 25850 517 25884
rect 552 25850 586 25884
rect 621 25850 655 25884
rect 690 25850 724 25884
rect 759 25850 793 25884
rect 828 25850 862 25884
rect 897 25850 931 25884
rect 966 25850 1000 25884
rect 1035 25850 1069 25884
rect 1104 25850 1138 25884
rect 1173 25850 1207 25884
rect 1242 25850 1276 25884
rect 1311 25850 1345 25884
rect 1380 25850 1414 25884
rect 1449 25850 1483 25884
rect 1518 25850 1552 25884
rect 1587 25850 1621 25884
rect 1656 25850 1690 25884
rect 1725 25850 1759 25884
rect 1794 25850 1828 25884
rect 1863 25850 1897 25884
rect 1932 25850 1966 25884
rect 2001 25850 2035 25884
rect 2070 25850 2104 25884
rect 2139 25850 2173 25884
rect 2208 25850 2242 25884
rect 2277 25850 2311 25884
rect 2346 25850 2380 25884
rect 2415 25850 2449 25884
rect 2484 25850 2518 25884
rect 2553 25850 2587 25884
rect 2622 25850 2656 25884
rect 2691 25850 2725 25884
rect 2760 25850 2794 25884
rect 2829 25850 2863 25884
rect 2898 25850 2932 25884
rect 2967 25850 3001 25884
rect 3036 25850 3070 25884
rect 3105 25850 3139 25884
rect 3174 25850 3208 25884
rect 3243 25850 3277 25884
rect 3312 25850 3346 25884
rect 3381 25850 3415 25884
rect 3450 25850 3484 25884
rect 3519 25850 3553 25884
rect 3588 25850 3622 25884
rect 3657 25850 3691 25884
rect 3726 25850 3760 25884
rect 3795 25850 3829 25884
rect 3864 25850 3898 25884
rect 3933 25850 3967 25884
rect 4002 25850 4036 25884
rect 4071 25850 4105 25884
rect 4140 25850 4174 25884
rect 4208 25850 4242 25884
rect 4276 25850 4310 25884
rect 4344 25850 4378 25884
rect 4412 25850 4446 25884
rect 4480 25850 4514 25884
rect 4548 25850 4582 25884
rect 4616 25850 4650 25884
rect 4684 25850 4718 25884
rect 4752 25850 4786 25884
rect 4820 25850 4854 25884
rect 4888 25850 4922 25884
rect 4956 25850 4990 25884
rect 5024 25850 5058 25884
rect 5092 25850 5126 25884
rect 5160 25850 5194 25884
rect 5228 25850 5262 25884
rect 5296 25850 5330 25884
rect 5364 25850 5398 25884
rect 5432 25850 5466 25884
rect 5500 25850 5534 25884
rect 5568 25850 5602 25884
rect 5636 25850 5670 25884
rect 5704 25850 5738 25884
rect 5772 25850 5806 25884
rect 5840 25850 5874 25884
rect 5908 25850 5942 25884
rect 5976 25850 6010 25884
rect 6044 25850 6078 25884
rect 6112 25850 6146 25884
rect 6180 25850 6214 25884
rect 6248 25850 6282 25884
rect 6316 25850 6350 25884
rect 6384 25850 6418 25884
rect 6452 25850 6486 25884
rect 6520 25850 6554 25884
rect 6588 25850 6622 25884
rect 6656 25850 6690 25884
rect 6724 25850 6758 25884
rect 6792 25850 6826 25884
rect 6860 25850 6894 25884
rect 6928 25850 6962 25884
rect 6996 25850 7030 25884
rect 7064 25850 7098 25884
rect 7132 25850 7166 25884
rect 7200 25850 7234 25884
rect 7268 25850 7302 25884
rect 7336 25850 7370 25884
rect 7404 25850 7438 25884
rect 7472 25850 7506 25884
rect 7540 25850 7574 25884
rect 7608 25850 7642 25884
rect 7676 25850 7710 25884
rect 7744 25850 7778 25884
rect 7812 25850 7846 25884
rect 7880 25850 7914 25884
rect 7948 25850 7982 25884
rect 8016 25850 8050 25884
rect 8084 25850 8118 25884
rect 8152 25850 8186 25884
rect 8220 25850 8254 25884
rect 8288 25850 8322 25884
rect 8356 25850 8390 25884
rect 8424 25850 8458 25884
rect 8492 25850 8526 25884
rect 8560 25850 8594 25884
rect 8628 25850 8662 25884
rect 8696 25850 8730 25884
rect 8764 25850 8798 25884
rect 8832 25850 8866 25884
rect 8900 25850 8934 25884
rect 8968 25850 9002 25884
rect 9036 25850 9070 25884
rect 9104 25850 9138 25884
rect 9172 25850 9206 25884
rect 9240 25850 9274 25884
rect 9308 25850 9342 25884
rect 9376 25850 9410 25884
rect 9444 25850 9478 25884
rect 9512 25850 9546 25884
rect 9580 25850 9614 25884
rect 9648 25850 9682 25884
rect 9716 25850 9750 25884
rect 9784 25850 9818 25884
rect 9852 25850 9886 25884
rect 9920 25850 9954 25884
rect 9988 25850 10022 25884
rect 10056 25850 10090 25884
rect 10124 25850 10158 25884
rect 10192 25850 10226 25884
rect 10260 25850 10294 25884
rect 10328 25850 10362 25884
rect 10396 25850 10430 25884
rect 10464 25850 10498 25884
rect 10532 25850 10566 25884
rect 10600 25850 10634 25884
rect 10668 25850 10702 25884
rect 10736 25850 10770 25884
rect 10804 25850 10838 25884
rect 10872 25850 10906 25884
rect 10940 25850 10974 25884
rect 11008 25850 11042 25884
rect 11076 25850 11110 25884
rect 11144 25850 11178 25884
rect 11212 25850 11246 25884
rect 11280 25850 11314 25884
rect 11348 25850 11382 25884
rect 11416 25850 11450 25884
rect 11484 25850 11518 25884
rect 11552 25850 11586 25884
rect 11620 25850 11654 25884
rect 11688 25850 11722 25884
rect 11756 25850 11790 25884
rect 11824 25850 11858 25884
rect 11892 25850 11926 25884
rect 11960 25850 11994 25884
rect 12028 25850 12062 25884
rect 12096 25850 12130 25884
rect 12164 25850 12198 25884
rect 12232 25850 12266 25884
rect 12300 25850 12334 25884
rect 12368 25850 12402 25884
rect 12436 25850 12470 25884
rect 12504 25850 12538 25884
rect 12572 25850 12606 25884
rect 12640 25850 12674 25884
rect 12708 25850 12742 25884
rect 12776 25850 12810 25884
rect 12844 25850 12878 25884
rect 12912 25850 12946 25884
rect 12980 25850 13014 25884
rect 13048 25850 13082 25884
rect 13116 25850 13150 25884
rect 13184 25850 13218 25884
rect 13252 25850 13286 25884
rect 13320 25850 13354 25884
rect 13388 25850 13422 25884
rect 13456 25850 13490 25884
rect 13524 25850 13558 25884
rect 13592 25850 13626 25884
rect 13660 25850 13694 25884
rect 13728 25850 13762 25884
rect 13796 25850 13830 25884
rect 13864 25850 13898 25884
rect 13932 25850 13966 25884
rect 14000 25850 14034 25884
rect 14068 25850 14102 25884
rect 14136 25850 14170 25884
rect 14204 25850 14238 25884
rect 14272 25850 14306 25884
rect 14340 25850 14374 25884
rect 14408 25850 14442 25884
rect 14476 25850 14510 25884
rect 14544 25850 14578 25884
rect 14612 25850 14646 25884
rect 14680 25850 14714 25884
rect 14748 25850 14782 25884
rect 14816 25850 14850 25884
rect 14884 25850 14918 25884
rect 69 25778 103 25812
rect 138 25778 172 25812
rect 207 25778 241 25812
rect 276 25778 310 25812
rect 345 25778 379 25812
rect 414 25778 448 25812
rect 483 25778 517 25812
rect 552 25778 586 25812
rect 621 25778 655 25812
rect 690 25778 724 25812
rect 759 25778 793 25812
rect 828 25778 862 25812
rect 897 25778 931 25812
rect 966 25778 1000 25812
rect 1035 25778 1069 25812
rect 1104 25778 1138 25812
rect 1173 25778 1207 25812
rect 1242 25778 1276 25812
rect 1311 25778 1345 25812
rect 1380 25778 1414 25812
rect 1449 25778 1483 25812
rect 1518 25778 1552 25812
rect 1587 25778 1621 25812
rect 1656 25778 1690 25812
rect 1725 25778 1759 25812
rect 1794 25778 1828 25812
rect 1863 25778 1897 25812
rect 1932 25778 1966 25812
rect 2001 25778 2035 25812
rect 2070 25778 2104 25812
rect 2139 25778 2173 25812
rect 2208 25778 2242 25812
rect 2277 25778 2311 25812
rect 2346 25778 2380 25812
rect 2415 25778 2449 25812
rect 2484 25778 2518 25812
rect 2553 25778 2587 25812
rect 2622 25778 2656 25812
rect 2691 25778 2725 25812
rect 2760 25778 2794 25812
rect 2829 25778 2863 25812
rect 2898 25778 2932 25812
rect 2967 25778 3001 25812
rect 3036 25778 3070 25812
rect 3105 25778 3139 25812
rect 3174 25778 3208 25812
rect 3243 25778 3277 25812
rect 3312 25778 3346 25812
rect 3381 25778 3415 25812
rect 3450 25778 3484 25812
rect 3519 25778 3553 25812
rect 3588 25778 3622 25812
rect 3657 25778 3691 25812
rect 3726 25778 3760 25812
rect 3795 25778 3829 25812
rect 3864 25778 3898 25812
rect 3933 25778 3967 25812
rect 4002 25778 4036 25812
rect 4071 25778 4105 25812
rect 4140 25778 4174 25812
rect 4208 25778 4242 25812
rect 4276 25778 4310 25812
rect 4344 25778 4378 25812
rect 4412 25778 4446 25812
rect 4480 25778 4514 25812
rect 4548 25778 4582 25812
rect 4616 25778 4650 25812
rect 4684 25778 4718 25812
rect 4752 25778 4786 25812
rect 4820 25778 4854 25812
rect 4888 25778 4922 25812
rect 4956 25778 4990 25812
rect 5024 25778 5058 25812
rect 5092 25778 5126 25812
rect 5160 25778 5194 25812
rect 5228 25778 5262 25812
rect 5296 25778 5330 25812
rect 5364 25778 5398 25812
rect 5432 25778 5466 25812
rect 5500 25778 5534 25812
rect 5568 25778 5602 25812
rect 5636 25778 5670 25812
rect 5704 25778 5738 25812
rect 5772 25778 5806 25812
rect 5840 25778 5874 25812
rect 5908 25778 5942 25812
rect 5976 25778 6010 25812
rect 6044 25778 6078 25812
rect 6112 25778 6146 25812
rect 6180 25778 6214 25812
rect 6248 25778 6282 25812
rect 6316 25778 6350 25812
rect 6384 25778 6418 25812
rect 6452 25778 6486 25812
rect 6520 25778 6554 25812
rect 6588 25778 6622 25812
rect 6656 25778 6690 25812
rect 6724 25778 6758 25812
rect 6792 25778 6826 25812
rect 6860 25778 6894 25812
rect 6928 25778 6962 25812
rect 6996 25778 7030 25812
rect 7064 25778 7098 25812
rect 7132 25778 7166 25812
rect 7200 25778 7234 25812
rect 7268 25778 7302 25812
rect 7336 25778 7370 25812
rect 7404 25778 7438 25812
rect 7472 25778 7506 25812
rect 7540 25778 7574 25812
rect 7608 25778 7642 25812
rect 7676 25778 7710 25812
rect 7744 25778 7778 25812
rect 7812 25778 7846 25812
rect 7880 25778 7914 25812
rect 7948 25778 7982 25812
rect 8016 25778 8050 25812
rect 8084 25778 8118 25812
rect 8152 25778 8186 25812
rect 8220 25778 8254 25812
rect 8288 25778 8322 25812
rect 8356 25778 8390 25812
rect 8424 25778 8458 25812
rect 8492 25778 8526 25812
rect 8560 25778 8594 25812
rect 8628 25778 8662 25812
rect 8696 25778 8730 25812
rect 8764 25778 8798 25812
rect 8832 25778 8866 25812
rect 8900 25778 8934 25812
rect 8968 25778 9002 25812
rect 9036 25778 9070 25812
rect 9104 25778 9138 25812
rect 9172 25778 9206 25812
rect 9240 25778 9274 25812
rect 9308 25778 9342 25812
rect 9376 25778 9410 25812
rect 9444 25778 9478 25812
rect 9512 25778 9546 25812
rect 9580 25778 9614 25812
rect 9648 25778 9682 25812
rect 9716 25778 9750 25812
rect 9784 25778 9818 25812
rect 9852 25778 9886 25812
rect 9920 25778 9954 25812
rect 9988 25778 10022 25812
rect 10056 25778 10090 25812
rect 10124 25778 10158 25812
rect 10192 25778 10226 25812
rect 10260 25778 10294 25812
rect 10328 25778 10362 25812
rect 10396 25778 10430 25812
rect 10464 25778 10498 25812
rect 10532 25778 10566 25812
rect 10600 25778 10634 25812
rect 10668 25778 10702 25812
rect 10736 25778 10770 25812
rect 10804 25778 10838 25812
rect 10872 25778 10906 25812
rect 10940 25778 10974 25812
rect 11008 25778 11042 25812
rect 11076 25778 11110 25812
rect 11144 25778 11178 25812
rect 11212 25778 11246 25812
rect 11280 25778 11314 25812
rect 11348 25778 11382 25812
rect 11416 25778 11450 25812
rect 11484 25778 11518 25812
rect 11552 25778 11586 25812
rect 11620 25778 11654 25812
rect 11688 25778 11722 25812
rect 11756 25778 11790 25812
rect 11824 25778 11858 25812
rect 11892 25778 11926 25812
rect 11960 25778 11994 25812
rect 12028 25778 12062 25812
rect 12096 25778 12130 25812
rect 12164 25778 12198 25812
rect 12232 25778 12266 25812
rect 12300 25778 12334 25812
rect 12368 25778 12402 25812
rect 12436 25778 12470 25812
rect 12504 25778 12538 25812
rect 12572 25778 12606 25812
rect 12640 25778 12674 25812
rect 12708 25778 12742 25812
rect 12776 25778 12810 25812
rect 12844 25778 12878 25812
rect 12912 25778 12946 25812
rect 12980 25778 13014 25812
rect 13048 25778 13082 25812
rect 13116 25778 13150 25812
rect 13184 25778 13218 25812
rect 13252 25778 13286 25812
rect 13320 25778 13354 25812
rect 13388 25778 13422 25812
rect 13456 25778 13490 25812
rect 13524 25778 13558 25812
rect 13592 25778 13626 25812
rect 13660 25778 13694 25812
rect 13728 25778 13762 25812
rect 13796 25778 13830 25812
rect 13864 25778 13898 25812
rect 13932 25778 13966 25812
rect 14000 25778 14034 25812
rect 14068 25778 14102 25812
rect 14136 25778 14170 25812
rect 14204 25778 14238 25812
rect 14272 25778 14306 25812
rect 14340 25778 14374 25812
rect 14408 25778 14442 25812
rect 14476 25778 14510 25812
rect 14544 25778 14578 25812
rect 14612 25778 14646 25812
rect 14680 25778 14714 25812
rect 14748 25778 14782 25812
rect 14816 25778 14850 25812
rect 14884 25778 14918 25812
rect 69 25706 103 25740
rect 138 25706 172 25740
rect 207 25706 241 25740
rect 276 25706 310 25740
rect 345 25706 379 25740
rect 414 25706 448 25740
rect 483 25706 517 25740
rect 552 25706 586 25740
rect 621 25706 655 25740
rect 690 25706 724 25740
rect 759 25706 793 25740
rect 828 25706 862 25740
rect 897 25706 931 25740
rect 966 25706 1000 25740
rect 1035 25706 1069 25740
rect 1104 25706 1138 25740
rect 1173 25706 1207 25740
rect 1242 25706 1276 25740
rect 1311 25706 1345 25740
rect 1380 25706 1414 25740
rect 1449 25706 1483 25740
rect 1518 25706 1552 25740
rect 1587 25706 1621 25740
rect 1656 25706 1690 25740
rect 1725 25706 1759 25740
rect 1794 25706 1828 25740
rect 1863 25706 1897 25740
rect 1932 25706 1966 25740
rect 2001 25706 2035 25740
rect 2070 25706 2104 25740
rect 2139 25706 2173 25740
rect 2208 25706 2242 25740
rect 2277 25706 2311 25740
rect 2346 25706 2380 25740
rect 2415 25706 2449 25740
rect 2484 25706 2518 25740
rect 2553 25706 2587 25740
rect 2622 25706 2656 25740
rect 2691 25706 2725 25740
rect 2760 25706 2794 25740
rect 2829 25706 2863 25740
rect 2898 25706 2932 25740
rect 2967 25706 3001 25740
rect 3036 25706 3070 25740
rect 3105 25706 3139 25740
rect 3174 25706 3208 25740
rect 3243 25706 3277 25740
rect 3312 25706 3346 25740
rect 3381 25706 3415 25740
rect 3450 25706 3484 25740
rect 3519 25706 3553 25740
rect 3588 25706 3622 25740
rect 3657 25706 3691 25740
rect 3726 25706 3760 25740
rect 3795 25706 3829 25740
rect 3864 25706 3898 25740
rect 3933 25706 3967 25740
rect 4002 25706 4036 25740
rect 4071 25706 4105 25740
rect 4140 25706 4174 25740
rect 4208 25706 4242 25740
rect 4276 25706 4310 25740
rect 4344 25706 4378 25740
rect 4412 25706 4446 25740
rect 4480 25706 4514 25740
rect 4548 25706 4582 25740
rect 4616 25706 4650 25740
rect 4684 25706 4718 25740
rect 4752 25706 4786 25740
rect 4820 25706 4854 25740
rect 4888 25706 4922 25740
rect 4956 25706 4990 25740
rect 5024 25706 5058 25740
rect 5092 25706 5126 25740
rect 5160 25706 5194 25740
rect 5228 25706 5262 25740
rect 5296 25706 5330 25740
rect 5364 25706 5398 25740
rect 5432 25706 5466 25740
rect 5500 25706 5534 25740
rect 5568 25706 5602 25740
rect 5636 25706 5670 25740
rect 5704 25706 5738 25740
rect 5772 25706 5806 25740
rect 5840 25706 5874 25740
rect 5908 25706 5942 25740
rect 5976 25706 6010 25740
rect 6044 25706 6078 25740
rect 6112 25706 6146 25740
rect 6180 25706 6214 25740
rect 6248 25706 6282 25740
rect 6316 25706 6350 25740
rect 6384 25706 6418 25740
rect 6452 25706 6486 25740
rect 6520 25706 6554 25740
rect 6588 25706 6622 25740
rect 6656 25706 6690 25740
rect 6724 25706 6758 25740
rect 6792 25706 6826 25740
rect 6860 25706 6894 25740
rect 6928 25706 6962 25740
rect 6996 25706 7030 25740
rect 7064 25706 7098 25740
rect 7132 25706 7166 25740
rect 7200 25706 7234 25740
rect 7268 25706 7302 25740
rect 7336 25706 7370 25740
rect 7404 25706 7438 25740
rect 7472 25706 7506 25740
rect 7540 25706 7574 25740
rect 7608 25706 7642 25740
rect 7676 25706 7710 25740
rect 7744 25706 7778 25740
rect 7812 25706 7846 25740
rect 7880 25706 7914 25740
rect 7948 25706 7982 25740
rect 8016 25706 8050 25740
rect 8084 25706 8118 25740
rect 8152 25706 8186 25740
rect 8220 25706 8254 25740
rect 8288 25706 8322 25740
rect 8356 25706 8390 25740
rect 8424 25706 8458 25740
rect 8492 25706 8526 25740
rect 8560 25706 8594 25740
rect 8628 25706 8662 25740
rect 8696 25706 8730 25740
rect 8764 25706 8798 25740
rect 8832 25706 8866 25740
rect 8900 25706 8934 25740
rect 8968 25706 9002 25740
rect 9036 25706 9070 25740
rect 9104 25706 9138 25740
rect 9172 25706 9206 25740
rect 9240 25706 9274 25740
rect 9308 25706 9342 25740
rect 9376 25706 9410 25740
rect 9444 25706 9478 25740
rect 9512 25706 9546 25740
rect 9580 25706 9614 25740
rect 9648 25706 9682 25740
rect 9716 25706 9750 25740
rect 9784 25706 9818 25740
rect 9852 25706 9886 25740
rect 9920 25706 9954 25740
rect 9988 25706 10022 25740
rect 10056 25706 10090 25740
rect 10124 25706 10158 25740
rect 10192 25706 10226 25740
rect 10260 25706 10294 25740
rect 10328 25706 10362 25740
rect 10396 25706 10430 25740
rect 10464 25706 10498 25740
rect 10532 25706 10566 25740
rect 10600 25706 10634 25740
rect 10668 25706 10702 25740
rect 10736 25706 10770 25740
rect 10804 25706 10838 25740
rect 10872 25706 10906 25740
rect 10940 25706 10974 25740
rect 11008 25706 11042 25740
rect 11076 25706 11110 25740
rect 11144 25706 11178 25740
rect 11212 25706 11246 25740
rect 11280 25706 11314 25740
rect 11348 25706 11382 25740
rect 11416 25706 11450 25740
rect 11484 25706 11518 25740
rect 11552 25706 11586 25740
rect 11620 25706 11654 25740
rect 11688 25706 11722 25740
rect 11756 25706 11790 25740
rect 11824 25706 11858 25740
rect 11892 25706 11926 25740
rect 11960 25706 11994 25740
rect 12028 25706 12062 25740
rect 12096 25706 12130 25740
rect 12164 25706 12198 25740
rect 12232 25706 12266 25740
rect 12300 25706 12334 25740
rect 12368 25706 12402 25740
rect 12436 25706 12470 25740
rect 12504 25706 12538 25740
rect 12572 25706 12606 25740
rect 12640 25706 12674 25740
rect 12708 25706 12742 25740
rect 12776 25706 12810 25740
rect 12844 25706 12878 25740
rect 12912 25706 12946 25740
rect 12980 25706 13014 25740
rect 13048 25706 13082 25740
rect 13116 25706 13150 25740
rect 13184 25706 13218 25740
rect 13252 25706 13286 25740
rect 13320 25706 13354 25740
rect 13388 25706 13422 25740
rect 13456 25706 13490 25740
rect 13524 25706 13558 25740
rect 13592 25706 13626 25740
rect 13660 25706 13694 25740
rect 13728 25706 13762 25740
rect 13796 25706 13830 25740
rect 13864 25706 13898 25740
rect 13932 25706 13966 25740
rect 14000 25706 14034 25740
rect 14068 25706 14102 25740
rect 14136 25706 14170 25740
rect 14204 25706 14238 25740
rect 14272 25706 14306 25740
rect 14340 25706 14374 25740
rect 14408 25706 14442 25740
rect 14476 25706 14510 25740
rect 14544 25706 14578 25740
rect 14612 25706 14646 25740
rect 14680 25706 14714 25740
rect 14748 25706 14782 25740
rect 14816 25706 14850 25740
rect 14884 25706 14918 25740
rect 69 25634 103 25668
rect 138 25634 172 25668
rect 207 25634 241 25668
rect 276 25634 310 25668
rect 345 25634 379 25668
rect 414 25634 448 25668
rect 483 25634 517 25668
rect 552 25634 586 25668
rect 621 25634 655 25668
rect 690 25634 724 25668
rect 759 25634 793 25668
rect 828 25634 862 25668
rect 897 25634 931 25668
rect 966 25634 1000 25668
rect 1035 25634 1069 25668
rect 1104 25634 1138 25668
rect 1173 25634 1207 25668
rect 1242 25634 1276 25668
rect 1311 25634 1345 25668
rect 1380 25634 1414 25668
rect 1449 25634 1483 25668
rect 1518 25634 1552 25668
rect 1587 25634 1621 25668
rect 1656 25634 1690 25668
rect 1725 25634 1759 25668
rect 1794 25634 1828 25668
rect 1863 25634 1897 25668
rect 1932 25634 1966 25668
rect 2001 25634 2035 25668
rect 2070 25634 2104 25668
rect 2139 25634 2173 25668
rect 2208 25634 2242 25668
rect 2277 25634 2311 25668
rect 2346 25634 2380 25668
rect 2415 25634 2449 25668
rect 2484 25634 2518 25668
rect 2553 25634 2587 25668
rect 2622 25634 2656 25668
rect 2691 25634 2725 25668
rect 2760 25634 2794 25668
rect 2829 25634 2863 25668
rect 2898 25634 2932 25668
rect 2967 25634 3001 25668
rect 3036 25634 3070 25668
rect 3105 25634 3139 25668
rect 3174 25634 3208 25668
rect 3243 25634 3277 25668
rect 3312 25634 3346 25668
rect 3381 25634 3415 25668
rect 3450 25634 3484 25668
rect 3519 25634 3553 25668
rect 3588 25634 3622 25668
rect 3657 25634 3691 25668
rect 3726 25634 3760 25668
rect 3795 25634 3829 25668
rect 3864 25634 3898 25668
rect 3933 25634 3967 25668
rect 4002 25634 4036 25668
rect 4071 25634 4105 25668
rect 4140 25634 4174 25668
rect 4208 25634 4242 25668
rect 4276 25634 4310 25668
rect 4344 25634 4378 25668
rect 4412 25634 4446 25668
rect 4480 25634 4514 25668
rect 4548 25634 4582 25668
rect 4616 25634 4650 25668
rect 4684 25634 4718 25668
rect 4752 25634 4786 25668
rect 4820 25634 4854 25668
rect 4888 25634 4922 25668
rect 4956 25634 4990 25668
rect 5024 25634 5058 25668
rect 5092 25634 5126 25668
rect 5160 25634 5194 25668
rect 5228 25634 5262 25668
rect 5296 25634 5330 25668
rect 5364 25634 5398 25668
rect 5432 25634 5466 25668
rect 5500 25634 5534 25668
rect 5568 25634 5602 25668
rect 5636 25634 5670 25668
rect 5704 25634 5738 25668
rect 5772 25634 5806 25668
rect 5840 25634 5874 25668
rect 5908 25634 5942 25668
rect 5976 25634 6010 25668
rect 6044 25634 6078 25668
rect 6112 25634 6146 25668
rect 6180 25634 6214 25668
rect 6248 25634 6282 25668
rect 6316 25634 6350 25668
rect 6384 25634 6418 25668
rect 6452 25634 6486 25668
rect 6520 25634 6554 25668
rect 6588 25634 6622 25668
rect 6656 25634 6690 25668
rect 6724 25634 6758 25668
rect 6792 25634 6826 25668
rect 6860 25634 6894 25668
rect 6928 25634 6962 25668
rect 6996 25634 7030 25668
rect 7064 25634 7098 25668
rect 7132 25634 7166 25668
rect 7200 25634 7234 25668
rect 7268 25634 7302 25668
rect 7336 25634 7370 25668
rect 7404 25634 7438 25668
rect 7472 25634 7506 25668
rect 7540 25634 7574 25668
rect 7608 25634 7642 25668
rect 7676 25634 7710 25668
rect 7744 25634 7778 25668
rect 7812 25634 7846 25668
rect 7880 25634 7914 25668
rect 7948 25634 7982 25668
rect 8016 25634 8050 25668
rect 8084 25634 8118 25668
rect 8152 25634 8186 25668
rect 8220 25634 8254 25668
rect 8288 25634 8322 25668
rect 8356 25634 8390 25668
rect 8424 25634 8458 25668
rect 8492 25634 8526 25668
rect 8560 25634 8594 25668
rect 8628 25634 8662 25668
rect 8696 25634 8730 25668
rect 8764 25634 8798 25668
rect 8832 25634 8866 25668
rect 8900 25634 8934 25668
rect 8968 25634 9002 25668
rect 9036 25634 9070 25668
rect 9104 25634 9138 25668
rect 9172 25634 9206 25668
rect 9240 25634 9274 25668
rect 9308 25634 9342 25668
rect 9376 25634 9410 25668
rect 9444 25634 9478 25668
rect 9512 25634 9546 25668
rect 9580 25634 9614 25668
rect 9648 25634 9682 25668
rect 9716 25634 9750 25668
rect 9784 25634 9818 25668
rect 9852 25634 9886 25668
rect 9920 25634 9954 25668
rect 9988 25634 10022 25668
rect 10056 25634 10090 25668
rect 10124 25634 10158 25668
rect 10192 25634 10226 25668
rect 10260 25634 10294 25668
rect 10328 25634 10362 25668
rect 10396 25634 10430 25668
rect 10464 25634 10498 25668
rect 10532 25634 10566 25668
rect 10600 25634 10634 25668
rect 10668 25634 10702 25668
rect 10736 25634 10770 25668
rect 10804 25634 10838 25668
rect 10872 25634 10906 25668
rect 10940 25634 10974 25668
rect 11008 25634 11042 25668
rect 11076 25634 11110 25668
rect 11144 25634 11178 25668
rect 11212 25634 11246 25668
rect 11280 25634 11314 25668
rect 11348 25634 11382 25668
rect 11416 25634 11450 25668
rect 11484 25634 11518 25668
rect 11552 25634 11586 25668
rect 11620 25634 11654 25668
rect 11688 25634 11722 25668
rect 11756 25634 11790 25668
rect 11824 25634 11858 25668
rect 11892 25634 11926 25668
rect 11960 25634 11994 25668
rect 12028 25634 12062 25668
rect 12096 25634 12130 25668
rect 12164 25634 12198 25668
rect 12232 25634 12266 25668
rect 12300 25634 12334 25668
rect 12368 25634 12402 25668
rect 12436 25634 12470 25668
rect 12504 25634 12538 25668
rect 12572 25634 12606 25668
rect 12640 25634 12674 25668
rect 12708 25634 12742 25668
rect 12776 25634 12810 25668
rect 12844 25634 12878 25668
rect 12912 25634 12946 25668
rect 12980 25634 13014 25668
rect 13048 25634 13082 25668
rect 13116 25634 13150 25668
rect 13184 25634 13218 25668
rect 13252 25634 13286 25668
rect 13320 25634 13354 25668
rect 13388 25634 13422 25668
rect 13456 25634 13490 25668
rect 13524 25634 13558 25668
rect 13592 25634 13626 25668
rect 13660 25634 13694 25668
rect 13728 25634 13762 25668
rect 13796 25634 13830 25668
rect 13864 25634 13898 25668
rect 13932 25634 13966 25668
rect 14000 25634 14034 25668
rect 14068 25634 14102 25668
rect 14136 25634 14170 25668
rect 14204 25634 14238 25668
rect 14272 25634 14306 25668
rect 14340 25634 14374 25668
rect 14408 25634 14442 25668
rect 14476 25634 14510 25668
rect 14544 25634 14578 25668
rect 14612 25634 14646 25668
rect 14680 25634 14714 25668
rect 14748 25634 14782 25668
rect 14816 25634 14850 25668
rect 14884 25634 14918 25668
<< locali >>
rect 59 28283 14882 28289
rect 59 28249 121 28283
rect 155 28249 190 28283
rect 224 28249 259 28283
rect 293 28249 328 28283
rect 362 28249 397 28283
rect 431 28249 466 28283
rect 500 28249 535 28283
rect 569 28249 604 28283
rect 638 28249 673 28283
rect 707 28249 742 28283
rect 776 28249 811 28283
rect 845 28249 880 28283
rect 914 28249 949 28283
rect 983 28249 1018 28283
rect 1052 28249 1087 28283
rect 1121 28249 1156 28283
rect 59 28215 1156 28249
rect 59 28181 121 28215
rect 155 28181 190 28215
rect 224 28181 259 28215
rect 293 28181 328 28215
rect 362 28181 397 28215
rect 431 28181 466 28215
rect 500 28181 535 28215
rect 569 28181 604 28215
rect 638 28181 673 28215
rect 707 28181 742 28215
rect 776 28181 811 28215
rect 845 28181 880 28215
rect 914 28181 949 28215
rect 983 28181 1018 28215
rect 1052 28181 1087 28215
rect 1121 28181 1156 28215
rect 59 28147 1156 28181
rect 59 28122 121 28147
rect 155 28122 190 28147
rect 224 28122 259 28147
rect 59 28088 112 28122
rect 155 28113 185 28122
rect 224 28113 258 28122
rect 293 28113 328 28147
rect 362 28122 397 28147
rect 431 28122 466 28147
rect 500 28122 535 28147
rect 569 28122 604 28147
rect 638 28122 673 28147
rect 707 28122 742 28147
rect 776 28122 811 28147
rect 845 28122 880 28147
rect 365 28113 397 28122
rect 438 28113 466 28122
rect 511 28113 535 28122
rect 584 28113 604 28122
rect 657 28113 673 28122
rect 730 28113 742 28122
rect 803 28113 811 28122
rect 876 28113 880 28122
rect 914 28122 949 28147
rect 914 28113 915 28122
rect 146 28088 185 28113
rect 219 28088 258 28113
rect 292 28088 331 28113
rect 365 28088 404 28113
rect 438 28088 477 28113
rect 511 28088 550 28113
rect 584 28088 623 28113
rect 657 28088 696 28113
rect 730 28088 769 28113
rect 803 28088 842 28113
rect 876 28088 915 28113
rect 983 28122 1018 28147
rect 1052 28122 1087 28147
rect 1121 28122 1156 28147
rect 983 28113 988 28122
rect 1052 28113 1061 28122
rect 1121 28113 1134 28122
rect 949 28088 988 28113
rect 1022 28088 1061 28113
rect 1095 28088 1134 28113
rect 59 28079 1156 28088
rect 59 28045 121 28079
rect 155 28045 190 28079
rect 224 28045 259 28079
rect 293 28045 328 28079
rect 362 28045 397 28079
rect 431 28045 466 28079
rect 500 28045 535 28079
rect 569 28045 604 28079
rect 638 28045 673 28079
rect 707 28045 742 28079
rect 776 28045 811 28079
rect 845 28045 880 28079
rect 914 28045 949 28079
rect 983 28045 1018 28079
rect 1052 28045 1087 28079
rect 1121 28045 1156 28079
rect 59 28040 1156 28045
rect 59 28006 112 28040
rect 146 28011 185 28040
rect 219 28011 258 28040
rect 292 28011 331 28040
rect 365 28011 404 28040
rect 438 28011 477 28040
rect 511 28011 550 28040
rect 584 28011 623 28040
rect 657 28011 696 28040
rect 730 28011 769 28040
rect 803 28011 842 28040
rect 876 28011 915 28040
rect 155 28006 185 28011
rect 224 28006 258 28011
rect 59 27977 121 28006
rect 155 27977 190 28006
rect 224 27977 259 28006
rect 293 27977 328 28011
rect 365 28006 397 28011
rect 438 28006 466 28011
rect 511 28006 535 28011
rect 584 28006 604 28011
rect 657 28006 673 28011
rect 730 28006 742 28011
rect 803 28006 811 28011
rect 876 28006 880 28011
rect 362 27977 397 28006
rect 431 27977 466 28006
rect 500 27977 535 28006
rect 569 27977 604 28006
rect 638 27977 673 28006
rect 707 27977 742 28006
rect 776 27977 811 28006
rect 845 27977 880 28006
rect 914 28006 915 28011
rect 949 28011 988 28040
rect 1022 28011 1061 28040
rect 1095 28011 1134 28040
rect 914 27977 949 28006
rect 983 28006 988 28011
rect 1052 28006 1061 28011
rect 1121 28006 1134 28011
rect 983 27977 1018 28006
rect 1052 27977 1087 28006
rect 1121 27977 1156 28006
rect 59 27958 1156 27977
rect 59 27924 112 27958
rect 146 27943 185 27958
rect 219 27943 258 27958
rect 292 27943 331 27958
rect 365 27943 404 27958
rect 438 27943 477 27958
rect 511 27943 550 27958
rect 584 27943 623 27958
rect 657 27943 696 27958
rect 730 27943 769 27958
rect 803 27943 842 27958
rect 876 27943 915 27958
rect 155 27924 185 27943
rect 224 27924 258 27943
rect 59 27909 121 27924
rect 155 27909 190 27924
rect 224 27909 259 27924
rect 293 27909 328 27943
rect 365 27924 397 27943
rect 438 27924 466 27943
rect 511 27924 535 27943
rect 584 27924 604 27943
rect 657 27924 673 27943
rect 730 27924 742 27943
rect 803 27924 811 27943
rect 876 27924 880 27943
rect 362 27909 397 27924
rect 431 27909 466 27924
rect 500 27909 535 27924
rect 569 27909 604 27924
rect 638 27909 673 27924
rect 707 27909 742 27924
rect 776 27909 811 27924
rect 845 27909 880 27924
rect 914 27924 915 27943
rect 949 27943 988 27958
rect 1022 27943 1061 27958
rect 1095 27943 1134 27958
rect 914 27909 949 27924
rect 983 27924 988 27943
rect 1052 27924 1061 27943
rect 1121 27924 1134 27943
rect 983 27909 1018 27924
rect 1052 27909 1087 27924
rect 1121 27909 1156 27924
rect 59 27876 1156 27909
rect 59 27842 112 27876
rect 146 27875 185 27876
rect 219 27875 258 27876
rect 292 27875 331 27876
rect 365 27875 404 27876
rect 438 27875 477 27876
rect 511 27875 550 27876
rect 584 27875 623 27876
rect 657 27875 696 27876
rect 730 27875 769 27876
rect 803 27875 842 27876
rect 876 27875 915 27876
rect 155 27842 185 27875
rect 224 27842 258 27875
rect 59 27841 121 27842
rect 155 27841 190 27842
rect 224 27841 259 27842
rect 293 27841 328 27875
rect 365 27842 397 27875
rect 438 27842 466 27875
rect 511 27842 535 27875
rect 584 27842 604 27875
rect 657 27842 673 27875
rect 730 27842 742 27875
rect 803 27842 811 27875
rect 876 27842 880 27875
rect 362 27841 397 27842
rect 431 27841 466 27842
rect 500 27841 535 27842
rect 569 27841 604 27842
rect 638 27841 673 27842
rect 707 27841 742 27842
rect 776 27841 811 27842
rect 845 27841 880 27842
rect 914 27842 915 27875
rect 949 27875 988 27876
rect 1022 27875 1061 27876
rect 1095 27875 1134 27876
rect 914 27841 949 27842
rect 983 27842 988 27875
rect 1052 27842 1061 27875
rect 1121 27842 1134 27875
rect 983 27841 1018 27842
rect 1052 27841 1087 27842
rect 1121 27841 1156 27842
rect 59 27807 1156 27841
rect 59 27794 121 27807
rect 155 27794 190 27807
rect 224 27794 259 27807
rect 59 27760 112 27794
rect 155 27773 185 27794
rect 224 27773 258 27794
rect 293 27773 328 27807
rect 362 27794 397 27807
rect 431 27794 466 27807
rect 500 27794 535 27807
rect 569 27794 604 27807
rect 638 27794 673 27807
rect 707 27794 742 27807
rect 776 27794 811 27807
rect 845 27794 880 27807
rect 365 27773 397 27794
rect 438 27773 466 27794
rect 511 27773 535 27794
rect 584 27773 604 27794
rect 657 27773 673 27794
rect 730 27773 742 27794
rect 803 27773 811 27794
rect 876 27773 880 27794
rect 914 27794 949 27807
rect 914 27773 915 27794
rect 146 27760 185 27773
rect 219 27760 258 27773
rect 292 27760 331 27773
rect 365 27760 404 27773
rect 438 27760 477 27773
rect 511 27760 550 27773
rect 584 27760 623 27773
rect 657 27760 696 27773
rect 730 27760 769 27773
rect 803 27760 842 27773
rect 876 27760 915 27773
rect 983 27794 1018 27807
rect 1052 27794 1087 27807
rect 1121 27794 1156 27807
rect 983 27773 988 27794
rect 1052 27773 1061 27794
rect 1121 27773 1134 27794
rect 949 27760 988 27773
rect 1022 27760 1061 27773
rect 1095 27760 1134 27773
rect 59 27739 1156 27760
rect 59 27712 121 27739
rect 155 27712 190 27739
rect 224 27712 259 27739
rect 59 27678 112 27712
rect 155 27705 185 27712
rect 224 27705 258 27712
rect 293 27705 328 27739
rect 362 27712 397 27739
rect 431 27712 466 27739
rect 500 27712 535 27739
rect 569 27712 604 27739
rect 638 27712 673 27739
rect 707 27712 742 27739
rect 776 27712 811 27739
rect 845 27712 880 27739
rect 365 27705 397 27712
rect 438 27705 466 27712
rect 511 27705 535 27712
rect 584 27705 604 27712
rect 657 27705 673 27712
rect 730 27705 742 27712
rect 803 27705 811 27712
rect 876 27705 880 27712
rect 914 27712 949 27739
rect 914 27705 915 27712
rect 146 27678 185 27705
rect 219 27678 258 27705
rect 292 27678 331 27705
rect 365 27678 404 27705
rect 438 27678 477 27705
rect 511 27678 550 27705
rect 584 27678 623 27705
rect 657 27678 696 27705
rect 730 27678 769 27705
rect 803 27678 842 27705
rect 876 27678 915 27705
rect 983 27712 1018 27739
rect 1052 27712 1087 27739
rect 1121 27712 1156 27739
rect 983 27705 988 27712
rect 1052 27705 1061 27712
rect 1121 27705 1134 27712
rect 949 27678 988 27705
rect 1022 27678 1061 27705
rect 1095 27678 1134 27705
rect 59 27671 1156 27678
rect 59 27637 121 27671
rect 155 27637 190 27671
rect 224 27637 259 27671
rect 293 27637 328 27671
rect 362 27637 397 27671
rect 431 27637 466 27671
rect 500 27637 535 27671
rect 569 27637 604 27671
rect 638 27637 673 27671
rect 707 27637 742 27671
rect 776 27637 811 27671
rect 845 27637 880 27671
rect 914 27637 949 27671
rect 983 27637 1018 27671
rect 1052 27637 1087 27671
rect 1121 27637 1156 27671
rect 59 27603 1156 27637
rect 59 27569 121 27603
rect 155 27569 190 27603
rect 224 27569 259 27603
rect 293 27569 328 27603
rect 362 27569 397 27603
rect 431 27569 466 27603
rect 500 27569 535 27603
rect 569 27569 604 27603
rect 638 27569 673 27603
rect 707 27569 742 27603
rect 776 27569 811 27603
rect 845 27569 880 27603
rect 914 27569 949 27603
rect 983 27569 1018 27603
rect 1052 27569 1087 27603
rect 1121 27569 1156 27603
rect 14858 27569 14882 28283
rect 59 27563 14882 27569
rect 57 27376 14962 27410
rect 57 27342 83 27376
rect 117 27342 152 27376
rect 186 27355 221 27376
rect 255 27355 290 27376
rect 324 27355 359 27376
rect 393 27355 428 27376
rect 462 27355 497 27376
rect 197 27342 221 27355
rect 271 27342 290 27355
rect 345 27342 359 27355
rect 419 27342 428 27355
rect 493 27342 497 27355
rect 531 27355 566 27376
rect 600 27355 635 27376
rect 669 27355 704 27376
rect 738 27355 773 27376
rect 807 27362 842 27376
rect 876 27362 911 27376
rect 945 27362 980 27376
rect 1014 27362 1049 27376
rect 1083 27362 1118 27376
rect 531 27342 533 27355
rect 600 27342 606 27355
rect 669 27342 679 27355
rect 738 27342 752 27355
rect 807 27342 827 27362
rect 876 27342 899 27362
rect 945 27342 971 27362
rect 1014 27342 1043 27362
rect 1083 27342 1115 27362
rect 1152 27342 1187 27376
rect 1221 27342 1256 27376
rect 1290 27362 1325 27376
rect 1359 27362 1394 27376
rect 1428 27362 1463 27376
rect 1497 27362 1532 27376
rect 1566 27362 1601 27376
rect 1635 27362 1670 27376
rect 1704 27362 1739 27376
rect 1773 27362 1808 27376
rect 1842 27362 1877 27376
rect 1911 27362 1946 27376
rect 1293 27342 1325 27362
rect 1365 27342 1394 27362
rect 1437 27342 1463 27362
rect 1509 27342 1532 27362
rect 1581 27342 1601 27362
rect 1653 27342 1670 27362
rect 1725 27342 1739 27362
rect 1798 27342 1808 27362
rect 1871 27342 1877 27362
rect 1944 27342 1946 27362
rect 1980 27362 2014 27376
rect 2048 27362 2082 27376
rect 1980 27342 1983 27362
rect 2048 27342 2056 27362
rect 2116 27355 2150 27376
rect 2116 27342 2142 27355
rect 2184 27342 2218 27376
rect 2252 27355 2286 27376
rect 2320 27355 2354 27376
rect 2388 27355 2422 27376
rect 2255 27342 2286 27355
rect 2334 27342 2354 27355
rect 2413 27342 2422 27355
rect 2456 27355 2490 27376
rect 2524 27355 2558 27376
rect 2592 27355 2626 27376
rect 2660 27355 2694 27376
rect 2456 27342 2458 27355
rect 2524 27342 2536 27355
rect 2592 27342 2614 27355
rect 2660 27342 2692 27355
rect 2728 27342 2762 27376
rect 2796 27372 14962 27376
rect 2796 27355 2848 27372
rect 57 27321 163 27342
rect 197 27321 237 27342
rect 271 27321 311 27342
rect 345 27321 385 27342
rect 419 27321 459 27342
rect 493 27321 533 27342
rect 567 27321 606 27342
rect 640 27321 679 27342
rect 713 27321 752 27342
rect 786 27328 827 27342
rect 861 27328 899 27342
rect 933 27328 971 27342
rect 1005 27328 1043 27342
rect 1077 27328 1115 27342
rect 1149 27328 1187 27342
rect 1221 27328 1259 27342
rect 1293 27328 1331 27342
rect 1365 27328 1403 27342
rect 1437 27328 1475 27342
rect 1509 27328 1547 27342
rect 1581 27328 1619 27342
rect 1653 27328 1691 27342
rect 1725 27328 1764 27342
rect 1798 27328 1837 27342
rect 1871 27328 1910 27342
rect 1944 27328 1983 27342
rect 2017 27328 2056 27342
rect 2090 27328 2142 27342
rect 786 27321 2142 27328
rect 2176 27321 2221 27342
rect 2255 27321 2300 27342
rect 2334 27321 2379 27342
rect 2413 27321 2458 27342
rect 2492 27321 2536 27342
rect 2570 27321 2614 27342
rect 2648 27321 2692 27342
rect 2726 27321 2770 27342
rect 2804 27321 2848 27355
rect 2882 27338 2916 27372
rect 2950 27355 2984 27372
rect 2960 27338 2984 27355
rect 3018 27338 3052 27372
rect 3086 27338 3120 27372
rect 3154 27338 3188 27372
rect 3222 27338 3256 27372
rect 3290 27338 3324 27372
rect 3358 27338 3392 27372
rect 3426 27338 3460 27372
rect 3494 27362 3528 27372
rect 3562 27362 3596 27372
rect 3630 27362 3664 27372
rect 3698 27362 3732 27372
rect 3766 27362 3800 27372
rect 3834 27362 3868 27372
rect 3499 27338 3528 27362
rect 3572 27338 3596 27362
rect 3645 27338 3664 27362
rect 3718 27338 3732 27362
rect 3791 27338 3800 27362
rect 3864 27338 3868 27362
rect 3902 27362 3936 27372
rect 3970 27362 4004 27372
rect 4038 27362 4072 27372
rect 4106 27362 4140 27372
rect 4174 27362 4208 27372
rect 4242 27362 4276 27372
rect 4310 27362 4344 27372
rect 4378 27362 4412 27372
rect 3902 27338 3903 27362
rect 3970 27338 3976 27362
rect 4038 27338 4049 27362
rect 4106 27338 4122 27362
rect 4174 27338 4194 27362
rect 4242 27338 4266 27362
rect 4310 27338 4338 27362
rect 4378 27338 4410 27362
rect 4446 27338 4480 27372
rect 4514 27362 4548 27372
rect 4582 27362 4616 27372
rect 4650 27362 4684 27372
rect 4718 27362 4752 27372
rect 4786 27362 4820 27372
rect 4854 27362 4888 27372
rect 4922 27362 4956 27372
rect 4990 27362 5024 27372
rect 4516 27338 4548 27362
rect 4588 27338 4616 27362
rect 4660 27338 4684 27362
rect 4732 27338 4752 27362
rect 4804 27338 4820 27362
rect 4876 27338 4888 27362
rect 4948 27338 4956 27362
rect 5020 27338 5024 27362
rect 5058 27362 5092 27372
rect 2882 27321 2926 27338
rect 2960 27328 3392 27338
rect 3426 27328 3465 27338
rect 3499 27328 3538 27338
rect 3572 27328 3611 27338
rect 3645 27328 3684 27338
rect 3718 27328 3757 27338
rect 3791 27328 3830 27338
rect 3864 27328 3903 27338
rect 3937 27328 3976 27338
rect 4010 27328 4049 27338
rect 4083 27328 4122 27338
rect 4156 27328 4194 27338
rect 4228 27328 4266 27338
rect 4300 27328 4338 27338
rect 4372 27328 4410 27338
rect 4444 27328 4482 27338
rect 4516 27328 4554 27338
rect 4588 27328 4626 27338
rect 4660 27328 4698 27338
rect 4732 27328 4770 27338
rect 4804 27328 4842 27338
rect 4876 27328 4914 27338
rect 4948 27328 4986 27338
rect 5020 27328 5058 27338
rect 5126 27362 5160 27372
rect 5194 27362 5228 27372
rect 5262 27362 5296 27372
rect 5330 27362 5364 27372
rect 5398 27362 5432 27372
rect 5466 27362 5500 27372
rect 5534 27362 5568 27372
rect 5602 27362 5636 27372
rect 5126 27338 5130 27362
rect 5194 27338 5202 27362
rect 5262 27338 5274 27362
rect 5330 27338 5346 27362
rect 5398 27338 5418 27362
rect 5466 27338 5490 27362
rect 5534 27338 5562 27362
rect 5602 27338 5634 27362
rect 5670 27338 5704 27372
rect 5738 27362 5772 27372
rect 5806 27362 5840 27372
rect 5874 27362 5908 27372
rect 5942 27362 5976 27372
rect 6010 27362 6044 27372
rect 6078 27362 6112 27372
rect 6146 27362 6180 27372
rect 6214 27362 6248 27372
rect 5740 27338 5772 27362
rect 5812 27338 5840 27362
rect 5884 27338 5908 27362
rect 5956 27338 5976 27362
rect 6028 27338 6044 27362
rect 6100 27338 6112 27362
rect 6172 27338 6180 27362
rect 6244 27338 6248 27362
rect 6282 27362 6316 27372
rect 5092 27328 5130 27338
rect 5164 27328 5202 27338
rect 5236 27328 5274 27338
rect 5308 27328 5346 27338
rect 5380 27328 5418 27338
rect 5452 27328 5490 27338
rect 5524 27328 5562 27338
rect 5596 27328 5634 27338
rect 5668 27328 5706 27338
rect 5740 27328 5778 27338
rect 5812 27328 5850 27338
rect 5884 27328 5922 27338
rect 5956 27328 5994 27338
rect 6028 27328 6066 27338
rect 6100 27328 6138 27338
rect 6172 27328 6210 27338
rect 6244 27328 6282 27338
rect 6350 27362 6384 27372
rect 6418 27362 6452 27372
rect 6486 27362 6520 27372
rect 6554 27362 6588 27372
rect 6622 27362 6656 27372
rect 6690 27362 6724 27372
rect 6758 27362 6792 27372
rect 6826 27362 6860 27372
rect 6350 27338 6354 27362
rect 6418 27338 6426 27362
rect 6486 27338 6498 27362
rect 6554 27338 6570 27362
rect 6622 27338 6642 27362
rect 6690 27338 6714 27362
rect 6758 27338 6786 27362
rect 6826 27338 6858 27362
rect 6894 27338 6928 27372
rect 6962 27362 6996 27372
rect 7030 27362 7064 27372
rect 7098 27362 7132 27372
rect 7166 27362 7200 27372
rect 7234 27362 7268 27372
rect 7302 27362 7336 27372
rect 7370 27362 7404 27372
rect 7438 27362 7472 27372
rect 6964 27338 6996 27362
rect 7036 27338 7064 27362
rect 7108 27338 7132 27362
rect 7180 27338 7200 27362
rect 7252 27338 7268 27362
rect 7324 27338 7336 27362
rect 7396 27338 7404 27362
rect 7468 27338 7472 27362
rect 7506 27362 7540 27372
rect 6316 27328 6354 27338
rect 6388 27328 6426 27338
rect 6460 27328 6498 27338
rect 6532 27328 6570 27338
rect 6604 27328 6642 27338
rect 6676 27328 6714 27338
rect 6748 27328 6786 27338
rect 6820 27328 6858 27338
rect 6892 27328 6930 27338
rect 6964 27328 7002 27338
rect 7036 27328 7074 27338
rect 7108 27328 7146 27338
rect 7180 27328 7218 27338
rect 7252 27328 7290 27338
rect 7324 27328 7362 27338
rect 7396 27328 7434 27338
rect 7468 27328 7506 27338
rect 7574 27362 7608 27372
rect 7642 27362 7676 27372
rect 7710 27362 7744 27372
rect 7778 27362 7812 27372
rect 7846 27362 7880 27372
rect 7914 27362 7948 27372
rect 7982 27362 8016 27372
rect 8050 27362 8084 27372
rect 7574 27338 7578 27362
rect 7642 27338 7650 27362
rect 7710 27338 7722 27362
rect 7778 27338 7794 27362
rect 7846 27338 7866 27362
rect 7914 27338 7938 27362
rect 7982 27338 8010 27362
rect 8050 27338 8082 27362
rect 8118 27338 8152 27372
rect 8186 27362 8220 27372
rect 8254 27362 8288 27372
rect 8322 27362 8356 27372
rect 8390 27362 8424 27372
rect 8458 27362 8492 27372
rect 8526 27362 8560 27372
rect 8594 27362 8628 27372
rect 8662 27362 8696 27372
rect 8188 27338 8220 27362
rect 8260 27338 8288 27362
rect 8332 27338 8356 27362
rect 8404 27338 8424 27362
rect 8476 27338 8492 27362
rect 8548 27338 8560 27362
rect 8620 27338 8628 27362
rect 8692 27338 8696 27362
rect 8730 27362 8764 27372
rect 7540 27328 7578 27338
rect 7612 27328 7650 27338
rect 7684 27328 7722 27338
rect 7756 27328 7794 27338
rect 7828 27328 7866 27338
rect 7900 27328 7938 27338
rect 7972 27328 8010 27338
rect 8044 27328 8082 27338
rect 8116 27328 8154 27338
rect 8188 27328 8226 27338
rect 8260 27328 8298 27338
rect 8332 27328 8370 27338
rect 8404 27328 8442 27338
rect 8476 27328 8514 27338
rect 8548 27328 8586 27338
rect 8620 27328 8658 27338
rect 8692 27328 8730 27338
rect 8798 27362 8832 27372
rect 8866 27362 8900 27372
rect 8934 27362 8968 27372
rect 9002 27362 9036 27372
rect 9070 27362 9104 27372
rect 9138 27362 9172 27372
rect 9206 27362 9240 27372
rect 9274 27362 9308 27372
rect 8798 27338 8802 27362
rect 8866 27338 8874 27362
rect 8934 27338 8946 27362
rect 9002 27338 9018 27362
rect 9070 27338 9090 27362
rect 9138 27338 9162 27362
rect 9206 27338 9234 27362
rect 9274 27338 9306 27362
rect 9342 27338 9376 27372
rect 9410 27362 9444 27372
rect 9478 27362 9512 27372
rect 9546 27362 9580 27372
rect 9614 27362 9648 27372
rect 9682 27362 9716 27372
rect 9750 27362 9784 27372
rect 9818 27362 9852 27372
rect 9886 27362 9920 27372
rect 9412 27338 9444 27362
rect 9484 27338 9512 27362
rect 9556 27338 9580 27362
rect 9628 27338 9648 27362
rect 9700 27338 9716 27362
rect 9772 27338 9784 27362
rect 9844 27338 9852 27362
rect 9916 27338 9920 27362
rect 9954 27362 9988 27372
rect 8764 27328 8802 27338
rect 8836 27328 8874 27338
rect 8908 27328 8946 27338
rect 8980 27328 9018 27338
rect 9052 27328 9090 27338
rect 9124 27328 9162 27338
rect 9196 27328 9234 27338
rect 9268 27328 9306 27338
rect 9340 27328 9378 27338
rect 9412 27328 9450 27338
rect 9484 27328 9522 27338
rect 9556 27328 9594 27338
rect 9628 27328 9666 27338
rect 9700 27328 9738 27338
rect 9772 27328 9810 27338
rect 9844 27328 9882 27338
rect 9916 27328 9954 27338
rect 10022 27362 10056 27372
rect 10090 27362 10124 27372
rect 10158 27362 10192 27372
rect 10226 27362 10260 27372
rect 10294 27362 10328 27372
rect 10362 27362 10396 27372
rect 10430 27362 10464 27372
rect 10498 27362 10532 27372
rect 10022 27338 10026 27362
rect 10090 27338 10098 27362
rect 10158 27338 10170 27362
rect 10226 27338 10242 27362
rect 10294 27338 10314 27362
rect 10362 27338 10386 27362
rect 10430 27338 10458 27362
rect 10498 27338 10530 27362
rect 10566 27338 10600 27372
rect 10634 27362 10668 27372
rect 10702 27362 10736 27372
rect 10770 27362 10804 27372
rect 10838 27362 10872 27372
rect 10906 27362 10940 27372
rect 10974 27362 11008 27372
rect 11042 27362 11076 27372
rect 11110 27362 11144 27372
rect 10636 27338 10668 27362
rect 10708 27338 10736 27362
rect 10780 27338 10804 27362
rect 10852 27338 10872 27362
rect 10924 27338 10940 27362
rect 10996 27338 11008 27362
rect 11068 27338 11076 27362
rect 11140 27338 11144 27362
rect 11178 27362 11212 27372
rect 9988 27328 10026 27338
rect 10060 27328 10098 27338
rect 10132 27328 10170 27338
rect 10204 27328 10242 27338
rect 10276 27328 10314 27338
rect 10348 27328 10386 27338
rect 10420 27328 10458 27338
rect 10492 27328 10530 27338
rect 10564 27328 10602 27338
rect 10636 27328 10674 27338
rect 10708 27328 10746 27338
rect 10780 27328 10818 27338
rect 10852 27328 10890 27338
rect 10924 27328 10962 27338
rect 10996 27328 11034 27338
rect 11068 27328 11106 27338
rect 11140 27328 11178 27338
rect 11246 27362 11280 27372
rect 11314 27362 11348 27372
rect 11382 27362 11416 27372
rect 11450 27362 11484 27372
rect 11518 27362 11552 27372
rect 11586 27362 11620 27372
rect 11654 27362 11688 27372
rect 11722 27362 11756 27372
rect 11246 27338 11250 27362
rect 11314 27338 11322 27362
rect 11382 27338 11394 27362
rect 11450 27338 11466 27362
rect 11518 27338 11538 27362
rect 11586 27338 11610 27362
rect 11654 27338 11682 27362
rect 11722 27338 11754 27362
rect 11790 27338 11824 27372
rect 11858 27362 11892 27372
rect 11926 27362 11960 27372
rect 11994 27362 12028 27372
rect 12062 27362 12096 27372
rect 12130 27362 12164 27372
rect 12198 27362 12232 27372
rect 12266 27362 12300 27372
rect 12334 27362 12368 27372
rect 11860 27338 11892 27362
rect 11932 27338 11960 27362
rect 12004 27338 12028 27362
rect 12076 27338 12096 27362
rect 12148 27338 12164 27362
rect 12220 27338 12232 27362
rect 12292 27338 12300 27362
rect 12364 27338 12368 27362
rect 12402 27362 12436 27372
rect 11212 27328 11250 27338
rect 11284 27328 11322 27338
rect 11356 27328 11394 27338
rect 11428 27328 11466 27338
rect 11500 27328 11538 27338
rect 11572 27328 11610 27338
rect 11644 27328 11682 27338
rect 11716 27328 11754 27338
rect 11788 27328 11826 27338
rect 11860 27328 11898 27338
rect 11932 27328 11970 27338
rect 12004 27328 12042 27338
rect 12076 27328 12114 27338
rect 12148 27328 12186 27338
rect 12220 27328 12258 27338
rect 12292 27328 12330 27338
rect 12364 27328 12402 27338
rect 12470 27362 12504 27372
rect 12538 27362 12572 27372
rect 12606 27362 12640 27372
rect 12674 27362 12708 27372
rect 12742 27362 12776 27372
rect 12810 27362 12844 27372
rect 12878 27362 12912 27372
rect 12946 27362 12980 27372
rect 12470 27338 12474 27362
rect 12538 27338 12546 27362
rect 12606 27338 12618 27362
rect 12674 27338 12690 27362
rect 12742 27338 12762 27362
rect 12810 27338 12834 27362
rect 12878 27338 12906 27362
rect 12946 27338 12978 27362
rect 13014 27338 13048 27372
rect 13082 27362 13116 27372
rect 13150 27362 13184 27372
rect 13218 27362 13252 27372
rect 13286 27362 13320 27372
rect 13354 27362 13388 27372
rect 13422 27362 13456 27372
rect 13490 27362 13524 27372
rect 13558 27362 13592 27372
rect 13084 27338 13116 27362
rect 13156 27338 13184 27362
rect 13228 27338 13252 27362
rect 13300 27338 13320 27362
rect 13372 27338 13388 27362
rect 13444 27338 13456 27362
rect 13516 27338 13524 27362
rect 13588 27338 13592 27362
rect 13626 27362 13660 27372
rect 12436 27328 12474 27338
rect 12508 27328 12546 27338
rect 12580 27328 12618 27338
rect 12652 27328 12690 27338
rect 12724 27328 12762 27338
rect 12796 27328 12834 27338
rect 12868 27328 12906 27338
rect 12940 27328 12978 27338
rect 13012 27328 13050 27338
rect 13084 27328 13122 27338
rect 13156 27328 13194 27338
rect 13228 27328 13266 27338
rect 13300 27328 13338 27338
rect 13372 27328 13410 27338
rect 13444 27328 13482 27338
rect 13516 27328 13554 27338
rect 13588 27328 13626 27338
rect 13694 27362 13728 27372
rect 13762 27362 13796 27372
rect 13830 27362 13864 27372
rect 13898 27362 13932 27372
rect 13966 27362 14000 27372
rect 14034 27362 14068 27372
rect 14102 27362 14136 27372
rect 14170 27362 14204 27372
rect 13694 27338 13698 27362
rect 13762 27338 13770 27362
rect 13830 27338 13842 27362
rect 13898 27338 13914 27362
rect 13966 27338 13986 27362
rect 14034 27338 14058 27362
rect 14102 27338 14130 27362
rect 14170 27338 14202 27362
rect 14238 27338 14272 27372
rect 14306 27362 14340 27372
rect 14374 27362 14408 27372
rect 14442 27362 14476 27372
rect 14510 27362 14544 27372
rect 14578 27362 14612 27372
rect 14646 27362 14680 27372
rect 14714 27362 14748 27372
rect 14782 27362 14816 27372
rect 14308 27338 14340 27362
rect 14380 27338 14408 27362
rect 14452 27338 14476 27362
rect 14524 27338 14544 27362
rect 14596 27338 14612 27362
rect 14668 27338 14680 27362
rect 14740 27338 14748 27362
rect 14812 27338 14816 27362
rect 14850 27362 14884 27372
rect 13660 27328 13698 27338
rect 13732 27328 13770 27338
rect 13804 27328 13842 27338
rect 13876 27328 13914 27338
rect 13948 27328 13986 27338
rect 14020 27328 14058 27338
rect 14092 27328 14130 27338
rect 14164 27328 14202 27338
rect 14236 27328 14274 27338
rect 14308 27328 14346 27338
rect 14380 27328 14418 27338
rect 14452 27328 14490 27338
rect 14524 27328 14562 27338
rect 14596 27328 14634 27338
rect 14668 27328 14706 27338
rect 14740 27328 14778 27338
rect 14812 27328 14850 27338
rect 14918 27338 14962 27372
rect 14884 27328 14962 27338
rect 2960 27321 14962 27328
rect 57 27302 14962 27321
rect 57 27268 83 27302
rect 117 27268 152 27302
rect 186 27268 221 27302
rect 255 27268 290 27302
rect 324 27268 359 27302
rect 393 27268 428 27302
rect 462 27268 497 27302
rect 531 27268 566 27302
rect 600 27268 635 27302
rect 669 27268 704 27302
rect 738 27268 773 27302
rect 807 27268 842 27302
rect 876 27268 911 27302
rect 945 27268 980 27302
rect 1014 27268 1049 27302
rect 1083 27268 1118 27302
rect 1152 27268 1187 27302
rect 1221 27268 1256 27302
rect 1290 27268 1325 27302
rect 1359 27268 1394 27302
rect 1428 27268 1463 27302
rect 1497 27268 1532 27302
rect 1566 27268 1601 27302
rect 1635 27268 1670 27302
rect 1704 27268 1739 27302
rect 1773 27268 1808 27302
rect 1842 27268 1877 27302
rect 1911 27268 1946 27302
rect 1980 27268 2014 27302
rect 2048 27268 2082 27302
rect 2116 27268 2150 27302
rect 2184 27268 2218 27302
rect 2252 27268 2286 27302
rect 2320 27268 2354 27302
rect 2388 27268 2422 27302
rect 2456 27268 2490 27302
rect 2524 27268 2558 27302
rect 2592 27268 2626 27302
rect 2660 27268 2694 27302
rect 2728 27268 2762 27302
rect 2796 27268 2848 27302
rect 2882 27268 2916 27302
rect 2950 27268 2984 27302
rect 3018 27268 3052 27302
rect 3086 27268 3120 27302
rect 3154 27268 3188 27302
rect 3222 27268 3256 27302
rect 3290 27268 3324 27302
rect 3358 27268 3392 27302
rect 3426 27268 3460 27302
rect 3494 27268 3528 27302
rect 3562 27268 3596 27302
rect 3630 27268 3664 27302
rect 3698 27268 3732 27302
rect 3766 27268 3800 27302
rect 3834 27268 3868 27302
rect 3902 27268 3936 27302
rect 3970 27268 4004 27302
rect 4038 27268 4072 27302
rect 4106 27268 4140 27302
rect 4174 27268 4208 27302
rect 4242 27268 4276 27302
rect 4310 27268 4344 27302
rect 4378 27268 4412 27302
rect 4446 27268 4480 27302
rect 4514 27268 4548 27302
rect 4582 27268 4616 27302
rect 4650 27268 4684 27302
rect 4718 27268 4752 27302
rect 4786 27268 4820 27302
rect 4854 27268 4888 27302
rect 4922 27268 4956 27302
rect 4990 27268 5024 27302
rect 5058 27268 5092 27302
rect 5126 27268 5160 27302
rect 5194 27268 5228 27302
rect 5262 27268 5296 27302
rect 5330 27268 5364 27302
rect 5398 27268 5432 27302
rect 5466 27268 5500 27302
rect 5534 27268 5568 27302
rect 5602 27268 5636 27302
rect 5670 27268 5704 27302
rect 5738 27268 5772 27302
rect 5806 27268 5840 27302
rect 5874 27268 5908 27302
rect 5942 27268 5976 27302
rect 6010 27268 6044 27302
rect 6078 27268 6112 27302
rect 6146 27268 6180 27302
rect 6214 27268 6248 27302
rect 6282 27268 6316 27302
rect 6350 27268 6384 27302
rect 6418 27268 6452 27302
rect 6486 27268 6520 27302
rect 6554 27268 6588 27302
rect 6622 27268 6656 27302
rect 6690 27268 6724 27302
rect 6758 27268 6792 27302
rect 6826 27268 6860 27302
rect 6894 27268 6928 27302
rect 6962 27268 6996 27302
rect 7030 27268 7064 27302
rect 7098 27268 7132 27302
rect 7166 27268 7200 27302
rect 7234 27268 7268 27302
rect 7302 27268 7336 27302
rect 7370 27268 7404 27302
rect 7438 27268 7472 27302
rect 7506 27268 7540 27302
rect 7574 27268 7608 27302
rect 7642 27268 7676 27302
rect 7710 27268 7744 27302
rect 7778 27268 7812 27302
rect 7846 27268 7880 27302
rect 7914 27268 7948 27302
rect 7982 27268 8016 27302
rect 8050 27268 8084 27302
rect 8118 27268 8152 27302
rect 8186 27268 8220 27302
rect 8254 27268 8288 27302
rect 8322 27268 8356 27302
rect 8390 27268 8424 27302
rect 8458 27268 8492 27302
rect 8526 27268 8560 27302
rect 8594 27268 8628 27302
rect 8662 27268 8696 27302
rect 8730 27268 8764 27302
rect 8798 27268 8832 27302
rect 8866 27268 8900 27302
rect 8934 27268 8968 27302
rect 9002 27268 9036 27302
rect 9070 27268 9104 27302
rect 9138 27268 9172 27302
rect 9206 27268 9240 27302
rect 9274 27268 9308 27302
rect 9342 27268 9376 27302
rect 9410 27268 9444 27302
rect 9478 27268 9512 27302
rect 9546 27268 9580 27302
rect 9614 27268 9648 27302
rect 9682 27268 9716 27302
rect 9750 27268 9784 27302
rect 9818 27268 9852 27302
rect 9886 27268 9920 27302
rect 9954 27268 9988 27302
rect 10022 27268 10056 27302
rect 10090 27268 10124 27302
rect 10158 27268 10192 27302
rect 10226 27268 10260 27302
rect 10294 27268 10328 27302
rect 10362 27268 10396 27302
rect 10430 27268 10464 27302
rect 10498 27268 10532 27302
rect 10566 27268 10600 27302
rect 10634 27268 10668 27302
rect 10702 27268 10736 27302
rect 10770 27268 10804 27302
rect 10838 27268 10872 27302
rect 10906 27268 10940 27302
rect 10974 27268 11008 27302
rect 11042 27268 11076 27302
rect 11110 27268 11144 27302
rect 11178 27268 11212 27302
rect 11246 27268 11280 27302
rect 11314 27268 11348 27302
rect 11382 27268 11416 27302
rect 11450 27268 11484 27302
rect 11518 27268 11552 27302
rect 11586 27268 11620 27302
rect 11654 27268 11688 27302
rect 11722 27268 11756 27302
rect 11790 27268 11824 27302
rect 11858 27268 11892 27302
rect 11926 27268 11960 27302
rect 11994 27268 12028 27302
rect 12062 27268 12096 27302
rect 12130 27268 12164 27302
rect 12198 27268 12232 27302
rect 12266 27268 12300 27302
rect 12334 27268 12368 27302
rect 12402 27268 12436 27302
rect 12470 27268 12504 27302
rect 12538 27268 12572 27302
rect 12606 27268 12640 27302
rect 12674 27268 12708 27302
rect 12742 27268 12776 27302
rect 12810 27268 12844 27302
rect 12878 27268 12912 27302
rect 12946 27268 12980 27302
rect 13014 27268 13048 27302
rect 13082 27268 13116 27302
rect 13150 27268 13184 27302
rect 13218 27268 13252 27302
rect 13286 27268 13320 27302
rect 13354 27268 13388 27302
rect 13422 27268 13456 27302
rect 13490 27268 13524 27302
rect 13558 27268 13592 27302
rect 13626 27268 13660 27302
rect 13694 27268 13728 27302
rect 13762 27268 13796 27302
rect 13830 27268 13864 27302
rect 13898 27268 13932 27302
rect 13966 27268 14000 27302
rect 14034 27268 14068 27302
rect 14102 27268 14136 27302
rect 14170 27268 14204 27302
rect 14238 27268 14272 27302
rect 14306 27268 14340 27302
rect 14374 27268 14408 27302
rect 14442 27268 14476 27302
rect 14510 27268 14544 27302
rect 14578 27268 14612 27302
rect 14646 27268 14680 27302
rect 14714 27268 14748 27302
rect 14782 27268 14816 27302
rect 14850 27268 14884 27302
rect 14918 27268 14962 27302
rect 57 27238 14962 27268
rect 57 27228 827 27238
rect 861 27228 899 27238
rect 933 27228 971 27238
rect 1005 27228 1043 27238
rect 1077 27228 1115 27238
rect 1149 27228 1187 27238
rect 1221 27228 1259 27238
rect 1293 27228 1331 27238
rect 1365 27228 1403 27238
rect 1437 27228 1475 27238
rect 1509 27228 1547 27238
rect 1581 27228 1619 27238
rect 1653 27228 1691 27238
rect 1725 27228 1764 27238
rect 1798 27228 1837 27238
rect 1871 27228 1910 27238
rect 1944 27228 1983 27238
rect 2017 27228 2056 27238
rect 2090 27232 3392 27238
rect 3426 27232 3465 27238
rect 3499 27232 3538 27238
rect 3572 27232 3611 27238
rect 3645 27232 3684 27238
rect 3718 27232 3757 27238
rect 3791 27232 3830 27238
rect 3864 27232 3903 27238
rect 3937 27232 3976 27238
rect 4010 27232 4049 27238
rect 4083 27232 4122 27238
rect 4156 27232 4194 27238
rect 4228 27232 4266 27238
rect 4300 27232 4338 27238
rect 4372 27232 4410 27238
rect 4444 27232 4482 27238
rect 4516 27232 4554 27238
rect 4588 27232 4626 27238
rect 4660 27232 4698 27238
rect 4732 27232 4770 27238
rect 4804 27232 4842 27238
rect 4876 27232 4914 27238
rect 4948 27232 4986 27238
rect 5020 27232 5058 27238
rect 2090 27228 2848 27232
rect 57 27194 83 27228
rect 117 27194 152 27228
rect 186 27194 221 27228
rect 255 27194 290 27228
rect 324 27194 359 27228
rect 393 27194 428 27228
rect 462 27194 497 27228
rect 531 27194 566 27228
rect 600 27194 635 27228
rect 669 27194 704 27228
rect 738 27194 773 27228
rect 807 27204 827 27228
rect 876 27204 899 27228
rect 945 27204 971 27228
rect 1014 27204 1043 27228
rect 1083 27204 1115 27228
rect 807 27194 842 27204
rect 876 27194 911 27204
rect 945 27194 980 27204
rect 1014 27194 1049 27204
rect 1083 27194 1118 27204
rect 1152 27194 1187 27228
rect 1221 27194 1256 27228
rect 1293 27204 1325 27228
rect 1365 27204 1394 27228
rect 1437 27204 1463 27228
rect 1509 27204 1532 27228
rect 1581 27204 1601 27228
rect 1653 27204 1670 27228
rect 1725 27204 1739 27228
rect 1798 27204 1808 27228
rect 1871 27204 1877 27228
rect 1944 27204 1946 27228
rect 1290 27194 1325 27204
rect 1359 27194 1394 27204
rect 1428 27194 1463 27204
rect 1497 27194 1532 27204
rect 1566 27194 1601 27204
rect 1635 27194 1670 27204
rect 1704 27194 1739 27204
rect 1773 27194 1808 27204
rect 1842 27194 1877 27204
rect 1911 27194 1946 27204
rect 1980 27204 1983 27228
rect 2048 27204 2056 27228
rect 1980 27194 2014 27204
rect 2048 27194 2082 27204
rect 2116 27194 2150 27228
rect 2184 27194 2218 27228
rect 2252 27194 2286 27228
rect 2320 27194 2354 27228
rect 2388 27194 2422 27228
rect 2456 27194 2490 27228
rect 2524 27194 2558 27228
rect 2592 27194 2626 27228
rect 2660 27194 2694 27228
rect 2728 27194 2762 27228
rect 2796 27198 2848 27228
rect 2882 27198 2916 27232
rect 2950 27198 2984 27232
rect 3018 27198 3052 27232
rect 3086 27198 3120 27232
rect 3154 27198 3188 27232
rect 3222 27198 3256 27232
rect 3290 27198 3324 27232
rect 3358 27198 3392 27232
rect 3426 27198 3460 27232
rect 3499 27204 3528 27232
rect 3572 27204 3596 27232
rect 3645 27204 3664 27232
rect 3718 27204 3732 27232
rect 3791 27204 3800 27232
rect 3864 27204 3868 27232
rect 3494 27198 3528 27204
rect 3562 27198 3596 27204
rect 3630 27198 3664 27204
rect 3698 27198 3732 27204
rect 3766 27198 3800 27204
rect 3834 27198 3868 27204
rect 3902 27204 3903 27232
rect 3970 27204 3976 27232
rect 4038 27204 4049 27232
rect 4106 27204 4122 27232
rect 4174 27204 4194 27232
rect 4242 27204 4266 27232
rect 4310 27204 4338 27232
rect 4378 27204 4410 27232
rect 3902 27198 3936 27204
rect 3970 27198 4004 27204
rect 4038 27198 4072 27204
rect 4106 27198 4140 27204
rect 4174 27198 4208 27204
rect 4242 27198 4276 27204
rect 4310 27198 4344 27204
rect 4378 27198 4412 27204
rect 4446 27198 4480 27232
rect 4516 27204 4548 27232
rect 4588 27204 4616 27232
rect 4660 27204 4684 27232
rect 4732 27204 4752 27232
rect 4804 27204 4820 27232
rect 4876 27204 4888 27232
rect 4948 27204 4956 27232
rect 5020 27204 5024 27232
rect 4514 27198 4548 27204
rect 4582 27198 4616 27204
rect 4650 27198 4684 27204
rect 4718 27198 4752 27204
rect 4786 27198 4820 27204
rect 4854 27198 4888 27204
rect 4922 27198 4956 27204
rect 4990 27198 5024 27204
rect 5092 27232 5130 27238
rect 5164 27232 5202 27238
rect 5236 27232 5274 27238
rect 5308 27232 5346 27238
rect 5380 27232 5418 27238
rect 5452 27232 5490 27238
rect 5524 27232 5562 27238
rect 5596 27232 5634 27238
rect 5668 27232 5706 27238
rect 5740 27232 5778 27238
rect 5812 27232 5850 27238
rect 5884 27232 5922 27238
rect 5956 27232 5994 27238
rect 6028 27232 6066 27238
rect 6100 27232 6138 27238
rect 6172 27232 6210 27238
rect 6244 27232 6282 27238
rect 5058 27198 5092 27204
rect 5126 27204 5130 27232
rect 5194 27204 5202 27232
rect 5262 27204 5274 27232
rect 5330 27204 5346 27232
rect 5398 27204 5418 27232
rect 5466 27204 5490 27232
rect 5534 27204 5562 27232
rect 5602 27204 5634 27232
rect 5126 27198 5160 27204
rect 5194 27198 5228 27204
rect 5262 27198 5296 27204
rect 5330 27198 5364 27204
rect 5398 27198 5432 27204
rect 5466 27198 5500 27204
rect 5534 27198 5568 27204
rect 5602 27198 5636 27204
rect 5670 27198 5704 27232
rect 5740 27204 5772 27232
rect 5812 27204 5840 27232
rect 5884 27204 5908 27232
rect 5956 27204 5976 27232
rect 6028 27204 6044 27232
rect 6100 27204 6112 27232
rect 6172 27204 6180 27232
rect 6244 27204 6248 27232
rect 5738 27198 5772 27204
rect 5806 27198 5840 27204
rect 5874 27198 5908 27204
rect 5942 27198 5976 27204
rect 6010 27198 6044 27204
rect 6078 27198 6112 27204
rect 6146 27198 6180 27204
rect 6214 27198 6248 27204
rect 6316 27232 6354 27238
rect 6388 27232 6426 27238
rect 6460 27232 6498 27238
rect 6532 27232 6570 27238
rect 6604 27232 6642 27238
rect 6676 27232 6714 27238
rect 6748 27232 6786 27238
rect 6820 27232 6858 27238
rect 6892 27232 6930 27238
rect 6964 27232 7002 27238
rect 7036 27232 7074 27238
rect 7108 27232 7146 27238
rect 7180 27232 7218 27238
rect 7252 27232 7290 27238
rect 7324 27232 7362 27238
rect 7396 27232 7434 27238
rect 7468 27232 7506 27238
rect 6282 27198 6316 27204
rect 6350 27204 6354 27232
rect 6418 27204 6426 27232
rect 6486 27204 6498 27232
rect 6554 27204 6570 27232
rect 6622 27204 6642 27232
rect 6690 27204 6714 27232
rect 6758 27204 6786 27232
rect 6826 27204 6858 27232
rect 6350 27198 6384 27204
rect 6418 27198 6452 27204
rect 6486 27198 6520 27204
rect 6554 27198 6588 27204
rect 6622 27198 6656 27204
rect 6690 27198 6724 27204
rect 6758 27198 6792 27204
rect 6826 27198 6860 27204
rect 6894 27198 6928 27232
rect 6964 27204 6996 27232
rect 7036 27204 7064 27232
rect 7108 27204 7132 27232
rect 7180 27204 7200 27232
rect 7252 27204 7268 27232
rect 7324 27204 7336 27232
rect 7396 27204 7404 27232
rect 7468 27204 7472 27232
rect 6962 27198 6996 27204
rect 7030 27198 7064 27204
rect 7098 27198 7132 27204
rect 7166 27198 7200 27204
rect 7234 27198 7268 27204
rect 7302 27198 7336 27204
rect 7370 27198 7404 27204
rect 7438 27198 7472 27204
rect 7540 27232 7578 27238
rect 7612 27232 7650 27238
rect 7684 27232 7722 27238
rect 7756 27232 7794 27238
rect 7828 27232 7866 27238
rect 7900 27232 7938 27238
rect 7972 27232 8010 27238
rect 8044 27232 8082 27238
rect 8116 27232 8154 27238
rect 8188 27232 8226 27238
rect 8260 27232 8298 27238
rect 8332 27232 8370 27238
rect 8404 27232 8442 27238
rect 8476 27232 8514 27238
rect 8548 27232 8586 27238
rect 8620 27232 8658 27238
rect 8692 27232 8730 27238
rect 7506 27198 7540 27204
rect 7574 27204 7578 27232
rect 7642 27204 7650 27232
rect 7710 27204 7722 27232
rect 7778 27204 7794 27232
rect 7846 27204 7866 27232
rect 7914 27204 7938 27232
rect 7982 27204 8010 27232
rect 8050 27204 8082 27232
rect 7574 27198 7608 27204
rect 7642 27198 7676 27204
rect 7710 27198 7744 27204
rect 7778 27198 7812 27204
rect 7846 27198 7880 27204
rect 7914 27198 7948 27204
rect 7982 27198 8016 27204
rect 8050 27198 8084 27204
rect 8118 27198 8152 27232
rect 8188 27204 8220 27232
rect 8260 27204 8288 27232
rect 8332 27204 8356 27232
rect 8404 27204 8424 27232
rect 8476 27204 8492 27232
rect 8548 27204 8560 27232
rect 8620 27204 8628 27232
rect 8692 27204 8696 27232
rect 8186 27198 8220 27204
rect 8254 27198 8288 27204
rect 8322 27198 8356 27204
rect 8390 27198 8424 27204
rect 8458 27198 8492 27204
rect 8526 27198 8560 27204
rect 8594 27198 8628 27204
rect 8662 27198 8696 27204
rect 8764 27232 8802 27238
rect 8836 27232 8874 27238
rect 8908 27232 8946 27238
rect 8980 27232 9018 27238
rect 9052 27232 9090 27238
rect 9124 27232 9162 27238
rect 9196 27232 9234 27238
rect 9268 27232 9306 27238
rect 9340 27232 9378 27238
rect 9412 27232 9450 27238
rect 9484 27232 9522 27238
rect 9556 27232 9594 27238
rect 9628 27232 9666 27238
rect 9700 27232 9738 27238
rect 9772 27232 9810 27238
rect 9844 27232 9882 27238
rect 9916 27232 9954 27238
rect 8730 27198 8764 27204
rect 8798 27204 8802 27232
rect 8866 27204 8874 27232
rect 8934 27204 8946 27232
rect 9002 27204 9018 27232
rect 9070 27204 9090 27232
rect 9138 27204 9162 27232
rect 9206 27204 9234 27232
rect 9274 27204 9306 27232
rect 8798 27198 8832 27204
rect 8866 27198 8900 27204
rect 8934 27198 8968 27204
rect 9002 27198 9036 27204
rect 9070 27198 9104 27204
rect 9138 27198 9172 27204
rect 9206 27198 9240 27204
rect 9274 27198 9308 27204
rect 9342 27198 9376 27232
rect 9412 27204 9444 27232
rect 9484 27204 9512 27232
rect 9556 27204 9580 27232
rect 9628 27204 9648 27232
rect 9700 27204 9716 27232
rect 9772 27204 9784 27232
rect 9844 27204 9852 27232
rect 9916 27204 9920 27232
rect 9410 27198 9444 27204
rect 9478 27198 9512 27204
rect 9546 27198 9580 27204
rect 9614 27198 9648 27204
rect 9682 27198 9716 27204
rect 9750 27198 9784 27204
rect 9818 27198 9852 27204
rect 9886 27198 9920 27204
rect 9988 27232 10026 27238
rect 10060 27232 10098 27238
rect 10132 27232 10170 27238
rect 10204 27232 10242 27238
rect 10276 27232 10314 27238
rect 10348 27232 10386 27238
rect 10420 27232 10458 27238
rect 10492 27232 10530 27238
rect 10564 27232 10602 27238
rect 10636 27232 10674 27238
rect 10708 27232 10746 27238
rect 10780 27232 10818 27238
rect 10852 27232 10890 27238
rect 10924 27232 10962 27238
rect 10996 27232 11034 27238
rect 11068 27232 11106 27238
rect 11140 27232 11178 27238
rect 9954 27198 9988 27204
rect 10022 27204 10026 27232
rect 10090 27204 10098 27232
rect 10158 27204 10170 27232
rect 10226 27204 10242 27232
rect 10294 27204 10314 27232
rect 10362 27204 10386 27232
rect 10430 27204 10458 27232
rect 10498 27204 10530 27232
rect 10022 27198 10056 27204
rect 10090 27198 10124 27204
rect 10158 27198 10192 27204
rect 10226 27198 10260 27204
rect 10294 27198 10328 27204
rect 10362 27198 10396 27204
rect 10430 27198 10464 27204
rect 10498 27198 10532 27204
rect 10566 27198 10600 27232
rect 10636 27204 10668 27232
rect 10708 27204 10736 27232
rect 10780 27204 10804 27232
rect 10852 27204 10872 27232
rect 10924 27204 10940 27232
rect 10996 27204 11008 27232
rect 11068 27204 11076 27232
rect 11140 27204 11144 27232
rect 10634 27198 10668 27204
rect 10702 27198 10736 27204
rect 10770 27198 10804 27204
rect 10838 27198 10872 27204
rect 10906 27198 10940 27204
rect 10974 27198 11008 27204
rect 11042 27198 11076 27204
rect 11110 27198 11144 27204
rect 11212 27232 11250 27238
rect 11284 27232 11322 27238
rect 11356 27232 11394 27238
rect 11428 27232 11466 27238
rect 11500 27232 11538 27238
rect 11572 27232 11610 27238
rect 11644 27232 11682 27238
rect 11716 27232 11754 27238
rect 11788 27232 11826 27238
rect 11860 27232 11898 27238
rect 11932 27232 11970 27238
rect 12004 27232 12042 27238
rect 12076 27232 12114 27238
rect 12148 27232 12186 27238
rect 12220 27232 12258 27238
rect 12292 27232 12330 27238
rect 12364 27232 12402 27238
rect 11178 27198 11212 27204
rect 11246 27204 11250 27232
rect 11314 27204 11322 27232
rect 11382 27204 11394 27232
rect 11450 27204 11466 27232
rect 11518 27204 11538 27232
rect 11586 27204 11610 27232
rect 11654 27204 11682 27232
rect 11722 27204 11754 27232
rect 11246 27198 11280 27204
rect 11314 27198 11348 27204
rect 11382 27198 11416 27204
rect 11450 27198 11484 27204
rect 11518 27198 11552 27204
rect 11586 27198 11620 27204
rect 11654 27198 11688 27204
rect 11722 27198 11756 27204
rect 11790 27198 11824 27232
rect 11860 27204 11892 27232
rect 11932 27204 11960 27232
rect 12004 27204 12028 27232
rect 12076 27204 12096 27232
rect 12148 27204 12164 27232
rect 12220 27204 12232 27232
rect 12292 27204 12300 27232
rect 12364 27204 12368 27232
rect 11858 27198 11892 27204
rect 11926 27198 11960 27204
rect 11994 27198 12028 27204
rect 12062 27198 12096 27204
rect 12130 27198 12164 27204
rect 12198 27198 12232 27204
rect 12266 27198 12300 27204
rect 12334 27198 12368 27204
rect 12436 27232 12474 27238
rect 12508 27232 12546 27238
rect 12580 27232 12618 27238
rect 12652 27232 12690 27238
rect 12724 27232 12762 27238
rect 12796 27232 12834 27238
rect 12868 27232 12906 27238
rect 12940 27232 12978 27238
rect 13012 27232 13050 27238
rect 13084 27232 13122 27238
rect 13156 27232 13194 27238
rect 13228 27232 13266 27238
rect 13300 27232 13338 27238
rect 13372 27232 13410 27238
rect 13444 27232 13482 27238
rect 13516 27232 13554 27238
rect 13588 27232 13626 27238
rect 12402 27198 12436 27204
rect 12470 27204 12474 27232
rect 12538 27204 12546 27232
rect 12606 27204 12618 27232
rect 12674 27204 12690 27232
rect 12742 27204 12762 27232
rect 12810 27204 12834 27232
rect 12878 27204 12906 27232
rect 12946 27204 12978 27232
rect 12470 27198 12504 27204
rect 12538 27198 12572 27204
rect 12606 27198 12640 27204
rect 12674 27198 12708 27204
rect 12742 27198 12776 27204
rect 12810 27198 12844 27204
rect 12878 27198 12912 27204
rect 12946 27198 12980 27204
rect 13014 27198 13048 27232
rect 13084 27204 13116 27232
rect 13156 27204 13184 27232
rect 13228 27204 13252 27232
rect 13300 27204 13320 27232
rect 13372 27204 13388 27232
rect 13444 27204 13456 27232
rect 13516 27204 13524 27232
rect 13588 27204 13592 27232
rect 13082 27198 13116 27204
rect 13150 27198 13184 27204
rect 13218 27198 13252 27204
rect 13286 27198 13320 27204
rect 13354 27198 13388 27204
rect 13422 27198 13456 27204
rect 13490 27198 13524 27204
rect 13558 27198 13592 27204
rect 13660 27232 13698 27238
rect 13732 27232 13770 27238
rect 13804 27232 13842 27238
rect 13876 27232 13914 27238
rect 13948 27232 13986 27238
rect 14020 27232 14058 27238
rect 14092 27232 14130 27238
rect 14164 27232 14202 27238
rect 14236 27232 14274 27238
rect 14308 27232 14346 27238
rect 14380 27232 14418 27238
rect 14452 27232 14490 27238
rect 14524 27232 14562 27238
rect 14596 27232 14634 27238
rect 14668 27232 14706 27238
rect 14740 27232 14778 27238
rect 14812 27232 14850 27238
rect 13626 27198 13660 27204
rect 13694 27204 13698 27232
rect 13762 27204 13770 27232
rect 13830 27204 13842 27232
rect 13898 27204 13914 27232
rect 13966 27204 13986 27232
rect 14034 27204 14058 27232
rect 14102 27204 14130 27232
rect 14170 27204 14202 27232
rect 13694 27198 13728 27204
rect 13762 27198 13796 27204
rect 13830 27198 13864 27204
rect 13898 27198 13932 27204
rect 13966 27198 14000 27204
rect 14034 27198 14068 27204
rect 14102 27198 14136 27204
rect 14170 27198 14204 27204
rect 14238 27198 14272 27232
rect 14308 27204 14340 27232
rect 14380 27204 14408 27232
rect 14452 27204 14476 27232
rect 14524 27204 14544 27232
rect 14596 27204 14612 27232
rect 14668 27204 14680 27232
rect 14740 27204 14748 27232
rect 14812 27204 14816 27232
rect 14306 27198 14340 27204
rect 14374 27198 14408 27204
rect 14442 27198 14476 27204
rect 14510 27198 14544 27204
rect 14578 27198 14612 27204
rect 14646 27198 14680 27204
rect 14714 27198 14748 27204
rect 14782 27198 14816 27204
rect 14884 27232 14962 27238
rect 14850 27198 14884 27204
rect 14918 27198 14962 27232
rect 2796 27194 14962 27198
rect 57 27162 14962 27194
rect 57 27154 2848 27162
rect 57 27120 83 27154
rect 117 27120 152 27154
rect 186 27120 221 27154
rect 255 27120 290 27154
rect 324 27120 359 27154
rect 393 27120 428 27154
rect 462 27120 497 27154
rect 531 27120 566 27154
rect 600 27120 635 27154
rect 669 27120 704 27154
rect 738 27120 773 27154
rect 807 27120 842 27154
rect 876 27120 911 27154
rect 945 27120 980 27154
rect 1014 27120 1049 27154
rect 1083 27120 1118 27154
rect 1152 27120 1187 27154
rect 1221 27120 1256 27154
rect 1290 27120 1325 27154
rect 1359 27120 1394 27154
rect 1428 27120 1463 27154
rect 1497 27120 1532 27154
rect 1566 27120 1601 27154
rect 1635 27120 1670 27154
rect 1704 27120 1739 27154
rect 1773 27120 1808 27154
rect 1842 27120 1877 27154
rect 1911 27120 1946 27154
rect 1980 27120 2014 27154
rect 2048 27120 2082 27154
rect 2116 27120 2150 27154
rect 2184 27120 2218 27154
rect 2252 27120 2286 27154
rect 2320 27120 2354 27154
rect 2388 27120 2422 27154
rect 2456 27120 2490 27154
rect 2524 27120 2558 27154
rect 2592 27120 2626 27154
rect 2660 27120 2694 27154
rect 2728 27120 2762 27154
rect 2796 27128 2848 27154
rect 2882 27128 2916 27162
rect 2950 27128 2984 27162
rect 3018 27128 3052 27162
rect 3086 27128 3120 27162
rect 3154 27128 3188 27162
rect 3222 27128 3256 27162
rect 3290 27128 3324 27162
rect 3358 27128 3392 27162
rect 3426 27128 3460 27162
rect 3494 27128 3528 27162
rect 3562 27128 3596 27162
rect 3630 27128 3664 27162
rect 3698 27128 3732 27162
rect 3766 27128 3800 27162
rect 3834 27128 3868 27162
rect 3902 27128 3936 27162
rect 3970 27128 4004 27162
rect 4038 27128 4072 27162
rect 4106 27128 4140 27162
rect 4174 27128 4208 27162
rect 4242 27128 4276 27162
rect 4310 27128 4344 27162
rect 4378 27128 4412 27162
rect 4446 27128 4480 27162
rect 4514 27128 4548 27162
rect 4582 27128 4616 27162
rect 4650 27128 4684 27162
rect 4718 27128 4752 27162
rect 4786 27128 4820 27162
rect 4854 27128 4888 27162
rect 4922 27128 4956 27162
rect 4990 27128 5024 27162
rect 5058 27128 5092 27162
rect 5126 27128 5160 27162
rect 5194 27128 5228 27162
rect 5262 27128 5296 27162
rect 5330 27128 5364 27162
rect 5398 27128 5432 27162
rect 5466 27128 5500 27162
rect 5534 27128 5568 27162
rect 5602 27128 5636 27162
rect 5670 27128 5704 27162
rect 5738 27128 5772 27162
rect 5806 27128 5840 27162
rect 5874 27128 5908 27162
rect 5942 27128 5976 27162
rect 6010 27128 6044 27162
rect 6078 27128 6112 27162
rect 6146 27128 6180 27162
rect 6214 27128 6248 27162
rect 6282 27128 6316 27162
rect 6350 27128 6384 27162
rect 6418 27128 6452 27162
rect 6486 27128 6520 27162
rect 6554 27128 6588 27162
rect 6622 27128 6656 27162
rect 6690 27128 6724 27162
rect 6758 27128 6792 27162
rect 6826 27128 6860 27162
rect 6894 27128 6928 27162
rect 6962 27128 6996 27162
rect 7030 27128 7064 27162
rect 7098 27128 7132 27162
rect 7166 27128 7200 27162
rect 7234 27128 7268 27162
rect 7302 27128 7336 27162
rect 7370 27128 7404 27162
rect 7438 27128 7472 27162
rect 7506 27128 7540 27162
rect 7574 27128 7608 27162
rect 7642 27128 7676 27162
rect 7710 27128 7744 27162
rect 7778 27128 7812 27162
rect 7846 27128 7880 27162
rect 7914 27128 7948 27162
rect 7982 27128 8016 27162
rect 8050 27128 8084 27162
rect 8118 27128 8152 27162
rect 8186 27128 8220 27162
rect 8254 27128 8288 27162
rect 8322 27128 8356 27162
rect 8390 27128 8424 27162
rect 8458 27128 8492 27162
rect 8526 27128 8560 27162
rect 8594 27128 8628 27162
rect 8662 27128 8696 27162
rect 8730 27128 8764 27162
rect 8798 27128 8832 27162
rect 8866 27128 8900 27162
rect 8934 27128 8968 27162
rect 9002 27128 9036 27162
rect 9070 27128 9104 27162
rect 9138 27128 9172 27162
rect 9206 27128 9240 27162
rect 9274 27128 9308 27162
rect 9342 27128 9376 27162
rect 9410 27128 9444 27162
rect 9478 27128 9512 27162
rect 9546 27128 9580 27162
rect 9614 27128 9648 27162
rect 9682 27128 9716 27162
rect 9750 27128 9784 27162
rect 9818 27128 9852 27162
rect 9886 27128 9920 27162
rect 9954 27128 9988 27162
rect 10022 27128 10056 27162
rect 10090 27128 10124 27162
rect 10158 27128 10192 27162
rect 10226 27128 10260 27162
rect 10294 27128 10328 27162
rect 10362 27128 10396 27162
rect 10430 27128 10464 27162
rect 10498 27128 10532 27162
rect 10566 27128 10600 27162
rect 10634 27128 10668 27162
rect 10702 27128 10736 27162
rect 10770 27128 10804 27162
rect 10838 27128 10872 27162
rect 10906 27128 10940 27162
rect 10974 27128 11008 27162
rect 11042 27128 11076 27162
rect 11110 27128 11144 27162
rect 11178 27128 11212 27162
rect 11246 27128 11280 27162
rect 11314 27128 11348 27162
rect 11382 27128 11416 27162
rect 11450 27128 11484 27162
rect 11518 27128 11552 27162
rect 11586 27128 11620 27162
rect 11654 27128 11688 27162
rect 11722 27128 11756 27162
rect 11790 27128 11824 27162
rect 11858 27128 11892 27162
rect 11926 27128 11960 27162
rect 11994 27128 12028 27162
rect 12062 27128 12096 27162
rect 12130 27128 12164 27162
rect 12198 27128 12232 27162
rect 12266 27128 12300 27162
rect 12334 27128 12368 27162
rect 12402 27128 12436 27162
rect 12470 27128 12504 27162
rect 12538 27128 12572 27162
rect 12606 27128 12640 27162
rect 12674 27128 12708 27162
rect 12742 27128 12776 27162
rect 12810 27128 12844 27162
rect 12878 27128 12912 27162
rect 12946 27128 12980 27162
rect 13014 27128 13048 27162
rect 13082 27128 13116 27162
rect 13150 27128 13184 27162
rect 13218 27128 13252 27162
rect 13286 27128 13320 27162
rect 13354 27128 13388 27162
rect 13422 27128 13456 27162
rect 13490 27128 13524 27162
rect 13558 27128 13592 27162
rect 13626 27128 13660 27162
rect 13694 27128 13728 27162
rect 13762 27128 13796 27162
rect 13830 27128 13864 27162
rect 13898 27128 13932 27162
rect 13966 27128 14000 27162
rect 14034 27128 14068 27162
rect 14102 27128 14136 27162
rect 14170 27128 14204 27162
rect 14238 27128 14272 27162
rect 14306 27128 14340 27162
rect 14374 27128 14408 27162
rect 14442 27128 14476 27162
rect 14510 27128 14544 27162
rect 14578 27128 14612 27162
rect 14646 27128 14680 27162
rect 14714 27128 14748 27162
rect 14782 27128 14816 27162
rect 14850 27128 14884 27162
rect 14918 27128 14962 27162
rect 2796 27120 14962 27128
rect 57 27092 14962 27120
rect 57 27086 2848 27092
rect 49 26794 151 27086
rect 2822 27058 2848 27086
rect 2882 27058 2916 27092
rect 2950 27058 2984 27092
rect 3018 27058 3052 27092
rect 3086 27058 3120 27092
rect 3154 27058 3188 27092
rect 3222 27058 3256 27092
rect 3290 27058 3324 27092
rect 3358 27058 3392 27092
rect 3426 27058 3460 27092
rect 3494 27058 3528 27092
rect 3562 27058 3596 27092
rect 3630 27058 3664 27092
rect 3698 27058 3732 27092
rect 3766 27058 3800 27092
rect 3834 27058 3868 27092
rect 3902 27058 3936 27092
rect 3970 27058 4004 27092
rect 4038 27058 4072 27092
rect 4106 27058 4140 27092
rect 4174 27058 4208 27092
rect 4242 27058 4276 27092
rect 4310 27058 4344 27092
rect 4378 27058 4412 27092
rect 4446 27058 4480 27092
rect 4514 27058 4548 27092
rect 4582 27058 4616 27092
rect 4650 27058 4684 27092
rect 4718 27058 4752 27092
rect 4786 27058 4820 27092
rect 4854 27058 4888 27092
rect 4922 27058 4956 27092
rect 4990 27058 5024 27092
rect 5058 27058 5092 27092
rect 5126 27058 5160 27092
rect 5194 27058 5228 27092
rect 5262 27058 5296 27092
rect 5330 27058 5364 27092
rect 5398 27058 5432 27092
rect 5466 27058 5500 27092
rect 5534 27058 5568 27092
rect 5602 27058 5636 27092
rect 5670 27058 5704 27092
rect 5738 27058 5772 27092
rect 5806 27058 5840 27092
rect 5874 27058 5908 27092
rect 5942 27058 5976 27092
rect 6010 27058 6044 27092
rect 6078 27058 6112 27092
rect 6146 27058 6180 27092
rect 6214 27058 6248 27092
rect 6282 27058 6316 27092
rect 6350 27058 6384 27092
rect 6418 27058 6452 27092
rect 6486 27058 6520 27092
rect 6554 27058 6588 27092
rect 6622 27058 6656 27092
rect 6690 27058 6724 27092
rect 6758 27058 6792 27092
rect 6826 27058 6860 27092
rect 6894 27058 6928 27092
rect 6962 27058 6996 27092
rect 7030 27058 7064 27092
rect 7098 27058 7132 27092
rect 7166 27058 7200 27092
rect 7234 27058 7268 27092
rect 7302 27058 7336 27092
rect 7370 27058 7404 27092
rect 7438 27058 7472 27092
rect 7506 27058 7540 27092
rect 7574 27058 7608 27092
rect 7642 27058 7676 27092
rect 7710 27058 7744 27092
rect 7778 27058 7812 27092
rect 7846 27058 7880 27092
rect 7914 27058 7948 27092
rect 7982 27058 8016 27092
rect 8050 27058 8084 27092
rect 8118 27058 8152 27092
rect 8186 27058 8220 27092
rect 8254 27058 8288 27092
rect 8322 27058 8356 27092
rect 8390 27058 8424 27092
rect 8458 27058 8492 27092
rect 8526 27058 8560 27092
rect 8594 27058 8628 27092
rect 8662 27058 8696 27092
rect 8730 27058 8764 27092
rect 8798 27058 8832 27092
rect 8866 27058 8900 27092
rect 8934 27058 8968 27092
rect 9002 27058 9036 27092
rect 9070 27058 9104 27092
rect 9138 27058 9172 27092
rect 9206 27058 9240 27092
rect 9274 27058 9308 27092
rect 9342 27058 9376 27092
rect 9410 27058 9444 27092
rect 9478 27058 9512 27092
rect 9546 27058 9580 27092
rect 9614 27058 9648 27092
rect 9682 27058 9716 27092
rect 9750 27058 9784 27092
rect 9818 27058 9852 27092
rect 9886 27058 9920 27092
rect 9954 27058 9988 27092
rect 10022 27058 10056 27092
rect 10090 27058 10124 27092
rect 10158 27058 10192 27092
rect 10226 27058 10260 27092
rect 10294 27058 10328 27092
rect 10362 27058 10396 27092
rect 10430 27058 10464 27092
rect 10498 27058 10532 27092
rect 10566 27058 10600 27092
rect 10634 27058 10668 27092
rect 10702 27058 10736 27092
rect 10770 27058 10804 27092
rect 10838 27058 10872 27092
rect 10906 27058 10940 27092
rect 10974 27058 11008 27092
rect 11042 27058 11076 27092
rect 11110 27058 11144 27092
rect 11178 27058 11212 27092
rect 11246 27058 11280 27092
rect 11314 27058 11348 27092
rect 11382 27058 11416 27092
rect 11450 27058 11484 27092
rect 11518 27058 11552 27092
rect 11586 27058 11620 27092
rect 11654 27058 11688 27092
rect 11722 27058 11756 27092
rect 11790 27058 11824 27092
rect 11858 27058 11892 27092
rect 11926 27058 11960 27092
rect 11994 27058 12028 27092
rect 12062 27058 12096 27092
rect 12130 27058 12164 27092
rect 12198 27058 12232 27092
rect 12266 27058 12300 27092
rect 12334 27058 12368 27092
rect 12402 27058 12436 27092
rect 12470 27058 12504 27092
rect 12538 27058 12572 27092
rect 12606 27058 12640 27092
rect 12674 27058 12708 27092
rect 12742 27058 12776 27092
rect 12810 27058 12844 27092
rect 12878 27058 12912 27092
rect 12946 27058 12980 27092
rect 13014 27058 13048 27092
rect 13082 27058 13116 27092
rect 13150 27058 13184 27092
rect 13218 27058 13252 27092
rect 13286 27058 13320 27092
rect 13354 27058 13388 27092
rect 13422 27058 13456 27092
rect 13490 27058 13524 27092
rect 13558 27058 13592 27092
rect 13626 27058 13660 27092
rect 13694 27058 13728 27092
rect 13762 27058 13796 27092
rect 13830 27058 13864 27092
rect 13898 27058 13932 27092
rect 13966 27058 14000 27092
rect 14034 27058 14068 27092
rect 14102 27058 14136 27092
rect 14170 27058 14204 27092
rect 14238 27058 14272 27092
rect 14306 27058 14340 27092
rect 14374 27058 14408 27092
rect 14442 27058 14476 27092
rect 14510 27058 14544 27092
rect 14578 27058 14612 27092
rect 14646 27058 14680 27092
rect 14714 27058 14748 27092
rect 14782 27058 14816 27092
rect 14850 27058 14884 27092
rect 14918 27058 14962 27092
rect 2822 27022 14962 27058
rect 2822 26988 2848 27022
rect 2882 26988 2916 27022
rect 2950 26988 2984 27022
rect 3018 26988 3052 27022
rect 3086 26988 3120 27022
rect 3154 26988 3188 27022
rect 3222 26988 3256 27022
rect 3290 26988 3324 27022
rect 3358 26988 3392 27022
rect 3426 26988 3460 27022
rect 3494 26988 3528 27022
rect 3562 26988 3596 27022
rect 3630 26988 3664 27022
rect 3698 26988 3732 27022
rect 3766 26988 3800 27022
rect 3834 26988 3868 27022
rect 3902 26988 3936 27022
rect 3970 26988 4004 27022
rect 4038 26988 4072 27022
rect 4106 26988 4140 27022
rect 4174 26988 4208 27022
rect 4242 26988 4276 27022
rect 4310 26988 4344 27022
rect 4378 26988 4412 27022
rect 4446 26988 4480 27022
rect 4514 26988 4548 27022
rect 4582 26988 4616 27022
rect 4650 26988 4684 27022
rect 4718 26988 4752 27022
rect 4786 26988 4820 27022
rect 4854 26988 4888 27022
rect 4922 26988 4956 27022
rect 4990 26988 5024 27022
rect 5058 26988 5092 27022
rect 5126 26988 5160 27022
rect 5194 26988 5228 27022
rect 5262 26988 5296 27022
rect 5330 26988 5364 27022
rect 5398 26988 5432 27022
rect 5466 26988 5500 27022
rect 5534 26988 5568 27022
rect 5602 26988 5636 27022
rect 5670 26988 5704 27022
rect 5738 26988 5772 27022
rect 5806 26988 5840 27022
rect 5874 26988 5908 27022
rect 5942 26988 5976 27022
rect 6010 26988 6044 27022
rect 6078 26988 6112 27022
rect 6146 26988 6180 27022
rect 6214 26988 6248 27022
rect 6282 26988 6316 27022
rect 6350 26988 6384 27022
rect 6418 26988 6452 27022
rect 6486 26988 6520 27022
rect 6554 26988 6588 27022
rect 6622 26988 6656 27022
rect 6690 26988 6724 27022
rect 6758 26988 6792 27022
rect 6826 26988 6860 27022
rect 6894 26988 6928 27022
rect 6962 26988 6996 27022
rect 7030 26988 7064 27022
rect 7098 26988 7132 27022
rect 7166 26988 7200 27022
rect 7234 26988 7268 27022
rect 7302 26988 7336 27022
rect 7370 26988 7404 27022
rect 7438 26988 7472 27022
rect 7506 26988 7540 27022
rect 7574 26988 7608 27022
rect 7642 26988 7676 27022
rect 7710 26988 7744 27022
rect 7778 26988 7812 27022
rect 7846 26988 7880 27022
rect 7914 26988 7948 27022
rect 7982 26988 8016 27022
rect 8050 26988 8084 27022
rect 8118 26988 8152 27022
rect 8186 26988 8220 27022
rect 8254 26988 8288 27022
rect 8322 26988 8356 27022
rect 8390 26988 8424 27022
rect 8458 26988 8492 27022
rect 8526 26988 8560 27022
rect 8594 26988 8628 27022
rect 8662 26988 8696 27022
rect 8730 26988 8764 27022
rect 8798 26988 8832 27022
rect 8866 26988 8900 27022
rect 8934 26988 8968 27022
rect 9002 26988 9036 27022
rect 9070 26988 9104 27022
rect 9138 26988 9172 27022
rect 9206 26988 9240 27022
rect 9274 26988 9308 27022
rect 9342 26988 9376 27022
rect 9410 26988 9444 27022
rect 9478 26988 9512 27022
rect 9546 26988 9580 27022
rect 9614 26988 9648 27022
rect 9682 26988 9716 27022
rect 9750 26988 9784 27022
rect 9818 26988 9852 27022
rect 9886 26988 9920 27022
rect 9954 26988 9988 27022
rect 10022 26988 10056 27022
rect 10090 26988 10124 27022
rect 10158 26988 10192 27022
rect 10226 26988 10260 27022
rect 10294 26988 10328 27022
rect 10362 26988 10396 27022
rect 10430 26988 10464 27022
rect 10498 26988 10532 27022
rect 10566 26988 10600 27022
rect 10634 26988 10668 27022
rect 10702 26988 10736 27022
rect 10770 26988 10804 27022
rect 10838 26988 10872 27022
rect 10906 26988 10940 27022
rect 10974 26988 11008 27022
rect 11042 26988 11076 27022
rect 11110 26988 11144 27022
rect 11178 26988 11212 27022
rect 11246 26988 11280 27022
rect 11314 26988 11348 27022
rect 11382 26988 11416 27022
rect 11450 26988 11484 27022
rect 11518 26988 11552 27022
rect 11586 26988 11620 27022
rect 11654 26988 11688 27022
rect 11722 26988 11756 27022
rect 11790 26988 11824 27022
rect 11858 26988 11892 27022
rect 11926 26988 11960 27022
rect 11994 26988 12028 27022
rect 12062 26988 12096 27022
rect 12130 26988 12164 27022
rect 12198 26988 12232 27022
rect 12266 26988 12300 27022
rect 12334 26988 12368 27022
rect 12402 26988 12436 27022
rect 12470 26988 12504 27022
rect 12538 26988 12572 27022
rect 12606 26988 12640 27022
rect 12674 26988 12708 27022
rect 12742 26988 12776 27022
rect 12810 26988 12844 27022
rect 12878 26988 12912 27022
rect 12946 26988 12980 27022
rect 13014 26988 13048 27022
rect 13082 26988 13116 27022
rect 13150 26988 13184 27022
rect 13218 26988 13252 27022
rect 13286 26988 13320 27022
rect 13354 26988 13388 27022
rect 13422 26988 13456 27022
rect 13490 26988 13524 27022
rect 13558 26988 13592 27022
rect 13626 26988 13660 27022
rect 13694 26988 13728 27022
rect 13762 26988 13796 27022
rect 13830 26988 13864 27022
rect 13898 26988 13932 27022
rect 13966 26988 14000 27022
rect 14034 26988 14068 27022
rect 14102 26988 14136 27022
rect 14170 26988 14204 27022
rect 14238 26988 14272 27022
rect 14306 26988 14340 27022
rect 14374 26988 14408 27022
rect 14442 26988 14476 27022
rect 14510 26988 14544 27022
rect 14578 26988 14612 27022
rect 14646 26988 14680 27022
rect 14714 26988 14748 27022
rect 14782 26988 14816 27022
rect 14850 26988 14884 27022
rect 14918 26988 14962 27022
rect 2822 26952 14962 26988
rect 2822 26918 2848 26952
rect 2882 26918 2916 26952
rect 2950 26918 2984 26952
rect 3018 26918 3052 26952
rect 3086 26918 3120 26952
rect 3154 26918 3188 26952
rect 3222 26918 3256 26952
rect 3290 26918 3324 26952
rect 3358 26918 3392 26952
rect 3426 26918 3460 26952
rect 3494 26918 3528 26952
rect 3562 26918 3596 26952
rect 3630 26918 3664 26952
rect 3698 26918 3732 26952
rect 3766 26918 3800 26952
rect 3834 26918 3868 26952
rect 3902 26918 3936 26952
rect 3970 26918 4004 26952
rect 4038 26918 4072 26952
rect 4106 26918 4140 26952
rect 4174 26918 4208 26952
rect 4242 26918 4276 26952
rect 4310 26918 4344 26952
rect 4378 26918 4412 26952
rect 4446 26918 4480 26952
rect 4514 26918 4548 26952
rect 4582 26918 4616 26952
rect 4650 26918 4684 26952
rect 4718 26918 4752 26952
rect 4786 26918 4820 26952
rect 4854 26918 4888 26952
rect 4922 26918 4956 26952
rect 4990 26918 5024 26952
rect 5058 26918 5092 26952
rect 5126 26918 5160 26952
rect 5194 26918 5228 26952
rect 5262 26918 5296 26952
rect 5330 26918 5364 26952
rect 5398 26918 5432 26952
rect 5466 26918 5500 26952
rect 5534 26918 5568 26952
rect 5602 26918 5636 26952
rect 5670 26918 5704 26952
rect 5738 26918 5772 26952
rect 5806 26918 5840 26952
rect 5874 26918 5908 26952
rect 5942 26918 5976 26952
rect 6010 26918 6044 26952
rect 6078 26918 6112 26952
rect 6146 26918 6180 26952
rect 6214 26918 6248 26952
rect 6282 26918 6316 26952
rect 6350 26918 6384 26952
rect 6418 26918 6452 26952
rect 6486 26918 6520 26952
rect 6554 26918 6588 26952
rect 6622 26918 6656 26952
rect 6690 26918 6724 26952
rect 6758 26918 6792 26952
rect 6826 26918 6860 26952
rect 6894 26918 6928 26952
rect 6962 26918 6996 26952
rect 7030 26918 7064 26952
rect 7098 26918 7132 26952
rect 7166 26918 7200 26952
rect 7234 26918 7268 26952
rect 7302 26918 7336 26952
rect 7370 26918 7404 26952
rect 7438 26918 7472 26952
rect 7506 26918 7540 26952
rect 7574 26918 7608 26952
rect 7642 26918 7676 26952
rect 7710 26918 7744 26952
rect 7778 26918 7812 26952
rect 7846 26918 7880 26952
rect 7914 26918 7948 26952
rect 7982 26918 8016 26952
rect 8050 26918 8084 26952
rect 8118 26918 8152 26952
rect 8186 26918 8220 26952
rect 8254 26918 8288 26952
rect 8322 26918 8356 26952
rect 8390 26918 8424 26952
rect 8458 26918 8492 26952
rect 8526 26918 8560 26952
rect 8594 26918 8628 26952
rect 8662 26918 8696 26952
rect 8730 26918 8764 26952
rect 8798 26918 8832 26952
rect 8866 26918 8900 26952
rect 8934 26918 8968 26952
rect 9002 26918 9036 26952
rect 9070 26918 9104 26952
rect 9138 26918 9172 26952
rect 9206 26918 9240 26952
rect 9274 26918 9308 26952
rect 9342 26918 9376 26952
rect 9410 26918 9444 26952
rect 9478 26918 9512 26952
rect 9546 26918 9580 26952
rect 9614 26918 9648 26952
rect 9682 26918 9716 26952
rect 9750 26918 9784 26952
rect 9818 26918 9852 26952
rect 9886 26918 9920 26952
rect 9954 26918 9988 26952
rect 10022 26918 10056 26952
rect 10090 26918 10124 26952
rect 10158 26918 10192 26952
rect 10226 26918 10260 26952
rect 10294 26918 10328 26952
rect 10362 26918 10396 26952
rect 10430 26918 10464 26952
rect 10498 26918 10532 26952
rect 10566 26918 10600 26952
rect 10634 26918 10668 26952
rect 10702 26918 10736 26952
rect 10770 26918 10804 26952
rect 10838 26918 10872 26952
rect 10906 26918 10940 26952
rect 10974 26918 11008 26952
rect 11042 26918 11076 26952
rect 11110 26918 11144 26952
rect 11178 26918 11212 26952
rect 11246 26918 11280 26952
rect 11314 26918 11348 26952
rect 11382 26918 11416 26952
rect 11450 26918 11484 26952
rect 11518 26918 11552 26952
rect 11586 26918 11620 26952
rect 11654 26918 11688 26952
rect 11722 26918 11756 26952
rect 11790 26918 11824 26952
rect 11858 26918 11892 26952
rect 11926 26918 11960 26952
rect 11994 26918 12028 26952
rect 12062 26918 12096 26952
rect 12130 26918 12164 26952
rect 12198 26918 12232 26952
rect 12266 26918 12300 26952
rect 12334 26918 12368 26952
rect 12402 26918 12436 26952
rect 12470 26918 12504 26952
rect 12538 26918 12572 26952
rect 12606 26918 12640 26952
rect 12674 26918 12708 26952
rect 12742 26918 12776 26952
rect 12810 26918 12844 26952
rect 12878 26918 12912 26952
rect 12946 26918 12980 26952
rect 13014 26918 13048 26952
rect 13082 26918 13116 26952
rect 13150 26918 13184 26952
rect 13218 26918 13252 26952
rect 13286 26918 13320 26952
rect 13354 26918 13388 26952
rect 13422 26918 13456 26952
rect 13490 26918 13524 26952
rect 13558 26918 13592 26952
rect 13626 26918 13660 26952
rect 13694 26918 13728 26952
rect 13762 26918 13796 26952
rect 13830 26918 13864 26952
rect 13898 26918 13932 26952
rect 13966 26918 14000 26952
rect 14034 26918 14068 26952
rect 14102 26918 14136 26952
rect 14170 26918 14204 26952
rect 14238 26918 14272 26952
rect 14306 26918 14340 26952
rect 14374 26918 14408 26952
rect 14442 26918 14476 26952
rect 14510 26918 14544 26952
rect 14578 26918 14612 26952
rect 14646 26918 14680 26952
rect 14714 26918 14748 26952
rect 14782 26918 14816 26952
rect 14850 26918 14884 26952
rect 14918 26918 14962 26952
rect 2822 26882 14962 26918
rect 2822 26848 2848 26882
rect 2882 26848 2916 26882
rect 2950 26848 2984 26882
rect 3018 26848 3052 26882
rect 3086 26848 3120 26882
rect 3154 26848 3188 26882
rect 3222 26848 3256 26882
rect 3290 26848 3324 26882
rect 3358 26848 3392 26882
rect 3426 26848 3460 26882
rect 3494 26848 3528 26882
rect 3562 26848 3596 26882
rect 3630 26848 3664 26882
rect 3698 26848 3732 26882
rect 3766 26848 3800 26882
rect 3834 26848 3868 26882
rect 3902 26848 3936 26882
rect 3970 26848 4004 26882
rect 4038 26848 4072 26882
rect 4106 26848 4140 26882
rect 4174 26848 4208 26882
rect 4242 26848 4276 26882
rect 4310 26848 4344 26882
rect 4378 26848 4412 26882
rect 4446 26848 4480 26882
rect 4514 26848 4548 26882
rect 4582 26848 4616 26882
rect 4650 26848 4684 26882
rect 4718 26848 4752 26882
rect 4786 26848 4820 26882
rect 4854 26848 4888 26882
rect 4922 26848 4956 26882
rect 4990 26848 5024 26882
rect 5058 26848 5092 26882
rect 5126 26848 5160 26882
rect 5194 26848 5228 26882
rect 5262 26848 5296 26882
rect 5330 26848 5364 26882
rect 5398 26848 5432 26882
rect 5466 26848 5500 26882
rect 5534 26848 5568 26882
rect 5602 26848 5636 26882
rect 5670 26848 5704 26882
rect 5738 26848 5772 26882
rect 5806 26848 5840 26882
rect 5874 26848 5908 26882
rect 5942 26848 5976 26882
rect 6010 26848 6044 26882
rect 6078 26848 6112 26882
rect 6146 26848 6180 26882
rect 6214 26848 6248 26882
rect 6282 26848 6316 26882
rect 6350 26848 6384 26882
rect 6418 26848 6452 26882
rect 6486 26848 6520 26882
rect 6554 26848 6588 26882
rect 6622 26848 6656 26882
rect 6690 26848 6724 26882
rect 6758 26848 6792 26882
rect 6826 26848 6860 26882
rect 6894 26848 6928 26882
rect 6962 26848 6996 26882
rect 7030 26848 7064 26882
rect 7098 26848 7132 26882
rect 7166 26848 7200 26882
rect 7234 26848 7268 26882
rect 7302 26848 7336 26882
rect 7370 26848 7404 26882
rect 7438 26848 7472 26882
rect 7506 26848 7540 26882
rect 7574 26848 7608 26882
rect 7642 26848 7676 26882
rect 7710 26848 7744 26882
rect 7778 26848 7812 26882
rect 7846 26848 7880 26882
rect 7914 26848 7948 26882
rect 7982 26848 8016 26882
rect 8050 26848 8084 26882
rect 8118 26848 8152 26882
rect 8186 26848 8220 26882
rect 8254 26848 8288 26882
rect 8322 26848 8356 26882
rect 8390 26848 8424 26882
rect 8458 26848 8492 26882
rect 8526 26848 8560 26882
rect 8594 26848 8628 26882
rect 8662 26848 8696 26882
rect 8730 26848 8764 26882
rect 8798 26848 8832 26882
rect 8866 26848 8900 26882
rect 8934 26848 8968 26882
rect 9002 26848 9036 26882
rect 9070 26848 9104 26882
rect 9138 26848 9172 26882
rect 9206 26848 9240 26882
rect 9274 26848 9308 26882
rect 9342 26848 9376 26882
rect 9410 26848 9444 26882
rect 9478 26848 9512 26882
rect 9546 26848 9580 26882
rect 9614 26848 9648 26882
rect 9682 26848 9716 26882
rect 9750 26848 9784 26882
rect 9818 26848 9852 26882
rect 9886 26848 9920 26882
rect 9954 26848 9988 26882
rect 10022 26848 10056 26882
rect 10090 26848 10124 26882
rect 10158 26848 10192 26882
rect 10226 26848 10260 26882
rect 10294 26848 10328 26882
rect 10362 26848 10396 26882
rect 10430 26848 10464 26882
rect 10498 26848 10532 26882
rect 10566 26848 10600 26882
rect 10634 26848 10668 26882
rect 10702 26848 10736 26882
rect 10770 26848 10804 26882
rect 10838 26848 10872 26882
rect 10906 26848 10940 26882
rect 10974 26848 11008 26882
rect 11042 26848 11076 26882
rect 11110 26848 11144 26882
rect 11178 26848 11212 26882
rect 11246 26848 11280 26882
rect 11314 26848 11348 26882
rect 11382 26848 11416 26882
rect 11450 26848 11484 26882
rect 11518 26848 11552 26882
rect 11586 26848 11620 26882
rect 11654 26848 11688 26882
rect 11722 26848 11756 26882
rect 11790 26848 11824 26882
rect 11858 26848 11892 26882
rect 11926 26848 11960 26882
rect 11994 26848 12028 26882
rect 12062 26848 12096 26882
rect 12130 26848 12164 26882
rect 12198 26848 12232 26882
rect 12266 26848 12300 26882
rect 12334 26848 12368 26882
rect 12402 26848 12436 26882
rect 12470 26848 12504 26882
rect 12538 26848 12572 26882
rect 12606 26848 12640 26882
rect 12674 26848 12708 26882
rect 12742 26848 12776 26882
rect 12810 26848 12844 26882
rect 12878 26848 12912 26882
rect 12946 26848 12980 26882
rect 13014 26848 13048 26882
rect 13082 26848 13116 26882
rect 13150 26848 13184 26882
rect 13218 26848 13252 26882
rect 13286 26848 13320 26882
rect 13354 26848 13388 26882
rect 13422 26848 13456 26882
rect 13490 26848 13524 26882
rect 13558 26848 13592 26882
rect 13626 26848 13660 26882
rect 13694 26848 13728 26882
rect 13762 26848 13796 26882
rect 13830 26848 13864 26882
rect 13898 26848 13932 26882
rect 13966 26848 14000 26882
rect 14034 26848 14068 26882
rect 14102 26848 14136 26882
rect 14170 26848 14204 26882
rect 14238 26848 14272 26882
rect 14306 26848 14340 26882
rect 14374 26848 14408 26882
rect 14442 26848 14476 26882
rect 14510 26848 14544 26882
rect 14578 26848 14612 26882
rect 14646 26848 14680 26882
rect 14714 26848 14748 26882
rect 14782 26848 14816 26882
rect 14850 26848 14884 26882
rect 14918 26848 14962 26882
rect 2822 26812 14962 26848
rect 2822 26794 2848 26812
rect 49 26778 2848 26794
rect 2882 26778 2916 26812
rect 2950 26778 2984 26812
rect 3018 26778 3052 26812
rect 3086 26778 3120 26812
rect 3154 26778 3188 26812
rect 3222 26778 3256 26812
rect 3290 26778 3324 26812
rect 3358 26778 3392 26812
rect 3426 26778 3460 26812
rect 3494 26778 3528 26812
rect 3562 26778 3596 26812
rect 3630 26778 3664 26812
rect 3698 26778 3732 26812
rect 3766 26778 3800 26812
rect 3834 26778 3868 26812
rect 3902 26778 3936 26812
rect 3970 26778 4004 26812
rect 4038 26778 4072 26812
rect 4106 26778 4140 26812
rect 4174 26778 4208 26812
rect 4242 26778 4276 26812
rect 4310 26778 4344 26812
rect 4378 26778 4412 26812
rect 4446 26778 4480 26812
rect 4514 26778 4548 26812
rect 4582 26778 4616 26812
rect 4650 26778 4684 26812
rect 4718 26778 4752 26812
rect 4786 26778 4820 26812
rect 4854 26778 4888 26812
rect 4922 26778 4956 26812
rect 4990 26778 5024 26812
rect 5058 26778 5092 26812
rect 5126 26778 5160 26812
rect 5194 26778 5228 26812
rect 5262 26778 5296 26812
rect 5330 26778 5364 26812
rect 5398 26778 5432 26812
rect 5466 26778 5500 26812
rect 5534 26778 5568 26812
rect 5602 26778 5636 26812
rect 5670 26778 5704 26812
rect 5738 26778 5772 26812
rect 5806 26778 5840 26812
rect 5874 26778 5908 26812
rect 5942 26778 5976 26812
rect 6010 26778 6044 26812
rect 6078 26778 6112 26812
rect 6146 26778 6180 26812
rect 6214 26778 6248 26812
rect 6282 26778 6316 26812
rect 6350 26778 6384 26812
rect 6418 26778 6452 26812
rect 6486 26778 6520 26812
rect 6554 26778 6588 26812
rect 6622 26778 6656 26812
rect 6690 26778 6724 26812
rect 6758 26778 6792 26812
rect 6826 26778 6860 26812
rect 6894 26778 6928 26812
rect 6962 26778 6996 26812
rect 7030 26778 7064 26812
rect 7098 26778 7132 26812
rect 7166 26778 7200 26812
rect 7234 26778 7268 26812
rect 7302 26778 7336 26812
rect 7370 26778 7404 26812
rect 7438 26778 7472 26812
rect 7506 26778 7540 26812
rect 7574 26778 7608 26812
rect 7642 26778 7676 26812
rect 7710 26778 7744 26812
rect 7778 26778 7812 26812
rect 7846 26778 7880 26812
rect 7914 26778 7948 26812
rect 7982 26778 8016 26812
rect 8050 26778 8084 26812
rect 8118 26778 8152 26812
rect 8186 26778 8220 26812
rect 8254 26778 8288 26812
rect 8322 26778 8356 26812
rect 8390 26778 8424 26812
rect 8458 26778 8492 26812
rect 8526 26778 8560 26812
rect 8594 26778 8628 26812
rect 8662 26778 8696 26812
rect 8730 26778 8764 26812
rect 8798 26778 8832 26812
rect 8866 26778 8900 26812
rect 8934 26778 8968 26812
rect 9002 26778 9036 26812
rect 9070 26778 9104 26812
rect 9138 26778 9172 26812
rect 9206 26778 9240 26812
rect 9274 26778 9308 26812
rect 9342 26778 9376 26812
rect 9410 26778 9444 26812
rect 9478 26778 9512 26812
rect 9546 26778 9580 26812
rect 9614 26778 9648 26812
rect 9682 26778 9716 26812
rect 9750 26778 9784 26812
rect 9818 26778 9852 26812
rect 9886 26778 9920 26812
rect 9954 26778 9988 26812
rect 10022 26778 10056 26812
rect 10090 26778 10124 26812
rect 10158 26778 10192 26812
rect 10226 26778 10260 26812
rect 10294 26778 10328 26812
rect 10362 26778 10396 26812
rect 10430 26778 10464 26812
rect 10498 26778 10532 26812
rect 10566 26778 10600 26812
rect 10634 26778 10668 26812
rect 10702 26778 10736 26812
rect 10770 26778 10804 26812
rect 10838 26778 10872 26812
rect 10906 26778 10940 26812
rect 10974 26778 11008 26812
rect 11042 26778 11076 26812
rect 11110 26778 11144 26812
rect 11178 26778 11212 26812
rect 11246 26778 11280 26812
rect 11314 26778 11348 26812
rect 11382 26778 11416 26812
rect 11450 26778 11484 26812
rect 11518 26778 11552 26812
rect 11586 26778 11620 26812
rect 11654 26778 11688 26812
rect 11722 26778 11756 26812
rect 11790 26778 11824 26812
rect 11858 26778 11892 26812
rect 11926 26778 11960 26812
rect 11994 26778 12028 26812
rect 12062 26778 12096 26812
rect 12130 26778 12164 26812
rect 12198 26778 12232 26812
rect 12266 26778 12300 26812
rect 12334 26778 12368 26812
rect 12402 26778 12436 26812
rect 12470 26778 12504 26812
rect 12538 26778 12572 26812
rect 12606 26778 12640 26812
rect 12674 26778 12708 26812
rect 12742 26778 12776 26812
rect 12810 26778 12844 26812
rect 12878 26778 12912 26812
rect 12946 26778 12980 26812
rect 13014 26778 13048 26812
rect 13082 26778 13116 26812
rect 13150 26778 13184 26812
rect 13218 26778 13252 26812
rect 13286 26778 13320 26812
rect 13354 26778 13388 26812
rect 13422 26778 13456 26812
rect 13490 26778 13524 26812
rect 13558 26778 13592 26812
rect 13626 26778 13660 26812
rect 13694 26778 13728 26812
rect 13762 26778 13796 26812
rect 13830 26778 13864 26812
rect 13898 26778 13932 26812
rect 13966 26778 14000 26812
rect 14034 26778 14068 26812
rect 14102 26778 14136 26812
rect 14170 26778 14204 26812
rect 14238 26778 14272 26812
rect 14306 26778 14340 26812
rect 14374 26778 14408 26812
rect 14442 26778 14476 26812
rect 14510 26778 14544 26812
rect 14578 26778 14612 26812
rect 14646 26778 14680 26812
rect 14714 26778 14748 26812
rect 14782 26778 14816 26812
rect 14850 26778 14884 26812
rect 14918 26778 14962 26812
rect 49 26757 14962 26778
rect 49 26723 83 26757
rect 117 26723 152 26757
rect 186 26723 221 26757
rect 255 26723 290 26757
rect 324 26723 359 26757
rect 393 26723 428 26757
rect 462 26723 497 26757
rect 531 26723 566 26757
rect 600 26723 635 26757
rect 669 26723 704 26757
rect 738 26723 773 26757
rect 807 26723 842 26757
rect 876 26723 911 26757
rect 945 26723 980 26757
rect 1014 26723 1049 26757
rect 1083 26723 1118 26757
rect 1152 26723 1187 26757
rect 1221 26723 1256 26757
rect 1290 26723 1325 26757
rect 1359 26723 1394 26757
rect 1428 26723 1463 26757
rect 1497 26723 1532 26757
rect 1566 26723 1601 26757
rect 1635 26723 1670 26757
rect 1704 26723 1739 26757
rect 1773 26723 1808 26757
rect 1842 26723 1877 26757
rect 1911 26723 1946 26757
rect 1980 26723 2014 26757
rect 2048 26723 2082 26757
rect 2116 26723 2150 26757
rect 2184 26723 2218 26757
rect 2252 26723 2286 26757
rect 2320 26723 2354 26757
rect 2388 26723 2422 26757
rect 2456 26723 2490 26757
rect 2524 26723 2558 26757
rect 2592 26723 2626 26757
rect 2660 26723 2694 26757
rect 2728 26723 2762 26757
rect 2796 26742 14962 26757
rect 2796 26723 2848 26742
rect 49 26708 2848 26723
rect 2882 26708 2916 26742
rect 2950 26708 2984 26742
rect 3018 26708 3052 26742
rect 3086 26708 3120 26742
rect 3154 26708 3188 26742
rect 3222 26708 3256 26742
rect 3290 26708 3324 26742
rect 3358 26708 3392 26742
rect 3426 26708 3460 26742
rect 3494 26708 3528 26742
rect 3562 26708 3596 26742
rect 3630 26708 3664 26742
rect 3698 26708 3732 26742
rect 3766 26708 3800 26742
rect 3834 26708 3868 26742
rect 3902 26708 3936 26742
rect 3970 26708 4004 26742
rect 4038 26708 4072 26742
rect 4106 26708 4140 26742
rect 4174 26708 4208 26742
rect 4242 26708 4276 26742
rect 4310 26708 4344 26742
rect 4378 26708 4412 26742
rect 4446 26708 4480 26742
rect 4514 26708 4548 26742
rect 4582 26708 4616 26742
rect 4650 26708 4684 26742
rect 4718 26708 4752 26742
rect 4786 26708 4820 26742
rect 4854 26708 4888 26742
rect 4922 26708 4956 26742
rect 4990 26708 5024 26742
rect 5058 26708 5092 26742
rect 5126 26708 5160 26742
rect 5194 26708 5228 26742
rect 5262 26708 5296 26742
rect 5330 26708 5364 26742
rect 5398 26708 5432 26742
rect 5466 26708 5500 26742
rect 5534 26708 5568 26742
rect 5602 26708 5636 26742
rect 5670 26708 5704 26742
rect 5738 26708 5772 26742
rect 5806 26708 5840 26742
rect 5874 26708 5908 26742
rect 5942 26708 5976 26742
rect 6010 26708 6044 26742
rect 6078 26708 6112 26742
rect 6146 26708 6180 26742
rect 6214 26708 6248 26742
rect 6282 26708 6316 26742
rect 6350 26708 6384 26742
rect 6418 26708 6452 26742
rect 6486 26708 6520 26742
rect 6554 26708 6588 26742
rect 6622 26708 6656 26742
rect 6690 26708 6724 26742
rect 6758 26708 6792 26742
rect 6826 26708 6860 26742
rect 6894 26708 6928 26742
rect 6962 26708 6996 26742
rect 7030 26708 7064 26742
rect 7098 26708 7132 26742
rect 7166 26708 7200 26742
rect 7234 26708 7268 26742
rect 7302 26708 7336 26742
rect 7370 26708 7404 26742
rect 7438 26708 7472 26742
rect 7506 26708 7540 26742
rect 7574 26708 7608 26742
rect 7642 26708 7676 26742
rect 7710 26708 7744 26742
rect 7778 26708 7812 26742
rect 7846 26708 7880 26742
rect 7914 26708 7948 26742
rect 7982 26708 8016 26742
rect 8050 26708 8084 26742
rect 8118 26708 8152 26742
rect 8186 26708 8220 26742
rect 8254 26708 8288 26742
rect 8322 26708 8356 26742
rect 8390 26708 8424 26742
rect 8458 26708 8492 26742
rect 8526 26708 8560 26742
rect 8594 26708 8628 26742
rect 8662 26708 8696 26742
rect 8730 26708 8764 26742
rect 8798 26708 8832 26742
rect 8866 26708 8900 26742
rect 8934 26708 8968 26742
rect 9002 26708 9036 26742
rect 9070 26708 9104 26742
rect 9138 26708 9172 26742
rect 9206 26708 9240 26742
rect 9274 26708 9308 26742
rect 9342 26708 9376 26742
rect 9410 26708 9444 26742
rect 9478 26708 9512 26742
rect 9546 26708 9580 26742
rect 9614 26708 9648 26742
rect 9682 26708 9716 26742
rect 9750 26708 9784 26742
rect 9818 26708 9852 26742
rect 9886 26708 9920 26742
rect 9954 26708 9988 26742
rect 10022 26708 10056 26742
rect 10090 26708 10124 26742
rect 10158 26708 10192 26742
rect 10226 26708 10260 26742
rect 10294 26708 10328 26742
rect 10362 26708 10396 26742
rect 10430 26708 10464 26742
rect 10498 26708 10532 26742
rect 10566 26708 10600 26742
rect 10634 26708 10668 26742
rect 10702 26708 10736 26742
rect 10770 26708 10804 26742
rect 10838 26708 10872 26742
rect 10906 26708 10940 26742
rect 10974 26708 11008 26742
rect 11042 26708 11076 26742
rect 11110 26708 11144 26742
rect 11178 26708 11212 26742
rect 11246 26708 11280 26742
rect 11314 26708 11348 26742
rect 11382 26708 11416 26742
rect 11450 26708 11484 26742
rect 11518 26708 11552 26742
rect 11586 26708 11620 26742
rect 11654 26708 11688 26742
rect 11722 26708 11756 26742
rect 11790 26708 11824 26742
rect 11858 26708 11892 26742
rect 11926 26708 11960 26742
rect 11994 26708 12028 26742
rect 12062 26708 12096 26742
rect 12130 26708 12164 26742
rect 12198 26708 12232 26742
rect 12266 26708 12300 26742
rect 12334 26708 12368 26742
rect 12402 26708 12436 26742
rect 12470 26708 12504 26742
rect 12538 26708 12572 26742
rect 12606 26708 12640 26742
rect 12674 26708 12708 26742
rect 12742 26708 12776 26742
rect 12810 26708 12844 26742
rect 12878 26708 12912 26742
rect 12946 26708 12980 26742
rect 13014 26708 13048 26742
rect 13082 26708 13116 26742
rect 13150 26708 13184 26742
rect 13218 26708 13252 26742
rect 13286 26708 13320 26742
rect 13354 26708 13388 26742
rect 13422 26708 13456 26742
rect 13490 26708 13524 26742
rect 13558 26708 13592 26742
rect 13626 26708 13660 26742
rect 13694 26708 13728 26742
rect 13762 26708 13796 26742
rect 13830 26708 13864 26742
rect 13898 26708 13932 26742
rect 13966 26708 14000 26742
rect 14034 26708 14068 26742
rect 14102 26708 14136 26742
rect 14170 26708 14204 26742
rect 14238 26708 14272 26742
rect 14306 26708 14340 26742
rect 14374 26708 14408 26742
rect 14442 26708 14476 26742
rect 14510 26708 14544 26742
rect 14578 26708 14612 26742
rect 14646 26708 14680 26742
rect 14714 26708 14748 26742
rect 14782 26708 14816 26742
rect 14850 26708 14884 26742
rect 14918 26708 14962 26742
rect 49 26683 14962 26708
rect 49 26649 83 26683
rect 117 26649 152 26683
rect 186 26649 221 26683
rect 255 26649 290 26683
rect 324 26649 359 26683
rect 393 26649 428 26683
rect 462 26649 497 26683
rect 531 26649 566 26683
rect 600 26649 635 26683
rect 669 26649 704 26683
rect 738 26649 773 26683
rect 807 26649 842 26683
rect 876 26649 911 26683
rect 945 26649 980 26683
rect 1014 26649 1049 26683
rect 1083 26649 1118 26683
rect 1152 26649 1187 26683
rect 1221 26649 1256 26683
rect 1290 26649 1325 26683
rect 1359 26649 1394 26683
rect 1428 26649 1463 26683
rect 1497 26649 1532 26683
rect 1566 26649 1601 26683
rect 1635 26649 1670 26683
rect 1704 26649 1739 26683
rect 1773 26649 1808 26683
rect 1842 26649 1877 26683
rect 1911 26649 1946 26683
rect 1980 26649 2014 26683
rect 2048 26649 2082 26683
rect 2116 26649 2150 26683
rect 2184 26649 2218 26683
rect 2252 26649 2286 26683
rect 2320 26649 2354 26683
rect 2388 26649 2422 26683
rect 2456 26649 2490 26683
rect 2524 26649 2558 26683
rect 2592 26649 2626 26683
rect 2660 26649 2694 26683
rect 2728 26649 2762 26683
rect 2796 26672 14962 26683
rect 2796 26649 2848 26672
rect 49 26638 2848 26649
rect 2882 26638 2916 26672
rect 2950 26638 2984 26672
rect 3018 26638 3052 26672
rect 3086 26638 3120 26672
rect 3154 26638 3188 26672
rect 3222 26638 3256 26672
rect 3290 26638 3324 26672
rect 3358 26638 3392 26672
rect 3426 26638 3460 26672
rect 3494 26638 3528 26672
rect 3562 26638 3596 26672
rect 3630 26638 3664 26672
rect 3698 26638 3732 26672
rect 3766 26638 3800 26672
rect 3834 26638 3868 26672
rect 3902 26638 3936 26672
rect 3970 26638 4004 26672
rect 4038 26638 4072 26672
rect 4106 26638 4140 26672
rect 4174 26638 4208 26672
rect 4242 26638 4276 26672
rect 4310 26638 4344 26672
rect 4378 26638 4412 26672
rect 4446 26638 4480 26672
rect 4514 26638 4548 26672
rect 4582 26638 4616 26672
rect 4650 26638 4684 26672
rect 4718 26638 4752 26672
rect 4786 26638 4820 26672
rect 4854 26638 4888 26672
rect 4922 26638 4956 26672
rect 4990 26638 5024 26672
rect 5058 26638 5092 26672
rect 5126 26638 5160 26672
rect 5194 26638 5228 26672
rect 5262 26638 5296 26672
rect 5330 26638 5364 26672
rect 5398 26638 5432 26672
rect 5466 26638 5500 26672
rect 5534 26638 5568 26672
rect 5602 26638 5636 26672
rect 5670 26638 5704 26672
rect 5738 26638 5772 26672
rect 5806 26638 5840 26672
rect 5874 26638 5908 26672
rect 5942 26638 5976 26672
rect 6010 26638 6044 26672
rect 6078 26638 6112 26672
rect 6146 26638 6180 26672
rect 6214 26638 6248 26672
rect 6282 26638 6316 26672
rect 6350 26638 6384 26672
rect 6418 26638 6452 26672
rect 6486 26638 6520 26672
rect 6554 26638 6588 26672
rect 6622 26638 6656 26672
rect 6690 26638 6724 26672
rect 6758 26638 6792 26672
rect 6826 26638 6860 26672
rect 6894 26638 6928 26672
rect 6962 26638 6996 26672
rect 7030 26638 7064 26672
rect 7098 26638 7132 26672
rect 7166 26638 7200 26672
rect 7234 26638 7268 26672
rect 7302 26638 7336 26672
rect 7370 26638 7404 26672
rect 7438 26638 7472 26672
rect 7506 26638 7540 26672
rect 7574 26638 7608 26672
rect 7642 26638 7676 26672
rect 7710 26638 7744 26672
rect 7778 26638 7812 26672
rect 7846 26638 7880 26672
rect 7914 26638 7948 26672
rect 7982 26638 8016 26672
rect 8050 26638 8084 26672
rect 8118 26638 8152 26672
rect 8186 26638 8220 26672
rect 8254 26638 8288 26672
rect 8322 26638 8356 26672
rect 8390 26638 8424 26672
rect 8458 26638 8492 26672
rect 8526 26638 8560 26672
rect 8594 26638 8628 26672
rect 8662 26638 8696 26672
rect 8730 26638 8764 26672
rect 8798 26638 8832 26672
rect 8866 26638 8900 26672
rect 8934 26638 8968 26672
rect 9002 26638 9036 26672
rect 9070 26638 9104 26672
rect 9138 26638 9172 26672
rect 9206 26638 9240 26672
rect 9274 26638 9308 26672
rect 9342 26638 9376 26672
rect 9410 26638 9444 26672
rect 9478 26638 9512 26672
rect 9546 26638 9580 26672
rect 9614 26638 9648 26672
rect 9682 26638 9716 26672
rect 9750 26638 9784 26672
rect 9818 26638 9852 26672
rect 9886 26638 9920 26672
rect 9954 26638 9988 26672
rect 10022 26638 10056 26672
rect 10090 26638 10124 26672
rect 10158 26638 10192 26672
rect 10226 26638 10260 26672
rect 10294 26638 10328 26672
rect 10362 26638 10396 26672
rect 10430 26638 10464 26672
rect 10498 26638 10532 26672
rect 10566 26638 10600 26672
rect 10634 26638 10668 26672
rect 10702 26638 10736 26672
rect 10770 26638 10804 26672
rect 10838 26638 10872 26672
rect 10906 26638 10940 26672
rect 10974 26638 11008 26672
rect 11042 26638 11076 26672
rect 11110 26638 11144 26672
rect 11178 26638 11212 26672
rect 11246 26638 11280 26672
rect 11314 26638 11348 26672
rect 11382 26638 11416 26672
rect 11450 26638 11484 26672
rect 11518 26638 11552 26672
rect 11586 26638 11620 26672
rect 11654 26638 11688 26672
rect 11722 26638 11756 26672
rect 11790 26638 11824 26672
rect 11858 26638 11892 26672
rect 11926 26638 11960 26672
rect 11994 26638 12028 26672
rect 12062 26638 12096 26672
rect 12130 26638 12164 26672
rect 12198 26638 12232 26672
rect 12266 26638 12300 26672
rect 12334 26638 12368 26672
rect 12402 26638 12436 26672
rect 12470 26638 12504 26672
rect 12538 26638 12572 26672
rect 12606 26638 12640 26672
rect 12674 26638 12708 26672
rect 12742 26638 12776 26672
rect 12810 26638 12844 26672
rect 12878 26638 12912 26672
rect 12946 26638 12980 26672
rect 13014 26638 13048 26672
rect 13082 26638 13116 26672
rect 13150 26638 13184 26672
rect 13218 26638 13252 26672
rect 13286 26638 13320 26672
rect 13354 26638 13388 26672
rect 13422 26638 13456 26672
rect 13490 26638 13524 26672
rect 13558 26638 13592 26672
rect 13626 26638 13660 26672
rect 13694 26638 13728 26672
rect 13762 26638 13796 26672
rect 13830 26638 13864 26672
rect 13898 26638 13932 26672
rect 13966 26638 14000 26672
rect 14034 26638 14068 26672
rect 14102 26638 14136 26672
rect 14170 26638 14204 26672
rect 14238 26638 14272 26672
rect 14306 26638 14340 26672
rect 14374 26638 14408 26672
rect 14442 26638 14476 26672
rect 14510 26638 14544 26672
rect 14578 26638 14612 26672
rect 14646 26638 14680 26672
rect 14714 26638 14748 26672
rect 14782 26638 14816 26672
rect 14850 26638 14884 26672
rect 14918 26638 14962 26672
rect 49 26609 14962 26638
rect 49 26575 83 26609
rect 117 26575 152 26609
rect 186 26575 221 26609
rect 255 26575 290 26609
rect 324 26575 359 26609
rect 393 26575 428 26609
rect 462 26575 497 26609
rect 531 26575 566 26609
rect 600 26575 635 26609
rect 669 26575 704 26609
rect 738 26575 773 26609
rect 807 26575 842 26609
rect 876 26575 911 26609
rect 945 26575 980 26609
rect 1014 26575 1049 26609
rect 1083 26575 1118 26609
rect 1152 26575 1187 26609
rect 1221 26575 1256 26609
rect 1290 26575 1325 26609
rect 1359 26575 1394 26609
rect 1428 26575 1463 26609
rect 1497 26575 1532 26609
rect 1566 26575 1601 26609
rect 1635 26575 1670 26609
rect 1704 26575 1739 26609
rect 1773 26575 1808 26609
rect 1842 26575 1877 26609
rect 1911 26575 1946 26609
rect 1980 26575 2014 26609
rect 2048 26575 2082 26609
rect 2116 26575 2150 26609
rect 2184 26575 2218 26609
rect 2252 26575 2286 26609
rect 2320 26575 2354 26609
rect 2388 26575 2422 26609
rect 2456 26575 2490 26609
rect 2524 26575 2558 26609
rect 2592 26575 2626 26609
rect 2660 26575 2694 26609
rect 2728 26575 2762 26609
rect 2796 26602 14962 26609
rect 2796 26575 2848 26602
rect 49 26568 2848 26575
rect 2882 26568 2916 26602
rect 2950 26568 2984 26602
rect 3018 26568 3052 26602
rect 3086 26568 3120 26602
rect 3154 26568 3188 26602
rect 3222 26568 3256 26602
rect 3290 26568 3324 26602
rect 3358 26568 3392 26602
rect 3426 26568 3460 26602
rect 3494 26568 3528 26602
rect 3562 26568 3596 26602
rect 3630 26568 3664 26602
rect 3698 26568 3732 26602
rect 3766 26568 3800 26602
rect 3834 26568 3868 26602
rect 3902 26568 3936 26602
rect 3970 26568 4004 26602
rect 4038 26568 4072 26602
rect 4106 26568 4140 26602
rect 4174 26568 4208 26602
rect 4242 26568 4276 26602
rect 4310 26568 4344 26602
rect 4378 26568 4412 26602
rect 4446 26568 4480 26602
rect 4514 26568 4548 26602
rect 4582 26568 4616 26602
rect 4650 26568 4684 26602
rect 4718 26568 4752 26602
rect 4786 26568 4820 26602
rect 4854 26568 4888 26602
rect 4922 26568 4956 26602
rect 4990 26568 5024 26602
rect 5058 26568 5092 26602
rect 5126 26568 5160 26602
rect 5194 26568 5228 26602
rect 5262 26568 5296 26602
rect 5330 26568 5364 26602
rect 5398 26568 5432 26602
rect 5466 26568 5500 26602
rect 5534 26568 5568 26602
rect 5602 26568 5636 26602
rect 5670 26568 5704 26602
rect 5738 26568 5772 26602
rect 5806 26568 5840 26602
rect 5874 26568 5908 26602
rect 5942 26568 5976 26602
rect 6010 26568 6044 26602
rect 6078 26568 6112 26602
rect 6146 26568 6180 26602
rect 6214 26568 6248 26602
rect 6282 26568 6316 26602
rect 6350 26568 6384 26602
rect 6418 26568 6452 26602
rect 6486 26568 6520 26602
rect 6554 26568 6588 26602
rect 6622 26568 6656 26602
rect 6690 26568 6724 26602
rect 6758 26568 6792 26602
rect 6826 26568 6860 26602
rect 6894 26568 6928 26602
rect 6962 26568 6996 26602
rect 7030 26568 7064 26602
rect 7098 26568 7132 26602
rect 7166 26568 7200 26602
rect 7234 26568 7268 26602
rect 7302 26568 7336 26602
rect 7370 26568 7404 26602
rect 7438 26568 7472 26602
rect 7506 26568 7540 26602
rect 7574 26568 7608 26602
rect 7642 26568 7676 26602
rect 7710 26568 7744 26602
rect 7778 26568 7812 26602
rect 7846 26568 7880 26602
rect 7914 26568 7948 26602
rect 7982 26568 8016 26602
rect 8050 26568 8084 26602
rect 8118 26568 8152 26602
rect 8186 26568 8220 26602
rect 8254 26568 8288 26602
rect 8322 26568 8356 26602
rect 8390 26568 8424 26602
rect 8458 26568 8492 26602
rect 8526 26568 8560 26602
rect 8594 26568 8628 26602
rect 8662 26568 8696 26602
rect 8730 26568 8764 26602
rect 8798 26568 8832 26602
rect 8866 26568 8900 26602
rect 8934 26568 8968 26602
rect 9002 26568 9036 26602
rect 9070 26568 9104 26602
rect 9138 26568 9172 26602
rect 9206 26568 9240 26602
rect 9274 26568 9308 26602
rect 9342 26568 9376 26602
rect 9410 26568 9444 26602
rect 9478 26568 9512 26602
rect 9546 26568 9580 26602
rect 9614 26568 9648 26602
rect 9682 26568 9716 26602
rect 9750 26568 9784 26602
rect 9818 26568 9852 26602
rect 9886 26568 9920 26602
rect 9954 26568 9988 26602
rect 10022 26568 10056 26602
rect 10090 26568 10124 26602
rect 10158 26568 10192 26602
rect 10226 26568 10260 26602
rect 10294 26568 10328 26602
rect 10362 26568 10396 26602
rect 10430 26568 10464 26602
rect 10498 26568 10532 26602
rect 10566 26568 10600 26602
rect 10634 26568 10668 26602
rect 10702 26568 10736 26602
rect 10770 26568 10804 26602
rect 10838 26568 10872 26602
rect 10906 26568 10940 26602
rect 10974 26568 11008 26602
rect 11042 26568 11076 26602
rect 11110 26568 11144 26602
rect 11178 26568 11212 26602
rect 11246 26568 11280 26602
rect 11314 26568 11348 26602
rect 11382 26568 11416 26602
rect 11450 26568 11484 26602
rect 11518 26568 11552 26602
rect 11586 26568 11620 26602
rect 11654 26568 11688 26602
rect 11722 26568 11756 26602
rect 11790 26568 11824 26602
rect 11858 26568 11892 26602
rect 11926 26568 11960 26602
rect 11994 26568 12028 26602
rect 12062 26568 12096 26602
rect 12130 26568 12164 26602
rect 12198 26568 12232 26602
rect 12266 26568 12300 26602
rect 12334 26568 12368 26602
rect 12402 26568 12436 26602
rect 12470 26568 12504 26602
rect 12538 26568 12572 26602
rect 12606 26568 12640 26602
rect 12674 26568 12708 26602
rect 12742 26568 12776 26602
rect 12810 26568 12844 26602
rect 12878 26568 12912 26602
rect 12946 26568 12980 26602
rect 13014 26568 13048 26602
rect 13082 26568 13116 26602
rect 13150 26568 13184 26602
rect 13218 26568 13252 26602
rect 13286 26568 13320 26602
rect 13354 26568 13388 26602
rect 13422 26568 13456 26602
rect 13490 26568 13524 26602
rect 13558 26568 13592 26602
rect 13626 26568 13660 26602
rect 13694 26568 13728 26602
rect 13762 26568 13796 26602
rect 13830 26568 13864 26602
rect 13898 26568 13932 26602
rect 13966 26568 14000 26602
rect 14034 26568 14068 26602
rect 14102 26568 14136 26602
rect 14170 26568 14204 26602
rect 14238 26568 14272 26602
rect 14306 26568 14340 26602
rect 14374 26568 14408 26602
rect 14442 26568 14476 26602
rect 14510 26568 14544 26602
rect 14578 26568 14612 26602
rect 14646 26568 14680 26602
rect 14714 26568 14748 26602
rect 14782 26568 14816 26602
rect 14850 26568 14884 26602
rect 14918 26568 14962 26602
rect 49 26535 14962 26568
rect 49 26501 83 26535
rect 117 26501 152 26535
rect 186 26501 221 26535
rect 255 26501 290 26535
rect 324 26501 359 26535
rect 393 26501 428 26535
rect 462 26501 497 26535
rect 531 26501 566 26535
rect 600 26501 635 26535
rect 669 26501 704 26535
rect 738 26501 773 26535
rect 807 26501 842 26535
rect 876 26501 911 26535
rect 945 26501 980 26535
rect 1014 26501 1049 26535
rect 1083 26501 1118 26535
rect 1152 26501 1187 26535
rect 1221 26501 1256 26535
rect 1290 26501 1325 26535
rect 1359 26501 1394 26535
rect 1428 26501 1463 26535
rect 1497 26501 1532 26535
rect 1566 26501 1601 26535
rect 1635 26501 1670 26535
rect 1704 26501 1739 26535
rect 1773 26501 1808 26535
rect 1842 26501 1877 26535
rect 1911 26501 1946 26535
rect 1980 26501 2014 26535
rect 2048 26501 2082 26535
rect 2116 26501 2150 26535
rect 2184 26501 2218 26535
rect 2252 26501 2286 26535
rect 2320 26501 2354 26535
rect 2388 26501 2422 26535
rect 2456 26501 2490 26535
rect 2524 26501 2558 26535
rect 2592 26501 2626 26535
rect 2660 26501 2694 26535
rect 2728 26501 2762 26535
rect 2796 26532 14962 26535
rect 2796 26501 2848 26532
rect 49 26498 2848 26501
rect 2882 26498 2916 26532
rect 2950 26498 2984 26532
rect 3018 26498 3052 26532
rect 3086 26498 3120 26532
rect 3154 26498 3188 26532
rect 3222 26498 3256 26532
rect 3290 26498 3324 26532
rect 3358 26498 3392 26532
rect 3426 26498 3460 26532
rect 3494 26498 3528 26532
rect 3562 26498 3596 26532
rect 3630 26498 3664 26532
rect 3698 26498 3732 26532
rect 3766 26498 3800 26532
rect 3834 26498 3868 26532
rect 3902 26498 3936 26532
rect 3970 26498 4004 26532
rect 4038 26498 4072 26532
rect 4106 26498 4140 26532
rect 4174 26498 4208 26532
rect 4242 26498 4276 26532
rect 4310 26498 4344 26532
rect 4378 26498 4412 26532
rect 4446 26498 4480 26532
rect 4514 26498 4548 26532
rect 4582 26498 4616 26532
rect 4650 26498 4684 26532
rect 4718 26498 4752 26532
rect 4786 26498 4820 26532
rect 4854 26498 4888 26532
rect 4922 26498 4956 26532
rect 4990 26498 5024 26532
rect 5058 26498 5092 26532
rect 5126 26498 5160 26532
rect 5194 26498 5228 26532
rect 5262 26498 5296 26532
rect 5330 26498 5364 26532
rect 5398 26498 5432 26532
rect 5466 26498 5500 26532
rect 5534 26498 5568 26532
rect 5602 26498 5636 26532
rect 5670 26498 5704 26532
rect 5738 26498 5772 26532
rect 5806 26498 5840 26532
rect 5874 26498 5908 26532
rect 5942 26498 5976 26532
rect 6010 26498 6044 26532
rect 6078 26498 6112 26532
rect 6146 26498 6180 26532
rect 6214 26498 6248 26532
rect 6282 26498 6316 26532
rect 6350 26498 6384 26532
rect 6418 26498 6452 26532
rect 6486 26498 6520 26532
rect 6554 26498 6588 26532
rect 6622 26498 6656 26532
rect 6690 26498 6724 26532
rect 6758 26498 6792 26532
rect 6826 26498 6860 26532
rect 6894 26498 6928 26532
rect 6962 26498 6996 26532
rect 7030 26498 7064 26532
rect 7098 26498 7132 26532
rect 7166 26498 7200 26532
rect 7234 26498 7268 26532
rect 7302 26498 7336 26532
rect 7370 26498 7404 26532
rect 7438 26498 7472 26532
rect 7506 26498 7540 26532
rect 7574 26498 7608 26532
rect 7642 26498 7676 26532
rect 7710 26498 7744 26532
rect 7778 26498 7812 26532
rect 7846 26498 7880 26532
rect 7914 26498 7948 26532
rect 7982 26498 8016 26532
rect 8050 26498 8084 26532
rect 8118 26498 8152 26532
rect 8186 26498 8220 26532
rect 8254 26498 8288 26532
rect 8322 26498 8356 26532
rect 8390 26498 8424 26532
rect 8458 26498 8492 26532
rect 8526 26498 8560 26532
rect 8594 26498 8628 26532
rect 8662 26498 8696 26532
rect 8730 26498 8764 26532
rect 8798 26498 8832 26532
rect 8866 26498 8900 26532
rect 8934 26498 8968 26532
rect 9002 26498 9036 26532
rect 9070 26498 9104 26532
rect 9138 26498 9172 26532
rect 9206 26498 9240 26532
rect 9274 26498 9308 26532
rect 9342 26498 9376 26532
rect 9410 26498 9444 26532
rect 9478 26498 9512 26532
rect 9546 26498 9580 26532
rect 9614 26498 9648 26532
rect 9682 26498 9716 26532
rect 9750 26498 9784 26532
rect 9818 26498 9852 26532
rect 9886 26498 9920 26532
rect 9954 26498 9988 26532
rect 10022 26498 10056 26532
rect 10090 26498 10124 26532
rect 10158 26498 10192 26532
rect 10226 26498 10260 26532
rect 10294 26498 10328 26532
rect 10362 26498 10396 26532
rect 10430 26498 10464 26532
rect 10498 26498 10532 26532
rect 10566 26498 10600 26532
rect 10634 26498 10668 26532
rect 10702 26498 10736 26532
rect 10770 26498 10804 26532
rect 10838 26498 10872 26532
rect 10906 26498 10940 26532
rect 10974 26498 11008 26532
rect 11042 26498 11076 26532
rect 11110 26498 11144 26532
rect 11178 26498 11212 26532
rect 11246 26498 11280 26532
rect 11314 26498 11348 26532
rect 11382 26498 11416 26532
rect 11450 26498 11484 26532
rect 11518 26498 11552 26532
rect 11586 26498 11620 26532
rect 11654 26498 11688 26532
rect 11722 26498 11756 26532
rect 11790 26498 11824 26532
rect 11858 26498 11892 26532
rect 11926 26498 11960 26532
rect 11994 26498 12028 26532
rect 12062 26498 12096 26532
rect 12130 26498 12164 26532
rect 12198 26498 12232 26532
rect 12266 26498 12300 26532
rect 12334 26498 12368 26532
rect 12402 26498 12436 26532
rect 12470 26498 12504 26532
rect 12538 26498 12572 26532
rect 12606 26498 12640 26532
rect 12674 26498 12708 26532
rect 12742 26498 12776 26532
rect 12810 26498 12844 26532
rect 12878 26498 12912 26532
rect 12946 26498 12980 26532
rect 13014 26498 13048 26532
rect 13082 26498 13116 26532
rect 13150 26498 13184 26532
rect 13218 26498 13252 26532
rect 13286 26498 13320 26532
rect 13354 26498 13388 26532
rect 13422 26498 13456 26532
rect 13490 26498 13524 26532
rect 13558 26498 13592 26532
rect 13626 26498 13660 26532
rect 13694 26498 13728 26532
rect 13762 26498 13796 26532
rect 13830 26498 13864 26532
rect 13898 26498 13932 26532
rect 13966 26498 14000 26532
rect 14034 26498 14068 26532
rect 14102 26498 14136 26532
rect 14170 26498 14204 26532
rect 14238 26498 14272 26532
rect 14306 26498 14340 26532
rect 14374 26498 14408 26532
rect 14442 26498 14476 26532
rect 14510 26498 14544 26532
rect 14578 26498 14612 26532
rect 14646 26498 14680 26532
rect 14714 26498 14748 26532
rect 14782 26498 14816 26532
rect 14850 26498 14884 26532
rect 14918 26498 14962 26532
rect 49 26462 14962 26498
rect 49 26461 2848 26462
rect 49 26427 83 26461
rect 117 26427 152 26461
rect 186 26427 221 26461
rect 255 26427 290 26461
rect 324 26427 359 26461
rect 393 26427 428 26461
rect 462 26427 497 26461
rect 531 26427 566 26461
rect 600 26427 635 26461
rect 669 26427 704 26461
rect 738 26427 773 26461
rect 807 26427 842 26461
rect 876 26427 911 26461
rect 945 26427 980 26461
rect 1014 26427 1049 26461
rect 1083 26427 1118 26461
rect 1152 26427 1187 26461
rect 1221 26427 1256 26461
rect 1290 26427 1325 26461
rect 1359 26427 1394 26461
rect 1428 26427 1463 26461
rect 1497 26427 1532 26461
rect 1566 26427 1601 26461
rect 1635 26427 1670 26461
rect 1704 26427 1739 26461
rect 1773 26427 1808 26461
rect 1842 26427 1877 26461
rect 1911 26427 1946 26461
rect 1980 26427 2014 26461
rect 2048 26427 2082 26461
rect 2116 26427 2150 26461
rect 2184 26427 2218 26461
rect 2252 26427 2286 26461
rect 2320 26427 2354 26461
rect 2388 26427 2422 26461
rect 2456 26427 2490 26461
rect 2524 26427 2558 26461
rect 2592 26427 2626 26461
rect 2660 26427 2694 26461
rect 2728 26427 2762 26461
rect 2796 26428 2848 26461
rect 2882 26428 2916 26462
rect 2950 26428 2984 26462
rect 3018 26428 3052 26462
rect 3086 26428 3120 26462
rect 3154 26428 3188 26462
rect 3222 26428 3256 26462
rect 3290 26428 3324 26462
rect 3358 26428 3392 26462
rect 3426 26428 3460 26462
rect 3494 26428 3528 26462
rect 3562 26428 3596 26462
rect 3630 26428 3664 26462
rect 3698 26428 3732 26462
rect 3766 26428 3800 26462
rect 3834 26428 3868 26462
rect 3902 26428 3936 26462
rect 3970 26428 4004 26462
rect 4038 26428 4072 26462
rect 4106 26428 4140 26462
rect 4174 26428 4208 26462
rect 4242 26428 4276 26462
rect 4310 26428 4344 26462
rect 4378 26428 4412 26462
rect 4446 26428 4480 26462
rect 4514 26428 4548 26462
rect 4582 26428 4616 26462
rect 4650 26428 4684 26462
rect 4718 26428 4752 26462
rect 4786 26428 4820 26462
rect 4854 26428 4888 26462
rect 4922 26428 4956 26462
rect 4990 26428 5024 26462
rect 5058 26428 5092 26462
rect 5126 26428 5160 26462
rect 5194 26428 5228 26462
rect 5262 26428 5296 26462
rect 5330 26428 5364 26462
rect 5398 26428 5432 26462
rect 5466 26428 5500 26462
rect 5534 26428 5568 26462
rect 5602 26428 5636 26462
rect 5670 26428 5704 26462
rect 5738 26428 5772 26462
rect 5806 26428 5840 26462
rect 5874 26428 5908 26462
rect 5942 26428 5976 26462
rect 6010 26428 6044 26462
rect 6078 26428 6112 26462
rect 6146 26428 6180 26462
rect 6214 26428 6248 26462
rect 6282 26428 6316 26462
rect 6350 26428 6384 26462
rect 6418 26428 6452 26462
rect 6486 26428 6520 26462
rect 6554 26428 6588 26462
rect 6622 26428 6656 26462
rect 6690 26428 6724 26462
rect 6758 26428 6792 26462
rect 6826 26428 6860 26462
rect 6894 26428 6928 26462
rect 6962 26428 6996 26462
rect 7030 26428 7064 26462
rect 7098 26428 7132 26462
rect 7166 26428 7200 26462
rect 7234 26428 7268 26462
rect 7302 26428 7336 26462
rect 7370 26428 7404 26462
rect 7438 26428 7472 26462
rect 7506 26428 7540 26462
rect 7574 26428 7608 26462
rect 7642 26428 7676 26462
rect 7710 26428 7744 26462
rect 7778 26428 7812 26462
rect 7846 26428 7880 26462
rect 7914 26428 7948 26462
rect 7982 26428 8016 26462
rect 8050 26428 8084 26462
rect 8118 26428 8152 26462
rect 8186 26428 8220 26462
rect 8254 26428 8288 26462
rect 8322 26428 8356 26462
rect 8390 26428 8424 26462
rect 8458 26428 8492 26462
rect 8526 26428 8560 26462
rect 8594 26428 8628 26462
rect 8662 26428 8696 26462
rect 8730 26428 8764 26462
rect 8798 26428 8832 26462
rect 8866 26428 8900 26462
rect 8934 26428 8968 26462
rect 9002 26428 9036 26462
rect 9070 26428 9104 26462
rect 9138 26428 9172 26462
rect 9206 26428 9240 26462
rect 9274 26428 9308 26462
rect 9342 26428 9376 26462
rect 9410 26428 9444 26462
rect 9478 26428 9512 26462
rect 9546 26428 9580 26462
rect 9614 26428 9648 26462
rect 9682 26428 9716 26462
rect 9750 26428 9784 26462
rect 9818 26428 9852 26462
rect 9886 26428 9920 26462
rect 9954 26428 9988 26462
rect 10022 26428 10056 26462
rect 10090 26428 10124 26462
rect 10158 26428 10192 26462
rect 10226 26428 10260 26462
rect 10294 26428 10328 26462
rect 10362 26428 10396 26462
rect 10430 26428 10464 26462
rect 10498 26428 10532 26462
rect 10566 26428 10600 26462
rect 10634 26428 10668 26462
rect 10702 26428 10736 26462
rect 10770 26428 10804 26462
rect 10838 26428 10872 26462
rect 10906 26428 10940 26462
rect 10974 26428 11008 26462
rect 11042 26428 11076 26462
rect 11110 26428 11144 26462
rect 11178 26428 11212 26462
rect 11246 26428 11280 26462
rect 11314 26428 11348 26462
rect 11382 26428 11416 26462
rect 11450 26428 11484 26462
rect 11518 26428 11552 26462
rect 11586 26428 11620 26462
rect 11654 26428 11688 26462
rect 11722 26428 11756 26462
rect 11790 26428 11824 26462
rect 11858 26428 11892 26462
rect 11926 26428 11960 26462
rect 11994 26428 12028 26462
rect 12062 26428 12096 26462
rect 12130 26428 12164 26462
rect 12198 26428 12232 26462
rect 12266 26428 12300 26462
rect 12334 26428 12368 26462
rect 12402 26428 12436 26462
rect 12470 26428 12504 26462
rect 12538 26428 12572 26462
rect 12606 26428 12640 26462
rect 12674 26428 12708 26462
rect 12742 26428 12776 26462
rect 12810 26428 12844 26462
rect 12878 26428 12912 26462
rect 12946 26428 12980 26462
rect 13014 26428 13048 26462
rect 13082 26428 13116 26462
rect 13150 26428 13184 26462
rect 13218 26428 13252 26462
rect 13286 26428 13320 26462
rect 13354 26428 13388 26462
rect 13422 26428 13456 26462
rect 13490 26428 13524 26462
rect 13558 26428 13592 26462
rect 13626 26428 13660 26462
rect 13694 26428 13728 26462
rect 13762 26428 13796 26462
rect 13830 26428 13864 26462
rect 13898 26428 13932 26462
rect 13966 26428 14000 26462
rect 14034 26428 14068 26462
rect 14102 26428 14136 26462
rect 14170 26428 14204 26462
rect 14238 26428 14272 26462
rect 14306 26428 14340 26462
rect 14374 26428 14408 26462
rect 14442 26428 14476 26462
rect 14510 26428 14544 26462
rect 14578 26428 14612 26462
rect 14646 26428 14680 26462
rect 14714 26428 14748 26462
rect 14782 26428 14816 26462
rect 14850 26428 14884 26462
rect 14918 26428 14962 26462
rect 2796 26427 14962 26428
rect 49 26351 14962 26427
rect 49 26317 83 26351
rect 117 26317 152 26351
rect 186 26317 221 26351
rect 255 26317 290 26351
rect 324 26317 359 26351
rect 393 26317 428 26351
rect 462 26317 497 26351
rect 531 26317 566 26351
rect 600 26317 635 26351
rect 669 26317 704 26351
rect 738 26317 773 26351
rect 807 26317 842 26351
rect 876 26317 911 26351
rect 945 26317 980 26351
rect 1014 26317 1049 26351
rect 1083 26317 1118 26351
rect 1152 26317 1187 26351
rect 1221 26317 1256 26351
rect 1290 26317 1325 26351
rect 1359 26317 1394 26351
rect 1428 26317 1463 26351
rect 1497 26317 1532 26351
rect 1566 26317 1601 26351
rect 1635 26317 1670 26351
rect 1704 26317 1739 26351
rect 1773 26317 1808 26351
rect 1842 26317 1877 26351
rect 1911 26317 1946 26351
rect 1980 26317 2015 26351
rect 2049 26317 2084 26351
rect 2118 26317 2153 26351
rect 2187 26317 2222 26351
rect 2256 26317 2291 26351
rect 2325 26317 2360 26351
rect 2394 26317 2429 26351
rect 2463 26317 2498 26351
rect 2532 26317 2567 26351
rect 2601 26317 2636 26351
rect 2670 26317 2705 26351
rect 2739 26317 2774 26351
rect 2808 26317 2843 26351
rect 2877 26317 2912 26351
rect 2946 26317 2981 26351
rect 3015 26317 3050 26351
rect 3084 26317 3119 26351
rect 3153 26317 3188 26351
rect 3222 26317 3256 26351
rect 3290 26317 3324 26351
rect 3358 26317 3392 26351
rect 3426 26317 3460 26351
rect 3494 26317 3528 26351
rect 3562 26317 3596 26351
rect 3630 26317 3664 26351
rect 3698 26317 3732 26351
rect 3766 26317 3800 26351
rect 3834 26317 3868 26351
rect 3902 26317 3936 26351
rect 3970 26317 4004 26351
rect 4038 26317 4072 26351
rect 4106 26317 4140 26351
rect 4174 26317 4208 26351
rect 4242 26317 4276 26351
rect 4310 26317 4344 26351
rect 4378 26317 4412 26351
rect 4446 26317 4480 26351
rect 4514 26317 4548 26351
rect 4582 26317 4616 26351
rect 4650 26317 4684 26351
rect 4718 26317 4752 26351
rect 4786 26317 4820 26351
rect 4854 26317 4888 26351
rect 4922 26317 4956 26351
rect 4990 26317 5024 26351
rect 5058 26317 5092 26351
rect 5126 26317 5160 26351
rect 5194 26317 5228 26351
rect 5262 26317 5296 26351
rect 5330 26317 5364 26351
rect 5398 26317 5432 26351
rect 5466 26317 5500 26351
rect 5534 26317 5568 26351
rect 5602 26317 5636 26351
rect 5670 26317 5704 26351
rect 5738 26317 5772 26351
rect 5806 26317 5840 26351
rect 5874 26317 5908 26351
rect 5942 26317 5976 26351
rect 6010 26317 6044 26351
rect 6078 26317 6112 26351
rect 6146 26317 6180 26351
rect 6214 26317 6248 26351
rect 6282 26317 6316 26351
rect 6350 26317 6384 26351
rect 6418 26317 6452 26351
rect 6486 26317 6520 26351
rect 6554 26317 6588 26351
rect 6622 26317 6656 26351
rect 6690 26317 6724 26351
rect 6758 26317 6792 26351
rect 6826 26317 6860 26351
rect 6894 26317 6928 26351
rect 6962 26317 6996 26351
rect 7030 26317 7064 26351
rect 7098 26317 7132 26351
rect 7166 26317 7200 26351
rect 7234 26317 7268 26351
rect 7302 26317 7336 26351
rect 7370 26317 7404 26351
rect 7438 26317 7472 26351
rect 7506 26317 7540 26351
rect 7574 26317 7608 26351
rect 7642 26317 7676 26351
rect 7710 26317 7744 26351
rect 7778 26317 7812 26351
rect 7846 26317 7880 26351
rect 7914 26317 7948 26351
rect 7982 26317 8016 26351
rect 8050 26317 8084 26351
rect 8118 26317 8152 26351
rect 8186 26317 8220 26351
rect 8254 26317 8288 26351
rect 8322 26317 8356 26351
rect 8390 26317 8424 26351
rect 8458 26317 8492 26351
rect 8526 26317 8560 26351
rect 8594 26317 8628 26351
rect 8662 26317 8696 26351
rect 8730 26317 8764 26351
rect 8798 26317 8832 26351
rect 8866 26317 8900 26351
rect 8934 26317 8968 26351
rect 9002 26317 9036 26351
rect 9070 26317 9104 26351
rect 9138 26317 9172 26351
rect 9206 26317 9240 26351
rect 9274 26317 9308 26351
rect 9342 26317 9376 26351
rect 9410 26317 9444 26351
rect 9478 26317 9512 26351
rect 9546 26317 9580 26351
rect 9614 26317 9648 26351
rect 9682 26317 9716 26351
rect 9750 26317 9784 26351
rect 9818 26317 9852 26351
rect 9886 26317 9920 26351
rect 9954 26317 9988 26351
rect 10022 26317 10056 26351
rect 10090 26317 10124 26351
rect 10158 26317 10192 26351
rect 10226 26317 10260 26351
rect 10294 26317 10328 26351
rect 10362 26317 10396 26351
rect 10430 26317 10464 26351
rect 10498 26317 10532 26351
rect 10566 26317 10600 26351
rect 10634 26317 10668 26351
rect 10702 26317 10736 26351
rect 10770 26317 10804 26351
rect 10838 26317 10872 26351
rect 10906 26317 10940 26351
rect 10974 26317 11008 26351
rect 11042 26317 11076 26351
rect 11110 26317 11144 26351
rect 11178 26317 11212 26351
rect 11246 26317 11280 26351
rect 11314 26317 11348 26351
rect 11382 26317 11416 26351
rect 11450 26317 11484 26351
rect 11518 26317 11552 26351
rect 11586 26317 11620 26351
rect 11654 26317 11688 26351
rect 11722 26317 11756 26351
rect 11790 26317 11824 26351
rect 11858 26317 11892 26351
rect 11926 26317 11960 26351
rect 11994 26317 12028 26351
rect 12062 26317 12096 26351
rect 12130 26317 12164 26351
rect 12198 26317 12232 26351
rect 12266 26317 12300 26351
rect 12334 26317 12368 26351
rect 12402 26317 12436 26351
rect 12470 26317 12504 26351
rect 12538 26317 12572 26351
rect 12606 26317 12640 26351
rect 12674 26317 12708 26351
rect 12742 26317 12776 26351
rect 12810 26317 12844 26351
rect 12878 26317 12912 26351
rect 12946 26317 12980 26351
rect 13014 26317 13048 26351
rect 13082 26317 13116 26351
rect 13150 26317 13184 26351
rect 13218 26317 13252 26351
rect 13286 26317 13320 26351
rect 13354 26317 13388 26351
rect 13422 26317 13456 26351
rect 13490 26317 13524 26351
rect 13558 26317 13592 26351
rect 13626 26317 13660 26351
rect 13694 26317 13728 26351
rect 13762 26317 13796 26351
rect 13830 26317 13864 26351
rect 13898 26317 13932 26351
rect 13966 26317 14000 26351
rect 14034 26317 14068 26351
rect 14102 26317 14136 26351
rect 14170 26317 14204 26351
rect 14238 26317 14272 26351
rect 14306 26317 14340 26351
rect 14374 26317 14408 26351
rect 14442 26317 14476 26351
rect 14510 26317 14544 26351
rect 14578 26317 14612 26351
rect 14646 26317 14680 26351
rect 14714 26317 14748 26351
rect 14782 26317 14816 26351
rect 14850 26317 14884 26351
rect 14918 26317 14962 26351
rect 49 26244 14962 26317
rect 49 26210 69 26244
rect 103 26210 138 26244
rect 172 26210 207 26244
rect 241 26210 276 26244
rect 310 26210 345 26244
rect 379 26210 414 26244
rect 448 26210 483 26244
rect 517 26210 552 26244
rect 586 26210 621 26244
rect 655 26210 690 26244
rect 724 26210 759 26244
rect 793 26210 828 26244
rect 862 26210 897 26244
rect 931 26210 966 26244
rect 1000 26210 1035 26244
rect 1069 26210 1104 26244
rect 1138 26210 1173 26244
rect 1207 26210 1242 26244
rect 1276 26210 1311 26244
rect 1345 26210 1380 26244
rect 1414 26210 1449 26244
rect 1483 26210 1518 26244
rect 1552 26210 1587 26244
rect 1621 26210 1656 26244
rect 1690 26210 1725 26244
rect 1759 26210 1794 26244
rect 1828 26210 1863 26244
rect 1897 26210 1932 26244
rect 1966 26210 2001 26244
rect 2035 26210 2070 26244
rect 2104 26210 2139 26244
rect 2173 26210 2208 26244
rect 2242 26210 2277 26244
rect 2311 26210 2346 26244
rect 2380 26210 2415 26244
rect 2449 26210 2484 26244
rect 2518 26210 2553 26244
rect 2587 26210 2622 26244
rect 2656 26210 2691 26244
rect 2725 26210 2760 26244
rect 2794 26210 2829 26244
rect 2863 26210 2898 26244
rect 2932 26210 2967 26244
rect 3001 26210 3036 26244
rect 3070 26210 3105 26244
rect 3139 26210 3174 26244
rect 3208 26210 3243 26244
rect 3277 26210 3312 26244
rect 3346 26210 3381 26244
rect 3415 26210 3450 26244
rect 3484 26210 3519 26244
rect 3553 26210 3588 26244
rect 3622 26210 3657 26244
rect 3691 26210 3726 26244
rect 3760 26210 3795 26244
rect 3829 26210 3864 26244
rect 3898 26210 3933 26244
rect 3967 26210 4002 26244
rect 4036 26210 4071 26244
rect 4105 26210 4140 26244
rect 4174 26210 4208 26244
rect 4242 26210 4276 26244
rect 4310 26210 4344 26244
rect 4378 26210 4412 26244
rect 4446 26210 4480 26244
rect 4514 26210 4548 26244
rect 4582 26210 4616 26244
rect 4650 26210 4684 26244
rect 4718 26210 4752 26244
rect 4786 26210 4820 26244
rect 4854 26210 4888 26244
rect 4922 26210 4956 26244
rect 4990 26210 5024 26244
rect 5058 26210 5092 26244
rect 5126 26210 5160 26244
rect 5194 26210 5228 26244
rect 5262 26210 5296 26244
rect 5330 26210 5364 26244
rect 5398 26210 5432 26244
rect 5466 26210 5500 26244
rect 5534 26210 5568 26244
rect 5602 26210 5636 26244
rect 5670 26210 5704 26244
rect 5738 26210 5772 26244
rect 5806 26210 5840 26244
rect 5874 26210 5908 26244
rect 5942 26210 5976 26244
rect 6010 26210 6044 26244
rect 6078 26210 6112 26244
rect 6146 26210 6180 26244
rect 6214 26210 6248 26244
rect 6282 26210 6316 26244
rect 6350 26210 6384 26244
rect 6418 26210 6452 26244
rect 6486 26210 6520 26244
rect 6554 26210 6588 26244
rect 6622 26210 6656 26244
rect 6690 26210 6724 26244
rect 6758 26210 6792 26244
rect 6826 26210 6860 26244
rect 6894 26210 6928 26244
rect 6962 26210 6996 26244
rect 7030 26210 7064 26244
rect 7098 26210 7132 26244
rect 7166 26210 7200 26244
rect 7234 26210 7268 26244
rect 7302 26210 7336 26244
rect 7370 26210 7404 26244
rect 7438 26210 7472 26244
rect 7506 26210 7540 26244
rect 7574 26210 7608 26244
rect 7642 26210 7676 26244
rect 7710 26210 7744 26244
rect 7778 26210 7812 26244
rect 7846 26210 7880 26244
rect 7914 26210 7948 26244
rect 7982 26210 8016 26244
rect 8050 26210 8084 26244
rect 8118 26210 8152 26244
rect 8186 26210 8220 26244
rect 8254 26210 8288 26244
rect 8322 26210 8356 26244
rect 8390 26210 8424 26244
rect 8458 26210 8492 26244
rect 8526 26210 8560 26244
rect 8594 26210 8628 26244
rect 8662 26210 8696 26244
rect 8730 26210 8764 26244
rect 8798 26210 8832 26244
rect 8866 26210 8900 26244
rect 8934 26210 8968 26244
rect 9002 26210 9036 26244
rect 9070 26210 9104 26244
rect 9138 26210 9172 26244
rect 9206 26210 9240 26244
rect 9274 26210 9308 26244
rect 9342 26210 9376 26244
rect 9410 26210 9444 26244
rect 9478 26210 9512 26244
rect 9546 26210 9580 26244
rect 9614 26210 9648 26244
rect 9682 26210 9716 26244
rect 9750 26210 9784 26244
rect 9818 26210 9852 26244
rect 9886 26210 9920 26244
rect 9954 26210 9988 26244
rect 10022 26210 10056 26244
rect 10090 26210 10124 26244
rect 10158 26210 10192 26244
rect 10226 26210 10260 26244
rect 10294 26210 10328 26244
rect 10362 26210 10396 26244
rect 10430 26210 10464 26244
rect 10498 26210 10532 26244
rect 10566 26210 10600 26244
rect 10634 26210 10668 26244
rect 10702 26210 10736 26244
rect 10770 26210 10804 26244
rect 10838 26210 10872 26244
rect 10906 26210 10940 26244
rect 10974 26210 11008 26244
rect 11042 26210 11076 26244
rect 11110 26210 11144 26244
rect 11178 26210 11212 26244
rect 11246 26210 11280 26244
rect 11314 26210 11348 26244
rect 11382 26210 11416 26244
rect 11450 26210 11484 26244
rect 11518 26210 11552 26244
rect 11586 26210 11620 26244
rect 11654 26210 11688 26244
rect 11722 26210 11756 26244
rect 11790 26210 11824 26244
rect 11858 26210 11892 26244
rect 11926 26210 11960 26244
rect 11994 26210 12028 26244
rect 12062 26210 12096 26244
rect 12130 26210 12164 26244
rect 12198 26210 12232 26244
rect 12266 26210 12300 26244
rect 12334 26210 12368 26244
rect 12402 26210 12436 26244
rect 12470 26210 12504 26244
rect 12538 26210 12572 26244
rect 12606 26210 12640 26244
rect 12674 26210 12708 26244
rect 12742 26210 12776 26244
rect 12810 26210 12844 26244
rect 12878 26210 12912 26244
rect 12946 26210 12980 26244
rect 13014 26210 13048 26244
rect 13082 26210 13116 26244
rect 13150 26210 13184 26244
rect 13218 26210 13252 26244
rect 13286 26210 13320 26244
rect 13354 26210 13388 26244
rect 13422 26210 13456 26244
rect 13490 26210 13524 26244
rect 13558 26210 13592 26244
rect 13626 26210 13660 26244
rect 13694 26210 13728 26244
rect 13762 26210 13796 26244
rect 13830 26210 13864 26244
rect 13898 26210 13932 26244
rect 13966 26210 14000 26244
rect 14034 26210 14068 26244
rect 14102 26210 14136 26244
rect 14170 26210 14204 26244
rect 14238 26210 14272 26244
rect 14306 26210 14340 26244
rect 14374 26210 14408 26244
rect 14442 26210 14476 26244
rect 14510 26210 14544 26244
rect 14578 26210 14612 26244
rect 14646 26210 14680 26244
rect 14714 26210 14748 26244
rect 14782 26210 14816 26244
rect 14850 26210 14884 26244
rect 14918 26210 14962 26244
rect 49 26185 14962 26210
rect 49 26172 243 26185
rect 277 26172 316 26185
rect 350 26172 389 26185
rect 423 26172 462 26185
rect 496 26172 535 26185
rect 569 26172 608 26185
rect 642 26172 681 26185
rect 715 26172 754 26185
rect 788 26172 827 26185
rect 861 26172 900 26185
rect 934 26172 973 26185
rect 1007 26172 1046 26185
rect 1080 26172 1119 26185
rect 1153 26172 1192 26185
rect 1226 26172 1265 26185
rect 1299 26172 1338 26185
rect 1372 26172 1411 26185
rect 1445 26172 1484 26185
rect 49 26138 69 26172
rect 103 26138 138 26172
rect 172 26138 207 26172
rect 241 26151 243 26172
rect 310 26151 316 26172
rect 379 26151 389 26172
rect 448 26151 462 26172
rect 517 26151 535 26172
rect 586 26151 608 26172
rect 655 26151 681 26172
rect 724 26151 754 26172
rect 793 26151 827 26172
rect 241 26138 276 26151
rect 310 26138 345 26151
rect 379 26138 414 26151
rect 448 26138 483 26151
rect 517 26138 552 26151
rect 586 26138 621 26151
rect 655 26138 690 26151
rect 724 26138 759 26151
rect 793 26138 828 26151
rect 862 26138 897 26172
rect 934 26151 966 26172
rect 1007 26151 1035 26172
rect 1080 26151 1104 26172
rect 1153 26151 1173 26172
rect 1226 26151 1242 26172
rect 1299 26151 1311 26172
rect 1372 26151 1380 26172
rect 1445 26151 1449 26172
rect 931 26138 966 26151
rect 1000 26138 1035 26151
rect 1069 26138 1104 26151
rect 1138 26138 1173 26151
rect 1207 26138 1242 26151
rect 1276 26138 1311 26151
rect 1345 26138 1380 26151
rect 1414 26138 1449 26151
rect 1483 26151 1484 26172
rect 1518 26172 1557 26185
rect 1591 26172 1630 26185
rect 1664 26172 1703 26185
rect 1737 26172 1776 26185
rect 1810 26172 1849 26185
rect 1883 26172 1922 26185
rect 1956 26172 1995 26185
rect 2029 26172 2068 26185
rect 2102 26172 2141 26185
rect 2175 26172 2214 26185
rect 2248 26172 2287 26185
rect 2321 26172 2360 26185
rect 2394 26172 2433 26185
rect 2467 26172 2506 26185
rect 2540 26172 2579 26185
rect 2613 26172 2652 26185
rect 2686 26172 2725 26185
rect 1483 26138 1518 26151
rect 1552 26151 1557 26172
rect 1621 26151 1630 26172
rect 1690 26151 1703 26172
rect 1759 26151 1776 26172
rect 1828 26151 1849 26172
rect 1897 26151 1922 26172
rect 1966 26151 1995 26172
rect 2035 26151 2068 26172
rect 1552 26138 1587 26151
rect 1621 26138 1656 26151
rect 1690 26138 1725 26151
rect 1759 26138 1794 26151
rect 1828 26138 1863 26151
rect 1897 26138 1932 26151
rect 1966 26138 2001 26151
rect 2035 26138 2070 26151
rect 2104 26138 2139 26172
rect 2175 26151 2208 26172
rect 2248 26151 2277 26172
rect 2321 26151 2346 26172
rect 2394 26151 2415 26172
rect 2467 26151 2484 26172
rect 2540 26151 2553 26172
rect 2613 26151 2622 26172
rect 2686 26151 2691 26172
rect 2173 26138 2208 26151
rect 2242 26138 2277 26151
rect 2311 26138 2346 26151
rect 2380 26138 2415 26151
rect 2449 26138 2484 26151
rect 2518 26138 2553 26151
rect 2587 26138 2622 26151
rect 2656 26138 2691 26151
rect 2759 26172 2798 26185
rect 2832 26172 2871 26185
rect 2905 26172 2944 26185
rect 2978 26172 3017 26185
rect 3051 26172 3090 26185
rect 3124 26172 3163 26185
rect 3197 26172 3236 26185
rect 3270 26172 3309 26185
rect 3343 26172 3382 26185
rect 3416 26172 3455 26185
rect 3489 26172 3528 26185
rect 3562 26172 3601 26185
rect 3635 26172 3674 26185
rect 3708 26172 3746 26185
rect 3780 26172 3818 26185
rect 3852 26172 3890 26185
rect 3924 26172 3962 26185
rect 3996 26172 4034 26185
rect 4068 26172 4106 26185
rect 2759 26151 2760 26172
rect 2725 26138 2760 26151
rect 2794 26151 2798 26172
rect 2863 26151 2871 26172
rect 2932 26151 2944 26172
rect 3001 26151 3017 26172
rect 3070 26151 3090 26172
rect 3139 26151 3163 26172
rect 3208 26151 3236 26172
rect 3277 26151 3309 26172
rect 2794 26138 2829 26151
rect 2863 26138 2898 26151
rect 2932 26138 2967 26151
rect 3001 26138 3036 26151
rect 3070 26138 3105 26151
rect 3139 26138 3174 26151
rect 3208 26138 3243 26151
rect 3277 26138 3312 26151
rect 3346 26138 3381 26172
rect 3416 26151 3450 26172
rect 3489 26151 3519 26172
rect 3562 26151 3588 26172
rect 3635 26151 3657 26172
rect 3708 26151 3726 26172
rect 3780 26151 3795 26172
rect 3852 26151 3864 26172
rect 3924 26151 3933 26172
rect 3996 26151 4002 26172
rect 4068 26151 4071 26172
rect 3415 26138 3450 26151
rect 3484 26138 3519 26151
rect 3553 26138 3588 26151
rect 3622 26138 3657 26151
rect 3691 26138 3726 26151
rect 3760 26138 3795 26151
rect 3829 26138 3864 26151
rect 3898 26138 3933 26151
rect 3967 26138 4002 26151
rect 4036 26138 4071 26151
rect 4105 26151 4106 26172
rect 4140 26172 4178 26185
rect 4212 26172 4250 26185
rect 4284 26172 4322 26185
rect 4356 26172 4394 26185
rect 4428 26172 4466 26185
rect 4500 26172 4538 26185
rect 4572 26172 4610 26185
rect 4644 26172 4682 26185
rect 4716 26172 4754 26185
rect 4788 26172 4826 26185
rect 4860 26172 4898 26185
rect 4932 26172 4970 26185
rect 5004 26172 5042 26185
rect 5076 26172 5114 26185
rect 5148 26172 5186 26185
rect 5220 26172 5258 26185
rect 5292 26172 5330 26185
rect 4105 26138 4140 26151
rect 4174 26151 4178 26172
rect 4242 26151 4250 26172
rect 4310 26151 4322 26172
rect 4378 26151 4394 26172
rect 4446 26151 4466 26172
rect 4514 26151 4538 26172
rect 4582 26151 4610 26172
rect 4650 26151 4682 26172
rect 4174 26138 4208 26151
rect 4242 26138 4276 26151
rect 4310 26138 4344 26151
rect 4378 26138 4412 26151
rect 4446 26138 4480 26151
rect 4514 26138 4548 26151
rect 4582 26138 4616 26151
rect 4650 26138 4684 26151
rect 4718 26138 4752 26172
rect 4788 26151 4820 26172
rect 4860 26151 4888 26172
rect 4932 26151 4956 26172
rect 5004 26151 5024 26172
rect 5076 26151 5092 26172
rect 5148 26151 5160 26172
rect 5220 26151 5228 26172
rect 5292 26151 5296 26172
rect 4786 26138 4820 26151
rect 4854 26138 4888 26151
rect 4922 26138 4956 26151
rect 4990 26138 5024 26151
rect 5058 26138 5092 26151
rect 5126 26138 5160 26151
rect 5194 26138 5228 26151
rect 5262 26138 5296 26151
rect 5364 26172 5402 26185
rect 5436 26172 5474 26185
rect 5508 26172 5546 26185
rect 5580 26172 5618 26185
rect 5652 26172 5690 26185
rect 5724 26172 5762 26185
rect 5796 26172 5834 26185
rect 5868 26172 5906 26185
rect 5940 26172 5978 26185
rect 6012 26172 6050 26185
rect 6084 26172 6122 26185
rect 6156 26172 6194 26185
rect 6228 26172 6266 26185
rect 6300 26172 6338 26185
rect 6372 26172 6410 26185
rect 6444 26172 6482 26185
rect 6516 26172 6554 26185
rect 5330 26138 5364 26151
rect 5398 26151 5402 26172
rect 5466 26151 5474 26172
rect 5534 26151 5546 26172
rect 5602 26151 5618 26172
rect 5670 26151 5690 26172
rect 5738 26151 5762 26172
rect 5806 26151 5834 26172
rect 5874 26151 5906 26172
rect 5398 26138 5432 26151
rect 5466 26138 5500 26151
rect 5534 26138 5568 26151
rect 5602 26138 5636 26151
rect 5670 26138 5704 26151
rect 5738 26138 5772 26151
rect 5806 26138 5840 26151
rect 5874 26138 5908 26151
rect 5942 26138 5976 26172
rect 6012 26151 6044 26172
rect 6084 26151 6112 26172
rect 6156 26151 6180 26172
rect 6228 26151 6248 26172
rect 6300 26151 6316 26172
rect 6372 26151 6384 26172
rect 6444 26151 6452 26172
rect 6516 26151 6520 26172
rect 6010 26138 6044 26151
rect 6078 26138 6112 26151
rect 6146 26138 6180 26151
rect 6214 26138 6248 26151
rect 6282 26138 6316 26151
rect 6350 26138 6384 26151
rect 6418 26138 6452 26151
rect 6486 26138 6520 26151
rect 6588 26172 6626 26185
rect 6660 26172 6698 26185
rect 6732 26172 6770 26185
rect 6804 26172 6842 26185
rect 6876 26172 6914 26185
rect 6948 26172 6986 26185
rect 7020 26172 7058 26185
rect 7092 26172 7130 26185
rect 7164 26172 7202 26185
rect 7236 26172 7274 26185
rect 7308 26172 7346 26185
rect 7380 26172 7418 26185
rect 7452 26172 7490 26185
rect 7524 26172 7562 26185
rect 7596 26172 7634 26185
rect 7668 26172 7706 26185
rect 7740 26172 7778 26185
rect 6554 26138 6588 26151
rect 6622 26151 6626 26172
rect 6690 26151 6698 26172
rect 6758 26151 6770 26172
rect 6826 26151 6842 26172
rect 6894 26151 6914 26172
rect 6962 26151 6986 26172
rect 7030 26151 7058 26172
rect 7098 26151 7130 26172
rect 6622 26138 6656 26151
rect 6690 26138 6724 26151
rect 6758 26138 6792 26151
rect 6826 26138 6860 26151
rect 6894 26138 6928 26151
rect 6962 26138 6996 26151
rect 7030 26138 7064 26151
rect 7098 26138 7132 26151
rect 7166 26138 7200 26172
rect 7236 26151 7268 26172
rect 7308 26151 7336 26172
rect 7380 26151 7404 26172
rect 7452 26151 7472 26172
rect 7524 26151 7540 26172
rect 7596 26151 7608 26172
rect 7668 26151 7676 26172
rect 7740 26151 7744 26172
rect 7234 26138 7268 26151
rect 7302 26138 7336 26151
rect 7370 26138 7404 26151
rect 7438 26138 7472 26151
rect 7506 26138 7540 26151
rect 7574 26138 7608 26151
rect 7642 26138 7676 26151
rect 7710 26138 7744 26151
rect 7812 26172 7850 26185
rect 7884 26172 7922 26185
rect 7956 26172 7994 26185
rect 8028 26172 8066 26185
rect 8100 26172 8138 26185
rect 8172 26172 8210 26185
rect 8244 26172 8282 26185
rect 8316 26172 8354 26185
rect 8388 26172 8426 26185
rect 8460 26172 8498 26185
rect 8532 26172 8570 26185
rect 8604 26172 8642 26185
rect 8676 26172 8714 26185
rect 8748 26172 8786 26185
rect 8820 26172 8858 26185
rect 8892 26172 8930 26185
rect 8964 26172 9002 26185
rect 7778 26138 7812 26151
rect 7846 26151 7850 26172
rect 7914 26151 7922 26172
rect 7982 26151 7994 26172
rect 8050 26151 8066 26172
rect 8118 26151 8138 26172
rect 8186 26151 8210 26172
rect 8254 26151 8282 26172
rect 8322 26151 8354 26172
rect 7846 26138 7880 26151
rect 7914 26138 7948 26151
rect 7982 26138 8016 26151
rect 8050 26138 8084 26151
rect 8118 26138 8152 26151
rect 8186 26138 8220 26151
rect 8254 26138 8288 26151
rect 8322 26138 8356 26151
rect 8390 26138 8424 26172
rect 8460 26151 8492 26172
rect 8532 26151 8560 26172
rect 8604 26151 8628 26172
rect 8676 26151 8696 26172
rect 8748 26151 8764 26172
rect 8820 26151 8832 26172
rect 8892 26151 8900 26172
rect 8964 26151 8968 26172
rect 8458 26138 8492 26151
rect 8526 26138 8560 26151
rect 8594 26138 8628 26151
rect 8662 26138 8696 26151
rect 8730 26138 8764 26151
rect 8798 26138 8832 26151
rect 8866 26138 8900 26151
rect 8934 26138 8968 26151
rect 9036 26172 9074 26185
rect 9108 26172 9146 26185
rect 9180 26172 9218 26185
rect 9252 26172 9290 26185
rect 9324 26172 9362 26185
rect 9396 26172 9434 26185
rect 9468 26172 9506 26185
rect 9540 26172 9578 26185
rect 9612 26172 9650 26185
rect 9684 26172 9722 26185
rect 9756 26172 9794 26185
rect 9828 26172 9866 26185
rect 9900 26172 9938 26185
rect 9972 26172 10010 26185
rect 10044 26172 10082 26185
rect 10116 26172 10154 26185
rect 10188 26172 10226 26185
rect 9002 26138 9036 26151
rect 9070 26151 9074 26172
rect 9138 26151 9146 26172
rect 9206 26151 9218 26172
rect 9274 26151 9290 26172
rect 9342 26151 9362 26172
rect 9410 26151 9434 26172
rect 9478 26151 9506 26172
rect 9546 26151 9578 26172
rect 9070 26138 9104 26151
rect 9138 26138 9172 26151
rect 9206 26138 9240 26151
rect 9274 26138 9308 26151
rect 9342 26138 9376 26151
rect 9410 26138 9444 26151
rect 9478 26138 9512 26151
rect 9546 26138 9580 26151
rect 9614 26138 9648 26172
rect 9684 26151 9716 26172
rect 9756 26151 9784 26172
rect 9828 26151 9852 26172
rect 9900 26151 9920 26172
rect 9972 26151 9988 26172
rect 10044 26151 10056 26172
rect 10116 26151 10124 26172
rect 10188 26151 10192 26172
rect 9682 26138 9716 26151
rect 9750 26138 9784 26151
rect 9818 26138 9852 26151
rect 9886 26138 9920 26151
rect 9954 26138 9988 26151
rect 10022 26138 10056 26151
rect 10090 26138 10124 26151
rect 10158 26138 10192 26151
rect 10260 26172 10298 26185
rect 10332 26172 10370 26185
rect 10404 26172 10442 26185
rect 10476 26172 10514 26185
rect 10548 26172 10586 26185
rect 10620 26172 10658 26185
rect 10692 26172 10730 26185
rect 10764 26172 10802 26185
rect 10836 26172 10874 26185
rect 10908 26172 10946 26185
rect 10980 26172 11018 26185
rect 11052 26172 11090 26185
rect 11124 26172 11162 26185
rect 11196 26172 11234 26185
rect 11268 26172 11306 26185
rect 11340 26172 11378 26185
rect 11412 26172 11450 26185
rect 10226 26138 10260 26151
rect 10294 26151 10298 26172
rect 10362 26151 10370 26172
rect 10430 26151 10442 26172
rect 10498 26151 10514 26172
rect 10566 26151 10586 26172
rect 10634 26151 10658 26172
rect 10702 26151 10730 26172
rect 10770 26151 10802 26172
rect 10294 26138 10328 26151
rect 10362 26138 10396 26151
rect 10430 26138 10464 26151
rect 10498 26138 10532 26151
rect 10566 26138 10600 26151
rect 10634 26138 10668 26151
rect 10702 26138 10736 26151
rect 10770 26138 10804 26151
rect 10838 26138 10872 26172
rect 10908 26151 10940 26172
rect 10980 26151 11008 26172
rect 11052 26151 11076 26172
rect 11124 26151 11144 26172
rect 11196 26151 11212 26172
rect 11268 26151 11280 26172
rect 11340 26151 11348 26172
rect 11412 26151 11416 26172
rect 10906 26138 10940 26151
rect 10974 26138 11008 26151
rect 11042 26138 11076 26151
rect 11110 26138 11144 26151
rect 11178 26138 11212 26151
rect 11246 26138 11280 26151
rect 11314 26138 11348 26151
rect 11382 26138 11416 26151
rect 11484 26172 11522 26185
rect 11556 26172 11594 26185
rect 11628 26172 11666 26185
rect 11700 26172 11738 26185
rect 11772 26172 11810 26185
rect 11844 26172 11882 26185
rect 11916 26172 11954 26185
rect 11988 26172 12026 26185
rect 12060 26172 12098 26185
rect 12132 26172 12170 26185
rect 12204 26172 12242 26185
rect 12276 26172 12314 26185
rect 12348 26172 12386 26185
rect 12420 26172 12458 26185
rect 12492 26172 12530 26185
rect 12564 26172 12602 26185
rect 12636 26172 12674 26185
rect 11450 26138 11484 26151
rect 11518 26151 11522 26172
rect 11586 26151 11594 26172
rect 11654 26151 11666 26172
rect 11722 26151 11738 26172
rect 11790 26151 11810 26172
rect 11858 26151 11882 26172
rect 11926 26151 11954 26172
rect 11994 26151 12026 26172
rect 11518 26138 11552 26151
rect 11586 26138 11620 26151
rect 11654 26138 11688 26151
rect 11722 26138 11756 26151
rect 11790 26138 11824 26151
rect 11858 26138 11892 26151
rect 11926 26138 11960 26151
rect 11994 26138 12028 26151
rect 12062 26138 12096 26172
rect 12132 26151 12164 26172
rect 12204 26151 12232 26172
rect 12276 26151 12300 26172
rect 12348 26151 12368 26172
rect 12420 26151 12436 26172
rect 12492 26151 12504 26172
rect 12564 26151 12572 26172
rect 12636 26151 12640 26172
rect 12130 26138 12164 26151
rect 12198 26138 12232 26151
rect 12266 26138 12300 26151
rect 12334 26138 12368 26151
rect 12402 26138 12436 26151
rect 12470 26138 12504 26151
rect 12538 26138 12572 26151
rect 12606 26138 12640 26151
rect 12708 26172 12746 26185
rect 12780 26172 12818 26185
rect 12852 26172 12890 26185
rect 12924 26172 12962 26185
rect 12996 26172 13034 26185
rect 13068 26172 13106 26185
rect 13140 26172 13178 26185
rect 13212 26172 13250 26185
rect 13284 26172 13322 26185
rect 13356 26172 13394 26185
rect 13428 26172 13466 26185
rect 13500 26172 13538 26185
rect 13572 26172 13610 26185
rect 13644 26172 13682 26185
rect 13716 26172 13754 26185
rect 13788 26172 13826 26185
rect 13860 26172 13898 26185
rect 12674 26138 12708 26151
rect 12742 26151 12746 26172
rect 12810 26151 12818 26172
rect 12878 26151 12890 26172
rect 12946 26151 12962 26172
rect 13014 26151 13034 26172
rect 13082 26151 13106 26172
rect 13150 26151 13178 26172
rect 13218 26151 13250 26172
rect 12742 26138 12776 26151
rect 12810 26138 12844 26151
rect 12878 26138 12912 26151
rect 12946 26138 12980 26151
rect 13014 26138 13048 26151
rect 13082 26138 13116 26151
rect 13150 26138 13184 26151
rect 13218 26138 13252 26151
rect 13286 26138 13320 26172
rect 13356 26151 13388 26172
rect 13428 26151 13456 26172
rect 13500 26151 13524 26172
rect 13572 26151 13592 26172
rect 13644 26151 13660 26172
rect 13716 26151 13728 26172
rect 13788 26151 13796 26172
rect 13860 26151 13864 26172
rect 13354 26138 13388 26151
rect 13422 26138 13456 26151
rect 13490 26138 13524 26151
rect 13558 26138 13592 26151
rect 13626 26138 13660 26151
rect 13694 26138 13728 26151
rect 13762 26138 13796 26151
rect 13830 26138 13864 26151
rect 13932 26172 13970 26185
rect 14004 26172 14042 26185
rect 14076 26172 14114 26185
rect 14148 26172 14186 26185
rect 14220 26172 14258 26185
rect 14292 26172 14330 26185
rect 14364 26172 14402 26185
rect 14436 26172 14474 26185
rect 14508 26172 14546 26185
rect 14580 26172 14618 26185
rect 14652 26172 14690 26185
rect 14724 26172 14962 26185
rect 13898 26138 13932 26151
rect 13966 26151 13970 26172
rect 14034 26151 14042 26172
rect 14102 26151 14114 26172
rect 14170 26151 14186 26172
rect 14238 26151 14258 26172
rect 14306 26151 14330 26172
rect 14374 26151 14402 26172
rect 14442 26151 14474 26172
rect 13966 26138 14000 26151
rect 14034 26138 14068 26151
rect 14102 26138 14136 26151
rect 14170 26138 14204 26151
rect 14238 26138 14272 26151
rect 14306 26138 14340 26151
rect 14374 26138 14408 26151
rect 14442 26138 14476 26151
rect 14510 26138 14544 26172
rect 14580 26151 14612 26172
rect 14652 26151 14680 26172
rect 14724 26151 14748 26172
rect 14578 26138 14612 26151
rect 14646 26138 14680 26151
rect 14714 26138 14748 26151
rect 14782 26138 14816 26172
rect 14850 26138 14884 26172
rect 14918 26138 14962 26172
rect 49 26111 14962 26138
rect 49 26100 243 26111
rect 277 26100 316 26111
rect 350 26100 389 26111
rect 423 26100 462 26111
rect 496 26100 535 26111
rect 569 26100 608 26111
rect 642 26100 681 26111
rect 715 26100 754 26111
rect 788 26100 827 26111
rect 861 26100 900 26111
rect 934 26100 973 26111
rect 1007 26100 1046 26111
rect 1080 26100 1119 26111
rect 1153 26100 1192 26111
rect 1226 26100 1265 26111
rect 1299 26100 1338 26111
rect 1372 26100 1411 26111
rect 1445 26100 1484 26111
rect 49 26066 69 26100
rect 103 26066 138 26100
rect 172 26066 207 26100
rect 241 26077 243 26100
rect 310 26077 316 26100
rect 379 26077 389 26100
rect 448 26077 462 26100
rect 517 26077 535 26100
rect 586 26077 608 26100
rect 655 26077 681 26100
rect 724 26077 754 26100
rect 793 26077 827 26100
rect 241 26066 276 26077
rect 310 26066 345 26077
rect 379 26066 414 26077
rect 448 26066 483 26077
rect 517 26066 552 26077
rect 586 26066 621 26077
rect 655 26066 690 26077
rect 724 26066 759 26077
rect 793 26066 828 26077
rect 862 26066 897 26100
rect 934 26077 966 26100
rect 1007 26077 1035 26100
rect 1080 26077 1104 26100
rect 1153 26077 1173 26100
rect 1226 26077 1242 26100
rect 1299 26077 1311 26100
rect 1372 26077 1380 26100
rect 1445 26077 1449 26100
rect 931 26066 966 26077
rect 1000 26066 1035 26077
rect 1069 26066 1104 26077
rect 1138 26066 1173 26077
rect 1207 26066 1242 26077
rect 1276 26066 1311 26077
rect 1345 26066 1380 26077
rect 1414 26066 1449 26077
rect 1483 26077 1484 26100
rect 1518 26100 1557 26111
rect 1591 26100 1630 26111
rect 1664 26100 1703 26111
rect 1737 26100 1776 26111
rect 1810 26100 1849 26111
rect 1883 26100 1922 26111
rect 1956 26100 1995 26111
rect 2029 26100 2068 26111
rect 2102 26100 2141 26111
rect 2175 26100 2214 26111
rect 2248 26100 2287 26111
rect 2321 26100 2360 26111
rect 2394 26100 2433 26111
rect 2467 26100 2506 26111
rect 2540 26100 2579 26111
rect 2613 26100 2652 26111
rect 2686 26100 2725 26111
rect 1483 26066 1518 26077
rect 1552 26077 1557 26100
rect 1621 26077 1630 26100
rect 1690 26077 1703 26100
rect 1759 26077 1776 26100
rect 1828 26077 1849 26100
rect 1897 26077 1922 26100
rect 1966 26077 1995 26100
rect 2035 26077 2068 26100
rect 1552 26066 1587 26077
rect 1621 26066 1656 26077
rect 1690 26066 1725 26077
rect 1759 26066 1794 26077
rect 1828 26066 1863 26077
rect 1897 26066 1932 26077
rect 1966 26066 2001 26077
rect 2035 26066 2070 26077
rect 2104 26066 2139 26100
rect 2175 26077 2208 26100
rect 2248 26077 2277 26100
rect 2321 26077 2346 26100
rect 2394 26077 2415 26100
rect 2467 26077 2484 26100
rect 2540 26077 2553 26100
rect 2613 26077 2622 26100
rect 2686 26077 2691 26100
rect 2173 26066 2208 26077
rect 2242 26066 2277 26077
rect 2311 26066 2346 26077
rect 2380 26066 2415 26077
rect 2449 26066 2484 26077
rect 2518 26066 2553 26077
rect 2587 26066 2622 26077
rect 2656 26066 2691 26077
rect 2759 26100 2798 26111
rect 2832 26100 2871 26111
rect 2905 26100 2944 26111
rect 2978 26100 3017 26111
rect 3051 26100 3090 26111
rect 3124 26100 3163 26111
rect 3197 26100 3236 26111
rect 3270 26100 3309 26111
rect 3343 26100 3382 26111
rect 3416 26100 3455 26111
rect 3489 26100 3528 26111
rect 3562 26100 3601 26111
rect 3635 26100 3674 26111
rect 3708 26100 3746 26111
rect 3780 26100 3818 26111
rect 3852 26100 3890 26111
rect 3924 26100 3962 26111
rect 3996 26100 4034 26111
rect 4068 26100 4106 26111
rect 2759 26077 2760 26100
rect 2725 26066 2760 26077
rect 2794 26077 2798 26100
rect 2863 26077 2871 26100
rect 2932 26077 2944 26100
rect 3001 26077 3017 26100
rect 3070 26077 3090 26100
rect 3139 26077 3163 26100
rect 3208 26077 3236 26100
rect 3277 26077 3309 26100
rect 2794 26066 2829 26077
rect 2863 26066 2898 26077
rect 2932 26066 2967 26077
rect 3001 26066 3036 26077
rect 3070 26066 3105 26077
rect 3139 26066 3174 26077
rect 3208 26066 3243 26077
rect 3277 26066 3312 26077
rect 3346 26066 3381 26100
rect 3416 26077 3450 26100
rect 3489 26077 3519 26100
rect 3562 26077 3588 26100
rect 3635 26077 3657 26100
rect 3708 26077 3726 26100
rect 3780 26077 3795 26100
rect 3852 26077 3864 26100
rect 3924 26077 3933 26100
rect 3996 26077 4002 26100
rect 4068 26077 4071 26100
rect 3415 26066 3450 26077
rect 3484 26066 3519 26077
rect 3553 26066 3588 26077
rect 3622 26066 3657 26077
rect 3691 26066 3726 26077
rect 3760 26066 3795 26077
rect 3829 26066 3864 26077
rect 3898 26066 3933 26077
rect 3967 26066 4002 26077
rect 4036 26066 4071 26077
rect 4105 26077 4106 26100
rect 4140 26100 4178 26111
rect 4212 26100 4250 26111
rect 4284 26100 4322 26111
rect 4356 26100 4394 26111
rect 4428 26100 4466 26111
rect 4500 26100 4538 26111
rect 4572 26100 4610 26111
rect 4644 26100 4682 26111
rect 4716 26100 4754 26111
rect 4788 26100 4826 26111
rect 4860 26100 4898 26111
rect 4932 26100 4970 26111
rect 5004 26100 5042 26111
rect 5076 26100 5114 26111
rect 5148 26100 5186 26111
rect 5220 26100 5258 26111
rect 5292 26100 5330 26111
rect 4105 26066 4140 26077
rect 4174 26077 4178 26100
rect 4242 26077 4250 26100
rect 4310 26077 4322 26100
rect 4378 26077 4394 26100
rect 4446 26077 4466 26100
rect 4514 26077 4538 26100
rect 4582 26077 4610 26100
rect 4650 26077 4682 26100
rect 4174 26066 4208 26077
rect 4242 26066 4276 26077
rect 4310 26066 4344 26077
rect 4378 26066 4412 26077
rect 4446 26066 4480 26077
rect 4514 26066 4548 26077
rect 4582 26066 4616 26077
rect 4650 26066 4684 26077
rect 4718 26066 4752 26100
rect 4788 26077 4820 26100
rect 4860 26077 4888 26100
rect 4932 26077 4956 26100
rect 5004 26077 5024 26100
rect 5076 26077 5092 26100
rect 5148 26077 5160 26100
rect 5220 26077 5228 26100
rect 5292 26077 5296 26100
rect 4786 26066 4820 26077
rect 4854 26066 4888 26077
rect 4922 26066 4956 26077
rect 4990 26066 5024 26077
rect 5058 26066 5092 26077
rect 5126 26066 5160 26077
rect 5194 26066 5228 26077
rect 5262 26066 5296 26077
rect 5364 26100 5402 26111
rect 5436 26100 5474 26111
rect 5508 26100 5546 26111
rect 5580 26100 5618 26111
rect 5652 26100 5690 26111
rect 5724 26100 5762 26111
rect 5796 26100 5834 26111
rect 5868 26100 5906 26111
rect 5940 26100 5978 26111
rect 6012 26100 6050 26111
rect 6084 26100 6122 26111
rect 6156 26100 6194 26111
rect 6228 26100 6266 26111
rect 6300 26100 6338 26111
rect 6372 26100 6410 26111
rect 6444 26100 6482 26111
rect 6516 26100 6554 26111
rect 5330 26066 5364 26077
rect 5398 26077 5402 26100
rect 5466 26077 5474 26100
rect 5534 26077 5546 26100
rect 5602 26077 5618 26100
rect 5670 26077 5690 26100
rect 5738 26077 5762 26100
rect 5806 26077 5834 26100
rect 5874 26077 5906 26100
rect 5398 26066 5432 26077
rect 5466 26066 5500 26077
rect 5534 26066 5568 26077
rect 5602 26066 5636 26077
rect 5670 26066 5704 26077
rect 5738 26066 5772 26077
rect 5806 26066 5840 26077
rect 5874 26066 5908 26077
rect 5942 26066 5976 26100
rect 6012 26077 6044 26100
rect 6084 26077 6112 26100
rect 6156 26077 6180 26100
rect 6228 26077 6248 26100
rect 6300 26077 6316 26100
rect 6372 26077 6384 26100
rect 6444 26077 6452 26100
rect 6516 26077 6520 26100
rect 6010 26066 6044 26077
rect 6078 26066 6112 26077
rect 6146 26066 6180 26077
rect 6214 26066 6248 26077
rect 6282 26066 6316 26077
rect 6350 26066 6384 26077
rect 6418 26066 6452 26077
rect 6486 26066 6520 26077
rect 6588 26100 6626 26111
rect 6660 26100 6698 26111
rect 6732 26100 6770 26111
rect 6804 26100 6842 26111
rect 6876 26100 6914 26111
rect 6948 26100 6986 26111
rect 7020 26100 7058 26111
rect 7092 26100 7130 26111
rect 7164 26100 7202 26111
rect 7236 26100 7274 26111
rect 7308 26100 7346 26111
rect 7380 26100 7418 26111
rect 7452 26100 7490 26111
rect 7524 26100 7562 26111
rect 7596 26100 7634 26111
rect 7668 26100 7706 26111
rect 7740 26100 7778 26111
rect 6554 26066 6588 26077
rect 6622 26077 6626 26100
rect 6690 26077 6698 26100
rect 6758 26077 6770 26100
rect 6826 26077 6842 26100
rect 6894 26077 6914 26100
rect 6962 26077 6986 26100
rect 7030 26077 7058 26100
rect 7098 26077 7130 26100
rect 6622 26066 6656 26077
rect 6690 26066 6724 26077
rect 6758 26066 6792 26077
rect 6826 26066 6860 26077
rect 6894 26066 6928 26077
rect 6962 26066 6996 26077
rect 7030 26066 7064 26077
rect 7098 26066 7132 26077
rect 7166 26066 7200 26100
rect 7236 26077 7268 26100
rect 7308 26077 7336 26100
rect 7380 26077 7404 26100
rect 7452 26077 7472 26100
rect 7524 26077 7540 26100
rect 7596 26077 7608 26100
rect 7668 26077 7676 26100
rect 7740 26077 7744 26100
rect 7234 26066 7268 26077
rect 7302 26066 7336 26077
rect 7370 26066 7404 26077
rect 7438 26066 7472 26077
rect 7506 26066 7540 26077
rect 7574 26066 7608 26077
rect 7642 26066 7676 26077
rect 7710 26066 7744 26077
rect 7812 26100 7850 26111
rect 7884 26100 7922 26111
rect 7956 26100 7994 26111
rect 8028 26100 8066 26111
rect 8100 26100 8138 26111
rect 8172 26100 8210 26111
rect 8244 26100 8282 26111
rect 8316 26100 8354 26111
rect 8388 26100 8426 26111
rect 8460 26100 8498 26111
rect 8532 26100 8570 26111
rect 8604 26100 8642 26111
rect 8676 26100 8714 26111
rect 8748 26100 8786 26111
rect 8820 26100 8858 26111
rect 8892 26100 8930 26111
rect 8964 26100 9002 26111
rect 7778 26066 7812 26077
rect 7846 26077 7850 26100
rect 7914 26077 7922 26100
rect 7982 26077 7994 26100
rect 8050 26077 8066 26100
rect 8118 26077 8138 26100
rect 8186 26077 8210 26100
rect 8254 26077 8282 26100
rect 8322 26077 8354 26100
rect 7846 26066 7880 26077
rect 7914 26066 7948 26077
rect 7982 26066 8016 26077
rect 8050 26066 8084 26077
rect 8118 26066 8152 26077
rect 8186 26066 8220 26077
rect 8254 26066 8288 26077
rect 8322 26066 8356 26077
rect 8390 26066 8424 26100
rect 8460 26077 8492 26100
rect 8532 26077 8560 26100
rect 8604 26077 8628 26100
rect 8676 26077 8696 26100
rect 8748 26077 8764 26100
rect 8820 26077 8832 26100
rect 8892 26077 8900 26100
rect 8964 26077 8968 26100
rect 8458 26066 8492 26077
rect 8526 26066 8560 26077
rect 8594 26066 8628 26077
rect 8662 26066 8696 26077
rect 8730 26066 8764 26077
rect 8798 26066 8832 26077
rect 8866 26066 8900 26077
rect 8934 26066 8968 26077
rect 9036 26100 9074 26111
rect 9108 26100 9146 26111
rect 9180 26100 9218 26111
rect 9252 26100 9290 26111
rect 9324 26100 9362 26111
rect 9396 26100 9434 26111
rect 9468 26100 9506 26111
rect 9540 26100 9578 26111
rect 9612 26100 9650 26111
rect 9684 26100 9722 26111
rect 9756 26100 9794 26111
rect 9828 26100 9866 26111
rect 9900 26100 9938 26111
rect 9972 26100 10010 26111
rect 10044 26100 10082 26111
rect 10116 26100 10154 26111
rect 10188 26100 10226 26111
rect 9002 26066 9036 26077
rect 9070 26077 9074 26100
rect 9138 26077 9146 26100
rect 9206 26077 9218 26100
rect 9274 26077 9290 26100
rect 9342 26077 9362 26100
rect 9410 26077 9434 26100
rect 9478 26077 9506 26100
rect 9546 26077 9578 26100
rect 9070 26066 9104 26077
rect 9138 26066 9172 26077
rect 9206 26066 9240 26077
rect 9274 26066 9308 26077
rect 9342 26066 9376 26077
rect 9410 26066 9444 26077
rect 9478 26066 9512 26077
rect 9546 26066 9580 26077
rect 9614 26066 9648 26100
rect 9684 26077 9716 26100
rect 9756 26077 9784 26100
rect 9828 26077 9852 26100
rect 9900 26077 9920 26100
rect 9972 26077 9988 26100
rect 10044 26077 10056 26100
rect 10116 26077 10124 26100
rect 10188 26077 10192 26100
rect 9682 26066 9716 26077
rect 9750 26066 9784 26077
rect 9818 26066 9852 26077
rect 9886 26066 9920 26077
rect 9954 26066 9988 26077
rect 10022 26066 10056 26077
rect 10090 26066 10124 26077
rect 10158 26066 10192 26077
rect 10260 26100 10298 26111
rect 10332 26100 10370 26111
rect 10404 26100 10442 26111
rect 10476 26100 10514 26111
rect 10548 26100 10586 26111
rect 10620 26100 10658 26111
rect 10692 26100 10730 26111
rect 10764 26100 10802 26111
rect 10836 26100 10874 26111
rect 10908 26100 10946 26111
rect 10980 26100 11018 26111
rect 11052 26100 11090 26111
rect 11124 26100 11162 26111
rect 11196 26100 11234 26111
rect 11268 26100 11306 26111
rect 11340 26100 11378 26111
rect 11412 26100 11450 26111
rect 10226 26066 10260 26077
rect 10294 26077 10298 26100
rect 10362 26077 10370 26100
rect 10430 26077 10442 26100
rect 10498 26077 10514 26100
rect 10566 26077 10586 26100
rect 10634 26077 10658 26100
rect 10702 26077 10730 26100
rect 10770 26077 10802 26100
rect 10294 26066 10328 26077
rect 10362 26066 10396 26077
rect 10430 26066 10464 26077
rect 10498 26066 10532 26077
rect 10566 26066 10600 26077
rect 10634 26066 10668 26077
rect 10702 26066 10736 26077
rect 10770 26066 10804 26077
rect 10838 26066 10872 26100
rect 10908 26077 10940 26100
rect 10980 26077 11008 26100
rect 11052 26077 11076 26100
rect 11124 26077 11144 26100
rect 11196 26077 11212 26100
rect 11268 26077 11280 26100
rect 11340 26077 11348 26100
rect 11412 26077 11416 26100
rect 10906 26066 10940 26077
rect 10974 26066 11008 26077
rect 11042 26066 11076 26077
rect 11110 26066 11144 26077
rect 11178 26066 11212 26077
rect 11246 26066 11280 26077
rect 11314 26066 11348 26077
rect 11382 26066 11416 26077
rect 11484 26100 11522 26111
rect 11556 26100 11594 26111
rect 11628 26100 11666 26111
rect 11700 26100 11738 26111
rect 11772 26100 11810 26111
rect 11844 26100 11882 26111
rect 11916 26100 11954 26111
rect 11988 26100 12026 26111
rect 12060 26100 12098 26111
rect 12132 26100 12170 26111
rect 12204 26100 12242 26111
rect 12276 26100 12314 26111
rect 12348 26100 12386 26111
rect 12420 26100 12458 26111
rect 12492 26100 12530 26111
rect 12564 26100 12602 26111
rect 12636 26100 12674 26111
rect 11450 26066 11484 26077
rect 11518 26077 11522 26100
rect 11586 26077 11594 26100
rect 11654 26077 11666 26100
rect 11722 26077 11738 26100
rect 11790 26077 11810 26100
rect 11858 26077 11882 26100
rect 11926 26077 11954 26100
rect 11994 26077 12026 26100
rect 11518 26066 11552 26077
rect 11586 26066 11620 26077
rect 11654 26066 11688 26077
rect 11722 26066 11756 26077
rect 11790 26066 11824 26077
rect 11858 26066 11892 26077
rect 11926 26066 11960 26077
rect 11994 26066 12028 26077
rect 12062 26066 12096 26100
rect 12132 26077 12164 26100
rect 12204 26077 12232 26100
rect 12276 26077 12300 26100
rect 12348 26077 12368 26100
rect 12420 26077 12436 26100
rect 12492 26077 12504 26100
rect 12564 26077 12572 26100
rect 12636 26077 12640 26100
rect 12130 26066 12164 26077
rect 12198 26066 12232 26077
rect 12266 26066 12300 26077
rect 12334 26066 12368 26077
rect 12402 26066 12436 26077
rect 12470 26066 12504 26077
rect 12538 26066 12572 26077
rect 12606 26066 12640 26077
rect 12708 26100 12746 26111
rect 12780 26100 12818 26111
rect 12852 26100 12890 26111
rect 12924 26100 12962 26111
rect 12996 26100 13034 26111
rect 13068 26100 13106 26111
rect 13140 26100 13178 26111
rect 13212 26100 13250 26111
rect 13284 26100 13322 26111
rect 13356 26100 13394 26111
rect 13428 26100 13466 26111
rect 13500 26100 13538 26111
rect 13572 26100 13610 26111
rect 13644 26100 13682 26111
rect 13716 26100 13754 26111
rect 13788 26100 13826 26111
rect 13860 26100 13898 26111
rect 12674 26066 12708 26077
rect 12742 26077 12746 26100
rect 12810 26077 12818 26100
rect 12878 26077 12890 26100
rect 12946 26077 12962 26100
rect 13014 26077 13034 26100
rect 13082 26077 13106 26100
rect 13150 26077 13178 26100
rect 13218 26077 13250 26100
rect 12742 26066 12776 26077
rect 12810 26066 12844 26077
rect 12878 26066 12912 26077
rect 12946 26066 12980 26077
rect 13014 26066 13048 26077
rect 13082 26066 13116 26077
rect 13150 26066 13184 26077
rect 13218 26066 13252 26077
rect 13286 26066 13320 26100
rect 13356 26077 13388 26100
rect 13428 26077 13456 26100
rect 13500 26077 13524 26100
rect 13572 26077 13592 26100
rect 13644 26077 13660 26100
rect 13716 26077 13728 26100
rect 13788 26077 13796 26100
rect 13860 26077 13864 26100
rect 13354 26066 13388 26077
rect 13422 26066 13456 26077
rect 13490 26066 13524 26077
rect 13558 26066 13592 26077
rect 13626 26066 13660 26077
rect 13694 26066 13728 26077
rect 13762 26066 13796 26077
rect 13830 26066 13864 26077
rect 13932 26100 13970 26111
rect 14004 26100 14042 26111
rect 14076 26100 14114 26111
rect 14148 26100 14186 26111
rect 14220 26100 14258 26111
rect 14292 26100 14330 26111
rect 14364 26100 14402 26111
rect 14436 26100 14474 26111
rect 14508 26100 14546 26111
rect 14580 26100 14618 26111
rect 14652 26100 14690 26111
rect 14724 26100 14962 26111
rect 13898 26066 13932 26077
rect 13966 26077 13970 26100
rect 14034 26077 14042 26100
rect 14102 26077 14114 26100
rect 14170 26077 14186 26100
rect 14238 26077 14258 26100
rect 14306 26077 14330 26100
rect 14374 26077 14402 26100
rect 14442 26077 14474 26100
rect 13966 26066 14000 26077
rect 14034 26066 14068 26077
rect 14102 26066 14136 26077
rect 14170 26066 14204 26077
rect 14238 26066 14272 26077
rect 14306 26066 14340 26077
rect 14374 26066 14408 26077
rect 14442 26066 14476 26077
rect 14510 26066 14544 26100
rect 14580 26077 14612 26100
rect 14652 26077 14680 26100
rect 14724 26077 14748 26100
rect 14578 26066 14612 26077
rect 14646 26066 14680 26077
rect 14714 26066 14748 26077
rect 14782 26066 14816 26100
rect 14850 26066 14884 26100
rect 14918 26066 14962 26100
rect 49 26037 14962 26066
rect 49 26028 243 26037
rect 277 26028 316 26037
rect 350 26028 389 26037
rect 423 26028 462 26037
rect 496 26028 535 26037
rect 569 26028 608 26037
rect 642 26028 681 26037
rect 715 26028 754 26037
rect 788 26028 827 26037
rect 861 26028 900 26037
rect 934 26028 973 26037
rect 1007 26028 1046 26037
rect 1080 26028 1119 26037
rect 1153 26028 1192 26037
rect 1226 26028 1265 26037
rect 1299 26028 1338 26037
rect 1372 26028 1411 26037
rect 1445 26028 1484 26037
rect 49 25994 69 26028
rect 103 25994 138 26028
rect 172 25994 207 26028
rect 241 26003 243 26028
rect 310 26003 316 26028
rect 379 26003 389 26028
rect 448 26003 462 26028
rect 517 26003 535 26028
rect 586 26003 608 26028
rect 655 26003 681 26028
rect 724 26003 754 26028
rect 793 26003 827 26028
rect 241 25994 276 26003
rect 310 25994 345 26003
rect 379 25994 414 26003
rect 448 25994 483 26003
rect 517 25994 552 26003
rect 586 25994 621 26003
rect 655 25994 690 26003
rect 724 25994 759 26003
rect 793 25994 828 26003
rect 862 25994 897 26028
rect 934 26003 966 26028
rect 1007 26003 1035 26028
rect 1080 26003 1104 26028
rect 1153 26003 1173 26028
rect 1226 26003 1242 26028
rect 1299 26003 1311 26028
rect 1372 26003 1380 26028
rect 1445 26003 1449 26028
rect 931 25994 966 26003
rect 1000 25994 1035 26003
rect 1069 25994 1104 26003
rect 1138 25994 1173 26003
rect 1207 25994 1242 26003
rect 1276 25994 1311 26003
rect 1345 25994 1380 26003
rect 1414 25994 1449 26003
rect 1483 26003 1484 26028
rect 1518 26028 1557 26037
rect 1591 26028 1630 26037
rect 1664 26028 1703 26037
rect 1737 26028 1776 26037
rect 1810 26028 1849 26037
rect 1883 26028 1922 26037
rect 1956 26028 1995 26037
rect 2029 26028 2068 26037
rect 2102 26028 2141 26037
rect 2175 26028 2214 26037
rect 2248 26028 2287 26037
rect 2321 26028 2360 26037
rect 2394 26028 2433 26037
rect 2467 26028 2506 26037
rect 2540 26028 2579 26037
rect 2613 26028 2652 26037
rect 2686 26028 2725 26037
rect 1483 25994 1518 26003
rect 1552 26003 1557 26028
rect 1621 26003 1630 26028
rect 1690 26003 1703 26028
rect 1759 26003 1776 26028
rect 1828 26003 1849 26028
rect 1897 26003 1922 26028
rect 1966 26003 1995 26028
rect 2035 26003 2068 26028
rect 1552 25994 1587 26003
rect 1621 25994 1656 26003
rect 1690 25994 1725 26003
rect 1759 25994 1794 26003
rect 1828 25994 1863 26003
rect 1897 25994 1932 26003
rect 1966 25994 2001 26003
rect 2035 25994 2070 26003
rect 2104 25994 2139 26028
rect 2175 26003 2208 26028
rect 2248 26003 2277 26028
rect 2321 26003 2346 26028
rect 2394 26003 2415 26028
rect 2467 26003 2484 26028
rect 2540 26003 2553 26028
rect 2613 26003 2622 26028
rect 2686 26003 2691 26028
rect 2173 25994 2208 26003
rect 2242 25994 2277 26003
rect 2311 25994 2346 26003
rect 2380 25994 2415 26003
rect 2449 25994 2484 26003
rect 2518 25994 2553 26003
rect 2587 25994 2622 26003
rect 2656 25994 2691 26003
rect 2759 26028 2798 26037
rect 2832 26028 2871 26037
rect 2905 26028 2944 26037
rect 2978 26028 3017 26037
rect 3051 26028 3090 26037
rect 3124 26028 3163 26037
rect 3197 26028 3236 26037
rect 3270 26028 3309 26037
rect 3343 26028 3382 26037
rect 3416 26028 3455 26037
rect 3489 26028 3528 26037
rect 3562 26028 3601 26037
rect 3635 26028 3674 26037
rect 3708 26028 3746 26037
rect 3780 26028 3818 26037
rect 3852 26028 3890 26037
rect 3924 26028 3962 26037
rect 3996 26028 4034 26037
rect 4068 26028 4106 26037
rect 2759 26003 2760 26028
rect 2725 25994 2760 26003
rect 2794 26003 2798 26028
rect 2863 26003 2871 26028
rect 2932 26003 2944 26028
rect 3001 26003 3017 26028
rect 3070 26003 3090 26028
rect 3139 26003 3163 26028
rect 3208 26003 3236 26028
rect 3277 26003 3309 26028
rect 2794 25994 2829 26003
rect 2863 25994 2898 26003
rect 2932 25994 2967 26003
rect 3001 25994 3036 26003
rect 3070 25994 3105 26003
rect 3139 25994 3174 26003
rect 3208 25994 3243 26003
rect 3277 25994 3312 26003
rect 3346 25994 3381 26028
rect 3416 26003 3450 26028
rect 3489 26003 3519 26028
rect 3562 26003 3588 26028
rect 3635 26003 3657 26028
rect 3708 26003 3726 26028
rect 3780 26003 3795 26028
rect 3852 26003 3864 26028
rect 3924 26003 3933 26028
rect 3996 26003 4002 26028
rect 4068 26003 4071 26028
rect 3415 25994 3450 26003
rect 3484 25994 3519 26003
rect 3553 25994 3588 26003
rect 3622 25994 3657 26003
rect 3691 25994 3726 26003
rect 3760 25994 3795 26003
rect 3829 25994 3864 26003
rect 3898 25994 3933 26003
rect 3967 25994 4002 26003
rect 4036 25994 4071 26003
rect 4105 26003 4106 26028
rect 4140 26028 4178 26037
rect 4212 26028 4250 26037
rect 4284 26028 4322 26037
rect 4356 26028 4394 26037
rect 4428 26028 4466 26037
rect 4500 26028 4538 26037
rect 4572 26028 4610 26037
rect 4644 26028 4682 26037
rect 4716 26028 4754 26037
rect 4788 26028 4826 26037
rect 4860 26028 4898 26037
rect 4932 26028 4970 26037
rect 5004 26028 5042 26037
rect 5076 26028 5114 26037
rect 5148 26028 5186 26037
rect 5220 26028 5258 26037
rect 5292 26028 5330 26037
rect 4105 25994 4140 26003
rect 4174 26003 4178 26028
rect 4242 26003 4250 26028
rect 4310 26003 4322 26028
rect 4378 26003 4394 26028
rect 4446 26003 4466 26028
rect 4514 26003 4538 26028
rect 4582 26003 4610 26028
rect 4650 26003 4682 26028
rect 4174 25994 4208 26003
rect 4242 25994 4276 26003
rect 4310 25994 4344 26003
rect 4378 25994 4412 26003
rect 4446 25994 4480 26003
rect 4514 25994 4548 26003
rect 4582 25994 4616 26003
rect 4650 25994 4684 26003
rect 4718 25994 4752 26028
rect 4788 26003 4820 26028
rect 4860 26003 4888 26028
rect 4932 26003 4956 26028
rect 5004 26003 5024 26028
rect 5076 26003 5092 26028
rect 5148 26003 5160 26028
rect 5220 26003 5228 26028
rect 5292 26003 5296 26028
rect 4786 25994 4820 26003
rect 4854 25994 4888 26003
rect 4922 25994 4956 26003
rect 4990 25994 5024 26003
rect 5058 25994 5092 26003
rect 5126 25994 5160 26003
rect 5194 25994 5228 26003
rect 5262 25994 5296 26003
rect 5364 26028 5402 26037
rect 5436 26028 5474 26037
rect 5508 26028 5546 26037
rect 5580 26028 5618 26037
rect 5652 26028 5690 26037
rect 5724 26028 5762 26037
rect 5796 26028 5834 26037
rect 5868 26028 5906 26037
rect 5940 26028 5978 26037
rect 6012 26028 6050 26037
rect 6084 26028 6122 26037
rect 6156 26028 6194 26037
rect 6228 26028 6266 26037
rect 6300 26028 6338 26037
rect 6372 26028 6410 26037
rect 6444 26028 6482 26037
rect 6516 26028 6554 26037
rect 5330 25994 5364 26003
rect 5398 26003 5402 26028
rect 5466 26003 5474 26028
rect 5534 26003 5546 26028
rect 5602 26003 5618 26028
rect 5670 26003 5690 26028
rect 5738 26003 5762 26028
rect 5806 26003 5834 26028
rect 5874 26003 5906 26028
rect 5398 25994 5432 26003
rect 5466 25994 5500 26003
rect 5534 25994 5568 26003
rect 5602 25994 5636 26003
rect 5670 25994 5704 26003
rect 5738 25994 5772 26003
rect 5806 25994 5840 26003
rect 5874 25994 5908 26003
rect 5942 25994 5976 26028
rect 6012 26003 6044 26028
rect 6084 26003 6112 26028
rect 6156 26003 6180 26028
rect 6228 26003 6248 26028
rect 6300 26003 6316 26028
rect 6372 26003 6384 26028
rect 6444 26003 6452 26028
rect 6516 26003 6520 26028
rect 6010 25994 6044 26003
rect 6078 25994 6112 26003
rect 6146 25994 6180 26003
rect 6214 25994 6248 26003
rect 6282 25994 6316 26003
rect 6350 25994 6384 26003
rect 6418 25994 6452 26003
rect 6486 25994 6520 26003
rect 6588 26028 6626 26037
rect 6660 26028 6698 26037
rect 6732 26028 6770 26037
rect 6804 26028 6842 26037
rect 6876 26028 6914 26037
rect 6948 26028 6986 26037
rect 7020 26028 7058 26037
rect 7092 26028 7130 26037
rect 7164 26028 7202 26037
rect 7236 26028 7274 26037
rect 7308 26028 7346 26037
rect 7380 26028 7418 26037
rect 7452 26028 7490 26037
rect 7524 26028 7562 26037
rect 7596 26028 7634 26037
rect 7668 26028 7706 26037
rect 7740 26028 7778 26037
rect 6554 25994 6588 26003
rect 6622 26003 6626 26028
rect 6690 26003 6698 26028
rect 6758 26003 6770 26028
rect 6826 26003 6842 26028
rect 6894 26003 6914 26028
rect 6962 26003 6986 26028
rect 7030 26003 7058 26028
rect 7098 26003 7130 26028
rect 6622 25994 6656 26003
rect 6690 25994 6724 26003
rect 6758 25994 6792 26003
rect 6826 25994 6860 26003
rect 6894 25994 6928 26003
rect 6962 25994 6996 26003
rect 7030 25994 7064 26003
rect 7098 25994 7132 26003
rect 7166 25994 7200 26028
rect 7236 26003 7268 26028
rect 7308 26003 7336 26028
rect 7380 26003 7404 26028
rect 7452 26003 7472 26028
rect 7524 26003 7540 26028
rect 7596 26003 7608 26028
rect 7668 26003 7676 26028
rect 7740 26003 7744 26028
rect 7234 25994 7268 26003
rect 7302 25994 7336 26003
rect 7370 25994 7404 26003
rect 7438 25994 7472 26003
rect 7506 25994 7540 26003
rect 7574 25994 7608 26003
rect 7642 25994 7676 26003
rect 7710 25994 7744 26003
rect 7812 26028 7850 26037
rect 7884 26028 7922 26037
rect 7956 26028 7994 26037
rect 8028 26028 8066 26037
rect 8100 26028 8138 26037
rect 8172 26028 8210 26037
rect 8244 26028 8282 26037
rect 8316 26028 8354 26037
rect 8388 26028 8426 26037
rect 8460 26028 8498 26037
rect 8532 26028 8570 26037
rect 8604 26028 8642 26037
rect 8676 26028 8714 26037
rect 8748 26028 8786 26037
rect 8820 26028 8858 26037
rect 8892 26028 8930 26037
rect 8964 26028 9002 26037
rect 7778 25994 7812 26003
rect 7846 26003 7850 26028
rect 7914 26003 7922 26028
rect 7982 26003 7994 26028
rect 8050 26003 8066 26028
rect 8118 26003 8138 26028
rect 8186 26003 8210 26028
rect 8254 26003 8282 26028
rect 8322 26003 8354 26028
rect 7846 25994 7880 26003
rect 7914 25994 7948 26003
rect 7982 25994 8016 26003
rect 8050 25994 8084 26003
rect 8118 25994 8152 26003
rect 8186 25994 8220 26003
rect 8254 25994 8288 26003
rect 8322 25994 8356 26003
rect 8390 25994 8424 26028
rect 8460 26003 8492 26028
rect 8532 26003 8560 26028
rect 8604 26003 8628 26028
rect 8676 26003 8696 26028
rect 8748 26003 8764 26028
rect 8820 26003 8832 26028
rect 8892 26003 8900 26028
rect 8964 26003 8968 26028
rect 8458 25994 8492 26003
rect 8526 25994 8560 26003
rect 8594 25994 8628 26003
rect 8662 25994 8696 26003
rect 8730 25994 8764 26003
rect 8798 25994 8832 26003
rect 8866 25994 8900 26003
rect 8934 25994 8968 26003
rect 9036 26028 9074 26037
rect 9108 26028 9146 26037
rect 9180 26028 9218 26037
rect 9252 26028 9290 26037
rect 9324 26028 9362 26037
rect 9396 26028 9434 26037
rect 9468 26028 9506 26037
rect 9540 26028 9578 26037
rect 9612 26028 9650 26037
rect 9684 26028 9722 26037
rect 9756 26028 9794 26037
rect 9828 26028 9866 26037
rect 9900 26028 9938 26037
rect 9972 26028 10010 26037
rect 10044 26028 10082 26037
rect 10116 26028 10154 26037
rect 10188 26028 10226 26037
rect 9002 25994 9036 26003
rect 9070 26003 9074 26028
rect 9138 26003 9146 26028
rect 9206 26003 9218 26028
rect 9274 26003 9290 26028
rect 9342 26003 9362 26028
rect 9410 26003 9434 26028
rect 9478 26003 9506 26028
rect 9546 26003 9578 26028
rect 9070 25994 9104 26003
rect 9138 25994 9172 26003
rect 9206 25994 9240 26003
rect 9274 25994 9308 26003
rect 9342 25994 9376 26003
rect 9410 25994 9444 26003
rect 9478 25994 9512 26003
rect 9546 25994 9580 26003
rect 9614 25994 9648 26028
rect 9684 26003 9716 26028
rect 9756 26003 9784 26028
rect 9828 26003 9852 26028
rect 9900 26003 9920 26028
rect 9972 26003 9988 26028
rect 10044 26003 10056 26028
rect 10116 26003 10124 26028
rect 10188 26003 10192 26028
rect 9682 25994 9716 26003
rect 9750 25994 9784 26003
rect 9818 25994 9852 26003
rect 9886 25994 9920 26003
rect 9954 25994 9988 26003
rect 10022 25994 10056 26003
rect 10090 25994 10124 26003
rect 10158 25994 10192 26003
rect 10260 26028 10298 26037
rect 10332 26028 10370 26037
rect 10404 26028 10442 26037
rect 10476 26028 10514 26037
rect 10548 26028 10586 26037
rect 10620 26028 10658 26037
rect 10692 26028 10730 26037
rect 10764 26028 10802 26037
rect 10836 26028 10874 26037
rect 10908 26028 10946 26037
rect 10980 26028 11018 26037
rect 11052 26028 11090 26037
rect 11124 26028 11162 26037
rect 11196 26028 11234 26037
rect 11268 26028 11306 26037
rect 11340 26028 11378 26037
rect 11412 26028 11450 26037
rect 10226 25994 10260 26003
rect 10294 26003 10298 26028
rect 10362 26003 10370 26028
rect 10430 26003 10442 26028
rect 10498 26003 10514 26028
rect 10566 26003 10586 26028
rect 10634 26003 10658 26028
rect 10702 26003 10730 26028
rect 10770 26003 10802 26028
rect 10294 25994 10328 26003
rect 10362 25994 10396 26003
rect 10430 25994 10464 26003
rect 10498 25994 10532 26003
rect 10566 25994 10600 26003
rect 10634 25994 10668 26003
rect 10702 25994 10736 26003
rect 10770 25994 10804 26003
rect 10838 25994 10872 26028
rect 10908 26003 10940 26028
rect 10980 26003 11008 26028
rect 11052 26003 11076 26028
rect 11124 26003 11144 26028
rect 11196 26003 11212 26028
rect 11268 26003 11280 26028
rect 11340 26003 11348 26028
rect 11412 26003 11416 26028
rect 10906 25994 10940 26003
rect 10974 25994 11008 26003
rect 11042 25994 11076 26003
rect 11110 25994 11144 26003
rect 11178 25994 11212 26003
rect 11246 25994 11280 26003
rect 11314 25994 11348 26003
rect 11382 25994 11416 26003
rect 11484 26028 11522 26037
rect 11556 26028 11594 26037
rect 11628 26028 11666 26037
rect 11700 26028 11738 26037
rect 11772 26028 11810 26037
rect 11844 26028 11882 26037
rect 11916 26028 11954 26037
rect 11988 26028 12026 26037
rect 12060 26028 12098 26037
rect 12132 26028 12170 26037
rect 12204 26028 12242 26037
rect 12276 26028 12314 26037
rect 12348 26028 12386 26037
rect 12420 26028 12458 26037
rect 12492 26028 12530 26037
rect 12564 26028 12602 26037
rect 12636 26028 12674 26037
rect 11450 25994 11484 26003
rect 11518 26003 11522 26028
rect 11586 26003 11594 26028
rect 11654 26003 11666 26028
rect 11722 26003 11738 26028
rect 11790 26003 11810 26028
rect 11858 26003 11882 26028
rect 11926 26003 11954 26028
rect 11994 26003 12026 26028
rect 11518 25994 11552 26003
rect 11586 25994 11620 26003
rect 11654 25994 11688 26003
rect 11722 25994 11756 26003
rect 11790 25994 11824 26003
rect 11858 25994 11892 26003
rect 11926 25994 11960 26003
rect 11994 25994 12028 26003
rect 12062 25994 12096 26028
rect 12132 26003 12164 26028
rect 12204 26003 12232 26028
rect 12276 26003 12300 26028
rect 12348 26003 12368 26028
rect 12420 26003 12436 26028
rect 12492 26003 12504 26028
rect 12564 26003 12572 26028
rect 12636 26003 12640 26028
rect 12130 25994 12164 26003
rect 12198 25994 12232 26003
rect 12266 25994 12300 26003
rect 12334 25994 12368 26003
rect 12402 25994 12436 26003
rect 12470 25994 12504 26003
rect 12538 25994 12572 26003
rect 12606 25994 12640 26003
rect 12708 26028 12746 26037
rect 12780 26028 12818 26037
rect 12852 26028 12890 26037
rect 12924 26028 12962 26037
rect 12996 26028 13034 26037
rect 13068 26028 13106 26037
rect 13140 26028 13178 26037
rect 13212 26028 13250 26037
rect 13284 26028 13322 26037
rect 13356 26028 13394 26037
rect 13428 26028 13466 26037
rect 13500 26028 13538 26037
rect 13572 26028 13610 26037
rect 13644 26028 13682 26037
rect 13716 26028 13754 26037
rect 13788 26028 13826 26037
rect 13860 26028 13898 26037
rect 12674 25994 12708 26003
rect 12742 26003 12746 26028
rect 12810 26003 12818 26028
rect 12878 26003 12890 26028
rect 12946 26003 12962 26028
rect 13014 26003 13034 26028
rect 13082 26003 13106 26028
rect 13150 26003 13178 26028
rect 13218 26003 13250 26028
rect 12742 25994 12776 26003
rect 12810 25994 12844 26003
rect 12878 25994 12912 26003
rect 12946 25994 12980 26003
rect 13014 25994 13048 26003
rect 13082 25994 13116 26003
rect 13150 25994 13184 26003
rect 13218 25994 13252 26003
rect 13286 25994 13320 26028
rect 13356 26003 13388 26028
rect 13428 26003 13456 26028
rect 13500 26003 13524 26028
rect 13572 26003 13592 26028
rect 13644 26003 13660 26028
rect 13716 26003 13728 26028
rect 13788 26003 13796 26028
rect 13860 26003 13864 26028
rect 13354 25994 13388 26003
rect 13422 25994 13456 26003
rect 13490 25994 13524 26003
rect 13558 25994 13592 26003
rect 13626 25994 13660 26003
rect 13694 25994 13728 26003
rect 13762 25994 13796 26003
rect 13830 25994 13864 26003
rect 13932 26028 13970 26037
rect 14004 26028 14042 26037
rect 14076 26028 14114 26037
rect 14148 26028 14186 26037
rect 14220 26028 14258 26037
rect 14292 26028 14330 26037
rect 14364 26028 14402 26037
rect 14436 26028 14474 26037
rect 14508 26028 14546 26037
rect 14580 26028 14618 26037
rect 14652 26028 14690 26037
rect 14724 26028 14962 26037
rect 13898 25994 13932 26003
rect 13966 26003 13970 26028
rect 14034 26003 14042 26028
rect 14102 26003 14114 26028
rect 14170 26003 14186 26028
rect 14238 26003 14258 26028
rect 14306 26003 14330 26028
rect 14374 26003 14402 26028
rect 14442 26003 14474 26028
rect 13966 25994 14000 26003
rect 14034 25994 14068 26003
rect 14102 25994 14136 26003
rect 14170 25994 14204 26003
rect 14238 25994 14272 26003
rect 14306 25994 14340 26003
rect 14374 25994 14408 26003
rect 14442 25994 14476 26003
rect 14510 25994 14544 26028
rect 14580 26003 14612 26028
rect 14652 26003 14680 26028
rect 14724 26003 14748 26028
rect 14578 25994 14612 26003
rect 14646 25994 14680 26003
rect 14714 25994 14748 26003
rect 14782 25994 14816 26028
rect 14850 25994 14884 26028
rect 14918 25994 14962 26028
rect 49 25963 14962 25994
rect 49 25956 243 25963
rect 277 25956 316 25963
rect 350 25956 389 25963
rect 423 25956 462 25963
rect 496 25956 535 25963
rect 569 25956 608 25963
rect 642 25956 681 25963
rect 715 25956 754 25963
rect 788 25956 827 25963
rect 861 25956 900 25963
rect 934 25956 973 25963
rect 1007 25956 1046 25963
rect 1080 25956 1119 25963
rect 1153 25956 1192 25963
rect 1226 25956 1265 25963
rect 1299 25956 1338 25963
rect 1372 25956 1411 25963
rect 1445 25956 1484 25963
rect 49 25922 69 25956
rect 103 25922 138 25956
rect 172 25922 207 25956
rect 241 25929 243 25956
rect 310 25929 316 25956
rect 379 25929 389 25956
rect 448 25929 462 25956
rect 517 25929 535 25956
rect 586 25929 608 25956
rect 655 25929 681 25956
rect 724 25929 754 25956
rect 793 25929 827 25956
rect 241 25922 276 25929
rect 310 25922 345 25929
rect 379 25922 414 25929
rect 448 25922 483 25929
rect 517 25922 552 25929
rect 586 25922 621 25929
rect 655 25922 690 25929
rect 724 25922 759 25929
rect 793 25922 828 25929
rect 862 25922 897 25956
rect 934 25929 966 25956
rect 1007 25929 1035 25956
rect 1080 25929 1104 25956
rect 1153 25929 1173 25956
rect 1226 25929 1242 25956
rect 1299 25929 1311 25956
rect 1372 25929 1380 25956
rect 1445 25929 1449 25956
rect 931 25922 966 25929
rect 1000 25922 1035 25929
rect 1069 25922 1104 25929
rect 1138 25922 1173 25929
rect 1207 25922 1242 25929
rect 1276 25922 1311 25929
rect 1345 25922 1380 25929
rect 1414 25922 1449 25929
rect 1483 25929 1484 25956
rect 1518 25956 1557 25963
rect 1591 25956 1630 25963
rect 1664 25956 1703 25963
rect 1737 25956 1776 25963
rect 1810 25956 1849 25963
rect 1883 25956 1922 25963
rect 1956 25956 1995 25963
rect 2029 25956 2068 25963
rect 2102 25956 2141 25963
rect 2175 25956 2214 25963
rect 2248 25956 2287 25963
rect 2321 25956 2360 25963
rect 2394 25956 2433 25963
rect 2467 25956 2506 25963
rect 2540 25956 2579 25963
rect 2613 25956 2652 25963
rect 2686 25956 2725 25963
rect 1483 25922 1518 25929
rect 1552 25929 1557 25956
rect 1621 25929 1630 25956
rect 1690 25929 1703 25956
rect 1759 25929 1776 25956
rect 1828 25929 1849 25956
rect 1897 25929 1922 25956
rect 1966 25929 1995 25956
rect 2035 25929 2068 25956
rect 1552 25922 1587 25929
rect 1621 25922 1656 25929
rect 1690 25922 1725 25929
rect 1759 25922 1794 25929
rect 1828 25922 1863 25929
rect 1897 25922 1932 25929
rect 1966 25922 2001 25929
rect 2035 25922 2070 25929
rect 2104 25922 2139 25956
rect 2175 25929 2208 25956
rect 2248 25929 2277 25956
rect 2321 25929 2346 25956
rect 2394 25929 2415 25956
rect 2467 25929 2484 25956
rect 2540 25929 2553 25956
rect 2613 25929 2622 25956
rect 2686 25929 2691 25956
rect 2173 25922 2208 25929
rect 2242 25922 2277 25929
rect 2311 25922 2346 25929
rect 2380 25922 2415 25929
rect 2449 25922 2484 25929
rect 2518 25922 2553 25929
rect 2587 25922 2622 25929
rect 2656 25922 2691 25929
rect 2759 25956 2798 25963
rect 2832 25956 2871 25963
rect 2905 25956 2944 25963
rect 2978 25956 3017 25963
rect 3051 25956 3090 25963
rect 3124 25956 3163 25963
rect 3197 25956 3236 25963
rect 3270 25956 3309 25963
rect 3343 25956 3382 25963
rect 3416 25956 3455 25963
rect 3489 25956 3528 25963
rect 3562 25956 3601 25963
rect 3635 25956 3674 25963
rect 3708 25956 3746 25963
rect 3780 25956 3818 25963
rect 3852 25956 3890 25963
rect 3924 25956 3962 25963
rect 3996 25956 4034 25963
rect 4068 25956 4106 25963
rect 2759 25929 2760 25956
rect 2725 25922 2760 25929
rect 2794 25929 2798 25956
rect 2863 25929 2871 25956
rect 2932 25929 2944 25956
rect 3001 25929 3017 25956
rect 3070 25929 3090 25956
rect 3139 25929 3163 25956
rect 3208 25929 3236 25956
rect 3277 25929 3309 25956
rect 2794 25922 2829 25929
rect 2863 25922 2898 25929
rect 2932 25922 2967 25929
rect 3001 25922 3036 25929
rect 3070 25922 3105 25929
rect 3139 25922 3174 25929
rect 3208 25922 3243 25929
rect 3277 25922 3312 25929
rect 3346 25922 3381 25956
rect 3416 25929 3450 25956
rect 3489 25929 3519 25956
rect 3562 25929 3588 25956
rect 3635 25929 3657 25956
rect 3708 25929 3726 25956
rect 3780 25929 3795 25956
rect 3852 25929 3864 25956
rect 3924 25929 3933 25956
rect 3996 25929 4002 25956
rect 4068 25929 4071 25956
rect 3415 25922 3450 25929
rect 3484 25922 3519 25929
rect 3553 25922 3588 25929
rect 3622 25922 3657 25929
rect 3691 25922 3726 25929
rect 3760 25922 3795 25929
rect 3829 25922 3864 25929
rect 3898 25922 3933 25929
rect 3967 25922 4002 25929
rect 4036 25922 4071 25929
rect 4105 25929 4106 25956
rect 4140 25956 4178 25963
rect 4212 25956 4250 25963
rect 4284 25956 4322 25963
rect 4356 25956 4394 25963
rect 4428 25956 4466 25963
rect 4500 25956 4538 25963
rect 4572 25956 4610 25963
rect 4644 25956 4682 25963
rect 4716 25956 4754 25963
rect 4788 25956 4826 25963
rect 4860 25956 4898 25963
rect 4932 25956 4970 25963
rect 5004 25956 5042 25963
rect 5076 25956 5114 25963
rect 5148 25956 5186 25963
rect 5220 25956 5258 25963
rect 5292 25956 5330 25963
rect 4105 25922 4140 25929
rect 4174 25929 4178 25956
rect 4242 25929 4250 25956
rect 4310 25929 4322 25956
rect 4378 25929 4394 25956
rect 4446 25929 4466 25956
rect 4514 25929 4538 25956
rect 4582 25929 4610 25956
rect 4650 25929 4682 25956
rect 4174 25922 4208 25929
rect 4242 25922 4276 25929
rect 4310 25922 4344 25929
rect 4378 25922 4412 25929
rect 4446 25922 4480 25929
rect 4514 25922 4548 25929
rect 4582 25922 4616 25929
rect 4650 25922 4684 25929
rect 4718 25922 4752 25956
rect 4788 25929 4820 25956
rect 4860 25929 4888 25956
rect 4932 25929 4956 25956
rect 5004 25929 5024 25956
rect 5076 25929 5092 25956
rect 5148 25929 5160 25956
rect 5220 25929 5228 25956
rect 5292 25929 5296 25956
rect 4786 25922 4820 25929
rect 4854 25922 4888 25929
rect 4922 25922 4956 25929
rect 4990 25922 5024 25929
rect 5058 25922 5092 25929
rect 5126 25922 5160 25929
rect 5194 25922 5228 25929
rect 5262 25922 5296 25929
rect 5364 25956 5402 25963
rect 5436 25956 5474 25963
rect 5508 25956 5546 25963
rect 5580 25956 5618 25963
rect 5652 25956 5690 25963
rect 5724 25956 5762 25963
rect 5796 25956 5834 25963
rect 5868 25956 5906 25963
rect 5940 25956 5978 25963
rect 6012 25956 6050 25963
rect 6084 25956 6122 25963
rect 6156 25956 6194 25963
rect 6228 25956 6266 25963
rect 6300 25956 6338 25963
rect 6372 25956 6410 25963
rect 6444 25956 6482 25963
rect 6516 25956 6554 25963
rect 5330 25922 5364 25929
rect 5398 25929 5402 25956
rect 5466 25929 5474 25956
rect 5534 25929 5546 25956
rect 5602 25929 5618 25956
rect 5670 25929 5690 25956
rect 5738 25929 5762 25956
rect 5806 25929 5834 25956
rect 5874 25929 5906 25956
rect 5398 25922 5432 25929
rect 5466 25922 5500 25929
rect 5534 25922 5568 25929
rect 5602 25922 5636 25929
rect 5670 25922 5704 25929
rect 5738 25922 5772 25929
rect 5806 25922 5840 25929
rect 5874 25922 5908 25929
rect 5942 25922 5976 25956
rect 6012 25929 6044 25956
rect 6084 25929 6112 25956
rect 6156 25929 6180 25956
rect 6228 25929 6248 25956
rect 6300 25929 6316 25956
rect 6372 25929 6384 25956
rect 6444 25929 6452 25956
rect 6516 25929 6520 25956
rect 6010 25922 6044 25929
rect 6078 25922 6112 25929
rect 6146 25922 6180 25929
rect 6214 25922 6248 25929
rect 6282 25922 6316 25929
rect 6350 25922 6384 25929
rect 6418 25922 6452 25929
rect 6486 25922 6520 25929
rect 6588 25956 6626 25963
rect 6660 25956 6698 25963
rect 6732 25956 6770 25963
rect 6804 25956 6842 25963
rect 6876 25956 6914 25963
rect 6948 25956 6986 25963
rect 7020 25956 7058 25963
rect 7092 25956 7130 25963
rect 7164 25956 7202 25963
rect 7236 25956 7274 25963
rect 7308 25956 7346 25963
rect 7380 25956 7418 25963
rect 7452 25956 7490 25963
rect 7524 25956 7562 25963
rect 7596 25956 7634 25963
rect 7668 25956 7706 25963
rect 7740 25956 7778 25963
rect 6554 25922 6588 25929
rect 6622 25929 6626 25956
rect 6690 25929 6698 25956
rect 6758 25929 6770 25956
rect 6826 25929 6842 25956
rect 6894 25929 6914 25956
rect 6962 25929 6986 25956
rect 7030 25929 7058 25956
rect 7098 25929 7130 25956
rect 6622 25922 6656 25929
rect 6690 25922 6724 25929
rect 6758 25922 6792 25929
rect 6826 25922 6860 25929
rect 6894 25922 6928 25929
rect 6962 25922 6996 25929
rect 7030 25922 7064 25929
rect 7098 25922 7132 25929
rect 7166 25922 7200 25956
rect 7236 25929 7268 25956
rect 7308 25929 7336 25956
rect 7380 25929 7404 25956
rect 7452 25929 7472 25956
rect 7524 25929 7540 25956
rect 7596 25929 7608 25956
rect 7668 25929 7676 25956
rect 7740 25929 7744 25956
rect 7234 25922 7268 25929
rect 7302 25922 7336 25929
rect 7370 25922 7404 25929
rect 7438 25922 7472 25929
rect 7506 25922 7540 25929
rect 7574 25922 7608 25929
rect 7642 25922 7676 25929
rect 7710 25922 7744 25929
rect 7812 25956 7850 25963
rect 7884 25956 7922 25963
rect 7956 25956 7994 25963
rect 8028 25956 8066 25963
rect 8100 25956 8138 25963
rect 8172 25956 8210 25963
rect 8244 25956 8282 25963
rect 8316 25956 8354 25963
rect 8388 25956 8426 25963
rect 8460 25956 8498 25963
rect 8532 25956 8570 25963
rect 8604 25956 8642 25963
rect 8676 25956 8714 25963
rect 8748 25956 8786 25963
rect 8820 25956 8858 25963
rect 8892 25956 8930 25963
rect 8964 25956 9002 25963
rect 7778 25922 7812 25929
rect 7846 25929 7850 25956
rect 7914 25929 7922 25956
rect 7982 25929 7994 25956
rect 8050 25929 8066 25956
rect 8118 25929 8138 25956
rect 8186 25929 8210 25956
rect 8254 25929 8282 25956
rect 8322 25929 8354 25956
rect 7846 25922 7880 25929
rect 7914 25922 7948 25929
rect 7982 25922 8016 25929
rect 8050 25922 8084 25929
rect 8118 25922 8152 25929
rect 8186 25922 8220 25929
rect 8254 25922 8288 25929
rect 8322 25922 8356 25929
rect 8390 25922 8424 25956
rect 8460 25929 8492 25956
rect 8532 25929 8560 25956
rect 8604 25929 8628 25956
rect 8676 25929 8696 25956
rect 8748 25929 8764 25956
rect 8820 25929 8832 25956
rect 8892 25929 8900 25956
rect 8964 25929 8968 25956
rect 8458 25922 8492 25929
rect 8526 25922 8560 25929
rect 8594 25922 8628 25929
rect 8662 25922 8696 25929
rect 8730 25922 8764 25929
rect 8798 25922 8832 25929
rect 8866 25922 8900 25929
rect 8934 25922 8968 25929
rect 9036 25956 9074 25963
rect 9108 25956 9146 25963
rect 9180 25956 9218 25963
rect 9252 25956 9290 25963
rect 9324 25956 9362 25963
rect 9396 25956 9434 25963
rect 9468 25956 9506 25963
rect 9540 25956 9578 25963
rect 9612 25956 9650 25963
rect 9684 25956 9722 25963
rect 9756 25956 9794 25963
rect 9828 25956 9866 25963
rect 9900 25956 9938 25963
rect 9972 25956 10010 25963
rect 10044 25956 10082 25963
rect 10116 25956 10154 25963
rect 10188 25956 10226 25963
rect 9002 25922 9036 25929
rect 9070 25929 9074 25956
rect 9138 25929 9146 25956
rect 9206 25929 9218 25956
rect 9274 25929 9290 25956
rect 9342 25929 9362 25956
rect 9410 25929 9434 25956
rect 9478 25929 9506 25956
rect 9546 25929 9578 25956
rect 9070 25922 9104 25929
rect 9138 25922 9172 25929
rect 9206 25922 9240 25929
rect 9274 25922 9308 25929
rect 9342 25922 9376 25929
rect 9410 25922 9444 25929
rect 9478 25922 9512 25929
rect 9546 25922 9580 25929
rect 9614 25922 9648 25956
rect 9684 25929 9716 25956
rect 9756 25929 9784 25956
rect 9828 25929 9852 25956
rect 9900 25929 9920 25956
rect 9972 25929 9988 25956
rect 10044 25929 10056 25956
rect 10116 25929 10124 25956
rect 10188 25929 10192 25956
rect 9682 25922 9716 25929
rect 9750 25922 9784 25929
rect 9818 25922 9852 25929
rect 9886 25922 9920 25929
rect 9954 25922 9988 25929
rect 10022 25922 10056 25929
rect 10090 25922 10124 25929
rect 10158 25922 10192 25929
rect 10260 25956 10298 25963
rect 10332 25956 10370 25963
rect 10404 25956 10442 25963
rect 10476 25956 10514 25963
rect 10548 25956 10586 25963
rect 10620 25956 10658 25963
rect 10692 25956 10730 25963
rect 10764 25956 10802 25963
rect 10836 25956 10874 25963
rect 10908 25956 10946 25963
rect 10980 25956 11018 25963
rect 11052 25956 11090 25963
rect 11124 25956 11162 25963
rect 11196 25956 11234 25963
rect 11268 25956 11306 25963
rect 11340 25956 11378 25963
rect 11412 25956 11450 25963
rect 10226 25922 10260 25929
rect 10294 25929 10298 25956
rect 10362 25929 10370 25956
rect 10430 25929 10442 25956
rect 10498 25929 10514 25956
rect 10566 25929 10586 25956
rect 10634 25929 10658 25956
rect 10702 25929 10730 25956
rect 10770 25929 10802 25956
rect 10294 25922 10328 25929
rect 10362 25922 10396 25929
rect 10430 25922 10464 25929
rect 10498 25922 10532 25929
rect 10566 25922 10600 25929
rect 10634 25922 10668 25929
rect 10702 25922 10736 25929
rect 10770 25922 10804 25929
rect 10838 25922 10872 25956
rect 10908 25929 10940 25956
rect 10980 25929 11008 25956
rect 11052 25929 11076 25956
rect 11124 25929 11144 25956
rect 11196 25929 11212 25956
rect 11268 25929 11280 25956
rect 11340 25929 11348 25956
rect 11412 25929 11416 25956
rect 10906 25922 10940 25929
rect 10974 25922 11008 25929
rect 11042 25922 11076 25929
rect 11110 25922 11144 25929
rect 11178 25922 11212 25929
rect 11246 25922 11280 25929
rect 11314 25922 11348 25929
rect 11382 25922 11416 25929
rect 11484 25956 11522 25963
rect 11556 25956 11594 25963
rect 11628 25956 11666 25963
rect 11700 25956 11738 25963
rect 11772 25956 11810 25963
rect 11844 25956 11882 25963
rect 11916 25956 11954 25963
rect 11988 25956 12026 25963
rect 12060 25956 12098 25963
rect 12132 25956 12170 25963
rect 12204 25956 12242 25963
rect 12276 25956 12314 25963
rect 12348 25956 12386 25963
rect 12420 25956 12458 25963
rect 12492 25956 12530 25963
rect 12564 25956 12602 25963
rect 12636 25956 12674 25963
rect 11450 25922 11484 25929
rect 11518 25929 11522 25956
rect 11586 25929 11594 25956
rect 11654 25929 11666 25956
rect 11722 25929 11738 25956
rect 11790 25929 11810 25956
rect 11858 25929 11882 25956
rect 11926 25929 11954 25956
rect 11994 25929 12026 25956
rect 11518 25922 11552 25929
rect 11586 25922 11620 25929
rect 11654 25922 11688 25929
rect 11722 25922 11756 25929
rect 11790 25922 11824 25929
rect 11858 25922 11892 25929
rect 11926 25922 11960 25929
rect 11994 25922 12028 25929
rect 12062 25922 12096 25956
rect 12132 25929 12164 25956
rect 12204 25929 12232 25956
rect 12276 25929 12300 25956
rect 12348 25929 12368 25956
rect 12420 25929 12436 25956
rect 12492 25929 12504 25956
rect 12564 25929 12572 25956
rect 12636 25929 12640 25956
rect 12130 25922 12164 25929
rect 12198 25922 12232 25929
rect 12266 25922 12300 25929
rect 12334 25922 12368 25929
rect 12402 25922 12436 25929
rect 12470 25922 12504 25929
rect 12538 25922 12572 25929
rect 12606 25922 12640 25929
rect 12708 25956 12746 25963
rect 12780 25956 12818 25963
rect 12852 25956 12890 25963
rect 12924 25956 12962 25963
rect 12996 25956 13034 25963
rect 13068 25956 13106 25963
rect 13140 25956 13178 25963
rect 13212 25956 13250 25963
rect 13284 25956 13322 25963
rect 13356 25956 13394 25963
rect 13428 25956 13466 25963
rect 13500 25956 13538 25963
rect 13572 25956 13610 25963
rect 13644 25956 13682 25963
rect 13716 25956 13754 25963
rect 13788 25956 13826 25963
rect 13860 25956 13898 25963
rect 12674 25922 12708 25929
rect 12742 25929 12746 25956
rect 12810 25929 12818 25956
rect 12878 25929 12890 25956
rect 12946 25929 12962 25956
rect 13014 25929 13034 25956
rect 13082 25929 13106 25956
rect 13150 25929 13178 25956
rect 13218 25929 13250 25956
rect 12742 25922 12776 25929
rect 12810 25922 12844 25929
rect 12878 25922 12912 25929
rect 12946 25922 12980 25929
rect 13014 25922 13048 25929
rect 13082 25922 13116 25929
rect 13150 25922 13184 25929
rect 13218 25922 13252 25929
rect 13286 25922 13320 25956
rect 13356 25929 13388 25956
rect 13428 25929 13456 25956
rect 13500 25929 13524 25956
rect 13572 25929 13592 25956
rect 13644 25929 13660 25956
rect 13716 25929 13728 25956
rect 13788 25929 13796 25956
rect 13860 25929 13864 25956
rect 13354 25922 13388 25929
rect 13422 25922 13456 25929
rect 13490 25922 13524 25929
rect 13558 25922 13592 25929
rect 13626 25922 13660 25929
rect 13694 25922 13728 25929
rect 13762 25922 13796 25929
rect 13830 25922 13864 25929
rect 13932 25956 13970 25963
rect 14004 25956 14042 25963
rect 14076 25956 14114 25963
rect 14148 25956 14186 25963
rect 14220 25956 14258 25963
rect 14292 25956 14330 25963
rect 14364 25956 14402 25963
rect 14436 25956 14474 25963
rect 14508 25956 14546 25963
rect 14580 25956 14618 25963
rect 14652 25956 14690 25963
rect 14724 25956 14962 25963
rect 13898 25922 13932 25929
rect 13966 25929 13970 25956
rect 14034 25929 14042 25956
rect 14102 25929 14114 25956
rect 14170 25929 14186 25956
rect 14238 25929 14258 25956
rect 14306 25929 14330 25956
rect 14374 25929 14402 25956
rect 14442 25929 14474 25956
rect 13966 25922 14000 25929
rect 14034 25922 14068 25929
rect 14102 25922 14136 25929
rect 14170 25922 14204 25929
rect 14238 25922 14272 25929
rect 14306 25922 14340 25929
rect 14374 25922 14408 25929
rect 14442 25922 14476 25929
rect 14510 25922 14544 25956
rect 14580 25929 14612 25956
rect 14652 25929 14680 25956
rect 14724 25929 14748 25956
rect 14578 25922 14612 25929
rect 14646 25922 14680 25929
rect 14714 25922 14748 25929
rect 14782 25922 14816 25956
rect 14850 25922 14884 25956
rect 14918 25922 14962 25956
rect 49 25889 14962 25922
rect 49 25884 243 25889
rect 277 25884 316 25889
rect 350 25884 389 25889
rect 423 25884 462 25889
rect 496 25884 535 25889
rect 569 25884 608 25889
rect 642 25884 681 25889
rect 715 25884 754 25889
rect 788 25884 827 25889
rect 861 25884 900 25889
rect 934 25884 973 25889
rect 1007 25884 1046 25889
rect 1080 25884 1119 25889
rect 1153 25884 1192 25889
rect 1226 25884 1265 25889
rect 1299 25884 1338 25889
rect 1372 25884 1411 25889
rect 1445 25884 1484 25889
rect 49 25850 69 25884
rect 103 25850 138 25884
rect 172 25850 207 25884
rect 241 25855 243 25884
rect 310 25855 316 25884
rect 379 25855 389 25884
rect 448 25855 462 25884
rect 517 25855 535 25884
rect 586 25855 608 25884
rect 655 25855 681 25884
rect 724 25855 754 25884
rect 793 25855 827 25884
rect 241 25850 276 25855
rect 310 25850 345 25855
rect 379 25850 414 25855
rect 448 25850 483 25855
rect 517 25850 552 25855
rect 586 25850 621 25855
rect 655 25850 690 25855
rect 724 25850 759 25855
rect 793 25850 828 25855
rect 862 25850 897 25884
rect 934 25855 966 25884
rect 1007 25855 1035 25884
rect 1080 25855 1104 25884
rect 1153 25855 1173 25884
rect 1226 25855 1242 25884
rect 1299 25855 1311 25884
rect 1372 25855 1380 25884
rect 1445 25855 1449 25884
rect 931 25850 966 25855
rect 1000 25850 1035 25855
rect 1069 25850 1104 25855
rect 1138 25850 1173 25855
rect 1207 25850 1242 25855
rect 1276 25850 1311 25855
rect 1345 25850 1380 25855
rect 1414 25850 1449 25855
rect 1483 25855 1484 25884
rect 1518 25884 1557 25889
rect 1591 25884 1630 25889
rect 1664 25884 1703 25889
rect 1737 25884 1776 25889
rect 1810 25884 1849 25889
rect 1883 25884 1922 25889
rect 1956 25884 1995 25889
rect 2029 25884 2068 25889
rect 2102 25884 2141 25889
rect 2175 25884 2214 25889
rect 2248 25884 2287 25889
rect 2321 25884 2360 25889
rect 2394 25884 2433 25889
rect 2467 25884 2506 25889
rect 2540 25884 2579 25889
rect 2613 25884 2652 25889
rect 2686 25884 2725 25889
rect 1483 25850 1518 25855
rect 1552 25855 1557 25884
rect 1621 25855 1630 25884
rect 1690 25855 1703 25884
rect 1759 25855 1776 25884
rect 1828 25855 1849 25884
rect 1897 25855 1922 25884
rect 1966 25855 1995 25884
rect 2035 25855 2068 25884
rect 1552 25850 1587 25855
rect 1621 25850 1656 25855
rect 1690 25850 1725 25855
rect 1759 25850 1794 25855
rect 1828 25850 1863 25855
rect 1897 25850 1932 25855
rect 1966 25850 2001 25855
rect 2035 25850 2070 25855
rect 2104 25850 2139 25884
rect 2175 25855 2208 25884
rect 2248 25855 2277 25884
rect 2321 25855 2346 25884
rect 2394 25855 2415 25884
rect 2467 25855 2484 25884
rect 2540 25855 2553 25884
rect 2613 25855 2622 25884
rect 2686 25855 2691 25884
rect 2173 25850 2208 25855
rect 2242 25850 2277 25855
rect 2311 25850 2346 25855
rect 2380 25850 2415 25855
rect 2449 25850 2484 25855
rect 2518 25850 2553 25855
rect 2587 25850 2622 25855
rect 2656 25850 2691 25855
rect 2759 25884 2798 25889
rect 2832 25884 2871 25889
rect 2905 25884 2944 25889
rect 2978 25884 3017 25889
rect 3051 25884 3090 25889
rect 3124 25884 3163 25889
rect 3197 25884 3236 25889
rect 3270 25884 3309 25889
rect 3343 25884 3382 25889
rect 3416 25884 3455 25889
rect 3489 25884 3528 25889
rect 3562 25884 3601 25889
rect 3635 25884 3674 25889
rect 3708 25884 3746 25889
rect 3780 25884 3818 25889
rect 3852 25884 3890 25889
rect 3924 25884 3962 25889
rect 3996 25884 4034 25889
rect 4068 25884 4106 25889
rect 2759 25855 2760 25884
rect 2725 25850 2760 25855
rect 2794 25855 2798 25884
rect 2863 25855 2871 25884
rect 2932 25855 2944 25884
rect 3001 25855 3017 25884
rect 3070 25855 3090 25884
rect 3139 25855 3163 25884
rect 3208 25855 3236 25884
rect 3277 25855 3309 25884
rect 2794 25850 2829 25855
rect 2863 25850 2898 25855
rect 2932 25850 2967 25855
rect 3001 25850 3036 25855
rect 3070 25850 3105 25855
rect 3139 25850 3174 25855
rect 3208 25850 3243 25855
rect 3277 25850 3312 25855
rect 3346 25850 3381 25884
rect 3416 25855 3450 25884
rect 3489 25855 3519 25884
rect 3562 25855 3588 25884
rect 3635 25855 3657 25884
rect 3708 25855 3726 25884
rect 3780 25855 3795 25884
rect 3852 25855 3864 25884
rect 3924 25855 3933 25884
rect 3996 25855 4002 25884
rect 4068 25855 4071 25884
rect 3415 25850 3450 25855
rect 3484 25850 3519 25855
rect 3553 25850 3588 25855
rect 3622 25850 3657 25855
rect 3691 25850 3726 25855
rect 3760 25850 3795 25855
rect 3829 25850 3864 25855
rect 3898 25850 3933 25855
rect 3967 25850 4002 25855
rect 4036 25850 4071 25855
rect 4105 25855 4106 25884
rect 4140 25884 4178 25889
rect 4212 25884 4250 25889
rect 4284 25884 4322 25889
rect 4356 25884 4394 25889
rect 4428 25884 4466 25889
rect 4500 25884 4538 25889
rect 4572 25884 4610 25889
rect 4644 25884 4682 25889
rect 4716 25884 4754 25889
rect 4788 25884 4826 25889
rect 4860 25884 4898 25889
rect 4932 25884 4970 25889
rect 5004 25884 5042 25889
rect 5076 25884 5114 25889
rect 5148 25884 5186 25889
rect 5220 25884 5258 25889
rect 5292 25884 5330 25889
rect 4105 25850 4140 25855
rect 4174 25855 4178 25884
rect 4242 25855 4250 25884
rect 4310 25855 4322 25884
rect 4378 25855 4394 25884
rect 4446 25855 4466 25884
rect 4514 25855 4538 25884
rect 4582 25855 4610 25884
rect 4650 25855 4682 25884
rect 4174 25850 4208 25855
rect 4242 25850 4276 25855
rect 4310 25850 4344 25855
rect 4378 25850 4412 25855
rect 4446 25850 4480 25855
rect 4514 25850 4548 25855
rect 4582 25850 4616 25855
rect 4650 25850 4684 25855
rect 4718 25850 4752 25884
rect 4788 25855 4820 25884
rect 4860 25855 4888 25884
rect 4932 25855 4956 25884
rect 5004 25855 5024 25884
rect 5076 25855 5092 25884
rect 5148 25855 5160 25884
rect 5220 25855 5228 25884
rect 5292 25855 5296 25884
rect 4786 25850 4820 25855
rect 4854 25850 4888 25855
rect 4922 25850 4956 25855
rect 4990 25850 5024 25855
rect 5058 25850 5092 25855
rect 5126 25850 5160 25855
rect 5194 25850 5228 25855
rect 5262 25850 5296 25855
rect 5364 25884 5402 25889
rect 5436 25884 5474 25889
rect 5508 25884 5546 25889
rect 5580 25884 5618 25889
rect 5652 25884 5690 25889
rect 5724 25884 5762 25889
rect 5796 25884 5834 25889
rect 5868 25884 5906 25889
rect 5940 25884 5978 25889
rect 6012 25884 6050 25889
rect 6084 25884 6122 25889
rect 6156 25884 6194 25889
rect 6228 25884 6266 25889
rect 6300 25884 6338 25889
rect 6372 25884 6410 25889
rect 6444 25884 6482 25889
rect 6516 25884 6554 25889
rect 5330 25850 5364 25855
rect 5398 25855 5402 25884
rect 5466 25855 5474 25884
rect 5534 25855 5546 25884
rect 5602 25855 5618 25884
rect 5670 25855 5690 25884
rect 5738 25855 5762 25884
rect 5806 25855 5834 25884
rect 5874 25855 5906 25884
rect 5398 25850 5432 25855
rect 5466 25850 5500 25855
rect 5534 25850 5568 25855
rect 5602 25850 5636 25855
rect 5670 25850 5704 25855
rect 5738 25850 5772 25855
rect 5806 25850 5840 25855
rect 5874 25850 5908 25855
rect 5942 25850 5976 25884
rect 6012 25855 6044 25884
rect 6084 25855 6112 25884
rect 6156 25855 6180 25884
rect 6228 25855 6248 25884
rect 6300 25855 6316 25884
rect 6372 25855 6384 25884
rect 6444 25855 6452 25884
rect 6516 25855 6520 25884
rect 6010 25850 6044 25855
rect 6078 25850 6112 25855
rect 6146 25850 6180 25855
rect 6214 25850 6248 25855
rect 6282 25850 6316 25855
rect 6350 25850 6384 25855
rect 6418 25850 6452 25855
rect 6486 25850 6520 25855
rect 6588 25884 6626 25889
rect 6660 25884 6698 25889
rect 6732 25884 6770 25889
rect 6804 25884 6842 25889
rect 6876 25884 6914 25889
rect 6948 25884 6986 25889
rect 7020 25884 7058 25889
rect 7092 25884 7130 25889
rect 7164 25884 7202 25889
rect 7236 25884 7274 25889
rect 7308 25884 7346 25889
rect 7380 25884 7418 25889
rect 7452 25884 7490 25889
rect 7524 25884 7562 25889
rect 7596 25884 7634 25889
rect 7668 25884 7706 25889
rect 7740 25884 7778 25889
rect 6554 25850 6588 25855
rect 6622 25855 6626 25884
rect 6690 25855 6698 25884
rect 6758 25855 6770 25884
rect 6826 25855 6842 25884
rect 6894 25855 6914 25884
rect 6962 25855 6986 25884
rect 7030 25855 7058 25884
rect 7098 25855 7130 25884
rect 6622 25850 6656 25855
rect 6690 25850 6724 25855
rect 6758 25850 6792 25855
rect 6826 25850 6860 25855
rect 6894 25850 6928 25855
rect 6962 25850 6996 25855
rect 7030 25850 7064 25855
rect 7098 25850 7132 25855
rect 7166 25850 7200 25884
rect 7236 25855 7268 25884
rect 7308 25855 7336 25884
rect 7380 25855 7404 25884
rect 7452 25855 7472 25884
rect 7524 25855 7540 25884
rect 7596 25855 7608 25884
rect 7668 25855 7676 25884
rect 7740 25855 7744 25884
rect 7234 25850 7268 25855
rect 7302 25850 7336 25855
rect 7370 25850 7404 25855
rect 7438 25850 7472 25855
rect 7506 25850 7540 25855
rect 7574 25850 7608 25855
rect 7642 25850 7676 25855
rect 7710 25850 7744 25855
rect 7812 25884 7850 25889
rect 7884 25884 7922 25889
rect 7956 25884 7994 25889
rect 8028 25884 8066 25889
rect 8100 25884 8138 25889
rect 8172 25884 8210 25889
rect 8244 25884 8282 25889
rect 8316 25884 8354 25889
rect 8388 25884 8426 25889
rect 8460 25884 8498 25889
rect 8532 25884 8570 25889
rect 8604 25884 8642 25889
rect 8676 25884 8714 25889
rect 8748 25884 8786 25889
rect 8820 25884 8858 25889
rect 8892 25884 8930 25889
rect 8964 25884 9002 25889
rect 7778 25850 7812 25855
rect 7846 25855 7850 25884
rect 7914 25855 7922 25884
rect 7982 25855 7994 25884
rect 8050 25855 8066 25884
rect 8118 25855 8138 25884
rect 8186 25855 8210 25884
rect 8254 25855 8282 25884
rect 8322 25855 8354 25884
rect 7846 25850 7880 25855
rect 7914 25850 7948 25855
rect 7982 25850 8016 25855
rect 8050 25850 8084 25855
rect 8118 25850 8152 25855
rect 8186 25850 8220 25855
rect 8254 25850 8288 25855
rect 8322 25850 8356 25855
rect 8390 25850 8424 25884
rect 8460 25855 8492 25884
rect 8532 25855 8560 25884
rect 8604 25855 8628 25884
rect 8676 25855 8696 25884
rect 8748 25855 8764 25884
rect 8820 25855 8832 25884
rect 8892 25855 8900 25884
rect 8964 25855 8968 25884
rect 8458 25850 8492 25855
rect 8526 25850 8560 25855
rect 8594 25850 8628 25855
rect 8662 25850 8696 25855
rect 8730 25850 8764 25855
rect 8798 25850 8832 25855
rect 8866 25850 8900 25855
rect 8934 25850 8968 25855
rect 9036 25884 9074 25889
rect 9108 25884 9146 25889
rect 9180 25884 9218 25889
rect 9252 25884 9290 25889
rect 9324 25884 9362 25889
rect 9396 25884 9434 25889
rect 9468 25884 9506 25889
rect 9540 25884 9578 25889
rect 9612 25884 9650 25889
rect 9684 25884 9722 25889
rect 9756 25884 9794 25889
rect 9828 25884 9866 25889
rect 9900 25884 9938 25889
rect 9972 25884 10010 25889
rect 10044 25884 10082 25889
rect 10116 25884 10154 25889
rect 10188 25884 10226 25889
rect 9002 25850 9036 25855
rect 9070 25855 9074 25884
rect 9138 25855 9146 25884
rect 9206 25855 9218 25884
rect 9274 25855 9290 25884
rect 9342 25855 9362 25884
rect 9410 25855 9434 25884
rect 9478 25855 9506 25884
rect 9546 25855 9578 25884
rect 9070 25850 9104 25855
rect 9138 25850 9172 25855
rect 9206 25850 9240 25855
rect 9274 25850 9308 25855
rect 9342 25850 9376 25855
rect 9410 25850 9444 25855
rect 9478 25850 9512 25855
rect 9546 25850 9580 25855
rect 9614 25850 9648 25884
rect 9684 25855 9716 25884
rect 9756 25855 9784 25884
rect 9828 25855 9852 25884
rect 9900 25855 9920 25884
rect 9972 25855 9988 25884
rect 10044 25855 10056 25884
rect 10116 25855 10124 25884
rect 10188 25855 10192 25884
rect 9682 25850 9716 25855
rect 9750 25850 9784 25855
rect 9818 25850 9852 25855
rect 9886 25850 9920 25855
rect 9954 25850 9988 25855
rect 10022 25850 10056 25855
rect 10090 25850 10124 25855
rect 10158 25850 10192 25855
rect 10260 25884 10298 25889
rect 10332 25884 10370 25889
rect 10404 25884 10442 25889
rect 10476 25884 10514 25889
rect 10548 25884 10586 25889
rect 10620 25884 10658 25889
rect 10692 25884 10730 25889
rect 10764 25884 10802 25889
rect 10836 25884 10874 25889
rect 10908 25884 10946 25889
rect 10980 25884 11018 25889
rect 11052 25884 11090 25889
rect 11124 25884 11162 25889
rect 11196 25884 11234 25889
rect 11268 25884 11306 25889
rect 11340 25884 11378 25889
rect 11412 25884 11450 25889
rect 10226 25850 10260 25855
rect 10294 25855 10298 25884
rect 10362 25855 10370 25884
rect 10430 25855 10442 25884
rect 10498 25855 10514 25884
rect 10566 25855 10586 25884
rect 10634 25855 10658 25884
rect 10702 25855 10730 25884
rect 10770 25855 10802 25884
rect 10294 25850 10328 25855
rect 10362 25850 10396 25855
rect 10430 25850 10464 25855
rect 10498 25850 10532 25855
rect 10566 25850 10600 25855
rect 10634 25850 10668 25855
rect 10702 25850 10736 25855
rect 10770 25850 10804 25855
rect 10838 25850 10872 25884
rect 10908 25855 10940 25884
rect 10980 25855 11008 25884
rect 11052 25855 11076 25884
rect 11124 25855 11144 25884
rect 11196 25855 11212 25884
rect 11268 25855 11280 25884
rect 11340 25855 11348 25884
rect 11412 25855 11416 25884
rect 10906 25850 10940 25855
rect 10974 25850 11008 25855
rect 11042 25850 11076 25855
rect 11110 25850 11144 25855
rect 11178 25850 11212 25855
rect 11246 25850 11280 25855
rect 11314 25850 11348 25855
rect 11382 25850 11416 25855
rect 11484 25884 11522 25889
rect 11556 25884 11594 25889
rect 11628 25884 11666 25889
rect 11700 25884 11738 25889
rect 11772 25884 11810 25889
rect 11844 25884 11882 25889
rect 11916 25884 11954 25889
rect 11988 25884 12026 25889
rect 12060 25884 12098 25889
rect 12132 25884 12170 25889
rect 12204 25884 12242 25889
rect 12276 25884 12314 25889
rect 12348 25884 12386 25889
rect 12420 25884 12458 25889
rect 12492 25884 12530 25889
rect 12564 25884 12602 25889
rect 12636 25884 12674 25889
rect 11450 25850 11484 25855
rect 11518 25855 11522 25884
rect 11586 25855 11594 25884
rect 11654 25855 11666 25884
rect 11722 25855 11738 25884
rect 11790 25855 11810 25884
rect 11858 25855 11882 25884
rect 11926 25855 11954 25884
rect 11994 25855 12026 25884
rect 11518 25850 11552 25855
rect 11586 25850 11620 25855
rect 11654 25850 11688 25855
rect 11722 25850 11756 25855
rect 11790 25850 11824 25855
rect 11858 25850 11892 25855
rect 11926 25850 11960 25855
rect 11994 25850 12028 25855
rect 12062 25850 12096 25884
rect 12132 25855 12164 25884
rect 12204 25855 12232 25884
rect 12276 25855 12300 25884
rect 12348 25855 12368 25884
rect 12420 25855 12436 25884
rect 12492 25855 12504 25884
rect 12564 25855 12572 25884
rect 12636 25855 12640 25884
rect 12130 25850 12164 25855
rect 12198 25850 12232 25855
rect 12266 25850 12300 25855
rect 12334 25850 12368 25855
rect 12402 25850 12436 25855
rect 12470 25850 12504 25855
rect 12538 25850 12572 25855
rect 12606 25850 12640 25855
rect 12708 25884 12746 25889
rect 12780 25884 12818 25889
rect 12852 25884 12890 25889
rect 12924 25884 12962 25889
rect 12996 25884 13034 25889
rect 13068 25884 13106 25889
rect 13140 25884 13178 25889
rect 13212 25884 13250 25889
rect 13284 25884 13322 25889
rect 13356 25884 13394 25889
rect 13428 25884 13466 25889
rect 13500 25884 13538 25889
rect 13572 25884 13610 25889
rect 13644 25884 13682 25889
rect 13716 25884 13754 25889
rect 13788 25884 13826 25889
rect 13860 25884 13898 25889
rect 12674 25850 12708 25855
rect 12742 25855 12746 25884
rect 12810 25855 12818 25884
rect 12878 25855 12890 25884
rect 12946 25855 12962 25884
rect 13014 25855 13034 25884
rect 13082 25855 13106 25884
rect 13150 25855 13178 25884
rect 13218 25855 13250 25884
rect 12742 25850 12776 25855
rect 12810 25850 12844 25855
rect 12878 25850 12912 25855
rect 12946 25850 12980 25855
rect 13014 25850 13048 25855
rect 13082 25850 13116 25855
rect 13150 25850 13184 25855
rect 13218 25850 13252 25855
rect 13286 25850 13320 25884
rect 13356 25855 13388 25884
rect 13428 25855 13456 25884
rect 13500 25855 13524 25884
rect 13572 25855 13592 25884
rect 13644 25855 13660 25884
rect 13716 25855 13728 25884
rect 13788 25855 13796 25884
rect 13860 25855 13864 25884
rect 13354 25850 13388 25855
rect 13422 25850 13456 25855
rect 13490 25850 13524 25855
rect 13558 25850 13592 25855
rect 13626 25850 13660 25855
rect 13694 25850 13728 25855
rect 13762 25850 13796 25855
rect 13830 25850 13864 25855
rect 13932 25884 13970 25889
rect 14004 25884 14042 25889
rect 14076 25884 14114 25889
rect 14148 25884 14186 25889
rect 14220 25884 14258 25889
rect 14292 25884 14330 25889
rect 14364 25884 14402 25889
rect 14436 25884 14474 25889
rect 14508 25884 14546 25889
rect 14580 25884 14618 25889
rect 14652 25884 14690 25889
rect 14724 25884 14962 25889
rect 13898 25850 13932 25855
rect 13966 25855 13970 25884
rect 14034 25855 14042 25884
rect 14102 25855 14114 25884
rect 14170 25855 14186 25884
rect 14238 25855 14258 25884
rect 14306 25855 14330 25884
rect 14374 25855 14402 25884
rect 14442 25855 14474 25884
rect 13966 25850 14000 25855
rect 14034 25850 14068 25855
rect 14102 25850 14136 25855
rect 14170 25850 14204 25855
rect 14238 25850 14272 25855
rect 14306 25850 14340 25855
rect 14374 25850 14408 25855
rect 14442 25850 14476 25855
rect 14510 25850 14544 25884
rect 14580 25855 14612 25884
rect 14652 25855 14680 25884
rect 14724 25855 14748 25884
rect 14578 25850 14612 25855
rect 14646 25850 14680 25855
rect 14714 25850 14748 25855
rect 14782 25850 14816 25884
rect 14850 25850 14884 25884
rect 14918 25850 14962 25884
rect 49 25815 14962 25850
rect 49 25812 243 25815
rect 277 25812 316 25815
rect 350 25812 389 25815
rect 423 25812 462 25815
rect 496 25812 535 25815
rect 569 25812 608 25815
rect 642 25812 681 25815
rect 715 25812 754 25815
rect 788 25812 827 25815
rect 861 25812 900 25815
rect 934 25812 973 25815
rect 1007 25812 1046 25815
rect 1080 25812 1119 25815
rect 1153 25812 1192 25815
rect 1226 25812 1265 25815
rect 1299 25812 1338 25815
rect 1372 25812 1411 25815
rect 1445 25812 1484 25815
rect 49 25778 69 25812
rect 103 25778 138 25812
rect 172 25778 207 25812
rect 241 25781 243 25812
rect 310 25781 316 25812
rect 379 25781 389 25812
rect 448 25781 462 25812
rect 517 25781 535 25812
rect 586 25781 608 25812
rect 655 25781 681 25812
rect 724 25781 754 25812
rect 793 25781 827 25812
rect 241 25778 276 25781
rect 310 25778 345 25781
rect 379 25778 414 25781
rect 448 25778 483 25781
rect 517 25778 552 25781
rect 586 25778 621 25781
rect 655 25778 690 25781
rect 724 25778 759 25781
rect 793 25778 828 25781
rect 862 25778 897 25812
rect 934 25781 966 25812
rect 1007 25781 1035 25812
rect 1080 25781 1104 25812
rect 1153 25781 1173 25812
rect 1226 25781 1242 25812
rect 1299 25781 1311 25812
rect 1372 25781 1380 25812
rect 1445 25781 1449 25812
rect 931 25778 966 25781
rect 1000 25778 1035 25781
rect 1069 25778 1104 25781
rect 1138 25778 1173 25781
rect 1207 25778 1242 25781
rect 1276 25778 1311 25781
rect 1345 25778 1380 25781
rect 1414 25778 1449 25781
rect 1483 25781 1484 25812
rect 1518 25812 1557 25815
rect 1591 25812 1630 25815
rect 1664 25812 1703 25815
rect 1737 25812 1776 25815
rect 1810 25812 1849 25815
rect 1883 25812 1922 25815
rect 1956 25812 1995 25815
rect 2029 25812 2068 25815
rect 2102 25812 2141 25815
rect 2175 25812 2214 25815
rect 2248 25812 2287 25815
rect 2321 25812 2360 25815
rect 2394 25812 2433 25815
rect 2467 25812 2506 25815
rect 2540 25812 2579 25815
rect 2613 25812 2652 25815
rect 2686 25812 2725 25815
rect 1483 25778 1518 25781
rect 1552 25781 1557 25812
rect 1621 25781 1630 25812
rect 1690 25781 1703 25812
rect 1759 25781 1776 25812
rect 1828 25781 1849 25812
rect 1897 25781 1922 25812
rect 1966 25781 1995 25812
rect 2035 25781 2068 25812
rect 1552 25778 1587 25781
rect 1621 25778 1656 25781
rect 1690 25778 1725 25781
rect 1759 25778 1794 25781
rect 1828 25778 1863 25781
rect 1897 25778 1932 25781
rect 1966 25778 2001 25781
rect 2035 25778 2070 25781
rect 2104 25778 2139 25812
rect 2175 25781 2208 25812
rect 2248 25781 2277 25812
rect 2321 25781 2346 25812
rect 2394 25781 2415 25812
rect 2467 25781 2484 25812
rect 2540 25781 2553 25812
rect 2613 25781 2622 25812
rect 2686 25781 2691 25812
rect 2173 25778 2208 25781
rect 2242 25778 2277 25781
rect 2311 25778 2346 25781
rect 2380 25778 2415 25781
rect 2449 25778 2484 25781
rect 2518 25778 2553 25781
rect 2587 25778 2622 25781
rect 2656 25778 2691 25781
rect 2759 25812 2798 25815
rect 2832 25812 2871 25815
rect 2905 25812 2944 25815
rect 2978 25812 3017 25815
rect 3051 25812 3090 25815
rect 3124 25812 3163 25815
rect 3197 25812 3236 25815
rect 3270 25812 3309 25815
rect 3343 25812 3382 25815
rect 3416 25812 3455 25815
rect 3489 25812 3528 25815
rect 3562 25812 3601 25815
rect 3635 25812 3674 25815
rect 3708 25812 3746 25815
rect 3780 25812 3818 25815
rect 3852 25812 3890 25815
rect 3924 25812 3962 25815
rect 3996 25812 4034 25815
rect 4068 25812 4106 25815
rect 2759 25781 2760 25812
rect 2725 25778 2760 25781
rect 2794 25781 2798 25812
rect 2863 25781 2871 25812
rect 2932 25781 2944 25812
rect 3001 25781 3017 25812
rect 3070 25781 3090 25812
rect 3139 25781 3163 25812
rect 3208 25781 3236 25812
rect 3277 25781 3309 25812
rect 2794 25778 2829 25781
rect 2863 25778 2898 25781
rect 2932 25778 2967 25781
rect 3001 25778 3036 25781
rect 3070 25778 3105 25781
rect 3139 25778 3174 25781
rect 3208 25778 3243 25781
rect 3277 25778 3312 25781
rect 3346 25778 3381 25812
rect 3416 25781 3450 25812
rect 3489 25781 3519 25812
rect 3562 25781 3588 25812
rect 3635 25781 3657 25812
rect 3708 25781 3726 25812
rect 3780 25781 3795 25812
rect 3852 25781 3864 25812
rect 3924 25781 3933 25812
rect 3996 25781 4002 25812
rect 4068 25781 4071 25812
rect 3415 25778 3450 25781
rect 3484 25778 3519 25781
rect 3553 25778 3588 25781
rect 3622 25778 3657 25781
rect 3691 25778 3726 25781
rect 3760 25778 3795 25781
rect 3829 25778 3864 25781
rect 3898 25778 3933 25781
rect 3967 25778 4002 25781
rect 4036 25778 4071 25781
rect 4105 25781 4106 25812
rect 4140 25812 4178 25815
rect 4212 25812 4250 25815
rect 4284 25812 4322 25815
rect 4356 25812 4394 25815
rect 4428 25812 4466 25815
rect 4500 25812 4538 25815
rect 4572 25812 4610 25815
rect 4644 25812 4682 25815
rect 4716 25812 4754 25815
rect 4788 25812 4826 25815
rect 4860 25812 4898 25815
rect 4932 25812 4970 25815
rect 5004 25812 5042 25815
rect 5076 25812 5114 25815
rect 5148 25812 5186 25815
rect 5220 25812 5258 25815
rect 5292 25812 5330 25815
rect 4105 25778 4140 25781
rect 4174 25781 4178 25812
rect 4242 25781 4250 25812
rect 4310 25781 4322 25812
rect 4378 25781 4394 25812
rect 4446 25781 4466 25812
rect 4514 25781 4538 25812
rect 4582 25781 4610 25812
rect 4650 25781 4682 25812
rect 4174 25778 4208 25781
rect 4242 25778 4276 25781
rect 4310 25778 4344 25781
rect 4378 25778 4412 25781
rect 4446 25778 4480 25781
rect 4514 25778 4548 25781
rect 4582 25778 4616 25781
rect 4650 25778 4684 25781
rect 4718 25778 4752 25812
rect 4788 25781 4820 25812
rect 4860 25781 4888 25812
rect 4932 25781 4956 25812
rect 5004 25781 5024 25812
rect 5076 25781 5092 25812
rect 5148 25781 5160 25812
rect 5220 25781 5228 25812
rect 5292 25781 5296 25812
rect 4786 25778 4820 25781
rect 4854 25778 4888 25781
rect 4922 25778 4956 25781
rect 4990 25778 5024 25781
rect 5058 25778 5092 25781
rect 5126 25778 5160 25781
rect 5194 25778 5228 25781
rect 5262 25778 5296 25781
rect 5364 25812 5402 25815
rect 5436 25812 5474 25815
rect 5508 25812 5546 25815
rect 5580 25812 5618 25815
rect 5652 25812 5690 25815
rect 5724 25812 5762 25815
rect 5796 25812 5834 25815
rect 5868 25812 5906 25815
rect 5940 25812 5978 25815
rect 6012 25812 6050 25815
rect 6084 25812 6122 25815
rect 6156 25812 6194 25815
rect 6228 25812 6266 25815
rect 6300 25812 6338 25815
rect 6372 25812 6410 25815
rect 6444 25812 6482 25815
rect 6516 25812 6554 25815
rect 5330 25778 5364 25781
rect 5398 25781 5402 25812
rect 5466 25781 5474 25812
rect 5534 25781 5546 25812
rect 5602 25781 5618 25812
rect 5670 25781 5690 25812
rect 5738 25781 5762 25812
rect 5806 25781 5834 25812
rect 5874 25781 5906 25812
rect 5398 25778 5432 25781
rect 5466 25778 5500 25781
rect 5534 25778 5568 25781
rect 5602 25778 5636 25781
rect 5670 25778 5704 25781
rect 5738 25778 5772 25781
rect 5806 25778 5840 25781
rect 5874 25778 5908 25781
rect 5942 25778 5976 25812
rect 6012 25781 6044 25812
rect 6084 25781 6112 25812
rect 6156 25781 6180 25812
rect 6228 25781 6248 25812
rect 6300 25781 6316 25812
rect 6372 25781 6384 25812
rect 6444 25781 6452 25812
rect 6516 25781 6520 25812
rect 6010 25778 6044 25781
rect 6078 25778 6112 25781
rect 6146 25778 6180 25781
rect 6214 25778 6248 25781
rect 6282 25778 6316 25781
rect 6350 25778 6384 25781
rect 6418 25778 6452 25781
rect 6486 25778 6520 25781
rect 6588 25812 6626 25815
rect 6660 25812 6698 25815
rect 6732 25812 6770 25815
rect 6804 25812 6842 25815
rect 6876 25812 6914 25815
rect 6948 25812 6986 25815
rect 7020 25812 7058 25815
rect 7092 25812 7130 25815
rect 7164 25812 7202 25815
rect 7236 25812 7274 25815
rect 7308 25812 7346 25815
rect 7380 25812 7418 25815
rect 7452 25812 7490 25815
rect 7524 25812 7562 25815
rect 7596 25812 7634 25815
rect 7668 25812 7706 25815
rect 7740 25812 7778 25815
rect 6554 25778 6588 25781
rect 6622 25781 6626 25812
rect 6690 25781 6698 25812
rect 6758 25781 6770 25812
rect 6826 25781 6842 25812
rect 6894 25781 6914 25812
rect 6962 25781 6986 25812
rect 7030 25781 7058 25812
rect 7098 25781 7130 25812
rect 6622 25778 6656 25781
rect 6690 25778 6724 25781
rect 6758 25778 6792 25781
rect 6826 25778 6860 25781
rect 6894 25778 6928 25781
rect 6962 25778 6996 25781
rect 7030 25778 7064 25781
rect 7098 25778 7132 25781
rect 7166 25778 7200 25812
rect 7236 25781 7268 25812
rect 7308 25781 7336 25812
rect 7380 25781 7404 25812
rect 7452 25781 7472 25812
rect 7524 25781 7540 25812
rect 7596 25781 7608 25812
rect 7668 25781 7676 25812
rect 7740 25781 7744 25812
rect 7234 25778 7268 25781
rect 7302 25778 7336 25781
rect 7370 25778 7404 25781
rect 7438 25778 7472 25781
rect 7506 25778 7540 25781
rect 7574 25778 7608 25781
rect 7642 25778 7676 25781
rect 7710 25778 7744 25781
rect 7812 25812 7850 25815
rect 7884 25812 7922 25815
rect 7956 25812 7994 25815
rect 8028 25812 8066 25815
rect 8100 25812 8138 25815
rect 8172 25812 8210 25815
rect 8244 25812 8282 25815
rect 8316 25812 8354 25815
rect 8388 25812 8426 25815
rect 8460 25812 8498 25815
rect 8532 25812 8570 25815
rect 8604 25812 8642 25815
rect 8676 25812 8714 25815
rect 8748 25812 8786 25815
rect 8820 25812 8858 25815
rect 8892 25812 8930 25815
rect 8964 25812 9002 25815
rect 7778 25778 7812 25781
rect 7846 25781 7850 25812
rect 7914 25781 7922 25812
rect 7982 25781 7994 25812
rect 8050 25781 8066 25812
rect 8118 25781 8138 25812
rect 8186 25781 8210 25812
rect 8254 25781 8282 25812
rect 8322 25781 8354 25812
rect 7846 25778 7880 25781
rect 7914 25778 7948 25781
rect 7982 25778 8016 25781
rect 8050 25778 8084 25781
rect 8118 25778 8152 25781
rect 8186 25778 8220 25781
rect 8254 25778 8288 25781
rect 8322 25778 8356 25781
rect 8390 25778 8424 25812
rect 8460 25781 8492 25812
rect 8532 25781 8560 25812
rect 8604 25781 8628 25812
rect 8676 25781 8696 25812
rect 8748 25781 8764 25812
rect 8820 25781 8832 25812
rect 8892 25781 8900 25812
rect 8964 25781 8968 25812
rect 8458 25778 8492 25781
rect 8526 25778 8560 25781
rect 8594 25778 8628 25781
rect 8662 25778 8696 25781
rect 8730 25778 8764 25781
rect 8798 25778 8832 25781
rect 8866 25778 8900 25781
rect 8934 25778 8968 25781
rect 9036 25812 9074 25815
rect 9108 25812 9146 25815
rect 9180 25812 9218 25815
rect 9252 25812 9290 25815
rect 9324 25812 9362 25815
rect 9396 25812 9434 25815
rect 9468 25812 9506 25815
rect 9540 25812 9578 25815
rect 9612 25812 9650 25815
rect 9684 25812 9722 25815
rect 9756 25812 9794 25815
rect 9828 25812 9866 25815
rect 9900 25812 9938 25815
rect 9972 25812 10010 25815
rect 10044 25812 10082 25815
rect 10116 25812 10154 25815
rect 10188 25812 10226 25815
rect 9002 25778 9036 25781
rect 9070 25781 9074 25812
rect 9138 25781 9146 25812
rect 9206 25781 9218 25812
rect 9274 25781 9290 25812
rect 9342 25781 9362 25812
rect 9410 25781 9434 25812
rect 9478 25781 9506 25812
rect 9546 25781 9578 25812
rect 9070 25778 9104 25781
rect 9138 25778 9172 25781
rect 9206 25778 9240 25781
rect 9274 25778 9308 25781
rect 9342 25778 9376 25781
rect 9410 25778 9444 25781
rect 9478 25778 9512 25781
rect 9546 25778 9580 25781
rect 9614 25778 9648 25812
rect 9684 25781 9716 25812
rect 9756 25781 9784 25812
rect 9828 25781 9852 25812
rect 9900 25781 9920 25812
rect 9972 25781 9988 25812
rect 10044 25781 10056 25812
rect 10116 25781 10124 25812
rect 10188 25781 10192 25812
rect 9682 25778 9716 25781
rect 9750 25778 9784 25781
rect 9818 25778 9852 25781
rect 9886 25778 9920 25781
rect 9954 25778 9988 25781
rect 10022 25778 10056 25781
rect 10090 25778 10124 25781
rect 10158 25778 10192 25781
rect 10260 25812 10298 25815
rect 10332 25812 10370 25815
rect 10404 25812 10442 25815
rect 10476 25812 10514 25815
rect 10548 25812 10586 25815
rect 10620 25812 10658 25815
rect 10692 25812 10730 25815
rect 10764 25812 10802 25815
rect 10836 25812 10874 25815
rect 10908 25812 10946 25815
rect 10980 25812 11018 25815
rect 11052 25812 11090 25815
rect 11124 25812 11162 25815
rect 11196 25812 11234 25815
rect 11268 25812 11306 25815
rect 11340 25812 11378 25815
rect 11412 25812 11450 25815
rect 10226 25778 10260 25781
rect 10294 25781 10298 25812
rect 10362 25781 10370 25812
rect 10430 25781 10442 25812
rect 10498 25781 10514 25812
rect 10566 25781 10586 25812
rect 10634 25781 10658 25812
rect 10702 25781 10730 25812
rect 10770 25781 10802 25812
rect 10294 25778 10328 25781
rect 10362 25778 10396 25781
rect 10430 25778 10464 25781
rect 10498 25778 10532 25781
rect 10566 25778 10600 25781
rect 10634 25778 10668 25781
rect 10702 25778 10736 25781
rect 10770 25778 10804 25781
rect 10838 25778 10872 25812
rect 10908 25781 10940 25812
rect 10980 25781 11008 25812
rect 11052 25781 11076 25812
rect 11124 25781 11144 25812
rect 11196 25781 11212 25812
rect 11268 25781 11280 25812
rect 11340 25781 11348 25812
rect 11412 25781 11416 25812
rect 10906 25778 10940 25781
rect 10974 25778 11008 25781
rect 11042 25778 11076 25781
rect 11110 25778 11144 25781
rect 11178 25778 11212 25781
rect 11246 25778 11280 25781
rect 11314 25778 11348 25781
rect 11382 25778 11416 25781
rect 11484 25812 11522 25815
rect 11556 25812 11594 25815
rect 11628 25812 11666 25815
rect 11700 25812 11738 25815
rect 11772 25812 11810 25815
rect 11844 25812 11882 25815
rect 11916 25812 11954 25815
rect 11988 25812 12026 25815
rect 12060 25812 12098 25815
rect 12132 25812 12170 25815
rect 12204 25812 12242 25815
rect 12276 25812 12314 25815
rect 12348 25812 12386 25815
rect 12420 25812 12458 25815
rect 12492 25812 12530 25815
rect 12564 25812 12602 25815
rect 12636 25812 12674 25815
rect 11450 25778 11484 25781
rect 11518 25781 11522 25812
rect 11586 25781 11594 25812
rect 11654 25781 11666 25812
rect 11722 25781 11738 25812
rect 11790 25781 11810 25812
rect 11858 25781 11882 25812
rect 11926 25781 11954 25812
rect 11994 25781 12026 25812
rect 11518 25778 11552 25781
rect 11586 25778 11620 25781
rect 11654 25778 11688 25781
rect 11722 25778 11756 25781
rect 11790 25778 11824 25781
rect 11858 25778 11892 25781
rect 11926 25778 11960 25781
rect 11994 25778 12028 25781
rect 12062 25778 12096 25812
rect 12132 25781 12164 25812
rect 12204 25781 12232 25812
rect 12276 25781 12300 25812
rect 12348 25781 12368 25812
rect 12420 25781 12436 25812
rect 12492 25781 12504 25812
rect 12564 25781 12572 25812
rect 12636 25781 12640 25812
rect 12130 25778 12164 25781
rect 12198 25778 12232 25781
rect 12266 25778 12300 25781
rect 12334 25778 12368 25781
rect 12402 25778 12436 25781
rect 12470 25778 12504 25781
rect 12538 25778 12572 25781
rect 12606 25778 12640 25781
rect 12708 25812 12746 25815
rect 12780 25812 12818 25815
rect 12852 25812 12890 25815
rect 12924 25812 12962 25815
rect 12996 25812 13034 25815
rect 13068 25812 13106 25815
rect 13140 25812 13178 25815
rect 13212 25812 13250 25815
rect 13284 25812 13322 25815
rect 13356 25812 13394 25815
rect 13428 25812 13466 25815
rect 13500 25812 13538 25815
rect 13572 25812 13610 25815
rect 13644 25812 13682 25815
rect 13716 25812 13754 25815
rect 13788 25812 13826 25815
rect 13860 25812 13898 25815
rect 12674 25778 12708 25781
rect 12742 25781 12746 25812
rect 12810 25781 12818 25812
rect 12878 25781 12890 25812
rect 12946 25781 12962 25812
rect 13014 25781 13034 25812
rect 13082 25781 13106 25812
rect 13150 25781 13178 25812
rect 13218 25781 13250 25812
rect 12742 25778 12776 25781
rect 12810 25778 12844 25781
rect 12878 25778 12912 25781
rect 12946 25778 12980 25781
rect 13014 25778 13048 25781
rect 13082 25778 13116 25781
rect 13150 25778 13184 25781
rect 13218 25778 13252 25781
rect 13286 25778 13320 25812
rect 13356 25781 13388 25812
rect 13428 25781 13456 25812
rect 13500 25781 13524 25812
rect 13572 25781 13592 25812
rect 13644 25781 13660 25812
rect 13716 25781 13728 25812
rect 13788 25781 13796 25812
rect 13860 25781 13864 25812
rect 13354 25778 13388 25781
rect 13422 25778 13456 25781
rect 13490 25778 13524 25781
rect 13558 25778 13592 25781
rect 13626 25778 13660 25781
rect 13694 25778 13728 25781
rect 13762 25778 13796 25781
rect 13830 25778 13864 25781
rect 13932 25812 13970 25815
rect 14004 25812 14042 25815
rect 14076 25812 14114 25815
rect 14148 25812 14186 25815
rect 14220 25812 14258 25815
rect 14292 25812 14330 25815
rect 14364 25812 14402 25815
rect 14436 25812 14474 25815
rect 14508 25812 14546 25815
rect 14580 25812 14618 25815
rect 14652 25812 14690 25815
rect 14724 25812 14962 25815
rect 13898 25778 13932 25781
rect 13966 25781 13970 25812
rect 14034 25781 14042 25812
rect 14102 25781 14114 25812
rect 14170 25781 14186 25812
rect 14238 25781 14258 25812
rect 14306 25781 14330 25812
rect 14374 25781 14402 25812
rect 14442 25781 14474 25812
rect 13966 25778 14000 25781
rect 14034 25778 14068 25781
rect 14102 25778 14136 25781
rect 14170 25778 14204 25781
rect 14238 25778 14272 25781
rect 14306 25778 14340 25781
rect 14374 25778 14408 25781
rect 14442 25778 14476 25781
rect 14510 25778 14544 25812
rect 14580 25781 14612 25812
rect 14652 25781 14680 25812
rect 14724 25781 14748 25812
rect 14578 25778 14612 25781
rect 14646 25778 14680 25781
rect 14714 25778 14748 25781
rect 14782 25778 14816 25812
rect 14850 25778 14884 25812
rect 14918 25778 14962 25812
rect 49 25741 14962 25778
rect 49 25740 243 25741
rect 277 25740 316 25741
rect 350 25740 389 25741
rect 423 25740 462 25741
rect 496 25740 535 25741
rect 569 25740 608 25741
rect 642 25740 681 25741
rect 715 25740 754 25741
rect 788 25740 827 25741
rect 861 25740 900 25741
rect 934 25740 973 25741
rect 1007 25740 1046 25741
rect 1080 25740 1119 25741
rect 1153 25740 1192 25741
rect 1226 25740 1265 25741
rect 1299 25740 1338 25741
rect 1372 25740 1411 25741
rect 1445 25740 1484 25741
rect 49 25706 69 25740
rect 103 25706 138 25740
rect 172 25706 207 25740
rect 241 25707 243 25740
rect 310 25707 316 25740
rect 379 25707 389 25740
rect 448 25707 462 25740
rect 517 25707 535 25740
rect 586 25707 608 25740
rect 655 25707 681 25740
rect 724 25707 754 25740
rect 793 25707 827 25740
rect 241 25706 276 25707
rect 310 25706 345 25707
rect 379 25706 414 25707
rect 448 25706 483 25707
rect 517 25706 552 25707
rect 586 25706 621 25707
rect 655 25706 690 25707
rect 724 25706 759 25707
rect 793 25706 828 25707
rect 862 25706 897 25740
rect 934 25707 966 25740
rect 1007 25707 1035 25740
rect 1080 25707 1104 25740
rect 1153 25707 1173 25740
rect 1226 25707 1242 25740
rect 1299 25707 1311 25740
rect 1372 25707 1380 25740
rect 1445 25707 1449 25740
rect 931 25706 966 25707
rect 1000 25706 1035 25707
rect 1069 25706 1104 25707
rect 1138 25706 1173 25707
rect 1207 25706 1242 25707
rect 1276 25706 1311 25707
rect 1345 25706 1380 25707
rect 1414 25706 1449 25707
rect 1483 25707 1484 25740
rect 1518 25740 1557 25741
rect 1591 25740 1630 25741
rect 1664 25740 1703 25741
rect 1737 25740 1776 25741
rect 1810 25740 1849 25741
rect 1883 25740 1922 25741
rect 1956 25740 1995 25741
rect 2029 25740 2068 25741
rect 2102 25740 2141 25741
rect 2175 25740 2214 25741
rect 2248 25740 2287 25741
rect 2321 25740 2360 25741
rect 2394 25740 2433 25741
rect 2467 25740 2506 25741
rect 2540 25740 2579 25741
rect 2613 25740 2652 25741
rect 2686 25740 2725 25741
rect 1483 25706 1518 25707
rect 1552 25707 1557 25740
rect 1621 25707 1630 25740
rect 1690 25707 1703 25740
rect 1759 25707 1776 25740
rect 1828 25707 1849 25740
rect 1897 25707 1922 25740
rect 1966 25707 1995 25740
rect 2035 25707 2068 25740
rect 1552 25706 1587 25707
rect 1621 25706 1656 25707
rect 1690 25706 1725 25707
rect 1759 25706 1794 25707
rect 1828 25706 1863 25707
rect 1897 25706 1932 25707
rect 1966 25706 2001 25707
rect 2035 25706 2070 25707
rect 2104 25706 2139 25740
rect 2175 25707 2208 25740
rect 2248 25707 2277 25740
rect 2321 25707 2346 25740
rect 2394 25707 2415 25740
rect 2467 25707 2484 25740
rect 2540 25707 2553 25740
rect 2613 25707 2622 25740
rect 2686 25707 2691 25740
rect 2173 25706 2208 25707
rect 2242 25706 2277 25707
rect 2311 25706 2346 25707
rect 2380 25706 2415 25707
rect 2449 25706 2484 25707
rect 2518 25706 2553 25707
rect 2587 25706 2622 25707
rect 2656 25706 2691 25707
rect 2759 25740 2798 25741
rect 2832 25740 2871 25741
rect 2905 25740 2944 25741
rect 2978 25740 3017 25741
rect 3051 25740 3090 25741
rect 3124 25740 3163 25741
rect 3197 25740 3236 25741
rect 3270 25740 3309 25741
rect 3343 25740 3382 25741
rect 3416 25740 3455 25741
rect 3489 25740 3528 25741
rect 3562 25740 3601 25741
rect 3635 25740 3674 25741
rect 3708 25740 3746 25741
rect 3780 25740 3818 25741
rect 3852 25740 3890 25741
rect 3924 25740 3962 25741
rect 3996 25740 4034 25741
rect 4068 25740 4106 25741
rect 2759 25707 2760 25740
rect 2725 25706 2760 25707
rect 2794 25707 2798 25740
rect 2863 25707 2871 25740
rect 2932 25707 2944 25740
rect 3001 25707 3017 25740
rect 3070 25707 3090 25740
rect 3139 25707 3163 25740
rect 3208 25707 3236 25740
rect 3277 25707 3309 25740
rect 2794 25706 2829 25707
rect 2863 25706 2898 25707
rect 2932 25706 2967 25707
rect 3001 25706 3036 25707
rect 3070 25706 3105 25707
rect 3139 25706 3174 25707
rect 3208 25706 3243 25707
rect 3277 25706 3312 25707
rect 3346 25706 3381 25740
rect 3416 25707 3450 25740
rect 3489 25707 3519 25740
rect 3562 25707 3588 25740
rect 3635 25707 3657 25740
rect 3708 25707 3726 25740
rect 3780 25707 3795 25740
rect 3852 25707 3864 25740
rect 3924 25707 3933 25740
rect 3996 25707 4002 25740
rect 4068 25707 4071 25740
rect 3415 25706 3450 25707
rect 3484 25706 3519 25707
rect 3553 25706 3588 25707
rect 3622 25706 3657 25707
rect 3691 25706 3726 25707
rect 3760 25706 3795 25707
rect 3829 25706 3864 25707
rect 3898 25706 3933 25707
rect 3967 25706 4002 25707
rect 4036 25706 4071 25707
rect 4105 25707 4106 25740
rect 4140 25740 4178 25741
rect 4212 25740 4250 25741
rect 4284 25740 4322 25741
rect 4356 25740 4394 25741
rect 4428 25740 4466 25741
rect 4500 25740 4538 25741
rect 4572 25740 4610 25741
rect 4644 25740 4682 25741
rect 4716 25740 4754 25741
rect 4788 25740 4826 25741
rect 4860 25740 4898 25741
rect 4932 25740 4970 25741
rect 5004 25740 5042 25741
rect 5076 25740 5114 25741
rect 5148 25740 5186 25741
rect 5220 25740 5258 25741
rect 5292 25740 5330 25741
rect 4105 25706 4140 25707
rect 4174 25707 4178 25740
rect 4242 25707 4250 25740
rect 4310 25707 4322 25740
rect 4378 25707 4394 25740
rect 4446 25707 4466 25740
rect 4514 25707 4538 25740
rect 4582 25707 4610 25740
rect 4650 25707 4682 25740
rect 4174 25706 4208 25707
rect 4242 25706 4276 25707
rect 4310 25706 4344 25707
rect 4378 25706 4412 25707
rect 4446 25706 4480 25707
rect 4514 25706 4548 25707
rect 4582 25706 4616 25707
rect 4650 25706 4684 25707
rect 4718 25706 4752 25740
rect 4788 25707 4820 25740
rect 4860 25707 4888 25740
rect 4932 25707 4956 25740
rect 5004 25707 5024 25740
rect 5076 25707 5092 25740
rect 5148 25707 5160 25740
rect 5220 25707 5228 25740
rect 5292 25707 5296 25740
rect 4786 25706 4820 25707
rect 4854 25706 4888 25707
rect 4922 25706 4956 25707
rect 4990 25706 5024 25707
rect 5058 25706 5092 25707
rect 5126 25706 5160 25707
rect 5194 25706 5228 25707
rect 5262 25706 5296 25707
rect 5364 25740 5402 25741
rect 5436 25740 5474 25741
rect 5508 25740 5546 25741
rect 5580 25740 5618 25741
rect 5652 25740 5690 25741
rect 5724 25740 5762 25741
rect 5796 25740 5834 25741
rect 5868 25740 5906 25741
rect 5940 25740 5978 25741
rect 6012 25740 6050 25741
rect 6084 25740 6122 25741
rect 6156 25740 6194 25741
rect 6228 25740 6266 25741
rect 6300 25740 6338 25741
rect 6372 25740 6410 25741
rect 6444 25740 6482 25741
rect 6516 25740 6554 25741
rect 5330 25706 5364 25707
rect 5398 25707 5402 25740
rect 5466 25707 5474 25740
rect 5534 25707 5546 25740
rect 5602 25707 5618 25740
rect 5670 25707 5690 25740
rect 5738 25707 5762 25740
rect 5806 25707 5834 25740
rect 5874 25707 5906 25740
rect 5398 25706 5432 25707
rect 5466 25706 5500 25707
rect 5534 25706 5568 25707
rect 5602 25706 5636 25707
rect 5670 25706 5704 25707
rect 5738 25706 5772 25707
rect 5806 25706 5840 25707
rect 5874 25706 5908 25707
rect 5942 25706 5976 25740
rect 6012 25707 6044 25740
rect 6084 25707 6112 25740
rect 6156 25707 6180 25740
rect 6228 25707 6248 25740
rect 6300 25707 6316 25740
rect 6372 25707 6384 25740
rect 6444 25707 6452 25740
rect 6516 25707 6520 25740
rect 6010 25706 6044 25707
rect 6078 25706 6112 25707
rect 6146 25706 6180 25707
rect 6214 25706 6248 25707
rect 6282 25706 6316 25707
rect 6350 25706 6384 25707
rect 6418 25706 6452 25707
rect 6486 25706 6520 25707
rect 6588 25740 6626 25741
rect 6660 25740 6698 25741
rect 6732 25740 6770 25741
rect 6804 25740 6842 25741
rect 6876 25740 6914 25741
rect 6948 25740 6986 25741
rect 7020 25740 7058 25741
rect 7092 25740 7130 25741
rect 7164 25740 7202 25741
rect 7236 25740 7274 25741
rect 7308 25740 7346 25741
rect 7380 25740 7418 25741
rect 7452 25740 7490 25741
rect 7524 25740 7562 25741
rect 7596 25740 7634 25741
rect 7668 25740 7706 25741
rect 7740 25740 7778 25741
rect 6554 25706 6588 25707
rect 6622 25707 6626 25740
rect 6690 25707 6698 25740
rect 6758 25707 6770 25740
rect 6826 25707 6842 25740
rect 6894 25707 6914 25740
rect 6962 25707 6986 25740
rect 7030 25707 7058 25740
rect 7098 25707 7130 25740
rect 6622 25706 6656 25707
rect 6690 25706 6724 25707
rect 6758 25706 6792 25707
rect 6826 25706 6860 25707
rect 6894 25706 6928 25707
rect 6962 25706 6996 25707
rect 7030 25706 7064 25707
rect 7098 25706 7132 25707
rect 7166 25706 7200 25740
rect 7236 25707 7268 25740
rect 7308 25707 7336 25740
rect 7380 25707 7404 25740
rect 7452 25707 7472 25740
rect 7524 25707 7540 25740
rect 7596 25707 7608 25740
rect 7668 25707 7676 25740
rect 7740 25707 7744 25740
rect 7234 25706 7268 25707
rect 7302 25706 7336 25707
rect 7370 25706 7404 25707
rect 7438 25706 7472 25707
rect 7506 25706 7540 25707
rect 7574 25706 7608 25707
rect 7642 25706 7676 25707
rect 7710 25706 7744 25707
rect 7812 25740 7850 25741
rect 7884 25740 7922 25741
rect 7956 25740 7994 25741
rect 8028 25740 8066 25741
rect 8100 25740 8138 25741
rect 8172 25740 8210 25741
rect 8244 25740 8282 25741
rect 8316 25740 8354 25741
rect 8388 25740 8426 25741
rect 8460 25740 8498 25741
rect 8532 25740 8570 25741
rect 8604 25740 8642 25741
rect 8676 25740 8714 25741
rect 8748 25740 8786 25741
rect 8820 25740 8858 25741
rect 8892 25740 8930 25741
rect 8964 25740 9002 25741
rect 7778 25706 7812 25707
rect 7846 25707 7850 25740
rect 7914 25707 7922 25740
rect 7982 25707 7994 25740
rect 8050 25707 8066 25740
rect 8118 25707 8138 25740
rect 8186 25707 8210 25740
rect 8254 25707 8282 25740
rect 8322 25707 8354 25740
rect 7846 25706 7880 25707
rect 7914 25706 7948 25707
rect 7982 25706 8016 25707
rect 8050 25706 8084 25707
rect 8118 25706 8152 25707
rect 8186 25706 8220 25707
rect 8254 25706 8288 25707
rect 8322 25706 8356 25707
rect 8390 25706 8424 25740
rect 8460 25707 8492 25740
rect 8532 25707 8560 25740
rect 8604 25707 8628 25740
rect 8676 25707 8696 25740
rect 8748 25707 8764 25740
rect 8820 25707 8832 25740
rect 8892 25707 8900 25740
rect 8964 25707 8968 25740
rect 8458 25706 8492 25707
rect 8526 25706 8560 25707
rect 8594 25706 8628 25707
rect 8662 25706 8696 25707
rect 8730 25706 8764 25707
rect 8798 25706 8832 25707
rect 8866 25706 8900 25707
rect 8934 25706 8968 25707
rect 9036 25740 9074 25741
rect 9108 25740 9146 25741
rect 9180 25740 9218 25741
rect 9252 25740 9290 25741
rect 9324 25740 9362 25741
rect 9396 25740 9434 25741
rect 9468 25740 9506 25741
rect 9540 25740 9578 25741
rect 9612 25740 9650 25741
rect 9684 25740 9722 25741
rect 9756 25740 9794 25741
rect 9828 25740 9866 25741
rect 9900 25740 9938 25741
rect 9972 25740 10010 25741
rect 10044 25740 10082 25741
rect 10116 25740 10154 25741
rect 10188 25740 10226 25741
rect 9002 25706 9036 25707
rect 9070 25707 9074 25740
rect 9138 25707 9146 25740
rect 9206 25707 9218 25740
rect 9274 25707 9290 25740
rect 9342 25707 9362 25740
rect 9410 25707 9434 25740
rect 9478 25707 9506 25740
rect 9546 25707 9578 25740
rect 9070 25706 9104 25707
rect 9138 25706 9172 25707
rect 9206 25706 9240 25707
rect 9274 25706 9308 25707
rect 9342 25706 9376 25707
rect 9410 25706 9444 25707
rect 9478 25706 9512 25707
rect 9546 25706 9580 25707
rect 9614 25706 9648 25740
rect 9684 25707 9716 25740
rect 9756 25707 9784 25740
rect 9828 25707 9852 25740
rect 9900 25707 9920 25740
rect 9972 25707 9988 25740
rect 10044 25707 10056 25740
rect 10116 25707 10124 25740
rect 10188 25707 10192 25740
rect 9682 25706 9716 25707
rect 9750 25706 9784 25707
rect 9818 25706 9852 25707
rect 9886 25706 9920 25707
rect 9954 25706 9988 25707
rect 10022 25706 10056 25707
rect 10090 25706 10124 25707
rect 10158 25706 10192 25707
rect 10260 25740 10298 25741
rect 10332 25740 10370 25741
rect 10404 25740 10442 25741
rect 10476 25740 10514 25741
rect 10548 25740 10586 25741
rect 10620 25740 10658 25741
rect 10692 25740 10730 25741
rect 10764 25740 10802 25741
rect 10836 25740 10874 25741
rect 10908 25740 10946 25741
rect 10980 25740 11018 25741
rect 11052 25740 11090 25741
rect 11124 25740 11162 25741
rect 11196 25740 11234 25741
rect 11268 25740 11306 25741
rect 11340 25740 11378 25741
rect 11412 25740 11450 25741
rect 10226 25706 10260 25707
rect 10294 25707 10298 25740
rect 10362 25707 10370 25740
rect 10430 25707 10442 25740
rect 10498 25707 10514 25740
rect 10566 25707 10586 25740
rect 10634 25707 10658 25740
rect 10702 25707 10730 25740
rect 10770 25707 10802 25740
rect 10294 25706 10328 25707
rect 10362 25706 10396 25707
rect 10430 25706 10464 25707
rect 10498 25706 10532 25707
rect 10566 25706 10600 25707
rect 10634 25706 10668 25707
rect 10702 25706 10736 25707
rect 10770 25706 10804 25707
rect 10838 25706 10872 25740
rect 10908 25707 10940 25740
rect 10980 25707 11008 25740
rect 11052 25707 11076 25740
rect 11124 25707 11144 25740
rect 11196 25707 11212 25740
rect 11268 25707 11280 25740
rect 11340 25707 11348 25740
rect 11412 25707 11416 25740
rect 10906 25706 10940 25707
rect 10974 25706 11008 25707
rect 11042 25706 11076 25707
rect 11110 25706 11144 25707
rect 11178 25706 11212 25707
rect 11246 25706 11280 25707
rect 11314 25706 11348 25707
rect 11382 25706 11416 25707
rect 11484 25740 11522 25741
rect 11556 25740 11594 25741
rect 11628 25740 11666 25741
rect 11700 25740 11738 25741
rect 11772 25740 11810 25741
rect 11844 25740 11882 25741
rect 11916 25740 11954 25741
rect 11988 25740 12026 25741
rect 12060 25740 12098 25741
rect 12132 25740 12170 25741
rect 12204 25740 12242 25741
rect 12276 25740 12314 25741
rect 12348 25740 12386 25741
rect 12420 25740 12458 25741
rect 12492 25740 12530 25741
rect 12564 25740 12602 25741
rect 12636 25740 12674 25741
rect 11450 25706 11484 25707
rect 11518 25707 11522 25740
rect 11586 25707 11594 25740
rect 11654 25707 11666 25740
rect 11722 25707 11738 25740
rect 11790 25707 11810 25740
rect 11858 25707 11882 25740
rect 11926 25707 11954 25740
rect 11994 25707 12026 25740
rect 11518 25706 11552 25707
rect 11586 25706 11620 25707
rect 11654 25706 11688 25707
rect 11722 25706 11756 25707
rect 11790 25706 11824 25707
rect 11858 25706 11892 25707
rect 11926 25706 11960 25707
rect 11994 25706 12028 25707
rect 12062 25706 12096 25740
rect 12132 25707 12164 25740
rect 12204 25707 12232 25740
rect 12276 25707 12300 25740
rect 12348 25707 12368 25740
rect 12420 25707 12436 25740
rect 12492 25707 12504 25740
rect 12564 25707 12572 25740
rect 12636 25707 12640 25740
rect 12130 25706 12164 25707
rect 12198 25706 12232 25707
rect 12266 25706 12300 25707
rect 12334 25706 12368 25707
rect 12402 25706 12436 25707
rect 12470 25706 12504 25707
rect 12538 25706 12572 25707
rect 12606 25706 12640 25707
rect 12708 25740 12746 25741
rect 12780 25740 12818 25741
rect 12852 25740 12890 25741
rect 12924 25740 12962 25741
rect 12996 25740 13034 25741
rect 13068 25740 13106 25741
rect 13140 25740 13178 25741
rect 13212 25740 13250 25741
rect 13284 25740 13322 25741
rect 13356 25740 13394 25741
rect 13428 25740 13466 25741
rect 13500 25740 13538 25741
rect 13572 25740 13610 25741
rect 13644 25740 13682 25741
rect 13716 25740 13754 25741
rect 13788 25740 13826 25741
rect 13860 25740 13898 25741
rect 12674 25706 12708 25707
rect 12742 25707 12746 25740
rect 12810 25707 12818 25740
rect 12878 25707 12890 25740
rect 12946 25707 12962 25740
rect 13014 25707 13034 25740
rect 13082 25707 13106 25740
rect 13150 25707 13178 25740
rect 13218 25707 13250 25740
rect 12742 25706 12776 25707
rect 12810 25706 12844 25707
rect 12878 25706 12912 25707
rect 12946 25706 12980 25707
rect 13014 25706 13048 25707
rect 13082 25706 13116 25707
rect 13150 25706 13184 25707
rect 13218 25706 13252 25707
rect 13286 25706 13320 25740
rect 13356 25707 13388 25740
rect 13428 25707 13456 25740
rect 13500 25707 13524 25740
rect 13572 25707 13592 25740
rect 13644 25707 13660 25740
rect 13716 25707 13728 25740
rect 13788 25707 13796 25740
rect 13860 25707 13864 25740
rect 13354 25706 13388 25707
rect 13422 25706 13456 25707
rect 13490 25706 13524 25707
rect 13558 25706 13592 25707
rect 13626 25706 13660 25707
rect 13694 25706 13728 25707
rect 13762 25706 13796 25707
rect 13830 25706 13864 25707
rect 13932 25740 13970 25741
rect 14004 25740 14042 25741
rect 14076 25740 14114 25741
rect 14148 25740 14186 25741
rect 14220 25740 14258 25741
rect 14292 25740 14330 25741
rect 14364 25740 14402 25741
rect 14436 25740 14474 25741
rect 14508 25740 14546 25741
rect 14580 25740 14618 25741
rect 14652 25740 14690 25741
rect 14724 25740 14962 25741
rect 13898 25706 13932 25707
rect 13966 25707 13970 25740
rect 14034 25707 14042 25740
rect 14102 25707 14114 25740
rect 14170 25707 14186 25740
rect 14238 25707 14258 25740
rect 14306 25707 14330 25740
rect 14374 25707 14402 25740
rect 14442 25707 14474 25740
rect 13966 25706 14000 25707
rect 14034 25706 14068 25707
rect 14102 25706 14136 25707
rect 14170 25706 14204 25707
rect 14238 25706 14272 25707
rect 14306 25706 14340 25707
rect 14374 25706 14408 25707
rect 14442 25706 14476 25707
rect 14510 25706 14544 25740
rect 14580 25707 14612 25740
rect 14652 25707 14680 25740
rect 14724 25707 14748 25740
rect 14578 25706 14612 25707
rect 14646 25706 14680 25707
rect 14714 25706 14748 25707
rect 14782 25706 14816 25740
rect 14850 25706 14884 25740
rect 14918 25706 14962 25740
rect 49 25668 14962 25706
rect 49 25634 69 25668
rect 103 25634 138 25668
rect 172 25634 207 25668
rect 241 25667 276 25668
rect 310 25667 345 25668
rect 379 25667 414 25668
rect 448 25667 483 25668
rect 517 25667 552 25668
rect 586 25667 621 25668
rect 655 25667 690 25668
rect 724 25667 759 25668
rect 793 25667 828 25668
rect 241 25634 243 25667
rect 310 25634 316 25667
rect 379 25634 389 25667
rect 448 25634 462 25667
rect 517 25634 535 25667
rect 586 25634 608 25667
rect 655 25634 681 25667
rect 724 25634 754 25667
rect 793 25634 827 25667
rect 862 25634 897 25668
rect 931 25667 966 25668
rect 1000 25667 1035 25668
rect 1069 25667 1104 25668
rect 1138 25667 1173 25668
rect 1207 25667 1242 25668
rect 1276 25667 1311 25668
rect 1345 25667 1380 25668
rect 1414 25667 1449 25668
rect 934 25634 966 25667
rect 1007 25634 1035 25667
rect 1080 25634 1104 25667
rect 1153 25634 1173 25667
rect 1226 25634 1242 25667
rect 1299 25634 1311 25667
rect 1372 25634 1380 25667
rect 1445 25634 1449 25667
rect 1483 25667 1518 25668
rect 1483 25634 1484 25667
rect 49 25633 243 25634
rect 277 25633 316 25634
rect 350 25633 389 25634
rect 423 25633 462 25634
rect 496 25633 535 25634
rect 569 25633 608 25634
rect 642 25633 681 25634
rect 715 25633 754 25634
rect 788 25633 827 25634
rect 861 25633 900 25634
rect 934 25633 973 25634
rect 1007 25633 1046 25634
rect 1080 25633 1119 25634
rect 1153 25633 1192 25634
rect 1226 25633 1265 25634
rect 1299 25633 1338 25634
rect 1372 25633 1411 25634
rect 1445 25633 1484 25634
rect 1552 25667 1587 25668
rect 1621 25667 1656 25668
rect 1690 25667 1725 25668
rect 1759 25667 1794 25668
rect 1828 25667 1863 25668
rect 1897 25667 1932 25668
rect 1966 25667 2001 25668
rect 2035 25667 2070 25668
rect 1552 25634 1557 25667
rect 1621 25634 1630 25667
rect 1690 25634 1703 25667
rect 1759 25634 1776 25667
rect 1828 25634 1849 25667
rect 1897 25634 1922 25667
rect 1966 25634 1995 25667
rect 2035 25634 2068 25667
rect 2104 25634 2139 25668
rect 2173 25667 2208 25668
rect 2242 25667 2277 25668
rect 2311 25667 2346 25668
rect 2380 25667 2415 25668
rect 2449 25667 2484 25668
rect 2518 25667 2553 25668
rect 2587 25667 2622 25668
rect 2656 25667 2691 25668
rect 2175 25634 2208 25667
rect 2248 25634 2277 25667
rect 2321 25634 2346 25667
rect 2394 25634 2415 25667
rect 2467 25634 2484 25667
rect 2540 25634 2553 25667
rect 2613 25634 2622 25667
rect 2686 25634 2691 25667
rect 2725 25667 2760 25668
rect 1518 25633 1557 25634
rect 1591 25633 1630 25634
rect 1664 25633 1703 25634
rect 1737 25633 1776 25634
rect 1810 25633 1849 25634
rect 1883 25633 1922 25634
rect 1956 25633 1995 25634
rect 2029 25633 2068 25634
rect 2102 25633 2141 25634
rect 2175 25633 2214 25634
rect 2248 25633 2287 25634
rect 2321 25633 2360 25634
rect 2394 25633 2433 25634
rect 2467 25633 2506 25634
rect 2540 25633 2579 25634
rect 2613 25633 2652 25634
rect 2686 25633 2725 25634
rect 2759 25634 2760 25667
rect 2794 25667 2829 25668
rect 2863 25667 2898 25668
rect 2932 25667 2967 25668
rect 3001 25667 3036 25668
rect 3070 25667 3105 25668
rect 3139 25667 3174 25668
rect 3208 25667 3243 25668
rect 3277 25667 3312 25668
rect 2794 25634 2798 25667
rect 2863 25634 2871 25667
rect 2932 25634 2944 25667
rect 3001 25634 3017 25667
rect 3070 25634 3090 25667
rect 3139 25634 3163 25667
rect 3208 25634 3236 25667
rect 3277 25634 3309 25667
rect 3346 25634 3381 25668
rect 3415 25667 3450 25668
rect 3484 25667 3519 25668
rect 3553 25667 3588 25668
rect 3622 25667 3657 25668
rect 3691 25667 3726 25668
rect 3760 25667 3795 25668
rect 3829 25667 3864 25668
rect 3898 25667 3933 25668
rect 3967 25667 4002 25668
rect 4036 25667 4071 25668
rect 3416 25634 3450 25667
rect 3489 25634 3519 25667
rect 3562 25634 3588 25667
rect 3635 25634 3657 25667
rect 3708 25634 3726 25667
rect 3780 25634 3795 25667
rect 3852 25634 3864 25667
rect 3924 25634 3933 25667
rect 3996 25634 4002 25667
rect 4068 25634 4071 25667
rect 4105 25667 4140 25668
rect 4105 25634 4106 25667
rect 2759 25633 2798 25634
rect 2832 25633 2871 25634
rect 2905 25633 2944 25634
rect 2978 25633 3017 25634
rect 3051 25633 3090 25634
rect 3124 25633 3163 25634
rect 3197 25633 3236 25634
rect 3270 25633 3309 25634
rect 3343 25633 3382 25634
rect 3416 25633 3455 25634
rect 3489 25633 3528 25634
rect 3562 25633 3601 25634
rect 3635 25633 3674 25634
rect 3708 25633 3746 25634
rect 3780 25633 3818 25634
rect 3852 25633 3890 25634
rect 3924 25633 3962 25634
rect 3996 25633 4034 25634
rect 4068 25633 4106 25634
rect 4174 25667 4208 25668
rect 4242 25667 4276 25668
rect 4310 25667 4344 25668
rect 4378 25667 4412 25668
rect 4446 25667 4480 25668
rect 4514 25667 4548 25668
rect 4582 25667 4616 25668
rect 4650 25667 4684 25668
rect 4174 25634 4178 25667
rect 4242 25634 4250 25667
rect 4310 25634 4322 25667
rect 4378 25634 4394 25667
rect 4446 25634 4466 25667
rect 4514 25634 4538 25667
rect 4582 25634 4610 25667
rect 4650 25634 4682 25667
rect 4718 25634 4752 25668
rect 4786 25667 4820 25668
rect 4854 25667 4888 25668
rect 4922 25667 4956 25668
rect 4990 25667 5024 25668
rect 5058 25667 5092 25668
rect 5126 25667 5160 25668
rect 5194 25667 5228 25668
rect 5262 25667 5296 25668
rect 4788 25634 4820 25667
rect 4860 25634 4888 25667
rect 4932 25634 4956 25667
rect 5004 25634 5024 25667
rect 5076 25634 5092 25667
rect 5148 25634 5160 25667
rect 5220 25634 5228 25667
rect 5292 25634 5296 25667
rect 5330 25667 5364 25668
rect 4140 25633 4178 25634
rect 4212 25633 4250 25634
rect 4284 25633 4322 25634
rect 4356 25633 4394 25634
rect 4428 25633 4466 25634
rect 4500 25633 4538 25634
rect 4572 25633 4610 25634
rect 4644 25633 4682 25634
rect 4716 25633 4754 25634
rect 4788 25633 4826 25634
rect 4860 25633 4898 25634
rect 4932 25633 4970 25634
rect 5004 25633 5042 25634
rect 5076 25633 5114 25634
rect 5148 25633 5186 25634
rect 5220 25633 5258 25634
rect 5292 25633 5330 25634
rect 5398 25667 5432 25668
rect 5466 25667 5500 25668
rect 5534 25667 5568 25668
rect 5602 25667 5636 25668
rect 5670 25667 5704 25668
rect 5738 25667 5772 25668
rect 5806 25667 5840 25668
rect 5874 25667 5908 25668
rect 5398 25634 5402 25667
rect 5466 25634 5474 25667
rect 5534 25634 5546 25667
rect 5602 25634 5618 25667
rect 5670 25634 5690 25667
rect 5738 25634 5762 25667
rect 5806 25634 5834 25667
rect 5874 25634 5906 25667
rect 5942 25634 5976 25668
rect 6010 25667 6044 25668
rect 6078 25667 6112 25668
rect 6146 25667 6180 25668
rect 6214 25667 6248 25668
rect 6282 25667 6316 25668
rect 6350 25667 6384 25668
rect 6418 25667 6452 25668
rect 6486 25667 6520 25668
rect 6012 25634 6044 25667
rect 6084 25634 6112 25667
rect 6156 25634 6180 25667
rect 6228 25634 6248 25667
rect 6300 25634 6316 25667
rect 6372 25634 6384 25667
rect 6444 25634 6452 25667
rect 6516 25634 6520 25667
rect 6554 25667 6588 25668
rect 5364 25633 5402 25634
rect 5436 25633 5474 25634
rect 5508 25633 5546 25634
rect 5580 25633 5618 25634
rect 5652 25633 5690 25634
rect 5724 25633 5762 25634
rect 5796 25633 5834 25634
rect 5868 25633 5906 25634
rect 5940 25633 5978 25634
rect 6012 25633 6050 25634
rect 6084 25633 6122 25634
rect 6156 25633 6194 25634
rect 6228 25633 6266 25634
rect 6300 25633 6338 25634
rect 6372 25633 6410 25634
rect 6444 25633 6482 25634
rect 6516 25633 6554 25634
rect 6622 25667 6656 25668
rect 6690 25667 6724 25668
rect 6758 25667 6792 25668
rect 6826 25667 6860 25668
rect 6894 25667 6928 25668
rect 6962 25667 6996 25668
rect 7030 25667 7064 25668
rect 7098 25667 7132 25668
rect 6622 25634 6626 25667
rect 6690 25634 6698 25667
rect 6758 25634 6770 25667
rect 6826 25634 6842 25667
rect 6894 25634 6914 25667
rect 6962 25634 6986 25667
rect 7030 25634 7058 25667
rect 7098 25634 7130 25667
rect 7166 25634 7200 25668
rect 7234 25667 7268 25668
rect 7302 25667 7336 25668
rect 7370 25667 7404 25668
rect 7438 25667 7472 25668
rect 7506 25667 7540 25668
rect 7574 25667 7608 25668
rect 7642 25667 7676 25668
rect 7710 25667 7744 25668
rect 7236 25634 7268 25667
rect 7308 25634 7336 25667
rect 7380 25634 7404 25667
rect 7452 25634 7472 25667
rect 7524 25634 7540 25667
rect 7596 25634 7608 25667
rect 7668 25634 7676 25667
rect 7740 25634 7744 25667
rect 7778 25667 7812 25668
rect 6588 25633 6626 25634
rect 6660 25633 6698 25634
rect 6732 25633 6770 25634
rect 6804 25633 6842 25634
rect 6876 25633 6914 25634
rect 6948 25633 6986 25634
rect 7020 25633 7058 25634
rect 7092 25633 7130 25634
rect 7164 25633 7202 25634
rect 7236 25633 7274 25634
rect 7308 25633 7346 25634
rect 7380 25633 7418 25634
rect 7452 25633 7490 25634
rect 7524 25633 7562 25634
rect 7596 25633 7634 25634
rect 7668 25633 7706 25634
rect 7740 25633 7778 25634
rect 7846 25667 7880 25668
rect 7914 25667 7948 25668
rect 7982 25667 8016 25668
rect 8050 25667 8084 25668
rect 8118 25667 8152 25668
rect 8186 25667 8220 25668
rect 8254 25667 8288 25668
rect 8322 25667 8356 25668
rect 7846 25634 7850 25667
rect 7914 25634 7922 25667
rect 7982 25634 7994 25667
rect 8050 25634 8066 25667
rect 8118 25634 8138 25667
rect 8186 25634 8210 25667
rect 8254 25634 8282 25667
rect 8322 25634 8354 25667
rect 8390 25634 8424 25668
rect 8458 25667 8492 25668
rect 8526 25667 8560 25668
rect 8594 25667 8628 25668
rect 8662 25667 8696 25668
rect 8730 25667 8764 25668
rect 8798 25667 8832 25668
rect 8866 25667 8900 25668
rect 8934 25667 8968 25668
rect 8460 25634 8492 25667
rect 8532 25634 8560 25667
rect 8604 25634 8628 25667
rect 8676 25634 8696 25667
rect 8748 25634 8764 25667
rect 8820 25634 8832 25667
rect 8892 25634 8900 25667
rect 8964 25634 8968 25667
rect 9002 25667 9036 25668
rect 7812 25633 7850 25634
rect 7884 25633 7922 25634
rect 7956 25633 7994 25634
rect 8028 25633 8066 25634
rect 8100 25633 8138 25634
rect 8172 25633 8210 25634
rect 8244 25633 8282 25634
rect 8316 25633 8354 25634
rect 8388 25633 8426 25634
rect 8460 25633 8498 25634
rect 8532 25633 8570 25634
rect 8604 25633 8642 25634
rect 8676 25633 8714 25634
rect 8748 25633 8786 25634
rect 8820 25633 8858 25634
rect 8892 25633 8930 25634
rect 8964 25633 9002 25634
rect 9070 25667 9104 25668
rect 9138 25667 9172 25668
rect 9206 25667 9240 25668
rect 9274 25667 9308 25668
rect 9342 25667 9376 25668
rect 9410 25667 9444 25668
rect 9478 25667 9512 25668
rect 9546 25667 9580 25668
rect 9070 25634 9074 25667
rect 9138 25634 9146 25667
rect 9206 25634 9218 25667
rect 9274 25634 9290 25667
rect 9342 25634 9362 25667
rect 9410 25634 9434 25667
rect 9478 25634 9506 25667
rect 9546 25634 9578 25667
rect 9614 25634 9648 25668
rect 9682 25667 9716 25668
rect 9750 25667 9784 25668
rect 9818 25667 9852 25668
rect 9886 25667 9920 25668
rect 9954 25667 9988 25668
rect 10022 25667 10056 25668
rect 10090 25667 10124 25668
rect 10158 25667 10192 25668
rect 9684 25634 9716 25667
rect 9756 25634 9784 25667
rect 9828 25634 9852 25667
rect 9900 25634 9920 25667
rect 9972 25634 9988 25667
rect 10044 25634 10056 25667
rect 10116 25634 10124 25667
rect 10188 25634 10192 25667
rect 10226 25667 10260 25668
rect 9036 25633 9074 25634
rect 9108 25633 9146 25634
rect 9180 25633 9218 25634
rect 9252 25633 9290 25634
rect 9324 25633 9362 25634
rect 9396 25633 9434 25634
rect 9468 25633 9506 25634
rect 9540 25633 9578 25634
rect 9612 25633 9650 25634
rect 9684 25633 9722 25634
rect 9756 25633 9794 25634
rect 9828 25633 9866 25634
rect 9900 25633 9938 25634
rect 9972 25633 10010 25634
rect 10044 25633 10082 25634
rect 10116 25633 10154 25634
rect 10188 25633 10226 25634
rect 10294 25667 10328 25668
rect 10362 25667 10396 25668
rect 10430 25667 10464 25668
rect 10498 25667 10532 25668
rect 10566 25667 10600 25668
rect 10634 25667 10668 25668
rect 10702 25667 10736 25668
rect 10770 25667 10804 25668
rect 10294 25634 10298 25667
rect 10362 25634 10370 25667
rect 10430 25634 10442 25667
rect 10498 25634 10514 25667
rect 10566 25634 10586 25667
rect 10634 25634 10658 25667
rect 10702 25634 10730 25667
rect 10770 25634 10802 25667
rect 10838 25634 10872 25668
rect 10906 25667 10940 25668
rect 10974 25667 11008 25668
rect 11042 25667 11076 25668
rect 11110 25667 11144 25668
rect 11178 25667 11212 25668
rect 11246 25667 11280 25668
rect 11314 25667 11348 25668
rect 11382 25667 11416 25668
rect 10908 25634 10940 25667
rect 10980 25634 11008 25667
rect 11052 25634 11076 25667
rect 11124 25634 11144 25667
rect 11196 25634 11212 25667
rect 11268 25634 11280 25667
rect 11340 25634 11348 25667
rect 11412 25634 11416 25667
rect 11450 25667 11484 25668
rect 10260 25633 10298 25634
rect 10332 25633 10370 25634
rect 10404 25633 10442 25634
rect 10476 25633 10514 25634
rect 10548 25633 10586 25634
rect 10620 25633 10658 25634
rect 10692 25633 10730 25634
rect 10764 25633 10802 25634
rect 10836 25633 10874 25634
rect 10908 25633 10946 25634
rect 10980 25633 11018 25634
rect 11052 25633 11090 25634
rect 11124 25633 11162 25634
rect 11196 25633 11234 25634
rect 11268 25633 11306 25634
rect 11340 25633 11378 25634
rect 11412 25633 11450 25634
rect 11518 25667 11552 25668
rect 11586 25667 11620 25668
rect 11654 25667 11688 25668
rect 11722 25667 11756 25668
rect 11790 25667 11824 25668
rect 11858 25667 11892 25668
rect 11926 25667 11960 25668
rect 11994 25667 12028 25668
rect 11518 25634 11522 25667
rect 11586 25634 11594 25667
rect 11654 25634 11666 25667
rect 11722 25634 11738 25667
rect 11790 25634 11810 25667
rect 11858 25634 11882 25667
rect 11926 25634 11954 25667
rect 11994 25634 12026 25667
rect 12062 25634 12096 25668
rect 12130 25667 12164 25668
rect 12198 25667 12232 25668
rect 12266 25667 12300 25668
rect 12334 25667 12368 25668
rect 12402 25667 12436 25668
rect 12470 25667 12504 25668
rect 12538 25667 12572 25668
rect 12606 25667 12640 25668
rect 12132 25634 12164 25667
rect 12204 25634 12232 25667
rect 12276 25634 12300 25667
rect 12348 25634 12368 25667
rect 12420 25634 12436 25667
rect 12492 25634 12504 25667
rect 12564 25634 12572 25667
rect 12636 25634 12640 25667
rect 12674 25667 12708 25668
rect 11484 25633 11522 25634
rect 11556 25633 11594 25634
rect 11628 25633 11666 25634
rect 11700 25633 11738 25634
rect 11772 25633 11810 25634
rect 11844 25633 11882 25634
rect 11916 25633 11954 25634
rect 11988 25633 12026 25634
rect 12060 25633 12098 25634
rect 12132 25633 12170 25634
rect 12204 25633 12242 25634
rect 12276 25633 12314 25634
rect 12348 25633 12386 25634
rect 12420 25633 12458 25634
rect 12492 25633 12530 25634
rect 12564 25633 12602 25634
rect 12636 25633 12674 25634
rect 12742 25667 12776 25668
rect 12810 25667 12844 25668
rect 12878 25667 12912 25668
rect 12946 25667 12980 25668
rect 13014 25667 13048 25668
rect 13082 25667 13116 25668
rect 13150 25667 13184 25668
rect 13218 25667 13252 25668
rect 12742 25634 12746 25667
rect 12810 25634 12818 25667
rect 12878 25634 12890 25667
rect 12946 25634 12962 25667
rect 13014 25634 13034 25667
rect 13082 25634 13106 25667
rect 13150 25634 13178 25667
rect 13218 25634 13250 25667
rect 13286 25634 13320 25668
rect 13354 25667 13388 25668
rect 13422 25667 13456 25668
rect 13490 25667 13524 25668
rect 13558 25667 13592 25668
rect 13626 25667 13660 25668
rect 13694 25667 13728 25668
rect 13762 25667 13796 25668
rect 13830 25667 13864 25668
rect 13356 25634 13388 25667
rect 13428 25634 13456 25667
rect 13500 25634 13524 25667
rect 13572 25634 13592 25667
rect 13644 25634 13660 25667
rect 13716 25634 13728 25667
rect 13788 25634 13796 25667
rect 13860 25634 13864 25667
rect 13898 25667 13932 25668
rect 12708 25633 12746 25634
rect 12780 25633 12818 25634
rect 12852 25633 12890 25634
rect 12924 25633 12962 25634
rect 12996 25633 13034 25634
rect 13068 25633 13106 25634
rect 13140 25633 13178 25634
rect 13212 25633 13250 25634
rect 13284 25633 13322 25634
rect 13356 25633 13394 25634
rect 13428 25633 13466 25634
rect 13500 25633 13538 25634
rect 13572 25633 13610 25634
rect 13644 25633 13682 25634
rect 13716 25633 13754 25634
rect 13788 25633 13826 25634
rect 13860 25633 13898 25634
rect 13966 25667 14000 25668
rect 14034 25667 14068 25668
rect 14102 25667 14136 25668
rect 14170 25667 14204 25668
rect 14238 25667 14272 25668
rect 14306 25667 14340 25668
rect 14374 25667 14408 25668
rect 14442 25667 14476 25668
rect 13966 25634 13970 25667
rect 14034 25634 14042 25667
rect 14102 25634 14114 25667
rect 14170 25634 14186 25667
rect 14238 25634 14258 25667
rect 14306 25634 14330 25667
rect 14374 25634 14402 25667
rect 14442 25634 14474 25667
rect 14510 25634 14544 25668
rect 14578 25667 14612 25668
rect 14646 25667 14680 25668
rect 14714 25667 14748 25668
rect 14580 25634 14612 25667
rect 14652 25634 14680 25667
rect 14724 25634 14748 25667
rect 14782 25634 14816 25668
rect 14850 25634 14884 25668
rect 14918 25634 14962 25668
rect 13932 25633 13970 25634
rect 14004 25633 14042 25634
rect 14076 25633 14114 25634
rect 14148 25633 14186 25634
rect 14220 25633 14258 25634
rect 14292 25633 14330 25634
rect 14364 25633 14402 25634
rect 14436 25633 14474 25634
rect 14508 25633 14546 25634
rect 14580 25633 14618 25634
rect 14652 25633 14690 25634
rect 14724 25633 14962 25634
rect 49 25599 14962 25633
rect -41 25444 8304 25445
rect -41 25410 77 25444
rect 111 25410 146 25444
rect 180 25410 215 25444
rect 249 25410 284 25444
rect 318 25410 353 25444
rect 387 25410 422 25444
rect 456 25410 491 25444
rect 525 25410 560 25444
rect 594 25410 629 25444
rect 663 25410 698 25444
rect 732 25410 766 25444
rect 800 25410 834 25444
rect 868 25410 902 25444
rect 936 25410 970 25444
rect 1004 25410 1038 25444
rect 1072 25410 1106 25444
rect 1140 25410 1174 25444
rect 1208 25410 1242 25444
rect 1276 25410 1310 25444
rect 1344 25410 1378 25444
rect 1412 25410 1446 25444
rect 1480 25410 1514 25444
rect 1548 25410 1582 25444
rect 1616 25410 1650 25444
rect 1684 25410 1718 25444
rect 1752 25410 1786 25444
rect 1820 25410 1854 25444
rect 1888 25410 1922 25444
rect 1956 25410 1990 25444
rect 2024 25410 2058 25444
rect 2092 25410 2126 25444
rect 2160 25410 2194 25444
rect 2228 25410 2262 25444
rect 2296 25410 2330 25444
rect 2364 25410 2398 25444
rect 2432 25410 2466 25444
rect 2500 25410 2534 25444
rect 2568 25410 2602 25444
rect 2636 25410 2670 25444
rect 2704 25410 2738 25444
rect 2772 25410 2806 25444
rect 2840 25410 2874 25444
rect 2908 25410 2942 25444
rect 2976 25410 3010 25444
rect 3044 25410 3078 25444
rect 3112 25410 3146 25444
rect 3180 25410 3214 25444
rect 3248 25410 3282 25444
rect 3316 25410 3350 25444
rect 3384 25410 3418 25444
rect 3452 25410 3486 25444
rect 3520 25410 3554 25444
rect 3588 25410 3622 25444
rect 3656 25410 3690 25444
rect 3724 25410 3758 25444
rect 3792 25410 3826 25444
rect 3860 25410 3894 25444
rect 3928 25410 3962 25444
rect 3996 25410 4030 25444
rect 4064 25410 4098 25444
rect 4132 25410 4166 25444
rect 4200 25410 4234 25444
rect 4268 25410 4302 25444
rect 4336 25410 4370 25444
rect 4404 25410 4438 25444
rect 4472 25410 4506 25444
rect 4540 25410 4574 25444
rect 4608 25410 4642 25444
rect 4676 25410 4710 25444
rect 4744 25410 4778 25444
rect 4812 25410 4846 25444
rect 4880 25410 4914 25444
rect 4948 25410 4982 25444
rect 5016 25410 5050 25444
rect 5084 25410 5118 25444
rect 5152 25410 5186 25444
rect 5220 25410 5254 25444
rect 5288 25410 5322 25444
rect 5356 25410 5390 25444
rect 5424 25410 5458 25444
rect 5492 25410 5526 25444
rect 5560 25410 5594 25444
rect 5628 25410 5662 25444
rect 5696 25410 5730 25444
rect 5764 25410 5798 25444
rect 5832 25410 5866 25444
rect 5900 25410 5934 25444
rect 5968 25410 6002 25444
rect 6036 25410 6070 25444
rect 6104 25410 6138 25444
rect 6172 25410 6206 25444
rect 6240 25410 6274 25444
rect 6308 25410 6342 25444
rect 6376 25410 6410 25444
rect 6444 25410 6478 25444
rect 6512 25410 6546 25444
rect 6580 25410 6614 25444
rect 6648 25410 6682 25444
rect 6716 25410 6750 25444
rect 6784 25410 6818 25444
rect 6852 25410 6886 25444
rect 6920 25410 6954 25444
rect 6988 25410 7022 25444
rect 7056 25410 7090 25444
rect 7124 25410 7158 25444
rect 7192 25410 7226 25444
rect 7260 25410 7294 25444
rect 7328 25410 7362 25444
rect 7396 25410 7430 25444
rect 7464 25410 7498 25444
rect 7532 25410 7566 25444
rect 7600 25410 7634 25444
rect 7668 25410 7702 25444
rect 7736 25410 7770 25444
rect 7804 25410 7838 25444
rect 7872 25410 7906 25444
rect 7940 25410 7974 25444
rect 8008 25410 8042 25444
rect 8076 25410 8110 25444
rect 8144 25410 8178 25444
rect 8212 25410 8246 25444
rect 8280 25410 8304 25444
rect -41 25358 8304 25410
rect -41 25324 77 25358
rect 111 25324 146 25358
rect 180 25324 215 25358
rect 249 25324 284 25358
rect 318 25324 353 25358
rect 387 25324 422 25358
rect 456 25324 491 25358
rect 525 25324 560 25358
rect 594 25324 629 25358
rect 663 25324 698 25358
rect 732 25324 766 25358
rect 800 25324 834 25358
rect 868 25324 902 25358
rect 936 25324 970 25358
rect 1004 25324 1038 25358
rect 1072 25324 1106 25358
rect 1140 25324 1174 25358
rect 1208 25324 1242 25358
rect 1276 25324 1310 25358
rect 1344 25324 1378 25358
rect 1412 25324 1446 25358
rect 1480 25324 1514 25358
rect 1548 25324 1582 25358
rect 1616 25324 1650 25358
rect 1684 25324 1718 25358
rect 1752 25324 1786 25358
rect 1820 25324 1854 25358
rect 1888 25324 1922 25358
rect 1956 25324 1990 25358
rect 2024 25324 2058 25358
rect 2092 25324 2126 25358
rect 2160 25324 2194 25358
rect 2228 25324 2262 25358
rect 2296 25324 2330 25358
rect 2364 25324 2398 25358
rect 2432 25324 2466 25358
rect 2500 25324 2534 25358
rect 2568 25324 2602 25358
rect 2636 25324 2670 25358
rect 2704 25324 2738 25358
rect 2772 25324 2806 25358
rect 2840 25324 2874 25358
rect 2908 25324 2942 25358
rect 2976 25324 3010 25358
rect 3044 25324 3078 25358
rect 3112 25324 3146 25358
rect 3180 25324 3214 25358
rect 3248 25324 3282 25358
rect 3316 25324 3350 25358
rect 3384 25324 3418 25358
rect 3452 25324 3486 25358
rect 3520 25324 3554 25358
rect 3588 25324 3622 25358
rect 3656 25324 3690 25358
rect 3724 25324 3758 25358
rect 3792 25324 3826 25358
rect 3860 25324 3894 25358
rect 3928 25324 3962 25358
rect 3996 25324 4030 25358
rect 4064 25324 4098 25358
rect 4132 25324 4166 25358
rect 4200 25324 4234 25358
rect 4268 25324 4302 25358
rect 4336 25324 4370 25358
rect 4404 25324 4438 25358
rect 4472 25324 4506 25358
rect 4540 25324 4574 25358
rect 4608 25324 4642 25358
rect 4676 25324 4710 25358
rect 4744 25324 4778 25358
rect 4812 25324 4846 25358
rect 4880 25324 4914 25358
rect 4948 25324 4982 25358
rect 5016 25324 5050 25358
rect 5084 25324 5118 25358
rect 5152 25324 5186 25358
rect 5220 25324 5254 25358
rect 5288 25324 5322 25358
rect 5356 25324 5390 25358
rect 5424 25324 5458 25358
rect 5492 25324 5526 25358
rect 5560 25324 5594 25358
rect 5628 25324 5662 25358
rect 5696 25324 5730 25358
rect 5764 25324 5798 25358
rect 5832 25324 5866 25358
rect 5900 25324 5934 25358
rect 5968 25324 6002 25358
rect 6036 25324 6070 25358
rect 6104 25324 6138 25358
rect 6172 25324 6206 25358
rect 6240 25324 6274 25358
rect 6308 25324 6342 25358
rect 6376 25324 6410 25358
rect 6444 25324 6478 25358
rect 6512 25324 6546 25358
rect 6580 25324 6614 25358
rect 6648 25324 6682 25358
rect 6716 25324 6750 25358
rect 6784 25324 6818 25358
rect 6852 25324 6886 25358
rect 6920 25324 6954 25358
rect 6988 25324 7022 25358
rect 7056 25324 7090 25358
rect 7124 25324 7158 25358
rect 7192 25324 7226 25358
rect 7260 25324 7294 25358
rect 7328 25324 7362 25358
rect 7396 25324 7430 25358
rect 7464 25324 7498 25358
rect 7532 25324 7566 25358
rect 7600 25324 7634 25358
rect 7668 25324 7702 25358
rect 7736 25324 7770 25358
rect 7804 25324 7838 25358
rect 7872 25324 7906 25358
rect 7940 25324 7974 25358
rect 8008 25324 8042 25358
rect 8076 25324 8110 25358
rect 8144 25324 8178 25358
rect 8212 25324 8246 25358
rect 8280 25324 8304 25358
rect -41 25272 8304 25324
rect -41 25238 77 25272
rect 111 25238 146 25272
rect 180 25238 215 25272
rect 249 25238 284 25272
rect 318 25238 353 25272
rect 387 25238 422 25272
rect 456 25238 491 25272
rect 525 25238 560 25272
rect 594 25238 629 25272
rect 663 25238 698 25272
rect 732 25238 766 25272
rect 800 25238 834 25272
rect 868 25238 902 25272
rect 936 25238 970 25272
rect 1004 25238 1038 25272
rect 1072 25238 1106 25272
rect 1140 25238 1174 25272
rect 1208 25238 1242 25272
rect 1276 25238 1310 25272
rect 1344 25238 1378 25272
rect 1412 25238 1446 25272
rect 1480 25238 1514 25272
rect 1548 25238 1582 25272
rect 1616 25238 1650 25272
rect 1684 25238 1718 25272
rect 1752 25238 1786 25272
rect 1820 25238 1854 25272
rect 1888 25238 1922 25272
rect 1956 25238 1990 25272
rect 2024 25238 2058 25272
rect 2092 25238 2126 25272
rect 2160 25238 2194 25272
rect 2228 25238 2262 25272
rect 2296 25238 2330 25272
rect 2364 25238 2398 25272
rect 2432 25238 2466 25272
rect 2500 25238 2534 25272
rect 2568 25238 2602 25272
rect 2636 25238 2670 25272
rect 2704 25238 2738 25272
rect 2772 25238 2806 25272
rect 2840 25238 2874 25272
rect 2908 25238 2942 25272
rect 2976 25238 3010 25272
rect 3044 25238 3078 25272
rect 3112 25238 3146 25272
rect 3180 25238 3214 25272
rect 3248 25238 3282 25272
rect 3316 25238 3350 25272
rect 3384 25238 3418 25272
rect 3452 25238 3486 25272
rect 3520 25238 3554 25272
rect 3588 25238 3622 25272
rect 3656 25238 3690 25272
rect 3724 25238 3758 25272
rect 3792 25238 3826 25272
rect 3860 25238 3894 25272
rect 3928 25238 3962 25272
rect 3996 25238 4030 25272
rect 4064 25238 4098 25272
rect 4132 25238 4166 25272
rect 4200 25238 4234 25272
rect 4268 25238 4302 25272
rect 4336 25238 4370 25272
rect 4404 25238 4438 25272
rect 4472 25238 4506 25272
rect 4540 25238 4574 25272
rect 4608 25238 4642 25272
rect 4676 25238 4710 25272
rect 4744 25238 4778 25272
rect 4812 25238 4846 25272
rect 4880 25238 4914 25272
rect 4948 25238 4982 25272
rect 5016 25238 5050 25272
rect 5084 25238 5118 25272
rect 5152 25238 5186 25272
rect 5220 25238 5254 25272
rect 5288 25238 5322 25272
rect 5356 25238 5390 25272
rect 5424 25238 5458 25272
rect 5492 25238 5526 25272
rect 5560 25238 5594 25272
rect 5628 25238 5662 25272
rect 5696 25238 5730 25272
rect 5764 25238 5798 25272
rect 5832 25238 5866 25272
rect 5900 25238 5934 25272
rect 5968 25238 6002 25272
rect 6036 25238 6070 25272
rect 6104 25238 6138 25272
rect 6172 25238 6206 25272
rect 6240 25238 6274 25272
rect 6308 25238 6342 25272
rect 6376 25238 6410 25272
rect 6444 25238 6478 25272
rect 6512 25238 6546 25272
rect 6580 25238 6614 25272
rect 6648 25238 6682 25272
rect 6716 25238 6750 25272
rect 6784 25238 6818 25272
rect 6852 25238 6886 25272
rect 6920 25238 6954 25272
rect 6988 25238 7022 25272
rect 7056 25238 7090 25272
rect 7124 25238 7158 25272
rect 7192 25238 7226 25272
rect 7260 25238 7294 25272
rect 7328 25238 7362 25272
rect 7396 25238 7430 25272
rect 7464 25238 7498 25272
rect 7532 25238 7566 25272
rect 7600 25238 7634 25272
rect 7668 25238 7702 25272
rect 7736 25238 7770 25272
rect 7804 25238 7838 25272
rect 7872 25238 7906 25272
rect 7940 25238 7974 25272
rect 8008 25238 8042 25272
rect 8076 25238 8110 25272
rect 8144 25238 8178 25272
rect 8212 25238 8246 25272
rect 8280 25238 8304 25272
rect -41 25180 8304 25238
rect 12408 25444 14882 25445
rect 12408 25410 12432 25444
rect 12466 25410 12501 25444
rect 12535 25410 12570 25444
rect 12604 25410 12639 25444
rect 12673 25410 12708 25444
rect 12742 25410 12777 25444
rect 12811 25410 12846 25444
rect 12880 25410 12915 25444
rect 12949 25410 12984 25444
rect 13018 25410 13053 25444
rect 13087 25410 13122 25444
rect 13156 25410 13191 25444
rect 13225 25410 13260 25444
rect 13294 25410 13328 25444
rect 13362 25410 13396 25444
rect 13430 25410 13464 25444
rect 13498 25410 13532 25444
rect 13566 25410 13600 25444
rect 13634 25410 13668 25444
rect 13702 25410 13736 25444
rect 13770 25410 13804 25444
rect 13838 25410 13872 25444
rect 13906 25410 13940 25444
rect 13974 25410 14008 25444
rect 14042 25410 14076 25444
rect 14110 25410 14144 25444
rect 14178 25410 14212 25444
rect 14246 25410 14280 25444
rect 14314 25410 14348 25444
rect 14382 25410 14416 25444
rect 14450 25410 14484 25444
rect 14518 25410 14552 25444
rect 14586 25410 14620 25444
rect 14654 25410 14688 25444
rect 14722 25410 14756 25444
rect 14790 25410 14824 25444
rect 14858 25410 14983 25444
rect 12408 25358 14983 25410
rect 12408 25324 12432 25358
rect 12466 25324 12501 25358
rect 12535 25324 12570 25358
rect 12604 25324 12639 25358
rect 12673 25324 12708 25358
rect 12742 25324 12777 25358
rect 12811 25324 12846 25358
rect 12880 25324 12915 25358
rect 12949 25324 12984 25358
rect 13018 25324 13053 25358
rect 13087 25324 13122 25358
rect 13156 25324 13191 25358
rect 13225 25324 13260 25358
rect 13294 25324 13328 25358
rect 13362 25324 13396 25358
rect 13430 25324 13464 25358
rect 13498 25324 13532 25358
rect 13566 25324 13600 25358
rect 13634 25324 13668 25358
rect 13702 25324 13736 25358
rect 13770 25324 13804 25358
rect 13838 25324 13872 25358
rect 13906 25324 13940 25358
rect 13974 25324 14008 25358
rect 14042 25324 14076 25358
rect 14110 25324 14144 25358
rect 14178 25324 14212 25358
rect 14246 25324 14280 25358
rect 14314 25324 14348 25358
rect 14382 25324 14416 25358
rect 14450 25324 14484 25358
rect 14518 25324 14552 25358
rect 14586 25324 14620 25358
rect 14654 25324 14688 25358
rect 14722 25324 14756 25358
rect 14790 25324 14824 25358
rect 14858 25324 14983 25358
rect 12408 25272 14983 25324
rect 12408 25238 12432 25272
rect 12466 25238 12501 25272
rect 12535 25238 12570 25272
rect 12604 25238 12639 25272
rect 12673 25238 12708 25272
rect 12742 25238 12777 25272
rect 12811 25238 12846 25272
rect 12880 25238 12915 25272
rect 12949 25238 12984 25272
rect 13018 25238 13053 25272
rect 13087 25238 13122 25272
rect 13156 25238 13191 25272
rect 13225 25238 13260 25272
rect 13294 25238 13328 25272
rect 13362 25238 13396 25272
rect 13430 25238 13464 25272
rect 13498 25238 13532 25272
rect 13566 25238 13600 25272
rect 13634 25238 13668 25272
rect 13702 25238 13736 25272
rect 13770 25238 13804 25272
rect 13838 25238 13872 25272
rect 13906 25238 13940 25272
rect 13974 25238 14008 25272
rect 14042 25238 14076 25272
rect 14110 25238 14144 25272
rect 14178 25238 14212 25272
rect 14246 25238 14280 25272
rect 14314 25238 14348 25272
rect 14382 25238 14416 25272
rect 14450 25238 14484 25272
rect 14518 25238 14552 25272
rect 14586 25238 14620 25272
rect 14654 25238 14688 25272
rect 14722 25238 14756 25272
rect 14790 25238 14824 25272
rect 14858 25238 14983 25272
rect 12408 25180 14983 25238
rect -41 25178 14983 25180
rect -41 25144 124 25178
rect 158 25144 193 25178
rect 227 25144 262 25178
rect 296 25144 331 25178
rect 365 25144 400 25178
rect 434 25144 469 25178
rect 503 25144 538 25178
rect 572 25144 607 25178
rect 641 25144 676 25178
rect 710 25144 745 25178
rect 779 25144 814 25178
rect 848 25144 883 25178
rect 917 25144 952 25178
rect 986 25144 1020 25178
rect 1054 25144 1088 25178
rect 1122 25144 1156 25178
rect 1190 25144 1224 25178
rect 1258 25144 1292 25178
rect 1326 25144 1360 25178
rect 1394 25144 1428 25178
rect 1462 25144 1496 25178
rect 1530 25144 1564 25178
rect 1598 25144 1632 25178
rect 1666 25144 1700 25178
rect 1734 25144 1768 25178
rect 1802 25144 1836 25178
rect 1870 25144 1904 25178
rect 1938 25144 1972 25178
rect 2006 25144 2040 25178
rect 2074 25144 2108 25178
rect 2142 25144 2176 25178
rect 2210 25144 2244 25178
rect 2278 25144 2312 25178
rect 2346 25144 2380 25178
rect 2414 25144 2448 25178
rect 2482 25144 2516 25178
rect 2550 25144 2584 25178
rect 2618 25144 2652 25178
rect 2686 25144 2720 25178
rect 2754 25144 2788 25178
rect 2822 25144 2856 25178
rect 2890 25144 2924 25178
rect 2958 25144 2992 25178
rect 3026 25144 3060 25178
rect 3094 25144 3128 25178
rect 3162 25144 3196 25178
rect 3230 25144 3264 25178
rect 3298 25144 3332 25178
rect 3366 25144 3400 25178
rect 3434 25144 3468 25178
rect 3502 25144 3536 25178
rect 3570 25144 3604 25178
rect 3638 25144 3672 25178
rect 3706 25144 3740 25178
rect 3774 25144 3808 25178
rect 3842 25144 3876 25178
rect 3910 25144 3944 25178
rect 3978 25144 4012 25178
rect 4046 25144 4080 25178
rect 4114 25144 4148 25178
rect 4182 25144 4216 25178
rect 4250 25144 4284 25178
rect 4318 25144 4352 25178
rect 4386 25144 4420 25178
rect 4454 25144 4488 25178
rect 4522 25144 4556 25178
rect 4590 25144 4624 25178
rect 4658 25144 4692 25178
rect 4726 25144 4760 25178
rect 4794 25144 4828 25178
rect 4862 25144 4896 25178
rect 4930 25144 4964 25178
rect 4998 25144 5032 25178
rect 5066 25144 5100 25178
rect 5134 25144 5168 25178
rect 5202 25144 5236 25178
rect 5270 25144 5304 25178
rect 5338 25144 5372 25178
rect 5406 25144 5440 25178
rect 5474 25144 5508 25178
rect 5542 25144 5576 25178
rect 5610 25144 5644 25178
rect 5678 25144 5712 25178
rect 5746 25144 5780 25178
rect 5814 25144 5848 25178
rect 5882 25144 5916 25178
rect 5950 25144 5984 25178
rect 6018 25144 6052 25178
rect 6086 25144 6120 25178
rect 6154 25144 6188 25178
rect 6222 25144 6256 25178
rect 6290 25144 6324 25178
rect 6358 25144 6392 25178
rect 6426 25144 6460 25178
rect 6494 25144 6528 25178
rect 6562 25144 6596 25178
rect 6630 25144 6664 25178
rect 6698 25144 6732 25178
rect 6766 25144 6800 25178
rect 6834 25144 6868 25178
rect 6902 25144 6936 25178
rect 6970 25144 7004 25178
rect 7038 25144 7072 25178
rect 7106 25144 7140 25178
rect 7174 25144 7208 25178
rect 7242 25144 7276 25178
rect 7310 25144 7344 25178
rect 7378 25144 7412 25178
rect 7446 25144 7480 25178
rect 7514 25144 7548 25178
rect 7582 25144 7616 25178
rect 7650 25144 7684 25178
rect 7718 25144 7752 25178
rect 7786 25144 7820 25178
rect 7854 25144 7888 25178
rect 7922 25144 7956 25178
rect 7990 25144 8024 25178
rect 8058 25144 8092 25178
rect 8126 25144 8160 25178
rect 8194 25144 8228 25178
rect 8262 25144 8296 25178
rect 8330 25144 8364 25178
rect 8398 25144 8432 25178
rect 8466 25144 8500 25178
rect 8534 25144 8568 25178
rect 8602 25144 8636 25178
rect 8670 25144 8704 25178
rect 8738 25144 8772 25178
rect 8806 25144 8840 25178
rect 8874 25144 8908 25178
rect 8942 25144 8976 25178
rect 9010 25144 9044 25178
rect 9078 25144 9112 25178
rect 9146 25144 9180 25178
rect 9214 25144 9248 25178
rect 9282 25144 9316 25178
rect 9350 25144 9384 25178
rect 9418 25144 9452 25178
rect 9486 25144 9520 25178
rect 9554 25144 9588 25178
rect 9622 25144 9656 25178
rect 9690 25144 9724 25178
rect 9758 25144 9792 25178
rect 9826 25144 9860 25178
rect 9894 25144 9928 25178
rect 9962 25144 9996 25178
rect 10030 25144 10064 25178
rect 10098 25144 10132 25178
rect 10166 25144 10200 25178
rect 10234 25144 10268 25178
rect 10302 25144 10336 25178
rect 10370 25144 10404 25178
rect 10438 25144 10472 25178
rect 10506 25144 10540 25178
rect 10574 25144 10608 25178
rect 10642 25144 10676 25178
rect 10710 25144 10744 25178
rect 10778 25144 10812 25178
rect 10846 25144 10880 25178
rect 10914 25144 10948 25178
rect 10982 25144 11016 25178
rect 11050 25144 11084 25178
rect 11118 25144 11152 25178
rect 11186 25144 11220 25178
rect 11254 25144 11288 25178
rect 11322 25144 11356 25178
rect 11390 25144 11424 25178
rect 11458 25144 11492 25178
rect 11526 25144 11560 25178
rect 11594 25144 11628 25178
rect 11662 25144 11696 25178
rect 11730 25144 11764 25178
rect 11798 25144 11832 25178
rect 11866 25144 11900 25178
rect 11934 25144 11968 25178
rect 12002 25144 12036 25178
rect 12070 25144 12104 25178
rect 12138 25144 12172 25178
rect 12206 25144 12240 25178
rect 12274 25144 12308 25178
rect 12342 25144 12376 25178
rect 12410 25144 12444 25178
rect 12478 25144 12512 25178
rect 12546 25144 12580 25178
rect 12614 25144 12648 25178
rect 12682 25144 12716 25178
rect 12750 25144 12784 25178
rect 12818 25144 12852 25178
rect 12886 25144 12920 25178
rect 12954 25144 12988 25178
rect 13022 25144 13056 25178
rect 13090 25144 13124 25178
rect 13158 25144 13192 25178
rect 13226 25144 13260 25178
rect 13294 25144 13328 25178
rect 13362 25144 13396 25178
rect 13430 25144 13464 25178
rect 13498 25144 13532 25178
rect 13566 25144 13600 25178
rect 13634 25144 13668 25178
rect 13702 25144 13736 25178
rect 13770 25144 13804 25178
rect 13838 25144 13872 25178
rect 13906 25144 13940 25178
rect 13974 25144 14008 25178
rect 14042 25144 14076 25178
rect 14110 25144 14144 25178
rect 14178 25144 14212 25178
rect 14246 25144 14280 25178
rect 14314 25144 14348 25178
rect 14382 25144 14416 25178
rect 14450 25144 14484 25178
rect 14518 25144 14552 25178
rect 14586 25144 14620 25178
rect 14654 25144 14688 25178
rect 14722 25144 14756 25178
rect 14790 25144 14824 25178
rect 14858 25144 14983 25178
rect -41 25106 14983 25144
rect -41 25072 124 25106
rect 158 25072 193 25106
rect 227 25072 262 25106
rect 296 25072 331 25106
rect 365 25072 400 25106
rect 434 25072 469 25106
rect 503 25072 538 25106
rect 572 25072 607 25106
rect 641 25072 676 25106
rect 710 25072 745 25106
rect 779 25072 814 25106
rect 848 25072 883 25106
rect 917 25072 952 25106
rect 986 25072 1020 25106
rect 1054 25072 1088 25106
rect 1122 25072 1156 25106
rect 1190 25072 1224 25106
rect 1258 25072 1292 25106
rect 1326 25072 1360 25106
rect 1394 25072 1428 25106
rect 1462 25072 1496 25106
rect 1530 25072 1564 25106
rect 1598 25072 1632 25106
rect 1666 25072 1700 25106
rect 1734 25072 1768 25106
rect 1802 25072 1836 25106
rect 1870 25072 1904 25106
rect 1938 25072 1972 25106
rect 2006 25072 2040 25106
rect 2074 25072 2108 25106
rect 2142 25072 2176 25106
rect 2210 25072 2244 25106
rect 2278 25072 2312 25106
rect 2346 25072 2380 25106
rect 2414 25072 2448 25106
rect 2482 25072 2516 25106
rect 2550 25072 2584 25106
rect 2618 25072 2652 25106
rect 2686 25072 2720 25106
rect 2754 25072 2788 25106
rect 2822 25072 2856 25106
rect 2890 25072 2924 25106
rect 2958 25072 2992 25106
rect 3026 25072 3060 25106
rect 3094 25072 3128 25106
rect 3162 25072 3196 25106
rect 3230 25072 3264 25106
rect 3298 25072 3332 25106
rect 3366 25072 3400 25106
rect 3434 25072 3468 25106
rect 3502 25072 3536 25106
rect 3570 25072 3604 25106
rect 3638 25072 3672 25106
rect 3706 25072 3740 25106
rect 3774 25072 3808 25106
rect 3842 25072 3876 25106
rect 3910 25072 3944 25106
rect 3978 25072 4012 25106
rect 4046 25072 4080 25106
rect 4114 25072 4148 25106
rect 4182 25072 4216 25106
rect 4250 25072 4284 25106
rect 4318 25072 4352 25106
rect 4386 25072 4420 25106
rect 4454 25072 4488 25106
rect 4522 25072 4556 25106
rect 4590 25072 4624 25106
rect 4658 25072 4692 25106
rect 4726 25072 4760 25106
rect 4794 25072 4828 25106
rect 4862 25072 4896 25106
rect 4930 25072 4964 25106
rect 4998 25072 5032 25106
rect 5066 25072 5100 25106
rect 5134 25072 5168 25106
rect 5202 25072 5236 25106
rect 5270 25072 5304 25106
rect 5338 25072 5372 25106
rect 5406 25072 5440 25106
rect 5474 25072 5508 25106
rect 5542 25072 5576 25106
rect 5610 25072 5644 25106
rect 5678 25072 5712 25106
rect 5746 25072 5780 25106
rect 5814 25072 5848 25106
rect 5882 25072 5916 25106
rect 5950 25072 5984 25106
rect 6018 25072 6052 25106
rect 6086 25072 6120 25106
rect 6154 25072 6188 25106
rect 6222 25072 6256 25106
rect 6290 25072 6324 25106
rect 6358 25072 6392 25106
rect 6426 25072 6460 25106
rect 6494 25072 6528 25106
rect 6562 25072 6596 25106
rect 6630 25072 6664 25106
rect 6698 25072 6732 25106
rect 6766 25072 6800 25106
rect 6834 25072 6868 25106
rect 6902 25072 6936 25106
rect 6970 25072 7004 25106
rect 7038 25072 7072 25106
rect 7106 25072 7140 25106
rect 7174 25072 7208 25106
rect 7242 25072 7276 25106
rect 7310 25072 7344 25106
rect 7378 25072 7412 25106
rect 7446 25072 7480 25106
rect 7514 25072 7548 25106
rect 7582 25072 7616 25106
rect 7650 25072 7684 25106
rect 7718 25072 7752 25106
rect 7786 25072 7820 25106
rect 7854 25072 7888 25106
rect 7922 25072 7956 25106
rect 7990 25072 8024 25106
rect 8058 25072 8092 25106
rect 8126 25072 8160 25106
rect 8194 25072 8228 25106
rect 8262 25072 8296 25106
rect 8330 25072 8364 25106
rect 8398 25072 8432 25106
rect 8466 25072 8500 25106
rect 8534 25072 8568 25106
rect 8602 25072 8636 25106
rect 8670 25072 8704 25106
rect 8738 25072 8772 25106
rect 8806 25072 8840 25106
rect 8874 25072 8908 25106
rect 8942 25072 8976 25106
rect 9010 25072 9044 25106
rect 9078 25072 9112 25106
rect 9146 25072 9180 25106
rect 9214 25072 9248 25106
rect 9282 25072 9316 25106
rect 9350 25072 9384 25106
rect 9418 25072 9452 25106
rect 9486 25072 9520 25106
rect 9554 25072 9588 25106
rect 9622 25072 9656 25106
rect 9690 25072 9724 25106
rect 9758 25072 9792 25106
rect 9826 25072 9860 25106
rect 9894 25072 9928 25106
rect 9962 25072 9996 25106
rect 10030 25072 10064 25106
rect 10098 25072 10132 25106
rect 10166 25072 10200 25106
rect 10234 25072 10268 25106
rect 10302 25072 10336 25106
rect 10370 25072 10404 25106
rect 10438 25072 10472 25106
rect 10506 25072 10540 25106
rect 10574 25072 10608 25106
rect 10642 25072 10676 25106
rect 10710 25072 10744 25106
rect 10778 25072 10812 25106
rect 10846 25072 10880 25106
rect 10914 25072 10948 25106
rect 10982 25072 11016 25106
rect 11050 25072 11084 25106
rect 11118 25072 11152 25106
rect 11186 25072 11220 25106
rect 11254 25072 11288 25106
rect 11322 25072 11356 25106
rect 11390 25072 11424 25106
rect 11458 25072 11492 25106
rect 11526 25072 11560 25106
rect 11594 25072 11628 25106
rect 11662 25072 11696 25106
rect 11730 25072 11764 25106
rect 11798 25072 11832 25106
rect 11866 25072 11900 25106
rect 11934 25072 11968 25106
rect 12002 25072 12036 25106
rect 12070 25072 12104 25106
rect 12138 25072 12172 25106
rect 12206 25072 12240 25106
rect 12274 25072 12308 25106
rect 12342 25072 12376 25106
rect 12410 25072 12444 25106
rect 12478 25072 12512 25106
rect 12546 25072 12580 25106
rect 12614 25072 12648 25106
rect 12682 25072 12716 25106
rect 12750 25072 12784 25106
rect 12818 25072 12852 25106
rect 12886 25072 12920 25106
rect 12954 25072 12988 25106
rect 13022 25072 13056 25106
rect 13090 25072 13124 25106
rect 13158 25072 13192 25106
rect 13226 25072 13260 25106
rect 13294 25072 13328 25106
rect 13362 25072 13396 25106
rect 13430 25072 13464 25106
rect 13498 25072 13532 25106
rect 13566 25072 13600 25106
rect 13634 25072 13668 25106
rect 13702 25072 13736 25106
rect 13770 25072 13804 25106
rect 13838 25072 13872 25106
rect 13906 25072 13940 25106
rect 13974 25072 14008 25106
rect 14042 25072 14076 25106
rect 14110 25072 14144 25106
rect 14178 25072 14212 25106
rect 14246 25072 14280 25106
rect 14314 25072 14348 25106
rect 14382 25072 14416 25106
rect 14450 25072 14484 25106
rect 14518 25072 14552 25106
rect 14586 25072 14620 25106
rect 14654 25072 14688 25106
rect 14722 25072 14756 25106
rect 14790 25072 14824 25106
rect 14858 25072 14983 25106
rect -41 25041 14983 25072
rect -41 25007 88 25041
rect 122 25034 161 25041
rect 195 25034 234 25041
rect 268 25034 307 25041
rect 341 25034 380 25041
rect 414 25034 453 25041
rect 487 25034 526 25041
rect 560 25034 599 25041
rect 633 25034 672 25041
rect 706 25034 745 25041
rect 779 25034 818 25041
rect 852 25034 891 25041
rect 925 25034 964 25041
rect 998 25034 1037 25041
rect 1071 25034 1110 25041
rect 1144 25034 1183 25041
rect 1217 25034 1256 25041
rect 1290 25034 1329 25041
rect 1363 25034 1402 25041
rect 1436 25034 1475 25041
rect 1509 25034 1548 25041
rect 1582 25034 1621 25041
rect 1655 25034 1694 25041
rect 1728 25034 1767 25041
rect 1801 25034 1840 25041
rect 1874 25034 1913 25041
rect 1947 25034 1986 25041
rect 2020 25034 2059 25041
rect 2093 25034 2132 25041
rect 2166 25034 2205 25041
rect 2239 25034 2278 25041
rect 122 25007 124 25034
rect -41 25000 124 25007
rect 158 25007 161 25034
rect 227 25007 234 25034
rect 296 25007 307 25034
rect 365 25007 380 25034
rect 434 25007 453 25034
rect 503 25007 526 25034
rect 572 25007 599 25034
rect 641 25007 672 25034
rect 158 25000 193 25007
rect 227 25000 262 25007
rect 296 25000 331 25007
rect 365 25000 400 25007
rect 434 25000 469 25007
rect 503 25000 538 25007
rect 572 25000 607 25007
rect 641 25000 676 25007
rect 710 25000 745 25034
rect 779 25000 814 25034
rect 852 25007 883 25034
rect 925 25007 952 25034
rect 998 25007 1020 25034
rect 1071 25007 1088 25034
rect 1144 25007 1156 25034
rect 1217 25007 1224 25034
rect 1290 25007 1292 25034
rect 848 25000 883 25007
rect 917 25000 952 25007
rect 986 25000 1020 25007
rect 1054 25000 1088 25007
rect 1122 25000 1156 25007
rect 1190 25000 1224 25007
rect 1258 25000 1292 25007
rect 1326 25007 1329 25034
rect 1394 25007 1402 25034
rect 1462 25007 1475 25034
rect 1530 25007 1548 25034
rect 1598 25007 1621 25034
rect 1666 25007 1694 25034
rect 1734 25007 1767 25034
rect 1326 25000 1360 25007
rect 1394 25000 1428 25007
rect 1462 25000 1496 25007
rect 1530 25000 1564 25007
rect 1598 25000 1632 25007
rect 1666 25000 1700 25007
rect 1734 25000 1768 25007
rect 1802 25000 1836 25034
rect 1874 25007 1904 25034
rect 1947 25007 1972 25034
rect 2020 25007 2040 25034
rect 2093 25007 2108 25034
rect 2166 25007 2176 25034
rect 2239 25007 2244 25034
rect 1870 25000 1904 25007
rect 1938 25000 1972 25007
rect 2006 25000 2040 25007
rect 2074 25000 2108 25007
rect 2142 25000 2176 25007
rect 2210 25000 2244 25007
rect 2312 25034 2351 25041
rect 2385 25034 2424 25041
rect 2458 25034 2497 25041
rect 2531 25034 2570 25041
rect 2604 25034 2643 25041
rect 2677 25034 2716 25041
rect 2750 25034 2789 25041
rect 2823 25034 2862 25041
rect 2896 25034 2935 25041
rect 2969 25034 3008 25041
rect 3042 25034 3081 25041
rect 3115 25034 3154 25041
rect 3188 25034 3227 25041
rect 3261 25034 3300 25041
rect 3334 25034 3373 25041
rect 3407 25034 3446 25041
rect 3480 25034 3519 25041
rect 3553 25034 3592 25041
rect 3626 25034 3665 25041
rect 3699 25034 3738 25041
rect 3772 25034 3811 25041
rect 3845 25034 3884 25041
rect 3918 25034 3957 25041
rect 3991 25034 4030 25041
rect 4064 25034 4103 25041
rect 4137 25034 4176 25041
rect 4210 25034 4249 25041
rect 4283 25034 4322 25041
rect 4356 25034 4395 25041
rect 4429 25034 4468 25041
rect 2278 25000 2312 25007
rect 2346 25007 2351 25034
rect 2414 25007 2424 25034
rect 2482 25007 2497 25034
rect 2550 25007 2570 25034
rect 2618 25007 2643 25034
rect 2686 25007 2716 25034
rect 2346 25000 2380 25007
rect 2414 25000 2448 25007
rect 2482 25000 2516 25007
rect 2550 25000 2584 25007
rect 2618 25000 2652 25007
rect 2686 25000 2720 25007
rect 2754 25000 2788 25034
rect 2823 25007 2856 25034
rect 2896 25007 2924 25034
rect 2969 25007 2992 25034
rect 3042 25007 3060 25034
rect 3115 25007 3128 25034
rect 3188 25007 3196 25034
rect 3261 25007 3264 25034
rect 2822 25000 2856 25007
rect 2890 25000 2924 25007
rect 2958 25000 2992 25007
rect 3026 25000 3060 25007
rect 3094 25000 3128 25007
rect 3162 25000 3196 25007
rect 3230 25000 3264 25007
rect 3298 25007 3300 25034
rect 3366 25007 3373 25034
rect 3434 25007 3446 25034
rect 3502 25007 3519 25034
rect 3570 25007 3592 25034
rect 3638 25007 3665 25034
rect 3706 25007 3738 25034
rect 3298 25000 3332 25007
rect 3366 25000 3400 25007
rect 3434 25000 3468 25007
rect 3502 25000 3536 25007
rect 3570 25000 3604 25007
rect 3638 25000 3672 25007
rect 3706 25000 3740 25007
rect 3774 25000 3808 25034
rect 3845 25007 3876 25034
rect 3918 25007 3944 25034
rect 3991 25007 4012 25034
rect 4064 25007 4080 25034
rect 4137 25007 4148 25034
rect 4210 25007 4216 25034
rect 4283 25007 4284 25034
rect 3842 25000 3876 25007
rect 3910 25000 3944 25007
rect 3978 25000 4012 25007
rect 4046 25000 4080 25007
rect 4114 25000 4148 25007
rect 4182 25000 4216 25007
rect 4250 25000 4284 25007
rect 4318 25007 4322 25034
rect 4386 25007 4395 25034
rect 4318 25000 4352 25007
rect 4386 25000 4420 25007
rect 4454 25000 4468 25034
rect -41 24969 4468 25000
rect -41 24935 88 24969
rect 122 24962 161 24969
rect 195 24962 234 24969
rect 268 24962 307 24969
rect 341 24962 380 24969
rect 414 24962 453 24969
rect 487 24962 526 24969
rect 560 24962 599 24969
rect 633 24962 672 24969
rect 706 24962 745 24969
rect 779 24962 818 24969
rect 852 24962 891 24969
rect 925 24962 964 24969
rect 998 24962 1037 24969
rect 1071 24962 1110 24969
rect 1144 24962 1183 24969
rect 1217 24962 1256 24969
rect 1290 24962 1329 24969
rect 1363 24962 1402 24969
rect 1436 24962 1475 24969
rect 1509 24962 1548 24969
rect 1582 24962 1621 24969
rect 1655 24962 1694 24969
rect 1728 24962 1767 24969
rect 1801 24962 1840 24969
rect 1874 24962 1913 24969
rect 1947 24962 1986 24969
rect 2020 24962 2059 24969
rect 2093 24962 2132 24969
rect 2166 24962 2205 24969
rect 2239 24962 2278 24969
rect 122 24935 124 24962
rect -41 24928 124 24935
rect 158 24935 161 24962
rect 227 24935 234 24962
rect 296 24935 307 24962
rect 365 24935 380 24962
rect 434 24935 453 24962
rect 503 24935 526 24962
rect 572 24935 599 24962
rect 641 24935 672 24962
rect 158 24928 193 24935
rect 227 24928 262 24935
rect 296 24928 331 24935
rect 365 24928 400 24935
rect 434 24928 469 24935
rect 503 24928 538 24935
rect 572 24928 607 24935
rect 641 24928 676 24935
rect 710 24928 745 24962
rect 779 24928 814 24962
rect 852 24935 883 24962
rect 925 24935 952 24962
rect 998 24935 1020 24962
rect 1071 24935 1088 24962
rect 1144 24935 1156 24962
rect 1217 24935 1224 24962
rect 1290 24935 1292 24962
rect 848 24928 883 24935
rect 917 24928 952 24935
rect 986 24928 1020 24935
rect 1054 24928 1088 24935
rect 1122 24928 1156 24935
rect 1190 24928 1224 24935
rect 1258 24928 1292 24935
rect 1326 24935 1329 24962
rect 1394 24935 1402 24962
rect 1462 24935 1475 24962
rect 1530 24935 1548 24962
rect 1598 24935 1621 24962
rect 1666 24935 1694 24962
rect 1734 24935 1767 24962
rect 1326 24928 1360 24935
rect 1394 24928 1428 24935
rect 1462 24928 1496 24935
rect 1530 24928 1564 24935
rect 1598 24928 1632 24935
rect 1666 24928 1700 24935
rect 1734 24928 1768 24935
rect 1802 24928 1836 24962
rect 1874 24935 1904 24962
rect 1947 24935 1972 24962
rect 2020 24935 2040 24962
rect 2093 24935 2108 24962
rect 2166 24935 2176 24962
rect 2239 24935 2244 24962
rect 1870 24928 1904 24935
rect 1938 24928 1972 24935
rect 2006 24928 2040 24935
rect 2074 24928 2108 24935
rect 2142 24928 2176 24935
rect 2210 24928 2244 24935
rect 2312 24962 2351 24969
rect 2385 24962 2424 24969
rect 2458 24962 2497 24969
rect 2531 24962 2570 24969
rect 2604 24962 2643 24969
rect 2677 24962 2716 24969
rect 2750 24962 2789 24969
rect 2823 24962 2862 24969
rect 2896 24962 2935 24969
rect 2969 24962 3008 24969
rect 3042 24962 3081 24969
rect 3115 24962 3154 24969
rect 3188 24962 3227 24969
rect 3261 24962 3300 24969
rect 3334 24962 3373 24969
rect 3407 24962 3446 24969
rect 3480 24962 3519 24969
rect 3553 24962 3592 24969
rect 3626 24962 3665 24969
rect 3699 24962 3738 24969
rect 3772 24962 3811 24969
rect 3845 24962 3884 24969
rect 3918 24962 3957 24969
rect 3991 24962 4030 24969
rect 4064 24962 4103 24969
rect 4137 24962 4176 24969
rect 4210 24962 4249 24969
rect 4283 24962 4322 24969
rect 4356 24962 4395 24969
rect 4429 24962 4468 24969
rect 2278 24928 2312 24935
rect 2346 24935 2351 24962
rect 2414 24935 2424 24962
rect 2482 24935 2497 24962
rect 2550 24935 2570 24962
rect 2618 24935 2643 24962
rect 2686 24935 2716 24962
rect 2346 24928 2380 24935
rect 2414 24928 2448 24935
rect 2482 24928 2516 24935
rect 2550 24928 2584 24935
rect 2618 24928 2652 24935
rect 2686 24928 2720 24935
rect 2754 24928 2788 24962
rect 2823 24935 2856 24962
rect 2896 24935 2924 24962
rect 2969 24935 2992 24962
rect 3042 24935 3060 24962
rect 3115 24935 3128 24962
rect 3188 24935 3196 24962
rect 3261 24935 3264 24962
rect 2822 24928 2856 24935
rect 2890 24928 2924 24935
rect 2958 24928 2992 24935
rect 3026 24928 3060 24935
rect 3094 24928 3128 24935
rect 3162 24928 3196 24935
rect 3230 24928 3264 24935
rect 3298 24935 3300 24962
rect 3366 24935 3373 24962
rect 3434 24935 3446 24962
rect 3502 24935 3519 24962
rect 3570 24935 3592 24962
rect 3638 24935 3665 24962
rect 3706 24935 3738 24962
rect 3298 24928 3332 24935
rect 3366 24928 3400 24935
rect 3434 24928 3468 24935
rect 3502 24928 3536 24935
rect 3570 24928 3604 24935
rect 3638 24928 3672 24935
rect 3706 24928 3740 24935
rect 3774 24928 3808 24962
rect 3845 24935 3876 24962
rect 3918 24935 3944 24962
rect 3991 24935 4012 24962
rect 4064 24935 4080 24962
rect 4137 24935 4148 24962
rect 4210 24935 4216 24962
rect 4283 24935 4284 24962
rect 3842 24928 3876 24935
rect 3910 24928 3944 24935
rect 3978 24928 4012 24935
rect 4046 24928 4080 24935
rect 4114 24928 4148 24935
rect 4182 24928 4216 24935
rect 4250 24928 4284 24935
rect 4318 24935 4322 24962
rect 4386 24935 4395 24962
rect 4318 24928 4352 24935
rect 4386 24928 4420 24935
rect 4454 24928 4468 24962
rect -41 24897 4468 24928
rect -41 24863 88 24897
rect 122 24890 161 24897
rect 195 24890 234 24897
rect 268 24890 307 24897
rect 341 24890 380 24897
rect 414 24890 453 24897
rect 487 24890 526 24897
rect 560 24890 599 24897
rect 633 24890 672 24897
rect 706 24890 745 24897
rect 779 24890 818 24897
rect 852 24890 891 24897
rect 925 24890 964 24897
rect 998 24890 1037 24897
rect 1071 24890 1110 24897
rect 1144 24890 1183 24897
rect 1217 24890 1256 24897
rect 1290 24890 1329 24897
rect 1363 24890 1402 24897
rect 1436 24890 1475 24897
rect 1509 24890 1548 24897
rect 1582 24890 1621 24897
rect 1655 24890 1694 24897
rect 1728 24890 1767 24897
rect 1801 24890 1840 24897
rect 1874 24890 1913 24897
rect 1947 24890 1986 24897
rect 2020 24890 2059 24897
rect 2093 24890 2132 24897
rect 2166 24890 2205 24897
rect 2239 24890 2278 24897
rect 122 24863 124 24890
rect -41 24856 124 24863
rect 158 24863 161 24890
rect 227 24863 234 24890
rect 296 24863 307 24890
rect 365 24863 380 24890
rect 434 24863 453 24890
rect 503 24863 526 24890
rect 572 24863 599 24890
rect 641 24863 672 24890
rect 158 24856 193 24863
rect 227 24856 262 24863
rect 296 24856 331 24863
rect 365 24856 400 24863
rect 434 24856 469 24863
rect 503 24856 538 24863
rect 572 24856 607 24863
rect 641 24856 676 24863
rect 710 24856 745 24890
rect 779 24856 814 24890
rect 852 24863 883 24890
rect 925 24863 952 24890
rect 998 24863 1020 24890
rect 1071 24863 1088 24890
rect 1144 24863 1156 24890
rect 1217 24863 1224 24890
rect 1290 24863 1292 24890
rect 848 24856 883 24863
rect 917 24856 952 24863
rect 986 24856 1020 24863
rect 1054 24856 1088 24863
rect 1122 24856 1156 24863
rect 1190 24856 1224 24863
rect 1258 24856 1292 24863
rect 1326 24863 1329 24890
rect 1394 24863 1402 24890
rect 1462 24863 1475 24890
rect 1530 24863 1548 24890
rect 1598 24863 1621 24890
rect 1666 24863 1694 24890
rect 1734 24863 1767 24890
rect 1326 24856 1360 24863
rect 1394 24856 1428 24863
rect 1462 24856 1496 24863
rect 1530 24856 1564 24863
rect 1598 24856 1632 24863
rect 1666 24856 1700 24863
rect 1734 24856 1768 24863
rect 1802 24856 1836 24890
rect 1874 24863 1904 24890
rect 1947 24863 1972 24890
rect 2020 24863 2040 24890
rect 2093 24863 2108 24890
rect 2166 24863 2176 24890
rect 2239 24863 2244 24890
rect 1870 24856 1904 24863
rect 1938 24856 1972 24863
rect 2006 24856 2040 24863
rect 2074 24856 2108 24863
rect 2142 24856 2176 24863
rect 2210 24856 2244 24863
rect 2312 24890 2351 24897
rect 2385 24890 2424 24897
rect 2458 24890 2497 24897
rect 2531 24890 2570 24897
rect 2604 24890 2643 24897
rect 2677 24890 2716 24897
rect 2750 24890 2789 24897
rect 2823 24890 2862 24897
rect 2896 24890 2935 24897
rect 2969 24890 3008 24897
rect 3042 24890 3081 24897
rect 3115 24890 3154 24897
rect 3188 24890 3227 24897
rect 3261 24890 3300 24897
rect 3334 24890 3373 24897
rect 3407 24890 3446 24897
rect 3480 24890 3519 24897
rect 3553 24890 3592 24897
rect 3626 24890 3665 24897
rect 3699 24890 3738 24897
rect 3772 24890 3811 24897
rect 3845 24890 3884 24897
rect 3918 24890 3957 24897
rect 3991 24890 4030 24897
rect 4064 24890 4103 24897
rect 4137 24890 4176 24897
rect 4210 24890 4249 24897
rect 4283 24890 4322 24897
rect 4356 24890 4395 24897
rect 4429 24890 4468 24897
rect 2278 24856 2312 24863
rect 2346 24863 2351 24890
rect 2414 24863 2424 24890
rect 2482 24863 2497 24890
rect 2550 24863 2570 24890
rect 2618 24863 2643 24890
rect 2686 24863 2716 24890
rect 2346 24856 2380 24863
rect 2414 24856 2448 24863
rect 2482 24856 2516 24863
rect 2550 24856 2584 24863
rect 2618 24856 2652 24863
rect 2686 24856 2720 24863
rect 2754 24856 2788 24890
rect 2823 24863 2856 24890
rect 2896 24863 2924 24890
rect 2969 24863 2992 24890
rect 3042 24863 3060 24890
rect 3115 24863 3128 24890
rect 3188 24863 3196 24890
rect 3261 24863 3264 24890
rect 2822 24856 2856 24863
rect 2890 24856 2924 24863
rect 2958 24856 2992 24863
rect 3026 24856 3060 24863
rect 3094 24856 3128 24863
rect 3162 24856 3196 24863
rect 3230 24856 3264 24863
rect 3298 24863 3300 24890
rect 3366 24863 3373 24890
rect 3434 24863 3446 24890
rect 3502 24863 3519 24890
rect 3570 24863 3592 24890
rect 3638 24863 3665 24890
rect 3706 24863 3738 24890
rect 3298 24856 3332 24863
rect 3366 24856 3400 24863
rect 3434 24856 3468 24863
rect 3502 24856 3536 24863
rect 3570 24856 3604 24863
rect 3638 24856 3672 24863
rect 3706 24856 3740 24863
rect 3774 24856 3808 24890
rect 3845 24863 3876 24890
rect 3918 24863 3944 24890
rect 3991 24863 4012 24890
rect 4064 24863 4080 24890
rect 4137 24863 4148 24890
rect 4210 24863 4216 24890
rect 4283 24863 4284 24890
rect 3842 24856 3876 24863
rect 3910 24856 3944 24863
rect 3978 24856 4012 24863
rect 4046 24856 4080 24863
rect 4114 24856 4148 24863
rect 4182 24856 4216 24863
rect 4250 24856 4284 24863
rect 4318 24863 4322 24890
rect 4386 24863 4395 24890
rect 4318 24856 4352 24863
rect 4386 24856 4420 24863
rect 4454 24856 4468 24890
rect -41 24825 4468 24856
rect -41 24791 88 24825
rect 122 24818 161 24825
rect 195 24818 234 24825
rect 268 24818 307 24825
rect 341 24818 380 24825
rect 414 24818 453 24825
rect 487 24818 526 24825
rect 560 24818 599 24825
rect 633 24818 672 24825
rect 706 24818 745 24825
rect 779 24818 818 24825
rect 852 24818 891 24825
rect 925 24818 964 24825
rect 998 24818 1037 24825
rect 1071 24818 1110 24825
rect 1144 24818 1183 24825
rect 1217 24818 1256 24825
rect 1290 24818 1329 24825
rect 1363 24818 1402 24825
rect 1436 24818 1475 24825
rect 1509 24818 1548 24825
rect 1582 24818 1621 24825
rect 1655 24818 1694 24825
rect 1728 24818 1767 24825
rect 1801 24818 1840 24825
rect 1874 24818 1913 24825
rect 1947 24818 1986 24825
rect 2020 24818 2059 24825
rect 2093 24818 2132 24825
rect 2166 24818 2205 24825
rect 2239 24818 2278 24825
rect 122 24791 124 24818
rect -41 24784 124 24791
rect 158 24791 161 24818
rect 227 24791 234 24818
rect 296 24791 307 24818
rect 365 24791 380 24818
rect 434 24791 453 24818
rect 503 24791 526 24818
rect 572 24791 599 24818
rect 641 24791 672 24818
rect 158 24784 193 24791
rect 227 24784 262 24791
rect 296 24784 331 24791
rect 365 24784 400 24791
rect 434 24784 469 24791
rect 503 24784 538 24791
rect 572 24784 607 24791
rect 641 24784 676 24791
rect 710 24784 745 24818
rect 779 24784 814 24818
rect 852 24791 883 24818
rect 925 24791 952 24818
rect 998 24791 1020 24818
rect 1071 24791 1088 24818
rect 1144 24791 1156 24818
rect 1217 24791 1224 24818
rect 1290 24791 1292 24818
rect 848 24784 883 24791
rect 917 24784 952 24791
rect 986 24784 1020 24791
rect 1054 24784 1088 24791
rect 1122 24784 1156 24791
rect 1190 24784 1224 24791
rect 1258 24784 1292 24791
rect 1326 24791 1329 24818
rect 1394 24791 1402 24818
rect 1462 24791 1475 24818
rect 1530 24791 1548 24818
rect 1598 24791 1621 24818
rect 1666 24791 1694 24818
rect 1734 24791 1767 24818
rect 1326 24784 1360 24791
rect 1394 24784 1428 24791
rect 1462 24784 1496 24791
rect 1530 24784 1564 24791
rect 1598 24784 1632 24791
rect 1666 24784 1700 24791
rect 1734 24784 1768 24791
rect 1802 24784 1836 24818
rect 1874 24791 1904 24818
rect 1947 24791 1972 24818
rect 2020 24791 2040 24818
rect 2093 24791 2108 24818
rect 2166 24791 2176 24818
rect 2239 24791 2244 24818
rect 1870 24784 1904 24791
rect 1938 24784 1972 24791
rect 2006 24784 2040 24791
rect 2074 24784 2108 24791
rect 2142 24784 2176 24791
rect 2210 24784 2244 24791
rect 2312 24818 2351 24825
rect 2385 24818 2424 24825
rect 2458 24818 2497 24825
rect 2531 24818 2570 24825
rect 2604 24818 2643 24825
rect 2677 24818 2716 24825
rect 2750 24818 2789 24825
rect 2823 24818 2862 24825
rect 2896 24818 2935 24825
rect 2969 24818 3008 24825
rect 3042 24818 3081 24825
rect 3115 24818 3154 24825
rect 3188 24818 3227 24825
rect 3261 24818 3300 24825
rect 3334 24818 3373 24825
rect 3407 24818 3446 24825
rect 3480 24818 3519 24825
rect 3553 24818 3592 24825
rect 3626 24818 3665 24825
rect 3699 24818 3738 24825
rect 3772 24818 3811 24825
rect 3845 24818 3884 24825
rect 3918 24818 3957 24825
rect 3991 24818 4030 24825
rect 4064 24818 4103 24825
rect 4137 24818 4176 24825
rect 4210 24818 4249 24825
rect 4283 24818 4322 24825
rect 4356 24818 4395 24825
rect 4429 24818 4468 24825
rect 2278 24784 2312 24791
rect 2346 24791 2351 24818
rect 2414 24791 2424 24818
rect 2482 24791 2497 24818
rect 2550 24791 2570 24818
rect 2618 24791 2643 24818
rect 2686 24791 2716 24818
rect 2346 24784 2380 24791
rect 2414 24784 2448 24791
rect 2482 24784 2516 24791
rect 2550 24784 2584 24791
rect 2618 24784 2652 24791
rect 2686 24784 2720 24791
rect 2754 24784 2788 24818
rect 2823 24791 2856 24818
rect 2896 24791 2924 24818
rect 2969 24791 2992 24818
rect 3042 24791 3060 24818
rect 3115 24791 3128 24818
rect 3188 24791 3196 24818
rect 3261 24791 3264 24818
rect 2822 24784 2856 24791
rect 2890 24784 2924 24791
rect 2958 24784 2992 24791
rect 3026 24784 3060 24791
rect 3094 24784 3128 24791
rect 3162 24784 3196 24791
rect 3230 24784 3264 24791
rect 3298 24791 3300 24818
rect 3366 24791 3373 24818
rect 3434 24791 3446 24818
rect 3502 24791 3519 24818
rect 3570 24791 3592 24818
rect 3638 24791 3665 24818
rect 3706 24791 3738 24818
rect 3298 24784 3332 24791
rect 3366 24784 3400 24791
rect 3434 24784 3468 24791
rect 3502 24784 3536 24791
rect 3570 24784 3604 24791
rect 3638 24784 3672 24791
rect 3706 24784 3740 24791
rect 3774 24784 3808 24818
rect 3845 24791 3876 24818
rect 3918 24791 3944 24818
rect 3991 24791 4012 24818
rect 4064 24791 4080 24818
rect 4137 24791 4148 24818
rect 4210 24791 4216 24818
rect 4283 24791 4284 24818
rect 3842 24784 3876 24791
rect 3910 24784 3944 24791
rect 3978 24784 4012 24791
rect 4046 24784 4080 24791
rect 4114 24784 4148 24791
rect 4182 24784 4216 24791
rect 4250 24784 4284 24791
rect 4318 24791 4322 24818
rect 4386 24791 4395 24818
rect 4318 24784 4352 24791
rect 4386 24784 4420 24791
rect 4454 24784 4468 24818
rect -41 24753 4468 24784
rect -41 24719 88 24753
rect 122 24746 161 24753
rect 195 24746 234 24753
rect 268 24746 307 24753
rect 341 24746 380 24753
rect 414 24746 453 24753
rect 487 24746 526 24753
rect 560 24746 599 24753
rect 633 24746 672 24753
rect 706 24746 745 24753
rect 779 24746 818 24753
rect 852 24746 891 24753
rect 925 24746 964 24753
rect 998 24746 1037 24753
rect 1071 24746 1110 24753
rect 1144 24746 1183 24753
rect 1217 24746 1256 24753
rect 1290 24746 1329 24753
rect 1363 24746 1402 24753
rect 1436 24746 1475 24753
rect 1509 24746 1548 24753
rect 1582 24746 1621 24753
rect 1655 24746 1694 24753
rect 1728 24746 1767 24753
rect 1801 24746 1840 24753
rect 1874 24746 1913 24753
rect 1947 24746 1986 24753
rect 2020 24746 2059 24753
rect 2093 24746 2132 24753
rect 2166 24746 2205 24753
rect 2239 24746 2278 24753
rect 122 24719 124 24746
rect -41 24712 124 24719
rect 158 24719 161 24746
rect 227 24719 234 24746
rect 296 24719 307 24746
rect 365 24719 380 24746
rect 434 24719 453 24746
rect 503 24719 526 24746
rect 572 24719 599 24746
rect 641 24719 672 24746
rect 158 24712 193 24719
rect 227 24712 262 24719
rect 296 24712 331 24719
rect 365 24712 400 24719
rect 434 24712 469 24719
rect 503 24712 538 24719
rect 572 24712 607 24719
rect 641 24712 676 24719
rect 710 24712 745 24746
rect 779 24712 814 24746
rect 852 24719 883 24746
rect 925 24719 952 24746
rect 998 24719 1020 24746
rect 1071 24719 1088 24746
rect 1144 24719 1156 24746
rect 1217 24719 1224 24746
rect 1290 24719 1292 24746
rect 848 24712 883 24719
rect 917 24712 952 24719
rect 986 24712 1020 24719
rect 1054 24712 1088 24719
rect 1122 24712 1156 24719
rect 1190 24712 1224 24719
rect 1258 24712 1292 24719
rect 1326 24719 1329 24746
rect 1394 24719 1402 24746
rect 1462 24719 1475 24746
rect 1530 24719 1548 24746
rect 1598 24719 1621 24746
rect 1666 24719 1694 24746
rect 1734 24719 1767 24746
rect 1326 24712 1360 24719
rect 1394 24712 1428 24719
rect 1462 24712 1496 24719
rect 1530 24712 1564 24719
rect 1598 24712 1632 24719
rect 1666 24712 1700 24719
rect 1734 24712 1768 24719
rect 1802 24712 1836 24746
rect 1874 24719 1904 24746
rect 1947 24719 1972 24746
rect 2020 24719 2040 24746
rect 2093 24719 2108 24746
rect 2166 24719 2176 24746
rect 2239 24719 2244 24746
rect 1870 24712 1904 24719
rect 1938 24712 1972 24719
rect 2006 24712 2040 24719
rect 2074 24712 2108 24719
rect 2142 24712 2176 24719
rect 2210 24712 2244 24719
rect 2312 24746 2351 24753
rect 2385 24746 2424 24753
rect 2458 24746 2497 24753
rect 2531 24746 2570 24753
rect 2604 24746 2643 24753
rect 2677 24746 2716 24753
rect 2750 24746 2789 24753
rect 2823 24746 2862 24753
rect 2896 24746 2935 24753
rect 2969 24746 3008 24753
rect 3042 24746 3081 24753
rect 3115 24746 3154 24753
rect 3188 24746 3227 24753
rect 3261 24746 3300 24753
rect 3334 24746 3373 24753
rect 3407 24746 3446 24753
rect 3480 24746 3519 24753
rect 3553 24746 3592 24753
rect 3626 24746 3665 24753
rect 3699 24746 3738 24753
rect 3772 24746 3811 24753
rect 3845 24746 3884 24753
rect 3918 24746 3957 24753
rect 3991 24746 4030 24753
rect 4064 24746 4103 24753
rect 4137 24746 4176 24753
rect 4210 24746 4249 24753
rect 4283 24746 4322 24753
rect 4356 24746 4395 24753
rect 4429 24746 4468 24753
rect 2278 24712 2312 24719
rect 2346 24719 2351 24746
rect 2414 24719 2424 24746
rect 2482 24719 2497 24746
rect 2550 24719 2570 24746
rect 2618 24719 2643 24746
rect 2686 24719 2716 24746
rect 2346 24712 2380 24719
rect 2414 24712 2448 24719
rect 2482 24712 2516 24719
rect 2550 24712 2584 24719
rect 2618 24712 2652 24719
rect 2686 24712 2720 24719
rect 2754 24712 2788 24746
rect 2823 24719 2856 24746
rect 2896 24719 2924 24746
rect 2969 24719 2992 24746
rect 3042 24719 3060 24746
rect 3115 24719 3128 24746
rect 3188 24719 3196 24746
rect 3261 24719 3264 24746
rect 2822 24712 2856 24719
rect 2890 24712 2924 24719
rect 2958 24712 2992 24719
rect 3026 24712 3060 24719
rect 3094 24712 3128 24719
rect 3162 24712 3196 24719
rect 3230 24712 3264 24719
rect 3298 24719 3300 24746
rect 3366 24719 3373 24746
rect 3434 24719 3446 24746
rect 3502 24719 3519 24746
rect 3570 24719 3592 24746
rect 3638 24719 3665 24746
rect 3706 24719 3738 24746
rect 3298 24712 3332 24719
rect 3366 24712 3400 24719
rect 3434 24712 3468 24719
rect 3502 24712 3536 24719
rect 3570 24712 3604 24719
rect 3638 24712 3672 24719
rect 3706 24712 3740 24719
rect 3774 24712 3808 24746
rect 3845 24719 3876 24746
rect 3918 24719 3944 24746
rect 3991 24719 4012 24746
rect 4064 24719 4080 24746
rect 4137 24719 4148 24746
rect 4210 24719 4216 24746
rect 4283 24719 4284 24746
rect 3842 24712 3876 24719
rect 3910 24712 3944 24719
rect 3978 24712 4012 24719
rect 4046 24712 4080 24719
rect 4114 24712 4148 24719
rect 4182 24712 4216 24719
rect 4250 24712 4284 24719
rect 4318 24719 4322 24746
rect 4386 24719 4395 24746
rect 4454 24719 4468 24746
rect 14870 24719 14983 25041
rect 4318 24712 4352 24719
rect 4386 24712 4420 24719
rect 4454 24712 4488 24719
rect 4522 24712 4556 24719
rect 4590 24712 4624 24719
rect 4658 24712 4692 24719
rect 4726 24712 4760 24719
rect 4794 24712 4828 24719
rect 4862 24712 4896 24719
rect 4930 24712 4964 24719
rect 4998 24712 5032 24719
rect 5066 24712 5100 24719
rect 5134 24712 5168 24719
rect 5202 24712 5236 24719
rect 5270 24712 5304 24719
rect 5338 24712 5372 24719
rect 5406 24712 5440 24719
rect 5474 24712 5508 24719
rect 5542 24712 5576 24719
rect 5610 24712 5644 24719
rect 5678 24712 5712 24719
rect 5746 24712 5780 24719
rect 5814 24712 5848 24719
rect 5882 24712 5916 24719
rect 5950 24712 5984 24719
rect 6018 24712 6052 24719
rect 6086 24712 6120 24719
rect 6154 24712 6188 24719
rect 6222 24712 6256 24719
rect 6290 24712 6324 24719
rect 6358 24712 6392 24719
rect 6426 24712 6460 24719
rect 6494 24712 6528 24719
rect 6562 24712 6596 24719
rect 6630 24712 6664 24719
rect 6698 24712 6732 24719
rect 6766 24712 6800 24719
rect 6834 24712 6868 24719
rect 6902 24712 6936 24719
rect 6970 24712 7004 24719
rect 7038 24712 7072 24719
rect 7106 24712 7140 24719
rect 7174 24712 7208 24719
rect 7242 24712 7276 24719
rect 7310 24712 7344 24719
rect 7378 24712 7412 24719
rect 7446 24712 7480 24719
rect 7514 24712 7548 24719
rect 7582 24712 7616 24719
rect 7650 24712 7684 24719
rect 7718 24712 7752 24719
rect 7786 24712 7820 24719
rect 7854 24712 7888 24719
rect 7922 24712 7956 24719
rect 7990 24712 8024 24719
rect 8058 24712 8092 24719
rect 8126 24712 8160 24719
rect 8194 24712 8228 24719
rect 8262 24712 8296 24719
rect 8330 24712 8364 24719
rect 8398 24712 8432 24719
rect 8466 24712 8500 24719
rect 8534 24712 8568 24719
rect 8602 24712 8636 24719
rect 8670 24712 8704 24719
rect 8738 24712 8772 24719
rect 8806 24712 8840 24719
rect 8874 24712 8908 24719
rect 8942 24712 8976 24719
rect 9010 24712 9044 24719
rect 9078 24712 9112 24719
rect 9146 24712 9180 24719
rect 9214 24712 9248 24719
rect 9282 24712 9316 24719
rect 9350 24712 9384 24719
rect 9418 24712 9452 24719
rect 9486 24712 9520 24719
rect 9554 24712 9588 24719
rect 9622 24712 9656 24719
rect 9690 24712 9724 24719
rect 9758 24712 9792 24719
rect 9826 24712 9860 24719
rect 9894 24712 9928 24719
rect 9962 24712 9996 24719
rect 10030 24712 10064 24719
rect 10098 24712 10132 24719
rect 10166 24712 10200 24719
rect 10234 24712 10268 24719
rect 10302 24712 10336 24719
rect 10370 24712 10404 24719
rect 10438 24712 10472 24719
rect 10506 24712 10540 24719
rect 10574 24712 10608 24719
rect 10642 24712 10676 24719
rect 10710 24712 10744 24719
rect 10778 24712 10812 24719
rect 10846 24712 10880 24719
rect 10914 24712 10948 24719
rect 10982 24712 11016 24719
rect 11050 24712 11084 24719
rect 11118 24712 11152 24719
rect 11186 24712 11220 24719
rect 11254 24712 11288 24719
rect 11322 24712 11356 24719
rect 11390 24712 11424 24719
rect 11458 24712 11492 24719
rect 11526 24712 11560 24719
rect 11594 24712 11628 24719
rect 11662 24712 11696 24719
rect 11730 24712 11764 24719
rect 11798 24712 11832 24719
rect 11866 24712 11900 24719
rect 11934 24712 11968 24719
rect 12002 24712 12036 24719
rect 12070 24712 12104 24719
rect 12138 24712 12172 24719
rect 12206 24712 12240 24719
rect 12274 24712 12308 24719
rect 12342 24712 12376 24719
rect 12410 24712 12444 24719
rect 12478 24712 12512 24719
rect 12546 24712 12580 24719
rect 12614 24712 12648 24719
rect 12682 24712 12716 24719
rect 12750 24712 12784 24719
rect 12818 24712 12852 24719
rect 12886 24712 12920 24719
rect 12954 24712 12988 24719
rect 13022 24712 13056 24719
rect 13090 24712 13124 24719
rect 13158 24712 13192 24719
rect 13226 24712 13260 24719
rect 13294 24712 13328 24719
rect 13362 24712 13396 24719
rect 13430 24712 13464 24719
rect 13498 24712 13532 24719
rect 13566 24712 13600 24719
rect 13634 24712 13668 24719
rect 13702 24712 13736 24719
rect 13770 24712 13804 24719
rect 13838 24712 13872 24719
rect 13906 24712 13940 24719
rect 13974 24712 14008 24719
rect 14042 24712 14076 24719
rect 14110 24712 14144 24719
rect 14178 24712 14212 24719
rect 14246 24712 14280 24719
rect 14314 24712 14348 24719
rect 14382 24712 14416 24719
rect 14450 24712 14484 24719
rect 14518 24712 14552 24719
rect 14586 24712 14620 24719
rect 14654 24712 14688 24719
rect 14722 24712 14756 24719
rect 14790 24712 14824 24719
rect 14858 24712 14983 24719
rect -41 24648 14983 24712
rect 53 19884 261 24648
rect 12408 24523 14983 24648
rect -17 19879 6960 19884
rect 14739 19879 14983 24523
rect -41 19859 14983 19879
rect -41 19858 77 19859
rect 111 19858 146 19859
rect -41 19824 70 19858
rect 111 19825 143 19858
rect 180 19825 215 19859
rect 249 19858 284 19859
rect 318 19858 353 19859
rect 387 19858 422 19859
rect 456 19858 491 19859
rect 525 19858 560 19859
rect 594 19858 629 19859
rect 663 19858 698 19859
rect 732 19858 767 19859
rect 801 19858 836 19859
rect 250 19825 284 19858
rect 323 19825 353 19858
rect 396 19825 422 19858
rect 469 19825 491 19858
rect 542 19825 560 19858
rect 615 19825 629 19858
rect 688 19825 698 19858
rect 761 19825 767 19858
rect 834 19825 836 19858
rect 870 19858 905 19859
rect 939 19858 974 19859
rect 1008 19858 1043 19859
rect 1077 19858 1112 19859
rect 1146 19858 1181 19859
rect 1215 19858 1250 19859
rect 1284 19858 1319 19859
rect 1353 19858 1388 19859
rect 870 19825 873 19858
rect 939 19825 946 19858
rect 1008 19825 1019 19858
rect 1077 19825 1092 19858
rect 1146 19825 1165 19858
rect 1215 19825 1238 19858
rect 1284 19825 1311 19858
rect 1353 19825 1384 19858
rect 1422 19825 1457 19859
rect 1491 19825 1526 19859
rect 1560 19858 1595 19859
rect 1629 19858 1664 19859
rect 1698 19858 1733 19859
rect 1767 19858 1802 19859
rect 1836 19858 1871 19859
rect 1905 19858 1940 19859
rect 1974 19858 2009 19859
rect 2043 19858 2078 19859
rect 1564 19825 1595 19858
rect 1637 19825 1664 19858
rect 1710 19825 1733 19858
rect 1783 19825 1802 19858
rect 1856 19825 1871 19858
rect 1929 19825 1940 19858
rect 2002 19825 2009 19858
rect 2075 19825 2078 19858
rect 2112 19858 2147 19859
rect 2181 19858 2216 19859
rect 2250 19858 2285 19859
rect 2319 19858 2354 19859
rect 2388 19858 2423 19859
rect 2457 19858 2492 19859
rect 2526 19858 2561 19859
rect 2595 19858 2630 19859
rect 2664 19858 2699 19859
rect 2112 19825 2114 19858
rect 2181 19825 2187 19858
rect 2250 19825 2260 19858
rect 2319 19825 2333 19858
rect 2388 19825 2406 19858
rect 2457 19825 2479 19858
rect 2526 19825 2552 19858
rect 2595 19825 2625 19858
rect 2664 19825 2698 19858
rect 2733 19825 2768 19859
rect 2802 19858 2837 19859
rect 2871 19858 2906 19859
rect 2940 19858 2975 19859
rect 3009 19858 3044 19859
rect 3078 19858 3113 19859
rect 3147 19858 3182 19859
rect 14436 19858 14983 19859
rect 2805 19825 2837 19858
rect 2878 19825 2906 19858
rect 2951 19825 2975 19858
rect 3024 19825 3044 19858
rect 3097 19825 3113 19858
rect 104 19824 143 19825
rect 177 19824 216 19825
rect 250 19824 289 19825
rect 323 19824 362 19825
rect 396 19824 435 19825
rect 469 19824 508 19825
rect 542 19824 581 19825
rect 615 19824 654 19825
rect 688 19824 727 19825
rect 761 19824 800 19825
rect 834 19824 873 19825
rect 907 19824 946 19825
rect 980 19824 1019 19825
rect 1053 19824 1092 19825
rect 1126 19824 1165 19825
rect 1199 19824 1238 19825
rect 1272 19824 1311 19825
rect 1345 19824 1384 19825
rect 1418 19824 1457 19825
rect 1491 19824 1530 19825
rect 1564 19824 1603 19825
rect 1637 19824 1676 19825
rect 1710 19824 1749 19825
rect 1783 19824 1822 19825
rect 1856 19824 1895 19825
rect 1929 19824 1968 19825
rect 2002 19824 2041 19825
rect 2075 19824 2114 19825
rect 2148 19824 2187 19825
rect 2221 19824 2260 19825
rect 2294 19824 2333 19825
rect 2367 19824 2406 19825
rect 2440 19824 2479 19825
rect 2513 19824 2552 19825
rect 2586 19824 2625 19825
rect 2659 19824 2698 19825
rect 2732 19824 2771 19825
rect 2805 19824 2844 19825
rect 2878 19824 2917 19825
rect 2951 19824 2990 19825
rect 3024 19824 3063 19825
rect 3097 19824 3136 19825
rect 3170 19824 3182 19858
rect 14436 19824 14442 19858
rect 14476 19831 14514 19858
rect 14548 19831 14586 19858
rect 14620 19831 14658 19858
rect 14476 19824 14484 19831
rect 14548 19824 14567 19831
rect 14620 19824 14650 19831
rect 14692 19824 14730 19858
rect 14764 19831 14802 19858
rect 14836 19831 14874 19858
rect 14767 19824 14802 19831
rect 14850 19824 14874 19831
rect 14908 19839 14983 19858
rect 14908 19824 14959 19839
rect -41 19791 3182 19824
rect -41 19772 77 19791
rect 111 19772 146 19791
rect -41 19738 70 19772
rect 111 19757 143 19772
rect 180 19757 215 19791
rect 249 19772 284 19791
rect 318 19772 353 19791
rect 387 19772 422 19791
rect 456 19772 491 19791
rect 525 19772 560 19791
rect 594 19772 629 19791
rect 663 19772 698 19791
rect 732 19772 767 19791
rect 801 19772 836 19791
rect 250 19757 284 19772
rect 323 19757 353 19772
rect 396 19757 422 19772
rect 469 19757 491 19772
rect 542 19757 560 19772
rect 615 19757 629 19772
rect 688 19757 698 19772
rect 761 19757 767 19772
rect 834 19757 836 19772
rect 870 19772 905 19791
rect 939 19772 974 19791
rect 1008 19772 1043 19791
rect 1077 19772 1112 19791
rect 1146 19772 1181 19791
rect 1215 19772 1250 19791
rect 1284 19772 1319 19791
rect 1353 19772 1388 19791
rect 870 19757 873 19772
rect 939 19757 946 19772
rect 1008 19757 1019 19772
rect 1077 19757 1092 19772
rect 1146 19757 1165 19772
rect 1215 19757 1238 19772
rect 1284 19757 1311 19772
rect 1353 19757 1384 19772
rect 1422 19757 1457 19791
rect 1491 19757 1526 19791
rect 1560 19772 1595 19791
rect 1629 19772 1664 19791
rect 1698 19772 1733 19791
rect 1767 19772 1802 19791
rect 1836 19772 1871 19791
rect 1905 19772 1940 19791
rect 1974 19772 2009 19791
rect 2043 19772 2078 19791
rect 1564 19757 1595 19772
rect 1637 19757 1664 19772
rect 1710 19757 1733 19772
rect 1783 19757 1802 19772
rect 1856 19757 1871 19772
rect 1929 19757 1940 19772
rect 2002 19757 2009 19772
rect 2075 19757 2078 19772
rect 2112 19772 2147 19791
rect 2181 19772 2216 19791
rect 2250 19772 2285 19791
rect 2319 19772 2354 19791
rect 2388 19772 2423 19791
rect 2457 19772 2492 19791
rect 2526 19772 2561 19791
rect 2595 19772 2630 19791
rect 2664 19772 2699 19791
rect 2112 19757 2114 19772
rect 2181 19757 2187 19772
rect 2250 19757 2260 19772
rect 2319 19757 2333 19772
rect 2388 19757 2406 19772
rect 2457 19757 2479 19772
rect 2526 19757 2552 19772
rect 2595 19757 2625 19772
rect 2664 19757 2698 19772
rect 2733 19757 2768 19791
rect 2802 19772 2837 19791
rect 2871 19772 2906 19791
rect 2940 19772 2975 19791
rect 3009 19772 3044 19791
rect 3078 19772 3113 19791
rect 3147 19772 3182 19791
rect 14436 19797 14484 19824
rect 14518 19797 14567 19824
rect 14601 19797 14650 19824
rect 14684 19797 14733 19824
rect 14767 19797 14816 19824
rect 14850 19797 14959 19824
rect 14436 19772 14959 19797
rect 2805 19757 2837 19772
rect 2878 19757 2906 19772
rect 2951 19757 2975 19772
rect 3024 19757 3044 19772
rect 3097 19757 3113 19772
rect 104 19738 143 19757
rect 177 19738 216 19757
rect 250 19738 289 19757
rect 323 19738 362 19757
rect 396 19738 435 19757
rect 469 19738 508 19757
rect 542 19738 581 19757
rect 615 19738 654 19757
rect 688 19738 727 19757
rect 761 19738 800 19757
rect 834 19738 873 19757
rect 907 19738 946 19757
rect 980 19738 1019 19757
rect 1053 19738 1092 19757
rect 1126 19738 1165 19757
rect 1199 19738 1238 19757
rect 1272 19738 1311 19757
rect 1345 19738 1384 19757
rect 1418 19738 1457 19757
rect 1491 19738 1530 19757
rect 1564 19738 1603 19757
rect 1637 19738 1676 19757
rect 1710 19738 1749 19757
rect 1783 19738 1822 19757
rect 1856 19738 1895 19757
rect 1929 19738 1968 19757
rect 2002 19738 2041 19757
rect 2075 19738 2114 19757
rect 2148 19738 2187 19757
rect 2221 19738 2260 19757
rect 2294 19738 2333 19757
rect 2367 19738 2406 19757
rect 2440 19738 2479 19757
rect 2513 19738 2552 19757
rect 2586 19738 2625 19757
rect 2659 19738 2698 19757
rect 2732 19738 2771 19757
rect 2805 19738 2844 19757
rect 2878 19738 2917 19757
rect 2951 19738 2990 19757
rect 3024 19738 3063 19757
rect 3097 19738 3136 19757
rect 3170 19738 3182 19772
rect 14436 19738 14442 19772
rect 14476 19761 14514 19772
rect 14548 19761 14586 19772
rect 14620 19761 14658 19772
rect 14476 19738 14484 19761
rect 14548 19738 14567 19761
rect 14620 19738 14650 19761
rect 14692 19738 14730 19772
rect 14764 19761 14802 19772
rect 14836 19761 14874 19772
rect 14767 19738 14802 19761
rect 14850 19738 14874 19761
rect 14908 19738 14959 19772
rect -41 19723 3182 19738
rect -41 19689 77 19723
rect 111 19689 146 19723
rect 180 19689 215 19723
rect 249 19689 284 19723
rect 318 19689 353 19723
rect 387 19689 422 19723
rect 456 19689 491 19723
rect 525 19689 560 19723
rect 594 19689 629 19723
rect 663 19689 698 19723
rect 732 19689 767 19723
rect 801 19689 836 19723
rect 870 19689 905 19723
rect 939 19689 974 19723
rect 1008 19689 1043 19723
rect 1077 19689 1112 19723
rect 1146 19689 1181 19723
rect 1215 19689 1250 19723
rect 1284 19689 1319 19723
rect 1353 19689 1388 19723
rect 1422 19689 1457 19723
rect 1491 19689 1526 19723
rect 1560 19689 1595 19723
rect 1629 19689 1664 19723
rect 1698 19689 1733 19723
rect 1767 19689 1802 19723
rect 1836 19689 1871 19723
rect 1905 19689 1940 19723
rect 1974 19689 2009 19723
rect 2043 19689 2078 19723
rect 2112 19689 2147 19723
rect 2181 19689 2216 19723
rect 2250 19689 2285 19723
rect 2319 19689 2354 19723
rect 2388 19689 2423 19723
rect 2457 19689 2492 19723
rect 2526 19689 2561 19723
rect 2595 19689 2630 19723
rect 2664 19689 2699 19723
rect 2733 19689 2768 19723
rect 2802 19689 2837 19723
rect 2871 19689 2906 19723
rect 2940 19689 2975 19723
rect 3009 19689 3044 19723
rect 3078 19689 3113 19723
rect 3147 19689 3182 19723
rect -41 19686 3182 19689
rect 14436 19727 14484 19738
rect 14518 19727 14567 19738
rect 14601 19727 14650 19738
rect 14684 19727 14733 19738
rect 14767 19727 14816 19738
rect 14850 19727 14959 19738
rect 14436 19691 14959 19727
rect 14436 19686 14484 19691
rect 14518 19686 14567 19691
rect 14601 19686 14650 19691
rect 14684 19686 14733 19691
rect 14767 19686 14816 19691
rect 14850 19686 14959 19691
rect -41 19652 70 19686
rect 104 19655 143 19686
rect 177 19655 216 19686
rect 250 19655 289 19686
rect 323 19655 362 19686
rect 396 19655 435 19686
rect 469 19655 508 19686
rect 542 19655 581 19686
rect 615 19655 654 19686
rect 688 19655 727 19686
rect 761 19655 800 19686
rect 834 19655 873 19686
rect 907 19655 946 19686
rect 980 19655 1019 19686
rect 1053 19655 1092 19686
rect 1126 19655 1165 19686
rect 1199 19655 1238 19686
rect 1272 19655 1311 19686
rect 1345 19655 1384 19686
rect 1418 19655 1457 19686
rect 1491 19655 1530 19686
rect 1564 19655 1603 19686
rect 1637 19655 1676 19686
rect 1710 19655 1749 19686
rect 1783 19655 1822 19686
rect 1856 19655 1895 19686
rect 1929 19655 1968 19686
rect 2002 19655 2041 19686
rect 2075 19655 2114 19686
rect 2148 19655 2187 19686
rect 2221 19655 2260 19686
rect 2294 19655 2333 19686
rect 2367 19655 2406 19686
rect 2440 19655 2479 19686
rect 2513 19655 2552 19686
rect 2586 19655 2625 19686
rect 2659 19655 2698 19686
rect 2732 19655 2771 19686
rect 2805 19655 2844 19686
rect 2878 19655 2917 19686
rect 2951 19655 2990 19686
rect 3024 19655 3063 19686
rect 3097 19655 3136 19686
rect 111 19652 143 19655
rect -41 19621 77 19652
rect 111 19621 146 19652
rect 180 19621 215 19655
rect 250 19652 284 19655
rect 323 19652 353 19655
rect 396 19652 422 19655
rect 469 19652 491 19655
rect 542 19652 560 19655
rect 615 19652 629 19655
rect 688 19652 698 19655
rect 761 19652 767 19655
rect 834 19652 836 19655
rect 249 19621 284 19652
rect 318 19621 353 19652
rect 387 19621 422 19652
rect 456 19621 491 19652
rect 525 19621 560 19652
rect 594 19621 629 19652
rect 663 19621 698 19652
rect 732 19621 767 19652
rect 801 19621 836 19652
rect 870 19652 873 19655
rect 939 19652 946 19655
rect 1008 19652 1019 19655
rect 1077 19652 1092 19655
rect 1146 19652 1165 19655
rect 1215 19652 1238 19655
rect 1284 19652 1311 19655
rect 1353 19652 1384 19655
rect 870 19621 905 19652
rect 939 19621 974 19652
rect 1008 19621 1043 19652
rect 1077 19621 1112 19652
rect 1146 19621 1181 19652
rect 1215 19621 1250 19652
rect 1284 19621 1319 19652
rect 1353 19621 1388 19652
rect 1422 19621 1457 19655
rect 1491 19621 1526 19655
rect 1564 19652 1595 19655
rect 1637 19652 1664 19655
rect 1710 19652 1733 19655
rect 1783 19652 1802 19655
rect 1856 19652 1871 19655
rect 1929 19652 1940 19655
rect 2002 19652 2009 19655
rect 2075 19652 2078 19655
rect 1560 19621 1595 19652
rect 1629 19621 1664 19652
rect 1698 19621 1733 19652
rect 1767 19621 1802 19652
rect 1836 19621 1871 19652
rect 1905 19621 1940 19652
rect 1974 19621 2009 19652
rect 2043 19621 2078 19652
rect 2112 19652 2114 19655
rect 2181 19652 2187 19655
rect 2250 19652 2260 19655
rect 2319 19652 2333 19655
rect 2388 19652 2406 19655
rect 2457 19652 2479 19655
rect 2526 19652 2552 19655
rect 2595 19652 2625 19655
rect 2664 19652 2698 19655
rect 2112 19621 2147 19652
rect 2181 19621 2216 19652
rect 2250 19621 2285 19652
rect 2319 19621 2354 19652
rect 2388 19621 2423 19652
rect 2457 19621 2492 19652
rect 2526 19621 2561 19652
rect 2595 19621 2630 19652
rect 2664 19621 2699 19652
rect 2733 19621 2768 19655
rect 2805 19652 2837 19655
rect 2878 19652 2906 19655
rect 2951 19652 2975 19655
rect 3024 19652 3044 19655
rect 3097 19652 3113 19655
rect 3170 19652 3182 19686
rect 14436 19652 14442 19686
rect 14476 19657 14484 19686
rect 14548 19657 14567 19686
rect 14620 19657 14650 19686
rect 14476 19652 14514 19657
rect 14548 19652 14586 19657
rect 14620 19652 14658 19657
rect 14692 19652 14730 19686
rect 14767 19657 14802 19686
rect 14850 19657 14874 19686
rect 14764 19652 14802 19657
rect 14836 19652 14874 19657
rect 14908 19652 14959 19686
rect 2802 19621 2837 19652
rect 2871 19621 2906 19652
rect 2940 19621 2975 19652
rect 3009 19621 3044 19652
rect 3078 19621 3113 19652
rect 3147 19621 3182 19652
rect 14436 19621 14959 19652
rect -41 19600 14484 19621
rect 14518 19600 14567 19621
rect 14601 19600 14650 19621
rect 14684 19600 14733 19621
rect 14767 19600 14816 19621
rect 14850 19600 14959 19621
rect -41 19566 70 19600
rect 104 19585 143 19600
rect 177 19585 216 19600
rect 250 19585 289 19600
rect 323 19585 362 19600
rect 396 19585 435 19600
rect 469 19585 508 19600
rect 542 19585 581 19600
rect 615 19585 654 19600
rect 688 19585 727 19600
rect 761 19585 800 19600
rect 834 19585 873 19600
rect 907 19585 946 19600
rect 980 19585 1019 19600
rect 1053 19585 1092 19600
rect 1126 19585 1165 19600
rect 1199 19585 1238 19600
rect 1272 19585 1311 19600
rect 1345 19585 1384 19600
rect 1418 19585 1457 19600
rect 1491 19585 1530 19600
rect 1564 19585 1603 19600
rect 1637 19585 1676 19600
rect 1710 19585 1749 19600
rect 1783 19585 1822 19600
rect 1856 19585 1895 19600
rect 1929 19585 1968 19600
rect 2002 19585 2041 19600
rect 2075 19585 2114 19600
rect 2148 19585 2187 19600
rect 2221 19585 2260 19600
rect 2294 19585 2333 19600
rect 2367 19585 2406 19600
rect 2440 19585 2479 19600
rect 2513 19585 2552 19600
rect 2586 19585 2625 19600
rect 2659 19585 2698 19600
rect 2732 19585 2771 19600
rect 2805 19585 2844 19600
rect 2878 19585 2917 19600
rect 2951 19585 2990 19600
rect 3024 19585 3063 19600
rect 3097 19585 3136 19600
rect 3170 19585 3209 19600
rect 3243 19585 3282 19600
rect 3316 19585 3354 19600
rect 111 19566 143 19585
rect -41 19551 77 19566
rect 111 19551 146 19566
rect 180 19551 215 19585
rect 250 19566 284 19585
rect 323 19566 353 19585
rect 396 19566 422 19585
rect 469 19566 491 19585
rect 542 19566 560 19585
rect 615 19566 629 19585
rect 688 19566 698 19585
rect 761 19566 767 19585
rect 834 19566 836 19585
rect 249 19551 284 19566
rect 318 19551 353 19566
rect 387 19551 422 19566
rect 456 19551 491 19566
rect 525 19551 560 19566
rect 594 19551 629 19566
rect 663 19551 698 19566
rect 732 19551 767 19566
rect 801 19551 836 19566
rect 870 19566 873 19585
rect 939 19566 946 19585
rect 1008 19566 1019 19585
rect 1077 19566 1092 19585
rect 1146 19566 1165 19585
rect 1215 19566 1238 19585
rect 1284 19566 1311 19585
rect 1353 19566 1384 19585
rect 870 19551 905 19566
rect 939 19551 974 19566
rect 1008 19551 1043 19566
rect 1077 19551 1112 19566
rect 1146 19551 1181 19566
rect 1215 19551 1250 19566
rect 1284 19551 1319 19566
rect 1353 19551 1388 19566
rect 1422 19551 1457 19585
rect 1491 19551 1526 19585
rect 1564 19566 1595 19585
rect 1637 19566 1664 19585
rect 1710 19566 1733 19585
rect 1783 19566 1802 19585
rect 1856 19566 1871 19585
rect 1929 19566 1940 19585
rect 2002 19566 2009 19585
rect 2075 19566 2078 19585
rect 1560 19551 1595 19566
rect 1629 19551 1664 19566
rect 1698 19551 1733 19566
rect 1767 19551 1802 19566
rect 1836 19551 1871 19566
rect 1905 19551 1940 19566
rect 1974 19551 2009 19566
rect 2043 19551 2078 19566
rect 2112 19566 2114 19585
rect 2181 19566 2187 19585
rect 2250 19566 2260 19585
rect 2319 19566 2333 19585
rect 2388 19566 2406 19585
rect 2457 19566 2479 19585
rect 2526 19566 2552 19585
rect 2595 19566 2625 19585
rect 2664 19566 2698 19585
rect 2112 19551 2147 19566
rect 2181 19551 2216 19566
rect 2250 19551 2285 19566
rect 2319 19551 2354 19566
rect 2388 19551 2423 19566
rect 2457 19551 2492 19566
rect 2526 19551 2561 19566
rect 2595 19551 2630 19566
rect 2664 19551 2699 19566
rect 2733 19551 2768 19585
rect 2805 19566 2837 19585
rect 2878 19566 2906 19585
rect 2951 19566 2975 19585
rect 3024 19566 3044 19585
rect 3097 19566 3113 19585
rect 3170 19566 3182 19585
rect 3243 19566 3251 19585
rect 3316 19566 3320 19585
rect 2802 19551 2837 19566
rect 2871 19551 2906 19566
rect 2940 19551 2975 19566
rect 3009 19551 3044 19566
rect 3078 19551 3113 19566
rect 3147 19551 3182 19566
rect 3216 19551 3251 19566
rect 3285 19551 3320 19566
rect 3388 19585 3426 19600
rect 3460 19585 3498 19600
rect 3532 19585 3570 19600
rect 3604 19585 3642 19600
rect 3676 19585 3714 19600
rect 3748 19585 3786 19600
rect 3820 19585 3858 19600
rect 3892 19585 3930 19600
rect 3964 19585 4002 19600
rect 4036 19585 4074 19600
rect 4108 19585 4146 19600
rect 4180 19585 4218 19600
rect 4252 19585 4290 19600
rect 4324 19585 4362 19600
rect 4396 19585 4434 19600
rect 4468 19585 4506 19600
rect 4540 19585 4578 19600
rect 4612 19585 4650 19600
rect 4684 19585 4722 19600
rect 4756 19585 4794 19600
rect 4828 19585 4866 19600
rect 4900 19585 4938 19600
rect 4972 19585 5010 19600
rect 5044 19585 5082 19600
rect 5116 19585 5154 19600
rect 5188 19585 5226 19600
rect 5260 19585 5298 19600
rect 5332 19585 5370 19600
rect 5404 19585 5442 19600
rect 5476 19585 5514 19600
rect 5548 19585 5586 19600
rect 5620 19585 5658 19600
rect 5692 19585 5730 19600
rect 5764 19585 5802 19600
rect 5836 19585 5874 19600
rect 5908 19585 5946 19600
rect 5980 19585 6018 19600
rect 6052 19585 6090 19600
rect 6124 19585 6162 19600
rect 6196 19585 6234 19600
rect 6268 19585 6306 19600
rect 6340 19585 6378 19600
rect 6412 19585 6450 19600
rect 6484 19585 6522 19600
rect 6556 19585 6594 19600
rect 6628 19585 6666 19600
rect 6700 19585 6738 19600
rect 6772 19585 6810 19600
rect 6844 19585 6882 19600
rect 6916 19585 6954 19600
rect 6988 19585 7026 19600
rect 7060 19585 7098 19600
rect 7132 19585 7170 19600
rect 7204 19585 7242 19600
rect 7276 19585 7314 19600
rect 7348 19585 7386 19600
rect 7420 19585 7458 19600
rect 7492 19585 7530 19600
rect 7564 19585 7602 19600
rect 7636 19585 7674 19600
rect 7708 19585 7746 19600
rect 7780 19585 7818 19600
rect 7852 19585 7890 19600
rect 7924 19585 7962 19600
rect 7996 19585 8034 19600
rect 8068 19585 8106 19600
rect 8140 19585 8178 19600
rect 8212 19585 8250 19600
rect 8284 19585 8322 19600
rect 8356 19585 8394 19600
rect 8428 19585 8466 19600
rect 8500 19585 8538 19600
rect 8572 19585 8610 19600
rect 8644 19585 8682 19600
rect 8716 19585 8754 19600
rect 8788 19585 8826 19600
rect 8860 19585 8898 19600
rect 8932 19585 8970 19600
rect 9004 19585 9042 19600
rect 9076 19585 9114 19600
rect 9148 19585 9186 19600
rect 9220 19585 9258 19600
rect 9292 19585 9330 19600
rect 9364 19585 9402 19600
rect 9436 19585 9474 19600
rect 9508 19585 9546 19600
rect 9580 19585 9618 19600
rect 9652 19585 9690 19600
rect 9724 19585 9762 19600
rect 9796 19585 9834 19600
rect 9868 19585 9906 19600
rect 9940 19585 9978 19600
rect 10012 19585 10050 19600
rect 10084 19585 10122 19600
rect 10156 19585 10194 19600
rect 10228 19585 10266 19600
rect 10300 19585 10338 19600
rect 10372 19585 10410 19600
rect 10444 19585 10482 19600
rect 10516 19585 10554 19600
rect 10588 19585 10626 19600
rect 10660 19585 10698 19600
rect 10732 19585 10770 19600
rect 10804 19585 10842 19600
rect 10876 19585 10914 19600
rect 10948 19585 10986 19600
rect 11020 19585 11058 19600
rect 11092 19585 11130 19600
rect 11164 19585 11202 19600
rect 11236 19585 11274 19600
rect 11308 19585 11346 19600
rect 11380 19585 11418 19600
rect 11452 19585 11490 19600
rect 11524 19585 11562 19600
rect 11596 19585 11634 19600
rect 11668 19585 11706 19600
rect 3388 19566 3389 19585
rect 3354 19551 3389 19566
rect 3423 19566 3426 19585
rect 3492 19566 3498 19585
rect 3561 19566 3570 19585
rect 3630 19566 3642 19585
rect 3699 19566 3714 19585
rect 3767 19566 3786 19585
rect 3835 19566 3858 19585
rect 3903 19566 3930 19585
rect 3971 19566 4002 19585
rect 3423 19551 3458 19566
rect 3492 19551 3527 19566
rect 3561 19551 3596 19566
rect 3630 19551 3665 19566
rect 3699 19551 3733 19566
rect 3767 19551 3801 19566
rect 3835 19551 3869 19566
rect 3903 19551 3937 19566
rect 3971 19551 4005 19566
rect 4039 19551 4073 19585
rect 4108 19566 4141 19585
rect 4180 19566 4209 19585
rect 4252 19566 4277 19585
rect 4324 19566 4345 19585
rect 4396 19566 4413 19585
rect 4468 19566 4481 19585
rect 4540 19566 4549 19585
rect 4612 19566 4617 19585
rect 4684 19566 4685 19585
rect 4107 19551 4141 19566
rect 4175 19551 4209 19566
rect 4243 19551 4277 19566
rect 4311 19551 4345 19566
rect 4379 19551 4413 19566
rect 4447 19551 4481 19566
rect 4515 19551 4549 19566
rect 4583 19551 4617 19566
rect 4651 19551 4685 19566
rect 4719 19566 4722 19585
rect 4787 19566 4794 19585
rect 4855 19566 4866 19585
rect 4923 19566 4938 19585
rect 4991 19566 5010 19585
rect 5059 19566 5082 19585
rect 5127 19566 5154 19585
rect 5195 19566 5226 19585
rect 4719 19551 4753 19566
rect 4787 19551 4821 19566
rect 4855 19551 4889 19566
rect 4923 19551 4957 19566
rect 4991 19551 5025 19566
rect 5059 19551 5093 19566
rect 5127 19551 5161 19566
rect 5195 19551 5229 19566
rect 5263 19551 5297 19585
rect 5332 19566 5365 19585
rect 5404 19566 5433 19585
rect 5476 19566 5501 19585
rect 5548 19566 5569 19585
rect 5620 19566 5637 19585
rect 5692 19566 5705 19585
rect 5764 19566 5773 19585
rect 5836 19566 5841 19585
rect 5908 19566 5909 19585
rect 5331 19551 5365 19566
rect 5399 19551 5433 19566
rect 5467 19551 5501 19566
rect 5535 19551 5569 19566
rect 5603 19551 5637 19566
rect 5671 19551 5705 19566
rect 5739 19551 5773 19566
rect 5807 19551 5841 19566
rect 5875 19551 5909 19566
rect 5943 19566 5946 19585
rect 6011 19566 6018 19585
rect 6079 19566 6090 19585
rect 6147 19566 6162 19585
rect 6215 19566 6234 19585
rect 6283 19566 6306 19585
rect 6351 19566 6378 19585
rect 6419 19566 6450 19585
rect 5943 19551 5977 19566
rect 6011 19551 6045 19566
rect 6079 19551 6113 19566
rect 6147 19551 6181 19566
rect 6215 19551 6249 19566
rect 6283 19551 6317 19566
rect 6351 19551 6385 19566
rect 6419 19551 6453 19566
rect 6487 19551 6521 19585
rect 6556 19566 6589 19585
rect 6628 19566 6657 19585
rect 6700 19566 6725 19585
rect 6772 19566 6793 19585
rect 6844 19566 6861 19585
rect 6916 19566 6929 19585
rect 6988 19566 6997 19585
rect 7060 19566 7065 19585
rect 7132 19566 7133 19585
rect 6555 19551 6589 19566
rect 6623 19551 6657 19566
rect 6691 19551 6725 19566
rect 6759 19551 6793 19566
rect 6827 19551 6861 19566
rect 6895 19551 6929 19566
rect 6963 19551 6997 19566
rect 7031 19551 7065 19566
rect 7099 19551 7133 19566
rect 7167 19566 7170 19585
rect 7235 19566 7242 19585
rect 7303 19566 7314 19585
rect 7371 19566 7386 19585
rect 7439 19566 7458 19585
rect 7507 19566 7530 19585
rect 7575 19566 7602 19585
rect 7643 19566 7674 19585
rect 7167 19551 7201 19566
rect 7235 19551 7269 19566
rect 7303 19551 7337 19566
rect 7371 19551 7405 19566
rect 7439 19551 7473 19566
rect 7507 19551 7541 19566
rect 7575 19551 7609 19566
rect 7643 19551 7677 19566
rect 7711 19551 7745 19585
rect 7780 19566 7813 19585
rect 7852 19566 7881 19585
rect 7924 19566 7949 19585
rect 7996 19566 8017 19585
rect 8068 19566 8085 19585
rect 8140 19566 8153 19585
rect 8212 19566 8221 19585
rect 8284 19566 8289 19585
rect 8356 19566 8357 19585
rect 7779 19551 7813 19566
rect 7847 19551 7881 19566
rect 7915 19551 7949 19566
rect 7983 19551 8017 19566
rect 8051 19551 8085 19566
rect 8119 19551 8153 19566
rect 8187 19551 8221 19566
rect 8255 19551 8289 19566
rect 8323 19551 8357 19566
rect 8391 19566 8394 19585
rect 8459 19566 8466 19585
rect 8527 19566 8538 19585
rect 8595 19566 8610 19585
rect 8663 19566 8682 19585
rect 8731 19566 8754 19585
rect 8799 19566 8826 19585
rect 8867 19566 8898 19585
rect 8391 19551 8425 19566
rect 8459 19551 8493 19566
rect 8527 19551 8561 19566
rect 8595 19551 8629 19566
rect 8663 19551 8697 19566
rect 8731 19551 8765 19566
rect 8799 19551 8833 19566
rect 8867 19551 8901 19566
rect 8935 19551 8969 19585
rect 9004 19566 9037 19585
rect 9076 19566 9105 19585
rect 9148 19566 9173 19585
rect 9220 19566 9241 19585
rect 9292 19566 9309 19585
rect 9364 19566 9377 19585
rect 9436 19566 9445 19585
rect 9508 19566 9513 19585
rect 9580 19566 9581 19585
rect 9003 19551 9037 19566
rect 9071 19551 9105 19566
rect 9139 19551 9173 19566
rect 9207 19551 9241 19566
rect 9275 19551 9309 19566
rect 9343 19551 9377 19566
rect 9411 19551 9445 19566
rect 9479 19551 9513 19566
rect 9547 19551 9581 19566
rect 9615 19566 9618 19585
rect 9683 19566 9690 19585
rect 9751 19566 9762 19585
rect 9819 19566 9834 19585
rect 9887 19566 9906 19585
rect 9955 19566 9978 19585
rect 10023 19566 10050 19585
rect 10091 19566 10122 19585
rect 9615 19551 9649 19566
rect 9683 19551 9717 19566
rect 9751 19551 9785 19566
rect 9819 19551 9853 19566
rect 9887 19551 9921 19566
rect 9955 19551 9989 19566
rect 10023 19551 10057 19566
rect 10091 19551 10125 19566
rect 10159 19551 10193 19585
rect 10228 19566 10261 19585
rect 10300 19566 10329 19585
rect 10372 19566 10397 19585
rect 10444 19566 10465 19585
rect 10516 19566 10533 19585
rect 10588 19566 10601 19585
rect 10660 19566 10669 19585
rect 10732 19566 10737 19585
rect 10804 19566 10805 19585
rect 10227 19551 10261 19566
rect 10295 19551 10329 19566
rect 10363 19551 10397 19566
rect 10431 19551 10465 19566
rect 10499 19551 10533 19566
rect 10567 19551 10601 19566
rect 10635 19551 10669 19566
rect 10703 19551 10737 19566
rect 10771 19551 10805 19566
rect 10839 19566 10842 19585
rect 10907 19566 10914 19585
rect 10975 19566 10986 19585
rect 11043 19566 11058 19585
rect 11111 19566 11130 19585
rect 11179 19566 11202 19585
rect 11247 19566 11274 19585
rect 11315 19566 11346 19585
rect 10839 19551 10873 19566
rect 10907 19551 10941 19566
rect 10975 19551 11009 19566
rect 11043 19551 11077 19566
rect 11111 19551 11145 19566
rect 11179 19551 11213 19566
rect 11247 19551 11281 19566
rect 11315 19551 11349 19566
rect 11383 19551 11417 19585
rect 11452 19566 11485 19585
rect 11524 19566 11553 19585
rect 11596 19566 11621 19585
rect 11668 19566 11689 19585
rect 11740 19566 11778 19600
rect 11812 19566 11850 19600
rect 11884 19566 11922 19600
rect 11956 19566 11994 19600
rect 12028 19566 12066 19600
rect 12100 19566 12138 19600
rect 12172 19566 12210 19600
rect 12244 19566 12282 19600
rect 12316 19566 12354 19600
rect 12388 19566 12426 19600
rect 12460 19566 12498 19600
rect 12532 19566 12570 19600
rect 12604 19566 12642 19600
rect 12676 19566 12714 19600
rect 12748 19566 12786 19600
rect 12820 19566 12858 19600
rect 12892 19566 12930 19600
rect 12964 19566 13002 19600
rect 13036 19566 13074 19600
rect 13108 19566 13146 19600
rect 13180 19566 13218 19600
rect 13252 19566 13290 19600
rect 13324 19566 13362 19600
rect 13396 19566 13434 19600
rect 13468 19566 13506 19600
rect 13540 19566 13578 19600
rect 13612 19566 13650 19600
rect 13684 19566 13722 19600
rect 13756 19566 13794 19600
rect 13828 19566 13866 19600
rect 13900 19566 13938 19600
rect 13972 19566 14010 19600
rect 14044 19566 14082 19600
rect 14116 19566 14154 19600
rect 14188 19566 14226 19600
rect 14260 19566 14298 19600
rect 14332 19566 14370 19600
rect 14404 19566 14442 19600
rect 14476 19587 14484 19600
rect 14548 19587 14567 19600
rect 14620 19587 14650 19600
rect 14476 19566 14514 19587
rect 14548 19566 14586 19587
rect 14620 19566 14658 19587
rect 14692 19566 14730 19600
rect 14767 19587 14802 19600
rect 14850 19587 14874 19600
rect 14764 19566 14802 19587
rect 14836 19566 14874 19587
rect 14908 19566 14959 19600
rect 11451 19551 11485 19566
rect 11519 19551 11553 19566
rect 11587 19551 11621 19566
rect 11655 19551 11689 19566
rect 11723 19557 14952 19566
rect 11723 19551 11771 19557
rect -41 19523 11771 19551
rect 11805 19523 11841 19557
rect 11875 19523 11911 19557
rect 11945 19523 11981 19557
rect 12015 19523 12051 19557
rect 12085 19523 12121 19557
rect 12155 19523 12191 19557
rect 12225 19523 12261 19557
rect 12295 19523 12331 19557
rect 12365 19523 12401 19557
rect 12435 19523 12470 19557
rect 12504 19523 12539 19557
rect 12573 19523 12608 19557
rect 12642 19523 12677 19557
rect 12711 19523 12746 19557
rect 12780 19523 12815 19557
rect 12849 19523 12884 19557
rect 12918 19523 12953 19557
rect 12987 19523 13022 19557
rect 13056 19523 13091 19557
rect 13125 19523 13160 19557
rect 13194 19523 13229 19557
rect 13263 19523 13298 19557
rect 13332 19523 13367 19557
rect 13401 19523 13436 19557
rect 13470 19523 13505 19557
rect 13539 19523 13574 19557
rect 13608 19523 13643 19557
rect 13677 19523 13712 19557
rect 13746 19523 13781 19557
rect 13815 19523 13850 19557
rect 13884 19523 13919 19557
rect 13953 19523 13988 19557
rect 14022 19523 14057 19557
rect 14091 19523 14126 19557
rect 14160 19523 14195 19557
rect 14229 19523 14264 19557
rect 14298 19523 14333 19557
rect 14367 19523 14402 19557
rect 14436 19551 14952 19557
rect 14436 19523 14484 19551
rect -41 19517 14484 19523
rect 14518 19517 14567 19551
rect 14601 19517 14650 19551
rect 14684 19517 14733 19551
rect 14767 19517 14816 19551
rect 14850 19517 14952 19551
rect -41 19513 14952 19517
rect -41 19479 77 19513
rect 111 19479 146 19513
rect 180 19479 215 19513
rect 249 19479 284 19513
rect 318 19479 353 19513
rect 387 19479 422 19513
rect 456 19479 491 19513
rect 525 19479 560 19513
rect 594 19479 629 19513
rect 663 19479 698 19513
rect 732 19479 767 19513
rect 801 19479 836 19513
rect 870 19479 905 19513
rect 939 19479 974 19513
rect 1008 19479 1043 19513
rect 1077 19479 1112 19513
rect 1146 19479 1181 19513
rect 1215 19479 1250 19513
rect 1284 19479 1319 19513
rect 1353 19479 1388 19513
rect 1422 19479 1457 19513
rect 1491 19479 1526 19513
rect 1560 19479 1595 19513
rect 1629 19479 1664 19513
rect 1698 19479 1733 19513
rect 1767 19479 1802 19513
rect 1836 19479 1871 19513
rect 1905 19479 1940 19513
rect 1974 19479 2009 19513
rect 2043 19479 2078 19513
rect 2112 19479 2147 19513
rect 2181 19479 2216 19513
rect 2250 19479 2285 19513
rect 2319 19479 2354 19513
rect 2388 19479 2423 19513
rect 2457 19479 2492 19513
rect 2526 19479 2561 19513
rect 2595 19479 2630 19513
rect 2664 19479 2699 19513
rect 2733 19479 2768 19513
rect 2802 19479 2837 19513
rect 2871 19479 2906 19513
rect 2940 19479 2975 19513
rect 3009 19479 3044 19513
rect 3078 19479 3113 19513
rect 3147 19479 3182 19513
rect 3216 19479 3251 19513
rect 3285 19479 3320 19513
rect 3354 19479 3389 19513
rect 3423 19479 3458 19513
rect 3492 19479 3527 19513
rect 3561 19479 3596 19513
rect 3630 19479 3665 19513
rect 3699 19479 3733 19513
rect 3767 19479 3801 19513
rect 3835 19479 3869 19513
rect 3903 19479 3937 19513
rect 3971 19479 4005 19513
rect 4039 19479 4073 19513
rect 4107 19479 4141 19513
rect 4175 19479 4209 19513
rect 4243 19479 4277 19513
rect 4311 19479 4345 19513
rect 4379 19479 4413 19513
rect 4447 19479 4481 19513
rect 4515 19479 4549 19513
rect 4583 19479 4617 19513
rect 4651 19479 4685 19513
rect 4719 19479 4753 19513
rect 4787 19479 4821 19513
rect 4855 19479 4889 19513
rect 4923 19479 4957 19513
rect 4991 19479 5025 19513
rect 5059 19479 5093 19513
rect 5127 19479 5161 19513
rect 5195 19479 5229 19513
rect 5263 19479 5297 19513
rect 5331 19479 5365 19513
rect 5399 19479 5433 19513
rect 5467 19479 5501 19513
rect 5535 19479 5569 19513
rect 5603 19479 5637 19513
rect 5671 19479 5705 19513
rect 5739 19479 5773 19513
rect 5807 19479 5841 19513
rect 5875 19479 5909 19513
rect 5943 19479 5977 19513
rect 6011 19479 6045 19513
rect 6079 19479 6113 19513
rect 6147 19479 6181 19513
rect 6215 19479 6249 19513
rect 6283 19479 6317 19513
rect 6351 19479 6385 19513
rect 6419 19479 6453 19513
rect 6487 19479 6521 19513
rect 6555 19479 6589 19513
rect 6623 19479 6657 19513
rect 6691 19479 6725 19513
rect 6759 19479 6793 19513
rect 6827 19479 6861 19513
rect 6895 19479 6929 19513
rect 6963 19479 6997 19513
rect 7031 19479 7065 19513
rect 7099 19479 7133 19513
rect 7167 19479 7201 19513
rect 7235 19479 7269 19513
rect 7303 19479 7337 19513
rect 7371 19479 7405 19513
rect 7439 19479 7473 19513
rect 7507 19479 7541 19513
rect 7575 19479 7609 19513
rect 7643 19479 7677 19513
rect 7711 19479 7745 19513
rect 7779 19479 7813 19513
rect 7847 19479 7881 19513
rect 7915 19479 7949 19513
rect 7983 19479 8017 19513
rect 8051 19479 8085 19513
rect 8119 19479 8153 19513
rect 8187 19479 8221 19513
rect 8255 19479 8289 19513
rect 8323 19479 8357 19513
rect 8391 19479 8425 19513
rect 8459 19479 8493 19513
rect 8527 19479 8561 19513
rect 8595 19479 8629 19513
rect 8663 19479 8697 19513
rect 8731 19479 8765 19513
rect 8799 19479 8833 19513
rect 8867 19479 8901 19513
rect 8935 19479 8969 19513
rect 9003 19479 9037 19513
rect 9071 19479 9105 19513
rect 9139 19479 9173 19513
rect 9207 19479 9241 19513
rect 9275 19479 9309 19513
rect 9343 19479 9377 19513
rect 9411 19479 9445 19513
rect 9479 19479 9513 19513
rect 9547 19479 9581 19513
rect 9615 19479 9649 19513
rect 9683 19479 9717 19513
rect 9751 19479 9785 19513
rect 9819 19479 9853 19513
rect 9887 19479 9921 19513
rect 9955 19479 9989 19513
rect 10023 19479 10057 19513
rect 10091 19479 10125 19513
rect 10159 19479 10193 19513
rect 10227 19479 10261 19513
rect 10295 19479 10329 19513
rect 10363 19479 10397 19513
rect 10431 19479 10465 19513
rect 10499 19479 10533 19513
rect 10567 19479 10601 19513
rect 10635 19479 10669 19513
rect 10703 19479 10737 19513
rect 10771 19479 10805 19513
rect 10839 19479 10873 19513
rect 10907 19479 10941 19513
rect 10975 19479 11009 19513
rect 11043 19479 11077 19513
rect 11111 19479 11145 19513
rect 11179 19479 11213 19513
rect 11247 19479 11281 19513
rect 11315 19479 11349 19513
rect 11383 19479 11417 19513
rect 11451 19479 11485 19513
rect 11519 19479 11553 19513
rect 11587 19479 11621 19513
rect 11655 19479 11689 19513
rect 11723 19481 14952 19513
rect 11723 19479 14484 19481
rect -41 19477 14484 19479
rect -41 19443 11771 19477
rect 11805 19443 11841 19477
rect 11875 19443 11911 19477
rect 11945 19443 11981 19477
rect 12015 19443 12051 19477
rect 12085 19443 12121 19477
rect 12155 19443 12191 19477
rect 12225 19443 12261 19477
rect 12295 19443 12331 19477
rect 12365 19443 12401 19477
rect 12435 19443 12470 19477
rect 12504 19443 12539 19477
rect 12573 19443 12608 19477
rect 12642 19443 12677 19477
rect 12711 19443 12746 19477
rect 12780 19443 12815 19477
rect 12849 19443 12884 19477
rect 12918 19443 12953 19477
rect 12987 19443 13022 19477
rect 13056 19443 13091 19477
rect 13125 19443 13160 19477
rect 13194 19443 13229 19477
rect 13263 19443 13298 19477
rect 13332 19443 13367 19477
rect 13401 19443 13436 19477
rect 13470 19443 13505 19477
rect 13539 19443 13574 19477
rect 13608 19443 13643 19477
rect 13677 19443 13712 19477
rect 13746 19443 13781 19477
rect 13815 19443 13850 19477
rect 13884 19443 13919 19477
rect 13953 19443 13988 19477
rect 14022 19443 14057 19477
rect 14091 19443 14126 19477
rect 14160 19443 14195 19477
rect 14229 19443 14264 19477
rect 14298 19443 14333 19477
rect 14367 19443 14402 19477
rect 14436 19447 14484 19477
rect 14518 19447 14567 19481
rect 14601 19447 14650 19481
rect 14684 19447 14733 19481
rect 14767 19447 14816 19481
rect 14850 19447 14952 19481
rect 14436 19443 14952 19447
rect -41 19441 14952 19443
rect -41 19407 77 19441
rect 111 19407 146 19441
rect 180 19407 215 19441
rect 249 19407 284 19441
rect 318 19407 353 19441
rect 387 19407 422 19441
rect 456 19407 491 19441
rect 525 19407 560 19441
rect 594 19407 629 19441
rect 663 19407 698 19441
rect 732 19407 767 19441
rect 801 19407 836 19441
rect 870 19407 905 19441
rect 939 19407 974 19441
rect 1008 19407 1043 19441
rect 1077 19407 1112 19441
rect 1146 19407 1181 19441
rect 1215 19407 1250 19441
rect 1284 19407 1319 19441
rect 1353 19407 1388 19441
rect 1422 19407 1457 19441
rect 1491 19407 1526 19441
rect 1560 19407 1595 19441
rect 1629 19407 1664 19441
rect 1698 19407 1733 19441
rect 1767 19407 1802 19441
rect 1836 19407 1871 19441
rect 1905 19407 1940 19441
rect 1974 19407 2009 19441
rect 2043 19407 2078 19441
rect 2112 19407 2147 19441
rect 2181 19407 2216 19441
rect 2250 19407 2285 19441
rect 2319 19407 2354 19441
rect 2388 19407 2423 19441
rect 2457 19407 2492 19441
rect 2526 19407 2561 19441
rect 2595 19407 2630 19441
rect 2664 19407 2699 19441
rect 2733 19407 2768 19441
rect 2802 19407 2837 19441
rect 2871 19407 2906 19441
rect 2940 19407 2975 19441
rect 3009 19407 3044 19441
rect 3078 19407 3113 19441
rect 3147 19407 3182 19441
rect 3216 19407 3251 19441
rect 3285 19407 3320 19441
rect 3354 19407 3389 19441
rect 3423 19407 3458 19441
rect 3492 19407 3527 19441
rect 3561 19407 3596 19441
rect 3630 19407 3665 19441
rect 3699 19407 3733 19441
rect 3767 19407 3801 19441
rect 3835 19407 3869 19441
rect 3903 19407 3937 19441
rect 3971 19407 4005 19441
rect 4039 19407 4073 19441
rect 4107 19407 4141 19441
rect 4175 19407 4209 19441
rect 4243 19407 4277 19441
rect 4311 19407 4345 19441
rect 4379 19407 4413 19441
rect 4447 19407 4481 19441
rect 4515 19407 4549 19441
rect 4583 19407 4617 19441
rect 4651 19407 4685 19441
rect 4719 19407 4753 19441
rect 4787 19407 4821 19441
rect 4855 19407 4889 19441
rect 4923 19407 4957 19441
rect 4991 19407 5025 19441
rect 5059 19407 5093 19441
rect 5127 19407 5161 19441
rect 5195 19407 5229 19441
rect 5263 19407 5297 19441
rect 5331 19407 5365 19441
rect 5399 19407 5433 19441
rect 5467 19407 5501 19441
rect 5535 19407 5569 19441
rect 5603 19407 5637 19441
rect 5671 19407 5705 19441
rect 5739 19407 5773 19441
rect 5807 19407 5841 19441
rect 5875 19407 5909 19441
rect 5943 19407 5977 19441
rect 6011 19407 6045 19441
rect 6079 19407 6113 19441
rect 6147 19407 6181 19441
rect 6215 19407 6249 19441
rect 6283 19407 6317 19441
rect 6351 19407 6385 19441
rect 6419 19407 6453 19441
rect 6487 19407 6521 19441
rect 6555 19407 6589 19441
rect 6623 19407 6657 19441
rect 6691 19407 6725 19441
rect 6759 19407 6793 19441
rect 6827 19407 6861 19441
rect 6895 19407 6929 19441
rect 6963 19407 6997 19441
rect 7031 19407 7065 19441
rect 7099 19407 7133 19441
rect 7167 19407 7201 19441
rect 7235 19407 7269 19441
rect 7303 19407 7337 19441
rect 7371 19407 7405 19441
rect 7439 19407 7473 19441
rect 7507 19407 7541 19441
rect 7575 19407 7609 19441
rect 7643 19407 7677 19441
rect 7711 19407 7745 19441
rect 7779 19407 7813 19441
rect 7847 19407 7881 19441
rect 7915 19407 7949 19441
rect 7983 19407 8017 19441
rect 8051 19407 8085 19441
rect 8119 19407 8153 19441
rect 8187 19407 8221 19441
rect 8255 19407 8289 19441
rect 8323 19407 8357 19441
rect 8391 19407 8425 19441
rect 8459 19407 8493 19441
rect 8527 19407 8561 19441
rect 8595 19407 8629 19441
rect 8663 19407 8697 19441
rect 8731 19407 8765 19441
rect 8799 19407 8833 19441
rect 8867 19407 8901 19441
rect 8935 19407 8969 19441
rect 9003 19407 9037 19441
rect 9071 19407 9105 19441
rect 9139 19407 9173 19441
rect 9207 19407 9241 19441
rect 9275 19407 9309 19441
rect 9343 19407 9377 19441
rect 9411 19407 9445 19441
rect 9479 19407 9513 19441
rect 9547 19407 9581 19441
rect 9615 19407 9649 19441
rect 9683 19407 9717 19441
rect 9751 19407 9785 19441
rect 9819 19407 9853 19441
rect 9887 19407 9921 19441
rect 9955 19407 9989 19441
rect 10023 19407 10057 19441
rect 10091 19407 10125 19441
rect 10159 19407 10193 19441
rect 10227 19407 10261 19441
rect 10295 19407 10329 19441
rect 10363 19407 10397 19441
rect 10431 19407 10465 19441
rect 10499 19407 10533 19441
rect 10567 19407 10601 19441
rect 10635 19407 10669 19441
rect 10703 19407 10737 19441
rect 10771 19407 10805 19441
rect 10839 19407 10873 19441
rect 10907 19407 10941 19441
rect 10975 19407 11009 19441
rect 11043 19407 11077 19441
rect 11111 19407 11145 19441
rect 11179 19407 11213 19441
rect 11247 19407 11281 19441
rect 11315 19407 11349 19441
rect 11383 19407 11417 19441
rect 11451 19407 11485 19441
rect 11519 19407 11553 19441
rect 11587 19407 11621 19441
rect 11655 19407 11689 19441
rect 11723 19411 14952 19441
rect 11723 19407 14484 19411
rect -41 19397 14484 19407
rect -41 19369 11771 19397
rect -41 19335 77 19369
rect 111 19335 146 19369
rect 180 19335 215 19369
rect 249 19335 284 19369
rect 318 19335 353 19369
rect 387 19335 422 19369
rect 456 19335 491 19369
rect 525 19335 560 19369
rect 594 19335 629 19369
rect 663 19335 698 19369
rect 732 19335 767 19369
rect 801 19335 836 19369
rect 870 19335 905 19369
rect 939 19335 974 19369
rect 1008 19335 1043 19369
rect 1077 19335 1112 19369
rect 1146 19335 1181 19369
rect 1215 19335 1250 19369
rect 1284 19335 1319 19369
rect 1353 19335 1388 19369
rect 1422 19335 1457 19369
rect 1491 19335 1526 19369
rect 1560 19335 1595 19369
rect 1629 19335 1664 19369
rect 1698 19335 1733 19369
rect 1767 19335 1802 19369
rect 1836 19335 1871 19369
rect 1905 19335 1940 19369
rect 1974 19335 2009 19369
rect 2043 19335 2078 19369
rect 2112 19335 2147 19369
rect 2181 19335 2216 19369
rect 2250 19335 2285 19369
rect 2319 19335 2354 19369
rect 2388 19335 2423 19369
rect 2457 19335 2492 19369
rect 2526 19335 2561 19369
rect 2595 19335 2630 19369
rect 2664 19335 2699 19369
rect 2733 19335 2768 19369
rect 2802 19335 2837 19369
rect 2871 19335 2906 19369
rect 2940 19335 2975 19369
rect 3009 19335 3044 19369
rect 3078 19335 3113 19369
rect 3147 19335 3182 19369
rect 3216 19335 3251 19369
rect 3285 19335 3320 19369
rect 3354 19335 3389 19369
rect 3423 19335 3458 19369
rect 3492 19335 3527 19369
rect 3561 19335 3596 19369
rect 3630 19335 3665 19369
rect 3699 19335 3733 19369
rect 3767 19335 3801 19369
rect 3835 19335 3869 19369
rect 3903 19335 3937 19369
rect 3971 19335 4005 19369
rect 4039 19335 4073 19369
rect 4107 19335 4141 19369
rect 4175 19335 4209 19369
rect 4243 19335 4277 19369
rect 4311 19335 4345 19369
rect 4379 19335 4413 19369
rect 4447 19335 4481 19369
rect 4515 19335 4549 19369
rect 4583 19335 4617 19369
rect 4651 19335 4685 19369
rect 4719 19335 4753 19369
rect 4787 19335 4821 19369
rect 4855 19335 4889 19369
rect 4923 19335 4957 19369
rect 4991 19335 5025 19369
rect 5059 19335 5093 19369
rect 5127 19335 5161 19369
rect 5195 19335 5229 19369
rect 5263 19335 5297 19369
rect 5331 19335 5365 19369
rect 5399 19335 5433 19369
rect 5467 19335 5501 19369
rect 5535 19335 5569 19369
rect 5603 19335 5637 19369
rect 5671 19335 5705 19369
rect 5739 19335 5773 19369
rect 5807 19335 5841 19369
rect 5875 19335 5909 19369
rect 5943 19335 5977 19369
rect 6011 19335 6045 19369
rect 6079 19335 6113 19369
rect 6147 19335 6181 19369
rect 6215 19335 6249 19369
rect 6283 19335 6317 19369
rect 6351 19335 6385 19369
rect 6419 19335 6453 19369
rect 6487 19335 6521 19369
rect 6555 19335 6589 19369
rect 6623 19335 6657 19369
rect 6691 19335 6725 19369
rect 6759 19335 6793 19369
rect 6827 19335 6861 19369
rect 6895 19335 6929 19369
rect 6963 19335 6997 19369
rect 7031 19335 7065 19369
rect 7099 19335 7133 19369
rect 7167 19335 7201 19369
rect 7235 19335 7269 19369
rect 7303 19335 7337 19369
rect 7371 19335 7405 19369
rect 7439 19335 7473 19369
rect 7507 19335 7541 19369
rect 7575 19335 7609 19369
rect 7643 19335 7677 19369
rect 7711 19335 7745 19369
rect 7779 19335 7813 19369
rect 7847 19335 7881 19369
rect 7915 19335 7949 19369
rect 7983 19335 8017 19369
rect 8051 19335 8085 19369
rect 8119 19335 8153 19369
rect 8187 19335 8221 19369
rect 8255 19335 8289 19369
rect 8323 19335 8357 19369
rect 8391 19335 8425 19369
rect 8459 19335 8493 19369
rect 8527 19335 8561 19369
rect 8595 19335 8629 19369
rect 8663 19335 8697 19369
rect 8731 19335 8765 19369
rect 8799 19335 8833 19369
rect 8867 19335 8901 19369
rect 8935 19335 8969 19369
rect 9003 19335 9037 19369
rect 9071 19335 9105 19369
rect 9139 19335 9173 19369
rect 9207 19335 9241 19369
rect 9275 19335 9309 19369
rect 9343 19335 9377 19369
rect 9411 19335 9445 19369
rect 9479 19335 9513 19369
rect 9547 19335 9581 19369
rect 9615 19335 9649 19369
rect 9683 19335 9717 19369
rect 9751 19335 9785 19369
rect 9819 19335 9853 19369
rect 9887 19335 9921 19369
rect 9955 19335 9989 19369
rect 10023 19335 10057 19369
rect 10091 19335 10125 19369
rect 10159 19335 10193 19369
rect 10227 19335 10261 19369
rect 10295 19335 10329 19369
rect 10363 19335 10397 19369
rect 10431 19335 10465 19369
rect 10499 19335 10533 19369
rect 10567 19335 10601 19369
rect 10635 19335 10669 19369
rect 10703 19335 10737 19369
rect 10771 19335 10805 19369
rect 10839 19335 10873 19369
rect 10907 19335 10941 19369
rect 10975 19335 11009 19369
rect 11043 19335 11077 19369
rect 11111 19335 11145 19369
rect 11179 19335 11213 19369
rect 11247 19335 11281 19369
rect 11315 19335 11349 19369
rect 11383 19335 11417 19369
rect 11451 19335 11485 19369
rect 11519 19335 11553 19369
rect 11587 19335 11621 19369
rect 11655 19335 11689 19369
rect 11723 19363 11771 19369
rect 11805 19363 11841 19397
rect 11875 19363 11911 19397
rect 11945 19363 11981 19397
rect 12015 19363 12051 19397
rect 12085 19363 12121 19397
rect 12155 19363 12191 19397
rect 12225 19363 12261 19397
rect 12295 19363 12331 19397
rect 12365 19363 12401 19397
rect 12435 19363 12470 19397
rect 12504 19363 12539 19397
rect 12573 19363 12608 19397
rect 12642 19363 12677 19397
rect 12711 19363 12746 19397
rect 12780 19363 12815 19397
rect 12849 19363 12884 19397
rect 12918 19363 12953 19397
rect 12987 19363 13022 19397
rect 13056 19363 13091 19397
rect 13125 19363 13160 19397
rect 13194 19363 13229 19397
rect 13263 19363 13298 19397
rect 13332 19363 13367 19397
rect 13401 19363 13436 19397
rect 13470 19363 13505 19397
rect 13539 19363 13574 19397
rect 13608 19363 13643 19397
rect 13677 19363 13712 19397
rect 13746 19363 13781 19397
rect 13815 19363 13850 19397
rect 13884 19363 13919 19397
rect 13953 19363 13988 19397
rect 14022 19363 14057 19397
rect 14091 19363 14126 19397
rect 14160 19363 14195 19397
rect 14229 19363 14264 19397
rect 14298 19363 14333 19397
rect 14367 19363 14402 19397
rect 14436 19377 14484 19397
rect 14518 19377 14567 19411
rect 14601 19377 14650 19411
rect 14684 19377 14733 19411
rect 14767 19377 14816 19411
rect 14850 19377 14952 19411
rect 14436 19363 14952 19377
rect 11723 19341 14952 19363
rect 11723 19335 14484 19341
rect -41 19330 14484 19335
rect -41 19297 11747 19330
rect -41 19263 77 19297
rect 111 19263 146 19297
rect 180 19263 215 19297
rect 249 19263 284 19297
rect 318 19263 353 19297
rect 387 19263 422 19297
rect 456 19263 491 19297
rect 525 19263 560 19297
rect 594 19263 629 19297
rect 663 19263 698 19297
rect 732 19263 767 19297
rect 801 19263 836 19297
rect 870 19263 905 19297
rect 939 19263 974 19297
rect 1008 19263 1043 19297
rect 1077 19263 1112 19297
rect 1146 19263 1181 19297
rect 1215 19263 1250 19297
rect 1284 19263 1319 19297
rect 1353 19263 1388 19297
rect 1422 19263 1457 19297
rect 1491 19263 1526 19297
rect 1560 19263 1595 19297
rect 1629 19263 1664 19297
rect 1698 19263 1733 19297
rect 1767 19263 1802 19297
rect 1836 19263 1871 19297
rect 1905 19263 1940 19297
rect 1974 19263 2009 19297
rect 2043 19263 2078 19297
rect 2112 19263 2147 19297
rect 2181 19263 2216 19297
rect 2250 19263 2285 19297
rect 2319 19263 2354 19297
rect 2388 19263 2423 19297
rect 2457 19263 2492 19297
rect 2526 19263 2561 19297
rect 2595 19263 2630 19297
rect 2664 19263 2699 19297
rect 2733 19263 2768 19297
rect 2802 19263 2837 19297
rect 2871 19263 2906 19297
rect 2940 19263 2975 19297
rect 3009 19263 3044 19297
rect 3078 19263 3113 19297
rect 3147 19263 3182 19297
rect 3216 19263 3251 19297
rect 3285 19263 3320 19297
rect 3354 19263 3389 19297
rect 3423 19263 3458 19297
rect 3492 19263 3527 19297
rect 3561 19263 3596 19297
rect 3630 19263 3665 19297
rect 3699 19263 3733 19297
rect 3767 19263 3801 19297
rect 3835 19263 3869 19297
rect 3903 19263 3937 19297
rect 3971 19263 4005 19297
rect 4039 19263 4073 19297
rect 4107 19263 4141 19297
rect 4175 19263 4209 19297
rect 4243 19263 4277 19297
rect 4311 19263 4345 19297
rect 4379 19263 4413 19297
rect 4447 19263 4481 19297
rect 4515 19263 4549 19297
rect 4583 19263 4617 19297
rect 4651 19263 4685 19297
rect 4719 19263 4753 19297
rect 4787 19263 4821 19297
rect 4855 19263 4889 19297
rect 4923 19263 4957 19297
rect 4991 19263 5025 19297
rect 5059 19263 5093 19297
rect 5127 19263 5161 19297
rect 5195 19263 5229 19297
rect 5263 19263 5297 19297
rect 5331 19263 5365 19297
rect 5399 19263 5433 19297
rect 5467 19263 5501 19297
rect 5535 19263 5569 19297
rect 5603 19263 5637 19297
rect 5671 19263 5705 19297
rect 5739 19263 5773 19297
rect 5807 19263 5841 19297
rect 5875 19263 5909 19297
rect 5943 19263 5977 19297
rect 6011 19263 6045 19297
rect 6079 19263 6113 19297
rect 6147 19263 6181 19297
rect 6215 19263 6249 19297
rect 6283 19263 6317 19297
rect 6351 19263 6385 19297
rect 6419 19263 6453 19297
rect 6487 19263 6521 19297
rect 6555 19263 6589 19297
rect 6623 19263 6657 19297
rect 6691 19263 6725 19297
rect 6759 19263 6793 19297
rect 6827 19263 6861 19297
rect 6895 19263 6929 19297
rect 6963 19263 6997 19297
rect 7031 19263 7065 19297
rect 7099 19263 7133 19297
rect 7167 19263 7201 19297
rect 7235 19263 7269 19297
rect 7303 19263 7337 19297
rect 7371 19263 7405 19297
rect 7439 19263 7473 19297
rect 7507 19263 7541 19297
rect 7575 19263 7609 19297
rect 7643 19263 7677 19297
rect 7711 19263 7745 19297
rect 7779 19263 7813 19297
rect 7847 19263 7881 19297
rect 7915 19263 7949 19297
rect 7983 19263 8017 19297
rect 8051 19263 8085 19297
rect 8119 19263 8153 19297
rect 8187 19263 8221 19297
rect 8255 19263 8289 19297
rect 8323 19263 8357 19297
rect 8391 19263 8425 19297
rect 8459 19263 8493 19297
rect 8527 19263 8561 19297
rect 8595 19263 8629 19297
rect 8663 19263 8697 19297
rect 8731 19263 8765 19297
rect 8799 19263 8833 19297
rect 8867 19263 8901 19297
rect 8935 19263 8969 19297
rect 9003 19263 9037 19297
rect 9071 19263 9105 19297
rect 9139 19263 9173 19297
rect 9207 19263 9241 19297
rect 9275 19263 9309 19297
rect 9343 19263 9377 19297
rect 9411 19263 9445 19297
rect 9479 19263 9513 19297
rect 9547 19263 9581 19297
rect 9615 19263 9649 19297
rect 9683 19263 9717 19297
rect 9751 19263 9785 19297
rect 9819 19263 9853 19297
rect 9887 19263 9921 19297
rect 9955 19263 9989 19297
rect 10023 19263 10057 19297
rect 10091 19263 10125 19297
rect 10159 19263 10193 19297
rect 10227 19263 10261 19297
rect 10295 19263 10329 19297
rect 10363 19263 10397 19297
rect 10431 19263 10465 19297
rect 10499 19263 10533 19297
rect 10567 19263 10601 19297
rect 10635 19263 10669 19297
rect 10703 19263 10737 19297
rect 10771 19263 10805 19297
rect 10839 19263 10873 19297
rect 10907 19263 10941 19297
rect 10975 19263 11009 19297
rect 11043 19263 11077 19297
rect 11111 19263 11145 19297
rect 11179 19263 11213 19297
rect 11247 19263 11281 19297
rect 11315 19263 11349 19297
rect 11383 19263 11417 19297
rect 11451 19263 11485 19297
rect 11519 19263 11553 19297
rect 11587 19263 11621 19297
rect 11655 19263 11689 19297
rect 11723 19263 11747 19297
rect -41 19225 11747 19263
rect -41 19191 77 19225
rect 111 19191 146 19225
rect 180 19191 215 19225
rect 249 19191 284 19225
rect 318 19191 353 19225
rect 387 19191 422 19225
rect 456 19191 491 19225
rect 525 19191 560 19225
rect 594 19191 629 19225
rect 663 19191 698 19225
rect 732 19191 767 19225
rect 801 19191 836 19225
rect 870 19191 905 19225
rect 939 19191 974 19225
rect 1008 19191 1043 19225
rect 1077 19191 1112 19225
rect 1146 19191 1181 19225
rect 1215 19191 1250 19225
rect 1284 19191 1319 19225
rect 1353 19191 1388 19225
rect 1422 19191 1457 19225
rect 1491 19191 1526 19225
rect 1560 19191 1595 19225
rect 1629 19191 1664 19225
rect 1698 19191 1733 19225
rect 1767 19191 1802 19225
rect 1836 19191 1871 19225
rect 1905 19191 1940 19225
rect 1974 19191 2009 19225
rect 2043 19191 2078 19225
rect 2112 19191 2147 19225
rect 2181 19191 2216 19225
rect 2250 19191 2285 19225
rect 2319 19191 2354 19225
rect 2388 19191 2423 19225
rect 2457 19191 2492 19225
rect 2526 19191 2561 19225
rect 2595 19191 2630 19225
rect 2664 19191 2699 19225
rect 2733 19191 2768 19225
rect 2802 19191 2837 19225
rect 2871 19191 2906 19225
rect 2940 19191 2975 19225
rect 3009 19191 3044 19225
rect 3078 19191 3113 19225
rect 3147 19191 3182 19225
rect 3216 19191 3251 19225
rect 3285 19191 3320 19225
rect 3354 19191 3389 19225
rect 3423 19191 3458 19225
rect 3492 19191 3527 19225
rect 3561 19191 3596 19225
rect 3630 19191 3665 19225
rect 3699 19191 3733 19225
rect 3767 19191 3801 19225
rect 3835 19191 3869 19225
rect 3903 19191 3937 19225
rect 3971 19191 4005 19225
rect 4039 19191 4073 19225
rect 4107 19191 4141 19225
rect 4175 19191 4209 19225
rect 4243 19191 4277 19225
rect 4311 19191 4345 19225
rect 4379 19191 4413 19225
rect 4447 19191 4481 19225
rect 4515 19191 4549 19225
rect 4583 19191 4617 19225
rect 4651 19191 4685 19225
rect 4719 19191 4753 19225
rect 4787 19191 4821 19225
rect 4855 19191 4889 19225
rect 4923 19191 4957 19225
rect 4991 19191 5025 19225
rect 5059 19191 5093 19225
rect 5127 19191 5161 19225
rect 5195 19191 5229 19225
rect 5263 19191 5297 19225
rect 5331 19191 5365 19225
rect 5399 19191 5433 19225
rect 5467 19191 5501 19225
rect 5535 19191 5569 19225
rect 5603 19191 5637 19225
rect 5671 19191 5705 19225
rect 5739 19191 5773 19225
rect 5807 19191 5841 19225
rect 5875 19191 5909 19225
rect 5943 19191 5977 19225
rect 6011 19191 6045 19225
rect 6079 19191 6113 19225
rect 6147 19191 6181 19225
rect 6215 19191 6249 19225
rect 6283 19191 6317 19225
rect 6351 19191 6385 19225
rect 6419 19191 6453 19225
rect 6487 19191 6521 19225
rect 6555 19191 6589 19225
rect 6623 19191 6657 19225
rect 6691 19191 6725 19225
rect 6759 19191 6793 19225
rect 6827 19191 6861 19225
rect 6895 19191 6929 19225
rect 6963 19191 6997 19225
rect 7031 19191 7065 19225
rect 7099 19191 7133 19225
rect 7167 19191 7201 19225
rect 7235 19191 7269 19225
rect 7303 19191 7337 19225
rect 7371 19191 7405 19225
rect 7439 19191 7473 19225
rect 7507 19191 7541 19225
rect 7575 19191 7609 19225
rect 7643 19191 7677 19225
rect 7711 19191 7745 19225
rect 7779 19191 7813 19225
rect 7847 19191 7881 19225
rect 7915 19191 7949 19225
rect 7983 19191 8017 19225
rect 8051 19191 8085 19225
rect 8119 19191 8153 19225
rect 8187 19191 8221 19225
rect 8255 19191 8289 19225
rect 8323 19191 8357 19225
rect 8391 19191 8425 19225
rect 8459 19191 8493 19225
rect 8527 19191 8561 19225
rect 8595 19191 8629 19225
rect 8663 19191 8697 19225
rect 8731 19191 8765 19225
rect 8799 19191 8833 19225
rect 8867 19191 8901 19225
rect 8935 19191 8969 19225
rect 9003 19191 9037 19225
rect 9071 19191 9105 19225
rect 9139 19191 9173 19225
rect 9207 19191 9241 19225
rect 9275 19191 9309 19225
rect 9343 19191 9377 19225
rect 9411 19191 9445 19225
rect 9479 19191 9513 19225
rect 9547 19191 9581 19225
rect 9615 19191 9649 19225
rect 9683 19191 9717 19225
rect 9751 19191 9785 19225
rect 9819 19191 9853 19225
rect 9887 19191 9921 19225
rect 9955 19191 9989 19225
rect 10023 19191 10057 19225
rect 10091 19191 10125 19225
rect 10159 19191 10193 19225
rect 10227 19191 10261 19225
rect 10295 19191 10329 19225
rect 10363 19191 10397 19225
rect 10431 19191 10465 19225
rect 10499 19191 10533 19225
rect 10567 19191 10601 19225
rect 10635 19191 10669 19225
rect 10703 19191 10737 19225
rect 10771 19191 10805 19225
rect 10839 19191 10873 19225
rect 10907 19191 10941 19225
rect 10975 19191 11009 19225
rect 11043 19191 11077 19225
rect 11111 19191 11145 19225
rect 11179 19191 11213 19225
rect 11247 19191 11281 19225
rect 11315 19191 11349 19225
rect 11383 19191 11417 19225
rect 11451 19191 11485 19225
rect 11519 19191 11553 19225
rect 11587 19191 11621 19225
rect 11655 19191 11689 19225
rect 11723 19191 11747 19225
rect -41 19153 11747 19191
rect -41 19119 77 19153
rect 111 19119 146 19153
rect 180 19119 215 19153
rect 249 19119 284 19153
rect 318 19119 353 19153
rect 387 19119 422 19153
rect 456 19119 491 19153
rect 525 19119 560 19153
rect 594 19119 629 19153
rect 663 19119 698 19153
rect 732 19119 767 19153
rect 801 19119 836 19153
rect 870 19119 905 19153
rect 939 19119 974 19153
rect 1008 19119 1043 19153
rect 1077 19119 1112 19153
rect 1146 19119 1181 19153
rect 1215 19119 1250 19153
rect 1284 19119 1319 19153
rect 1353 19119 1388 19153
rect 1422 19119 1457 19153
rect 1491 19119 1526 19153
rect 1560 19119 1595 19153
rect 1629 19119 1664 19153
rect 1698 19119 1733 19153
rect 1767 19119 1802 19153
rect 1836 19119 1871 19153
rect 1905 19119 1940 19153
rect 1974 19119 2009 19153
rect 2043 19119 2078 19153
rect 2112 19119 2147 19153
rect 2181 19119 2216 19153
rect 2250 19119 2285 19153
rect 2319 19119 2354 19153
rect 2388 19119 2423 19153
rect 2457 19119 2492 19153
rect 2526 19119 2561 19153
rect 2595 19119 2630 19153
rect 2664 19119 2699 19153
rect 2733 19119 2768 19153
rect 2802 19119 2837 19153
rect 2871 19119 2906 19153
rect 2940 19119 2975 19153
rect 3009 19119 3044 19153
rect 3078 19119 3113 19153
rect 3147 19119 3182 19153
rect 3216 19119 3251 19153
rect 3285 19119 3320 19153
rect 3354 19119 3389 19153
rect 3423 19119 3458 19153
rect 3492 19119 3527 19153
rect 3561 19119 3596 19153
rect 3630 19119 3665 19153
rect 3699 19119 3733 19153
rect 3767 19119 3801 19153
rect 3835 19119 3869 19153
rect 3903 19119 3937 19153
rect 3971 19119 4005 19153
rect 4039 19119 4073 19153
rect 4107 19119 4141 19153
rect 4175 19119 4209 19153
rect 4243 19119 4277 19153
rect 4311 19119 4345 19153
rect 4379 19119 4413 19153
rect 4447 19119 4481 19153
rect 4515 19119 4549 19153
rect 4583 19119 4617 19153
rect 4651 19119 4685 19153
rect 4719 19119 4753 19153
rect 4787 19119 4821 19153
rect 4855 19119 4889 19153
rect 4923 19119 4957 19153
rect 4991 19119 5025 19153
rect 5059 19119 5093 19153
rect 5127 19119 5161 19153
rect 5195 19119 5229 19153
rect 5263 19119 5297 19153
rect 5331 19119 5365 19153
rect 5399 19119 5433 19153
rect 5467 19119 5501 19153
rect 5535 19119 5569 19153
rect 5603 19119 5637 19153
rect 5671 19119 5705 19153
rect 5739 19119 5773 19153
rect 5807 19119 5841 19153
rect 5875 19119 5909 19153
rect 5943 19119 5977 19153
rect 6011 19119 6045 19153
rect 6079 19119 6113 19153
rect 6147 19119 6181 19153
rect 6215 19119 6249 19153
rect 6283 19119 6317 19153
rect 6351 19119 6385 19153
rect 6419 19119 6453 19153
rect 6487 19119 6521 19153
rect 6555 19119 6589 19153
rect 6623 19119 6657 19153
rect 6691 19119 6725 19153
rect 6759 19119 6793 19153
rect 6827 19119 6861 19153
rect 6895 19119 6929 19153
rect 6963 19119 6997 19153
rect 7031 19119 7065 19153
rect 7099 19119 7133 19153
rect 7167 19119 7201 19153
rect 7235 19119 7269 19153
rect 7303 19119 7337 19153
rect 7371 19119 7405 19153
rect 7439 19119 7473 19153
rect 7507 19119 7541 19153
rect 7575 19119 7609 19153
rect 7643 19119 7677 19153
rect 7711 19119 7745 19153
rect 7779 19119 7813 19153
rect 7847 19119 7881 19153
rect 7915 19119 7949 19153
rect 7983 19119 8017 19153
rect 8051 19119 8085 19153
rect 8119 19119 8153 19153
rect 8187 19119 8221 19153
rect 8255 19119 8289 19153
rect 8323 19119 8357 19153
rect 8391 19119 8425 19153
rect 8459 19119 8493 19153
rect 8527 19119 8561 19153
rect 8595 19119 8629 19153
rect 8663 19119 8697 19153
rect 8731 19119 8765 19153
rect 8799 19119 8833 19153
rect 8867 19119 8901 19153
rect 8935 19119 8969 19153
rect 9003 19119 9037 19153
rect 9071 19119 9105 19153
rect 9139 19119 9173 19153
rect 9207 19119 9241 19153
rect 9275 19119 9309 19153
rect 9343 19119 9377 19153
rect 9411 19119 9445 19153
rect 9479 19119 9513 19153
rect 9547 19119 9581 19153
rect 9615 19119 9649 19153
rect 9683 19119 9717 19153
rect 9751 19119 9785 19153
rect 9819 19119 9853 19153
rect 9887 19119 9921 19153
rect 9955 19119 9989 19153
rect 10023 19119 10057 19153
rect 10091 19119 10125 19153
rect 10159 19119 10193 19153
rect 10227 19119 10261 19153
rect 10295 19119 10329 19153
rect 10363 19119 10397 19153
rect 10431 19119 10465 19153
rect 10499 19119 10533 19153
rect 10567 19119 10601 19153
rect 10635 19119 10669 19153
rect 10703 19119 10737 19153
rect 10771 19119 10805 19153
rect 10839 19119 10873 19153
rect 10907 19119 10941 19153
rect 10975 19119 11009 19153
rect 11043 19119 11077 19153
rect 11111 19119 11145 19153
rect 11179 19119 11213 19153
rect 11247 19119 11281 19153
rect 11315 19119 11349 19153
rect 11383 19119 11417 19153
rect 11451 19119 11485 19153
rect 11519 19119 11553 19153
rect 11587 19119 11621 19153
rect 11655 19119 11689 19153
rect 11723 19119 11747 19153
rect -41 19081 11747 19119
rect -41 19047 77 19081
rect 111 19047 146 19081
rect 180 19047 215 19081
rect 249 19047 284 19081
rect 318 19047 353 19081
rect 387 19047 422 19081
rect 456 19047 491 19081
rect 525 19047 560 19081
rect 594 19047 629 19081
rect 663 19047 698 19081
rect 732 19047 767 19081
rect 801 19047 836 19081
rect 870 19047 905 19081
rect 939 19047 974 19081
rect 1008 19047 1043 19081
rect 1077 19047 1112 19081
rect 1146 19047 1181 19081
rect 1215 19047 1250 19081
rect 1284 19047 1319 19081
rect 1353 19047 1388 19081
rect 1422 19047 1457 19081
rect 1491 19047 1526 19081
rect 1560 19047 1595 19081
rect 1629 19047 1664 19081
rect 1698 19047 1733 19081
rect 1767 19047 1802 19081
rect 1836 19047 1871 19081
rect 1905 19047 1940 19081
rect 1974 19047 2009 19081
rect 2043 19047 2078 19081
rect 2112 19047 2147 19081
rect 2181 19047 2216 19081
rect 2250 19047 2285 19081
rect 2319 19047 2354 19081
rect 2388 19047 2423 19081
rect 2457 19047 2492 19081
rect 2526 19047 2561 19081
rect 2595 19047 2630 19081
rect 2664 19047 2699 19081
rect 2733 19047 2768 19081
rect 2802 19047 2837 19081
rect 2871 19047 2906 19081
rect 2940 19047 2975 19081
rect 3009 19047 3044 19081
rect 3078 19047 3113 19081
rect 3147 19047 3182 19081
rect 3216 19047 3251 19081
rect 3285 19047 3320 19081
rect 3354 19047 3389 19081
rect 3423 19047 3458 19081
rect 3492 19047 3527 19081
rect 3561 19047 3596 19081
rect 3630 19047 3665 19081
rect 3699 19047 3733 19081
rect 3767 19047 3801 19081
rect 3835 19047 3869 19081
rect 3903 19047 3937 19081
rect 3971 19047 4005 19081
rect 4039 19047 4073 19081
rect 4107 19047 4141 19081
rect 4175 19047 4209 19081
rect 4243 19047 4277 19081
rect 4311 19047 4345 19081
rect 4379 19047 4413 19081
rect 4447 19047 4481 19081
rect 4515 19047 4549 19081
rect 4583 19047 4617 19081
rect 4651 19047 4685 19081
rect 4719 19047 4753 19081
rect 4787 19047 4821 19081
rect 4855 19047 4889 19081
rect 4923 19047 4957 19081
rect 4991 19047 5025 19081
rect 5059 19047 5093 19081
rect 5127 19047 5161 19081
rect 5195 19047 5229 19081
rect 5263 19047 5297 19081
rect 5331 19047 5365 19081
rect 5399 19047 5433 19081
rect 5467 19047 5501 19081
rect 5535 19047 5569 19081
rect 5603 19047 5637 19081
rect 5671 19047 5705 19081
rect 5739 19047 5773 19081
rect 5807 19047 5841 19081
rect 5875 19047 5909 19081
rect 5943 19047 5977 19081
rect 6011 19047 6045 19081
rect 6079 19047 6113 19081
rect 6147 19047 6181 19081
rect 6215 19047 6249 19081
rect 6283 19047 6317 19081
rect 6351 19047 6385 19081
rect 6419 19047 6453 19081
rect 6487 19047 6521 19081
rect 6555 19047 6589 19081
rect 6623 19047 6657 19081
rect 6691 19047 6725 19081
rect 6759 19047 6793 19081
rect 6827 19047 6861 19081
rect 6895 19047 6929 19081
rect 6963 19047 6997 19081
rect 7031 19047 7065 19081
rect 7099 19047 7133 19081
rect 7167 19047 7201 19081
rect 7235 19047 7269 19081
rect 7303 19047 7337 19081
rect 7371 19047 7405 19081
rect 7439 19047 7473 19081
rect 7507 19047 7541 19081
rect 7575 19047 7609 19081
rect 7643 19047 7677 19081
rect 7711 19047 7745 19081
rect 7779 19047 7813 19081
rect 7847 19047 7881 19081
rect 7915 19047 7949 19081
rect 7983 19047 8017 19081
rect 8051 19047 8085 19081
rect 8119 19047 8153 19081
rect 8187 19047 8221 19081
rect 8255 19047 8289 19081
rect 8323 19047 8357 19081
rect 8391 19047 8425 19081
rect 8459 19047 8493 19081
rect 8527 19047 8561 19081
rect 8595 19047 8629 19081
rect 8663 19047 8697 19081
rect 8731 19047 8765 19081
rect 8799 19047 8833 19081
rect 8867 19047 8901 19081
rect 8935 19047 8969 19081
rect 9003 19047 9037 19081
rect 9071 19047 9105 19081
rect 9139 19047 9173 19081
rect 9207 19047 9241 19081
rect 9275 19047 9309 19081
rect 9343 19047 9377 19081
rect 9411 19047 9445 19081
rect 9479 19047 9513 19081
rect 9547 19047 9581 19081
rect 9615 19047 9649 19081
rect 9683 19047 9717 19081
rect 9751 19047 9785 19081
rect 9819 19047 9853 19081
rect 9887 19047 9921 19081
rect 9955 19047 9989 19081
rect 10023 19047 10057 19081
rect 10091 19047 10125 19081
rect 10159 19047 10193 19081
rect 10227 19047 10261 19081
rect 10295 19047 10329 19081
rect 10363 19047 10397 19081
rect 10431 19047 10465 19081
rect 10499 19047 10533 19081
rect 10567 19047 10601 19081
rect 10635 19047 10669 19081
rect 10703 19047 10737 19081
rect 10771 19047 10805 19081
rect 10839 19047 10873 19081
rect 10907 19047 10941 19081
rect 10975 19047 11009 19081
rect 11043 19047 11077 19081
rect 11111 19047 11145 19081
rect 11179 19047 11213 19081
rect 11247 19047 11281 19081
rect 11315 19047 11349 19081
rect 11383 19047 11417 19081
rect 11451 19047 11485 19081
rect 11519 19047 11553 19081
rect 11587 19047 11621 19081
rect 11655 19047 11689 19081
rect 11723 19047 11747 19081
rect -41 19009 11747 19047
rect -41 18975 77 19009
rect 111 18975 146 19009
rect 180 18975 215 19009
rect 249 18975 284 19009
rect 318 18975 353 19009
rect 387 18975 422 19009
rect 456 18975 491 19009
rect 525 18975 560 19009
rect 594 18975 629 19009
rect 663 18975 698 19009
rect 732 18975 767 19009
rect 801 18975 836 19009
rect 870 18975 905 19009
rect 939 18975 974 19009
rect 1008 18975 1043 19009
rect 1077 18975 1112 19009
rect 1146 18975 1181 19009
rect 1215 18975 1250 19009
rect 1284 18975 1319 19009
rect 1353 18975 1388 19009
rect 1422 18975 1457 19009
rect 1491 18975 1526 19009
rect 1560 18975 1595 19009
rect 1629 18975 1664 19009
rect 1698 18975 1733 19009
rect 1767 18975 1802 19009
rect 1836 18975 1871 19009
rect 1905 18975 1940 19009
rect 1974 18975 2009 19009
rect 2043 18975 2078 19009
rect 2112 18975 2147 19009
rect 2181 18975 2216 19009
rect 2250 18975 2285 19009
rect 2319 18975 2354 19009
rect 2388 18975 2423 19009
rect 2457 18975 2492 19009
rect 2526 18975 2561 19009
rect 2595 18975 2630 19009
rect 2664 18975 2699 19009
rect 2733 18975 2768 19009
rect 2802 18975 2837 19009
rect 2871 18975 2906 19009
rect 2940 18975 2975 19009
rect 3009 18975 3044 19009
rect 3078 18975 3113 19009
rect 3147 18975 3182 19009
rect 3216 18975 3251 19009
rect 3285 18975 3320 19009
rect 3354 18975 3389 19009
rect 3423 18975 3458 19009
rect 3492 18975 3527 19009
rect 3561 18975 3596 19009
rect 3630 18975 3665 19009
rect 3699 18975 3733 19009
rect 3767 18975 3801 19009
rect 3835 18975 3869 19009
rect 3903 18975 3937 19009
rect 3971 18975 4005 19009
rect 4039 18975 4073 19009
rect 4107 18975 4141 19009
rect 4175 18975 4209 19009
rect 4243 18975 4277 19009
rect 4311 18975 4345 19009
rect 4379 18975 4413 19009
rect 4447 18975 4481 19009
rect 4515 18975 4549 19009
rect 4583 18975 4617 19009
rect 4651 18975 4685 19009
rect 4719 18975 4753 19009
rect 4787 18975 4821 19009
rect 4855 18975 4889 19009
rect 4923 18975 4957 19009
rect 4991 18975 5025 19009
rect 5059 18975 5093 19009
rect 5127 18975 5161 19009
rect 5195 18975 5229 19009
rect 5263 18975 5297 19009
rect 5331 18975 5365 19009
rect 5399 18975 5433 19009
rect 5467 18975 5501 19009
rect 5535 18975 5569 19009
rect 5603 18975 5637 19009
rect 5671 18975 5705 19009
rect 5739 18975 5773 19009
rect 5807 18975 5841 19009
rect 5875 18975 5909 19009
rect 5943 18975 5977 19009
rect 6011 18975 6045 19009
rect 6079 18975 6113 19009
rect 6147 18975 6181 19009
rect 6215 18975 6249 19009
rect 6283 18975 6317 19009
rect 6351 18975 6385 19009
rect 6419 18975 6453 19009
rect 6487 18975 6521 19009
rect 6555 18975 6589 19009
rect 6623 18975 6657 19009
rect 6691 18975 6725 19009
rect 6759 18975 6793 19009
rect 6827 18975 6861 19009
rect 6895 18975 6929 19009
rect 6963 18975 6997 19009
rect 7031 18975 7065 19009
rect 7099 18975 7133 19009
rect 7167 18975 7201 19009
rect 7235 18975 7269 19009
rect 7303 18975 7337 19009
rect 7371 18975 7405 19009
rect 7439 18975 7473 19009
rect 7507 18975 7541 19009
rect 7575 18975 7609 19009
rect 7643 18975 7677 19009
rect 7711 18975 7745 19009
rect 7779 18975 7813 19009
rect 7847 18975 7881 19009
rect 7915 18975 7949 19009
rect 7983 18975 8017 19009
rect 8051 18975 8085 19009
rect 8119 18975 8153 19009
rect 8187 18975 8221 19009
rect 8255 18975 8289 19009
rect 8323 18975 8357 19009
rect 8391 18975 8425 19009
rect 8459 18975 8493 19009
rect 8527 18975 8561 19009
rect 8595 18975 8629 19009
rect 8663 18975 8697 19009
rect 8731 18975 8765 19009
rect 8799 18975 8833 19009
rect 8867 18975 8901 19009
rect 8935 18975 8969 19009
rect 9003 18975 9037 19009
rect 9071 18975 9105 19009
rect 9139 18975 9173 19009
rect 9207 18975 9241 19009
rect 9275 18975 9309 19009
rect 9343 18975 9377 19009
rect 9411 18975 9445 19009
rect 9479 18975 9513 19009
rect 9547 18975 9581 19009
rect 9615 18975 9649 19009
rect 9683 18975 9717 19009
rect 9751 18975 9785 19009
rect 9819 18975 9853 19009
rect 9887 18975 9921 19009
rect 9955 18975 9989 19009
rect 10023 18975 10057 19009
rect 10091 18975 10125 19009
rect 10159 18975 10193 19009
rect 10227 18975 10261 19009
rect 10295 18975 10329 19009
rect 10363 18975 10397 19009
rect 10431 18975 10465 19009
rect 10499 18975 10533 19009
rect 10567 18975 10601 19009
rect 10635 18975 10669 19009
rect 10703 18975 10737 19009
rect 10771 18975 10805 19009
rect 10839 18975 10873 19009
rect 10907 18975 10941 19009
rect 10975 18975 11009 19009
rect 11043 18975 11077 19009
rect 11111 18975 11145 19009
rect 11179 18975 11213 19009
rect 11247 18975 11281 19009
rect 11315 18975 11349 19009
rect 11383 18975 11417 19009
rect 11451 18975 11485 19009
rect 11519 18975 11553 19009
rect 11587 18975 11621 19009
rect 11655 18975 11689 19009
rect 11723 18975 11747 19009
rect -41 18915 11747 18975
rect 14460 19307 14484 19330
rect 14518 19307 14567 19341
rect 14601 19307 14650 19341
rect 14684 19307 14733 19341
rect 14767 19307 14816 19341
rect 14850 19307 14952 19341
rect 14460 19271 14952 19307
rect 14460 19237 14484 19271
rect 14518 19237 14567 19271
rect 14601 19237 14650 19271
rect 14684 19237 14733 19271
rect 14767 19237 14816 19271
rect 14850 19237 14952 19271
rect 14460 19201 14952 19237
rect 14460 19167 14484 19201
rect 14518 19167 14567 19201
rect 14601 19167 14650 19201
rect 14684 19167 14733 19201
rect 14767 19167 14816 19201
rect 14850 19167 14952 19201
rect 14460 19131 14952 19167
rect 14460 19097 14484 19131
rect 14518 19097 14567 19131
rect 14601 19097 14650 19131
rect 14684 19097 14733 19131
rect 14767 19097 14816 19131
rect 14850 19097 14952 19131
rect 14460 19061 14952 19097
rect 14460 19027 14484 19061
rect 14518 19027 14567 19061
rect 14601 19027 14650 19061
rect 14684 19027 14733 19061
rect 14767 19027 14816 19061
rect 14850 19027 14952 19061
rect 14460 18915 14952 19027
rect -41 18881 77 18915
rect 111 18881 146 18915
rect 180 18881 215 18915
rect 249 18881 284 18915
rect 318 18881 353 18915
rect 387 18881 422 18915
rect 456 18881 491 18915
rect 525 18881 560 18915
rect 594 18881 629 18915
rect 663 18881 698 18915
rect 732 18881 767 18915
rect 801 18881 836 18915
rect 870 18881 905 18915
rect 939 18881 974 18915
rect 1008 18881 1043 18915
rect 1077 18881 1112 18915
rect 1146 18881 1181 18915
rect 1215 18881 1250 18915
rect 1284 18881 1319 18915
rect 1353 18881 1388 18915
rect 1422 18881 1457 18915
rect 1491 18881 1526 18915
rect 1560 18881 1595 18915
rect 1629 18881 1664 18915
rect 1698 18881 1733 18915
rect 1767 18881 1802 18915
rect 1836 18881 1871 18915
rect 1905 18881 1940 18915
rect 1974 18881 2009 18915
rect 2043 18881 2078 18915
rect 2112 18881 2147 18915
rect 2181 18881 2216 18915
rect 2250 18881 2285 18915
rect 2319 18881 2354 18915
rect 2388 18881 2423 18915
rect 2457 18881 2492 18915
rect 2526 18881 2561 18915
rect 2595 18881 2630 18915
rect 2664 18881 2699 18915
rect 2733 18881 2768 18915
rect 2802 18881 2837 18915
rect 2871 18881 2906 18915
rect 2940 18881 2975 18915
rect 3009 18881 3044 18915
rect 3078 18881 3113 18915
rect 3147 18881 3182 18915
rect 3216 18881 3251 18915
rect 3285 18881 3320 18915
rect 3354 18881 3389 18915
rect 3423 18881 3458 18915
rect 3492 18881 3527 18915
rect 3561 18881 3596 18915
rect -41 18847 3596 18881
rect -41 18813 77 18847
rect 111 18813 146 18847
rect 180 18813 215 18847
rect 249 18813 284 18847
rect 318 18813 353 18847
rect 387 18813 422 18847
rect 456 18813 491 18847
rect 525 18813 560 18847
rect 594 18813 629 18847
rect 663 18813 698 18847
rect 732 18813 767 18847
rect 801 18813 836 18847
rect 870 18813 905 18847
rect 939 18813 974 18847
rect 1008 18813 1043 18847
rect 1077 18813 1112 18847
rect 1146 18813 1181 18847
rect 1215 18813 1250 18847
rect 1284 18813 1319 18847
rect 1353 18813 1388 18847
rect 1422 18813 1457 18847
rect 1491 18813 1526 18847
rect 1560 18813 1595 18847
rect 1629 18813 1664 18847
rect 1698 18813 1733 18847
rect 1767 18813 1802 18847
rect 1836 18813 1871 18847
rect 1905 18813 1940 18847
rect 1974 18813 2009 18847
rect 2043 18813 2078 18847
rect 2112 18813 2147 18847
rect 2181 18813 2216 18847
rect 2250 18813 2285 18847
rect 2319 18813 2354 18847
rect 2388 18813 2423 18847
rect 2457 18813 2492 18847
rect 2526 18813 2561 18847
rect 2595 18813 2630 18847
rect 2664 18813 2699 18847
rect 2733 18813 2768 18847
rect 2802 18813 2837 18847
rect 2871 18813 2906 18847
rect 2940 18813 2975 18847
rect 3009 18813 3044 18847
rect 3078 18813 3113 18847
rect 3147 18813 3182 18847
rect 3216 18813 3251 18847
rect 3285 18813 3320 18847
rect 3354 18813 3389 18847
rect 3423 18813 3458 18847
rect 3492 18813 3527 18847
rect 3561 18813 3596 18847
rect -41 18779 3596 18813
rect -41 18745 77 18779
rect 111 18745 146 18779
rect 180 18745 215 18779
rect 249 18745 284 18779
rect 318 18745 353 18779
rect 387 18745 422 18779
rect 456 18745 491 18779
rect 525 18745 560 18779
rect 594 18745 629 18779
rect 663 18745 698 18779
rect 732 18745 767 18779
rect 801 18745 836 18779
rect 870 18745 905 18779
rect 939 18745 974 18779
rect 1008 18745 1043 18779
rect 1077 18745 1112 18779
rect 1146 18745 1181 18779
rect 1215 18745 1250 18779
rect 1284 18745 1319 18779
rect 1353 18745 1388 18779
rect 1422 18745 1457 18779
rect 1491 18745 1526 18779
rect 1560 18745 1595 18779
rect 1629 18745 1664 18779
rect 1698 18745 1733 18779
rect 1767 18745 1802 18779
rect 1836 18745 1871 18779
rect 1905 18745 1940 18779
rect 1974 18745 2009 18779
rect 2043 18745 2078 18779
rect 2112 18745 2147 18779
rect 2181 18745 2216 18779
rect 2250 18745 2285 18779
rect 2319 18745 2354 18779
rect 2388 18745 2423 18779
rect 2457 18745 2492 18779
rect 2526 18745 2561 18779
rect 2595 18745 2630 18779
rect 2664 18745 2699 18779
rect 2733 18745 2768 18779
rect 2802 18745 2837 18779
rect 2871 18745 2906 18779
rect 2940 18745 2975 18779
rect 3009 18745 3044 18779
rect 3078 18745 3113 18779
rect 3147 18745 3182 18779
rect 3216 18745 3251 18779
rect 3285 18745 3320 18779
rect 3354 18745 3389 18779
rect 3423 18745 3458 18779
rect 3492 18745 3527 18779
rect 3561 18745 3596 18779
rect -41 18711 3596 18745
rect -41 18677 77 18711
rect 111 18677 146 18711
rect 180 18677 215 18711
rect 249 18677 284 18711
rect 318 18677 353 18711
rect 387 18677 422 18711
rect 456 18677 491 18711
rect 525 18677 560 18711
rect 594 18677 629 18711
rect 663 18677 698 18711
rect 732 18677 767 18711
rect 801 18677 836 18711
rect 870 18677 905 18711
rect 939 18677 974 18711
rect 1008 18677 1043 18711
rect 1077 18677 1112 18711
rect 1146 18677 1181 18711
rect 1215 18677 1250 18711
rect 1284 18677 1319 18711
rect 1353 18677 1388 18711
rect 1422 18677 1457 18711
rect 1491 18677 1526 18711
rect 1560 18677 1595 18711
rect 1629 18677 1664 18711
rect 1698 18677 1733 18711
rect 1767 18677 1802 18711
rect 1836 18677 1871 18711
rect 1905 18677 1940 18711
rect 1974 18677 2009 18711
rect 2043 18677 2078 18711
rect 2112 18677 2147 18711
rect 2181 18677 2216 18711
rect 2250 18677 2285 18711
rect 2319 18677 2354 18711
rect 2388 18677 2423 18711
rect 2457 18677 2492 18711
rect 2526 18677 2561 18711
rect 2595 18677 2630 18711
rect 2664 18677 2699 18711
rect 2733 18677 2768 18711
rect 2802 18677 2837 18711
rect 2871 18677 2906 18711
rect 2940 18677 2975 18711
rect 3009 18677 3044 18711
rect 3078 18677 3113 18711
rect 3147 18677 3182 18711
rect 3216 18677 3251 18711
rect 3285 18677 3320 18711
rect 3354 18677 3389 18711
rect 3423 18677 3458 18711
rect 3492 18677 3527 18711
rect 3561 18677 3596 18711
rect 14850 18677 14952 18915
rect -41 18589 14952 18677
rect 197 18555 221 18589
rect 255 18555 290 18589
rect 324 18555 359 18589
rect 393 18555 427 18589
rect 461 18555 495 18589
rect 529 18555 563 18589
rect 597 18555 631 18589
rect 665 18555 699 18589
rect 733 18555 767 18589
rect 801 18555 835 18589
rect 869 18555 903 18589
rect 937 18555 971 18589
rect 1005 18555 1039 18589
rect 1073 18555 1107 18589
rect 1141 18555 1175 18589
rect 1209 18555 1243 18589
rect 1277 18555 1311 18589
rect 1345 18555 1379 18589
rect 1413 18555 1447 18589
rect 1481 18555 1515 18589
rect 1549 18555 1583 18589
rect 1617 18555 1651 18589
rect 1685 18555 1719 18589
rect 1753 18555 1787 18589
rect 1821 18555 1855 18589
rect 1889 18555 1923 18589
rect 1957 18555 1991 18589
rect 2025 18555 2059 18589
rect 2093 18555 2127 18589
rect 2161 18555 2195 18589
rect 2229 18555 2263 18589
rect 2297 18555 2331 18589
rect 2365 18555 2399 18589
rect 2433 18555 2467 18589
rect 2501 18555 2535 18589
rect 2569 18555 2603 18589
rect 2637 18555 2671 18589
rect 2705 18555 2739 18589
rect 2773 18555 2807 18589
rect 2841 18555 2875 18589
rect 2909 18555 2943 18589
rect 2977 18555 3011 18589
rect 3045 18555 3079 18589
rect 3113 18555 3147 18589
rect 3181 18555 3215 18589
rect 3249 18555 3283 18589
rect 3317 18555 3351 18589
rect 3385 18555 3419 18589
rect 3453 18555 3487 18589
rect 3521 18555 3555 18589
rect 3589 18555 3623 18589
rect 3657 18555 3691 18589
rect 3725 18555 3759 18589
rect 3793 18555 3827 18589
rect 3861 18555 3895 18589
rect 3929 18555 3963 18589
rect 3997 18555 4031 18589
rect 4065 18555 4099 18589
rect 4133 18555 4167 18589
rect 4201 18555 4235 18589
rect 4269 18555 4303 18589
rect 4337 18555 4371 18589
rect 4405 18555 4439 18589
rect 4473 18555 4507 18589
rect 4541 18555 4575 18589
rect 4609 18555 4643 18589
rect 4677 18555 4711 18589
rect 4745 18555 4779 18589
rect 4813 18555 4847 18589
rect 4881 18555 4915 18589
rect 4949 18555 4983 18589
rect 5017 18555 5051 18589
rect 5085 18555 5119 18589
rect 5153 18555 5187 18589
rect 5221 18555 5255 18589
rect 5289 18555 5323 18589
rect 5357 18555 5391 18589
rect 5425 18555 5459 18589
rect 5493 18555 5527 18589
rect 5561 18555 5595 18589
rect 5629 18555 5663 18589
rect 5697 18555 5731 18589
rect 5765 18555 5799 18589
rect 5833 18555 5867 18589
rect 5901 18555 5935 18589
rect 5969 18555 6003 18589
rect 6037 18555 6071 18589
rect 6105 18555 6139 18589
rect 6173 18555 6207 18589
rect 6241 18555 6275 18589
rect 6309 18555 6343 18589
rect 6377 18555 6411 18589
rect 6445 18555 6479 18589
rect 6513 18555 6547 18589
rect 6581 18555 6615 18589
rect 6649 18555 6683 18589
rect 6717 18555 6751 18589
rect 6785 18555 6819 18589
rect 6853 18555 6887 18589
rect 6921 18555 6955 18589
rect 6989 18555 7023 18589
rect 7057 18555 7091 18589
rect 7125 18555 7159 18589
rect 7193 18555 7227 18589
rect 7261 18555 7295 18589
rect 7329 18555 7363 18589
rect 7397 18555 7431 18589
rect 7465 18555 7499 18589
rect 7533 18555 7567 18589
rect 7601 18555 7635 18589
rect 7669 18555 7703 18589
rect 7737 18555 7771 18589
rect 7805 18555 7839 18589
rect 7873 18555 7907 18589
rect 7941 18555 7975 18589
rect 8009 18555 8043 18589
rect 8077 18555 8111 18589
rect 8145 18555 8179 18589
rect 8213 18555 8247 18589
rect 8281 18555 8315 18589
rect 8349 18555 8383 18589
rect 8417 18555 8451 18589
rect 8485 18555 8519 18589
rect 8553 18555 8587 18589
rect 8621 18555 8655 18589
rect 8689 18555 8723 18589
rect 8757 18555 8791 18589
rect 8825 18555 8859 18589
rect 8893 18555 8927 18589
rect 8961 18555 8995 18589
rect 9029 18555 9063 18589
rect 9097 18555 9131 18589
rect 9165 18555 9199 18589
rect 9233 18555 9267 18589
rect 9301 18555 9335 18589
rect 9369 18555 9403 18589
rect 9437 18555 9471 18589
rect 9505 18555 9539 18589
rect 9573 18555 9607 18589
rect 9641 18555 9675 18589
rect 9709 18555 9743 18589
rect 9777 18555 9811 18589
rect 9845 18555 9879 18589
rect 9913 18555 9947 18589
rect 9981 18555 10015 18589
rect 10049 18555 10083 18589
rect 10117 18555 10151 18589
rect 10185 18555 10219 18589
rect 10253 18555 10287 18589
rect 10321 18555 10355 18589
rect 10389 18555 10423 18589
rect 10457 18555 10491 18589
rect 10525 18555 10559 18589
rect 10593 18555 10627 18589
rect 10661 18555 10695 18589
rect 10729 18555 10763 18589
rect 10797 18555 10831 18589
rect 10865 18555 10899 18589
rect 10933 18555 10967 18589
rect 11001 18555 11035 18589
rect 11069 18555 11103 18589
rect 11137 18555 11171 18589
rect 11205 18555 11239 18589
rect 11273 18555 11307 18589
rect 11341 18555 11375 18589
rect 11409 18555 11443 18589
rect 11477 18555 11511 18589
rect 11545 18555 11579 18589
rect 11613 18555 11647 18589
rect 11681 18555 11715 18589
rect 11749 18555 11783 18589
rect 11817 18555 11851 18589
rect 11885 18555 11919 18589
rect 11953 18555 11987 18589
rect 12021 18555 12055 18589
rect 12089 18555 12123 18589
rect 12157 18555 12191 18589
rect 12225 18555 12259 18589
rect 12293 18555 12327 18589
rect 12361 18555 12395 18589
rect 12429 18555 12463 18589
rect 12497 18555 12531 18589
rect 12565 18555 12599 18589
rect 12633 18555 12667 18589
rect 12701 18555 12735 18589
rect 12769 18555 12803 18589
rect 12837 18555 12871 18589
rect 12905 18555 12939 18589
rect 12973 18555 13007 18589
rect 13041 18555 13075 18589
rect 13109 18555 13143 18589
rect 13177 18555 13211 18589
rect 13245 18555 13279 18589
rect 13313 18555 13347 18589
rect 13381 18555 13415 18589
rect 13449 18555 13483 18589
rect 13517 18555 13551 18589
rect 13585 18555 13619 18589
rect 13653 18555 13687 18589
rect 13721 18555 13755 18589
rect 13789 18555 13823 18589
rect 13857 18555 13891 18589
rect 13925 18555 13959 18589
rect 13993 18555 14027 18589
rect 14061 18555 14095 18589
rect 14129 18555 14163 18589
rect 14197 18555 14231 18589
rect 14265 18555 14299 18589
rect 14333 18555 14367 18589
rect 14401 18555 14435 18589
rect 14469 18555 14503 18589
rect 14537 18555 14571 18589
rect 14605 18555 14639 18589
rect 14673 18555 14707 18589
rect 14741 18555 14772 18589
rect 197 18519 14772 18555
rect 197 18485 221 18519
rect 255 18485 290 18519
rect 324 18485 359 18519
rect 393 18485 427 18519
rect 461 18485 495 18519
rect 529 18485 563 18519
rect 597 18485 631 18519
rect 665 18485 699 18519
rect 733 18485 767 18519
rect 801 18485 835 18519
rect 869 18485 903 18519
rect 937 18485 971 18519
rect 1005 18485 1039 18519
rect 1073 18485 1107 18519
rect 1141 18485 1175 18519
rect 1209 18485 1243 18519
rect 1277 18485 1311 18519
rect 1345 18485 1379 18519
rect 1413 18485 1447 18519
rect 1481 18485 1515 18519
rect 1549 18485 1583 18519
rect 1617 18485 1651 18519
rect 1685 18485 1719 18519
rect 1753 18485 1787 18519
rect 1821 18485 1855 18519
rect 1889 18485 1923 18519
rect 1957 18485 1991 18519
rect 2025 18485 2059 18519
rect 2093 18485 2127 18519
rect 2161 18485 2195 18519
rect 2229 18485 2263 18519
rect 2297 18485 2331 18519
rect 2365 18485 2399 18519
rect 2433 18485 2467 18519
rect 2501 18485 2535 18519
rect 2569 18485 2603 18519
rect 2637 18485 2671 18519
rect 2705 18485 2739 18519
rect 2773 18485 2807 18519
rect 2841 18485 2875 18519
rect 2909 18485 2943 18519
rect 2977 18485 3011 18519
rect 3045 18485 3079 18519
rect 3113 18485 3147 18519
rect 3181 18485 3215 18519
rect 3249 18485 3283 18519
rect 3317 18485 3351 18519
rect 3385 18485 3419 18519
rect 3453 18485 3487 18519
rect 3521 18485 3555 18519
rect 3589 18485 3623 18519
rect 3657 18485 3691 18519
rect 3725 18485 3759 18519
rect 3793 18485 3827 18519
rect 3861 18485 3895 18519
rect 3929 18485 3963 18519
rect 3997 18485 4031 18519
rect 4065 18485 4099 18519
rect 4133 18485 4167 18519
rect 4201 18485 4235 18519
rect 4269 18485 4303 18519
rect 4337 18485 4371 18519
rect 4405 18485 4439 18519
rect 4473 18485 4507 18519
rect 4541 18485 4575 18519
rect 4609 18485 4643 18519
rect 4677 18485 4711 18519
rect 4745 18485 4779 18519
rect 4813 18485 4847 18519
rect 4881 18485 4915 18519
rect 4949 18485 4983 18519
rect 5017 18485 5051 18519
rect 5085 18485 5119 18519
rect 5153 18485 5187 18519
rect 5221 18485 5255 18519
rect 5289 18485 5323 18519
rect 5357 18485 5391 18519
rect 5425 18485 5459 18519
rect 5493 18485 5527 18519
rect 5561 18485 5595 18519
rect 5629 18485 5663 18519
rect 5697 18485 5731 18519
rect 5765 18485 5799 18519
rect 5833 18485 5867 18519
rect 5901 18485 5935 18519
rect 5969 18485 6003 18519
rect 6037 18485 6071 18519
rect 6105 18485 6139 18519
rect 6173 18485 6207 18519
rect 6241 18485 6275 18519
rect 6309 18485 6343 18519
rect 6377 18485 6411 18519
rect 6445 18485 6479 18519
rect 6513 18485 6547 18519
rect 6581 18485 6615 18519
rect 6649 18485 6683 18519
rect 6717 18485 6751 18519
rect 6785 18485 6819 18519
rect 6853 18485 6887 18519
rect 6921 18485 6955 18519
rect 6989 18485 7023 18519
rect 7057 18485 7091 18519
rect 7125 18485 7159 18519
rect 7193 18485 7227 18519
rect 7261 18485 7295 18519
rect 7329 18485 7363 18519
rect 7397 18485 7431 18519
rect 7465 18485 7499 18519
rect 7533 18485 7567 18519
rect 7601 18485 7635 18519
rect 7669 18485 7703 18519
rect 7737 18485 7771 18519
rect 7805 18485 7839 18519
rect 7873 18485 7907 18519
rect 7941 18485 7975 18519
rect 8009 18485 8043 18519
rect 8077 18485 8111 18519
rect 8145 18485 8179 18519
rect 8213 18485 8247 18519
rect 8281 18485 8315 18519
rect 8349 18485 8383 18519
rect 8417 18485 8451 18519
rect 8485 18485 8519 18519
rect 8553 18485 8587 18519
rect 8621 18485 8655 18519
rect 8689 18485 8723 18519
rect 8757 18485 8791 18519
rect 8825 18485 8859 18519
rect 8893 18485 8927 18519
rect 8961 18485 8995 18519
rect 9029 18485 9063 18519
rect 9097 18485 9131 18519
rect 9165 18485 9199 18519
rect 9233 18485 9267 18519
rect 9301 18485 9335 18519
rect 9369 18485 9403 18519
rect 9437 18485 9471 18519
rect 9505 18485 9539 18519
rect 9573 18485 9607 18519
rect 9641 18485 9675 18519
rect 9709 18485 9743 18519
rect 9777 18485 9811 18519
rect 9845 18485 9879 18519
rect 9913 18485 9947 18519
rect 9981 18485 10015 18519
rect 10049 18485 10083 18519
rect 10117 18485 10151 18519
rect 10185 18485 10219 18519
rect 10253 18485 10287 18519
rect 10321 18485 10355 18519
rect 10389 18485 10423 18519
rect 10457 18485 10491 18519
rect 10525 18485 10559 18519
rect 10593 18485 10627 18519
rect 10661 18485 10695 18519
rect 10729 18485 10763 18519
rect 10797 18485 10831 18519
rect 10865 18485 10899 18519
rect 10933 18485 10967 18519
rect 11001 18485 11035 18519
rect 11069 18485 11103 18519
rect 11137 18485 11171 18519
rect 11205 18485 11239 18519
rect 11273 18485 11307 18519
rect 11341 18485 11375 18519
rect 11409 18485 11443 18519
rect 11477 18485 11511 18519
rect 11545 18485 11579 18519
rect 11613 18485 11647 18519
rect 11681 18485 11715 18519
rect 11749 18485 11783 18519
rect 11817 18485 11851 18519
rect 11885 18485 11919 18519
rect 11953 18485 11987 18519
rect 12021 18485 12055 18519
rect 12089 18485 12123 18519
rect 12157 18485 12191 18519
rect 12225 18485 12259 18519
rect 12293 18485 12327 18519
rect 12361 18485 12395 18519
rect 12429 18485 12463 18519
rect 12497 18485 12531 18519
rect 12565 18485 12599 18519
rect 12633 18485 12667 18519
rect 12701 18485 12735 18519
rect 12769 18485 12803 18519
rect 12837 18485 12871 18519
rect 12905 18485 12939 18519
rect 12973 18485 13007 18519
rect 13041 18485 13075 18519
rect 13109 18485 13143 18519
rect 13177 18485 13211 18519
rect 13245 18485 13279 18519
rect 13313 18485 13347 18519
rect 13381 18485 13415 18519
rect 13449 18485 13483 18519
rect 13517 18485 13551 18519
rect 13585 18485 13619 18519
rect 13653 18485 13687 18519
rect 13721 18485 13755 18519
rect 13789 18485 13823 18519
rect 13857 18485 13891 18519
rect 13925 18485 13959 18519
rect 13993 18485 14027 18519
rect 14061 18485 14095 18519
rect 14129 18485 14163 18519
rect 14197 18485 14231 18519
rect 14265 18485 14299 18519
rect 14333 18485 14367 18519
rect 14401 18485 14435 18519
rect 14469 18485 14503 18519
rect 14537 18485 14571 18519
rect 14605 18485 14639 18519
rect 14673 18485 14707 18519
rect 14741 18485 14772 18519
rect 197 18449 14772 18485
rect 197 18415 221 18449
rect 255 18415 290 18449
rect 324 18415 359 18449
rect 393 18415 427 18449
rect 461 18415 495 18449
rect 529 18415 563 18449
rect 597 18415 631 18449
rect 665 18415 699 18449
rect 733 18415 767 18449
rect 801 18415 835 18449
rect 869 18415 903 18449
rect 937 18415 971 18449
rect 1005 18415 1039 18449
rect 1073 18415 1107 18449
rect 1141 18415 1175 18449
rect 1209 18415 1243 18449
rect 1277 18415 1311 18449
rect 1345 18415 1379 18449
rect 1413 18415 1447 18449
rect 1481 18415 1515 18449
rect 1549 18415 1583 18449
rect 1617 18415 1651 18449
rect 1685 18415 1719 18449
rect 1753 18415 1787 18449
rect 1821 18415 1855 18449
rect 1889 18415 1923 18449
rect 1957 18415 1991 18449
rect 2025 18415 2059 18449
rect 2093 18415 2127 18449
rect 2161 18415 2195 18449
rect 2229 18415 2263 18449
rect 2297 18415 2331 18449
rect 2365 18415 2399 18449
rect 2433 18415 2467 18449
rect 2501 18415 2535 18449
rect 2569 18415 2603 18449
rect 2637 18415 2671 18449
rect 2705 18415 2739 18449
rect 2773 18415 2807 18449
rect 2841 18415 2875 18449
rect 2909 18415 2943 18449
rect 2977 18415 3011 18449
rect 3045 18415 3079 18449
rect 3113 18415 3147 18449
rect 3181 18415 3215 18449
rect 3249 18415 3283 18449
rect 3317 18415 3351 18449
rect 3385 18415 3419 18449
rect 3453 18415 3487 18449
rect 3521 18415 3555 18449
rect 3589 18415 3623 18449
rect 3657 18415 3691 18449
rect 3725 18415 3759 18449
rect 3793 18415 3827 18449
rect 3861 18415 3895 18449
rect 3929 18415 3963 18449
rect 3997 18415 4031 18449
rect 4065 18415 4099 18449
rect 4133 18415 4167 18449
rect 4201 18415 4235 18449
rect 4269 18415 4303 18449
rect 4337 18415 4371 18449
rect 4405 18415 4439 18449
rect 4473 18415 4507 18449
rect 4541 18415 4575 18449
rect 4609 18415 4643 18449
rect 4677 18415 4711 18449
rect 4745 18415 4779 18449
rect 4813 18415 4847 18449
rect 4881 18415 4915 18449
rect 4949 18415 4983 18449
rect 5017 18415 5051 18449
rect 5085 18415 5119 18449
rect 5153 18415 5187 18449
rect 5221 18415 5255 18449
rect 5289 18415 5323 18449
rect 5357 18415 5391 18449
rect 5425 18415 5459 18449
rect 5493 18415 5527 18449
rect 5561 18415 5595 18449
rect 5629 18415 5663 18449
rect 5697 18415 5731 18449
rect 5765 18415 5799 18449
rect 5833 18415 5867 18449
rect 5901 18415 5935 18449
rect 5969 18415 6003 18449
rect 6037 18415 6071 18449
rect 6105 18415 6139 18449
rect 6173 18415 6207 18449
rect 6241 18415 6275 18449
rect 6309 18415 6343 18449
rect 6377 18415 6411 18449
rect 6445 18415 6479 18449
rect 6513 18415 6547 18449
rect 6581 18415 6615 18449
rect 6649 18415 6683 18449
rect 6717 18415 6751 18449
rect 6785 18415 6819 18449
rect 6853 18415 6887 18449
rect 6921 18415 6955 18449
rect 6989 18415 7023 18449
rect 7057 18415 7091 18449
rect 7125 18415 7159 18449
rect 7193 18415 7227 18449
rect 7261 18415 7295 18449
rect 7329 18415 7363 18449
rect 7397 18415 7431 18449
rect 7465 18415 7499 18449
rect 7533 18415 7567 18449
rect 7601 18415 7635 18449
rect 7669 18415 7703 18449
rect 7737 18415 7771 18449
rect 7805 18415 7839 18449
rect 7873 18415 7907 18449
rect 7941 18415 7975 18449
rect 8009 18415 8043 18449
rect 8077 18415 8111 18449
rect 8145 18415 8179 18449
rect 8213 18415 8247 18449
rect 8281 18415 8315 18449
rect 8349 18415 8383 18449
rect 8417 18415 8451 18449
rect 8485 18415 8519 18449
rect 8553 18415 8587 18449
rect 8621 18415 8655 18449
rect 8689 18415 8723 18449
rect 8757 18415 8791 18449
rect 8825 18415 8859 18449
rect 8893 18415 8927 18449
rect 8961 18415 8995 18449
rect 9029 18415 9063 18449
rect 9097 18415 9131 18449
rect 9165 18415 9199 18449
rect 9233 18415 9267 18449
rect 9301 18415 9335 18449
rect 9369 18415 9403 18449
rect 9437 18415 9471 18449
rect 9505 18415 9539 18449
rect 9573 18415 9607 18449
rect 9641 18415 9675 18449
rect 9709 18415 9743 18449
rect 9777 18415 9811 18449
rect 9845 18415 9879 18449
rect 9913 18415 9947 18449
rect 9981 18415 10015 18449
rect 10049 18415 10083 18449
rect 10117 18415 10151 18449
rect 10185 18415 10219 18449
rect 10253 18415 10287 18449
rect 10321 18415 10355 18449
rect 10389 18415 10423 18449
rect 10457 18415 10491 18449
rect 10525 18415 10559 18449
rect 10593 18415 10627 18449
rect 10661 18415 10695 18449
rect 10729 18415 10763 18449
rect 10797 18415 10831 18449
rect 10865 18415 10899 18449
rect 10933 18415 10967 18449
rect 11001 18415 11035 18449
rect 11069 18415 11103 18449
rect 11137 18415 11171 18449
rect 11205 18415 11239 18449
rect 11273 18415 11307 18449
rect 11341 18415 11375 18449
rect 11409 18415 11443 18449
rect 11477 18415 11511 18449
rect 11545 18415 11579 18449
rect 11613 18415 11647 18449
rect 11681 18415 11715 18449
rect 11749 18415 11783 18449
rect 11817 18415 11851 18449
rect 11885 18415 11919 18449
rect 11953 18415 11987 18449
rect 12021 18415 12055 18449
rect 12089 18415 12123 18449
rect 12157 18415 12191 18449
rect 12225 18415 12259 18449
rect 12293 18415 12327 18449
rect 12361 18415 12395 18449
rect 12429 18415 12463 18449
rect 12497 18415 12531 18449
rect 12565 18415 12599 18449
rect 12633 18415 12667 18449
rect 12701 18415 12735 18449
rect 12769 18415 12803 18449
rect 12837 18415 12871 18449
rect 12905 18415 12939 18449
rect 12973 18415 13007 18449
rect 13041 18415 13075 18449
rect 13109 18415 13143 18449
rect 13177 18415 13211 18449
rect 13245 18415 13279 18449
rect 13313 18415 13347 18449
rect 13381 18415 13415 18449
rect 13449 18415 13483 18449
rect 13517 18415 13551 18449
rect 13585 18415 13619 18449
rect 13653 18415 13687 18449
rect 13721 18415 13755 18449
rect 13789 18415 13823 18449
rect 13857 18415 13891 18449
rect 13925 18415 13959 18449
rect 13993 18415 14027 18449
rect 14061 18415 14095 18449
rect 14129 18415 14163 18449
rect 14197 18415 14231 18449
rect 14265 18415 14299 18449
rect 14333 18415 14367 18449
rect 14401 18415 14435 18449
rect 14469 18415 14503 18449
rect 14537 18415 14571 18449
rect 14605 18415 14639 18449
rect 14673 18415 14707 18449
rect 14741 18415 14772 18449
rect 197 18382 14772 18415
rect 197 18348 209 18382
rect 243 18379 282 18382
rect 316 18379 355 18382
rect 389 18379 428 18382
rect 462 18379 501 18382
rect 535 18379 574 18382
rect 608 18379 647 18382
rect 681 18379 720 18382
rect 754 18379 793 18382
rect 827 18379 866 18382
rect 900 18379 939 18382
rect 973 18379 1012 18382
rect 1046 18379 1085 18382
rect 1119 18379 1158 18382
rect 1192 18379 1231 18382
rect 1265 18379 1304 18382
rect 1338 18379 1377 18382
rect 1411 18379 1450 18382
rect 1484 18379 1523 18382
rect 1557 18379 1596 18382
rect 1630 18379 1669 18382
rect 1703 18379 1742 18382
rect 1776 18379 1815 18382
rect 1849 18379 1888 18382
rect 1922 18379 1961 18382
rect 1995 18379 2034 18382
rect 2068 18379 2107 18382
rect 2141 18379 2180 18382
rect 2214 18379 2253 18382
rect 2287 18379 2326 18382
rect 2360 18379 2399 18382
rect 2433 18379 2472 18382
rect 2506 18379 2545 18382
rect 2579 18379 2618 18382
rect 2652 18379 2691 18382
rect 2725 18379 2764 18382
rect 2798 18379 2837 18382
rect 2871 18379 2910 18382
rect 2944 18379 2983 18382
rect 3017 18379 3056 18382
rect 3090 18379 3129 18382
rect 3163 18379 3202 18382
rect 3236 18379 3275 18382
rect 3309 18379 3348 18382
rect 3382 18379 3421 18382
rect 3455 18379 3494 18382
rect 3528 18379 3566 18382
rect 3600 18379 3638 18382
rect 3672 18379 3710 18382
rect 3744 18379 3782 18382
rect 3816 18379 3854 18382
rect 3888 18379 3926 18382
rect 3960 18379 3998 18382
rect 4032 18379 4070 18382
rect 4104 18379 4142 18382
rect 4176 18379 4214 18382
rect 4248 18379 4286 18382
rect 4320 18379 4358 18382
rect 4392 18379 4430 18382
rect 4464 18379 4502 18382
rect 4536 18379 4574 18382
rect 4608 18379 4646 18382
rect 4680 18379 4718 18382
rect 4752 18379 4790 18382
rect 4824 18379 4862 18382
rect 4896 18379 4934 18382
rect 4968 18379 5006 18382
rect 5040 18379 5078 18382
rect 5112 18379 5150 18382
rect 5184 18379 5222 18382
rect 5256 18379 5294 18382
rect 5328 18379 5366 18382
rect 5400 18379 5438 18382
rect 5472 18379 5510 18382
rect 5544 18379 5582 18382
rect 5616 18379 5654 18382
rect 5688 18379 5726 18382
rect 5760 18379 5798 18382
rect 5832 18379 5870 18382
rect 5904 18379 5942 18382
rect 5976 18379 6014 18382
rect 6048 18379 6086 18382
rect 6120 18379 6158 18382
rect 6192 18379 6230 18382
rect 6264 18379 6302 18382
rect 6336 18379 6374 18382
rect 6408 18379 6446 18382
rect 6480 18379 6518 18382
rect 6552 18379 6590 18382
rect 6624 18379 6662 18382
rect 6696 18379 6734 18382
rect 6768 18379 6806 18382
rect 6840 18379 6878 18382
rect 6912 18379 6950 18382
rect 6984 18379 7022 18382
rect 7056 18379 7094 18382
rect 7128 18379 7166 18382
rect 7200 18379 7238 18382
rect 7272 18379 7310 18382
rect 7344 18379 7382 18382
rect 7416 18379 7454 18382
rect 7488 18379 7526 18382
rect 7560 18379 7598 18382
rect 7632 18379 7670 18382
rect 7704 18379 7742 18382
rect 7776 18379 7814 18382
rect 7848 18379 7886 18382
rect 7920 18379 7958 18382
rect 7992 18379 8030 18382
rect 8064 18379 8102 18382
rect 8136 18379 8174 18382
rect 8208 18379 8246 18382
rect 8280 18379 8318 18382
rect 8352 18379 8390 18382
rect 8424 18379 8462 18382
rect 8496 18379 8534 18382
rect 8568 18379 8606 18382
rect 8640 18379 8678 18382
rect 8712 18379 8750 18382
rect 8784 18379 8822 18382
rect 8856 18379 8894 18382
rect 8928 18379 8966 18382
rect 9000 18379 9038 18382
rect 9072 18379 9110 18382
rect 9144 18379 9182 18382
rect 9216 18379 9254 18382
rect 9288 18379 9326 18382
rect 9360 18379 9398 18382
rect 9432 18379 9470 18382
rect 9504 18379 9542 18382
rect 9576 18379 9614 18382
rect 9648 18379 9686 18382
rect 9720 18379 9758 18382
rect 9792 18379 9830 18382
rect 9864 18379 9902 18382
rect 9936 18379 9974 18382
rect 10008 18379 10046 18382
rect 10080 18379 10118 18382
rect 10152 18379 10190 18382
rect 10224 18379 10262 18382
rect 10296 18379 10334 18382
rect 10368 18379 10406 18382
rect 10440 18379 10478 18382
rect 10512 18379 10550 18382
rect 10584 18379 10622 18382
rect 10656 18379 10694 18382
rect 10728 18379 10766 18382
rect 10800 18379 10838 18382
rect 10872 18379 10910 18382
rect 10944 18379 10982 18382
rect 11016 18379 11054 18382
rect 11088 18379 11126 18382
rect 11160 18379 11198 18382
rect 11232 18379 11270 18382
rect 11304 18379 11342 18382
rect 11376 18379 11414 18382
rect 11448 18379 11486 18382
rect 11520 18379 11558 18382
rect 11592 18379 11630 18382
rect 11664 18379 11702 18382
rect 11736 18379 11774 18382
rect 11808 18379 11846 18382
rect 11880 18379 11918 18382
rect 11952 18379 11990 18382
rect 12024 18379 12062 18382
rect 12096 18379 12134 18382
rect 12168 18379 12206 18382
rect 12240 18379 12278 18382
rect 12312 18379 12350 18382
rect 12384 18379 12422 18382
rect 12456 18379 12494 18382
rect 12528 18379 12566 18382
rect 12600 18379 12638 18382
rect 12672 18379 12710 18382
rect 12744 18379 12782 18382
rect 12816 18379 12854 18382
rect 12888 18379 12926 18382
rect 12960 18379 12998 18382
rect 13032 18379 13070 18382
rect 13104 18379 13142 18382
rect 13176 18379 13214 18382
rect 13248 18379 13286 18382
rect 13320 18379 13358 18382
rect 13392 18379 13430 18382
rect 13464 18379 13502 18382
rect 13536 18379 13574 18382
rect 13608 18379 13646 18382
rect 13680 18379 13718 18382
rect 13752 18379 13790 18382
rect 13824 18379 13862 18382
rect 13896 18379 13934 18382
rect 13968 18379 14006 18382
rect 14040 18379 14078 18382
rect 14112 18379 14150 18382
rect 14184 18379 14222 18382
rect 14256 18379 14294 18382
rect 14328 18379 14366 18382
rect 14400 18379 14438 18382
rect 14472 18379 14510 18382
rect 14544 18379 14582 18382
rect 14616 18379 14654 18382
rect 14688 18379 14726 18382
rect 255 18348 282 18379
rect 324 18348 355 18379
rect 197 18345 221 18348
rect 255 18345 290 18348
rect 324 18345 359 18348
rect 393 18345 427 18379
rect 462 18348 495 18379
rect 535 18348 563 18379
rect 608 18348 631 18379
rect 681 18348 699 18379
rect 754 18348 767 18379
rect 827 18348 835 18379
rect 900 18348 903 18379
rect 461 18345 495 18348
rect 529 18345 563 18348
rect 597 18345 631 18348
rect 665 18345 699 18348
rect 733 18345 767 18348
rect 801 18345 835 18348
rect 869 18345 903 18348
rect 937 18348 939 18379
rect 1005 18348 1012 18379
rect 1073 18348 1085 18379
rect 1141 18348 1158 18379
rect 1209 18348 1231 18379
rect 1277 18348 1304 18379
rect 1345 18348 1377 18379
rect 937 18345 971 18348
rect 1005 18345 1039 18348
rect 1073 18345 1107 18348
rect 1141 18345 1175 18348
rect 1209 18345 1243 18348
rect 1277 18345 1311 18348
rect 1345 18345 1379 18348
rect 1413 18345 1447 18379
rect 1484 18348 1515 18379
rect 1557 18348 1583 18379
rect 1630 18348 1651 18379
rect 1703 18348 1719 18379
rect 1776 18348 1787 18379
rect 1849 18348 1855 18379
rect 1922 18348 1923 18379
rect 1481 18345 1515 18348
rect 1549 18345 1583 18348
rect 1617 18345 1651 18348
rect 1685 18345 1719 18348
rect 1753 18345 1787 18348
rect 1821 18345 1855 18348
rect 1889 18345 1923 18348
rect 1957 18348 1961 18379
rect 2025 18348 2034 18379
rect 2093 18348 2107 18379
rect 2161 18348 2180 18379
rect 2229 18348 2253 18379
rect 2297 18348 2326 18379
rect 1957 18345 1991 18348
rect 2025 18345 2059 18348
rect 2093 18345 2127 18348
rect 2161 18345 2195 18348
rect 2229 18345 2263 18348
rect 2297 18345 2331 18348
rect 2365 18345 2399 18379
rect 2433 18345 2467 18379
rect 2506 18348 2535 18379
rect 2579 18348 2603 18379
rect 2652 18348 2671 18379
rect 2725 18348 2739 18379
rect 2798 18348 2807 18379
rect 2871 18348 2875 18379
rect 2501 18345 2535 18348
rect 2569 18345 2603 18348
rect 2637 18345 2671 18348
rect 2705 18345 2739 18348
rect 2773 18345 2807 18348
rect 2841 18345 2875 18348
rect 2909 18348 2910 18379
rect 2977 18348 2983 18379
rect 3045 18348 3056 18379
rect 3113 18348 3129 18379
rect 3181 18348 3202 18379
rect 3249 18348 3275 18379
rect 3317 18348 3348 18379
rect 2909 18345 2943 18348
rect 2977 18345 3011 18348
rect 3045 18345 3079 18348
rect 3113 18345 3147 18348
rect 3181 18345 3215 18348
rect 3249 18345 3283 18348
rect 3317 18345 3351 18348
rect 3385 18345 3419 18379
rect 3455 18348 3487 18379
rect 3528 18348 3555 18379
rect 3600 18348 3623 18379
rect 3672 18348 3691 18379
rect 3744 18348 3759 18379
rect 3816 18348 3827 18379
rect 3888 18348 3895 18379
rect 3960 18348 3963 18379
rect 3453 18345 3487 18348
rect 3521 18345 3555 18348
rect 3589 18345 3623 18348
rect 3657 18345 3691 18348
rect 3725 18345 3759 18348
rect 3793 18345 3827 18348
rect 3861 18345 3895 18348
rect 3929 18345 3963 18348
rect 3997 18348 3998 18379
rect 4065 18348 4070 18379
rect 4133 18348 4142 18379
rect 4201 18348 4214 18379
rect 4269 18348 4286 18379
rect 4337 18348 4358 18379
rect 4405 18348 4430 18379
rect 4473 18348 4502 18379
rect 4541 18348 4574 18379
rect 3997 18345 4031 18348
rect 4065 18345 4099 18348
rect 4133 18345 4167 18348
rect 4201 18345 4235 18348
rect 4269 18345 4303 18348
rect 4337 18345 4371 18348
rect 4405 18345 4439 18348
rect 4473 18345 4507 18348
rect 4541 18345 4575 18348
rect 4609 18345 4643 18379
rect 4680 18348 4711 18379
rect 4752 18348 4779 18379
rect 4824 18348 4847 18379
rect 4896 18348 4915 18379
rect 4968 18348 4983 18379
rect 5040 18348 5051 18379
rect 5112 18348 5119 18379
rect 5184 18348 5187 18379
rect 4677 18345 4711 18348
rect 4745 18345 4779 18348
rect 4813 18345 4847 18348
rect 4881 18345 4915 18348
rect 4949 18345 4983 18348
rect 5017 18345 5051 18348
rect 5085 18345 5119 18348
rect 5153 18345 5187 18348
rect 5221 18348 5222 18379
rect 5289 18348 5294 18379
rect 5357 18348 5366 18379
rect 5425 18348 5438 18379
rect 5493 18348 5510 18379
rect 5561 18348 5582 18379
rect 5629 18348 5654 18379
rect 5697 18348 5726 18379
rect 5765 18348 5798 18379
rect 5221 18345 5255 18348
rect 5289 18345 5323 18348
rect 5357 18345 5391 18348
rect 5425 18345 5459 18348
rect 5493 18345 5527 18348
rect 5561 18345 5595 18348
rect 5629 18345 5663 18348
rect 5697 18345 5731 18348
rect 5765 18345 5799 18348
rect 5833 18345 5867 18379
rect 5904 18348 5935 18379
rect 5976 18348 6003 18379
rect 6048 18348 6071 18379
rect 6120 18348 6139 18379
rect 6192 18348 6207 18379
rect 6264 18348 6275 18379
rect 6336 18348 6343 18379
rect 6408 18348 6411 18379
rect 5901 18345 5935 18348
rect 5969 18345 6003 18348
rect 6037 18345 6071 18348
rect 6105 18345 6139 18348
rect 6173 18345 6207 18348
rect 6241 18345 6275 18348
rect 6309 18345 6343 18348
rect 6377 18345 6411 18348
rect 6445 18348 6446 18379
rect 6513 18348 6518 18379
rect 6581 18348 6590 18379
rect 6649 18348 6662 18379
rect 6717 18348 6734 18379
rect 6785 18348 6806 18379
rect 6853 18348 6878 18379
rect 6921 18348 6950 18379
rect 6989 18348 7022 18379
rect 6445 18345 6479 18348
rect 6513 18345 6547 18348
rect 6581 18345 6615 18348
rect 6649 18345 6683 18348
rect 6717 18345 6751 18348
rect 6785 18345 6819 18348
rect 6853 18345 6887 18348
rect 6921 18345 6955 18348
rect 6989 18345 7023 18348
rect 7057 18345 7091 18379
rect 7128 18348 7159 18379
rect 7200 18348 7227 18379
rect 7272 18348 7295 18379
rect 7344 18348 7363 18379
rect 7416 18348 7431 18379
rect 7488 18348 7499 18379
rect 7560 18348 7567 18379
rect 7632 18348 7635 18379
rect 7125 18345 7159 18348
rect 7193 18345 7227 18348
rect 7261 18345 7295 18348
rect 7329 18345 7363 18348
rect 7397 18345 7431 18348
rect 7465 18345 7499 18348
rect 7533 18345 7567 18348
rect 7601 18345 7635 18348
rect 7669 18348 7670 18379
rect 7737 18348 7742 18379
rect 7805 18348 7814 18379
rect 7873 18348 7886 18379
rect 7941 18348 7958 18379
rect 8009 18348 8030 18379
rect 8077 18348 8102 18379
rect 8145 18348 8174 18379
rect 8213 18348 8246 18379
rect 7669 18345 7703 18348
rect 7737 18345 7771 18348
rect 7805 18345 7839 18348
rect 7873 18345 7907 18348
rect 7941 18345 7975 18348
rect 8009 18345 8043 18348
rect 8077 18345 8111 18348
rect 8145 18345 8179 18348
rect 8213 18345 8247 18348
rect 8281 18345 8315 18379
rect 8352 18348 8383 18379
rect 8424 18348 8451 18379
rect 8496 18348 8519 18379
rect 8568 18348 8587 18379
rect 8640 18348 8655 18379
rect 8712 18348 8723 18379
rect 8784 18348 8791 18379
rect 8856 18348 8859 18379
rect 8349 18345 8383 18348
rect 8417 18345 8451 18348
rect 8485 18345 8519 18348
rect 8553 18345 8587 18348
rect 8621 18345 8655 18348
rect 8689 18345 8723 18348
rect 8757 18345 8791 18348
rect 8825 18345 8859 18348
rect 8893 18348 8894 18379
rect 8961 18348 8966 18379
rect 9029 18348 9038 18379
rect 9097 18348 9110 18379
rect 9165 18348 9182 18379
rect 9233 18348 9254 18379
rect 9301 18348 9326 18379
rect 9369 18348 9398 18379
rect 9437 18348 9470 18379
rect 8893 18345 8927 18348
rect 8961 18345 8995 18348
rect 9029 18345 9063 18348
rect 9097 18345 9131 18348
rect 9165 18345 9199 18348
rect 9233 18345 9267 18348
rect 9301 18345 9335 18348
rect 9369 18345 9403 18348
rect 9437 18345 9471 18348
rect 9505 18345 9539 18379
rect 9576 18348 9607 18379
rect 9648 18348 9675 18379
rect 9720 18348 9743 18379
rect 9792 18348 9811 18379
rect 9864 18348 9879 18379
rect 9936 18348 9947 18379
rect 10008 18348 10015 18379
rect 10080 18348 10083 18379
rect 9573 18345 9607 18348
rect 9641 18345 9675 18348
rect 9709 18345 9743 18348
rect 9777 18345 9811 18348
rect 9845 18345 9879 18348
rect 9913 18345 9947 18348
rect 9981 18345 10015 18348
rect 10049 18345 10083 18348
rect 10117 18348 10118 18379
rect 10185 18348 10190 18379
rect 10253 18348 10262 18379
rect 10321 18348 10334 18379
rect 10389 18348 10406 18379
rect 10457 18348 10478 18379
rect 10525 18348 10550 18379
rect 10593 18348 10622 18379
rect 10661 18348 10694 18379
rect 10117 18345 10151 18348
rect 10185 18345 10219 18348
rect 10253 18345 10287 18348
rect 10321 18345 10355 18348
rect 10389 18345 10423 18348
rect 10457 18345 10491 18348
rect 10525 18345 10559 18348
rect 10593 18345 10627 18348
rect 10661 18345 10695 18348
rect 10729 18345 10763 18379
rect 10800 18348 10831 18379
rect 10872 18348 10899 18379
rect 10944 18348 10967 18379
rect 11016 18348 11035 18379
rect 11088 18348 11103 18379
rect 11160 18348 11171 18379
rect 11232 18348 11239 18379
rect 11304 18348 11307 18379
rect 10797 18345 10831 18348
rect 10865 18345 10899 18348
rect 10933 18345 10967 18348
rect 11001 18345 11035 18348
rect 11069 18345 11103 18348
rect 11137 18345 11171 18348
rect 11205 18345 11239 18348
rect 11273 18345 11307 18348
rect 11341 18348 11342 18379
rect 11409 18348 11414 18379
rect 11477 18348 11486 18379
rect 11545 18348 11558 18379
rect 11613 18348 11630 18379
rect 11681 18348 11702 18379
rect 11749 18348 11774 18379
rect 11817 18348 11846 18379
rect 11885 18348 11918 18379
rect 11341 18345 11375 18348
rect 11409 18345 11443 18348
rect 11477 18345 11511 18348
rect 11545 18345 11579 18348
rect 11613 18345 11647 18348
rect 11681 18345 11715 18348
rect 11749 18345 11783 18348
rect 11817 18345 11851 18348
rect 11885 18345 11919 18348
rect 11953 18345 11987 18379
rect 12024 18348 12055 18379
rect 12096 18348 12123 18379
rect 12168 18348 12191 18379
rect 12240 18348 12259 18379
rect 12312 18348 12327 18379
rect 12384 18348 12395 18379
rect 12456 18348 12463 18379
rect 12528 18348 12531 18379
rect 12021 18345 12055 18348
rect 12089 18345 12123 18348
rect 12157 18345 12191 18348
rect 12225 18345 12259 18348
rect 12293 18345 12327 18348
rect 12361 18345 12395 18348
rect 12429 18345 12463 18348
rect 12497 18345 12531 18348
rect 12565 18348 12566 18379
rect 12633 18348 12638 18379
rect 12701 18348 12710 18379
rect 12769 18348 12782 18379
rect 12837 18348 12854 18379
rect 12905 18348 12926 18379
rect 12973 18348 12998 18379
rect 13041 18348 13070 18379
rect 13109 18348 13142 18379
rect 12565 18345 12599 18348
rect 12633 18345 12667 18348
rect 12701 18345 12735 18348
rect 12769 18345 12803 18348
rect 12837 18345 12871 18348
rect 12905 18345 12939 18348
rect 12973 18345 13007 18348
rect 13041 18345 13075 18348
rect 13109 18345 13143 18348
rect 13177 18345 13211 18379
rect 13248 18348 13279 18379
rect 13320 18348 13347 18379
rect 13392 18348 13415 18379
rect 13464 18348 13483 18379
rect 13536 18348 13551 18379
rect 13608 18348 13619 18379
rect 13680 18348 13687 18379
rect 13752 18348 13755 18379
rect 13245 18345 13279 18348
rect 13313 18345 13347 18348
rect 13381 18345 13415 18348
rect 13449 18345 13483 18348
rect 13517 18345 13551 18348
rect 13585 18345 13619 18348
rect 13653 18345 13687 18348
rect 13721 18345 13755 18348
rect 13789 18348 13790 18379
rect 13857 18348 13862 18379
rect 13925 18348 13934 18379
rect 13993 18348 14006 18379
rect 14061 18348 14078 18379
rect 14129 18348 14150 18379
rect 14197 18348 14222 18379
rect 14265 18348 14294 18379
rect 14333 18348 14366 18379
rect 13789 18345 13823 18348
rect 13857 18345 13891 18348
rect 13925 18345 13959 18348
rect 13993 18345 14027 18348
rect 14061 18345 14095 18348
rect 14129 18345 14163 18348
rect 14197 18345 14231 18348
rect 14265 18345 14299 18348
rect 14333 18345 14367 18348
rect 14401 18345 14435 18379
rect 14472 18348 14503 18379
rect 14544 18348 14571 18379
rect 14616 18348 14639 18379
rect 14688 18348 14707 18379
rect 14760 18348 14772 18382
rect 14469 18345 14503 18348
rect 14537 18345 14571 18348
rect 14605 18345 14639 18348
rect 14673 18345 14707 18348
rect 14741 18345 14772 18348
rect 197 18309 14772 18345
rect 197 18306 221 18309
rect 255 18306 290 18309
rect 324 18306 359 18309
rect 197 18272 209 18306
rect 255 18275 282 18306
rect 324 18275 355 18306
rect 393 18275 427 18309
rect 461 18306 495 18309
rect 529 18306 563 18309
rect 597 18306 631 18309
rect 665 18306 699 18309
rect 733 18306 767 18309
rect 801 18306 835 18309
rect 869 18306 903 18309
rect 462 18275 495 18306
rect 535 18275 563 18306
rect 608 18275 631 18306
rect 681 18275 699 18306
rect 754 18275 767 18306
rect 827 18275 835 18306
rect 900 18275 903 18306
rect 937 18306 971 18309
rect 1005 18306 1039 18309
rect 1073 18306 1107 18309
rect 1141 18306 1175 18309
rect 1209 18306 1243 18309
rect 1277 18306 1311 18309
rect 1345 18306 1379 18309
rect 937 18275 939 18306
rect 1005 18275 1012 18306
rect 1073 18275 1085 18306
rect 1141 18275 1158 18306
rect 1209 18275 1231 18306
rect 1277 18275 1304 18306
rect 1345 18275 1377 18306
rect 1413 18275 1447 18309
rect 1481 18306 1515 18309
rect 1549 18306 1583 18309
rect 1617 18306 1651 18309
rect 1685 18306 1719 18309
rect 1753 18306 1787 18309
rect 1821 18306 1855 18309
rect 1889 18306 1923 18309
rect 1484 18275 1515 18306
rect 1557 18275 1583 18306
rect 1630 18275 1651 18306
rect 1703 18275 1719 18306
rect 1776 18275 1787 18306
rect 1849 18275 1855 18306
rect 1922 18275 1923 18306
rect 1957 18306 1991 18309
rect 2025 18306 2059 18309
rect 2093 18306 2127 18309
rect 2161 18306 2195 18309
rect 2229 18306 2263 18309
rect 2297 18306 2331 18309
rect 1957 18275 1961 18306
rect 2025 18275 2034 18306
rect 2093 18275 2107 18306
rect 2161 18275 2180 18306
rect 2229 18275 2253 18306
rect 2297 18275 2326 18306
rect 2365 18275 2399 18309
rect 2433 18275 2467 18309
rect 2501 18306 2535 18309
rect 2569 18306 2603 18309
rect 2637 18306 2671 18309
rect 2705 18306 2739 18309
rect 2773 18306 2807 18309
rect 2841 18306 2875 18309
rect 2506 18275 2535 18306
rect 2579 18275 2603 18306
rect 2652 18275 2671 18306
rect 2725 18275 2739 18306
rect 2798 18275 2807 18306
rect 2871 18275 2875 18306
rect 2909 18306 2943 18309
rect 2977 18306 3011 18309
rect 3045 18306 3079 18309
rect 3113 18306 3147 18309
rect 3181 18306 3215 18309
rect 3249 18306 3283 18309
rect 3317 18306 3351 18309
rect 2909 18275 2910 18306
rect 2977 18275 2983 18306
rect 3045 18275 3056 18306
rect 3113 18275 3129 18306
rect 3181 18275 3202 18306
rect 3249 18275 3275 18306
rect 3317 18275 3348 18306
rect 3385 18275 3419 18309
rect 3453 18306 3487 18309
rect 3521 18306 3555 18309
rect 3589 18306 3623 18309
rect 3657 18306 3691 18309
rect 3725 18306 3759 18309
rect 3793 18306 3827 18309
rect 3861 18306 3895 18309
rect 3929 18306 3963 18309
rect 3455 18275 3487 18306
rect 3528 18275 3555 18306
rect 3600 18275 3623 18306
rect 3672 18275 3691 18306
rect 3744 18275 3759 18306
rect 3816 18275 3827 18306
rect 3888 18275 3895 18306
rect 3960 18275 3963 18306
rect 3997 18306 4031 18309
rect 4065 18306 4099 18309
rect 4133 18306 4167 18309
rect 4201 18306 4235 18309
rect 4269 18306 4303 18309
rect 4337 18306 4371 18309
rect 4405 18306 4439 18309
rect 4473 18306 4507 18309
rect 4541 18306 4575 18309
rect 3997 18275 3998 18306
rect 4065 18275 4070 18306
rect 4133 18275 4142 18306
rect 4201 18275 4214 18306
rect 4269 18275 4286 18306
rect 4337 18275 4358 18306
rect 4405 18275 4430 18306
rect 4473 18275 4502 18306
rect 4541 18275 4574 18306
rect 4609 18275 4643 18309
rect 4677 18306 4711 18309
rect 4745 18306 4779 18309
rect 4813 18306 4847 18309
rect 4881 18306 4915 18309
rect 4949 18306 4983 18309
rect 5017 18306 5051 18309
rect 5085 18306 5119 18309
rect 5153 18306 5187 18309
rect 4680 18275 4711 18306
rect 4752 18275 4779 18306
rect 4824 18275 4847 18306
rect 4896 18275 4915 18306
rect 4968 18275 4983 18306
rect 5040 18275 5051 18306
rect 5112 18275 5119 18306
rect 5184 18275 5187 18306
rect 5221 18306 5255 18309
rect 5289 18306 5323 18309
rect 5357 18306 5391 18309
rect 5425 18306 5459 18309
rect 5493 18306 5527 18309
rect 5561 18306 5595 18309
rect 5629 18306 5663 18309
rect 5697 18306 5731 18309
rect 5765 18306 5799 18309
rect 5221 18275 5222 18306
rect 5289 18275 5294 18306
rect 5357 18275 5366 18306
rect 5425 18275 5438 18306
rect 5493 18275 5510 18306
rect 5561 18275 5582 18306
rect 5629 18275 5654 18306
rect 5697 18275 5726 18306
rect 5765 18275 5798 18306
rect 5833 18275 5867 18309
rect 5901 18306 5935 18309
rect 5969 18306 6003 18309
rect 6037 18306 6071 18309
rect 6105 18306 6139 18309
rect 6173 18306 6207 18309
rect 6241 18306 6275 18309
rect 6309 18306 6343 18309
rect 6377 18306 6411 18309
rect 5904 18275 5935 18306
rect 5976 18275 6003 18306
rect 6048 18275 6071 18306
rect 6120 18275 6139 18306
rect 6192 18275 6207 18306
rect 6264 18275 6275 18306
rect 6336 18275 6343 18306
rect 6408 18275 6411 18306
rect 6445 18306 6479 18309
rect 6513 18306 6547 18309
rect 6581 18306 6615 18309
rect 6649 18306 6683 18309
rect 6717 18306 6751 18309
rect 6785 18306 6819 18309
rect 6853 18306 6887 18309
rect 6921 18306 6955 18309
rect 6989 18306 7023 18309
rect 6445 18275 6446 18306
rect 6513 18275 6518 18306
rect 6581 18275 6590 18306
rect 6649 18275 6662 18306
rect 6717 18275 6734 18306
rect 6785 18275 6806 18306
rect 6853 18275 6878 18306
rect 6921 18275 6950 18306
rect 6989 18275 7022 18306
rect 7057 18275 7091 18309
rect 7125 18306 7159 18309
rect 7193 18306 7227 18309
rect 7261 18306 7295 18309
rect 7329 18306 7363 18309
rect 7397 18306 7431 18309
rect 7465 18306 7499 18309
rect 7533 18306 7567 18309
rect 7601 18306 7635 18309
rect 7128 18275 7159 18306
rect 7200 18275 7227 18306
rect 7272 18275 7295 18306
rect 7344 18275 7363 18306
rect 7416 18275 7431 18306
rect 7488 18275 7499 18306
rect 7560 18275 7567 18306
rect 7632 18275 7635 18306
rect 7669 18306 7703 18309
rect 7737 18306 7771 18309
rect 7805 18306 7839 18309
rect 7873 18306 7907 18309
rect 7941 18306 7975 18309
rect 8009 18306 8043 18309
rect 8077 18306 8111 18309
rect 8145 18306 8179 18309
rect 8213 18306 8247 18309
rect 7669 18275 7670 18306
rect 7737 18275 7742 18306
rect 7805 18275 7814 18306
rect 7873 18275 7886 18306
rect 7941 18275 7958 18306
rect 8009 18275 8030 18306
rect 8077 18275 8102 18306
rect 8145 18275 8174 18306
rect 8213 18275 8246 18306
rect 8281 18275 8315 18309
rect 8349 18306 8383 18309
rect 8417 18306 8451 18309
rect 8485 18306 8519 18309
rect 8553 18306 8587 18309
rect 8621 18306 8655 18309
rect 8689 18306 8723 18309
rect 8757 18306 8791 18309
rect 8825 18306 8859 18309
rect 8352 18275 8383 18306
rect 8424 18275 8451 18306
rect 8496 18275 8519 18306
rect 8568 18275 8587 18306
rect 8640 18275 8655 18306
rect 8712 18275 8723 18306
rect 8784 18275 8791 18306
rect 8856 18275 8859 18306
rect 8893 18306 8927 18309
rect 8961 18306 8995 18309
rect 9029 18306 9063 18309
rect 9097 18306 9131 18309
rect 9165 18306 9199 18309
rect 9233 18306 9267 18309
rect 9301 18306 9335 18309
rect 9369 18306 9403 18309
rect 9437 18306 9471 18309
rect 8893 18275 8894 18306
rect 8961 18275 8966 18306
rect 9029 18275 9038 18306
rect 9097 18275 9110 18306
rect 9165 18275 9182 18306
rect 9233 18275 9254 18306
rect 9301 18275 9326 18306
rect 9369 18275 9398 18306
rect 9437 18275 9470 18306
rect 9505 18275 9539 18309
rect 9573 18306 9607 18309
rect 9641 18306 9675 18309
rect 9709 18306 9743 18309
rect 9777 18306 9811 18309
rect 9845 18306 9879 18309
rect 9913 18306 9947 18309
rect 9981 18306 10015 18309
rect 10049 18306 10083 18309
rect 9576 18275 9607 18306
rect 9648 18275 9675 18306
rect 9720 18275 9743 18306
rect 9792 18275 9811 18306
rect 9864 18275 9879 18306
rect 9936 18275 9947 18306
rect 10008 18275 10015 18306
rect 10080 18275 10083 18306
rect 10117 18306 10151 18309
rect 10185 18306 10219 18309
rect 10253 18306 10287 18309
rect 10321 18306 10355 18309
rect 10389 18306 10423 18309
rect 10457 18306 10491 18309
rect 10525 18306 10559 18309
rect 10593 18306 10627 18309
rect 10661 18306 10695 18309
rect 10117 18275 10118 18306
rect 10185 18275 10190 18306
rect 10253 18275 10262 18306
rect 10321 18275 10334 18306
rect 10389 18275 10406 18306
rect 10457 18275 10478 18306
rect 10525 18275 10550 18306
rect 10593 18275 10622 18306
rect 10661 18275 10694 18306
rect 10729 18275 10763 18309
rect 10797 18306 10831 18309
rect 10865 18306 10899 18309
rect 10933 18306 10967 18309
rect 11001 18306 11035 18309
rect 11069 18306 11103 18309
rect 11137 18306 11171 18309
rect 11205 18306 11239 18309
rect 11273 18306 11307 18309
rect 10800 18275 10831 18306
rect 10872 18275 10899 18306
rect 10944 18275 10967 18306
rect 11016 18275 11035 18306
rect 11088 18275 11103 18306
rect 11160 18275 11171 18306
rect 11232 18275 11239 18306
rect 11304 18275 11307 18306
rect 11341 18306 11375 18309
rect 11409 18306 11443 18309
rect 11477 18306 11511 18309
rect 11545 18306 11579 18309
rect 11613 18306 11647 18309
rect 11681 18306 11715 18309
rect 11749 18306 11783 18309
rect 11817 18306 11851 18309
rect 11885 18306 11919 18309
rect 11341 18275 11342 18306
rect 11409 18275 11414 18306
rect 11477 18275 11486 18306
rect 11545 18275 11558 18306
rect 11613 18275 11630 18306
rect 11681 18275 11702 18306
rect 11749 18275 11774 18306
rect 11817 18275 11846 18306
rect 11885 18275 11918 18306
rect 11953 18275 11987 18309
rect 12021 18306 12055 18309
rect 12089 18306 12123 18309
rect 12157 18306 12191 18309
rect 12225 18306 12259 18309
rect 12293 18306 12327 18309
rect 12361 18306 12395 18309
rect 12429 18306 12463 18309
rect 12497 18306 12531 18309
rect 12024 18275 12055 18306
rect 12096 18275 12123 18306
rect 12168 18275 12191 18306
rect 12240 18275 12259 18306
rect 12312 18275 12327 18306
rect 12384 18275 12395 18306
rect 12456 18275 12463 18306
rect 12528 18275 12531 18306
rect 12565 18306 12599 18309
rect 12633 18306 12667 18309
rect 12701 18306 12735 18309
rect 12769 18306 12803 18309
rect 12837 18306 12871 18309
rect 12905 18306 12939 18309
rect 12973 18306 13007 18309
rect 13041 18306 13075 18309
rect 13109 18306 13143 18309
rect 12565 18275 12566 18306
rect 12633 18275 12638 18306
rect 12701 18275 12710 18306
rect 12769 18275 12782 18306
rect 12837 18275 12854 18306
rect 12905 18275 12926 18306
rect 12973 18275 12998 18306
rect 13041 18275 13070 18306
rect 13109 18275 13142 18306
rect 13177 18275 13211 18309
rect 13245 18306 13279 18309
rect 13313 18306 13347 18309
rect 13381 18306 13415 18309
rect 13449 18306 13483 18309
rect 13517 18306 13551 18309
rect 13585 18306 13619 18309
rect 13653 18306 13687 18309
rect 13721 18306 13755 18309
rect 13248 18275 13279 18306
rect 13320 18275 13347 18306
rect 13392 18275 13415 18306
rect 13464 18275 13483 18306
rect 13536 18275 13551 18306
rect 13608 18275 13619 18306
rect 13680 18275 13687 18306
rect 13752 18275 13755 18306
rect 13789 18306 13823 18309
rect 13857 18306 13891 18309
rect 13925 18306 13959 18309
rect 13993 18306 14027 18309
rect 14061 18306 14095 18309
rect 14129 18306 14163 18309
rect 14197 18306 14231 18309
rect 14265 18306 14299 18309
rect 14333 18306 14367 18309
rect 13789 18275 13790 18306
rect 13857 18275 13862 18306
rect 13925 18275 13934 18306
rect 13993 18275 14006 18306
rect 14061 18275 14078 18306
rect 14129 18275 14150 18306
rect 14197 18275 14222 18306
rect 14265 18275 14294 18306
rect 14333 18275 14366 18306
rect 14401 18275 14435 18309
rect 14469 18306 14503 18309
rect 14537 18306 14571 18309
rect 14605 18306 14639 18309
rect 14673 18306 14707 18309
rect 14741 18306 14772 18309
rect 14472 18275 14503 18306
rect 14544 18275 14571 18306
rect 14616 18275 14639 18306
rect 14688 18275 14707 18306
rect 243 18272 282 18275
rect 316 18272 355 18275
rect 389 18272 428 18275
rect 462 18272 501 18275
rect 535 18272 574 18275
rect 608 18272 647 18275
rect 681 18272 720 18275
rect 754 18272 793 18275
rect 827 18272 866 18275
rect 900 18272 939 18275
rect 973 18272 1012 18275
rect 1046 18272 1085 18275
rect 1119 18272 1158 18275
rect 1192 18272 1231 18275
rect 1265 18272 1304 18275
rect 1338 18272 1377 18275
rect 1411 18272 1450 18275
rect 1484 18272 1523 18275
rect 1557 18272 1596 18275
rect 1630 18272 1669 18275
rect 1703 18272 1742 18275
rect 1776 18272 1815 18275
rect 1849 18272 1888 18275
rect 1922 18272 1961 18275
rect 1995 18272 2034 18275
rect 2068 18272 2107 18275
rect 2141 18272 2180 18275
rect 2214 18272 2253 18275
rect 2287 18272 2326 18275
rect 2360 18272 2399 18275
rect 2433 18272 2472 18275
rect 2506 18272 2545 18275
rect 2579 18272 2618 18275
rect 2652 18272 2691 18275
rect 2725 18272 2764 18275
rect 2798 18272 2837 18275
rect 2871 18272 2910 18275
rect 2944 18272 2983 18275
rect 3017 18272 3056 18275
rect 3090 18272 3129 18275
rect 3163 18272 3202 18275
rect 3236 18272 3275 18275
rect 3309 18272 3348 18275
rect 3382 18272 3421 18275
rect 3455 18272 3494 18275
rect 3528 18272 3566 18275
rect 3600 18272 3638 18275
rect 3672 18272 3710 18275
rect 3744 18272 3782 18275
rect 3816 18272 3854 18275
rect 3888 18272 3926 18275
rect 3960 18272 3998 18275
rect 4032 18272 4070 18275
rect 4104 18272 4142 18275
rect 4176 18272 4214 18275
rect 4248 18272 4286 18275
rect 4320 18272 4358 18275
rect 4392 18272 4430 18275
rect 4464 18272 4502 18275
rect 4536 18272 4574 18275
rect 4608 18272 4646 18275
rect 4680 18272 4718 18275
rect 4752 18272 4790 18275
rect 4824 18272 4862 18275
rect 4896 18272 4934 18275
rect 4968 18272 5006 18275
rect 5040 18272 5078 18275
rect 5112 18272 5150 18275
rect 5184 18272 5222 18275
rect 5256 18272 5294 18275
rect 5328 18272 5366 18275
rect 5400 18272 5438 18275
rect 5472 18272 5510 18275
rect 5544 18272 5582 18275
rect 5616 18272 5654 18275
rect 5688 18272 5726 18275
rect 5760 18272 5798 18275
rect 5832 18272 5870 18275
rect 5904 18272 5942 18275
rect 5976 18272 6014 18275
rect 6048 18272 6086 18275
rect 6120 18272 6158 18275
rect 6192 18272 6230 18275
rect 6264 18272 6302 18275
rect 6336 18272 6374 18275
rect 6408 18272 6446 18275
rect 6480 18272 6518 18275
rect 6552 18272 6590 18275
rect 6624 18272 6662 18275
rect 6696 18272 6734 18275
rect 6768 18272 6806 18275
rect 6840 18272 6878 18275
rect 6912 18272 6950 18275
rect 6984 18272 7022 18275
rect 7056 18272 7094 18275
rect 7128 18272 7166 18275
rect 7200 18272 7238 18275
rect 7272 18272 7310 18275
rect 7344 18272 7382 18275
rect 7416 18272 7454 18275
rect 7488 18272 7526 18275
rect 7560 18272 7598 18275
rect 7632 18272 7670 18275
rect 7704 18272 7742 18275
rect 7776 18272 7814 18275
rect 7848 18272 7886 18275
rect 7920 18272 7958 18275
rect 7992 18272 8030 18275
rect 8064 18272 8102 18275
rect 8136 18272 8174 18275
rect 8208 18272 8246 18275
rect 8280 18272 8318 18275
rect 8352 18272 8390 18275
rect 8424 18272 8462 18275
rect 8496 18272 8534 18275
rect 8568 18272 8606 18275
rect 8640 18272 8678 18275
rect 8712 18272 8750 18275
rect 8784 18272 8822 18275
rect 8856 18272 8894 18275
rect 8928 18272 8966 18275
rect 9000 18272 9038 18275
rect 9072 18272 9110 18275
rect 9144 18272 9182 18275
rect 9216 18272 9254 18275
rect 9288 18272 9326 18275
rect 9360 18272 9398 18275
rect 9432 18272 9470 18275
rect 9504 18272 9542 18275
rect 9576 18272 9614 18275
rect 9648 18272 9686 18275
rect 9720 18272 9758 18275
rect 9792 18272 9830 18275
rect 9864 18272 9902 18275
rect 9936 18272 9974 18275
rect 10008 18272 10046 18275
rect 10080 18272 10118 18275
rect 10152 18272 10190 18275
rect 10224 18272 10262 18275
rect 10296 18272 10334 18275
rect 10368 18272 10406 18275
rect 10440 18272 10478 18275
rect 10512 18272 10550 18275
rect 10584 18272 10622 18275
rect 10656 18272 10694 18275
rect 10728 18272 10766 18275
rect 10800 18272 10838 18275
rect 10872 18272 10910 18275
rect 10944 18272 10982 18275
rect 11016 18272 11054 18275
rect 11088 18272 11126 18275
rect 11160 18272 11198 18275
rect 11232 18272 11270 18275
rect 11304 18272 11342 18275
rect 11376 18272 11414 18275
rect 11448 18272 11486 18275
rect 11520 18272 11558 18275
rect 11592 18272 11630 18275
rect 11664 18272 11702 18275
rect 11736 18272 11774 18275
rect 11808 18272 11846 18275
rect 11880 18272 11918 18275
rect 11952 18272 11990 18275
rect 12024 18272 12062 18275
rect 12096 18272 12134 18275
rect 12168 18272 12206 18275
rect 12240 18272 12278 18275
rect 12312 18272 12350 18275
rect 12384 18272 12422 18275
rect 12456 18272 12494 18275
rect 12528 18272 12566 18275
rect 12600 18272 12638 18275
rect 12672 18272 12710 18275
rect 12744 18272 12782 18275
rect 12816 18272 12854 18275
rect 12888 18272 12926 18275
rect 12960 18272 12998 18275
rect 13032 18272 13070 18275
rect 13104 18272 13142 18275
rect 13176 18272 13214 18275
rect 13248 18272 13286 18275
rect 13320 18272 13358 18275
rect 13392 18272 13430 18275
rect 13464 18272 13502 18275
rect 13536 18272 13574 18275
rect 13608 18272 13646 18275
rect 13680 18272 13718 18275
rect 13752 18272 13790 18275
rect 13824 18272 13862 18275
rect 13896 18272 13934 18275
rect 13968 18272 14006 18275
rect 14040 18272 14078 18275
rect 14112 18272 14150 18275
rect 14184 18272 14222 18275
rect 14256 18272 14294 18275
rect 14328 18272 14366 18275
rect 14400 18272 14438 18275
rect 14472 18272 14510 18275
rect 14544 18272 14582 18275
rect 14616 18272 14654 18275
rect 14688 18272 14726 18275
rect 14760 18272 14772 18306
rect 197 18239 14772 18272
rect 197 18230 221 18239
rect 255 18230 290 18239
rect 324 18230 359 18239
rect 197 18196 209 18230
rect 255 18205 282 18230
rect 324 18205 355 18230
rect 393 18205 427 18239
rect 461 18230 495 18239
rect 529 18230 563 18239
rect 597 18230 631 18239
rect 665 18230 699 18239
rect 733 18230 767 18239
rect 801 18230 835 18239
rect 869 18230 903 18239
rect 462 18205 495 18230
rect 535 18205 563 18230
rect 608 18205 631 18230
rect 681 18205 699 18230
rect 754 18205 767 18230
rect 827 18205 835 18230
rect 900 18205 903 18230
rect 937 18230 971 18239
rect 1005 18230 1039 18239
rect 1073 18230 1107 18239
rect 1141 18230 1175 18239
rect 1209 18230 1243 18239
rect 1277 18230 1311 18239
rect 1345 18230 1379 18239
rect 937 18205 939 18230
rect 1005 18205 1012 18230
rect 1073 18205 1085 18230
rect 1141 18205 1158 18230
rect 1209 18205 1231 18230
rect 1277 18205 1304 18230
rect 1345 18205 1377 18230
rect 1413 18205 1447 18239
rect 1481 18230 1515 18239
rect 1549 18230 1583 18239
rect 1617 18230 1651 18239
rect 1685 18230 1719 18239
rect 1753 18230 1787 18239
rect 1821 18230 1855 18239
rect 1889 18230 1923 18239
rect 1484 18205 1515 18230
rect 1557 18205 1583 18230
rect 1630 18205 1651 18230
rect 1703 18205 1719 18230
rect 1776 18205 1787 18230
rect 1849 18205 1855 18230
rect 1922 18205 1923 18230
rect 1957 18230 1991 18239
rect 2025 18230 2059 18239
rect 2093 18230 2127 18239
rect 2161 18230 2195 18239
rect 2229 18230 2263 18239
rect 2297 18230 2331 18239
rect 1957 18205 1961 18230
rect 2025 18205 2034 18230
rect 2093 18205 2107 18230
rect 2161 18205 2180 18230
rect 2229 18205 2253 18230
rect 2297 18205 2326 18230
rect 2365 18205 2399 18239
rect 2433 18205 2467 18239
rect 2501 18230 2535 18239
rect 2569 18230 2603 18239
rect 2637 18230 2671 18239
rect 2705 18230 2739 18239
rect 2773 18230 2807 18239
rect 2841 18230 2875 18239
rect 2506 18205 2535 18230
rect 2579 18205 2603 18230
rect 2652 18205 2671 18230
rect 2725 18205 2739 18230
rect 2798 18205 2807 18230
rect 2871 18205 2875 18230
rect 2909 18230 2943 18239
rect 2977 18230 3011 18239
rect 3045 18230 3079 18239
rect 3113 18230 3147 18239
rect 3181 18230 3215 18239
rect 3249 18230 3283 18239
rect 3317 18230 3351 18239
rect 2909 18205 2910 18230
rect 2977 18205 2983 18230
rect 3045 18205 3056 18230
rect 3113 18205 3129 18230
rect 3181 18205 3202 18230
rect 3249 18205 3275 18230
rect 3317 18205 3348 18230
rect 3385 18205 3419 18239
rect 3453 18230 3487 18239
rect 3521 18230 3555 18239
rect 3589 18230 3623 18239
rect 3657 18230 3691 18239
rect 3725 18230 3759 18239
rect 3793 18230 3827 18239
rect 3861 18230 3895 18239
rect 3929 18230 3963 18239
rect 3455 18205 3487 18230
rect 3528 18205 3555 18230
rect 3600 18205 3623 18230
rect 3672 18205 3691 18230
rect 3744 18205 3759 18230
rect 3816 18205 3827 18230
rect 3888 18205 3895 18230
rect 3960 18205 3963 18230
rect 3997 18230 4031 18239
rect 4065 18230 4099 18239
rect 4133 18230 4167 18239
rect 4201 18230 4235 18239
rect 4269 18230 4303 18239
rect 4337 18230 4371 18239
rect 4405 18230 4439 18239
rect 4473 18230 4507 18239
rect 4541 18230 4575 18239
rect 3997 18205 3998 18230
rect 4065 18205 4070 18230
rect 4133 18205 4142 18230
rect 4201 18205 4214 18230
rect 4269 18205 4286 18230
rect 4337 18205 4358 18230
rect 4405 18205 4430 18230
rect 4473 18205 4502 18230
rect 4541 18205 4574 18230
rect 4609 18205 4643 18239
rect 4677 18230 4711 18239
rect 4745 18230 4779 18239
rect 4813 18230 4847 18239
rect 4881 18230 4915 18239
rect 4949 18230 4983 18239
rect 5017 18230 5051 18239
rect 5085 18230 5119 18239
rect 5153 18230 5187 18239
rect 4680 18205 4711 18230
rect 4752 18205 4779 18230
rect 4824 18205 4847 18230
rect 4896 18205 4915 18230
rect 4968 18205 4983 18230
rect 5040 18205 5051 18230
rect 5112 18205 5119 18230
rect 5184 18205 5187 18230
rect 5221 18230 5255 18239
rect 5289 18230 5323 18239
rect 5357 18230 5391 18239
rect 5425 18230 5459 18239
rect 5493 18230 5527 18239
rect 5561 18230 5595 18239
rect 5629 18230 5663 18239
rect 5697 18230 5731 18239
rect 5765 18230 5799 18239
rect 5221 18205 5222 18230
rect 5289 18205 5294 18230
rect 5357 18205 5366 18230
rect 5425 18205 5438 18230
rect 5493 18205 5510 18230
rect 5561 18205 5582 18230
rect 5629 18205 5654 18230
rect 5697 18205 5726 18230
rect 5765 18205 5798 18230
rect 5833 18205 5867 18239
rect 5901 18230 5935 18239
rect 5969 18230 6003 18239
rect 6037 18230 6071 18239
rect 6105 18230 6139 18239
rect 6173 18230 6207 18239
rect 6241 18230 6275 18239
rect 6309 18230 6343 18239
rect 6377 18230 6411 18239
rect 5904 18205 5935 18230
rect 5976 18205 6003 18230
rect 6048 18205 6071 18230
rect 6120 18205 6139 18230
rect 6192 18205 6207 18230
rect 6264 18205 6275 18230
rect 6336 18205 6343 18230
rect 6408 18205 6411 18230
rect 6445 18230 6479 18239
rect 6513 18230 6547 18239
rect 6581 18230 6615 18239
rect 6649 18230 6683 18239
rect 6717 18230 6751 18239
rect 6785 18230 6819 18239
rect 6853 18230 6887 18239
rect 6921 18230 6955 18239
rect 6989 18230 7023 18239
rect 6445 18205 6446 18230
rect 6513 18205 6518 18230
rect 6581 18205 6590 18230
rect 6649 18205 6662 18230
rect 6717 18205 6734 18230
rect 6785 18205 6806 18230
rect 6853 18205 6878 18230
rect 6921 18205 6950 18230
rect 6989 18205 7022 18230
rect 7057 18205 7091 18239
rect 7125 18230 7159 18239
rect 7193 18230 7227 18239
rect 7261 18230 7295 18239
rect 7329 18230 7363 18239
rect 7397 18230 7431 18239
rect 7465 18230 7499 18239
rect 7533 18230 7567 18239
rect 7601 18230 7635 18239
rect 7128 18205 7159 18230
rect 7200 18205 7227 18230
rect 7272 18205 7295 18230
rect 7344 18205 7363 18230
rect 7416 18205 7431 18230
rect 7488 18205 7499 18230
rect 7560 18205 7567 18230
rect 7632 18205 7635 18230
rect 7669 18230 7703 18239
rect 7737 18230 7771 18239
rect 7805 18230 7839 18239
rect 7873 18230 7907 18239
rect 7941 18230 7975 18239
rect 8009 18230 8043 18239
rect 8077 18230 8111 18239
rect 8145 18230 8179 18239
rect 8213 18230 8247 18239
rect 7669 18205 7670 18230
rect 7737 18205 7742 18230
rect 7805 18205 7814 18230
rect 7873 18205 7886 18230
rect 7941 18205 7958 18230
rect 8009 18205 8030 18230
rect 8077 18205 8102 18230
rect 8145 18205 8174 18230
rect 8213 18205 8246 18230
rect 8281 18205 8315 18239
rect 8349 18230 8383 18239
rect 8417 18230 8451 18239
rect 8485 18230 8519 18239
rect 8553 18230 8587 18239
rect 8621 18230 8655 18239
rect 8689 18230 8723 18239
rect 8757 18230 8791 18239
rect 8825 18230 8859 18239
rect 8352 18205 8383 18230
rect 8424 18205 8451 18230
rect 8496 18205 8519 18230
rect 8568 18205 8587 18230
rect 8640 18205 8655 18230
rect 8712 18205 8723 18230
rect 8784 18205 8791 18230
rect 8856 18205 8859 18230
rect 8893 18230 8927 18239
rect 8961 18230 8995 18239
rect 9029 18230 9063 18239
rect 9097 18230 9131 18239
rect 9165 18230 9199 18239
rect 9233 18230 9267 18239
rect 9301 18230 9335 18239
rect 9369 18230 9403 18239
rect 9437 18230 9471 18239
rect 8893 18205 8894 18230
rect 8961 18205 8966 18230
rect 9029 18205 9038 18230
rect 9097 18205 9110 18230
rect 9165 18205 9182 18230
rect 9233 18205 9254 18230
rect 9301 18205 9326 18230
rect 9369 18205 9398 18230
rect 9437 18205 9470 18230
rect 9505 18205 9539 18239
rect 9573 18230 9607 18239
rect 9641 18230 9675 18239
rect 9709 18230 9743 18239
rect 9777 18230 9811 18239
rect 9845 18230 9879 18239
rect 9913 18230 9947 18239
rect 9981 18230 10015 18239
rect 10049 18230 10083 18239
rect 9576 18205 9607 18230
rect 9648 18205 9675 18230
rect 9720 18205 9743 18230
rect 9792 18205 9811 18230
rect 9864 18205 9879 18230
rect 9936 18205 9947 18230
rect 10008 18205 10015 18230
rect 10080 18205 10083 18230
rect 10117 18230 10151 18239
rect 10185 18230 10219 18239
rect 10253 18230 10287 18239
rect 10321 18230 10355 18239
rect 10389 18230 10423 18239
rect 10457 18230 10491 18239
rect 10525 18230 10559 18239
rect 10593 18230 10627 18239
rect 10661 18230 10695 18239
rect 10117 18205 10118 18230
rect 10185 18205 10190 18230
rect 10253 18205 10262 18230
rect 10321 18205 10334 18230
rect 10389 18205 10406 18230
rect 10457 18205 10478 18230
rect 10525 18205 10550 18230
rect 10593 18205 10622 18230
rect 10661 18205 10694 18230
rect 10729 18205 10763 18239
rect 10797 18230 10831 18239
rect 10865 18230 10899 18239
rect 10933 18230 10967 18239
rect 11001 18230 11035 18239
rect 11069 18230 11103 18239
rect 11137 18230 11171 18239
rect 11205 18230 11239 18239
rect 11273 18230 11307 18239
rect 10800 18205 10831 18230
rect 10872 18205 10899 18230
rect 10944 18205 10967 18230
rect 11016 18205 11035 18230
rect 11088 18205 11103 18230
rect 11160 18205 11171 18230
rect 11232 18205 11239 18230
rect 11304 18205 11307 18230
rect 11341 18230 11375 18239
rect 11409 18230 11443 18239
rect 11477 18230 11511 18239
rect 11545 18230 11579 18239
rect 11613 18230 11647 18239
rect 11681 18230 11715 18239
rect 11749 18230 11783 18239
rect 11817 18230 11851 18239
rect 11885 18230 11919 18239
rect 11341 18205 11342 18230
rect 11409 18205 11414 18230
rect 11477 18205 11486 18230
rect 11545 18205 11558 18230
rect 11613 18205 11630 18230
rect 11681 18205 11702 18230
rect 11749 18205 11774 18230
rect 11817 18205 11846 18230
rect 11885 18205 11918 18230
rect 11953 18205 11987 18239
rect 12021 18230 12055 18239
rect 12089 18230 12123 18239
rect 12157 18230 12191 18239
rect 12225 18230 12259 18239
rect 12293 18230 12327 18239
rect 12361 18230 12395 18239
rect 12429 18230 12463 18239
rect 12497 18230 12531 18239
rect 12024 18205 12055 18230
rect 12096 18205 12123 18230
rect 12168 18205 12191 18230
rect 12240 18205 12259 18230
rect 12312 18205 12327 18230
rect 12384 18205 12395 18230
rect 12456 18205 12463 18230
rect 12528 18205 12531 18230
rect 12565 18230 12599 18239
rect 12633 18230 12667 18239
rect 12701 18230 12735 18239
rect 12769 18230 12803 18239
rect 12837 18230 12871 18239
rect 12905 18230 12939 18239
rect 12973 18230 13007 18239
rect 13041 18230 13075 18239
rect 13109 18230 13143 18239
rect 12565 18205 12566 18230
rect 12633 18205 12638 18230
rect 12701 18205 12710 18230
rect 12769 18205 12782 18230
rect 12837 18205 12854 18230
rect 12905 18205 12926 18230
rect 12973 18205 12998 18230
rect 13041 18205 13070 18230
rect 13109 18205 13142 18230
rect 13177 18205 13211 18239
rect 13245 18230 13279 18239
rect 13313 18230 13347 18239
rect 13381 18230 13415 18239
rect 13449 18230 13483 18239
rect 13517 18230 13551 18239
rect 13585 18230 13619 18239
rect 13653 18230 13687 18239
rect 13721 18230 13755 18239
rect 13248 18205 13279 18230
rect 13320 18205 13347 18230
rect 13392 18205 13415 18230
rect 13464 18205 13483 18230
rect 13536 18205 13551 18230
rect 13608 18205 13619 18230
rect 13680 18205 13687 18230
rect 13752 18205 13755 18230
rect 13789 18230 13823 18239
rect 13857 18230 13891 18239
rect 13925 18230 13959 18239
rect 13993 18230 14027 18239
rect 14061 18230 14095 18239
rect 14129 18230 14163 18239
rect 14197 18230 14231 18239
rect 14265 18230 14299 18239
rect 14333 18230 14367 18239
rect 13789 18205 13790 18230
rect 13857 18205 13862 18230
rect 13925 18205 13934 18230
rect 13993 18205 14006 18230
rect 14061 18205 14078 18230
rect 14129 18205 14150 18230
rect 14197 18205 14222 18230
rect 14265 18205 14294 18230
rect 14333 18205 14366 18230
rect 14401 18205 14435 18239
rect 14469 18230 14503 18239
rect 14537 18230 14571 18239
rect 14605 18230 14639 18239
rect 14673 18230 14707 18239
rect 14741 18230 14772 18239
rect 14472 18205 14503 18230
rect 14544 18205 14571 18230
rect 14616 18205 14639 18230
rect 14688 18205 14707 18230
rect 243 18196 282 18205
rect 316 18196 355 18205
rect 389 18196 428 18205
rect 462 18196 501 18205
rect 535 18196 574 18205
rect 608 18196 647 18205
rect 681 18196 720 18205
rect 754 18196 793 18205
rect 827 18196 866 18205
rect 900 18196 939 18205
rect 973 18196 1012 18205
rect 1046 18196 1085 18205
rect 1119 18196 1158 18205
rect 1192 18196 1231 18205
rect 1265 18196 1304 18205
rect 1338 18196 1377 18205
rect 1411 18196 1450 18205
rect 1484 18196 1523 18205
rect 1557 18196 1596 18205
rect 1630 18196 1669 18205
rect 1703 18196 1742 18205
rect 1776 18196 1815 18205
rect 1849 18196 1888 18205
rect 1922 18196 1961 18205
rect 1995 18196 2034 18205
rect 2068 18196 2107 18205
rect 2141 18196 2180 18205
rect 2214 18196 2253 18205
rect 2287 18196 2326 18205
rect 2360 18196 2399 18205
rect 2433 18196 2472 18205
rect 2506 18196 2545 18205
rect 2579 18196 2618 18205
rect 2652 18196 2691 18205
rect 2725 18196 2764 18205
rect 2798 18196 2837 18205
rect 2871 18196 2910 18205
rect 2944 18196 2983 18205
rect 3017 18196 3056 18205
rect 3090 18196 3129 18205
rect 3163 18196 3202 18205
rect 3236 18196 3275 18205
rect 3309 18196 3348 18205
rect 3382 18196 3421 18205
rect 3455 18196 3494 18205
rect 3528 18196 3566 18205
rect 3600 18196 3638 18205
rect 3672 18196 3710 18205
rect 3744 18196 3782 18205
rect 3816 18196 3854 18205
rect 3888 18196 3926 18205
rect 3960 18196 3998 18205
rect 4032 18196 4070 18205
rect 4104 18196 4142 18205
rect 4176 18196 4214 18205
rect 4248 18196 4286 18205
rect 4320 18196 4358 18205
rect 4392 18196 4430 18205
rect 4464 18196 4502 18205
rect 4536 18196 4574 18205
rect 4608 18196 4646 18205
rect 4680 18196 4718 18205
rect 4752 18196 4790 18205
rect 4824 18196 4862 18205
rect 4896 18196 4934 18205
rect 4968 18196 5006 18205
rect 5040 18196 5078 18205
rect 5112 18196 5150 18205
rect 5184 18196 5222 18205
rect 5256 18196 5294 18205
rect 5328 18196 5366 18205
rect 5400 18196 5438 18205
rect 5472 18196 5510 18205
rect 5544 18196 5582 18205
rect 5616 18196 5654 18205
rect 5688 18196 5726 18205
rect 5760 18196 5798 18205
rect 5832 18196 5870 18205
rect 5904 18196 5942 18205
rect 5976 18196 6014 18205
rect 6048 18196 6086 18205
rect 6120 18196 6158 18205
rect 6192 18196 6230 18205
rect 6264 18196 6302 18205
rect 6336 18196 6374 18205
rect 6408 18196 6446 18205
rect 6480 18196 6518 18205
rect 6552 18196 6590 18205
rect 6624 18196 6662 18205
rect 6696 18196 6734 18205
rect 6768 18196 6806 18205
rect 6840 18196 6878 18205
rect 6912 18196 6950 18205
rect 6984 18196 7022 18205
rect 7056 18196 7094 18205
rect 7128 18196 7166 18205
rect 7200 18196 7238 18205
rect 7272 18196 7310 18205
rect 7344 18196 7382 18205
rect 7416 18196 7454 18205
rect 7488 18196 7526 18205
rect 7560 18196 7598 18205
rect 7632 18196 7670 18205
rect 7704 18196 7742 18205
rect 7776 18196 7814 18205
rect 7848 18196 7886 18205
rect 7920 18196 7958 18205
rect 7992 18196 8030 18205
rect 8064 18196 8102 18205
rect 8136 18196 8174 18205
rect 8208 18196 8246 18205
rect 8280 18196 8318 18205
rect 8352 18196 8390 18205
rect 8424 18196 8462 18205
rect 8496 18196 8534 18205
rect 8568 18196 8606 18205
rect 8640 18196 8678 18205
rect 8712 18196 8750 18205
rect 8784 18196 8822 18205
rect 8856 18196 8894 18205
rect 8928 18196 8966 18205
rect 9000 18196 9038 18205
rect 9072 18196 9110 18205
rect 9144 18196 9182 18205
rect 9216 18196 9254 18205
rect 9288 18196 9326 18205
rect 9360 18196 9398 18205
rect 9432 18196 9470 18205
rect 9504 18196 9542 18205
rect 9576 18196 9614 18205
rect 9648 18196 9686 18205
rect 9720 18196 9758 18205
rect 9792 18196 9830 18205
rect 9864 18196 9902 18205
rect 9936 18196 9974 18205
rect 10008 18196 10046 18205
rect 10080 18196 10118 18205
rect 10152 18196 10190 18205
rect 10224 18196 10262 18205
rect 10296 18196 10334 18205
rect 10368 18196 10406 18205
rect 10440 18196 10478 18205
rect 10512 18196 10550 18205
rect 10584 18196 10622 18205
rect 10656 18196 10694 18205
rect 10728 18196 10766 18205
rect 10800 18196 10838 18205
rect 10872 18196 10910 18205
rect 10944 18196 10982 18205
rect 11016 18196 11054 18205
rect 11088 18196 11126 18205
rect 11160 18196 11198 18205
rect 11232 18196 11270 18205
rect 11304 18196 11342 18205
rect 11376 18196 11414 18205
rect 11448 18196 11486 18205
rect 11520 18196 11558 18205
rect 11592 18196 11630 18205
rect 11664 18196 11702 18205
rect 11736 18196 11774 18205
rect 11808 18196 11846 18205
rect 11880 18196 11918 18205
rect 11952 18196 11990 18205
rect 12024 18196 12062 18205
rect 12096 18196 12134 18205
rect 12168 18196 12206 18205
rect 12240 18196 12278 18205
rect 12312 18196 12350 18205
rect 12384 18196 12422 18205
rect 12456 18196 12494 18205
rect 12528 18196 12566 18205
rect 12600 18196 12638 18205
rect 12672 18196 12710 18205
rect 12744 18196 12782 18205
rect 12816 18196 12854 18205
rect 12888 18196 12926 18205
rect 12960 18196 12998 18205
rect 13032 18196 13070 18205
rect 13104 18196 13142 18205
rect 13176 18196 13214 18205
rect 13248 18196 13286 18205
rect 13320 18196 13358 18205
rect 13392 18196 13430 18205
rect 13464 18196 13502 18205
rect 13536 18196 13574 18205
rect 13608 18196 13646 18205
rect 13680 18196 13718 18205
rect 13752 18196 13790 18205
rect 13824 18196 13862 18205
rect 13896 18196 13934 18205
rect 13968 18196 14006 18205
rect 14040 18196 14078 18205
rect 14112 18196 14150 18205
rect 14184 18196 14222 18205
rect 14256 18196 14294 18205
rect 14328 18196 14366 18205
rect 14400 18196 14438 18205
rect 14472 18196 14510 18205
rect 14544 18196 14582 18205
rect 14616 18196 14654 18205
rect 14688 18196 14726 18205
rect 14760 18196 14772 18230
rect 197 18169 14772 18196
rect 197 18154 221 18169
rect 255 18154 290 18169
rect 324 18154 359 18169
rect 197 18120 209 18154
rect 255 18135 282 18154
rect 324 18135 355 18154
rect 393 18135 427 18169
rect 461 18154 495 18169
rect 529 18154 563 18169
rect 597 18154 631 18169
rect 665 18154 699 18169
rect 733 18154 767 18169
rect 801 18154 835 18169
rect 869 18154 903 18169
rect 462 18135 495 18154
rect 535 18135 563 18154
rect 608 18135 631 18154
rect 681 18135 699 18154
rect 754 18135 767 18154
rect 827 18135 835 18154
rect 900 18135 903 18154
rect 937 18154 971 18169
rect 1005 18154 1039 18169
rect 1073 18154 1107 18169
rect 1141 18154 1175 18169
rect 1209 18154 1243 18169
rect 1277 18154 1311 18169
rect 1345 18154 1379 18169
rect 937 18135 939 18154
rect 1005 18135 1012 18154
rect 1073 18135 1085 18154
rect 1141 18135 1158 18154
rect 1209 18135 1231 18154
rect 1277 18135 1304 18154
rect 1345 18135 1377 18154
rect 1413 18135 1447 18169
rect 1481 18154 1515 18169
rect 1549 18154 1583 18169
rect 1617 18154 1651 18169
rect 1685 18154 1719 18169
rect 1753 18154 1787 18169
rect 1821 18154 1855 18169
rect 1889 18154 1923 18169
rect 1484 18135 1515 18154
rect 1557 18135 1583 18154
rect 1630 18135 1651 18154
rect 1703 18135 1719 18154
rect 1776 18135 1787 18154
rect 1849 18135 1855 18154
rect 1922 18135 1923 18154
rect 1957 18154 1991 18169
rect 2025 18154 2059 18169
rect 2093 18154 2127 18169
rect 2161 18154 2195 18169
rect 2229 18154 2263 18169
rect 2297 18154 2331 18169
rect 1957 18135 1961 18154
rect 2025 18135 2034 18154
rect 2093 18135 2107 18154
rect 2161 18135 2180 18154
rect 2229 18135 2253 18154
rect 2297 18135 2326 18154
rect 2365 18135 2399 18169
rect 2433 18135 2467 18169
rect 2501 18154 2535 18169
rect 2569 18154 2603 18169
rect 2637 18154 2671 18169
rect 2705 18154 2739 18169
rect 2773 18154 2807 18169
rect 2841 18154 2875 18169
rect 2506 18135 2535 18154
rect 2579 18135 2603 18154
rect 2652 18135 2671 18154
rect 2725 18135 2739 18154
rect 2798 18135 2807 18154
rect 2871 18135 2875 18154
rect 2909 18154 2943 18169
rect 2977 18154 3011 18169
rect 3045 18154 3079 18169
rect 3113 18154 3147 18169
rect 3181 18154 3215 18169
rect 3249 18154 3283 18169
rect 3317 18154 3351 18169
rect 2909 18135 2910 18154
rect 2977 18135 2983 18154
rect 3045 18135 3056 18154
rect 3113 18135 3129 18154
rect 3181 18135 3202 18154
rect 3249 18135 3275 18154
rect 3317 18135 3348 18154
rect 3385 18135 3419 18169
rect 3453 18154 3487 18169
rect 3521 18154 3555 18169
rect 3589 18154 3623 18169
rect 3657 18154 3691 18169
rect 3725 18154 3759 18169
rect 3793 18154 3827 18169
rect 3861 18154 3895 18169
rect 3929 18154 3963 18169
rect 3455 18135 3487 18154
rect 3528 18135 3555 18154
rect 3600 18135 3623 18154
rect 3672 18135 3691 18154
rect 3744 18135 3759 18154
rect 3816 18135 3827 18154
rect 3888 18135 3895 18154
rect 3960 18135 3963 18154
rect 3997 18154 4031 18169
rect 4065 18154 4099 18169
rect 4133 18154 4167 18169
rect 4201 18154 4235 18169
rect 4269 18154 4303 18169
rect 4337 18154 4371 18169
rect 4405 18154 4439 18169
rect 4473 18154 4507 18169
rect 4541 18154 4575 18169
rect 3997 18135 3998 18154
rect 4065 18135 4070 18154
rect 4133 18135 4142 18154
rect 4201 18135 4214 18154
rect 4269 18135 4286 18154
rect 4337 18135 4358 18154
rect 4405 18135 4430 18154
rect 4473 18135 4502 18154
rect 4541 18135 4574 18154
rect 4609 18135 4643 18169
rect 4677 18154 4711 18169
rect 4745 18154 4779 18169
rect 4813 18154 4847 18169
rect 4881 18154 4915 18169
rect 4949 18154 4983 18169
rect 5017 18154 5051 18169
rect 5085 18154 5119 18169
rect 5153 18154 5187 18169
rect 4680 18135 4711 18154
rect 4752 18135 4779 18154
rect 4824 18135 4847 18154
rect 4896 18135 4915 18154
rect 4968 18135 4983 18154
rect 5040 18135 5051 18154
rect 5112 18135 5119 18154
rect 5184 18135 5187 18154
rect 5221 18154 5255 18169
rect 5289 18154 5323 18169
rect 5357 18154 5391 18169
rect 5425 18154 5459 18169
rect 5493 18154 5527 18169
rect 5561 18154 5595 18169
rect 5629 18154 5663 18169
rect 5697 18154 5731 18169
rect 5765 18154 5799 18169
rect 5221 18135 5222 18154
rect 5289 18135 5294 18154
rect 5357 18135 5366 18154
rect 5425 18135 5438 18154
rect 5493 18135 5510 18154
rect 5561 18135 5582 18154
rect 5629 18135 5654 18154
rect 5697 18135 5726 18154
rect 5765 18135 5798 18154
rect 5833 18135 5867 18169
rect 5901 18154 5935 18169
rect 5969 18154 6003 18169
rect 6037 18154 6071 18169
rect 6105 18154 6139 18169
rect 6173 18154 6207 18169
rect 6241 18154 6275 18169
rect 6309 18154 6343 18169
rect 6377 18154 6411 18169
rect 5904 18135 5935 18154
rect 5976 18135 6003 18154
rect 6048 18135 6071 18154
rect 6120 18135 6139 18154
rect 6192 18135 6207 18154
rect 6264 18135 6275 18154
rect 6336 18135 6343 18154
rect 6408 18135 6411 18154
rect 6445 18154 6479 18169
rect 6513 18154 6547 18169
rect 6581 18154 6615 18169
rect 6649 18154 6683 18169
rect 6717 18154 6751 18169
rect 6785 18154 6819 18169
rect 6853 18154 6887 18169
rect 6921 18154 6955 18169
rect 6989 18154 7023 18169
rect 6445 18135 6446 18154
rect 6513 18135 6518 18154
rect 6581 18135 6590 18154
rect 6649 18135 6662 18154
rect 6717 18135 6734 18154
rect 6785 18135 6806 18154
rect 6853 18135 6878 18154
rect 6921 18135 6950 18154
rect 6989 18135 7022 18154
rect 7057 18135 7091 18169
rect 7125 18154 7159 18169
rect 7193 18154 7227 18169
rect 7261 18154 7295 18169
rect 7329 18154 7363 18169
rect 7397 18154 7431 18169
rect 7465 18154 7499 18169
rect 7533 18154 7567 18169
rect 7601 18154 7635 18169
rect 7128 18135 7159 18154
rect 7200 18135 7227 18154
rect 7272 18135 7295 18154
rect 7344 18135 7363 18154
rect 7416 18135 7431 18154
rect 7488 18135 7499 18154
rect 7560 18135 7567 18154
rect 7632 18135 7635 18154
rect 7669 18154 7703 18169
rect 7737 18154 7771 18169
rect 7805 18154 7839 18169
rect 7873 18154 7907 18169
rect 7941 18154 7975 18169
rect 8009 18154 8043 18169
rect 8077 18154 8111 18169
rect 8145 18154 8179 18169
rect 8213 18154 8247 18169
rect 7669 18135 7670 18154
rect 7737 18135 7742 18154
rect 7805 18135 7814 18154
rect 7873 18135 7886 18154
rect 7941 18135 7958 18154
rect 8009 18135 8030 18154
rect 8077 18135 8102 18154
rect 8145 18135 8174 18154
rect 8213 18135 8246 18154
rect 8281 18135 8315 18169
rect 8349 18154 8383 18169
rect 8417 18154 8451 18169
rect 8485 18154 8519 18169
rect 8553 18154 8587 18169
rect 8621 18154 8655 18169
rect 8689 18154 8723 18169
rect 8757 18154 8791 18169
rect 8825 18154 8859 18169
rect 8352 18135 8383 18154
rect 8424 18135 8451 18154
rect 8496 18135 8519 18154
rect 8568 18135 8587 18154
rect 8640 18135 8655 18154
rect 8712 18135 8723 18154
rect 8784 18135 8791 18154
rect 8856 18135 8859 18154
rect 8893 18154 8927 18169
rect 8961 18154 8995 18169
rect 9029 18154 9063 18169
rect 9097 18154 9131 18169
rect 9165 18154 9199 18169
rect 9233 18154 9267 18169
rect 9301 18154 9335 18169
rect 9369 18154 9403 18169
rect 9437 18154 9471 18169
rect 8893 18135 8894 18154
rect 8961 18135 8966 18154
rect 9029 18135 9038 18154
rect 9097 18135 9110 18154
rect 9165 18135 9182 18154
rect 9233 18135 9254 18154
rect 9301 18135 9326 18154
rect 9369 18135 9398 18154
rect 9437 18135 9470 18154
rect 9505 18135 9539 18169
rect 9573 18154 9607 18169
rect 9641 18154 9675 18169
rect 9709 18154 9743 18169
rect 9777 18154 9811 18169
rect 9845 18154 9879 18169
rect 9913 18154 9947 18169
rect 9981 18154 10015 18169
rect 10049 18154 10083 18169
rect 9576 18135 9607 18154
rect 9648 18135 9675 18154
rect 9720 18135 9743 18154
rect 9792 18135 9811 18154
rect 9864 18135 9879 18154
rect 9936 18135 9947 18154
rect 10008 18135 10015 18154
rect 10080 18135 10083 18154
rect 10117 18154 10151 18169
rect 10185 18154 10219 18169
rect 10253 18154 10287 18169
rect 10321 18154 10355 18169
rect 10389 18154 10423 18169
rect 10457 18154 10491 18169
rect 10525 18154 10559 18169
rect 10593 18154 10627 18169
rect 10661 18154 10695 18169
rect 10117 18135 10118 18154
rect 10185 18135 10190 18154
rect 10253 18135 10262 18154
rect 10321 18135 10334 18154
rect 10389 18135 10406 18154
rect 10457 18135 10478 18154
rect 10525 18135 10550 18154
rect 10593 18135 10622 18154
rect 10661 18135 10694 18154
rect 10729 18135 10763 18169
rect 10797 18154 10831 18169
rect 10865 18154 10899 18169
rect 10933 18154 10967 18169
rect 11001 18154 11035 18169
rect 11069 18154 11103 18169
rect 11137 18154 11171 18169
rect 11205 18154 11239 18169
rect 11273 18154 11307 18169
rect 10800 18135 10831 18154
rect 10872 18135 10899 18154
rect 10944 18135 10967 18154
rect 11016 18135 11035 18154
rect 11088 18135 11103 18154
rect 11160 18135 11171 18154
rect 11232 18135 11239 18154
rect 11304 18135 11307 18154
rect 11341 18154 11375 18169
rect 11409 18154 11443 18169
rect 11477 18154 11511 18169
rect 11545 18154 11579 18169
rect 11613 18154 11647 18169
rect 11681 18154 11715 18169
rect 11749 18154 11783 18169
rect 11817 18154 11851 18169
rect 11885 18154 11919 18169
rect 11341 18135 11342 18154
rect 11409 18135 11414 18154
rect 11477 18135 11486 18154
rect 11545 18135 11558 18154
rect 11613 18135 11630 18154
rect 11681 18135 11702 18154
rect 11749 18135 11774 18154
rect 11817 18135 11846 18154
rect 11885 18135 11918 18154
rect 11953 18135 11987 18169
rect 12021 18154 12055 18169
rect 12089 18154 12123 18169
rect 12157 18154 12191 18169
rect 12225 18154 12259 18169
rect 12293 18154 12327 18169
rect 12361 18154 12395 18169
rect 12429 18154 12463 18169
rect 12497 18154 12531 18169
rect 12024 18135 12055 18154
rect 12096 18135 12123 18154
rect 12168 18135 12191 18154
rect 12240 18135 12259 18154
rect 12312 18135 12327 18154
rect 12384 18135 12395 18154
rect 12456 18135 12463 18154
rect 12528 18135 12531 18154
rect 12565 18154 12599 18169
rect 12633 18154 12667 18169
rect 12701 18154 12735 18169
rect 12769 18154 12803 18169
rect 12837 18154 12871 18169
rect 12905 18154 12939 18169
rect 12973 18154 13007 18169
rect 13041 18154 13075 18169
rect 13109 18154 13143 18169
rect 12565 18135 12566 18154
rect 12633 18135 12638 18154
rect 12701 18135 12710 18154
rect 12769 18135 12782 18154
rect 12837 18135 12854 18154
rect 12905 18135 12926 18154
rect 12973 18135 12998 18154
rect 13041 18135 13070 18154
rect 13109 18135 13142 18154
rect 13177 18135 13211 18169
rect 13245 18154 13279 18169
rect 13313 18154 13347 18169
rect 13381 18154 13415 18169
rect 13449 18154 13483 18169
rect 13517 18154 13551 18169
rect 13585 18154 13619 18169
rect 13653 18154 13687 18169
rect 13721 18154 13755 18169
rect 13248 18135 13279 18154
rect 13320 18135 13347 18154
rect 13392 18135 13415 18154
rect 13464 18135 13483 18154
rect 13536 18135 13551 18154
rect 13608 18135 13619 18154
rect 13680 18135 13687 18154
rect 13752 18135 13755 18154
rect 13789 18154 13823 18169
rect 13857 18154 13891 18169
rect 13925 18154 13959 18169
rect 13993 18154 14027 18169
rect 14061 18154 14095 18169
rect 14129 18154 14163 18169
rect 14197 18154 14231 18169
rect 14265 18154 14299 18169
rect 14333 18154 14367 18169
rect 13789 18135 13790 18154
rect 13857 18135 13862 18154
rect 13925 18135 13934 18154
rect 13993 18135 14006 18154
rect 14061 18135 14078 18154
rect 14129 18135 14150 18154
rect 14197 18135 14222 18154
rect 14265 18135 14294 18154
rect 14333 18135 14366 18154
rect 14401 18135 14435 18169
rect 14469 18154 14503 18169
rect 14537 18154 14571 18169
rect 14605 18154 14639 18169
rect 14673 18154 14707 18169
rect 14741 18154 14772 18169
rect 14472 18135 14503 18154
rect 14544 18135 14571 18154
rect 14616 18135 14639 18154
rect 14688 18135 14707 18154
rect 243 18120 282 18135
rect 316 18120 355 18135
rect 389 18120 428 18135
rect 462 18120 501 18135
rect 535 18120 574 18135
rect 608 18120 647 18135
rect 681 18120 720 18135
rect 754 18120 793 18135
rect 827 18120 866 18135
rect 900 18120 939 18135
rect 973 18120 1012 18135
rect 1046 18120 1085 18135
rect 1119 18120 1158 18135
rect 1192 18120 1231 18135
rect 1265 18120 1304 18135
rect 1338 18120 1377 18135
rect 1411 18120 1450 18135
rect 1484 18120 1523 18135
rect 1557 18120 1596 18135
rect 1630 18120 1669 18135
rect 1703 18120 1742 18135
rect 1776 18120 1815 18135
rect 1849 18120 1888 18135
rect 1922 18120 1961 18135
rect 1995 18120 2034 18135
rect 2068 18120 2107 18135
rect 2141 18120 2180 18135
rect 2214 18120 2253 18135
rect 2287 18120 2326 18135
rect 2360 18120 2399 18135
rect 2433 18120 2472 18135
rect 2506 18120 2545 18135
rect 2579 18120 2618 18135
rect 2652 18120 2691 18135
rect 2725 18120 2764 18135
rect 2798 18120 2837 18135
rect 2871 18120 2910 18135
rect 2944 18120 2983 18135
rect 3017 18120 3056 18135
rect 3090 18120 3129 18135
rect 3163 18120 3202 18135
rect 3236 18120 3275 18135
rect 3309 18120 3348 18135
rect 3382 18120 3421 18135
rect 3455 18120 3494 18135
rect 3528 18120 3566 18135
rect 3600 18120 3638 18135
rect 3672 18120 3710 18135
rect 3744 18120 3782 18135
rect 3816 18120 3854 18135
rect 3888 18120 3926 18135
rect 3960 18120 3998 18135
rect 4032 18120 4070 18135
rect 4104 18120 4142 18135
rect 4176 18120 4214 18135
rect 4248 18120 4286 18135
rect 4320 18120 4358 18135
rect 4392 18120 4430 18135
rect 4464 18120 4502 18135
rect 4536 18120 4574 18135
rect 4608 18120 4646 18135
rect 4680 18120 4718 18135
rect 4752 18120 4790 18135
rect 4824 18120 4862 18135
rect 4896 18120 4934 18135
rect 4968 18120 5006 18135
rect 5040 18120 5078 18135
rect 5112 18120 5150 18135
rect 5184 18120 5222 18135
rect 5256 18120 5294 18135
rect 5328 18120 5366 18135
rect 5400 18120 5438 18135
rect 5472 18120 5510 18135
rect 5544 18120 5582 18135
rect 5616 18120 5654 18135
rect 5688 18120 5726 18135
rect 5760 18120 5798 18135
rect 5832 18120 5870 18135
rect 5904 18120 5942 18135
rect 5976 18120 6014 18135
rect 6048 18120 6086 18135
rect 6120 18120 6158 18135
rect 6192 18120 6230 18135
rect 6264 18120 6302 18135
rect 6336 18120 6374 18135
rect 6408 18120 6446 18135
rect 6480 18120 6518 18135
rect 6552 18120 6590 18135
rect 6624 18120 6662 18135
rect 6696 18120 6734 18135
rect 6768 18120 6806 18135
rect 6840 18120 6878 18135
rect 6912 18120 6950 18135
rect 6984 18120 7022 18135
rect 7056 18120 7094 18135
rect 7128 18120 7166 18135
rect 7200 18120 7238 18135
rect 7272 18120 7310 18135
rect 7344 18120 7382 18135
rect 7416 18120 7454 18135
rect 7488 18120 7526 18135
rect 7560 18120 7598 18135
rect 7632 18120 7670 18135
rect 7704 18120 7742 18135
rect 7776 18120 7814 18135
rect 7848 18120 7886 18135
rect 7920 18120 7958 18135
rect 7992 18120 8030 18135
rect 8064 18120 8102 18135
rect 8136 18120 8174 18135
rect 8208 18120 8246 18135
rect 8280 18120 8318 18135
rect 8352 18120 8390 18135
rect 8424 18120 8462 18135
rect 8496 18120 8534 18135
rect 8568 18120 8606 18135
rect 8640 18120 8678 18135
rect 8712 18120 8750 18135
rect 8784 18120 8822 18135
rect 8856 18120 8894 18135
rect 8928 18120 8966 18135
rect 9000 18120 9038 18135
rect 9072 18120 9110 18135
rect 9144 18120 9182 18135
rect 9216 18120 9254 18135
rect 9288 18120 9326 18135
rect 9360 18120 9398 18135
rect 9432 18120 9470 18135
rect 9504 18120 9542 18135
rect 9576 18120 9614 18135
rect 9648 18120 9686 18135
rect 9720 18120 9758 18135
rect 9792 18120 9830 18135
rect 9864 18120 9902 18135
rect 9936 18120 9974 18135
rect 10008 18120 10046 18135
rect 10080 18120 10118 18135
rect 10152 18120 10190 18135
rect 10224 18120 10262 18135
rect 10296 18120 10334 18135
rect 10368 18120 10406 18135
rect 10440 18120 10478 18135
rect 10512 18120 10550 18135
rect 10584 18120 10622 18135
rect 10656 18120 10694 18135
rect 10728 18120 10766 18135
rect 10800 18120 10838 18135
rect 10872 18120 10910 18135
rect 10944 18120 10982 18135
rect 11016 18120 11054 18135
rect 11088 18120 11126 18135
rect 11160 18120 11198 18135
rect 11232 18120 11270 18135
rect 11304 18120 11342 18135
rect 11376 18120 11414 18135
rect 11448 18120 11486 18135
rect 11520 18120 11558 18135
rect 11592 18120 11630 18135
rect 11664 18120 11702 18135
rect 11736 18120 11774 18135
rect 11808 18120 11846 18135
rect 11880 18120 11918 18135
rect 11952 18120 11990 18135
rect 12024 18120 12062 18135
rect 12096 18120 12134 18135
rect 12168 18120 12206 18135
rect 12240 18120 12278 18135
rect 12312 18120 12350 18135
rect 12384 18120 12422 18135
rect 12456 18120 12494 18135
rect 12528 18120 12566 18135
rect 12600 18120 12638 18135
rect 12672 18120 12710 18135
rect 12744 18120 12782 18135
rect 12816 18120 12854 18135
rect 12888 18120 12926 18135
rect 12960 18120 12998 18135
rect 13032 18120 13070 18135
rect 13104 18120 13142 18135
rect 13176 18120 13214 18135
rect 13248 18120 13286 18135
rect 13320 18120 13358 18135
rect 13392 18120 13430 18135
rect 13464 18120 13502 18135
rect 13536 18120 13574 18135
rect 13608 18120 13646 18135
rect 13680 18120 13718 18135
rect 13752 18120 13790 18135
rect 13824 18120 13862 18135
rect 13896 18120 13934 18135
rect 13968 18120 14006 18135
rect 14040 18120 14078 18135
rect 14112 18120 14150 18135
rect 14184 18120 14222 18135
rect 14256 18120 14294 18135
rect 14328 18120 14366 18135
rect 14400 18120 14438 18135
rect 14472 18120 14510 18135
rect 14544 18120 14582 18135
rect 14616 18120 14654 18135
rect 14688 18120 14726 18135
rect 14760 18120 14772 18154
rect 197 18099 14772 18120
rect 197 18078 221 18099
rect 255 18078 290 18099
rect 324 18078 359 18099
rect 197 18044 209 18078
rect 255 18065 282 18078
rect 324 18065 355 18078
rect 393 18065 427 18099
rect 461 18078 495 18099
rect 529 18078 563 18099
rect 597 18078 631 18099
rect 665 18078 699 18099
rect 733 18078 767 18099
rect 801 18078 835 18099
rect 869 18078 903 18099
rect 462 18065 495 18078
rect 535 18065 563 18078
rect 608 18065 631 18078
rect 681 18065 699 18078
rect 754 18065 767 18078
rect 827 18065 835 18078
rect 900 18065 903 18078
rect 937 18078 971 18099
rect 1005 18078 1039 18099
rect 1073 18078 1107 18099
rect 1141 18078 1175 18099
rect 1209 18078 1243 18099
rect 1277 18078 1311 18099
rect 1345 18078 1379 18099
rect 937 18065 939 18078
rect 1005 18065 1012 18078
rect 1073 18065 1085 18078
rect 1141 18065 1158 18078
rect 1209 18065 1231 18078
rect 1277 18065 1304 18078
rect 1345 18065 1377 18078
rect 1413 18065 1447 18099
rect 1481 18078 1515 18099
rect 1549 18078 1583 18099
rect 1617 18078 1651 18099
rect 1685 18078 1719 18099
rect 1753 18078 1787 18099
rect 1821 18078 1855 18099
rect 1889 18078 1923 18099
rect 1484 18065 1515 18078
rect 1557 18065 1583 18078
rect 1630 18065 1651 18078
rect 1703 18065 1719 18078
rect 1776 18065 1787 18078
rect 1849 18065 1855 18078
rect 1922 18065 1923 18078
rect 1957 18078 1991 18099
rect 2025 18078 2059 18099
rect 2093 18078 2127 18099
rect 2161 18078 2195 18099
rect 2229 18078 2263 18099
rect 2297 18078 2331 18099
rect 1957 18065 1961 18078
rect 2025 18065 2034 18078
rect 2093 18065 2107 18078
rect 2161 18065 2180 18078
rect 2229 18065 2253 18078
rect 2297 18065 2326 18078
rect 2365 18065 2399 18099
rect 2433 18065 2467 18099
rect 2501 18078 2535 18099
rect 2569 18078 2603 18099
rect 2637 18078 2671 18099
rect 2705 18078 2739 18099
rect 2773 18078 2807 18099
rect 2841 18078 2875 18099
rect 2506 18065 2535 18078
rect 2579 18065 2603 18078
rect 2652 18065 2671 18078
rect 2725 18065 2739 18078
rect 2798 18065 2807 18078
rect 2871 18065 2875 18078
rect 2909 18078 2943 18099
rect 2977 18078 3011 18099
rect 3045 18078 3079 18099
rect 3113 18078 3147 18099
rect 3181 18078 3215 18099
rect 3249 18078 3283 18099
rect 3317 18078 3351 18099
rect 2909 18065 2910 18078
rect 2977 18065 2983 18078
rect 3045 18065 3056 18078
rect 3113 18065 3129 18078
rect 3181 18065 3202 18078
rect 3249 18065 3275 18078
rect 3317 18065 3348 18078
rect 3385 18065 3419 18099
rect 3453 18078 3487 18099
rect 3521 18078 3555 18099
rect 3589 18078 3623 18099
rect 3657 18078 3691 18099
rect 3725 18078 3759 18099
rect 3793 18078 3827 18099
rect 3861 18078 3895 18099
rect 3929 18078 3963 18099
rect 3455 18065 3487 18078
rect 3528 18065 3555 18078
rect 3600 18065 3623 18078
rect 3672 18065 3691 18078
rect 3744 18065 3759 18078
rect 3816 18065 3827 18078
rect 3888 18065 3895 18078
rect 3960 18065 3963 18078
rect 3997 18078 4031 18099
rect 4065 18078 4099 18099
rect 4133 18078 4167 18099
rect 4201 18078 4235 18099
rect 4269 18078 4303 18099
rect 4337 18078 4371 18099
rect 4405 18078 4439 18099
rect 4473 18078 4507 18099
rect 4541 18078 4575 18099
rect 3997 18065 3998 18078
rect 4065 18065 4070 18078
rect 4133 18065 4142 18078
rect 4201 18065 4214 18078
rect 4269 18065 4286 18078
rect 4337 18065 4358 18078
rect 4405 18065 4430 18078
rect 4473 18065 4502 18078
rect 4541 18065 4574 18078
rect 4609 18065 4643 18099
rect 4677 18078 4711 18099
rect 4745 18078 4779 18099
rect 4813 18078 4847 18099
rect 4881 18078 4915 18099
rect 4949 18078 4983 18099
rect 5017 18078 5051 18099
rect 5085 18078 5119 18099
rect 5153 18078 5187 18099
rect 4680 18065 4711 18078
rect 4752 18065 4779 18078
rect 4824 18065 4847 18078
rect 4896 18065 4915 18078
rect 4968 18065 4983 18078
rect 5040 18065 5051 18078
rect 5112 18065 5119 18078
rect 5184 18065 5187 18078
rect 5221 18078 5255 18099
rect 5289 18078 5323 18099
rect 5357 18078 5391 18099
rect 5425 18078 5459 18099
rect 5493 18078 5527 18099
rect 5561 18078 5595 18099
rect 5629 18078 5663 18099
rect 5697 18078 5731 18099
rect 5765 18078 5799 18099
rect 5221 18065 5222 18078
rect 5289 18065 5294 18078
rect 5357 18065 5366 18078
rect 5425 18065 5438 18078
rect 5493 18065 5510 18078
rect 5561 18065 5582 18078
rect 5629 18065 5654 18078
rect 5697 18065 5726 18078
rect 5765 18065 5798 18078
rect 5833 18065 5867 18099
rect 5901 18078 5935 18099
rect 5969 18078 6003 18099
rect 6037 18078 6071 18099
rect 6105 18078 6139 18099
rect 6173 18078 6207 18099
rect 6241 18078 6275 18099
rect 6309 18078 6343 18099
rect 6377 18078 6411 18099
rect 5904 18065 5935 18078
rect 5976 18065 6003 18078
rect 6048 18065 6071 18078
rect 6120 18065 6139 18078
rect 6192 18065 6207 18078
rect 6264 18065 6275 18078
rect 6336 18065 6343 18078
rect 6408 18065 6411 18078
rect 6445 18078 6479 18099
rect 6513 18078 6547 18099
rect 6581 18078 6615 18099
rect 6649 18078 6683 18099
rect 6717 18078 6751 18099
rect 6785 18078 6819 18099
rect 6853 18078 6887 18099
rect 6921 18078 6955 18099
rect 6989 18078 7023 18099
rect 6445 18065 6446 18078
rect 6513 18065 6518 18078
rect 6581 18065 6590 18078
rect 6649 18065 6662 18078
rect 6717 18065 6734 18078
rect 6785 18065 6806 18078
rect 6853 18065 6878 18078
rect 6921 18065 6950 18078
rect 6989 18065 7022 18078
rect 7057 18065 7091 18099
rect 7125 18078 7159 18099
rect 7193 18078 7227 18099
rect 7261 18078 7295 18099
rect 7329 18078 7363 18099
rect 7397 18078 7431 18099
rect 7465 18078 7499 18099
rect 7533 18078 7567 18099
rect 7601 18078 7635 18099
rect 7128 18065 7159 18078
rect 7200 18065 7227 18078
rect 7272 18065 7295 18078
rect 7344 18065 7363 18078
rect 7416 18065 7431 18078
rect 7488 18065 7499 18078
rect 7560 18065 7567 18078
rect 7632 18065 7635 18078
rect 7669 18078 7703 18099
rect 7737 18078 7771 18099
rect 7805 18078 7839 18099
rect 7873 18078 7907 18099
rect 7941 18078 7975 18099
rect 8009 18078 8043 18099
rect 8077 18078 8111 18099
rect 8145 18078 8179 18099
rect 8213 18078 8247 18099
rect 7669 18065 7670 18078
rect 7737 18065 7742 18078
rect 7805 18065 7814 18078
rect 7873 18065 7886 18078
rect 7941 18065 7958 18078
rect 8009 18065 8030 18078
rect 8077 18065 8102 18078
rect 8145 18065 8174 18078
rect 8213 18065 8246 18078
rect 8281 18065 8315 18099
rect 8349 18078 8383 18099
rect 8417 18078 8451 18099
rect 8485 18078 8519 18099
rect 8553 18078 8587 18099
rect 8621 18078 8655 18099
rect 8689 18078 8723 18099
rect 8757 18078 8791 18099
rect 8825 18078 8859 18099
rect 8352 18065 8383 18078
rect 8424 18065 8451 18078
rect 8496 18065 8519 18078
rect 8568 18065 8587 18078
rect 8640 18065 8655 18078
rect 8712 18065 8723 18078
rect 8784 18065 8791 18078
rect 8856 18065 8859 18078
rect 8893 18078 8927 18099
rect 8961 18078 8995 18099
rect 9029 18078 9063 18099
rect 9097 18078 9131 18099
rect 9165 18078 9199 18099
rect 9233 18078 9267 18099
rect 9301 18078 9335 18099
rect 9369 18078 9403 18099
rect 9437 18078 9471 18099
rect 8893 18065 8894 18078
rect 8961 18065 8966 18078
rect 9029 18065 9038 18078
rect 9097 18065 9110 18078
rect 9165 18065 9182 18078
rect 9233 18065 9254 18078
rect 9301 18065 9326 18078
rect 9369 18065 9398 18078
rect 9437 18065 9470 18078
rect 9505 18065 9539 18099
rect 9573 18078 9607 18099
rect 9641 18078 9675 18099
rect 9709 18078 9743 18099
rect 9777 18078 9811 18099
rect 9845 18078 9879 18099
rect 9913 18078 9947 18099
rect 9981 18078 10015 18099
rect 10049 18078 10083 18099
rect 9576 18065 9607 18078
rect 9648 18065 9675 18078
rect 9720 18065 9743 18078
rect 9792 18065 9811 18078
rect 9864 18065 9879 18078
rect 9936 18065 9947 18078
rect 10008 18065 10015 18078
rect 10080 18065 10083 18078
rect 10117 18078 10151 18099
rect 10185 18078 10219 18099
rect 10253 18078 10287 18099
rect 10321 18078 10355 18099
rect 10389 18078 10423 18099
rect 10457 18078 10491 18099
rect 10525 18078 10559 18099
rect 10593 18078 10627 18099
rect 10661 18078 10695 18099
rect 10117 18065 10118 18078
rect 10185 18065 10190 18078
rect 10253 18065 10262 18078
rect 10321 18065 10334 18078
rect 10389 18065 10406 18078
rect 10457 18065 10478 18078
rect 10525 18065 10550 18078
rect 10593 18065 10622 18078
rect 10661 18065 10694 18078
rect 10729 18065 10763 18099
rect 10797 18078 10831 18099
rect 10865 18078 10899 18099
rect 10933 18078 10967 18099
rect 11001 18078 11035 18099
rect 11069 18078 11103 18099
rect 11137 18078 11171 18099
rect 11205 18078 11239 18099
rect 11273 18078 11307 18099
rect 10800 18065 10831 18078
rect 10872 18065 10899 18078
rect 10944 18065 10967 18078
rect 11016 18065 11035 18078
rect 11088 18065 11103 18078
rect 11160 18065 11171 18078
rect 11232 18065 11239 18078
rect 11304 18065 11307 18078
rect 11341 18078 11375 18099
rect 11409 18078 11443 18099
rect 11477 18078 11511 18099
rect 11545 18078 11579 18099
rect 11613 18078 11647 18099
rect 11681 18078 11715 18099
rect 11749 18078 11783 18099
rect 11817 18078 11851 18099
rect 11885 18078 11919 18099
rect 11341 18065 11342 18078
rect 11409 18065 11414 18078
rect 11477 18065 11486 18078
rect 11545 18065 11558 18078
rect 11613 18065 11630 18078
rect 11681 18065 11702 18078
rect 11749 18065 11774 18078
rect 11817 18065 11846 18078
rect 11885 18065 11918 18078
rect 11953 18065 11987 18099
rect 12021 18078 12055 18099
rect 12089 18078 12123 18099
rect 12157 18078 12191 18099
rect 12225 18078 12259 18099
rect 12293 18078 12327 18099
rect 12361 18078 12395 18099
rect 12429 18078 12463 18099
rect 12497 18078 12531 18099
rect 12024 18065 12055 18078
rect 12096 18065 12123 18078
rect 12168 18065 12191 18078
rect 12240 18065 12259 18078
rect 12312 18065 12327 18078
rect 12384 18065 12395 18078
rect 12456 18065 12463 18078
rect 12528 18065 12531 18078
rect 12565 18078 12599 18099
rect 12633 18078 12667 18099
rect 12701 18078 12735 18099
rect 12769 18078 12803 18099
rect 12837 18078 12871 18099
rect 12905 18078 12939 18099
rect 12973 18078 13007 18099
rect 13041 18078 13075 18099
rect 13109 18078 13143 18099
rect 12565 18065 12566 18078
rect 12633 18065 12638 18078
rect 12701 18065 12710 18078
rect 12769 18065 12782 18078
rect 12837 18065 12854 18078
rect 12905 18065 12926 18078
rect 12973 18065 12998 18078
rect 13041 18065 13070 18078
rect 13109 18065 13142 18078
rect 13177 18065 13211 18099
rect 13245 18078 13279 18099
rect 13313 18078 13347 18099
rect 13381 18078 13415 18099
rect 13449 18078 13483 18099
rect 13517 18078 13551 18099
rect 13585 18078 13619 18099
rect 13653 18078 13687 18099
rect 13721 18078 13755 18099
rect 13248 18065 13279 18078
rect 13320 18065 13347 18078
rect 13392 18065 13415 18078
rect 13464 18065 13483 18078
rect 13536 18065 13551 18078
rect 13608 18065 13619 18078
rect 13680 18065 13687 18078
rect 13752 18065 13755 18078
rect 13789 18078 13823 18099
rect 13857 18078 13891 18099
rect 13925 18078 13959 18099
rect 13993 18078 14027 18099
rect 14061 18078 14095 18099
rect 14129 18078 14163 18099
rect 14197 18078 14231 18099
rect 14265 18078 14299 18099
rect 14333 18078 14367 18099
rect 13789 18065 13790 18078
rect 13857 18065 13862 18078
rect 13925 18065 13934 18078
rect 13993 18065 14006 18078
rect 14061 18065 14078 18078
rect 14129 18065 14150 18078
rect 14197 18065 14222 18078
rect 14265 18065 14294 18078
rect 14333 18065 14366 18078
rect 14401 18065 14435 18099
rect 14469 18078 14503 18099
rect 14537 18078 14571 18099
rect 14605 18078 14639 18099
rect 14673 18078 14707 18099
rect 14741 18078 14772 18099
rect 14472 18065 14503 18078
rect 14544 18065 14571 18078
rect 14616 18065 14639 18078
rect 14688 18065 14707 18078
rect 243 18044 282 18065
rect 316 18044 355 18065
rect 389 18044 428 18065
rect 462 18044 501 18065
rect 535 18044 574 18065
rect 608 18044 647 18065
rect 681 18044 720 18065
rect 754 18044 793 18065
rect 827 18044 866 18065
rect 900 18044 939 18065
rect 973 18044 1012 18065
rect 1046 18044 1085 18065
rect 1119 18044 1158 18065
rect 1192 18044 1231 18065
rect 1265 18044 1304 18065
rect 1338 18044 1377 18065
rect 1411 18044 1450 18065
rect 1484 18044 1523 18065
rect 1557 18044 1596 18065
rect 1630 18044 1669 18065
rect 1703 18044 1742 18065
rect 1776 18044 1815 18065
rect 1849 18044 1888 18065
rect 1922 18044 1961 18065
rect 1995 18044 2034 18065
rect 2068 18044 2107 18065
rect 2141 18044 2180 18065
rect 2214 18044 2253 18065
rect 2287 18044 2326 18065
rect 2360 18044 2399 18065
rect 2433 18044 2472 18065
rect 2506 18044 2545 18065
rect 2579 18044 2618 18065
rect 2652 18044 2691 18065
rect 2725 18044 2764 18065
rect 2798 18044 2837 18065
rect 2871 18044 2910 18065
rect 2944 18044 2983 18065
rect 3017 18044 3056 18065
rect 3090 18044 3129 18065
rect 3163 18044 3202 18065
rect 3236 18044 3275 18065
rect 3309 18044 3348 18065
rect 3382 18044 3421 18065
rect 3455 18044 3494 18065
rect 3528 18044 3566 18065
rect 3600 18044 3638 18065
rect 3672 18044 3710 18065
rect 3744 18044 3782 18065
rect 3816 18044 3854 18065
rect 3888 18044 3926 18065
rect 3960 18044 3998 18065
rect 4032 18044 4070 18065
rect 4104 18044 4142 18065
rect 4176 18044 4214 18065
rect 4248 18044 4286 18065
rect 4320 18044 4358 18065
rect 4392 18044 4430 18065
rect 4464 18044 4502 18065
rect 4536 18044 4574 18065
rect 4608 18044 4646 18065
rect 4680 18044 4718 18065
rect 4752 18044 4790 18065
rect 4824 18044 4862 18065
rect 4896 18044 4934 18065
rect 4968 18044 5006 18065
rect 5040 18044 5078 18065
rect 5112 18044 5150 18065
rect 5184 18044 5222 18065
rect 5256 18044 5294 18065
rect 5328 18044 5366 18065
rect 5400 18044 5438 18065
rect 5472 18044 5510 18065
rect 5544 18044 5582 18065
rect 5616 18044 5654 18065
rect 5688 18044 5726 18065
rect 5760 18044 5798 18065
rect 5832 18044 5870 18065
rect 5904 18044 5942 18065
rect 5976 18044 6014 18065
rect 6048 18044 6086 18065
rect 6120 18044 6158 18065
rect 6192 18044 6230 18065
rect 6264 18044 6302 18065
rect 6336 18044 6374 18065
rect 6408 18044 6446 18065
rect 6480 18044 6518 18065
rect 6552 18044 6590 18065
rect 6624 18044 6662 18065
rect 6696 18044 6734 18065
rect 6768 18044 6806 18065
rect 6840 18044 6878 18065
rect 6912 18044 6950 18065
rect 6984 18044 7022 18065
rect 7056 18044 7094 18065
rect 7128 18044 7166 18065
rect 7200 18044 7238 18065
rect 7272 18044 7310 18065
rect 7344 18044 7382 18065
rect 7416 18044 7454 18065
rect 7488 18044 7526 18065
rect 7560 18044 7598 18065
rect 7632 18044 7670 18065
rect 7704 18044 7742 18065
rect 7776 18044 7814 18065
rect 7848 18044 7886 18065
rect 7920 18044 7958 18065
rect 7992 18044 8030 18065
rect 8064 18044 8102 18065
rect 8136 18044 8174 18065
rect 8208 18044 8246 18065
rect 8280 18044 8318 18065
rect 8352 18044 8390 18065
rect 8424 18044 8462 18065
rect 8496 18044 8534 18065
rect 8568 18044 8606 18065
rect 8640 18044 8678 18065
rect 8712 18044 8750 18065
rect 8784 18044 8822 18065
rect 8856 18044 8894 18065
rect 8928 18044 8966 18065
rect 9000 18044 9038 18065
rect 9072 18044 9110 18065
rect 9144 18044 9182 18065
rect 9216 18044 9254 18065
rect 9288 18044 9326 18065
rect 9360 18044 9398 18065
rect 9432 18044 9470 18065
rect 9504 18044 9542 18065
rect 9576 18044 9614 18065
rect 9648 18044 9686 18065
rect 9720 18044 9758 18065
rect 9792 18044 9830 18065
rect 9864 18044 9902 18065
rect 9936 18044 9974 18065
rect 10008 18044 10046 18065
rect 10080 18044 10118 18065
rect 10152 18044 10190 18065
rect 10224 18044 10262 18065
rect 10296 18044 10334 18065
rect 10368 18044 10406 18065
rect 10440 18044 10478 18065
rect 10512 18044 10550 18065
rect 10584 18044 10622 18065
rect 10656 18044 10694 18065
rect 10728 18044 10766 18065
rect 10800 18044 10838 18065
rect 10872 18044 10910 18065
rect 10944 18044 10982 18065
rect 11016 18044 11054 18065
rect 11088 18044 11126 18065
rect 11160 18044 11198 18065
rect 11232 18044 11270 18065
rect 11304 18044 11342 18065
rect 11376 18044 11414 18065
rect 11448 18044 11486 18065
rect 11520 18044 11558 18065
rect 11592 18044 11630 18065
rect 11664 18044 11702 18065
rect 11736 18044 11774 18065
rect 11808 18044 11846 18065
rect 11880 18044 11918 18065
rect 11952 18044 11990 18065
rect 12024 18044 12062 18065
rect 12096 18044 12134 18065
rect 12168 18044 12206 18065
rect 12240 18044 12278 18065
rect 12312 18044 12350 18065
rect 12384 18044 12422 18065
rect 12456 18044 12494 18065
rect 12528 18044 12566 18065
rect 12600 18044 12638 18065
rect 12672 18044 12710 18065
rect 12744 18044 12782 18065
rect 12816 18044 12854 18065
rect 12888 18044 12926 18065
rect 12960 18044 12998 18065
rect 13032 18044 13070 18065
rect 13104 18044 13142 18065
rect 13176 18044 13214 18065
rect 13248 18044 13286 18065
rect 13320 18044 13358 18065
rect 13392 18044 13430 18065
rect 13464 18044 13502 18065
rect 13536 18044 13574 18065
rect 13608 18044 13646 18065
rect 13680 18044 13718 18065
rect 13752 18044 13790 18065
rect 13824 18044 13862 18065
rect 13896 18044 13934 18065
rect 13968 18044 14006 18065
rect 14040 18044 14078 18065
rect 14112 18044 14150 18065
rect 14184 18044 14222 18065
rect 14256 18044 14294 18065
rect 14328 18044 14366 18065
rect 14400 18044 14438 18065
rect 14472 18044 14510 18065
rect 14544 18044 14582 18065
rect 14616 18044 14654 18065
rect 14688 18044 14726 18065
rect 14760 18044 14772 18078
rect 197 18029 14772 18044
rect 197 18002 221 18029
rect 255 18002 290 18029
rect 324 18002 359 18029
rect 197 17968 209 18002
rect 255 17995 282 18002
rect 324 17995 355 18002
rect 393 17995 427 18029
rect 461 18002 495 18029
rect 529 18002 563 18029
rect 597 18002 631 18029
rect 665 18002 699 18029
rect 733 18002 767 18029
rect 801 18002 835 18029
rect 869 18002 903 18029
rect 462 17995 495 18002
rect 535 17995 563 18002
rect 608 17995 631 18002
rect 681 17995 699 18002
rect 754 17995 767 18002
rect 827 17995 835 18002
rect 900 17995 903 18002
rect 937 18002 971 18029
rect 1005 18002 1039 18029
rect 1073 18002 1107 18029
rect 1141 18002 1175 18029
rect 1209 18002 1243 18029
rect 1277 18002 1311 18029
rect 1345 18002 1379 18029
rect 937 17995 939 18002
rect 1005 17995 1012 18002
rect 1073 17995 1085 18002
rect 1141 17995 1158 18002
rect 1209 17995 1231 18002
rect 1277 17995 1304 18002
rect 1345 17995 1377 18002
rect 1413 17995 1447 18029
rect 1481 18002 1515 18029
rect 1549 18002 1583 18029
rect 1617 18002 1651 18029
rect 1685 18002 1719 18029
rect 1753 18002 1787 18029
rect 1821 18002 1855 18029
rect 1889 18002 1923 18029
rect 1484 17995 1515 18002
rect 1557 17995 1583 18002
rect 1630 17995 1651 18002
rect 1703 17995 1719 18002
rect 1776 17995 1787 18002
rect 1849 17995 1855 18002
rect 1922 17995 1923 18002
rect 1957 18002 1991 18029
rect 2025 18002 2059 18029
rect 2093 18002 2127 18029
rect 2161 18002 2195 18029
rect 2229 18002 2263 18029
rect 2297 18002 2331 18029
rect 1957 17995 1961 18002
rect 2025 17995 2034 18002
rect 2093 17995 2107 18002
rect 2161 17995 2180 18002
rect 2229 17995 2253 18002
rect 2297 17995 2326 18002
rect 2365 17995 2399 18029
rect 2433 17995 2467 18029
rect 2501 18002 2535 18029
rect 2569 18002 2603 18029
rect 2637 18002 2671 18029
rect 2705 18002 2739 18029
rect 2773 18002 2807 18029
rect 2841 18002 2875 18029
rect 2506 17995 2535 18002
rect 2579 17995 2603 18002
rect 2652 17995 2671 18002
rect 2725 17995 2739 18002
rect 2798 17995 2807 18002
rect 2871 17995 2875 18002
rect 2909 18002 2943 18029
rect 2977 18002 3011 18029
rect 3045 18002 3079 18029
rect 3113 18002 3147 18029
rect 3181 18002 3215 18029
rect 3249 18002 3283 18029
rect 3317 18002 3351 18029
rect 2909 17995 2910 18002
rect 2977 17995 2983 18002
rect 3045 17995 3056 18002
rect 3113 17995 3129 18002
rect 3181 17995 3202 18002
rect 3249 17995 3275 18002
rect 3317 17995 3348 18002
rect 3385 17995 3419 18029
rect 3453 18002 3487 18029
rect 3521 18002 3555 18029
rect 3589 18002 3623 18029
rect 3657 18002 3691 18029
rect 3725 18002 3759 18029
rect 3793 18002 3827 18029
rect 3861 18002 3895 18029
rect 3929 18002 3963 18029
rect 3455 17995 3487 18002
rect 3528 17995 3555 18002
rect 3600 17995 3623 18002
rect 3672 17995 3691 18002
rect 3744 17995 3759 18002
rect 3816 17995 3827 18002
rect 3888 17995 3895 18002
rect 3960 17995 3963 18002
rect 3997 18002 4031 18029
rect 4065 18002 4099 18029
rect 4133 18002 4167 18029
rect 4201 18002 4235 18029
rect 4269 18002 4303 18029
rect 4337 18002 4371 18029
rect 4405 18002 4439 18029
rect 4473 18002 4507 18029
rect 4541 18002 4575 18029
rect 3997 17995 3998 18002
rect 4065 17995 4070 18002
rect 4133 17995 4142 18002
rect 4201 17995 4214 18002
rect 4269 17995 4286 18002
rect 4337 17995 4358 18002
rect 4405 17995 4430 18002
rect 4473 17995 4502 18002
rect 4541 17995 4574 18002
rect 4609 17995 4643 18029
rect 4677 18002 4711 18029
rect 4745 18002 4779 18029
rect 4813 18002 4847 18029
rect 4881 18002 4915 18029
rect 4949 18002 4983 18029
rect 5017 18002 5051 18029
rect 5085 18002 5119 18029
rect 5153 18002 5187 18029
rect 4680 17995 4711 18002
rect 4752 17995 4779 18002
rect 4824 17995 4847 18002
rect 4896 17995 4915 18002
rect 4968 17995 4983 18002
rect 5040 17995 5051 18002
rect 5112 17995 5119 18002
rect 5184 17995 5187 18002
rect 5221 18002 5255 18029
rect 5289 18002 5323 18029
rect 5357 18002 5391 18029
rect 5425 18002 5459 18029
rect 5493 18002 5527 18029
rect 5561 18002 5595 18029
rect 5629 18002 5663 18029
rect 5697 18002 5731 18029
rect 5765 18002 5799 18029
rect 5221 17995 5222 18002
rect 5289 17995 5294 18002
rect 5357 17995 5366 18002
rect 5425 17995 5438 18002
rect 5493 17995 5510 18002
rect 5561 17995 5582 18002
rect 5629 17995 5654 18002
rect 5697 17995 5726 18002
rect 5765 17995 5798 18002
rect 5833 17995 5867 18029
rect 5901 18002 5935 18029
rect 5969 18002 6003 18029
rect 6037 18002 6071 18029
rect 6105 18002 6139 18029
rect 6173 18002 6207 18029
rect 6241 18002 6275 18029
rect 6309 18002 6343 18029
rect 6377 18002 6411 18029
rect 5904 17995 5935 18002
rect 5976 17995 6003 18002
rect 6048 17995 6071 18002
rect 6120 17995 6139 18002
rect 6192 17995 6207 18002
rect 6264 17995 6275 18002
rect 6336 17995 6343 18002
rect 6408 17995 6411 18002
rect 6445 18002 6479 18029
rect 6513 18002 6547 18029
rect 6581 18002 6615 18029
rect 6649 18002 6683 18029
rect 6717 18002 6751 18029
rect 6785 18002 6819 18029
rect 6853 18002 6887 18029
rect 6921 18002 6955 18029
rect 6989 18002 7023 18029
rect 6445 17995 6446 18002
rect 6513 17995 6518 18002
rect 6581 17995 6590 18002
rect 6649 17995 6662 18002
rect 6717 17995 6734 18002
rect 6785 17995 6806 18002
rect 6853 17995 6878 18002
rect 6921 17995 6950 18002
rect 6989 17995 7022 18002
rect 7057 17995 7091 18029
rect 7125 18002 7159 18029
rect 7193 18002 7227 18029
rect 7261 18002 7295 18029
rect 7329 18002 7363 18029
rect 7397 18002 7431 18029
rect 7465 18002 7499 18029
rect 7533 18002 7567 18029
rect 7601 18002 7635 18029
rect 7128 17995 7159 18002
rect 7200 17995 7227 18002
rect 7272 17995 7295 18002
rect 7344 17995 7363 18002
rect 7416 17995 7431 18002
rect 7488 17995 7499 18002
rect 7560 17995 7567 18002
rect 7632 17995 7635 18002
rect 7669 18002 7703 18029
rect 7737 18002 7771 18029
rect 7805 18002 7839 18029
rect 7873 18002 7907 18029
rect 7941 18002 7975 18029
rect 8009 18002 8043 18029
rect 8077 18002 8111 18029
rect 8145 18002 8179 18029
rect 8213 18002 8247 18029
rect 7669 17995 7670 18002
rect 7737 17995 7742 18002
rect 7805 17995 7814 18002
rect 7873 17995 7886 18002
rect 7941 17995 7958 18002
rect 8009 17995 8030 18002
rect 8077 17995 8102 18002
rect 8145 17995 8174 18002
rect 8213 17995 8246 18002
rect 8281 17995 8315 18029
rect 8349 18002 8383 18029
rect 8417 18002 8451 18029
rect 8485 18002 8519 18029
rect 8553 18002 8587 18029
rect 8621 18002 8655 18029
rect 8689 18002 8723 18029
rect 8757 18002 8791 18029
rect 8825 18002 8859 18029
rect 8352 17995 8383 18002
rect 8424 17995 8451 18002
rect 8496 17995 8519 18002
rect 8568 17995 8587 18002
rect 8640 17995 8655 18002
rect 8712 17995 8723 18002
rect 8784 17995 8791 18002
rect 8856 17995 8859 18002
rect 8893 18002 8927 18029
rect 8961 18002 8995 18029
rect 9029 18002 9063 18029
rect 9097 18002 9131 18029
rect 9165 18002 9199 18029
rect 9233 18002 9267 18029
rect 9301 18002 9335 18029
rect 9369 18002 9403 18029
rect 9437 18002 9471 18029
rect 8893 17995 8894 18002
rect 8961 17995 8966 18002
rect 9029 17995 9038 18002
rect 9097 17995 9110 18002
rect 9165 17995 9182 18002
rect 9233 17995 9254 18002
rect 9301 17995 9326 18002
rect 9369 17995 9398 18002
rect 9437 17995 9470 18002
rect 9505 17995 9539 18029
rect 9573 18002 9607 18029
rect 9641 18002 9675 18029
rect 9709 18002 9743 18029
rect 9777 18002 9811 18029
rect 9845 18002 9879 18029
rect 9913 18002 9947 18029
rect 9981 18002 10015 18029
rect 10049 18002 10083 18029
rect 9576 17995 9607 18002
rect 9648 17995 9675 18002
rect 9720 17995 9743 18002
rect 9792 17995 9811 18002
rect 9864 17995 9879 18002
rect 9936 17995 9947 18002
rect 10008 17995 10015 18002
rect 10080 17995 10083 18002
rect 10117 18002 10151 18029
rect 10185 18002 10219 18029
rect 10253 18002 10287 18029
rect 10321 18002 10355 18029
rect 10389 18002 10423 18029
rect 10457 18002 10491 18029
rect 10525 18002 10559 18029
rect 10593 18002 10627 18029
rect 10661 18002 10695 18029
rect 10117 17995 10118 18002
rect 10185 17995 10190 18002
rect 10253 17995 10262 18002
rect 10321 17995 10334 18002
rect 10389 17995 10406 18002
rect 10457 17995 10478 18002
rect 10525 17995 10550 18002
rect 10593 17995 10622 18002
rect 10661 17995 10694 18002
rect 10729 17995 10763 18029
rect 10797 18002 10831 18029
rect 10865 18002 10899 18029
rect 10933 18002 10967 18029
rect 11001 18002 11035 18029
rect 11069 18002 11103 18029
rect 11137 18002 11171 18029
rect 11205 18002 11239 18029
rect 11273 18002 11307 18029
rect 10800 17995 10831 18002
rect 10872 17995 10899 18002
rect 10944 17995 10967 18002
rect 11016 17995 11035 18002
rect 11088 17995 11103 18002
rect 11160 17995 11171 18002
rect 11232 17995 11239 18002
rect 11304 17995 11307 18002
rect 11341 18002 11375 18029
rect 11409 18002 11443 18029
rect 11477 18002 11511 18029
rect 11545 18002 11579 18029
rect 11613 18002 11647 18029
rect 11681 18002 11715 18029
rect 11749 18002 11783 18029
rect 11817 18002 11851 18029
rect 11885 18002 11919 18029
rect 11341 17995 11342 18002
rect 11409 17995 11414 18002
rect 11477 17995 11486 18002
rect 11545 17995 11558 18002
rect 11613 17995 11630 18002
rect 11681 17995 11702 18002
rect 11749 17995 11774 18002
rect 11817 17995 11846 18002
rect 11885 17995 11918 18002
rect 11953 17995 11987 18029
rect 12021 18002 12055 18029
rect 12089 18002 12123 18029
rect 12157 18002 12191 18029
rect 12225 18002 12259 18029
rect 12293 18002 12327 18029
rect 12361 18002 12395 18029
rect 12429 18002 12463 18029
rect 12497 18002 12531 18029
rect 12024 17995 12055 18002
rect 12096 17995 12123 18002
rect 12168 17995 12191 18002
rect 12240 17995 12259 18002
rect 12312 17995 12327 18002
rect 12384 17995 12395 18002
rect 12456 17995 12463 18002
rect 12528 17995 12531 18002
rect 12565 18002 12599 18029
rect 12633 18002 12667 18029
rect 12701 18002 12735 18029
rect 12769 18002 12803 18029
rect 12837 18002 12871 18029
rect 12905 18002 12939 18029
rect 12973 18002 13007 18029
rect 13041 18002 13075 18029
rect 13109 18002 13143 18029
rect 12565 17995 12566 18002
rect 12633 17995 12638 18002
rect 12701 17995 12710 18002
rect 12769 17995 12782 18002
rect 12837 17995 12854 18002
rect 12905 17995 12926 18002
rect 12973 17995 12998 18002
rect 13041 17995 13070 18002
rect 13109 17995 13142 18002
rect 13177 17995 13211 18029
rect 13245 18002 13279 18029
rect 13313 18002 13347 18029
rect 13381 18002 13415 18029
rect 13449 18002 13483 18029
rect 13517 18002 13551 18029
rect 13585 18002 13619 18029
rect 13653 18002 13687 18029
rect 13721 18002 13755 18029
rect 13248 17995 13279 18002
rect 13320 17995 13347 18002
rect 13392 17995 13415 18002
rect 13464 17995 13483 18002
rect 13536 17995 13551 18002
rect 13608 17995 13619 18002
rect 13680 17995 13687 18002
rect 13752 17995 13755 18002
rect 13789 18002 13823 18029
rect 13857 18002 13891 18029
rect 13925 18002 13959 18029
rect 13993 18002 14027 18029
rect 14061 18002 14095 18029
rect 14129 18002 14163 18029
rect 14197 18002 14231 18029
rect 14265 18002 14299 18029
rect 14333 18002 14367 18029
rect 13789 17995 13790 18002
rect 13857 17995 13862 18002
rect 13925 17995 13934 18002
rect 13993 17995 14006 18002
rect 14061 17995 14078 18002
rect 14129 17995 14150 18002
rect 14197 17995 14222 18002
rect 14265 17995 14294 18002
rect 14333 17995 14366 18002
rect 14401 17995 14435 18029
rect 14469 18002 14503 18029
rect 14537 18002 14571 18029
rect 14605 18002 14639 18029
rect 14673 18002 14707 18029
rect 14741 18002 14772 18029
rect 14472 17995 14503 18002
rect 14544 17995 14571 18002
rect 14616 17995 14639 18002
rect 14688 17995 14707 18002
rect 243 17968 282 17995
rect 316 17968 355 17995
rect 389 17968 428 17995
rect 462 17968 501 17995
rect 535 17968 574 17995
rect 608 17968 647 17995
rect 681 17968 720 17995
rect 754 17968 793 17995
rect 827 17968 866 17995
rect 900 17968 939 17995
rect 973 17968 1012 17995
rect 1046 17968 1085 17995
rect 1119 17968 1158 17995
rect 1192 17968 1231 17995
rect 1265 17968 1304 17995
rect 1338 17968 1377 17995
rect 1411 17968 1450 17995
rect 1484 17968 1523 17995
rect 1557 17968 1596 17995
rect 1630 17968 1669 17995
rect 1703 17968 1742 17995
rect 1776 17968 1815 17995
rect 1849 17968 1888 17995
rect 1922 17968 1961 17995
rect 1995 17968 2034 17995
rect 2068 17968 2107 17995
rect 2141 17968 2180 17995
rect 2214 17968 2253 17995
rect 2287 17968 2326 17995
rect 2360 17968 2399 17995
rect 2433 17968 2472 17995
rect 2506 17968 2545 17995
rect 2579 17968 2618 17995
rect 2652 17968 2691 17995
rect 2725 17968 2764 17995
rect 2798 17968 2837 17995
rect 2871 17968 2910 17995
rect 2944 17968 2983 17995
rect 3017 17968 3056 17995
rect 3090 17968 3129 17995
rect 3163 17968 3202 17995
rect 3236 17968 3275 17995
rect 3309 17968 3348 17995
rect 3382 17968 3421 17995
rect 3455 17968 3494 17995
rect 3528 17968 3566 17995
rect 3600 17968 3638 17995
rect 3672 17968 3710 17995
rect 3744 17968 3782 17995
rect 3816 17968 3854 17995
rect 3888 17968 3926 17995
rect 3960 17968 3998 17995
rect 4032 17968 4070 17995
rect 4104 17968 4142 17995
rect 4176 17968 4214 17995
rect 4248 17968 4286 17995
rect 4320 17968 4358 17995
rect 4392 17968 4430 17995
rect 4464 17968 4502 17995
rect 4536 17968 4574 17995
rect 4608 17968 4646 17995
rect 4680 17968 4718 17995
rect 4752 17968 4790 17995
rect 4824 17968 4862 17995
rect 4896 17968 4934 17995
rect 4968 17968 5006 17995
rect 5040 17968 5078 17995
rect 5112 17968 5150 17995
rect 5184 17968 5222 17995
rect 5256 17968 5294 17995
rect 5328 17968 5366 17995
rect 5400 17968 5438 17995
rect 5472 17968 5510 17995
rect 5544 17968 5582 17995
rect 5616 17968 5654 17995
rect 5688 17968 5726 17995
rect 5760 17968 5798 17995
rect 5832 17968 5870 17995
rect 5904 17968 5942 17995
rect 5976 17968 6014 17995
rect 6048 17968 6086 17995
rect 6120 17968 6158 17995
rect 6192 17968 6230 17995
rect 6264 17968 6302 17995
rect 6336 17968 6374 17995
rect 6408 17968 6446 17995
rect 6480 17968 6518 17995
rect 6552 17968 6590 17995
rect 6624 17968 6662 17995
rect 6696 17968 6734 17995
rect 6768 17968 6806 17995
rect 6840 17968 6878 17995
rect 6912 17968 6950 17995
rect 6984 17968 7022 17995
rect 7056 17968 7094 17995
rect 7128 17968 7166 17995
rect 7200 17968 7238 17995
rect 7272 17968 7310 17995
rect 7344 17968 7382 17995
rect 7416 17968 7454 17995
rect 7488 17968 7526 17995
rect 7560 17968 7598 17995
rect 7632 17968 7670 17995
rect 7704 17968 7742 17995
rect 7776 17968 7814 17995
rect 7848 17968 7886 17995
rect 7920 17968 7958 17995
rect 7992 17968 8030 17995
rect 8064 17968 8102 17995
rect 8136 17968 8174 17995
rect 8208 17968 8246 17995
rect 8280 17968 8318 17995
rect 8352 17968 8390 17995
rect 8424 17968 8462 17995
rect 8496 17968 8534 17995
rect 8568 17968 8606 17995
rect 8640 17968 8678 17995
rect 8712 17968 8750 17995
rect 8784 17968 8822 17995
rect 8856 17968 8894 17995
rect 8928 17968 8966 17995
rect 9000 17968 9038 17995
rect 9072 17968 9110 17995
rect 9144 17968 9182 17995
rect 9216 17968 9254 17995
rect 9288 17968 9326 17995
rect 9360 17968 9398 17995
rect 9432 17968 9470 17995
rect 9504 17968 9542 17995
rect 9576 17968 9614 17995
rect 9648 17968 9686 17995
rect 9720 17968 9758 17995
rect 9792 17968 9830 17995
rect 9864 17968 9902 17995
rect 9936 17968 9974 17995
rect 10008 17968 10046 17995
rect 10080 17968 10118 17995
rect 10152 17968 10190 17995
rect 10224 17968 10262 17995
rect 10296 17968 10334 17995
rect 10368 17968 10406 17995
rect 10440 17968 10478 17995
rect 10512 17968 10550 17995
rect 10584 17968 10622 17995
rect 10656 17968 10694 17995
rect 10728 17968 10766 17995
rect 10800 17968 10838 17995
rect 10872 17968 10910 17995
rect 10944 17968 10982 17995
rect 11016 17968 11054 17995
rect 11088 17968 11126 17995
rect 11160 17968 11198 17995
rect 11232 17968 11270 17995
rect 11304 17968 11342 17995
rect 11376 17968 11414 17995
rect 11448 17968 11486 17995
rect 11520 17968 11558 17995
rect 11592 17968 11630 17995
rect 11664 17968 11702 17995
rect 11736 17968 11774 17995
rect 11808 17968 11846 17995
rect 11880 17968 11918 17995
rect 11952 17968 11990 17995
rect 12024 17968 12062 17995
rect 12096 17968 12134 17995
rect 12168 17968 12206 17995
rect 12240 17968 12278 17995
rect 12312 17968 12350 17995
rect 12384 17968 12422 17995
rect 12456 17968 12494 17995
rect 12528 17968 12566 17995
rect 12600 17968 12638 17995
rect 12672 17968 12710 17995
rect 12744 17968 12782 17995
rect 12816 17968 12854 17995
rect 12888 17968 12926 17995
rect 12960 17968 12998 17995
rect 13032 17968 13070 17995
rect 13104 17968 13142 17995
rect 13176 17968 13214 17995
rect 13248 17968 13286 17995
rect 13320 17968 13358 17995
rect 13392 17968 13430 17995
rect 13464 17968 13502 17995
rect 13536 17968 13574 17995
rect 13608 17968 13646 17995
rect 13680 17968 13718 17995
rect 13752 17968 13790 17995
rect 13824 17968 13862 17995
rect 13896 17968 13934 17995
rect 13968 17968 14006 17995
rect 14040 17968 14078 17995
rect 14112 17968 14150 17995
rect 14184 17968 14222 17995
rect 14256 17968 14294 17995
rect 14328 17968 14366 17995
rect 14400 17968 14438 17995
rect 14472 17968 14510 17995
rect 14544 17968 14582 17995
rect 14616 17968 14654 17995
rect 14688 17968 14726 17995
rect 14760 17968 14772 18002
rect 197 17959 14772 17968
rect 197 17926 221 17959
rect 255 17926 290 17959
rect 324 17926 359 17959
rect 197 17892 209 17926
rect 255 17925 282 17926
rect 324 17925 355 17926
rect 393 17925 427 17959
rect 461 17926 495 17959
rect 529 17926 563 17959
rect 597 17926 631 17959
rect 665 17926 699 17959
rect 733 17926 767 17959
rect 801 17926 835 17959
rect 869 17926 903 17959
rect 462 17925 495 17926
rect 535 17925 563 17926
rect 608 17925 631 17926
rect 681 17925 699 17926
rect 754 17925 767 17926
rect 827 17925 835 17926
rect 900 17925 903 17926
rect 937 17926 971 17959
rect 1005 17926 1039 17959
rect 1073 17926 1107 17959
rect 1141 17926 1175 17959
rect 1209 17926 1243 17959
rect 1277 17926 1311 17959
rect 1345 17926 1379 17959
rect 937 17925 939 17926
rect 1005 17925 1012 17926
rect 1073 17925 1085 17926
rect 1141 17925 1158 17926
rect 1209 17925 1231 17926
rect 1277 17925 1304 17926
rect 1345 17925 1377 17926
rect 1413 17925 1447 17959
rect 1481 17926 1515 17959
rect 1549 17926 1583 17959
rect 1617 17926 1651 17959
rect 1685 17926 1719 17959
rect 1753 17926 1787 17959
rect 1821 17926 1855 17959
rect 1889 17926 1923 17959
rect 1484 17925 1515 17926
rect 1557 17925 1583 17926
rect 1630 17925 1651 17926
rect 1703 17925 1719 17926
rect 1776 17925 1787 17926
rect 1849 17925 1855 17926
rect 1922 17925 1923 17926
rect 1957 17926 1991 17959
rect 2025 17926 2059 17959
rect 2093 17926 2127 17959
rect 2161 17926 2195 17959
rect 2229 17926 2263 17959
rect 2297 17926 2331 17959
rect 1957 17925 1961 17926
rect 2025 17925 2034 17926
rect 2093 17925 2107 17926
rect 2161 17925 2180 17926
rect 2229 17925 2253 17926
rect 2297 17925 2326 17926
rect 2365 17925 2399 17959
rect 2433 17925 2467 17959
rect 2501 17926 2535 17959
rect 2569 17926 2603 17959
rect 2637 17926 2671 17959
rect 2705 17926 2739 17959
rect 2773 17926 2807 17959
rect 2841 17926 2875 17959
rect 2506 17925 2535 17926
rect 2579 17925 2603 17926
rect 2652 17925 2671 17926
rect 2725 17925 2739 17926
rect 2798 17925 2807 17926
rect 2871 17925 2875 17926
rect 2909 17926 2943 17959
rect 2977 17926 3011 17959
rect 3045 17926 3079 17959
rect 3113 17926 3147 17959
rect 3181 17926 3215 17959
rect 3249 17926 3283 17959
rect 3317 17926 3351 17959
rect 2909 17925 2910 17926
rect 2977 17925 2983 17926
rect 3045 17925 3056 17926
rect 3113 17925 3129 17926
rect 3181 17925 3202 17926
rect 3249 17925 3275 17926
rect 3317 17925 3348 17926
rect 3385 17925 3419 17959
rect 3453 17926 3487 17959
rect 3521 17926 3555 17959
rect 3589 17926 3623 17959
rect 3657 17926 3691 17959
rect 3725 17926 3759 17959
rect 3793 17926 3827 17959
rect 3861 17926 3895 17959
rect 3929 17926 3963 17959
rect 3455 17925 3487 17926
rect 3528 17925 3555 17926
rect 3600 17925 3623 17926
rect 3672 17925 3691 17926
rect 3744 17925 3759 17926
rect 3816 17925 3827 17926
rect 3888 17925 3895 17926
rect 3960 17925 3963 17926
rect 3997 17926 4031 17959
rect 4065 17926 4099 17959
rect 4133 17926 4167 17959
rect 4201 17926 4235 17959
rect 4269 17926 4303 17959
rect 4337 17926 4371 17959
rect 4405 17926 4439 17959
rect 4473 17926 4507 17959
rect 4541 17926 4575 17959
rect 3997 17925 3998 17926
rect 4065 17925 4070 17926
rect 4133 17925 4142 17926
rect 4201 17925 4214 17926
rect 4269 17925 4286 17926
rect 4337 17925 4358 17926
rect 4405 17925 4430 17926
rect 4473 17925 4502 17926
rect 4541 17925 4574 17926
rect 4609 17925 4643 17959
rect 4677 17926 4711 17959
rect 4745 17926 4779 17959
rect 4813 17926 4847 17959
rect 4881 17926 4915 17959
rect 4949 17926 4983 17959
rect 5017 17926 5051 17959
rect 5085 17926 5119 17959
rect 5153 17926 5187 17959
rect 4680 17925 4711 17926
rect 4752 17925 4779 17926
rect 4824 17925 4847 17926
rect 4896 17925 4915 17926
rect 4968 17925 4983 17926
rect 5040 17925 5051 17926
rect 5112 17925 5119 17926
rect 5184 17925 5187 17926
rect 5221 17926 5255 17959
rect 5289 17926 5323 17959
rect 5357 17926 5391 17959
rect 5425 17926 5459 17959
rect 5493 17926 5527 17959
rect 5561 17926 5595 17959
rect 5629 17926 5663 17959
rect 5697 17926 5731 17959
rect 5765 17926 5799 17959
rect 5221 17925 5222 17926
rect 5289 17925 5294 17926
rect 5357 17925 5366 17926
rect 5425 17925 5438 17926
rect 5493 17925 5510 17926
rect 5561 17925 5582 17926
rect 5629 17925 5654 17926
rect 5697 17925 5726 17926
rect 5765 17925 5798 17926
rect 5833 17925 5867 17959
rect 5901 17926 5935 17959
rect 5969 17926 6003 17959
rect 6037 17926 6071 17959
rect 6105 17926 6139 17959
rect 6173 17926 6207 17959
rect 6241 17926 6275 17959
rect 6309 17926 6343 17959
rect 6377 17926 6411 17959
rect 5904 17925 5935 17926
rect 5976 17925 6003 17926
rect 6048 17925 6071 17926
rect 6120 17925 6139 17926
rect 6192 17925 6207 17926
rect 6264 17925 6275 17926
rect 6336 17925 6343 17926
rect 6408 17925 6411 17926
rect 6445 17926 6479 17959
rect 6513 17926 6547 17959
rect 6581 17926 6615 17959
rect 6649 17926 6683 17959
rect 6717 17926 6751 17959
rect 6785 17926 6819 17959
rect 6853 17926 6887 17959
rect 6921 17926 6955 17959
rect 6989 17926 7023 17959
rect 6445 17925 6446 17926
rect 6513 17925 6518 17926
rect 6581 17925 6590 17926
rect 6649 17925 6662 17926
rect 6717 17925 6734 17926
rect 6785 17925 6806 17926
rect 6853 17925 6878 17926
rect 6921 17925 6950 17926
rect 6989 17925 7022 17926
rect 7057 17925 7091 17959
rect 7125 17926 7159 17959
rect 7193 17926 7227 17959
rect 7261 17926 7295 17959
rect 7329 17926 7363 17959
rect 7397 17926 7431 17959
rect 7465 17926 7499 17959
rect 7533 17926 7567 17959
rect 7601 17926 7635 17959
rect 7128 17925 7159 17926
rect 7200 17925 7227 17926
rect 7272 17925 7295 17926
rect 7344 17925 7363 17926
rect 7416 17925 7431 17926
rect 7488 17925 7499 17926
rect 7560 17925 7567 17926
rect 7632 17925 7635 17926
rect 7669 17926 7703 17959
rect 7737 17926 7771 17959
rect 7805 17926 7839 17959
rect 7873 17926 7907 17959
rect 7941 17926 7975 17959
rect 8009 17926 8043 17959
rect 8077 17926 8111 17959
rect 8145 17926 8179 17959
rect 8213 17926 8247 17959
rect 7669 17925 7670 17926
rect 7737 17925 7742 17926
rect 7805 17925 7814 17926
rect 7873 17925 7886 17926
rect 7941 17925 7958 17926
rect 8009 17925 8030 17926
rect 8077 17925 8102 17926
rect 8145 17925 8174 17926
rect 8213 17925 8246 17926
rect 8281 17925 8315 17959
rect 8349 17926 8383 17959
rect 8417 17926 8451 17959
rect 8485 17926 8519 17959
rect 8553 17926 8587 17959
rect 8621 17926 8655 17959
rect 8689 17926 8723 17959
rect 8757 17926 8791 17959
rect 8825 17926 8859 17959
rect 8352 17925 8383 17926
rect 8424 17925 8451 17926
rect 8496 17925 8519 17926
rect 8568 17925 8587 17926
rect 8640 17925 8655 17926
rect 8712 17925 8723 17926
rect 8784 17925 8791 17926
rect 8856 17925 8859 17926
rect 8893 17926 8927 17959
rect 8961 17926 8995 17959
rect 9029 17926 9063 17959
rect 9097 17926 9131 17959
rect 9165 17926 9199 17959
rect 9233 17926 9267 17959
rect 9301 17926 9335 17959
rect 9369 17926 9403 17959
rect 9437 17926 9471 17959
rect 8893 17925 8894 17926
rect 8961 17925 8966 17926
rect 9029 17925 9038 17926
rect 9097 17925 9110 17926
rect 9165 17925 9182 17926
rect 9233 17925 9254 17926
rect 9301 17925 9326 17926
rect 9369 17925 9398 17926
rect 9437 17925 9470 17926
rect 9505 17925 9539 17959
rect 9573 17926 9607 17959
rect 9641 17926 9675 17959
rect 9709 17926 9743 17959
rect 9777 17926 9811 17959
rect 9845 17926 9879 17959
rect 9913 17926 9947 17959
rect 9981 17926 10015 17959
rect 10049 17926 10083 17959
rect 9576 17925 9607 17926
rect 9648 17925 9675 17926
rect 9720 17925 9743 17926
rect 9792 17925 9811 17926
rect 9864 17925 9879 17926
rect 9936 17925 9947 17926
rect 10008 17925 10015 17926
rect 10080 17925 10083 17926
rect 10117 17926 10151 17959
rect 10185 17926 10219 17959
rect 10253 17926 10287 17959
rect 10321 17926 10355 17959
rect 10389 17926 10423 17959
rect 10457 17926 10491 17959
rect 10525 17926 10559 17959
rect 10593 17926 10627 17959
rect 10661 17926 10695 17959
rect 10117 17925 10118 17926
rect 10185 17925 10190 17926
rect 10253 17925 10262 17926
rect 10321 17925 10334 17926
rect 10389 17925 10406 17926
rect 10457 17925 10478 17926
rect 10525 17925 10550 17926
rect 10593 17925 10622 17926
rect 10661 17925 10694 17926
rect 10729 17925 10763 17959
rect 10797 17926 10831 17959
rect 10865 17926 10899 17959
rect 10933 17926 10967 17959
rect 11001 17926 11035 17959
rect 11069 17926 11103 17959
rect 11137 17926 11171 17959
rect 11205 17926 11239 17959
rect 11273 17926 11307 17959
rect 10800 17925 10831 17926
rect 10872 17925 10899 17926
rect 10944 17925 10967 17926
rect 11016 17925 11035 17926
rect 11088 17925 11103 17926
rect 11160 17925 11171 17926
rect 11232 17925 11239 17926
rect 11304 17925 11307 17926
rect 11341 17926 11375 17959
rect 11409 17926 11443 17959
rect 11477 17926 11511 17959
rect 11545 17926 11579 17959
rect 11613 17926 11647 17959
rect 11681 17926 11715 17959
rect 11749 17926 11783 17959
rect 11817 17926 11851 17959
rect 11885 17926 11919 17959
rect 11341 17925 11342 17926
rect 11409 17925 11414 17926
rect 11477 17925 11486 17926
rect 11545 17925 11558 17926
rect 11613 17925 11630 17926
rect 11681 17925 11702 17926
rect 11749 17925 11774 17926
rect 11817 17925 11846 17926
rect 11885 17925 11918 17926
rect 11953 17925 11987 17959
rect 12021 17926 12055 17959
rect 12089 17926 12123 17959
rect 12157 17926 12191 17959
rect 12225 17926 12259 17959
rect 12293 17926 12327 17959
rect 12361 17926 12395 17959
rect 12429 17926 12463 17959
rect 12497 17926 12531 17959
rect 12024 17925 12055 17926
rect 12096 17925 12123 17926
rect 12168 17925 12191 17926
rect 12240 17925 12259 17926
rect 12312 17925 12327 17926
rect 12384 17925 12395 17926
rect 12456 17925 12463 17926
rect 12528 17925 12531 17926
rect 12565 17926 12599 17959
rect 12633 17926 12667 17959
rect 12701 17926 12735 17959
rect 12769 17926 12803 17959
rect 12837 17926 12871 17959
rect 12905 17926 12939 17959
rect 12973 17926 13007 17959
rect 13041 17926 13075 17959
rect 13109 17926 13143 17959
rect 12565 17925 12566 17926
rect 12633 17925 12638 17926
rect 12701 17925 12710 17926
rect 12769 17925 12782 17926
rect 12837 17925 12854 17926
rect 12905 17925 12926 17926
rect 12973 17925 12998 17926
rect 13041 17925 13070 17926
rect 13109 17925 13142 17926
rect 13177 17925 13211 17959
rect 13245 17926 13279 17959
rect 13313 17926 13347 17959
rect 13381 17926 13415 17959
rect 13449 17926 13483 17959
rect 13517 17926 13551 17959
rect 13585 17926 13619 17959
rect 13653 17926 13687 17959
rect 13721 17926 13755 17959
rect 13248 17925 13279 17926
rect 13320 17925 13347 17926
rect 13392 17925 13415 17926
rect 13464 17925 13483 17926
rect 13536 17925 13551 17926
rect 13608 17925 13619 17926
rect 13680 17925 13687 17926
rect 13752 17925 13755 17926
rect 13789 17926 13823 17959
rect 13857 17926 13891 17959
rect 13925 17926 13959 17959
rect 13993 17926 14027 17959
rect 14061 17926 14095 17959
rect 14129 17926 14163 17959
rect 14197 17926 14231 17959
rect 14265 17926 14299 17959
rect 14333 17926 14367 17959
rect 13789 17925 13790 17926
rect 13857 17925 13862 17926
rect 13925 17925 13934 17926
rect 13993 17925 14006 17926
rect 14061 17925 14078 17926
rect 14129 17925 14150 17926
rect 14197 17925 14222 17926
rect 14265 17925 14294 17926
rect 14333 17925 14366 17926
rect 14401 17925 14435 17959
rect 14469 17926 14503 17959
rect 14537 17926 14571 17959
rect 14605 17926 14639 17959
rect 14673 17926 14707 17959
rect 14741 17926 14772 17959
rect 14472 17925 14503 17926
rect 14544 17925 14571 17926
rect 14616 17925 14639 17926
rect 14688 17925 14707 17926
rect 243 17892 282 17925
rect 316 17892 355 17925
rect 389 17892 428 17925
rect 462 17892 501 17925
rect 535 17892 574 17925
rect 608 17892 647 17925
rect 681 17892 720 17925
rect 754 17892 793 17925
rect 827 17892 866 17925
rect 900 17892 939 17925
rect 973 17892 1012 17925
rect 1046 17892 1085 17925
rect 1119 17892 1158 17925
rect 1192 17892 1231 17925
rect 1265 17892 1304 17925
rect 1338 17892 1377 17925
rect 1411 17892 1450 17925
rect 1484 17892 1523 17925
rect 1557 17892 1596 17925
rect 1630 17892 1669 17925
rect 1703 17892 1742 17925
rect 1776 17892 1815 17925
rect 1849 17892 1888 17925
rect 1922 17892 1961 17925
rect 1995 17892 2034 17925
rect 2068 17892 2107 17925
rect 2141 17892 2180 17925
rect 2214 17892 2253 17925
rect 2287 17892 2326 17925
rect 2360 17892 2399 17925
rect 2433 17892 2472 17925
rect 2506 17892 2545 17925
rect 2579 17892 2618 17925
rect 2652 17892 2691 17925
rect 2725 17892 2764 17925
rect 2798 17892 2837 17925
rect 2871 17892 2910 17925
rect 2944 17892 2983 17925
rect 3017 17892 3056 17925
rect 3090 17892 3129 17925
rect 3163 17892 3202 17925
rect 3236 17892 3275 17925
rect 3309 17892 3348 17925
rect 3382 17892 3421 17925
rect 3455 17892 3494 17925
rect 3528 17892 3566 17925
rect 3600 17892 3638 17925
rect 3672 17892 3710 17925
rect 3744 17892 3782 17925
rect 3816 17892 3854 17925
rect 3888 17892 3926 17925
rect 3960 17892 3998 17925
rect 4032 17892 4070 17925
rect 4104 17892 4142 17925
rect 4176 17892 4214 17925
rect 4248 17892 4286 17925
rect 4320 17892 4358 17925
rect 4392 17892 4430 17925
rect 4464 17892 4502 17925
rect 4536 17892 4574 17925
rect 4608 17892 4646 17925
rect 4680 17892 4718 17925
rect 4752 17892 4790 17925
rect 4824 17892 4862 17925
rect 4896 17892 4934 17925
rect 4968 17892 5006 17925
rect 5040 17892 5078 17925
rect 5112 17892 5150 17925
rect 5184 17892 5222 17925
rect 5256 17892 5294 17925
rect 5328 17892 5366 17925
rect 5400 17892 5438 17925
rect 5472 17892 5510 17925
rect 5544 17892 5582 17925
rect 5616 17892 5654 17925
rect 5688 17892 5726 17925
rect 5760 17892 5798 17925
rect 5832 17892 5870 17925
rect 5904 17892 5942 17925
rect 5976 17892 6014 17925
rect 6048 17892 6086 17925
rect 6120 17892 6158 17925
rect 6192 17892 6230 17925
rect 6264 17892 6302 17925
rect 6336 17892 6374 17925
rect 6408 17892 6446 17925
rect 6480 17892 6518 17925
rect 6552 17892 6590 17925
rect 6624 17892 6662 17925
rect 6696 17892 6734 17925
rect 6768 17892 6806 17925
rect 6840 17892 6878 17925
rect 6912 17892 6950 17925
rect 6984 17892 7022 17925
rect 7056 17892 7094 17925
rect 7128 17892 7166 17925
rect 7200 17892 7238 17925
rect 7272 17892 7310 17925
rect 7344 17892 7382 17925
rect 7416 17892 7454 17925
rect 7488 17892 7526 17925
rect 7560 17892 7598 17925
rect 7632 17892 7670 17925
rect 7704 17892 7742 17925
rect 7776 17892 7814 17925
rect 7848 17892 7886 17925
rect 7920 17892 7958 17925
rect 7992 17892 8030 17925
rect 8064 17892 8102 17925
rect 8136 17892 8174 17925
rect 8208 17892 8246 17925
rect 8280 17892 8318 17925
rect 8352 17892 8390 17925
rect 8424 17892 8462 17925
rect 8496 17892 8534 17925
rect 8568 17892 8606 17925
rect 8640 17892 8678 17925
rect 8712 17892 8750 17925
rect 8784 17892 8822 17925
rect 8856 17892 8894 17925
rect 8928 17892 8966 17925
rect 9000 17892 9038 17925
rect 9072 17892 9110 17925
rect 9144 17892 9182 17925
rect 9216 17892 9254 17925
rect 9288 17892 9326 17925
rect 9360 17892 9398 17925
rect 9432 17892 9470 17925
rect 9504 17892 9542 17925
rect 9576 17892 9614 17925
rect 9648 17892 9686 17925
rect 9720 17892 9758 17925
rect 9792 17892 9830 17925
rect 9864 17892 9902 17925
rect 9936 17892 9974 17925
rect 10008 17892 10046 17925
rect 10080 17892 10118 17925
rect 10152 17892 10190 17925
rect 10224 17892 10262 17925
rect 10296 17892 10334 17925
rect 10368 17892 10406 17925
rect 10440 17892 10478 17925
rect 10512 17892 10550 17925
rect 10584 17892 10622 17925
rect 10656 17892 10694 17925
rect 10728 17892 10766 17925
rect 10800 17892 10838 17925
rect 10872 17892 10910 17925
rect 10944 17892 10982 17925
rect 11016 17892 11054 17925
rect 11088 17892 11126 17925
rect 11160 17892 11198 17925
rect 11232 17892 11270 17925
rect 11304 17892 11342 17925
rect 11376 17892 11414 17925
rect 11448 17892 11486 17925
rect 11520 17892 11558 17925
rect 11592 17892 11630 17925
rect 11664 17892 11702 17925
rect 11736 17892 11774 17925
rect 11808 17892 11846 17925
rect 11880 17892 11918 17925
rect 11952 17892 11990 17925
rect 12024 17892 12062 17925
rect 12096 17892 12134 17925
rect 12168 17892 12206 17925
rect 12240 17892 12278 17925
rect 12312 17892 12350 17925
rect 12384 17892 12422 17925
rect 12456 17892 12494 17925
rect 12528 17892 12566 17925
rect 12600 17892 12638 17925
rect 12672 17892 12710 17925
rect 12744 17892 12782 17925
rect 12816 17892 12854 17925
rect 12888 17892 12926 17925
rect 12960 17892 12998 17925
rect 13032 17892 13070 17925
rect 13104 17892 13142 17925
rect 13176 17892 13214 17925
rect 13248 17892 13286 17925
rect 13320 17892 13358 17925
rect 13392 17892 13430 17925
rect 13464 17892 13502 17925
rect 13536 17892 13574 17925
rect 13608 17892 13646 17925
rect 13680 17892 13718 17925
rect 13752 17892 13790 17925
rect 13824 17892 13862 17925
rect 13896 17892 13934 17925
rect 13968 17892 14006 17925
rect 14040 17892 14078 17925
rect 14112 17892 14150 17925
rect 14184 17892 14222 17925
rect 14256 17892 14294 17925
rect 14328 17892 14366 17925
rect 14400 17892 14438 17925
rect 14472 17892 14510 17925
rect 14544 17892 14582 17925
rect 14616 17892 14654 17925
rect 14688 17892 14726 17925
rect 14760 17892 14772 17926
rect 197 17889 14772 17892
rect 197 17855 221 17889
rect 255 17855 290 17889
rect 324 17855 359 17889
rect 393 17855 427 17889
rect 461 17855 495 17889
rect 529 17855 563 17889
rect 597 17855 631 17889
rect 665 17855 699 17889
rect 733 17855 767 17889
rect 801 17855 835 17889
rect 869 17855 903 17889
rect 937 17855 971 17889
rect 1005 17855 1039 17889
rect 1073 17855 1107 17889
rect 1141 17855 1175 17889
rect 1209 17855 1243 17889
rect 1277 17855 1311 17889
rect 1345 17855 1379 17889
rect 1413 17855 1447 17889
rect 1481 17855 1515 17889
rect 1549 17855 1583 17889
rect 1617 17855 1651 17889
rect 1685 17855 1719 17889
rect 1753 17855 1787 17889
rect 1821 17855 1855 17889
rect 1889 17855 1923 17889
rect 1957 17855 1991 17889
rect 2025 17855 2059 17889
rect 2093 17855 2127 17889
rect 2161 17855 2195 17889
rect 2229 17855 2263 17889
rect 2297 17855 2331 17889
rect 2365 17855 2399 17889
rect 2433 17855 2467 17889
rect 2501 17855 2535 17889
rect 2569 17855 2603 17889
rect 2637 17855 2671 17889
rect 2705 17855 2739 17889
rect 2773 17855 2807 17889
rect 2841 17855 2875 17889
rect 2909 17855 2943 17889
rect 2977 17855 3011 17889
rect 3045 17855 3079 17889
rect 3113 17855 3147 17889
rect 3181 17855 3215 17889
rect 3249 17855 3283 17889
rect 3317 17855 3351 17889
rect 3385 17855 3419 17889
rect 3453 17855 3487 17889
rect 3521 17855 3555 17889
rect 3589 17855 3623 17889
rect 3657 17855 3691 17889
rect 3725 17855 3759 17889
rect 3793 17855 3827 17889
rect 3861 17855 3895 17889
rect 3929 17855 3963 17889
rect 3997 17855 4031 17889
rect 4065 17855 4099 17889
rect 4133 17855 4167 17889
rect 4201 17855 4235 17889
rect 4269 17855 4303 17889
rect 4337 17855 4371 17889
rect 4405 17855 4439 17889
rect 4473 17855 4507 17889
rect 4541 17855 4575 17889
rect 4609 17855 4643 17889
rect 4677 17855 4711 17889
rect 4745 17855 4779 17889
rect 4813 17855 4847 17889
rect 4881 17855 4915 17889
rect 4949 17855 4983 17889
rect 5017 17855 5051 17889
rect 5085 17855 5119 17889
rect 5153 17855 5187 17889
rect 5221 17855 5255 17889
rect 5289 17855 5323 17889
rect 5357 17855 5391 17889
rect 5425 17855 5459 17889
rect 5493 17855 5527 17889
rect 5561 17855 5595 17889
rect 5629 17855 5663 17889
rect 5697 17855 5731 17889
rect 5765 17855 5799 17889
rect 5833 17855 5867 17889
rect 5901 17855 5935 17889
rect 5969 17855 6003 17889
rect 6037 17855 6071 17889
rect 6105 17855 6139 17889
rect 6173 17855 6207 17889
rect 6241 17855 6275 17889
rect 6309 17855 6343 17889
rect 6377 17855 6411 17889
rect 6445 17855 6479 17889
rect 6513 17855 6547 17889
rect 6581 17855 6615 17889
rect 6649 17855 6683 17889
rect 6717 17855 6751 17889
rect 6785 17855 6819 17889
rect 6853 17855 6887 17889
rect 6921 17855 6955 17889
rect 6989 17855 7023 17889
rect 7057 17855 7091 17889
rect 7125 17855 7159 17889
rect 7193 17855 7227 17889
rect 7261 17855 7295 17889
rect 7329 17855 7363 17889
rect 7397 17855 7431 17889
rect 7465 17855 7499 17889
rect 7533 17855 7567 17889
rect 7601 17855 7635 17889
rect 7669 17855 7703 17889
rect 7737 17855 7771 17889
rect 7805 17855 7839 17889
rect 7873 17855 7907 17889
rect 7941 17855 7975 17889
rect 8009 17855 8043 17889
rect 8077 17855 8111 17889
rect 8145 17855 8179 17889
rect 8213 17855 8247 17889
rect 8281 17855 8315 17889
rect 8349 17855 8383 17889
rect 8417 17855 8451 17889
rect 8485 17855 8519 17889
rect 8553 17855 8587 17889
rect 8621 17855 8655 17889
rect 8689 17855 8723 17889
rect 8757 17855 8791 17889
rect 8825 17855 8859 17889
rect 8893 17855 8927 17889
rect 8961 17855 8995 17889
rect 9029 17855 9063 17889
rect 9097 17855 9131 17889
rect 9165 17855 9199 17889
rect 9233 17855 9267 17889
rect 9301 17855 9335 17889
rect 9369 17855 9403 17889
rect 9437 17855 9471 17889
rect 9505 17855 9539 17889
rect 9573 17855 9607 17889
rect 9641 17855 9675 17889
rect 9709 17855 9743 17889
rect 9777 17855 9811 17889
rect 9845 17855 9879 17889
rect 9913 17855 9947 17889
rect 9981 17855 10015 17889
rect 10049 17855 10083 17889
rect 10117 17855 10151 17889
rect 10185 17855 10219 17889
rect 10253 17855 10287 17889
rect 10321 17855 10355 17889
rect 10389 17855 10423 17889
rect 10457 17855 10491 17889
rect 10525 17855 10559 17889
rect 10593 17855 10627 17889
rect 10661 17855 10695 17889
rect 10729 17855 10763 17889
rect 10797 17855 10831 17889
rect 10865 17855 10899 17889
rect 10933 17855 10967 17889
rect 11001 17855 11035 17889
rect 11069 17855 11103 17889
rect 11137 17855 11171 17889
rect 11205 17855 11239 17889
rect 11273 17855 11307 17889
rect 11341 17855 11375 17889
rect 11409 17855 11443 17889
rect 11477 17855 11511 17889
rect 11545 17855 11579 17889
rect 11613 17855 11647 17889
rect 11681 17855 11715 17889
rect 11749 17855 11783 17889
rect 11817 17855 11851 17889
rect 11885 17855 11919 17889
rect 11953 17855 11987 17889
rect 12021 17855 12055 17889
rect 12089 17855 12123 17889
rect 12157 17855 12191 17889
rect 12225 17855 12259 17889
rect 12293 17855 12327 17889
rect 12361 17855 12395 17889
rect 12429 17855 12463 17889
rect 12497 17855 12531 17889
rect 12565 17855 12599 17889
rect 12633 17855 12667 17889
rect 12701 17855 12735 17889
rect 12769 17855 12803 17889
rect 12837 17855 12871 17889
rect 12905 17855 12939 17889
rect 12973 17855 13007 17889
rect 13041 17855 13075 17889
rect 13109 17855 13143 17889
rect 13177 17855 13211 17889
rect 13245 17855 13279 17889
rect 13313 17855 13347 17889
rect 13381 17855 13415 17889
rect 13449 17855 13483 17889
rect 13517 17855 13551 17889
rect 13585 17855 13619 17889
rect 13653 17855 13687 17889
rect 13721 17855 13755 17889
rect 13789 17855 13823 17889
rect 13857 17855 13891 17889
rect 13925 17855 13959 17889
rect 13993 17855 14027 17889
rect 14061 17855 14095 17889
rect 14129 17855 14163 17889
rect 14197 17855 14231 17889
rect 14265 17855 14299 17889
rect 14333 17855 14367 17889
rect 14401 17855 14435 17889
rect 14469 17855 14503 17889
rect 14537 17855 14571 17889
rect 14605 17855 14639 17889
rect 14673 17855 14707 17889
rect 14741 17855 14772 17889
<< viali >>
rect 112 28113 121 28122
rect 121 28113 146 28122
rect 185 28113 190 28122
rect 190 28113 219 28122
rect 258 28113 259 28122
rect 259 28113 292 28122
rect 331 28113 362 28122
rect 362 28113 365 28122
rect 404 28113 431 28122
rect 431 28113 438 28122
rect 477 28113 500 28122
rect 500 28113 511 28122
rect 550 28113 569 28122
rect 569 28113 584 28122
rect 623 28113 638 28122
rect 638 28113 657 28122
rect 696 28113 707 28122
rect 707 28113 730 28122
rect 769 28113 776 28122
rect 776 28113 803 28122
rect 842 28113 845 28122
rect 845 28113 876 28122
rect 112 28088 146 28113
rect 185 28088 219 28113
rect 258 28088 292 28113
rect 331 28088 365 28113
rect 404 28088 438 28113
rect 477 28088 511 28113
rect 550 28088 584 28113
rect 623 28088 657 28113
rect 696 28088 730 28113
rect 769 28088 803 28113
rect 842 28088 876 28113
rect 915 28088 949 28122
rect 988 28113 1018 28122
rect 1018 28113 1022 28122
rect 1061 28113 1087 28122
rect 1087 28113 1095 28122
rect 988 28088 1022 28113
rect 1061 28088 1095 28113
rect 1134 28088 1156 28122
rect 1156 28088 1168 28122
rect 1207 28088 1241 28122
rect 1280 28088 1314 28122
rect 1353 28088 1387 28122
rect 1426 28088 1460 28122
rect 1499 28088 1533 28122
rect 1571 28088 1605 28122
rect 1643 28088 1677 28122
rect 1715 28088 1749 28122
rect 1787 28088 1821 28122
rect 1859 28088 1893 28122
rect 1931 28088 1965 28122
rect 2003 28088 2037 28122
rect 2075 28088 2109 28122
rect 2147 28088 2181 28122
rect 2219 28088 2253 28122
rect 2291 28088 2325 28122
rect 2363 28088 2397 28122
rect 2435 28088 2469 28122
rect 2507 28088 2541 28122
rect 2579 28088 2613 28122
rect 2651 28088 2685 28122
rect 2723 28088 2757 28122
rect 2795 28088 2829 28122
rect 2867 28088 2901 28122
rect 2939 28088 2973 28122
rect 3011 28088 3045 28122
rect 3083 28088 3117 28122
rect 3155 28088 3189 28122
rect 3227 28088 3261 28122
rect 3299 28088 3333 28122
rect 3371 28088 3405 28122
rect 3443 28088 3477 28122
rect 3515 28088 3549 28122
rect 3587 28088 3621 28122
rect 3659 28088 3693 28122
rect 3731 28088 3765 28122
rect 3803 28088 3837 28122
rect 3875 28088 3909 28122
rect 3947 28088 3981 28122
rect 4019 28088 4053 28122
rect 4091 28088 4125 28122
rect 4163 28088 4197 28122
rect 4235 28088 4269 28122
rect 4307 28088 4341 28122
rect 4379 28088 4413 28122
rect 4451 28088 4485 28122
rect 4523 28088 4557 28122
rect 4595 28088 4629 28122
rect 4667 28088 4701 28122
rect 4739 28088 4773 28122
rect 4811 28088 4845 28122
rect 4883 28088 4917 28122
rect 4955 28088 4989 28122
rect 5027 28088 5061 28122
rect 5099 28088 5133 28122
rect 5171 28088 5205 28122
rect 5243 28088 5277 28122
rect 5315 28088 5349 28122
rect 5387 28088 5421 28122
rect 5459 28088 5493 28122
rect 5531 28088 5565 28122
rect 5603 28088 5637 28122
rect 5675 28088 5709 28122
rect 5747 28088 5781 28122
rect 5819 28088 5853 28122
rect 5891 28088 5925 28122
rect 5963 28088 5997 28122
rect 6035 28088 6069 28122
rect 6107 28088 6141 28122
rect 6179 28088 6213 28122
rect 6251 28088 6285 28122
rect 6323 28088 6357 28122
rect 6395 28088 6429 28122
rect 6467 28088 6501 28122
rect 6539 28088 6573 28122
rect 6611 28088 6645 28122
rect 6683 28088 6717 28122
rect 6755 28088 6789 28122
rect 6827 28088 6861 28122
rect 6899 28088 6933 28122
rect 6971 28088 7005 28122
rect 7043 28088 7077 28122
rect 7115 28088 7149 28122
rect 7187 28088 7221 28122
rect 7259 28088 7293 28122
rect 7331 28088 7365 28122
rect 7403 28088 7437 28122
rect 7475 28088 7509 28122
rect 7547 28088 7581 28122
rect 7619 28088 7653 28122
rect 7691 28088 7725 28122
rect 7763 28088 7797 28122
rect 7835 28088 7869 28122
rect 7907 28088 7941 28122
rect 7979 28088 8013 28122
rect 8051 28088 8085 28122
rect 8123 28088 8157 28122
rect 8195 28088 8229 28122
rect 8267 28088 8301 28122
rect 8339 28088 8373 28122
rect 8411 28088 8445 28122
rect 8483 28088 8517 28122
rect 8555 28088 8589 28122
rect 8627 28088 8661 28122
rect 8699 28088 8733 28122
rect 8771 28088 8805 28122
rect 8843 28088 8877 28122
rect 8915 28088 8949 28122
rect 8987 28088 9021 28122
rect 9059 28088 9093 28122
rect 9131 28088 9165 28122
rect 9203 28088 9237 28122
rect 9275 28088 9309 28122
rect 9347 28088 9381 28122
rect 9419 28088 9453 28122
rect 9491 28088 9525 28122
rect 9563 28088 9597 28122
rect 9635 28088 9669 28122
rect 9707 28088 9741 28122
rect 9779 28088 9813 28122
rect 9851 28088 9885 28122
rect 9923 28088 9957 28122
rect 9995 28088 10029 28122
rect 10067 28088 10101 28122
rect 10139 28088 10173 28122
rect 10211 28088 10245 28122
rect 10283 28088 10317 28122
rect 10355 28088 10389 28122
rect 10427 28088 10461 28122
rect 10499 28088 10533 28122
rect 10571 28088 10605 28122
rect 10643 28088 10677 28122
rect 10715 28088 10749 28122
rect 10787 28088 10821 28122
rect 10859 28088 10893 28122
rect 10931 28088 10965 28122
rect 11003 28088 11037 28122
rect 11075 28088 11109 28122
rect 11147 28088 11181 28122
rect 11219 28088 11253 28122
rect 11291 28088 11325 28122
rect 11363 28088 11397 28122
rect 11435 28088 11469 28122
rect 11507 28088 11541 28122
rect 11579 28088 11613 28122
rect 11651 28088 11685 28122
rect 11723 28088 11757 28122
rect 11795 28088 11829 28122
rect 11867 28088 11901 28122
rect 11939 28088 11973 28122
rect 12011 28088 12045 28122
rect 12083 28088 12117 28122
rect 12155 28088 12189 28122
rect 12227 28088 12261 28122
rect 12299 28088 12333 28122
rect 12371 28088 12405 28122
rect 12443 28088 12477 28122
rect 12515 28088 12549 28122
rect 12587 28088 12621 28122
rect 12659 28088 12693 28122
rect 12731 28088 12765 28122
rect 12803 28088 12837 28122
rect 12875 28088 12909 28122
rect 12947 28088 12981 28122
rect 13019 28088 13053 28122
rect 13091 28088 13125 28122
rect 13163 28088 13197 28122
rect 13235 28088 13269 28122
rect 13307 28088 13341 28122
rect 13379 28088 13413 28122
rect 13451 28088 13485 28122
rect 13523 28088 13557 28122
rect 13595 28088 13629 28122
rect 13667 28088 13701 28122
rect 13739 28088 13773 28122
rect 13811 28088 13845 28122
rect 13883 28088 13917 28122
rect 112 28011 146 28040
rect 185 28011 219 28040
rect 258 28011 292 28040
rect 331 28011 365 28040
rect 404 28011 438 28040
rect 477 28011 511 28040
rect 550 28011 584 28040
rect 623 28011 657 28040
rect 696 28011 730 28040
rect 769 28011 803 28040
rect 842 28011 876 28040
rect 112 28006 121 28011
rect 121 28006 146 28011
rect 185 28006 190 28011
rect 190 28006 219 28011
rect 258 28006 259 28011
rect 259 28006 292 28011
rect 331 28006 362 28011
rect 362 28006 365 28011
rect 404 28006 431 28011
rect 431 28006 438 28011
rect 477 28006 500 28011
rect 500 28006 511 28011
rect 550 28006 569 28011
rect 569 28006 584 28011
rect 623 28006 638 28011
rect 638 28006 657 28011
rect 696 28006 707 28011
rect 707 28006 730 28011
rect 769 28006 776 28011
rect 776 28006 803 28011
rect 842 28006 845 28011
rect 845 28006 876 28011
rect 915 28006 949 28040
rect 988 28011 1022 28040
rect 1061 28011 1095 28040
rect 988 28006 1018 28011
rect 1018 28006 1022 28011
rect 1061 28006 1087 28011
rect 1087 28006 1095 28011
rect 1134 28006 1156 28040
rect 1156 28006 1168 28040
rect 1207 28006 1241 28040
rect 1280 28006 1314 28040
rect 1353 28006 1387 28040
rect 1426 28006 1460 28040
rect 1499 28006 1533 28040
rect 1571 28006 1605 28040
rect 1643 28006 1677 28040
rect 1715 28006 1749 28040
rect 1787 28006 1821 28040
rect 1859 28006 1893 28040
rect 1931 28006 1965 28040
rect 2003 28006 2037 28040
rect 2075 28006 2109 28040
rect 2147 28006 2181 28040
rect 2219 28006 2253 28040
rect 2291 28006 2325 28040
rect 2363 28006 2397 28040
rect 2435 28006 2469 28040
rect 2507 28006 2541 28040
rect 2579 28006 2613 28040
rect 2651 28006 2685 28040
rect 2723 28006 2757 28040
rect 2795 28006 2829 28040
rect 2867 28006 2901 28040
rect 2939 28006 2973 28040
rect 3011 28006 3045 28040
rect 3083 28006 3117 28040
rect 3155 28006 3189 28040
rect 3227 28006 3261 28040
rect 3299 28006 3333 28040
rect 3371 28006 3405 28040
rect 3443 28006 3477 28040
rect 3515 28006 3549 28040
rect 3587 28006 3621 28040
rect 3659 28006 3693 28040
rect 3731 28006 3765 28040
rect 3803 28006 3837 28040
rect 3875 28006 3909 28040
rect 3947 28006 3981 28040
rect 4019 28006 4053 28040
rect 4091 28006 4125 28040
rect 4163 28006 4197 28040
rect 4235 28006 4269 28040
rect 4307 28006 4341 28040
rect 4379 28006 4413 28040
rect 4451 28006 4485 28040
rect 4523 28006 4557 28040
rect 4595 28006 4629 28040
rect 4667 28006 4701 28040
rect 4739 28006 4773 28040
rect 4811 28006 4845 28040
rect 4883 28006 4917 28040
rect 4955 28006 4989 28040
rect 5027 28006 5061 28040
rect 5099 28006 5133 28040
rect 5171 28006 5205 28040
rect 5243 28006 5277 28040
rect 5315 28006 5349 28040
rect 5387 28006 5421 28040
rect 5459 28006 5493 28040
rect 5531 28006 5565 28040
rect 5603 28006 5637 28040
rect 5675 28006 5709 28040
rect 5747 28006 5781 28040
rect 5819 28006 5853 28040
rect 5891 28006 5925 28040
rect 5963 28006 5997 28040
rect 6035 28006 6069 28040
rect 6107 28006 6141 28040
rect 6179 28006 6213 28040
rect 6251 28006 6285 28040
rect 6323 28006 6357 28040
rect 6395 28006 6429 28040
rect 6467 28006 6501 28040
rect 6539 28006 6573 28040
rect 6611 28006 6645 28040
rect 6683 28006 6717 28040
rect 6755 28006 6789 28040
rect 6827 28006 6861 28040
rect 6899 28006 6933 28040
rect 6971 28006 7005 28040
rect 7043 28006 7077 28040
rect 7115 28006 7149 28040
rect 7187 28006 7221 28040
rect 7259 28006 7293 28040
rect 7331 28006 7365 28040
rect 7403 28006 7437 28040
rect 7475 28006 7509 28040
rect 7547 28006 7581 28040
rect 7619 28006 7653 28040
rect 7691 28006 7725 28040
rect 7763 28006 7797 28040
rect 7835 28006 7869 28040
rect 7907 28006 7941 28040
rect 7979 28006 8013 28040
rect 8051 28006 8085 28040
rect 8123 28006 8157 28040
rect 8195 28006 8229 28040
rect 8267 28006 8301 28040
rect 8339 28006 8373 28040
rect 8411 28006 8445 28040
rect 8483 28006 8517 28040
rect 8555 28006 8589 28040
rect 8627 28006 8661 28040
rect 8699 28006 8733 28040
rect 8771 28006 8805 28040
rect 8843 28006 8877 28040
rect 8915 28006 8949 28040
rect 8987 28006 9021 28040
rect 9059 28006 9093 28040
rect 9131 28006 9165 28040
rect 9203 28006 9237 28040
rect 9275 28006 9309 28040
rect 9347 28006 9381 28040
rect 9419 28006 9453 28040
rect 9491 28006 9525 28040
rect 9563 28006 9597 28040
rect 9635 28006 9669 28040
rect 9707 28006 9741 28040
rect 9779 28006 9813 28040
rect 9851 28006 9885 28040
rect 9923 28006 9957 28040
rect 9995 28006 10029 28040
rect 10067 28006 10101 28040
rect 10139 28006 10173 28040
rect 10211 28006 10245 28040
rect 10283 28006 10317 28040
rect 10355 28006 10389 28040
rect 10427 28006 10461 28040
rect 10499 28006 10533 28040
rect 10571 28006 10605 28040
rect 10643 28006 10677 28040
rect 10715 28006 10749 28040
rect 10787 28006 10821 28040
rect 10859 28006 10893 28040
rect 10931 28006 10965 28040
rect 11003 28006 11037 28040
rect 11075 28006 11109 28040
rect 11147 28006 11181 28040
rect 11219 28006 11253 28040
rect 11291 28006 11325 28040
rect 11363 28006 11397 28040
rect 11435 28006 11469 28040
rect 11507 28006 11541 28040
rect 11579 28006 11613 28040
rect 11651 28006 11685 28040
rect 11723 28006 11757 28040
rect 11795 28006 11829 28040
rect 11867 28006 11901 28040
rect 11939 28006 11973 28040
rect 12011 28006 12045 28040
rect 12083 28006 12117 28040
rect 12155 28006 12189 28040
rect 12227 28006 12261 28040
rect 12299 28006 12333 28040
rect 12371 28006 12405 28040
rect 12443 28006 12477 28040
rect 12515 28006 12549 28040
rect 12587 28006 12621 28040
rect 12659 28006 12693 28040
rect 12731 28006 12765 28040
rect 12803 28006 12837 28040
rect 12875 28006 12909 28040
rect 12947 28006 12981 28040
rect 13019 28006 13053 28040
rect 13091 28006 13125 28040
rect 13163 28006 13197 28040
rect 13235 28006 13269 28040
rect 13307 28006 13341 28040
rect 13379 28006 13413 28040
rect 13451 28006 13485 28040
rect 13523 28006 13557 28040
rect 13595 28006 13629 28040
rect 13667 28006 13701 28040
rect 13739 28006 13773 28040
rect 13811 28006 13845 28040
rect 13883 28006 13917 28040
rect 112 27943 146 27958
rect 185 27943 219 27958
rect 258 27943 292 27958
rect 331 27943 365 27958
rect 404 27943 438 27958
rect 477 27943 511 27958
rect 550 27943 584 27958
rect 623 27943 657 27958
rect 696 27943 730 27958
rect 769 27943 803 27958
rect 842 27943 876 27958
rect 112 27924 121 27943
rect 121 27924 146 27943
rect 185 27924 190 27943
rect 190 27924 219 27943
rect 258 27924 259 27943
rect 259 27924 292 27943
rect 331 27924 362 27943
rect 362 27924 365 27943
rect 404 27924 431 27943
rect 431 27924 438 27943
rect 477 27924 500 27943
rect 500 27924 511 27943
rect 550 27924 569 27943
rect 569 27924 584 27943
rect 623 27924 638 27943
rect 638 27924 657 27943
rect 696 27924 707 27943
rect 707 27924 730 27943
rect 769 27924 776 27943
rect 776 27924 803 27943
rect 842 27924 845 27943
rect 845 27924 876 27943
rect 915 27924 949 27958
rect 988 27943 1022 27958
rect 1061 27943 1095 27958
rect 988 27924 1018 27943
rect 1018 27924 1022 27943
rect 1061 27924 1087 27943
rect 1087 27924 1095 27943
rect 1134 27924 1156 27958
rect 1156 27924 1168 27958
rect 1207 27924 1241 27958
rect 1280 27924 1314 27958
rect 1353 27924 1387 27958
rect 1426 27924 1460 27958
rect 1499 27924 1533 27958
rect 1571 27924 1605 27958
rect 1643 27924 1677 27958
rect 1715 27924 1749 27958
rect 1787 27924 1821 27958
rect 1859 27924 1893 27958
rect 1931 27924 1965 27958
rect 2003 27924 2037 27958
rect 2075 27924 2109 27958
rect 2147 27924 2181 27958
rect 2219 27924 2253 27958
rect 2291 27924 2325 27958
rect 2363 27924 2397 27958
rect 2435 27924 2469 27958
rect 2507 27924 2541 27958
rect 2579 27924 2613 27958
rect 2651 27924 2685 27958
rect 2723 27924 2757 27958
rect 2795 27924 2829 27958
rect 2867 27924 2901 27958
rect 2939 27924 2973 27958
rect 3011 27924 3045 27958
rect 3083 27924 3117 27958
rect 3155 27924 3189 27958
rect 3227 27924 3261 27958
rect 3299 27924 3333 27958
rect 3371 27924 3405 27958
rect 3443 27924 3477 27958
rect 3515 27924 3549 27958
rect 3587 27924 3621 27958
rect 3659 27924 3693 27958
rect 3731 27924 3765 27958
rect 3803 27924 3837 27958
rect 3875 27924 3909 27958
rect 3947 27924 3981 27958
rect 4019 27924 4053 27958
rect 4091 27924 4125 27958
rect 4163 27924 4197 27958
rect 4235 27924 4269 27958
rect 4307 27924 4341 27958
rect 4379 27924 4413 27958
rect 4451 27924 4485 27958
rect 4523 27924 4557 27958
rect 4595 27924 4629 27958
rect 4667 27924 4701 27958
rect 4739 27924 4773 27958
rect 4811 27924 4845 27958
rect 4883 27924 4917 27958
rect 4955 27924 4989 27958
rect 5027 27924 5061 27958
rect 5099 27924 5133 27958
rect 5171 27924 5205 27958
rect 5243 27924 5277 27958
rect 5315 27924 5349 27958
rect 5387 27924 5421 27958
rect 5459 27924 5493 27958
rect 5531 27924 5565 27958
rect 5603 27924 5637 27958
rect 5675 27924 5709 27958
rect 5747 27924 5781 27958
rect 5819 27924 5853 27958
rect 5891 27924 5925 27958
rect 5963 27924 5997 27958
rect 6035 27924 6069 27958
rect 6107 27924 6141 27958
rect 6179 27924 6213 27958
rect 6251 27924 6285 27958
rect 6323 27924 6357 27958
rect 6395 27924 6429 27958
rect 6467 27924 6501 27958
rect 6539 27924 6573 27958
rect 6611 27924 6645 27958
rect 6683 27924 6717 27958
rect 6755 27924 6789 27958
rect 6827 27924 6861 27958
rect 6899 27924 6933 27958
rect 6971 27924 7005 27958
rect 7043 27924 7077 27958
rect 7115 27924 7149 27958
rect 7187 27924 7221 27958
rect 7259 27924 7293 27958
rect 7331 27924 7365 27958
rect 7403 27924 7437 27958
rect 7475 27924 7509 27958
rect 7547 27924 7581 27958
rect 7619 27924 7653 27958
rect 7691 27924 7725 27958
rect 7763 27924 7797 27958
rect 7835 27924 7869 27958
rect 7907 27924 7941 27958
rect 7979 27924 8013 27958
rect 8051 27924 8085 27958
rect 8123 27924 8157 27958
rect 8195 27924 8229 27958
rect 8267 27924 8301 27958
rect 8339 27924 8373 27958
rect 8411 27924 8445 27958
rect 8483 27924 8517 27958
rect 8555 27924 8589 27958
rect 8627 27924 8661 27958
rect 8699 27924 8733 27958
rect 8771 27924 8805 27958
rect 8843 27924 8877 27958
rect 8915 27924 8949 27958
rect 8987 27924 9021 27958
rect 9059 27924 9093 27958
rect 9131 27924 9165 27958
rect 9203 27924 9237 27958
rect 9275 27924 9309 27958
rect 9347 27924 9381 27958
rect 9419 27924 9453 27958
rect 9491 27924 9525 27958
rect 9563 27924 9597 27958
rect 9635 27924 9669 27958
rect 9707 27924 9741 27958
rect 9779 27924 9813 27958
rect 9851 27924 9885 27958
rect 9923 27924 9957 27958
rect 9995 27924 10029 27958
rect 10067 27924 10101 27958
rect 10139 27924 10173 27958
rect 10211 27924 10245 27958
rect 10283 27924 10317 27958
rect 10355 27924 10389 27958
rect 10427 27924 10461 27958
rect 10499 27924 10533 27958
rect 10571 27924 10605 27958
rect 10643 27924 10677 27958
rect 10715 27924 10749 27958
rect 10787 27924 10821 27958
rect 10859 27924 10893 27958
rect 10931 27924 10965 27958
rect 11003 27924 11037 27958
rect 11075 27924 11109 27958
rect 11147 27924 11181 27958
rect 11219 27924 11253 27958
rect 11291 27924 11325 27958
rect 11363 27924 11397 27958
rect 11435 27924 11469 27958
rect 11507 27924 11541 27958
rect 11579 27924 11613 27958
rect 11651 27924 11685 27958
rect 11723 27924 11757 27958
rect 11795 27924 11829 27958
rect 11867 27924 11901 27958
rect 11939 27924 11973 27958
rect 12011 27924 12045 27958
rect 12083 27924 12117 27958
rect 12155 27924 12189 27958
rect 12227 27924 12261 27958
rect 12299 27924 12333 27958
rect 12371 27924 12405 27958
rect 12443 27924 12477 27958
rect 12515 27924 12549 27958
rect 12587 27924 12621 27958
rect 12659 27924 12693 27958
rect 12731 27924 12765 27958
rect 12803 27924 12837 27958
rect 12875 27924 12909 27958
rect 12947 27924 12981 27958
rect 13019 27924 13053 27958
rect 13091 27924 13125 27958
rect 13163 27924 13197 27958
rect 13235 27924 13269 27958
rect 13307 27924 13341 27958
rect 13379 27924 13413 27958
rect 13451 27924 13485 27958
rect 13523 27924 13557 27958
rect 13595 27924 13629 27958
rect 13667 27924 13701 27958
rect 13739 27924 13773 27958
rect 13811 27924 13845 27958
rect 13883 27924 13917 27958
rect 112 27875 146 27876
rect 185 27875 219 27876
rect 258 27875 292 27876
rect 331 27875 365 27876
rect 404 27875 438 27876
rect 477 27875 511 27876
rect 550 27875 584 27876
rect 623 27875 657 27876
rect 696 27875 730 27876
rect 769 27875 803 27876
rect 842 27875 876 27876
rect 112 27842 121 27875
rect 121 27842 146 27875
rect 185 27842 190 27875
rect 190 27842 219 27875
rect 258 27842 259 27875
rect 259 27842 292 27875
rect 331 27842 362 27875
rect 362 27842 365 27875
rect 404 27842 431 27875
rect 431 27842 438 27875
rect 477 27842 500 27875
rect 500 27842 511 27875
rect 550 27842 569 27875
rect 569 27842 584 27875
rect 623 27842 638 27875
rect 638 27842 657 27875
rect 696 27842 707 27875
rect 707 27842 730 27875
rect 769 27842 776 27875
rect 776 27842 803 27875
rect 842 27842 845 27875
rect 845 27842 876 27875
rect 915 27842 949 27876
rect 988 27875 1022 27876
rect 1061 27875 1095 27876
rect 988 27842 1018 27875
rect 1018 27842 1022 27875
rect 1061 27842 1087 27875
rect 1087 27842 1095 27875
rect 1134 27842 1156 27876
rect 1156 27842 1168 27876
rect 1207 27842 1241 27876
rect 1280 27842 1314 27876
rect 1353 27842 1387 27876
rect 1426 27842 1460 27876
rect 1499 27842 1533 27876
rect 1571 27842 1605 27876
rect 1643 27842 1677 27876
rect 1715 27842 1749 27876
rect 1787 27842 1821 27876
rect 1859 27842 1893 27876
rect 1931 27842 1965 27876
rect 2003 27842 2037 27876
rect 2075 27842 2109 27876
rect 2147 27842 2181 27876
rect 2219 27842 2253 27876
rect 2291 27842 2325 27876
rect 2363 27842 2397 27876
rect 2435 27842 2469 27876
rect 2507 27842 2541 27876
rect 2579 27842 2613 27876
rect 2651 27842 2685 27876
rect 2723 27842 2757 27876
rect 2795 27842 2829 27876
rect 2867 27842 2901 27876
rect 2939 27842 2973 27876
rect 3011 27842 3045 27876
rect 3083 27842 3117 27876
rect 3155 27842 3189 27876
rect 3227 27842 3261 27876
rect 3299 27842 3333 27876
rect 3371 27842 3405 27876
rect 3443 27842 3477 27876
rect 3515 27842 3549 27876
rect 3587 27842 3621 27876
rect 3659 27842 3693 27876
rect 3731 27842 3765 27876
rect 3803 27842 3837 27876
rect 3875 27842 3909 27876
rect 3947 27842 3981 27876
rect 4019 27842 4053 27876
rect 4091 27842 4125 27876
rect 4163 27842 4197 27876
rect 4235 27842 4269 27876
rect 4307 27842 4341 27876
rect 4379 27842 4413 27876
rect 4451 27842 4485 27876
rect 4523 27842 4557 27876
rect 4595 27842 4629 27876
rect 4667 27842 4701 27876
rect 4739 27842 4773 27876
rect 4811 27842 4845 27876
rect 4883 27842 4917 27876
rect 4955 27842 4989 27876
rect 5027 27842 5061 27876
rect 5099 27842 5133 27876
rect 5171 27842 5205 27876
rect 5243 27842 5277 27876
rect 5315 27842 5349 27876
rect 5387 27842 5421 27876
rect 5459 27842 5493 27876
rect 5531 27842 5565 27876
rect 5603 27842 5637 27876
rect 5675 27842 5709 27876
rect 5747 27842 5781 27876
rect 5819 27842 5853 27876
rect 5891 27842 5925 27876
rect 5963 27842 5997 27876
rect 6035 27842 6069 27876
rect 6107 27842 6141 27876
rect 6179 27842 6213 27876
rect 6251 27842 6285 27876
rect 6323 27842 6357 27876
rect 6395 27842 6429 27876
rect 6467 27842 6501 27876
rect 6539 27842 6573 27876
rect 6611 27842 6645 27876
rect 6683 27842 6717 27876
rect 6755 27842 6789 27876
rect 6827 27842 6861 27876
rect 6899 27842 6933 27876
rect 6971 27842 7005 27876
rect 7043 27842 7077 27876
rect 7115 27842 7149 27876
rect 7187 27842 7221 27876
rect 7259 27842 7293 27876
rect 7331 27842 7365 27876
rect 7403 27842 7437 27876
rect 7475 27842 7509 27876
rect 7547 27842 7581 27876
rect 7619 27842 7653 27876
rect 7691 27842 7725 27876
rect 7763 27842 7797 27876
rect 7835 27842 7869 27876
rect 7907 27842 7941 27876
rect 7979 27842 8013 27876
rect 8051 27842 8085 27876
rect 8123 27842 8157 27876
rect 8195 27842 8229 27876
rect 8267 27842 8301 27876
rect 8339 27842 8373 27876
rect 8411 27842 8445 27876
rect 8483 27842 8517 27876
rect 8555 27842 8589 27876
rect 8627 27842 8661 27876
rect 8699 27842 8733 27876
rect 8771 27842 8805 27876
rect 8843 27842 8877 27876
rect 8915 27842 8949 27876
rect 8987 27842 9021 27876
rect 9059 27842 9093 27876
rect 9131 27842 9165 27876
rect 9203 27842 9237 27876
rect 9275 27842 9309 27876
rect 9347 27842 9381 27876
rect 9419 27842 9453 27876
rect 9491 27842 9525 27876
rect 9563 27842 9597 27876
rect 9635 27842 9669 27876
rect 9707 27842 9741 27876
rect 9779 27842 9813 27876
rect 9851 27842 9885 27876
rect 9923 27842 9957 27876
rect 9995 27842 10029 27876
rect 10067 27842 10101 27876
rect 10139 27842 10173 27876
rect 10211 27842 10245 27876
rect 10283 27842 10317 27876
rect 10355 27842 10389 27876
rect 10427 27842 10461 27876
rect 10499 27842 10533 27876
rect 10571 27842 10605 27876
rect 10643 27842 10677 27876
rect 10715 27842 10749 27876
rect 10787 27842 10821 27876
rect 10859 27842 10893 27876
rect 10931 27842 10965 27876
rect 11003 27842 11037 27876
rect 11075 27842 11109 27876
rect 11147 27842 11181 27876
rect 11219 27842 11253 27876
rect 11291 27842 11325 27876
rect 11363 27842 11397 27876
rect 11435 27842 11469 27876
rect 11507 27842 11541 27876
rect 11579 27842 11613 27876
rect 11651 27842 11685 27876
rect 11723 27842 11757 27876
rect 11795 27842 11829 27876
rect 11867 27842 11901 27876
rect 11939 27842 11973 27876
rect 12011 27842 12045 27876
rect 12083 27842 12117 27876
rect 12155 27842 12189 27876
rect 12227 27842 12261 27876
rect 12299 27842 12333 27876
rect 12371 27842 12405 27876
rect 12443 27842 12477 27876
rect 12515 27842 12549 27876
rect 12587 27842 12621 27876
rect 12659 27842 12693 27876
rect 12731 27842 12765 27876
rect 12803 27842 12837 27876
rect 12875 27842 12909 27876
rect 12947 27842 12981 27876
rect 13019 27842 13053 27876
rect 13091 27842 13125 27876
rect 13163 27842 13197 27876
rect 13235 27842 13269 27876
rect 13307 27842 13341 27876
rect 13379 27842 13413 27876
rect 13451 27842 13485 27876
rect 13523 27842 13557 27876
rect 13595 27842 13629 27876
rect 13667 27842 13701 27876
rect 13739 27842 13773 27876
rect 13811 27842 13845 27876
rect 13883 27842 13917 27876
rect 112 27773 121 27794
rect 121 27773 146 27794
rect 185 27773 190 27794
rect 190 27773 219 27794
rect 258 27773 259 27794
rect 259 27773 292 27794
rect 331 27773 362 27794
rect 362 27773 365 27794
rect 404 27773 431 27794
rect 431 27773 438 27794
rect 477 27773 500 27794
rect 500 27773 511 27794
rect 550 27773 569 27794
rect 569 27773 584 27794
rect 623 27773 638 27794
rect 638 27773 657 27794
rect 696 27773 707 27794
rect 707 27773 730 27794
rect 769 27773 776 27794
rect 776 27773 803 27794
rect 842 27773 845 27794
rect 845 27773 876 27794
rect 112 27760 146 27773
rect 185 27760 219 27773
rect 258 27760 292 27773
rect 331 27760 365 27773
rect 404 27760 438 27773
rect 477 27760 511 27773
rect 550 27760 584 27773
rect 623 27760 657 27773
rect 696 27760 730 27773
rect 769 27760 803 27773
rect 842 27760 876 27773
rect 915 27760 949 27794
rect 988 27773 1018 27794
rect 1018 27773 1022 27794
rect 1061 27773 1087 27794
rect 1087 27773 1095 27794
rect 988 27760 1022 27773
rect 1061 27760 1095 27773
rect 1134 27760 1156 27794
rect 1156 27760 1168 27794
rect 1207 27760 1241 27794
rect 1280 27760 1314 27794
rect 1353 27760 1387 27794
rect 1426 27760 1460 27794
rect 1499 27760 1533 27794
rect 1571 27760 1605 27794
rect 1643 27760 1677 27794
rect 1715 27760 1749 27794
rect 1787 27760 1821 27794
rect 1859 27760 1893 27794
rect 1931 27760 1965 27794
rect 2003 27760 2037 27794
rect 2075 27760 2109 27794
rect 2147 27760 2181 27794
rect 2219 27760 2253 27794
rect 2291 27760 2325 27794
rect 2363 27760 2397 27794
rect 2435 27760 2469 27794
rect 2507 27760 2541 27794
rect 2579 27760 2613 27794
rect 2651 27760 2685 27794
rect 2723 27760 2757 27794
rect 2795 27760 2829 27794
rect 2867 27760 2901 27794
rect 2939 27760 2973 27794
rect 3011 27760 3045 27794
rect 3083 27760 3117 27794
rect 3155 27760 3189 27794
rect 3227 27760 3261 27794
rect 3299 27760 3333 27794
rect 3371 27760 3405 27794
rect 3443 27760 3477 27794
rect 3515 27760 3549 27794
rect 3587 27760 3621 27794
rect 3659 27760 3693 27794
rect 3731 27760 3765 27794
rect 3803 27760 3837 27794
rect 3875 27760 3909 27794
rect 3947 27760 3981 27794
rect 4019 27760 4053 27794
rect 4091 27760 4125 27794
rect 4163 27760 4197 27794
rect 4235 27760 4269 27794
rect 4307 27760 4341 27794
rect 4379 27760 4413 27794
rect 4451 27760 4485 27794
rect 4523 27760 4557 27794
rect 4595 27760 4629 27794
rect 4667 27760 4701 27794
rect 4739 27760 4773 27794
rect 4811 27760 4845 27794
rect 4883 27760 4917 27794
rect 4955 27760 4989 27794
rect 5027 27760 5061 27794
rect 5099 27760 5133 27794
rect 5171 27760 5205 27794
rect 5243 27760 5277 27794
rect 5315 27760 5349 27794
rect 5387 27760 5421 27794
rect 5459 27760 5493 27794
rect 5531 27760 5565 27794
rect 5603 27760 5637 27794
rect 5675 27760 5709 27794
rect 5747 27760 5781 27794
rect 5819 27760 5853 27794
rect 5891 27760 5925 27794
rect 5963 27760 5997 27794
rect 6035 27760 6069 27794
rect 6107 27760 6141 27794
rect 6179 27760 6213 27794
rect 6251 27760 6285 27794
rect 6323 27760 6357 27794
rect 6395 27760 6429 27794
rect 6467 27760 6501 27794
rect 6539 27760 6573 27794
rect 6611 27760 6645 27794
rect 6683 27760 6717 27794
rect 6755 27760 6789 27794
rect 6827 27760 6861 27794
rect 6899 27760 6933 27794
rect 6971 27760 7005 27794
rect 7043 27760 7077 27794
rect 7115 27760 7149 27794
rect 7187 27760 7221 27794
rect 7259 27760 7293 27794
rect 7331 27760 7365 27794
rect 7403 27760 7437 27794
rect 7475 27760 7509 27794
rect 7547 27760 7581 27794
rect 7619 27760 7653 27794
rect 7691 27760 7725 27794
rect 7763 27760 7797 27794
rect 7835 27760 7869 27794
rect 7907 27760 7941 27794
rect 7979 27760 8013 27794
rect 8051 27760 8085 27794
rect 8123 27760 8157 27794
rect 8195 27760 8229 27794
rect 8267 27760 8301 27794
rect 8339 27760 8373 27794
rect 8411 27760 8445 27794
rect 8483 27760 8517 27794
rect 8555 27760 8589 27794
rect 8627 27760 8661 27794
rect 8699 27760 8733 27794
rect 8771 27760 8805 27794
rect 8843 27760 8877 27794
rect 8915 27760 8949 27794
rect 8987 27760 9021 27794
rect 9059 27760 9093 27794
rect 9131 27760 9165 27794
rect 9203 27760 9237 27794
rect 9275 27760 9309 27794
rect 9347 27760 9381 27794
rect 9419 27760 9453 27794
rect 9491 27760 9525 27794
rect 9563 27760 9597 27794
rect 9635 27760 9669 27794
rect 9707 27760 9741 27794
rect 9779 27760 9813 27794
rect 9851 27760 9885 27794
rect 9923 27760 9957 27794
rect 9995 27760 10029 27794
rect 10067 27760 10101 27794
rect 10139 27760 10173 27794
rect 10211 27760 10245 27794
rect 10283 27760 10317 27794
rect 10355 27760 10389 27794
rect 10427 27760 10461 27794
rect 10499 27760 10533 27794
rect 10571 27760 10605 27794
rect 10643 27760 10677 27794
rect 10715 27760 10749 27794
rect 10787 27760 10821 27794
rect 10859 27760 10893 27794
rect 10931 27760 10965 27794
rect 11003 27760 11037 27794
rect 11075 27760 11109 27794
rect 11147 27760 11181 27794
rect 11219 27760 11253 27794
rect 11291 27760 11325 27794
rect 11363 27760 11397 27794
rect 11435 27760 11469 27794
rect 11507 27760 11541 27794
rect 11579 27760 11613 27794
rect 11651 27760 11685 27794
rect 11723 27760 11757 27794
rect 11795 27760 11829 27794
rect 11867 27760 11901 27794
rect 11939 27760 11973 27794
rect 12011 27760 12045 27794
rect 12083 27760 12117 27794
rect 12155 27760 12189 27794
rect 12227 27760 12261 27794
rect 12299 27760 12333 27794
rect 12371 27760 12405 27794
rect 12443 27760 12477 27794
rect 12515 27760 12549 27794
rect 12587 27760 12621 27794
rect 12659 27760 12693 27794
rect 12731 27760 12765 27794
rect 12803 27760 12837 27794
rect 12875 27760 12909 27794
rect 12947 27760 12981 27794
rect 13019 27760 13053 27794
rect 13091 27760 13125 27794
rect 13163 27760 13197 27794
rect 13235 27760 13269 27794
rect 13307 27760 13341 27794
rect 13379 27760 13413 27794
rect 13451 27760 13485 27794
rect 13523 27760 13557 27794
rect 13595 27760 13629 27794
rect 13667 27760 13701 27794
rect 13739 27760 13773 27794
rect 13811 27760 13845 27794
rect 13883 27760 13917 27794
rect 112 27705 121 27712
rect 121 27705 146 27712
rect 185 27705 190 27712
rect 190 27705 219 27712
rect 258 27705 259 27712
rect 259 27705 292 27712
rect 331 27705 362 27712
rect 362 27705 365 27712
rect 404 27705 431 27712
rect 431 27705 438 27712
rect 477 27705 500 27712
rect 500 27705 511 27712
rect 550 27705 569 27712
rect 569 27705 584 27712
rect 623 27705 638 27712
rect 638 27705 657 27712
rect 696 27705 707 27712
rect 707 27705 730 27712
rect 769 27705 776 27712
rect 776 27705 803 27712
rect 842 27705 845 27712
rect 845 27705 876 27712
rect 112 27678 146 27705
rect 185 27678 219 27705
rect 258 27678 292 27705
rect 331 27678 365 27705
rect 404 27678 438 27705
rect 477 27678 511 27705
rect 550 27678 584 27705
rect 623 27678 657 27705
rect 696 27678 730 27705
rect 769 27678 803 27705
rect 842 27678 876 27705
rect 915 27678 949 27712
rect 988 27705 1018 27712
rect 1018 27705 1022 27712
rect 1061 27705 1087 27712
rect 1087 27705 1095 27712
rect 988 27678 1022 27705
rect 1061 27678 1095 27705
rect 1134 27678 1156 27712
rect 1156 27678 1168 27712
rect 1207 27678 1241 27712
rect 1280 27678 1314 27712
rect 1353 27678 1387 27712
rect 1426 27678 1460 27712
rect 1499 27678 1533 27712
rect 1571 27678 1605 27712
rect 1643 27678 1677 27712
rect 1715 27678 1749 27712
rect 1787 27678 1821 27712
rect 1859 27678 1893 27712
rect 1931 27678 1965 27712
rect 2003 27678 2037 27712
rect 2075 27678 2109 27712
rect 2147 27678 2181 27712
rect 2219 27678 2253 27712
rect 2291 27678 2325 27712
rect 2363 27678 2397 27712
rect 2435 27678 2469 27712
rect 2507 27678 2541 27712
rect 2579 27678 2613 27712
rect 2651 27678 2685 27712
rect 2723 27678 2757 27712
rect 2795 27678 2829 27712
rect 2867 27678 2901 27712
rect 2939 27678 2973 27712
rect 3011 27678 3045 27712
rect 3083 27678 3117 27712
rect 3155 27678 3189 27712
rect 3227 27678 3261 27712
rect 3299 27678 3333 27712
rect 3371 27678 3405 27712
rect 3443 27678 3477 27712
rect 3515 27678 3549 27712
rect 3587 27678 3621 27712
rect 3659 27678 3693 27712
rect 3731 27678 3765 27712
rect 3803 27678 3837 27712
rect 3875 27678 3909 27712
rect 3947 27678 3981 27712
rect 4019 27678 4053 27712
rect 4091 27678 4125 27712
rect 4163 27678 4197 27712
rect 4235 27678 4269 27712
rect 4307 27678 4341 27712
rect 4379 27678 4413 27712
rect 4451 27678 4485 27712
rect 4523 27678 4557 27712
rect 4595 27678 4629 27712
rect 4667 27678 4701 27712
rect 4739 27678 4773 27712
rect 4811 27678 4845 27712
rect 4883 27678 4917 27712
rect 4955 27678 4989 27712
rect 5027 27678 5061 27712
rect 5099 27678 5133 27712
rect 5171 27678 5205 27712
rect 5243 27678 5277 27712
rect 5315 27678 5349 27712
rect 5387 27678 5421 27712
rect 5459 27678 5493 27712
rect 5531 27678 5565 27712
rect 5603 27678 5637 27712
rect 5675 27678 5709 27712
rect 5747 27678 5781 27712
rect 5819 27678 5853 27712
rect 5891 27678 5925 27712
rect 5963 27678 5997 27712
rect 6035 27678 6069 27712
rect 6107 27678 6141 27712
rect 6179 27678 6213 27712
rect 6251 27678 6285 27712
rect 6323 27678 6357 27712
rect 6395 27678 6429 27712
rect 6467 27678 6501 27712
rect 6539 27678 6573 27712
rect 6611 27678 6645 27712
rect 6683 27678 6717 27712
rect 6755 27678 6789 27712
rect 6827 27678 6861 27712
rect 6899 27678 6933 27712
rect 6971 27678 7005 27712
rect 7043 27678 7077 27712
rect 7115 27678 7149 27712
rect 7187 27678 7221 27712
rect 7259 27678 7293 27712
rect 7331 27678 7365 27712
rect 7403 27678 7437 27712
rect 7475 27678 7509 27712
rect 7547 27678 7581 27712
rect 7619 27678 7653 27712
rect 7691 27678 7725 27712
rect 7763 27678 7797 27712
rect 7835 27678 7869 27712
rect 7907 27678 7941 27712
rect 7979 27678 8013 27712
rect 8051 27678 8085 27712
rect 8123 27678 8157 27712
rect 8195 27678 8229 27712
rect 8267 27678 8301 27712
rect 8339 27678 8373 27712
rect 8411 27678 8445 27712
rect 8483 27678 8517 27712
rect 8555 27678 8589 27712
rect 8627 27678 8661 27712
rect 8699 27678 8733 27712
rect 8771 27678 8805 27712
rect 8843 27678 8877 27712
rect 8915 27678 8949 27712
rect 8987 27678 9021 27712
rect 9059 27678 9093 27712
rect 9131 27678 9165 27712
rect 9203 27678 9237 27712
rect 9275 27678 9309 27712
rect 9347 27678 9381 27712
rect 9419 27678 9453 27712
rect 9491 27678 9525 27712
rect 9563 27678 9597 27712
rect 9635 27678 9669 27712
rect 9707 27678 9741 27712
rect 9779 27678 9813 27712
rect 9851 27678 9885 27712
rect 9923 27678 9957 27712
rect 9995 27678 10029 27712
rect 10067 27678 10101 27712
rect 10139 27678 10173 27712
rect 10211 27678 10245 27712
rect 10283 27678 10317 27712
rect 10355 27678 10389 27712
rect 10427 27678 10461 27712
rect 10499 27678 10533 27712
rect 10571 27678 10605 27712
rect 10643 27678 10677 27712
rect 10715 27678 10749 27712
rect 10787 27678 10821 27712
rect 10859 27678 10893 27712
rect 10931 27678 10965 27712
rect 11003 27678 11037 27712
rect 11075 27678 11109 27712
rect 11147 27678 11181 27712
rect 11219 27678 11253 27712
rect 11291 27678 11325 27712
rect 11363 27678 11397 27712
rect 11435 27678 11469 27712
rect 11507 27678 11541 27712
rect 11579 27678 11613 27712
rect 11651 27678 11685 27712
rect 11723 27678 11757 27712
rect 11795 27678 11829 27712
rect 11867 27678 11901 27712
rect 11939 27678 11973 27712
rect 12011 27678 12045 27712
rect 12083 27678 12117 27712
rect 12155 27678 12189 27712
rect 12227 27678 12261 27712
rect 12299 27678 12333 27712
rect 12371 27678 12405 27712
rect 12443 27678 12477 27712
rect 12515 27678 12549 27712
rect 12587 27678 12621 27712
rect 12659 27678 12693 27712
rect 12731 27678 12765 27712
rect 12803 27678 12837 27712
rect 12875 27678 12909 27712
rect 12947 27678 12981 27712
rect 13019 27678 13053 27712
rect 13091 27678 13125 27712
rect 13163 27678 13197 27712
rect 13235 27678 13269 27712
rect 13307 27678 13341 27712
rect 13379 27678 13413 27712
rect 13451 27678 13485 27712
rect 13523 27678 13557 27712
rect 13595 27678 13629 27712
rect 13667 27678 13701 27712
rect 13739 27678 13773 27712
rect 13811 27678 13845 27712
rect 13883 27678 13917 27712
rect 163 27342 186 27355
rect 186 27342 197 27355
rect 237 27342 255 27355
rect 255 27342 271 27355
rect 311 27342 324 27355
rect 324 27342 345 27355
rect 385 27342 393 27355
rect 393 27342 419 27355
rect 459 27342 462 27355
rect 462 27342 493 27355
rect 533 27342 566 27355
rect 566 27342 567 27355
rect 606 27342 635 27355
rect 635 27342 640 27355
rect 679 27342 704 27355
rect 704 27342 713 27355
rect 752 27342 773 27355
rect 773 27342 786 27355
rect 827 27342 842 27362
rect 842 27342 861 27362
rect 899 27342 911 27362
rect 911 27342 933 27362
rect 971 27342 980 27362
rect 980 27342 1005 27362
rect 1043 27342 1049 27362
rect 1049 27342 1077 27362
rect 1115 27342 1118 27362
rect 1118 27342 1149 27362
rect 1187 27342 1221 27362
rect 1259 27342 1290 27362
rect 1290 27342 1293 27362
rect 1331 27342 1359 27362
rect 1359 27342 1365 27362
rect 1403 27342 1428 27362
rect 1428 27342 1437 27362
rect 1475 27342 1497 27362
rect 1497 27342 1509 27362
rect 1547 27342 1566 27362
rect 1566 27342 1581 27362
rect 1619 27342 1635 27362
rect 1635 27342 1653 27362
rect 1691 27342 1704 27362
rect 1704 27342 1725 27362
rect 1764 27342 1773 27362
rect 1773 27342 1798 27362
rect 1837 27342 1842 27362
rect 1842 27342 1871 27362
rect 1910 27342 1911 27362
rect 1911 27342 1944 27362
rect 1983 27342 2014 27362
rect 2014 27342 2017 27362
rect 2056 27342 2082 27362
rect 2082 27342 2090 27362
rect 2142 27342 2150 27355
rect 2150 27342 2176 27355
rect 2221 27342 2252 27355
rect 2252 27342 2255 27355
rect 2300 27342 2320 27355
rect 2320 27342 2334 27355
rect 2379 27342 2388 27355
rect 2388 27342 2413 27355
rect 2458 27342 2490 27355
rect 2490 27342 2492 27355
rect 2536 27342 2558 27355
rect 2558 27342 2570 27355
rect 2614 27342 2626 27355
rect 2626 27342 2648 27355
rect 2692 27342 2694 27355
rect 2694 27342 2726 27355
rect 2770 27342 2796 27355
rect 2796 27342 2804 27355
rect 163 27321 197 27342
rect 237 27321 271 27342
rect 311 27321 345 27342
rect 385 27321 419 27342
rect 459 27321 493 27342
rect 533 27321 567 27342
rect 606 27321 640 27342
rect 679 27321 713 27342
rect 752 27321 786 27342
rect 827 27328 861 27342
rect 899 27328 933 27342
rect 971 27328 1005 27342
rect 1043 27328 1077 27342
rect 1115 27328 1149 27342
rect 1187 27328 1221 27342
rect 1259 27328 1293 27342
rect 1331 27328 1365 27342
rect 1403 27328 1437 27342
rect 1475 27328 1509 27342
rect 1547 27328 1581 27342
rect 1619 27328 1653 27342
rect 1691 27328 1725 27342
rect 1764 27328 1798 27342
rect 1837 27328 1871 27342
rect 1910 27328 1944 27342
rect 1983 27328 2017 27342
rect 2056 27328 2090 27342
rect 2142 27321 2176 27342
rect 2221 27321 2255 27342
rect 2300 27321 2334 27342
rect 2379 27321 2413 27342
rect 2458 27321 2492 27342
rect 2536 27321 2570 27342
rect 2614 27321 2648 27342
rect 2692 27321 2726 27342
rect 2770 27321 2804 27342
rect 2848 27338 2882 27355
rect 2926 27338 2950 27355
rect 2950 27338 2960 27355
rect 3392 27338 3426 27362
rect 3465 27338 3494 27362
rect 3494 27338 3499 27362
rect 3538 27338 3562 27362
rect 3562 27338 3572 27362
rect 3611 27338 3630 27362
rect 3630 27338 3645 27362
rect 3684 27338 3698 27362
rect 3698 27338 3718 27362
rect 3757 27338 3766 27362
rect 3766 27338 3791 27362
rect 3830 27338 3834 27362
rect 3834 27338 3864 27362
rect 3903 27338 3936 27362
rect 3936 27338 3937 27362
rect 3976 27338 4004 27362
rect 4004 27338 4010 27362
rect 4049 27338 4072 27362
rect 4072 27338 4083 27362
rect 4122 27338 4140 27362
rect 4140 27338 4156 27362
rect 4194 27338 4208 27362
rect 4208 27338 4228 27362
rect 4266 27338 4276 27362
rect 4276 27338 4300 27362
rect 4338 27338 4344 27362
rect 4344 27338 4372 27362
rect 4410 27338 4412 27362
rect 4412 27338 4444 27362
rect 4482 27338 4514 27362
rect 4514 27338 4516 27362
rect 4554 27338 4582 27362
rect 4582 27338 4588 27362
rect 4626 27338 4650 27362
rect 4650 27338 4660 27362
rect 4698 27338 4718 27362
rect 4718 27338 4732 27362
rect 4770 27338 4786 27362
rect 4786 27338 4804 27362
rect 4842 27338 4854 27362
rect 4854 27338 4876 27362
rect 4914 27338 4922 27362
rect 4922 27338 4948 27362
rect 4986 27338 4990 27362
rect 4990 27338 5020 27362
rect 2848 27321 2882 27338
rect 2926 27321 2960 27338
rect 3392 27328 3426 27338
rect 3465 27328 3499 27338
rect 3538 27328 3572 27338
rect 3611 27328 3645 27338
rect 3684 27328 3718 27338
rect 3757 27328 3791 27338
rect 3830 27328 3864 27338
rect 3903 27328 3937 27338
rect 3976 27328 4010 27338
rect 4049 27328 4083 27338
rect 4122 27328 4156 27338
rect 4194 27328 4228 27338
rect 4266 27328 4300 27338
rect 4338 27328 4372 27338
rect 4410 27328 4444 27338
rect 4482 27328 4516 27338
rect 4554 27328 4588 27338
rect 4626 27328 4660 27338
rect 4698 27328 4732 27338
rect 4770 27328 4804 27338
rect 4842 27328 4876 27338
rect 4914 27328 4948 27338
rect 4986 27328 5020 27338
rect 5058 27328 5092 27362
rect 5130 27338 5160 27362
rect 5160 27338 5164 27362
rect 5202 27338 5228 27362
rect 5228 27338 5236 27362
rect 5274 27338 5296 27362
rect 5296 27338 5308 27362
rect 5346 27338 5364 27362
rect 5364 27338 5380 27362
rect 5418 27338 5432 27362
rect 5432 27338 5452 27362
rect 5490 27338 5500 27362
rect 5500 27338 5524 27362
rect 5562 27338 5568 27362
rect 5568 27338 5596 27362
rect 5634 27338 5636 27362
rect 5636 27338 5668 27362
rect 5706 27338 5738 27362
rect 5738 27338 5740 27362
rect 5778 27338 5806 27362
rect 5806 27338 5812 27362
rect 5850 27338 5874 27362
rect 5874 27338 5884 27362
rect 5922 27338 5942 27362
rect 5942 27338 5956 27362
rect 5994 27338 6010 27362
rect 6010 27338 6028 27362
rect 6066 27338 6078 27362
rect 6078 27338 6100 27362
rect 6138 27338 6146 27362
rect 6146 27338 6172 27362
rect 6210 27338 6214 27362
rect 6214 27338 6244 27362
rect 5130 27328 5164 27338
rect 5202 27328 5236 27338
rect 5274 27328 5308 27338
rect 5346 27328 5380 27338
rect 5418 27328 5452 27338
rect 5490 27328 5524 27338
rect 5562 27328 5596 27338
rect 5634 27328 5668 27338
rect 5706 27328 5740 27338
rect 5778 27328 5812 27338
rect 5850 27328 5884 27338
rect 5922 27328 5956 27338
rect 5994 27328 6028 27338
rect 6066 27328 6100 27338
rect 6138 27328 6172 27338
rect 6210 27328 6244 27338
rect 6282 27328 6316 27362
rect 6354 27338 6384 27362
rect 6384 27338 6388 27362
rect 6426 27338 6452 27362
rect 6452 27338 6460 27362
rect 6498 27338 6520 27362
rect 6520 27338 6532 27362
rect 6570 27338 6588 27362
rect 6588 27338 6604 27362
rect 6642 27338 6656 27362
rect 6656 27338 6676 27362
rect 6714 27338 6724 27362
rect 6724 27338 6748 27362
rect 6786 27338 6792 27362
rect 6792 27338 6820 27362
rect 6858 27338 6860 27362
rect 6860 27338 6892 27362
rect 6930 27338 6962 27362
rect 6962 27338 6964 27362
rect 7002 27338 7030 27362
rect 7030 27338 7036 27362
rect 7074 27338 7098 27362
rect 7098 27338 7108 27362
rect 7146 27338 7166 27362
rect 7166 27338 7180 27362
rect 7218 27338 7234 27362
rect 7234 27338 7252 27362
rect 7290 27338 7302 27362
rect 7302 27338 7324 27362
rect 7362 27338 7370 27362
rect 7370 27338 7396 27362
rect 7434 27338 7438 27362
rect 7438 27338 7468 27362
rect 6354 27328 6388 27338
rect 6426 27328 6460 27338
rect 6498 27328 6532 27338
rect 6570 27328 6604 27338
rect 6642 27328 6676 27338
rect 6714 27328 6748 27338
rect 6786 27328 6820 27338
rect 6858 27328 6892 27338
rect 6930 27328 6964 27338
rect 7002 27328 7036 27338
rect 7074 27328 7108 27338
rect 7146 27328 7180 27338
rect 7218 27328 7252 27338
rect 7290 27328 7324 27338
rect 7362 27328 7396 27338
rect 7434 27328 7468 27338
rect 7506 27328 7540 27362
rect 7578 27338 7608 27362
rect 7608 27338 7612 27362
rect 7650 27338 7676 27362
rect 7676 27338 7684 27362
rect 7722 27338 7744 27362
rect 7744 27338 7756 27362
rect 7794 27338 7812 27362
rect 7812 27338 7828 27362
rect 7866 27338 7880 27362
rect 7880 27338 7900 27362
rect 7938 27338 7948 27362
rect 7948 27338 7972 27362
rect 8010 27338 8016 27362
rect 8016 27338 8044 27362
rect 8082 27338 8084 27362
rect 8084 27338 8116 27362
rect 8154 27338 8186 27362
rect 8186 27338 8188 27362
rect 8226 27338 8254 27362
rect 8254 27338 8260 27362
rect 8298 27338 8322 27362
rect 8322 27338 8332 27362
rect 8370 27338 8390 27362
rect 8390 27338 8404 27362
rect 8442 27338 8458 27362
rect 8458 27338 8476 27362
rect 8514 27338 8526 27362
rect 8526 27338 8548 27362
rect 8586 27338 8594 27362
rect 8594 27338 8620 27362
rect 8658 27338 8662 27362
rect 8662 27338 8692 27362
rect 7578 27328 7612 27338
rect 7650 27328 7684 27338
rect 7722 27328 7756 27338
rect 7794 27328 7828 27338
rect 7866 27328 7900 27338
rect 7938 27328 7972 27338
rect 8010 27328 8044 27338
rect 8082 27328 8116 27338
rect 8154 27328 8188 27338
rect 8226 27328 8260 27338
rect 8298 27328 8332 27338
rect 8370 27328 8404 27338
rect 8442 27328 8476 27338
rect 8514 27328 8548 27338
rect 8586 27328 8620 27338
rect 8658 27328 8692 27338
rect 8730 27328 8764 27362
rect 8802 27338 8832 27362
rect 8832 27338 8836 27362
rect 8874 27338 8900 27362
rect 8900 27338 8908 27362
rect 8946 27338 8968 27362
rect 8968 27338 8980 27362
rect 9018 27338 9036 27362
rect 9036 27338 9052 27362
rect 9090 27338 9104 27362
rect 9104 27338 9124 27362
rect 9162 27338 9172 27362
rect 9172 27338 9196 27362
rect 9234 27338 9240 27362
rect 9240 27338 9268 27362
rect 9306 27338 9308 27362
rect 9308 27338 9340 27362
rect 9378 27338 9410 27362
rect 9410 27338 9412 27362
rect 9450 27338 9478 27362
rect 9478 27338 9484 27362
rect 9522 27338 9546 27362
rect 9546 27338 9556 27362
rect 9594 27338 9614 27362
rect 9614 27338 9628 27362
rect 9666 27338 9682 27362
rect 9682 27338 9700 27362
rect 9738 27338 9750 27362
rect 9750 27338 9772 27362
rect 9810 27338 9818 27362
rect 9818 27338 9844 27362
rect 9882 27338 9886 27362
rect 9886 27338 9916 27362
rect 8802 27328 8836 27338
rect 8874 27328 8908 27338
rect 8946 27328 8980 27338
rect 9018 27328 9052 27338
rect 9090 27328 9124 27338
rect 9162 27328 9196 27338
rect 9234 27328 9268 27338
rect 9306 27328 9340 27338
rect 9378 27328 9412 27338
rect 9450 27328 9484 27338
rect 9522 27328 9556 27338
rect 9594 27328 9628 27338
rect 9666 27328 9700 27338
rect 9738 27328 9772 27338
rect 9810 27328 9844 27338
rect 9882 27328 9916 27338
rect 9954 27328 9988 27362
rect 10026 27338 10056 27362
rect 10056 27338 10060 27362
rect 10098 27338 10124 27362
rect 10124 27338 10132 27362
rect 10170 27338 10192 27362
rect 10192 27338 10204 27362
rect 10242 27338 10260 27362
rect 10260 27338 10276 27362
rect 10314 27338 10328 27362
rect 10328 27338 10348 27362
rect 10386 27338 10396 27362
rect 10396 27338 10420 27362
rect 10458 27338 10464 27362
rect 10464 27338 10492 27362
rect 10530 27338 10532 27362
rect 10532 27338 10564 27362
rect 10602 27338 10634 27362
rect 10634 27338 10636 27362
rect 10674 27338 10702 27362
rect 10702 27338 10708 27362
rect 10746 27338 10770 27362
rect 10770 27338 10780 27362
rect 10818 27338 10838 27362
rect 10838 27338 10852 27362
rect 10890 27338 10906 27362
rect 10906 27338 10924 27362
rect 10962 27338 10974 27362
rect 10974 27338 10996 27362
rect 11034 27338 11042 27362
rect 11042 27338 11068 27362
rect 11106 27338 11110 27362
rect 11110 27338 11140 27362
rect 10026 27328 10060 27338
rect 10098 27328 10132 27338
rect 10170 27328 10204 27338
rect 10242 27328 10276 27338
rect 10314 27328 10348 27338
rect 10386 27328 10420 27338
rect 10458 27328 10492 27338
rect 10530 27328 10564 27338
rect 10602 27328 10636 27338
rect 10674 27328 10708 27338
rect 10746 27328 10780 27338
rect 10818 27328 10852 27338
rect 10890 27328 10924 27338
rect 10962 27328 10996 27338
rect 11034 27328 11068 27338
rect 11106 27328 11140 27338
rect 11178 27328 11212 27362
rect 11250 27338 11280 27362
rect 11280 27338 11284 27362
rect 11322 27338 11348 27362
rect 11348 27338 11356 27362
rect 11394 27338 11416 27362
rect 11416 27338 11428 27362
rect 11466 27338 11484 27362
rect 11484 27338 11500 27362
rect 11538 27338 11552 27362
rect 11552 27338 11572 27362
rect 11610 27338 11620 27362
rect 11620 27338 11644 27362
rect 11682 27338 11688 27362
rect 11688 27338 11716 27362
rect 11754 27338 11756 27362
rect 11756 27338 11788 27362
rect 11826 27338 11858 27362
rect 11858 27338 11860 27362
rect 11898 27338 11926 27362
rect 11926 27338 11932 27362
rect 11970 27338 11994 27362
rect 11994 27338 12004 27362
rect 12042 27338 12062 27362
rect 12062 27338 12076 27362
rect 12114 27338 12130 27362
rect 12130 27338 12148 27362
rect 12186 27338 12198 27362
rect 12198 27338 12220 27362
rect 12258 27338 12266 27362
rect 12266 27338 12292 27362
rect 12330 27338 12334 27362
rect 12334 27338 12364 27362
rect 11250 27328 11284 27338
rect 11322 27328 11356 27338
rect 11394 27328 11428 27338
rect 11466 27328 11500 27338
rect 11538 27328 11572 27338
rect 11610 27328 11644 27338
rect 11682 27328 11716 27338
rect 11754 27328 11788 27338
rect 11826 27328 11860 27338
rect 11898 27328 11932 27338
rect 11970 27328 12004 27338
rect 12042 27328 12076 27338
rect 12114 27328 12148 27338
rect 12186 27328 12220 27338
rect 12258 27328 12292 27338
rect 12330 27328 12364 27338
rect 12402 27328 12436 27362
rect 12474 27338 12504 27362
rect 12504 27338 12508 27362
rect 12546 27338 12572 27362
rect 12572 27338 12580 27362
rect 12618 27338 12640 27362
rect 12640 27338 12652 27362
rect 12690 27338 12708 27362
rect 12708 27338 12724 27362
rect 12762 27338 12776 27362
rect 12776 27338 12796 27362
rect 12834 27338 12844 27362
rect 12844 27338 12868 27362
rect 12906 27338 12912 27362
rect 12912 27338 12940 27362
rect 12978 27338 12980 27362
rect 12980 27338 13012 27362
rect 13050 27338 13082 27362
rect 13082 27338 13084 27362
rect 13122 27338 13150 27362
rect 13150 27338 13156 27362
rect 13194 27338 13218 27362
rect 13218 27338 13228 27362
rect 13266 27338 13286 27362
rect 13286 27338 13300 27362
rect 13338 27338 13354 27362
rect 13354 27338 13372 27362
rect 13410 27338 13422 27362
rect 13422 27338 13444 27362
rect 13482 27338 13490 27362
rect 13490 27338 13516 27362
rect 13554 27338 13558 27362
rect 13558 27338 13588 27362
rect 12474 27328 12508 27338
rect 12546 27328 12580 27338
rect 12618 27328 12652 27338
rect 12690 27328 12724 27338
rect 12762 27328 12796 27338
rect 12834 27328 12868 27338
rect 12906 27328 12940 27338
rect 12978 27328 13012 27338
rect 13050 27328 13084 27338
rect 13122 27328 13156 27338
rect 13194 27328 13228 27338
rect 13266 27328 13300 27338
rect 13338 27328 13372 27338
rect 13410 27328 13444 27338
rect 13482 27328 13516 27338
rect 13554 27328 13588 27338
rect 13626 27328 13660 27362
rect 13698 27338 13728 27362
rect 13728 27338 13732 27362
rect 13770 27338 13796 27362
rect 13796 27338 13804 27362
rect 13842 27338 13864 27362
rect 13864 27338 13876 27362
rect 13914 27338 13932 27362
rect 13932 27338 13948 27362
rect 13986 27338 14000 27362
rect 14000 27338 14020 27362
rect 14058 27338 14068 27362
rect 14068 27338 14092 27362
rect 14130 27338 14136 27362
rect 14136 27338 14164 27362
rect 14202 27338 14204 27362
rect 14204 27338 14236 27362
rect 14274 27338 14306 27362
rect 14306 27338 14308 27362
rect 14346 27338 14374 27362
rect 14374 27338 14380 27362
rect 14418 27338 14442 27362
rect 14442 27338 14452 27362
rect 14490 27338 14510 27362
rect 14510 27338 14524 27362
rect 14562 27338 14578 27362
rect 14578 27338 14596 27362
rect 14634 27338 14646 27362
rect 14646 27338 14668 27362
rect 14706 27338 14714 27362
rect 14714 27338 14740 27362
rect 14778 27338 14782 27362
rect 14782 27338 14812 27362
rect 13698 27328 13732 27338
rect 13770 27328 13804 27338
rect 13842 27328 13876 27338
rect 13914 27328 13948 27338
rect 13986 27328 14020 27338
rect 14058 27328 14092 27338
rect 14130 27328 14164 27338
rect 14202 27328 14236 27338
rect 14274 27328 14308 27338
rect 14346 27328 14380 27338
rect 14418 27328 14452 27338
rect 14490 27328 14524 27338
rect 14562 27328 14596 27338
rect 14634 27328 14668 27338
rect 14706 27328 14740 27338
rect 14778 27328 14812 27338
rect 14850 27328 14884 27362
rect 827 27228 861 27238
rect 899 27228 933 27238
rect 971 27228 1005 27238
rect 1043 27228 1077 27238
rect 1115 27228 1149 27238
rect 1187 27228 1221 27238
rect 1259 27228 1293 27238
rect 1331 27228 1365 27238
rect 1403 27228 1437 27238
rect 1475 27228 1509 27238
rect 1547 27228 1581 27238
rect 1619 27228 1653 27238
rect 1691 27228 1725 27238
rect 1764 27228 1798 27238
rect 1837 27228 1871 27238
rect 1910 27228 1944 27238
rect 1983 27228 2017 27238
rect 2056 27228 2090 27238
rect 3392 27232 3426 27238
rect 3465 27232 3499 27238
rect 3538 27232 3572 27238
rect 3611 27232 3645 27238
rect 3684 27232 3718 27238
rect 3757 27232 3791 27238
rect 3830 27232 3864 27238
rect 3903 27232 3937 27238
rect 3976 27232 4010 27238
rect 4049 27232 4083 27238
rect 4122 27232 4156 27238
rect 4194 27232 4228 27238
rect 4266 27232 4300 27238
rect 4338 27232 4372 27238
rect 4410 27232 4444 27238
rect 4482 27232 4516 27238
rect 4554 27232 4588 27238
rect 4626 27232 4660 27238
rect 4698 27232 4732 27238
rect 4770 27232 4804 27238
rect 4842 27232 4876 27238
rect 4914 27232 4948 27238
rect 4986 27232 5020 27238
rect 827 27204 842 27228
rect 842 27204 861 27228
rect 899 27204 911 27228
rect 911 27204 933 27228
rect 971 27204 980 27228
rect 980 27204 1005 27228
rect 1043 27204 1049 27228
rect 1049 27204 1077 27228
rect 1115 27204 1118 27228
rect 1118 27204 1149 27228
rect 1187 27204 1221 27228
rect 1259 27204 1290 27228
rect 1290 27204 1293 27228
rect 1331 27204 1359 27228
rect 1359 27204 1365 27228
rect 1403 27204 1428 27228
rect 1428 27204 1437 27228
rect 1475 27204 1497 27228
rect 1497 27204 1509 27228
rect 1547 27204 1566 27228
rect 1566 27204 1581 27228
rect 1619 27204 1635 27228
rect 1635 27204 1653 27228
rect 1691 27204 1704 27228
rect 1704 27204 1725 27228
rect 1764 27204 1773 27228
rect 1773 27204 1798 27228
rect 1837 27204 1842 27228
rect 1842 27204 1871 27228
rect 1910 27204 1911 27228
rect 1911 27204 1944 27228
rect 1983 27204 2014 27228
rect 2014 27204 2017 27228
rect 2056 27204 2082 27228
rect 2082 27204 2090 27228
rect 3392 27204 3426 27232
rect 3465 27204 3494 27232
rect 3494 27204 3499 27232
rect 3538 27204 3562 27232
rect 3562 27204 3572 27232
rect 3611 27204 3630 27232
rect 3630 27204 3645 27232
rect 3684 27204 3698 27232
rect 3698 27204 3718 27232
rect 3757 27204 3766 27232
rect 3766 27204 3791 27232
rect 3830 27204 3834 27232
rect 3834 27204 3864 27232
rect 3903 27204 3936 27232
rect 3936 27204 3937 27232
rect 3976 27204 4004 27232
rect 4004 27204 4010 27232
rect 4049 27204 4072 27232
rect 4072 27204 4083 27232
rect 4122 27204 4140 27232
rect 4140 27204 4156 27232
rect 4194 27204 4208 27232
rect 4208 27204 4228 27232
rect 4266 27204 4276 27232
rect 4276 27204 4300 27232
rect 4338 27204 4344 27232
rect 4344 27204 4372 27232
rect 4410 27204 4412 27232
rect 4412 27204 4444 27232
rect 4482 27204 4514 27232
rect 4514 27204 4516 27232
rect 4554 27204 4582 27232
rect 4582 27204 4588 27232
rect 4626 27204 4650 27232
rect 4650 27204 4660 27232
rect 4698 27204 4718 27232
rect 4718 27204 4732 27232
rect 4770 27204 4786 27232
rect 4786 27204 4804 27232
rect 4842 27204 4854 27232
rect 4854 27204 4876 27232
rect 4914 27204 4922 27232
rect 4922 27204 4948 27232
rect 4986 27204 4990 27232
rect 4990 27204 5020 27232
rect 5058 27204 5092 27238
rect 5130 27232 5164 27238
rect 5202 27232 5236 27238
rect 5274 27232 5308 27238
rect 5346 27232 5380 27238
rect 5418 27232 5452 27238
rect 5490 27232 5524 27238
rect 5562 27232 5596 27238
rect 5634 27232 5668 27238
rect 5706 27232 5740 27238
rect 5778 27232 5812 27238
rect 5850 27232 5884 27238
rect 5922 27232 5956 27238
rect 5994 27232 6028 27238
rect 6066 27232 6100 27238
rect 6138 27232 6172 27238
rect 6210 27232 6244 27238
rect 5130 27204 5160 27232
rect 5160 27204 5164 27232
rect 5202 27204 5228 27232
rect 5228 27204 5236 27232
rect 5274 27204 5296 27232
rect 5296 27204 5308 27232
rect 5346 27204 5364 27232
rect 5364 27204 5380 27232
rect 5418 27204 5432 27232
rect 5432 27204 5452 27232
rect 5490 27204 5500 27232
rect 5500 27204 5524 27232
rect 5562 27204 5568 27232
rect 5568 27204 5596 27232
rect 5634 27204 5636 27232
rect 5636 27204 5668 27232
rect 5706 27204 5738 27232
rect 5738 27204 5740 27232
rect 5778 27204 5806 27232
rect 5806 27204 5812 27232
rect 5850 27204 5874 27232
rect 5874 27204 5884 27232
rect 5922 27204 5942 27232
rect 5942 27204 5956 27232
rect 5994 27204 6010 27232
rect 6010 27204 6028 27232
rect 6066 27204 6078 27232
rect 6078 27204 6100 27232
rect 6138 27204 6146 27232
rect 6146 27204 6172 27232
rect 6210 27204 6214 27232
rect 6214 27204 6244 27232
rect 6282 27204 6316 27238
rect 6354 27232 6388 27238
rect 6426 27232 6460 27238
rect 6498 27232 6532 27238
rect 6570 27232 6604 27238
rect 6642 27232 6676 27238
rect 6714 27232 6748 27238
rect 6786 27232 6820 27238
rect 6858 27232 6892 27238
rect 6930 27232 6964 27238
rect 7002 27232 7036 27238
rect 7074 27232 7108 27238
rect 7146 27232 7180 27238
rect 7218 27232 7252 27238
rect 7290 27232 7324 27238
rect 7362 27232 7396 27238
rect 7434 27232 7468 27238
rect 6354 27204 6384 27232
rect 6384 27204 6388 27232
rect 6426 27204 6452 27232
rect 6452 27204 6460 27232
rect 6498 27204 6520 27232
rect 6520 27204 6532 27232
rect 6570 27204 6588 27232
rect 6588 27204 6604 27232
rect 6642 27204 6656 27232
rect 6656 27204 6676 27232
rect 6714 27204 6724 27232
rect 6724 27204 6748 27232
rect 6786 27204 6792 27232
rect 6792 27204 6820 27232
rect 6858 27204 6860 27232
rect 6860 27204 6892 27232
rect 6930 27204 6962 27232
rect 6962 27204 6964 27232
rect 7002 27204 7030 27232
rect 7030 27204 7036 27232
rect 7074 27204 7098 27232
rect 7098 27204 7108 27232
rect 7146 27204 7166 27232
rect 7166 27204 7180 27232
rect 7218 27204 7234 27232
rect 7234 27204 7252 27232
rect 7290 27204 7302 27232
rect 7302 27204 7324 27232
rect 7362 27204 7370 27232
rect 7370 27204 7396 27232
rect 7434 27204 7438 27232
rect 7438 27204 7468 27232
rect 7506 27204 7540 27238
rect 7578 27232 7612 27238
rect 7650 27232 7684 27238
rect 7722 27232 7756 27238
rect 7794 27232 7828 27238
rect 7866 27232 7900 27238
rect 7938 27232 7972 27238
rect 8010 27232 8044 27238
rect 8082 27232 8116 27238
rect 8154 27232 8188 27238
rect 8226 27232 8260 27238
rect 8298 27232 8332 27238
rect 8370 27232 8404 27238
rect 8442 27232 8476 27238
rect 8514 27232 8548 27238
rect 8586 27232 8620 27238
rect 8658 27232 8692 27238
rect 7578 27204 7608 27232
rect 7608 27204 7612 27232
rect 7650 27204 7676 27232
rect 7676 27204 7684 27232
rect 7722 27204 7744 27232
rect 7744 27204 7756 27232
rect 7794 27204 7812 27232
rect 7812 27204 7828 27232
rect 7866 27204 7880 27232
rect 7880 27204 7900 27232
rect 7938 27204 7948 27232
rect 7948 27204 7972 27232
rect 8010 27204 8016 27232
rect 8016 27204 8044 27232
rect 8082 27204 8084 27232
rect 8084 27204 8116 27232
rect 8154 27204 8186 27232
rect 8186 27204 8188 27232
rect 8226 27204 8254 27232
rect 8254 27204 8260 27232
rect 8298 27204 8322 27232
rect 8322 27204 8332 27232
rect 8370 27204 8390 27232
rect 8390 27204 8404 27232
rect 8442 27204 8458 27232
rect 8458 27204 8476 27232
rect 8514 27204 8526 27232
rect 8526 27204 8548 27232
rect 8586 27204 8594 27232
rect 8594 27204 8620 27232
rect 8658 27204 8662 27232
rect 8662 27204 8692 27232
rect 8730 27204 8764 27238
rect 8802 27232 8836 27238
rect 8874 27232 8908 27238
rect 8946 27232 8980 27238
rect 9018 27232 9052 27238
rect 9090 27232 9124 27238
rect 9162 27232 9196 27238
rect 9234 27232 9268 27238
rect 9306 27232 9340 27238
rect 9378 27232 9412 27238
rect 9450 27232 9484 27238
rect 9522 27232 9556 27238
rect 9594 27232 9628 27238
rect 9666 27232 9700 27238
rect 9738 27232 9772 27238
rect 9810 27232 9844 27238
rect 9882 27232 9916 27238
rect 8802 27204 8832 27232
rect 8832 27204 8836 27232
rect 8874 27204 8900 27232
rect 8900 27204 8908 27232
rect 8946 27204 8968 27232
rect 8968 27204 8980 27232
rect 9018 27204 9036 27232
rect 9036 27204 9052 27232
rect 9090 27204 9104 27232
rect 9104 27204 9124 27232
rect 9162 27204 9172 27232
rect 9172 27204 9196 27232
rect 9234 27204 9240 27232
rect 9240 27204 9268 27232
rect 9306 27204 9308 27232
rect 9308 27204 9340 27232
rect 9378 27204 9410 27232
rect 9410 27204 9412 27232
rect 9450 27204 9478 27232
rect 9478 27204 9484 27232
rect 9522 27204 9546 27232
rect 9546 27204 9556 27232
rect 9594 27204 9614 27232
rect 9614 27204 9628 27232
rect 9666 27204 9682 27232
rect 9682 27204 9700 27232
rect 9738 27204 9750 27232
rect 9750 27204 9772 27232
rect 9810 27204 9818 27232
rect 9818 27204 9844 27232
rect 9882 27204 9886 27232
rect 9886 27204 9916 27232
rect 9954 27204 9988 27238
rect 10026 27232 10060 27238
rect 10098 27232 10132 27238
rect 10170 27232 10204 27238
rect 10242 27232 10276 27238
rect 10314 27232 10348 27238
rect 10386 27232 10420 27238
rect 10458 27232 10492 27238
rect 10530 27232 10564 27238
rect 10602 27232 10636 27238
rect 10674 27232 10708 27238
rect 10746 27232 10780 27238
rect 10818 27232 10852 27238
rect 10890 27232 10924 27238
rect 10962 27232 10996 27238
rect 11034 27232 11068 27238
rect 11106 27232 11140 27238
rect 10026 27204 10056 27232
rect 10056 27204 10060 27232
rect 10098 27204 10124 27232
rect 10124 27204 10132 27232
rect 10170 27204 10192 27232
rect 10192 27204 10204 27232
rect 10242 27204 10260 27232
rect 10260 27204 10276 27232
rect 10314 27204 10328 27232
rect 10328 27204 10348 27232
rect 10386 27204 10396 27232
rect 10396 27204 10420 27232
rect 10458 27204 10464 27232
rect 10464 27204 10492 27232
rect 10530 27204 10532 27232
rect 10532 27204 10564 27232
rect 10602 27204 10634 27232
rect 10634 27204 10636 27232
rect 10674 27204 10702 27232
rect 10702 27204 10708 27232
rect 10746 27204 10770 27232
rect 10770 27204 10780 27232
rect 10818 27204 10838 27232
rect 10838 27204 10852 27232
rect 10890 27204 10906 27232
rect 10906 27204 10924 27232
rect 10962 27204 10974 27232
rect 10974 27204 10996 27232
rect 11034 27204 11042 27232
rect 11042 27204 11068 27232
rect 11106 27204 11110 27232
rect 11110 27204 11140 27232
rect 11178 27204 11212 27238
rect 11250 27232 11284 27238
rect 11322 27232 11356 27238
rect 11394 27232 11428 27238
rect 11466 27232 11500 27238
rect 11538 27232 11572 27238
rect 11610 27232 11644 27238
rect 11682 27232 11716 27238
rect 11754 27232 11788 27238
rect 11826 27232 11860 27238
rect 11898 27232 11932 27238
rect 11970 27232 12004 27238
rect 12042 27232 12076 27238
rect 12114 27232 12148 27238
rect 12186 27232 12220 27238
rect 12258 27232 12292 27238
rect 12330 27232 12364 27238
rect 11250 27204 11280 27232
rect 11280 27204 11284 27232
rect 11322 27204 11348 27232
rect 11348 27204 11356 27232
rect 11394 27204 11416 27232
rect 11416 27204 11428 27232
rect 11466 27204 11484 27232
rect 11484 27204 11500 27232
rect 11538 27204 11552 27232
rect 11552 27204 11572 27232
rect 11610 27204 11620 27232
rect 11620 27204 11644 27232
rect 11682 27204 11688 27232
rect 11688 27204 11716 27232
rect 11754 27204 11756 27232
rect 11756 27204 11788 27232
rect 11826 27204 11858 27232
rect 11858 27204 11860 27232
rect 11898 27204 11926 27232
rect 11926 27204 11932 27232
rect 11970 27204 11994 27232
rect 11994 27204 12004 27232
rect 12042 27204 12062 27232
rect 12062 27204 12076 27232
rect 12114 27204 12130 27232
rect 12130 27204 12148 27232
rect 12186 27204 12198 27232
rect 12198 27204 12220 27232
rect 12258 27204 12266 27232
rect 12266 27204 12292 27232
rect 12330 27204 12334 27232
rect 12334 27204 12364 27232
rect 12402 27204 12436 27238
rect 12474 27232 12508 27238
rect 12546 27232 12580 27238
rect 12618 27232 12652 27238
rect 12690 27232 12724 27238
rect 12762 27232 12796 27238
rect 12834 27232 12868 27238
rect 12906 27232 12940 27238
rect 12978 27232 13012 27238
rect 13050 27232 13084 27238
rect 13122 27232 13156 27238
rect 13194 27232 13228 27238
rect 13266 27232 13300 27238
rect 13338 27232 13372 27238
rect 13410 27232 13444 27238
rect 13482 27232 13516 27238
rect 13554 27232 13588 27238
rect 12474 27204 12504 27232
rect 12504 27204 12508 27232
rect 12546 27204 12572 27232
rect 12572 27204 12580 27232
rect 12618 27204 12640 27232
rect 12640 27204 12652 27232
rect 12690 27204 12708 27232
rect 12708 27204 12724 27232
rect 12762 27204 12776 27232
rect 12776 27204 12796 27232
rect 12834 27204 12844 27232
rect 12844 27204 12868 27232
rect 12906 27204 12912 27232
rect 12912 27204 12940 27232
rect 12978 27204 12980 27232
rect 12980 27204 13012 27232
rect 13050 27204 13082 27232
rect 13082 27204 13084 27232
rect 13122 27204 13150 27232
rect 13150 27204 13156 27232
rect 13194 27204 13218 27232
rect 13218 27204 13228 27232
rect 13266 27204 13286 27232
rect 13286 27204 13300 27232
rect 13338 27204 13354 27232
rect 13354 27204 13372 27232
rect 13410 27204 13422 27232
rect 13422 27204 13444 27232
rect 13482 27204 13490 27232
rect 13490 27204 13516 27232
rect 13554 27204 13558 27232
rect 13558 27204 13588 27232
rect 13626 27204 13660 27238
rect 13698 27232 13732 27238
rect 13770 27232 13804 27238
rect 13842 27232 13876 27238
rect 13914 27232 13948 27238
rect 13986 27232 14020 27238
rect 14058 27232 14092 27238
rect 14130 27232 14164 27238
rect 14202 27232 14236 27238
rect 14274 27232 14308 27238
rect 14346 27232 14380 27238
rect 14418 27232 14452 27238
rect 14490 27232 14524 27238
rect 14562 27232 14596 27238
rect 14634 27232 14668 27238
rect 14706 27232 14740 27238
rect 14778 27232 14812 27238
rect 13698 27204 13728 27232
rect 13728 27204 13732 27232
rect 13770 27204 13796 27232
rect 13796 27204 13804 27232
rect 13842 27204 13864 27232
rect 13864 27204 13876 27232
rect 13914 27204 13932 27232
rect 13932 27204 13948 27232
rect 13986 27204 14000 27232
rect 14000 27204 14020 27232
rect 14058 27204 14068 27232
rect 14068 27204 14092 27232
rect 14130 27204 14136 27232
rect 14136 27204 14164 27232
rect 14202 27204 14204 27232
rect 14204 27204 14236 27232
rect 14274 27204 14306 27232
rect 14306 27204 14308 27232
rect 14346 27204 14374 27232
rect 14374 27204 14380 27232
rect 14418 27204 14442 27232
rect 14442 27204 14452 27232
rect 14490 27204 14510 27232
rect 14510 27204 14524 27232
rect 14562 27204 14578 27232
rect 14578 27204 14596 27232
rect 14634 27204 14646 27232
rect 14646 27204 14668 27232
rect 14706 27204 14714 27232
rect 14714 27204 14740 27232
rect 14778 27204 14782 27232
rect 14782 27204 14812 27232
rect 14850 27204 14884 27238
rect 243 26172 277 26185
rect 316 26172 350 26185
rect 389 26172 423 26185
rect 462 26172 496 26185
rect 535 26172 569 26185
rect 608 26172 642 26185
rect 681 26172 715 26185
rect 754 26172 788 26185
rect 827 26172 861 26185
rect 900 26172 934 26185
rect 973 26172 1007 26185
rect 1046 26172 1080 26185
rect 1119 26172 1153 26185
rect 1192 26172 1226 26185
rect 1265 26172 1299 26185
rect 1338 26172 1372 26185
rect 1411 26172 1445 26185
rect 243 26151 276 26172
rect 276 26151 277 26172
rect 316 26151 345 26172
rect 345 26151 350 26172
rect 389 26151 414 26172
rect 414 26151 423 26172
rect 462 26151 483 26172
rect 483 26151 496 26172
rect 535 26151 552 26172
rect 552 26151 569 26172
rect 608 26151 621 26172
rect 621 26151 642 26172
rect 681 26151 690 26172
rect 690 26151 715 26172
rect 754 26151 759 26172
rect 759 26151 788 26172
rect 827 26151 828 26172
rect 828 26151 861 26172
rect 900 26151 931 26172
rect 931 26151 934 26172
rect 973 26151 1000 26172
rect 1000 26151 1007 26172
rect 1046 26151 1069 26172
rect 1069 26151 1080 26172
rect 1119 26151 1138 26172
rect 1138 26151 1153 26172
rect 1192 26151 1207 26172
rect 1207 26151 1226 26172
rect 1265 26151 1276 26172
rect 1276 26151 1299 26172
rect 1338 26151 1345 26172
rect 1345 26151 1372 26172
rect 1411 26151 1414 26172
rect 1414 26151 1445 26172
rect 1484 26151 1518 26185
rect 1557 26172 1591 26185
rect 1630 26172 1664 26185
rect 1703 26172 1737 26185
rect 1776 26172 1810 26185
rect 1849 26172 1883 26185
rect 1922 26172 1956 26185
rect 1995 26172 2029 26185
rect 2068 26172 2102 26185
rect 2141 26172 2175 26185
rect 2214 26172 2248 26185
rect 2287 26172 2321 26185
rect 2360 26172 2394 26185
rect 2433 26172 2467 26185
rect 2506 26172 2540 26185
rect 2579 26172 2613 26185
rect 2652 26172 2686 26185
rect 1557 26151 1587 26172
rect 1587 26151 1591 26172
rect 1630 26151 1656 26172
rect 1656 26151 1664 26172
rect 1703 26151 1725 26172
rect 1725 26151 1737 26172
rect 1776 26151 1794 26172
rect 1794 26151 1810 26172
rect 1849 26151 1863 26172
rect 1863 26151 1883 26172
rect 1922 26151 1932 26172
rect 1932 26151 1956 26172
rect 1995 26151 2001 26172
rect 2001 26151 2029 26172
rect 2068 26151 2070 26172
rect 2070 26151 2102 26172
rect 2141 26151 2173 26172
rect 2173 26151 2175 26172
rect 2214 26151 2242 26172
rect 2242 26151 2248 26172
rect 2287 26151 2311 26172
rect 2311 26151 2321 26172
rect 2360 26151 2380 26172
rect 2380 26151 2394 26172
rect 2433 26151 2449 26172
rect 2449 26151 2467 26172
rect 2506 26151 2518 26172
rect 2518 26151 2540 26172
rect 2579 26151 2587 26172
rect 2587 26151 2613 26172
rect 2652 26151 2656 26172
rect 2656 26151 2686 26172
rect 2725 26151 2759 26185
rect 2798 26172 2832 26185
rect 2871 26172 2905 26185
rect 2944 26172 2978 26185
rect 3017 26172 3051 26185
rect 3090 26172 3124 26185
rect 3163 26172 3197 26185
rect 3236 26172 3270 26185
rect 3309 26172 3343 26185
rect 3382 26172 3416 26185
rect 3455 26172 3489 26185
rect 3528 26172 3562 26185
rect 3601 26172 3635 26185
rect 3674 26172 3708 26185
rect 3746 26172 3780 26185
rect 3818 26172 3852 26185
rect 3890 26172 3924 26185
rect 3962 26172 3996 26185
rect 4034 26172 4068 26185
rect 2798 26151 2829 26172
rect 2829 26151 2832 26172
rect 2871 26151 2898 26172
rect 2898 26151 2905 26172
rect 2944 26151 2967 26172
rect 2967 26151 2978 26172
rect 3017 26151 3036 26172
rect 3036 26151 3051 26172
rect 3090 26151 3105 26172
rect 3105 26151 3124 26172
rect 3163 26151 3174 26172
rect 3174 26151 3197 26172
rect 3236 26151 3243 26172
rect 3243 26151 3270 26172
rect 3309 26151 3312 26172
rect 3312 26151 3343 26172
rect 3382 26151 3415 26172
rect 3415 26151 3416 26172
rect 3455 26151 3484 26172
rect 3484 26151 3489 26172
rect 3528 26151 3553 26172
rect 3553 26151 3562 26172
rect 3601 26151 3622 26172
rect 3622 26151 3635 26172
rect 3674 26151 3691 26172
rect 3691 26151 3708 26172
rect 3746 26151 3760 26172
rect 3760 26151 3780 26172
rect 3818 26151 3829 26172
rect 3829 26151 3852 26172
rect 3890 26151 3898 26172
rect 3898 26151 3924 26172
rect 3962 26151 3967 26172
rect 3967 26151 3996 26172
rect 4034 26151 4036 26172
rect 4036 26151 4068 26172
rect 4106 26151 4140 26185
rect 4178 26172 4212 26185
rect 4250 26172 4284 26185
rect 4322 26172 4356 26185
rect 4394 26172 4428 26185
rect 4466 26172 4500 26185
rect 4538 26172 4572 26185
rect 4610 26172 4644 26185
rect 4682 26172 4716 26185
rect 4754 26172 4788 26185
rect 4826 26172 4860 26185
rect 4898 26172 4932 26185
rect 4970 26172 5004 26185
rect 5042 26172 5076 26185
rect 5114 26172 5148 26185
rect 5186 26172 5220 26185
rect 5258 26172 5292 26185
rect 4178 26151 4208 26172
rect 4208 26151 4212 26172
rect 4250 26151 4276 26172
rect 4276 26151 4284 26172
rect 4322 26151 4344 26172
rect 4344 26151 4356 26172
rect 4394 26151 4412 26172
rect 4412 26151 4428 26172
rect 4466 26151 4480 26172
rect 4480 26151 4500 26172
rect 4538 26151 4548 26172
rect 4548 26151 4572 26172
rect 4610 26151 4616 26172
rect 4616 26151 4644 26172
rect 4682 26151 4684 26172
rect 4684 26151 4716 26172
rect 4754 26151 4786 26172
rect 4786 26151 4788 26172
rect 4826 26151 4854 26172
rect 4854 26151 4860 26172
rect 4898 26151 4922 26172
rect 4922 26151 4932 26172
rect 4970 26151 4990 26172
rect 4990 26151 5004 26172
rect 5042 26151 5058 26172
rect 5058 26151 5076 26172
rect 5114 26151 5126 26172
rect 5126 26151 5148 26172
rect 5186 26151 5194 26172
rect 5194 26151 5220 26172
rect 5258 26151 5262 26172
rect 5262 26151 5292 26172
rect 5330 26151 5364 26185
rect 5402 26172 5436 26185
rect 5474 26172 5508 26185
rect 5546 26172 5580 26185
rect 5618 26172 5652 26185
rect 5690 26172 5724 26185
rect 5762 26172 5796 26185
rect 5834 26172 5868 26185
rect 5906 26172 5940 26185
rect 5978 26172 6012 26185
rect 6050 26172 6084 26185
rect 6122 26172 6156 26185
rect 6194 26172 6228 26185
rect 6266 26172 6300 26185
rect 6338 26172 6372 26185
rect 6410 26172 6444 26185
rect 6482 26172 6516 26185
rect 5402 26151 5432 26172
rect 5432 26151 5436 26172
rect 5474 26151 5500 26172
rect 5500 26151 5508 26172
rect 5546 26151 5568 26172
rect 5568 26151 5580 26172
rect 5618 26151 5636 26172
rect 5636 26151 5652 26172
rect 5690 26151 5704 26172
rect 5704 26151 5724 26172
rect 5762 26151 5772 26172
rect 5772 26151 5796 26172
rect 5834 26151 5840 26172
rect 5840 26151 5868 26172
rect 5906 26151 5908 26172
rect 5908 26151 5940 26172
rect 5978 26151 6010 26172
rect 6010 26151 6012 26172
rect 6050 26151 6078 26172
rect 6078 26151 6084 26172
rect 6122 26151 6146 26172
rect 6146 26151 6156 26172
rect 6194 26151 6214 26172
rect 6214 26151 6228 26172
rect 6266 26151 6282 26172
rect 6282 26151 6300 26172
rect 6338 26151 6350 26172
rect 6350 26151 6372 26172
rect 6410 26151 6418 26172
rect 6418 26151 6444 26172
rect 6482 26151 6486 26172
rect 6486 26151 6516 26172
rect 6554 26151 6588 26185
rect 6626 26172 6660 26185
rect 6698 26172 6732 26185
rect 6770 26172 6804 26185
rect 6842 26172 6876 26185
rect 6914 26172 6948 26185
rect 6986 26172 7020 26185
rect 7058 26172 7092 26185
rect 7130 26172 7164 26185
rect 7202 26172 7236 26185
rect 7274 26172 7308 26185
rect 7346 26172 7380 26185
rect 7418 26172 7452 26185
rect 7490 26172 7524 26185
rect 7562 26172 7596 26185
rect 7634 26172 7668 26185
rect 7706 26172 7740 26185
rect 6626 26151 6656 26172
rect 6656 26151 6660 26172
rect 6698 26151 6724 26172
rect 6724 26151 6732 26172
rect 6770 26151 6792 26172
rect 6792 26151 6804 26172
rect 6842 26151 6860 26172
rect 6860 26151 6876 26172
rect 6914 26151 6928 26172
rect 6928 26151 6948 26172
rect 6986 26151 6996 26172
rect 6996 26151 7020 26172
rect 7058 26151 7064 26172
rect 7064 26151 7092 26172
rect 7130 26151 7132 26172
rect 7132 26151 7164 26172
rect 7202 26151 7234 26172
rect 7234 26151 7236 26172
rect 7274 26151 7302 26172
rect 7302 26151 7308 26172
rect 7346 26151 7370 26172
rect 7370 26151 7380 26172
rect 7418 26151 7438 26172
rect 7438 26151 7452 26172
rect 7490 26151 7506 26172
rect 7506 26151 7524 26172
rect 7562 26151 7574 26172
rect 7574 26151 7596 26172
rect 7634 26151 7642 26172
rect 7642 26151 7668 26172
rect 7706 26151 7710 26172
rect 7710 26151 7740 26172
rect 7778 26151 7812 26185
rect 7850 26172 7884 26185
rect 7922 26172 7956 26185
rect 7994 26172 8028 26185
rect 8066 26172 8100 26185
rect 8138 26172 8172 26185
rect 8210 26172 8244 26185
rect 8282 26172 8316 26185
rect 8354 26172 8388 26185
rect 8426 26172 8460 26185
rect 8498 26172 8532 26185
rect 8570 26172 8604 26185
rect 8642 26172 8676 26185
rect 8714 26172 8748 26185
rect 8786 26172 8820 26185
rect 8858 26172 8892 26185
rect 8930 26172 8964 26185
rect 7850 26151 7880 26172
rect 7880 26151 7884 26172
rect 7922 26151 7948 26172
rect 7948 26151 7956 26172
rect 7994 26151 8016 26172
rect 8016 26151 8028 26172
rect 8066 26151 8084 26172
rect 8084 26151 8100 26172
rect 8138 26151 8152 26172
rect 8152 26151 8172 26172
rect 8210 26151 8220 26172
rect 8220 26151 8244 26172
rect 8282 26151 8288 26172
rect 8288 26151 8316 26172
rect 8354 26151 8356 26172
rect 8356 26151 8388 26172
rect 8426 26151 8458 26172
rect 8458 26151 8460 26172
rect 8498 26151 8526 26172
rect 8526 26151 8532 26172
rect 8570 26151 8594 26172
rect 8594 26151 8604 26172
rect 8642 26151 8662 26172
rect 8662 26151 8676 26172
rect 8714 26151 8730 26172
rect 8730 26151 8748 26172
rect 8786 26151 8798 26172
rect 8798 26151 8820 26172
rect 8858 26151 8866 26172
rect 8866 26151 8892 26172
rect 8930 26151 8934 26172
rect 8934 26151 8964 26172
rect 9002 26151 9036 26185
rect 9074 26172 9108 26185
rect 9146 26172 9180 26185
rect 9218 26172 9252 26185
rect 9290 26172 9324 26185
rect 9362 26172 9396 26185
rect 9434 26172 9468 26185
rect 9506 26172 9540 26185
rect 9578 26172 9612 26185
rect 9650 26172 9684 26185
rect 9722 26172 9756 26185
rect 9794 26172 9828 26185
rect 9866 26172 9900 26185
rect 9938 26172 9972 26185
rect 10010 26172 10044 26185
rect 10082 26172 10116 26185
rect 10154 26172 10188 26185
rect 9074 26151 9104 26172
rect 9104 26151 9108 26172
rect 9146 26151 9172 26172
rect 9172 26151 9180 26172
rect 9218 26151 9240 26172
rect 9240 26151 9252 26172
rect 9290 26151 9308 26172
rect 9308 26151 9324 26172
rect 9362 26151 9376 26172
rect 9376 26151 9396 26172
rect 9434 26151 9444 26172
rect 9444 26151 9468 26172
rect 9506 26151 9512 26172
rect 9512 26151 9540 26172
rect 9578 26151 9580 26172
rect 9580 26151 9612 26172
rect 9650 26151 9682 26172
rect 9682 26151 9684 26172
rect 9722 26151 9750 26172
rect 9750 26151 9756 26172
rect 9794 26151 9818 26172
rect 9818 26151 9828 26172
rect 9866 26151 9886 26172
rect 9886 26151 9900 26172
rect 9938 26151 9954 26172
rect 9954 26151 9972 26172
rect 10010 26151 10022 26172
rect 10022 26151 10044 26172
rect 10082 26151 10090 26172
rect 10090 26151 10116 26172
rect 10154 26151 10158 26172
rect 10158 26151 10188 26172
rect 10226 26151 10260 26185
rect 10298 26172 10332 26185
rect 10370 26172 10404 26185
rect 10442 26172 10476 26185
rect 10514 26172 10548 26185
rect 10586 26172 10620 26185
rect 10658 26172 10692 26185
rect 10730 26172 10764 26185
rect 10802 26172 10836 26185
rect 10874 26172 10908 26185
rect 10946 26172 10980 26185
rect 11018 26172 11052 26185
rect 11090 26172 11124 26185
rect 11162 26172 11196 26185
rect 11234 26172 11268 26185
rect 11306 26172 11340 26185
rect 11378 26172 11412 26185
rect 10298 26151 10328 26172
rect 10328 26151 10332 26172
rect 10370 26151 10396 26172
rect 10396 26151 10404 26172
rect 10442 26151 10464 26172
rect 10464 26151 10476 26172
rect 10514 26151 10532 26172
rect 10532 26151 10548 26172
rect 10586 26151 10600 26172
rect 10600 26151 10620 26172
rect 10658 26151 10668 26172
rect 10668 26151 10692 26172
rect 10730 26151 10736 26172
rect 10736 26151 10764 26172
rect 10802 26151 10804 26172
rect 10804 26151 10836 26172
rect 10874 26151 10906 26172
rect 10906 26151 10908 26172
rect 10946 26151 10974 26172
rect 10974 26151 10980 26172
rect 11018 26151 11042 26172
rect 11042 26151 11052 26172
rect 11090 26151 11110 26172
rect 11110 26151 11124 26172
rect 11162 26151 11178 26172
rect 11178 26151 11196 26172
rect 11234 26151 11246 26172
rect 11246 26151 11268 26172
rect 11306 26151 11314 26172
rect 11314 26151 11340 26172
rect 11378 26151 11382 26172
rect 11382 26151 11412 26172
rect 11450 26151 11484 26185
rect 11522 26172 11556 26185
rect 11594 26172 11628 26185
rect 11666 26172 11700 26185
rect 11738 26172 11772 26185
rect 11810 26172 11844 26185
rect 11882 26172 11916 26185
rect 11954 26172 11988 26185
rect 12026 26172 12060 26185
rect 12098 26172 12132 26185
rect 12170 26172 12204 26185
rect 12242 26172 12276 26185
rect 12314 26172 12348 26185
rect 12386 26172 12420 26185
rect 12458 26172 12492 26185
rect 12530 26172 12564 26185
rect 12602 26172 12636 26185
rect 11522 26151 11552 26172
rect 11552 26151 11556 26172
rect 11594 26151 11620 26172
rect 11620 26151 11628 26172
rect 11666 26151 11688 26172
rect 11688 26151 11700 26172
rect 11738 26151 11756 26172
rect 11756 26151 11772 26172
rect 11810 26151 11824 26172
rect 11824 26151 11844 26172
rect 11882 26151 11892 26172
rect 11892 26151 11916 26172
rect 11954 26151 11960 26172
rect 11960 26151 11988 26172
rect 12026 26151 12028 26172
rect 12028 26151 12060 26172
rect 12098 26151 12130 26172
rect 12130 26151 12132 26172
rect 12170 26151 12198 26172
rect 12198 26151 12204 26172
rect 12242 26151 12266 26172
rect 12266 26151 12276 26172
rect 12314 26151 12334 26172
rect 12334 26151 12348 26172
rect 12386 26151 12402 26172
rect 12402 26151 12420 26172
rect 12458 26151 12470 26172
rect 12470 26151 12492 26172
rect 12530 26151 12538 26172
rect 12538 26151 12564 26172
rect 12602 26151 12606 26172
rect 12606 26151 12636 26172
rect 12674 26151 12708 26185
rect 12746 26172 12780 26185
rect 12818 26172 12852 26185
rect 12890 26172 12924 26185
rect 12962 26172 12996 26185
rect 13034 26172 13068 26185
rect 13106 26172 13140 26185
rect 13178 26172 13212 26185
rect 13250 26172 13284 26185
rect 13322 26172 13356 26185
rect 13394 26172 13428 26185
rect 13466 26172 13500 26185
rect 13538 26172 13572 26185
rect 13610 26172 13644 26185
rect 13682 26172 13716 26185
rect 13754 26172 13788 26185
rect 13826 26172 13860 26185
rect 12746 26151 12776 26172
rect 12776 26151 12780 26172
rect 12818 26151 12844 26172
rect 12844 26151 12852 26172
rect 12890 26151 12912 26172
rect 12912 26151 12924 26172
rect 12962 26151 12980 26172
rect 12980 26151 12996 26172
rect 13034 26151 13048 26172
rect 13048 26151 13068 26172
rect 13106 26151 13116 26172
rect 13116 26151 13140 26172
rect 13178 26151 13184 26172
rect 13184 26151 13212 26172
rect 13250 26151 13252 26172
rect 13252 26151 13284 26172
rect 13322 26151 13354 26172
rect 13354 26151 13356 26172
rect 13394 26151 13422 26172
rect 13422 26151 13428 26172
rect 13466 26151 13490 26172
rect 13490 26151 13500 26172
rect 13538 26151 13558 26172
rect 13558 26151 13572 26172
rect 13610 26151 13626 26172
rect 13626 26151 13644 26172
rect 13682 26151 13694 26172
rect 13694 26151 13716 26172
rect 13754 26151 13762 26172
rect 13762 26151 13788 26172
rect 13826 26151 13830 26172
rect 13830 26151 13860 26172
rect 13898 26151 13932 26185
rect 13970 26172 14004 26185
rect 14042 26172 14076 26185
rect 14114 26172 14148 26185
rect 14186 26172 14220 26185
rect 14258 26172 14292 26185
rect 14330 26172 14364 26185
rect 14402 26172 14436 26185
rect 14474 26172 14508 26185
rect 14546 26172 14580 26185
rect 14618 26172 14652 26185
rect 14690 26172 14724 26185
rect 13970 26151 14000 26172
rect 14000 26151 14004 26172
rect 14042 26151 14068 26172
rect 14068 26151 14076 26172
rect 14114 26151 14136 26172
rect 14136 26151 14148 26172
rect 14186 26151 14204 26172
rect 14204 26151 14220 26172
rect 14258 26151 14272 26172
rect 14272 26151 14292 26172
rect 14330 26151 14340 26172
rect 14340 26151 14364 26172
rect 14402 26151 14408 26172
rect 14408 26151 14436 26172
rect 14474 26151 14476 26172
rect 14476 26151 14508 26172
rect 14546 26151 14578 26172
rect 14578 26151 14580 26172
rect 14618 26151 14646 26172
rect 14646 26151 14652 26172
rect 14690 26151 14714 26172
rect 14714 26151 14724 26172
rect 243 26100 277 26111
rect 316 26100 350 26111
rect 389 26100 423 26111
rect 462 26100 496 26111
rect 535 26100 569 26111
rect 608 26100 642 26111
rect 681 26100 715 26111
rect 754 26100 788 26111
rect 827 26100 861 26111
rect 900 26100 934 26111
rect 973 26100 1007 26111
rect 1046 26100 1080 26111
rect 1119 26100 1153 26111
rect 1192 26100 1226 26111
rect 1265 26100 1299 26111
rect 1338 26100 1372 26111
rect 1411 26100 1445 26111
rect 243 26077 276 26100
rect 276 26077 277 26100
rect 316 26077 345 26100
rect 345 26077 350 26100
rect 389 26077 414 26100
rect 414 26077 423 26100
rect 462 26077 483 26100
rect 483 26077 496 26100
rect 535 26077 552 26100
rect 552 26077 569 26100
rect 608 26077 621 26100
rect 621 26077 642 26100
rect 681 26077 690 26100
rect 690 26077 715 26100
rect 754 26077 759 26100
rect 759 26077 788 26100
rect 827 26077 828 26100
rect 828 26077 861 26100
rect 900 26077 931 26100
rect 931 26077 934 26100
rect 973 26077 1000 26100
rect 1000 26077 1007 26100
rect 1046 26077 1069 26100
rect 1069 26077 1080 26100
rect 1119 26077 1138 26100
rect 1138 26077 1153 26100
rect 1192 26077 1207 26100
rect 1207 26077 1226 26100
rect 1265 26077 1276 26100
rect 1276 26077 1299 26100
rect 1338 26077 1345 26100
rect 1345 26077 1372 26100
rect 1411 26077 1414 26100
rect 1414 26077 1445 26100
rect 1484 26077 1518 26111
rect 1557 26100 1591 26111
rect 1630 26100 1664 26111
rect 1703 26100 1737 26111
rect 1776 26100 1810 26111
rect 1849 26100 1883 26111
rect 1922 26100 1956 26111
rect 1995 26100 2029 26111
rect 2068 26100 2102 26111
rect 2141 26100 2175 26111
rect 2214 26100 2248 26111
rect 2287 26100 2321 26111
rect 2360 26100 2394 26111
rect 2433 26100 2467 26111
rect 2506 26100 2540 26111
rect 2579 26100 2613 26111
rect 2652 26100 2686 26111
rect 1557 26077 1587 26100
rect 1587 26077 1591 26100
rect 1630 26077 1656 26100
rect 1656 26077 1664 26100
rect 1703 26077 1725 26100
rect 1725 26077 1737 26100
rect 1776 26077 1794 26100
rect 1794 26077 1810 26100
rect 1849 26077 1863 26100
rect 1863 26077 1883 26100
rect 1922 26077 1932 26100
rect 1932 26077 1956 26100
rect 1995 26077 2001 26100
rect 2001 26077 2029 26100
rect 2068 26077 2070 26100
rect 2070 26077 2102 26100
rect 2141 26077 2173 26100
rect 2173 26077 2175 26100
rect 2214 26077 2242 26100
rect 2242 26077 2248 26100
rect 2287 26077 2311 26100
rect 2311 26077 2321 26100
rect 2360 26077 2380 26100
rect 2380 26077 2394 26100
rect 2433 26077 2449 26100
rect 2449 26077 2467 26100
rect 2506 26077 2518 26100
rect 2518 26077 2540 26100
rect 2579 26077 2587 26100
rect 2587 26077 2613 26100
rect 2652 26077 2656 26100
rect 2656 26077 2686 26100
rect 2725 26077 2759 26111
rect 2798 26100 2832 26111
rect 2871 26100 2905 26111
rect 2944 26100 2978 26111
rect 3017 26100 3051 26111
rect 3090 26100 3124 26111
rect 3163 26100 3197 26111
rect 3236 26100 3270 26111
rect 3309 26100 3343 26111
rect 3382 26100 3416 26111
rect 3455 26100 3489 26111
rect 3528 26100 3562 26111
rect 3601 26100 3635 26111
rect 3674 26100 3708 26111
rect 3746 26100 3780 26111
rect 3818 26100 3852 26111
rect 3890 26100 3924 26111
rect 3962 26100 3996 26111
rect 4034 26100 4068 26111
rect 2798 26077 2829 26100
rect 2829 26077 2832 26100
rect 2871 26077 2898 26100
rect 2898 26077 2905 26100
rect 2944 26077 2967 26100
rect 2967 26077 2978 26100
rect 3017 26077 3036 26100
rect 3036 26077 3051 26100
rect 3090 26077 3105 26100
rect 3105 26077 3124 26100
rect 3163 26077 3174 26100
rect 3174 26077 3197 26100
rect 3236 26077 3243 26100
rect 3243 26077 3270 26100
rect 3309 26077 3312 26100
rect 3312 26077 3343 26100
rect 3382 26077 3415 26100
rect 3415 26077 3416 26100
rect 3455 26077 3484 26100
rect 3484 26077 3489 26100
rect 3528 26077 3553 26100
rect 3553 26077 3562 26100
rect 3601 26077 3622 26100
rect 3622 26077 3635 26100
rect 3674 26077 3691 26100
rect 3691 26077 3708 26100
rect 3746 26077 3760 26100
rect 3760 26077 3780 26100
rect 3818 26077 3829 26100
rect 3829 26077 3852 26100
rect 3890 26077 3898 26100
rect 3898 26077 3924 26100
rect 3962 26077 3967 26100
rect 3967 26077 3996 26100
rect 4034 26077 4036 26100
rect 4036 26077 4068 26100
rect 4106 26077 4140 26111
rect 4178 26100 4212 26111
rect 4250 26100 4284 26111
rect 4322 26100 4356 26111
rect 4394 26100 4428 26111
rect 4466 26100 4500 26111
rect 4538 26100 4572 26111
rect 4610 26100 4644 26111
rect 4682 26100 4716 26111
rect 4754 26100 4788 26111
rect 4826 26100 4860 26111
rect 4898 26100 4932 26111
rect 4970 26100 5004 26111
rect 5042 26100 5076 26111
rect 5114 26100 5148 26111
rect 5186 26100 5220 26111
rect 5258 26100 5292 26111
rect 4178 26077 4208 26100
rect 4208 26077 4212 26100
rect 4250 26077 4276 26100
rect 4276 26077 4284 26100
rect 4322 26077 4344 26100
rect 4344 26077 4356 26100
rect 4394 26077 4412 26100
rect 4412 26077 4428 26100
rect 4466 26077 4480 26100
rect 4480 26077 4500 26100
rect 4538 26077 4548 26100
rect 4548 26077 4572 26100
rect 4610 26077 4616 26100
rect 4616 26077 4644 26100
rect 4682 26077 4684 26100
rect 4684 26077 4716 26100
rect 4754 26077 4786 26100
rect 4786 26077 4788 26100
rect 4826 26077 4854 26100
rect 4854 26077 4860 26100
rect 4898 26077 4922 26100
rect 4922 26077 4932 26100
rect 4970 26077 4990 26100
rect 4990 26077 5004 26100
rect 5042 26077 5058 26100
rect 5058 26077 5076 26100
rect 5114 26077 5126 26100
rect 5126 26077 5148 26100
rect 5186 26077 5194 26100
rect 5194 26077 5220 26100
rect 5258 26077 5262 26100
rect 5262 26077 5292 26100
rect 5330 26077 5364 26111
rect 5402 26100 5436 26111
rect 5474 26100 5508 26111
rect 5546 26100 5580 26111
rect 5618 26100 5652 26111
rect 5690 26100 5724 26111
rect 5762 26100 5796 26111
rect 5834 26100 5868 26111
rect 5906 26100 5940 26111
rect 5978 26100 6012 26111
rect 6050 26100 6084 26111
rect 6122 26100 6156 26111
rect 6194 26100 6228 26111
rect 6266 26100 6300 26111
rect 6338 26100 6372 26111
rect 6410 26100 6444 26111
rect 6482 26100 6516 26111
rect 5402 26077 5432 26100
rect 5432 26077 5436 26100
rect 5474 26077 5500 26100
rect 5500 26077 5508 26100
rect 5546 26077 5568 26100
rect 5568 26077 5580 26100
rect 5618 26077 5636 26100
rect 5636 26077 5652 26100
rect 5690 26077 5704 26100
rect 5704 26077 5724 26100
rect 5762 26077 5772 26100
rect 5772 26077 5796 26100
rect 5834 26077 5840 26100
rect 5840 26077 5868 26100
rect 5906 26077 5908 26100
rect 5908 26077 5940 26100
rect 5978 26077 6010 26100
rect 6010 26077 6012 26100
rect 6050 26077 6078 26100
rect 6078 26077 6084 26100
rect 6122 26077 6146 26100
rect 6146 26077 6156 26100
rect 6194 26077 6214 26100
rect 6214 26077 6228 26100
rect 6266 26077 6282 26100
rect 6282 26077 6300 26100
rect 6338 26077 6350 26100
rect 6350 26077 6372 26100
rect 6410 26077 6418 26100
rect 6418 26077 6444 26100
rect 6482 26077 6486 26100
rect 6486 26077 6516 26100
rect 6554 26077 6588 26111
rect 6626 26100 6660 26111
rect 6698 26100 6732 26111
rect 6770 26100 6804 26111
rect 6842 26100 6876 26111
rect 6914 26100 6948 26111
rect 6986 26100 7020 26111
rect 7058 26100 7092 26111
rect 7130 26100 7164 26111
rect 7202 26100 7236 26111
rect 7274 26100 7308 26111
rect 7346 26100 7380 26111
rect 7418 26100 7452 26111
rect 7490 26100 7524 26111
rect 7562 26100 7596 26111
rect 7634 26100 7668 26111
rect 7706 26100 7740 26111
rect 6626 26077 6656 26100
rect 6656 26077 6660 26100
rect 6698 26077 6724 26100
rect 6724 26077 6732 26100
rect 6770 26077 6792 26100
rect 6792 26077 6804 26100
rect 6842 26077 6860 26100
rect 6860 26077 6876 26100
rect 6914 26077 6928 26100
rect 6928 26077 6948 26100
rect 6986 26077 6996 26100
rect 6996 26077 7020 26100
rect 7058 26077 7064 26100
rect 7064 26077 7092 26100
rect 7130 26077 7132 26100
rect 7132 26077 7164 26100
rect 7202 26077 7234 26100
rect 7234 26077 7236 26100
rect 7274 26077 7302 26100
rect 7302 26077 7308 26100
rect 7346 26077 7370 26100
rect 7370 26077 7380 26100
rect 7418 26077 7438 26100
rect 7438 26077 7452 26100
rect 7490 26077 7506 26100
rect 7506 26077 7524 26100
rect 7562 26077 7574 26100
rect 7574 26077 7596 26100
rect 7634 26077 7642 26100
rect 7642 26077 7668 26100
rect 7706 26077 7710 26100
rect 7710 26077 7740 26100
rect 7778 26077 7812 26111
rect 7850 26100 7884 26111
rect 7922 26100 7956 26111
rect 7994 26100 8028 26111
rect 8066 26100 8100 26111
rect 8138 26100 8172 26111
rect 8210 26100 8244 26111
rect 8282 26100 8316 26111
rect 8354 26100 8388 26111
rect 8426 26100 8460 26111
rect 8498 26100 8532 26111
rect 8570 26100 8604 26111
rect 8642 26100 8676 26111
rect 8714 26100 8748 26111
rect 8786 26100 8820 26111
rect 8858 26100 8892 26111
rect 8930 26100 8964 26111
rect 7850 26077 7880 26100
rect 7880 26077 7884 26100
rect 7922 26077 7948 26100
rect 7948 26077 7956 26100
rect 7994 26077 8016 26100
rect 8016 26077 8028 26100
rect 8066 26077 8084 26100
rect 8084 26077 8100 26100
rect 8138 26077 8152 26100
rect 8152 26077 8172 26100
rect 8210 26077 8220 26100
rect 8220 26077 8244 26100
rect 8282 26077 8288 26100
rect 8288 26077 8316 26100
rect 8354 26077 8356 26100
rect 8356 26077 8388 26100
rect 8426 26077 8458 26100
rect 8458 26077 8460 26100
rect 8498 26077 8526 26100
rect 8526 26077 8532 26100
rect 8570 26077 8594 26100
rect 8594 26077 8604 26100
rect 8642 26077 8662 26100
rect 8662 26077 8676 26100
rect 8714 26077 8730 26100
rect 8730 26077 8748 26100
rect 8786 26077 8798 26100
rect 8798 26077 8820 26100
rect 8858 26077 8866 26100
rect 8866 26077 8892 26100
rect 8930 26077 8934 26100
rect 8934 26077 8964 26100
rect 9002 26077 9036 26111
rect 9074 26100 9108 26111
rect 9146 26100 9180 26111
rect 9218 26100 9252 26111
rect 9290 26100 9324 26111
rect 9362 26100 9396 26111
rect 9434 26100 9468 26111
rect 9506 26100 9540 26111
rect 9578 26100 9612 26111
rect 9650 26100 9684 26111
rect 9722 26100 9756 26111
rect 9794 26100 9828 26111
rect 9866 26100 9900 26111
rect 9938 26100 9972 26111
rect 10010 26100 10044 26111
rect 10082 26100 10116 26111
rect 10154 26100 10188 26111
rect 9074 26077 9104 26100
rect 9104 26077 9108 26100
rect 9146 26077 9172 26100
rect 9172 26077 9180 26100
rect 9218 26077 9240 26100
rect 9240 26077 9252 26100
rect 9290 26077 9308 26100
rect 9308 26077 9324 26100
rect 9362 26077 9376 26100
rect 9376 26077 9396 26100
rect 9434 26077 9444 26100
rect 9444 26077 9468 26100
rect 9506 26077 9512 26100
rect 9512 26077 9540 26100
rect 9578 26077 9580 26100
rect 9580 26077 9612 26100
rect 9650 26077 9682 26100
rect 9682 26077 9684 26100
rect 9722 26077 9750 26100
rect 9750 26077 9756 26100
rect 9794 26077 9818 26100
rect 9818 26077 9828 26100
rect 9866 26077 9886 26100
rect 9886 26077 9900 26100
rect 9938 26077 9954 26100
rect 9954 26077 9972 26100
rect 10010 26077 10022 26100
rect 10022 26077 10044 26100
rect 10082 26077 10090 26100
rect 10090 26077 10116 26100
rect 10154 26077 10158 26100
rect 10158 26077 10188 26100
rect 10226 26077 10260 26111
rect 10298 26100 10332 26111
rect 10370 26100 10404 26111
rect 10442 26100 10476 26111
rect 10514 26100 10548 26111
rect 10586 26100 10620 26111
rect 10658 26100 10692 26111
rect 10730 26100 10764 26111
rect 10802 26100 10836 26111
rect 10874 26100 10908 26111
rect 10946 26100 10980 26111
rect 11018 26100 11052 26111
rect 11090 26100 11124 26111
rect 11162 26100 11196 26111
rect 11234 26100 11268 26111
rect 11306 26100 11340 26111
rect 11378 26100 11412 26111
rect 10298 26077 10328 26100
rect 10328 26077 10332 26100
rect 10370 26077 10396 26100
rect 10396 26077 10404 26100
rect 10442 26077 10464 26100
rect 10464 26077 10476 26100
rect 10514 26077 10532 26100
rect 10532 26077 10548 26100
rect 10586 26077 10600 26100
rect 10600 26077 10620 26100
rect 10658 26077 10668 26100
rect 10668 26077 10692 26100
rect 10730 26077 10736 26100
rect 10736 26077 10764 26100
rect 10802 26077 10804 26100
rect 10804 26077 10836 26100
rect 10874 26077 10906 26100
rect 10906 26077 10908 26100
rect 10946 26077 10974 26100
rect 10974 26077 10980 26100
rect 11018 26077 11042 26100
rect 11042 26077 11052 26100
rect 11090 26077 11110 26100
rect 11110 26077 11124 26100
rect 11162 26077 11178 26100
rect 11178 26077 11196 26100
rect 11234 26077 11246 26100
rect 11246 26077 11268 26100
rect 11306 26077 11314 26100
rect 11314 26077 11340 26100
rect 11378 26077 11382 26100
rect 11382 26077 11412 26100
rect 11450 26077 11484 26111
rect 11522 26100 11556 26111
rect 11594 26100 11628 26111
rect 11666 26100 11700 26111
rect 11738 26100 11772 26111
rect 11810 26100 11844 26111
rect 11882 26100 11916 26111
rect 11954 26100 11988 26111
rect 12026 26100 12060 26111
rect 12098 26100 12132 26111
rect 12170 26100 12204 26111
rect 12242 26100 12276 26111
rect 12314 26100 12348 26111
rect 12386 26100 12420 26111
rect 12458 26100 12492 26111
rect 12530 26100 12564 26111
rect 12602 26100 12636 26111
rect 11522 26077 11552 26100
rect 11552 26077 11556 26100
rect 11594 26077 11620 26100
rect 11620 26077 11628 26100
rect 11666 26077 11688 26100
rect 11688 26077 11700 26100
rect 11738 26077 11756 26100
rect 11756 26077 11772 26100
rect 11810 26077 11824 26100
rect 11824 26077 11844 26100
rect 11882 26077 11892 26100
rect 11892 26077 11916 26100
rect 11954 26077 11960 26100
rect 11960 26077 11988 26100
rect 12026 26077 12028 26100
rect 12028 26077 12060 26100
rect 12098 26077 12130 26100
rect 12130 26077 12132 26100
rect 12170 26077 12198 26100
rect 12198 26077 12204 26100
rect 12242 26077 12266 26100
rect 12266 26077 12276 26100
rect 12314 26077 12334 26100
rect 12334 26077 12348 26100
rect 12386 26077 12402 26100
rect 12402 26077 12420 26100
rect 12458 26077 12470 26100
rect 12470 26077 12492 26100
rect 12530 26077 12538 26100
rect 12538 26077 12564 26100
rect 12602 26077 12606 26100
rect 12606 26077 12636 26100
rect 12674 26077 12708 26111
rect 12746 26100 12780 26111
rect 12818 26100 12852 26111
rect 12890 26100 12924 26111
rect 12962 26100 12996 26111
rect 13034 26100 13068 26111
rect 13106 26100 13140 26111
rect 13178 26100 13212 26111
rect 13250 26100 13284 26111
rect 13322 26100 13356 26111
rect 13394 26100 13428 26111
rect 13466 26100 13500 26111
rect 13538 26100 13572 26111
rect 13610 26100 13644 26111
rect 13682 26100 13716 26111
rect 13754 26100 13788 26111
rect 13826 26100 13860 26111
rect 12746 26077 12776 26100
rect 12776 26077 12780 26100
rect 12818 26077 12844 26100
rect 12844 26077 12852 26100
rect 12890 26077 12912 26100
rect 12912 26077 12924 26100
rect 12962 26077 12980 26100
rect 12980 26077 12996 26100
rect 13034 26077 13048 26100
rect 13048 26077 13068 26100
rect 13106 26077 13116 26100
rect 13116 26077 13140 26100
rect 13178 26077 13184 26100
rect 13184 26077 13212 26100
rect 13250 26077 13252 26100
rect 13252 26077 13284 26100
rect 13322 26077 13354 26100
rect 13354 26077 13356 26100
rect 13394 26077 13422 26100
rect 13422 26077 13428 26100
rect 13466 26077 13490 26100
rect 13490 26077 13500 26100
rect 13538 26077 13558 26100
rect 13558 26077 13572 26100
rect 13610 26077 13626 26100
rect 13626 26077 13644 26100
rect 13682 26077 13694 26100
rect 13694 26077 13716 26100
rect 13754 26077 13762 26100
rect 13762 26077 13788 26100
rect 13826 26077 13830 26100
rect 13830 26077 13860 26100
rect 13898 26077 13932 26111
rect 13970 26100 14004 26111
rect 14042 26100 14076 26111
rect 14114 26100 14148 26111
rect 14186 26100 14220 26111
rect 14258 26100 14292 26111
rect 14330 26100 14364 26111
rect 14402 26100 14436 26111
rect 14474 26100 14508 26111
rect 14546 26100 14580 26111
rect 14618 26100 14652 26111
rect 14690 26100 14724 26111
rect 13970 26077 14000 26100
rect 14000 26077 14004 26100
rect 14042 26077 14068 26100
rect 14068 26077 14076 26100
rect 14114 26077 14136 26100
rect 14136 26077 14148 26100
rect 14186 26077 14204 26100
rect 14204 26077 14220 26100
rect 14258 26077 14272 26100
rect 14272 26077 14292 26100
rect 14330 26077 14340 26100
rect 14340 26077 14364 26100
rect 14402 26077 14408 26100
rect 14408 26077 14436 26100
rect 14474 26077 14476 26100
rect 14476 26077 14508 26100
rect 14546 26077 14578 26100
rect 14578 26077 14580 26100
rect 14618 26077 14646 26100
rect 14646 26077 14652 26100
rect 14690 26077 14714 26100
rect 14714 26077 14724 26100
rect 243 26028 277 26037
rect 316 26028 350 26037
rect 389 26028 423 26037
rect 462 26028 496 26037
rect 535 26028 569 26037
rect 608 26028 642 26037
rect 681 26028 715 26037
rect 754 26028 788 26037
rect 827 26028 861 26037
rect 900 26028 934 26037
rect 973 26028 1007 26037
rect 1046 26028 1080 26037
rect 1119 26028 1153 26037
rect 1192 26028 1226 26037
rect 1265 26028 1299 26037
rect 1338 26028 1372 26037
rect 1411 26028 1445 26037
rect 243 26003 276 26028
rect 276 26003 277 26028
rect 316 26003 345 26028
rect 345 26003 350 26028
rect 389 26003 414 26028
rect 414 26003 423 26028
rect 462 26003 483 26028
rect 483 26003 496 26028
rect 535 26003 552 26028
rect 552 26003 569 26028
rect 608 26003 621 26028
rect 621 26003 642 26028
rect 681 26003 690 26028
rect 690 26003 715 26028
rect 754 26003 759 26028
rect 759 26003 788 26028
rect 827 26003 828 26028
rect 828 26003 861 26028
rect 900 26003 931 26028
rect 931 26003 934 26028
rect 973 26003 1000 26028
rect 1000 26003 1007 26028
rect 1046 26003 1069 26028
rect 1069 26003 1080 26028
rect 1119 26003 1138 26028
rect 1138 26003 1153 26028
rect 1192 26003 1207 26028
rect 1207 26003 1226 26028
rect 1265 26003 1276 26028
rect 1276 26003 1299 26028
rect 1338 26003 1345 26028
rect 1345 26003 1372 26028
rect 1411 26003 1414 26028
rect 1414 26003 1445 26028
rect 1484 26003 1518 26037
rect 1557 26028 1591 26037
rect 1630 26028 1664 26037
rect 1703 26028 1737 26037
rect 1776 26028 1810 26037
rect 1849 26028 1883 26037
rect 1922 26028 1956 26037
rect 1995 26028 2029 26037
rect 2068 26028 2102 26037
rect 2141 26028 2175 26037
rect 2214 26028 2248 26037
rect 2287 26028 2321 26037
rect 2360 26028 2394 26037
rect 2433 26028 2467 26037
rect 2506 26028 2540 26037
rect 2579 26028 2613 26037
rect 2652 26028 2686 26037
rect 1557 26003 1587 26028
rect 1587 26003 1591 26028
rect 1630 26003 1656 26028
rect 1656 26003 1664 26028
rect 1703 26003 1725 26028
rect 1725 26003 1737 26028
rect 1776 26003 1794 26028
rect 1794 26003 1810 26028
rect 1849 26003 1863 26028
rect 1863 26003 1883 26028
rect 1922 26003 1932 26028
rect 1932 26003 1956 26028
rect 1995 26003 2001 26028
rect 2001 26003 2029 26028
rect 2068 26003 2070 26028
rect 2070 26003 2102 26028
rect 2141 26003 2173 26028
rect 2173 26003 2175 26028
rect 2214 26003 2242 26028
rect 2242 26003 2248 26028
rect 2287 26003 2311 26028
rect 2311 26003 2321 26028
rect 2360 26003 2380 26028
rect 2380 26003 2394 26028
rect 2433 26003 2449 26028
rect 2449 26003 2467 26028
rect 2506 26003 2518 26028
rect 2518 26003 2540 26028
rect 2579 26003 2587 26028
rect 2587 26003 2613 26028
rect 2652 26003 2656 26028
rect 2656 26003 2686 26028
rect 2725 26003 2759 26037
rect 2798 26028 2832 26037
rect 2871 26028 2905 26037
rect 2944 26028 2978 26037
rect 3017 26028 3051 26037
rect 3090 26028 3124 26037
rect 3163 26028 3197 26037
rect 3236 26028 3270 26037
rect 3309 26028 3343 26037
rect 3382 26028 3416 26037
rect 3455 26028 3489 26037
rect 3528 26028 3562 26037
rect 3601 26028 3635 26037
rect 3674 26028 3708 26037
rect 3746 26028 3780 26037
rect 3818 26028 3852 26037
rect 3890 26028 3924 26037
rect 3962 26028 3996 26037
rect 4034 26028 4068 26037
rect 2798 26003 2829 26028
rect 2829 26003 2832 26028
rect 2871 26003 2898 26028
rect 2898 26003 2905 26028
rect 2944 26003 2967 26028
rect 2967 26003 2978 26028
rect 3017 26003 3036 26028
rect 3036 26003 3051 26028
rect 3090 26003 3105 26028
rect 3105 26003 3124 26028
rect 3163 26003 3174 26028
rect 3174 26003 3197 26028
rect 3236 26003 3243 26028
rect 3243 26003 3270 26028
rect 3309 26003 3312 26028
rect 3312 26003 3343 26028
rect 3382 26003 3415 26028
rect 3415 26003 3416 26028
rect 3455 26003 3484 26028
rect 3484 26003 3489 26028
rect 3528 26003 3553 26028
rect 3553 26003 3562 26028
rect 3601 26003 3622 26028
rect 3622 26003 3635 26028
rect 3674 26003 3691 26028
rect 3691 26003 3708 26028
rect 3746 26003 3760 26028
rect 3760 26003 3780 26028
rect 3818 26003 3829 26028
rect 3829 26003 3852 26028
rect 3890 26003 3898 26028
rect 3898 26003 3924 26028
rect 3962 26003 3967 26028
rect 3967 26003 3996 26028
rect 4034 26003 4036 26028
rect 4036 26003 4068 26028
rect 4106 26003 4140 26037
rect 4178 26028 4212 26037
rect 4250 26028 4284 26037
rect 4322 26028 4356 26037
rect 4394 26028 4428 26037
rect 4466 26028 4500 26037
rect 4538 26028 4572 26037
rect 4610 26028 4644 26037
rect 4682 26028 4716 26037
rect 4754 26028 4788 26037
rect 4826 26028 4860 26037
rect 4898 26028 4932 26037
rect 4970 26028 5004 26037
rect 5042 26028 5076 26037
rect 5114 26028 5148 26037
rect 5186 26028 5220 26037
rect 5258 26028 5292 26037
rect 4178 26003 4208 26028
rect 4208 26003 4212 26028
rect 4250 26003 4276 26028
rect 4276 26003 4284 26028
rect 4322 26003 4344 26028
rect 4344 26003 4356 26028
rect 4394 26003 4412 26028
rect 4412 26003 4428 26028
rect 4466 26003 4480 26028
rect 4480 26003 4500 26028
rect 4538 26003 4548 26028
rect 4548 26003 4572 26028
rect 4610 26003 4616 26028
rect 4616 26003 4644 26028
rect 4682 26003 4684 26028
rect 4684 26003 4716 26028
rect 4754 26003 4786 26028
rect 4786 26003 4788 26028
rect 4826 26003 4854 26028
rect 4854 26003 4860 26028
rect 4898 26003 4922 26028
rect 4922 26003 4932 26028
rect 4970 26003 4990 26028
rect 4990 26003 5004 26028
rect 5042 26003 5058 26028
rect 5058 26003 5076 26028
rect 5114 26003 5126 26028
rect 5126 26003 5148 26028
rect 5186 26003 5194 26028
rect 5194 26003 5220 26028
rect 5258 26003 5262 26028
rect 5262 26003 5292 26028
rect 5330 26003 5364 26037
rect 5402 26028 5436 26037
rect 5474 26028 5508 26037
rect 5546 26028 5580 26037
rect 5618 26028 5652 26037
rect 5690 26028 5724 26037
rect 5762 26028 5796 26037
rect 5834 26028 5868 26037
rect 5906 26028 5940 26037
rect 5978 26028 6012 26037
rect 6050 26028 6084 26037
rect 6122 26028 6156 26037
rect 6194 26028 6228 26037
rect 6266 26028 6300 26037
rect 6338 26028 6372 26037
rect 6410 26028 6444 26037
rect 6482 26028 6516 26037
rect 5402 26003 5432 26028
rect 5432 26003 5436 26028
rect 5474 26003 5500 26028
rect 5500 26003 5508 26028
rect 5546 26003 5568 26028
rect 5568 26003 5580 26028
rect 5618 26003 5636 26028
rect 5636 26003 5652 26028
rect 5690 26003 5704 26028
rect 5704 26003 5724 26028
rect 5762 26003 5772 26028
rect 5772 26003 5796 26028
rect 5834 26003 5840 26028
rect 5840 26003 5868 26028
rect 5906 26003 5908 26028
rect 5908 26003 5940 26028
rect 5978 26003 6010 26028
rect 6010 26003 6012 26028
rect 6050 26003 6078 26028
rect 6078 26003 6084 26028
rect 6122 26003 6146 26028
rect 6146 26003 6156 26028
rect 6194 26003 6214 26028
rect 6214 26003 6228 26028
rect 6266 26003 6282 26028
rect 6282 26003 6300 26028
rect 6338 26003 6350 26028
rect 6350 26003 6372 26028
rect 6410 26003 6418 26028
rect 6418 26003 6444 26028
rect 6482 26003 6486 26028
rect 6486 26003 6516 26028
rect 6554 26003 6588 26037
rect 6626 26028 6660 26037
rect 6698 26028 6732 26037
rect 6770 26028 6804 26037
rect 6842 26028 6876 26037
rect 6914 26028 6948 26037
rect 6986 26028 7020 26037
rect 7058 26028 7092 26037
rect 7130 26028 7164 26037
rect 7202 26028 7236 26037
rect 7274 26028 7308 26037
rect 7346 26028 7380 26037
rect 7418 26028 7452 26037
rect 7490 26028 7524 26037
rect 7562 26028 7596 26037
rect 7634 26028 7668 26037
rect 7706 26028 7740 26037
rect 6626 26003 6656 26028
rect 6656 26003 6660 26028
rect 6698 26003 6724 26028
rect 6724 26003 6732 26028
rect 6770 26003 6792 26028
rect 6792 26003 6804 26028
rect 6842 26003 6860 26028
rect 6860 26003 6876 26028
rect 6914 26003 6928 26028
rect 6928 26003 6948 26028
rect 6986 26003 6996 26028
rect 6996 26003 7020 26028
rect 7058 26003 7064 26028
rect 7064 26003 7092 26028
rect 7130 26003 7132 26028
rect 7132 26003 7164 26028
rect 7202 26003 7234 26028
rect 7234 26003 7236 26028
rect 7274 26003 7302 26028
rect 7302 26003 7308 26028
rect 7346 26003 7370 26028
rect 7370 26003 7380 26028
rect 7418 26003 7438 26028
rect 7438 26003 7452 26028
rect 7490 26003 7506 26028
rect 7506 26003 7524 26028
rect 7562 26003 7574 26028
rect 7574 26003 7596 26028
rect 7634 26003 7642 26028
rect 7642 26003 7668 26028
rect 7706 26003 7710 26028
rect 7710 26003 7740 26028
rect 7778 26003 7812 26037
rect 7850 26028 7884 26037
rect 7922 26028 7956 26037
rect 7994 26028 8028 26037
rect 8066 26028 8100 26037
rect 8138 26028 8172 26037
rect 8210 26028 8244 26037
rect 8282 26028 8316 26037
rect 8354 26028 8388 26037
rect 8426 26028 8460 26037
rect 8498 26028 8532 26037
rect 8570 26028 8604 26037
rect 8642 26028 8676 26037
rect 8714 26028 8748 26037
rect 8786 26028 8820 26037
rect 8858 26028 8892 26037
rect 8930 26028 8964 26037
rect 7850 26003 7880 26028
rect 7880 26003 7884 26028
rect 7922 26003 7948 26028
rect 7948 26003 7956 26028
rect 7994 26003 8016 26028
rect 8016 26003 8028 26028
rect 8066 26003 8084 26028
rect 8084 26003 8100 26028
rect 8138 26003 8152 26028
rect 8152 26003 8172 26028
rect 8210 26003 8220 26028
rect 8220 26003 8244 26028
rect 8282 26003 8288 26028
rect 8288 26003 8316 26028
rect 8354 26003 8356 26028
rect 8356 26003 8388 26028
rect 8426 26003 8458 26028
rect 8458 26003 8460 26028
rect 8498 26003 8526 26028
rect 8526 26003 8532 26028
rect 8570 26003 8594 26028
rect 8594 26003 8604 26028
rect 8642 26003 8662 26028
rect 8662 26003 8676 26028
rect 8714 26003 8730 26028
rect 8730 26003 8748 26028
rect 8786 26003 8798 26028
rect 8798 26003 8820 26028
rect 8858 26003 8866 26028
rect 8866 26003 8892 26028
rect 8930 26003 8934 26028
rect 8934 26003 8964 26028
rect 9002 26003 9036 26037
rect 9074 26028 9108 26037
rect 9146 26028 9180 26037
rect 9218 26028 9252 26037
rect 9290 26028 9324 26037
rect 9362 26028 9396 26037
rect 9434 26028 9468 26037
rect 9506 26028 9540 26037
rect 9578 26028 9612 26037
rect 9650 26028 9684 26037
rect 9722 26028 9756 26037
rect 9794 26028 9828 26037
rect 9866 26028 9900 26037
rect 9938 26028 9972 26037
rect 10010 26028 10044 26037
rect 10082 26028 10116 26037
rect 10154 26028 10188 26037
rect 9074 26003 9104 26028
rect 9104 26003 9108 26028
rect 9146 26003 9172 26028
rect 9172 26003 9180 26028
rect 9218 26003 9240 26028
rect 9240 26003 9252 26028
rect 9290 26003 9308 26028
rect 9308 26003 9324 26028
rect 9362 26003 9376 26028
rect 9376 26003 9396 26028
rect 9434 26003 9444 26028
rect 9444 26003 9468 26028
rect 9506 26003 9512 26028
rect 9512 26003 9540 26028
rect 9578 26003 9580 26028
rect 9580 26003 9612 26028
rect 9650 26003 9682 26028
rect 9682 26003 9684 26028
rect 9722 26003 9750 26028
rect 9750 26003 9756 26028
rect 9794 26003 9818 26028
rect 9818 26003 9828 26028
rect 9866 26003 9886 26028
rect 9886 26003 9900 26028
rect 9938 26003 9954 26028
rect 9954 26003 9972 26028
rect 10010 26003 10022 26028
rect 10022 26003 10044 26028
rect 10082 26003 10090 26028
rect 10090 26003 10116 26028
rect 10154 26003 10158 26028
rect 10158 26003 10188 26028
rect 10226 26003 10260 26037
rect 10298 26028 10332 26037
rect 10370 26028 10404 26037
rect 10442 26028 10476 26037
rect 10514 26028 10548 26037
rect 10586 26028 10620 26037
rect 10658 26028 10692 26037
rect 10730 26028 10764 26037
rect 10802 26028 10836 26037
rect 10874 26028 10908 26037
rect 10946 26028 10980 26037
rect 11018 26028 11052 26037
rect 11090 26028 11124 26037
rect 11162 26028 11196 26037
rect 11234 26028 11268 26037
rect 11306 26028 11340 26037
rect 11378 26028 11412 26037
rect 10298 26003 10328 26028
rect 10328 26003 10332 26028
rect 10370 26003 10396 26028
rect 10396 26003 10404 26028
rect 10442 26003 10464 26028
rect 10464 26003 10476 26028
rect 10514 26003 10532 26028
rect 10532 26003 10548 26028
rect 10586 26003 10600 26028
rect 10600 26003 10620 26028
rect 10658 26003 10668 26028
rect 10668 26003 10692 26028
rect 10730 26003 10736 26028
rect 10736 26003 10764 26028
rect 10802 26003 10804 26028
rect 10804 26003 10836 26028
rect 10874 26003 10906 26028
rect 10906 26003 10908 26028
rect 10946 26003 10974 26028
rect 10974 26003 10980 26028
rect 11018 26003 11042 26028
rect 11042 26003 11052 26028
rect 11090 26003 11110 26028
rect 11110 26003 11124 26028
rect 11162 26003 11178 26028
rect 11178 26003 11196 26028
rect 11234 26003 11246 26028
rect 11246 26003 11268 26028
rect 11306 26003 11314 26028
rect 11314 26003 11340 26028
rect 11378 26003 11382 26028
rect 11382 26003 11412 26028
rect 11450 26003 11484 26037
rect 11522 26028 11556 26037
rect 11594 26028 11628 26037
rect 11666 26028 11700 26037
rect 11738 26028 11772 26037
rect 11810 26028 11844 26037
rect 11882 26028 11916 26037
rect 11954 26028 11988 26037
rect 12026 26028 12060 26037
rect 12098 26028 12132 26037
rect 12170 26028 12204 26037
rect 12242 26028 12276 26037
rect 12314 26028 12348 26037
rect 12386 26028 12420 26037
rect 12458 26028 12492 26037
rect 12530 26028 12564 26037
rect 12602 26028 12636 26037
rect 11522 26003 11552 26028
rect 11552 26003 11556 26028
rect 11594 26003 11620 26028
rect 11620 26003 11628 26028
rect 11666 26003 11688 26028
rect 11688 26003 11700 26028
rect 11738 26003 11756 26028
rect 11756 26003 11772 26028
rect 11810 26003 11824 26028
rect 11824 26003 11844 26028
rect 11882 26003 11892 26028
rect 11892 26003 11916 26028
rect 11954 26003 11960 26028
rect 11960 26003 11988 26028
rect 12026 26003 12028 26028
rect 12028 26003 12060 26028
rect 12098 26003 12130 26028
rect 12130 26003 12132 26028
rect 12170 26003 12198 26028
rect 12198 26003 12204 26028
rect 12242 26003 12266 26028
rect 12266 26003 12276 26028
rect 12314 26003 12334 26028
rect 12334 26003 12348 26028
rect 12386 26003 12402 26028
rect 12402 26003 12420 26028
rect 12458 26003 12470 26028
rect 12470 26003 12492 26028
rect 12530 26003 12538 26028
rect 12538 26003 12564 26028
rect 12602 26003 12606 26028
rect 12606 26003 12636 26028
rect 12674 26003 12708 26037
rect 12746 26028 12780 26037
rect 12818 26028 12852 26037
rect 12890 26028 12924 26037
rect 12962 26028 12996 26037
rect 13034 26028 13068 26037
rect 13106 26028 13140 26037
rect 13178 26028 13212 26037
rect 13250 26028 13284 26037
rect 13322 26028 13356 26037
rect 13394 26028 13428 26037
rect 13466 26028 13500 26037
rect 13538 26028 13572 26037
rect 13610 26028 13644 26037
rect 13682 26028 13716 26037
rect 13754 26028 13788 26037
rect 13826 26028 13860 26037
rect 12746 26003 12776 26028
rect 12776 26003 12780 26028
rect 12818 26003 12844 26028
rect 12844 26003 12852 26028
rect 12890 26003 12912 26028
rect 12912 26003 12924 26028
rect 12962 26003 12980 26028
rect 12980 26003 12996 26028
rect 13034 26003 13048 26028
rect 13048 26003 13068 26028
rect 13106 26003 13116 26028
rect 13116 26003 13140 26028
rect 13178 26003 13184 26028
rect 13184 26003 13212 26028
rect 13250 26003 13252 26028
rect 13252 26003 13284 26028
rect 13322 26003 13354 26028
rect 13354 26003 13356 26028
rect 13394 26003 13422 26028
rect 13422 26003 13428 26028
rect 13466 26003 13490 26028
rect 13490 26003 13500 26028
rect 13538 26003 13558 26028
rect 13558 26003 13572 26028
rect 13610 26003 13626 26028
rect 13626 26003 13644 26028
rect 13682 26003 13694 26028
rect 13694 26003 13716 26028
rect 13754 26003 13762 26028
rect 13762 26003 13788 26028
rect 13826 26003 13830 26028
rect 13830 26003 13860 26028
rect 13898 26003 13932 26037
rect 13970 26028 14004 26037
rect 14042 26028 14076 26037
rect 14114 26028 14148 26037
rect 14186 26028 14220 26037
rect 14258 26028 14292 26037
rect 14330 26028 14364 26037
rect 14402 26028 14436 26037
rect 14474 26028 14508 26037
rect 14546 26028 14580 26037
rect 14618 26028 14652 26037
rect 14690 26028 14724 26037
rect 13970 26003 14000 26028
rect 14000 26003 14004 26028
rect 14042 26003 14068 26028
rect 14068 26003 14076 26028
rect 14114 26003 14136 26028
rect 14136 26003 14148 26028
rect 14186 26003 14204 26028
rect 14204 26003 14220 26028
rect 14258 26003 14272 26028
rect 14272 26003 14292 26028
rect 14330 26003 14340 26028
rect 14340 26003 14364 26028
rect 14402 26003 14408 26028
rect 14408 26003 14436 26028
rect 14474 26003 14476 26028
rect 14476 26003 14508 26028
rect 14546 26003 14578 26028
rect 14578 26003 14580 26028
rect 14618 26003 14646 26028
rect 14646 26003 14652 26028
rect 14690 26003 14714 26028
rect 14714 26003 14724 26028
rect 243 25956 277 25963
rect 316 25956 350 25963
rect 389 25956 423 25963
rect 462 25956 496 25963
rect 535 25956 569 25963
rect 608 25956 642 25963
rect 681 25956 715 25963
rect 754 25956 788 25963
rect 827 25956 861 25963
rect 900 25956 934 25963
rect 973 25956 1007 25963
rect 1046 25956 1080 25963
rect 1119 25956 1153 25963
rect 1192 25956 1226 25963
rect 1265 25956 1299 25963
rect 1338 25956 1372 25963
rect 1411 25956 1445 25963
rect 243 25929 276 25956
rect 276 25929 277 25956
rect 316 25929 345 25956
rect 345 25929 350 25956
rect 389 25929 414 25956
rect 414 25929 423 25956
rect 462 25929 483 25956
rect 483 25929 496 25956
rect 535 25929 552 25956
rect 552 25929 569 25956
rect 608 25929 621 25956
rect 621 25929 642 25956
rect 681 25929 690 25956
rect 690 25929 715 25956
rect 754 25929 759 25956
rect 759 25929 788 25956
rect 827 25929 828 25956
rect 828 25929 861 25956
rect 900 25929 931 25956
rect 931 25929 934 25956
rect 973 25929 1000 25956
rect 1000 25929 1007 25956
rect 1046 25929 1069 25956
rect 1069 25929 1080 25956
rect 1119 25929 1138 25956
rect 1138 25929 1153 25956
rect 1192 25929 1207 25956
rect 1207 25929 1226 25956
rect 1265 25929 1276 25956
rect 1276 25929 1299 25956
rect 1338 25929 1345 25956
rect 1345 25929 1372 25956
rect 1411 25929 1414 25956
rect 1414 25929 1445 25956
rect 1484 25929 1518 25963
rect 1557 25956 1591 25963
rect 1630 25956 1664 25963
rect 1703 25956 1737 25963
rect 1776 25956 1810 25963
rect 1849 25956 1883 25963
rect 1922 25956 1956 25963
rect 1995 25956 2029 25963
rect 2068 25956 2102 25963
rect 2141 25956 2175 25963
rect 2214 25956 2248 25963
rect 2287 25956 2321 25963
rect 2360 25956 2394 25963
rect 2433 25956 2467 25963
rect 2506 25956 2540 25963
rect 2579 25956 2613 25963
rect 2652 25956 2686 25963
rect 1557 25929 1587 25956
rect 1587 25929 1591 25956
rect 1630 25929 1656 25956
rect 1656 25929 1664 25956
rect 1703 25929 1725 25956
rect 1725 25929 1737 25956
rect 1776 25929 1794 25956
rect 1794 25929 1810 25956
rect 1849 25929 1863 25956
rect 1863 25929 1883 25956
rect 1922 25929 1932 25956
rect 1932 25929 1956 25956
rect 1995 25929 2001 25956
rect 2001 25929 2029 25956
rect 2068 25929 2070 25956
rect 2070 25929 2102 25956
rect 2141 25929 2173 25956
rect 2173 25929 2175 25956
rect 2214 25929 2242 25956
rect 2242 25929 2248 25956
rect 2287 25929 2311 25956
rect 2311 25929 2321 25956
rect 2360 25929 2380 25956
rect 2380 25929 2394 25956
rect 2433 25929 2449 25956
rect 2449 25929 2467 25956
rect 2506 25929 2518 25956
rect 2518 25929 2540 25956
rect 2579 25929 2587 25956
rect 2587 25929 2613 25956
rect 2652 25929 2656 25956
rect 2656 25929 2686 25956
rect 2725 25929 2759 25963
rect 2798 25956 2832 25963
rect 2871 25956 2905 25963
rect 2944 25956 2978 25963
rect 3017 25956 3051 25963
rect 3090 25956 3124 25963
rect 3163 25956 3197 25963
rect 3236 25956 3270 25963
rect 3309 25956 3343 25963
rect 3382 25956 3416 25963
rect 3455 25956 3489 25963
rect 3528 25956 3562 25963
rect 3601 25956 3635 25963
rect 3674 25956 3708 25963
rect 3746 25956 3780 25963
rect 3818 25956 3852 25963
rect 3890 25956 3924 25963
rect 3962 25956 3996 25963
rect 4034 25956 4068 25963
rect 2798 25929 2829 25956
rect 2829 25929 2832 25956
rect 2871 25929 2898 25956
rect 2898 25929 2905 25956
rect 2944 25929 2967 25956
rect 2967 25929 2978 25956
rect 3017 25929 3036 25956
rect 3036 25929 3051 25956
rect 3090 25929 3105 25956
rect 3105 25929 3124 25956
rect 3163 25929 3174 25956
rect 3174 25929 3197 25956
rect 3236 25929 3243 25956
rect 3243 25929 3270 25956
rect 3309 25929 3312 25956
rect 3312 25929 3343 25956
rect 3382 25929 3415 25956
rect 3415 25929 3416 25956
rect 3455 25929 3484 25956
rect 3484 25929 3489 25956
rect 3528 25929 3553 25956
rect 3553 25929 3562 25956
rect 3601 25929 3622 25956
rect 3622 25929 3635 25956
rect 3674 25929 3691 25956
rect 3691 25929 3708 25956
rect 3746 25929 3760 25956
rect 3760 25929 3780 25956
rect 3818 25929 3829 25956
rect 3829 25929 3852 25956
rect 3890 25929 3898 25956
rect 3898 25929 3924 25956
rect 3962 25929 3967 25956
rect 3967 25929 3996 25956
rect 4034 25929 4036 25956
rect 4036 25929 4068 25956
rect 4106 25929 4140 25963
rect 4178 25956 4212 25963
rect 4250 25956 4284 25963
rect 4322 25956 4356 25963
rect 4394 25956 4428 25963
rect 4466 25956 4500 25963
rect 4538 25956 4572 25963
rect 4610 25956 4644 25963
rect 4682 25956 4716 25963
rect 4754 25956 4788 25963
rect 4826 25956 4860 25963
rect 4898 25956 4932 25963
rect 4970 25956 5004 25963
rect 5042 25956 5076 25963
rect 5114 25956 5148 25963
rect 5186 25956 5220 25963
rect 5258 25956 5292 25963
rect 4178 25929 4208 25956
rect 4208 25929 4212 25956
rect 4250 25929 4276 25956
rect 4276 25929 4284 25956
rect 4322 25929 4344 25956
rect 4344 25929 4356 25956
rect 4394 25929 4412 25956
rect 4412 25929 4428 25956
rect 4466 25929 4480 25956
rect 4480 25929 4500 25956
rect 4538 25929 4548 25956
rect 4548 25929 4572 25956
rect 4610 25929 4616 25956
rect 4616 25929 4644 25956
rect 4682 25929 4684 25956
rect 4684 25929 4716 25956
rect 4754 25929 4786 25956
rect 4786 25929 4788 25956
rect 4826 25929 4854 25956
rect 4854 25929 4860 25956
rect 4898 25929 4922 25956
rect 4922 25929 4932 25956
rect 4970 25929 4990 25956
rect 4990 25929 5004 25956
rect 5042 25929 5058 25956
rect 5058 25929 5076 25956
rect 5114 25929 5126 25956
rect 5126 25929 5148 25956
rect 5186 25929 5194 25956
rect 5194 25929 5220 25956
rect 5258 25929 5262 25956
rect 5262 25929 5292 25956
rect 5330 25929 5364 25963
rect 5402 25956 5436 25963
rect 5474 25956 5508 25963
rect 5546 25956 5580 25963
rect 5618 25956 5652 25963
rect 5690 25956 5724 25963
rect 5762 25956 5796 25963
rect 5834 25956 5868 25963
rect 5906 25956 5940 25963
rect 5978 25956 6012 25963
rect 6050 25956 6084 25963
rect 6122 25956 6156 25963
rect 6194 25956 6228 25963
rect 6266 25956 6300 25963
rect 6338 25956 6372 25963
rect 6410 25956 6444 25963
rect 6482 25956 6516 25963
rect 5402 25929 5432 25956
rect 5432 25929 5436 25956
rect 5474 25929 5500 25956
rect 5500 25929 5508 25956
rect 5546 25929 5568 25956
rect 5568 25929 5580 25956
rect 5618 25929 5636 25956
rect 5636 25929 5652 25956
rect 5690 25929 5704 25956
rect 5704 25929 5724 25956
rect 5762 25929 5772 25956
rect 5772 25929 5796 25956
rect 5834 25929 5840 25956
rect 5840 25929 5868 25956
rect 5906 25929 5908 25956
rect 5908 25929 5940 25956
rect 5978 25929 6010 25956
rect 6010 25929 6012 25956
rect 6050 25929 6078 25956
rect 6078 25929 6084 25956
rect 6122 25929 6146 25956
rect 6146 25929 6156 25956
rect 6194 25929 6214 25956
rect 6214 25929 6228 25956
rect 6266 25929 6282 25956
rect 6282 25929 6300 25956
rect 6338 25929 6350 25956
rect 6350 25929 6372 25956
rect 6410 25929 6418 25956
rect 6418 25929 6444 25956
rect 6482 25929 6486 25956
rect 6486 25929 6516 25956
rect 6554 25929 6588 25963
rect 6626 25956 6660 25963
rect 6698 25956 6732 25963
rect 6770 25956 6804 25963
rect 6842 25956 6876 25963
rect 6914 25956 6948 25963
rect 6986 25956 7020 25963
rect 7058 25956 7092 25963
rect 7130 25956 7164 25963
rect 7202 25956 7236 25963
rect 7274 25956 7308 25963
rect 7346 25956 7380 25963
rect 7418 25956 7452 25963
rect 7490 25956 7524 25963
rect 7562 25956 7596 25963
rect 7634 25956 7668 25963
rect 7706 25956 7740 25963
rect 6626 25929 6656 25956
rect 6656 25929 6660 25956
rect 6698 25929 6724 25956
rect 6724 25929 6732 25956
rect 6770 25929 6792 25956
rect 6792 25929 6804 25956
rect 6842 25929 6860 25956
rect 6860 25929 6876 25956
rect 6914 25929 6928 25956
rect 6928 25929 6948 25956
rect 6986 25929 6996 25956
rect 6996 25929 7020 25956
rect 7058 25929 7064 25956
rect 7064 25929 7092 25956
rect 7130 25929 7132 25956
rect 7132 25929 7164 25956
rect 7202 25929 7234 25956
rect 7234 25929 7236 25956
rect 7274 25929 7302 25956
rect 7302 25929 7308 25956
rect 7346 25929 7370 25956
rect 7370 25929 7380 25956
rect 7418 25929 7438 25956
rect 7438 25929 7452 25956
rect 7490 25929 7506 25956
rect 7506 25929 7524 25956
rect 7562 25929 7574 25956
rect 7574 25929 7596 25956
rect 7634 25929 7642 25956
rect 7642 25929 7668 25956
rect 7706 25929 7710 25956
rect 7710 25929 7740 25956
rect 7778 25929 7812 25963
rect 7850 25956 7884 25963
rect 7922 25956 7956 25963
rect 7994 25956 8028 25963
rect 8066 25956 8100 25963
rect 8138 25956 8172 25963
rect 8210 25956 8244 25963
rect 8282 25956 8316 25963
rect 8354 25956 8388 25963
rect 8426 25956 8460 25963
rect 8498 25956 8532 25963
rect 8570 25956 8604 25963
rect 8642 25956 8676 25963
rect 8714 25956 8748 25963
rect 8786 25956 8820 25963
rect 8858 25956 8892 25963
rect 8930 25956 8964 25963
rect 7850 25929 7880 25956
rect 7880 25929 7884 25956
rect 7922 25929 7948 25956
rect 7948 25929 7956 25956
rect 7994 25929 8016 25956
rect 8016 25929 8028 25956
rect 8066 25929 8084 25956
rect 8084 25929 8100 25956
rect 8138 25929 8152 25956
rect 8152 25929 8172 25956
rect 8210 25929 8220 25956
rect 8220 25929 8244 25956
rect 8282 25929 8288 25956
rect 8288 25929 8316 25956
rect 8354 25929 8356 25956
rect 8356 25929 8388 25956
rect 8426 25929 8458 25956
rect 8458 25929 8460 25956
rect 8498 25929 8526 25956
rect 8526 25929 8532 25956
rect 8570 25929 8594 25956
rect 8594 25929 8604 25956
rect 8642 25929 8662 25956
rect 8662 25929 8676 25956
rect 8714 25929 8730 25956
rect 8730 25929 8748 25956
rect 8786 25929 8798 25956
rect 8798 25929 8820 25956
rect 8858 25929 8866 25956
rect 8866 25929 8892 25956
rect 8930 25929 8934 25956
rect 8934 25929 8964 25956
rect 9002 25929 9036 25963
rect 9074 25956 9108 25963
rect 9146 25956 9180 25963
rect 9218 25956 9252 25963
rect 9290 25956 9324 25963
rect 9362 25956 9396 25963
rect 9434 25956 9468 25963
rect 9506 25956 9540 25963
rect 9578 25956 9612 25963
rect 9650 25956 9684 25963
rect 9722 25956 9756 25963
rect 9794 25956 9828 25963
rect 9866 25956 9900 25963
rect 9938 25956 9972 25963
rect 10010 25956 10044 25963
rect 10082 25956 10116 25963
rect 10154 25956 10188 25963
rect 9074 25929 9104 25956
rect 9104 25929 9108 25956
rect 9146 25929 9172 25956
rect 9172 25929 9180 25956
rect 9218 25929 9240 25956
rect 9240 25929 9252 25956
rect 9290 25929 9308 25956
rect 9308 25929 9324 25956
rect 9362 25929 9376 25956
rect 9376 25929 9396 25956
rect 9434 25929 9444 25956
rect 9444 25929 9468 25956
rect 9506 25929 9512 25956
rect 9512 25929 9540 25956
rect 9578 25929 9580 25956
rect 9580 25929 9612 25956
rect 9650 25929 9682 25956
rect 9682 25929 9684 25956
rect 9722 25929 9750 25956
rect 9750 25929 9756 25956
rect 9794 25929 9818 25956
rect 9818 25929 9828 25956
rect 9866 25929 9886 25956
rect 9886 25929 9900 25956
rect 9938 25929 9954 25956
rect 9954 25929 9972 25956
rect 10010 25929 10022 25956
rect 10022 25929 10044 25956
rect 10082 25929 10090 25956
rect 10090 25929 10116 25956
rect 10154 25929 10158 25956
rect 10158 25929 10188 25956
rect 10226 25929 10260 25963
rect 10298 25956 10332 25963
rect 10370 25956 10404 25963
rect 10442 25956 10476 25963
rect 10514 25956 10548 25963
rect 10586 25956 10620 25963
rect 10658 25956 10692 25963
rect 10730 25956 10764 25963
rect 10802 25956 10836 25963
rect 10874 25956 10908 25963
rect 10946 25956 10980 25963
rect 11018 25956 11052 25963
rect 11090 25956 11124 25963
rect 11162 25956 11196 25963
rect 11234 25956 11268 25963
rect 11306 25956 11340 25963
rect 11378 25956 11412 25963
rect 10298 25929 10328 25956
rect 10328 25929 10332 25956
rect 10370 25929 10396 25956
rect 10396 25929 10404 25956
rect 10442 25929 10464 25956
rect 10464 25929 10476 25956
rect 10514 25929 10532 25956
rect 10532 25929 10548 25956
rect 10586 25929 10600 25956
rect 10600 25929 10620 25956
rect 10658 25929 10668 25956
rect 10668 25929 10692 25956
rect 10730 25929 10736 25956
rect 10736 25929 10764 25956
rect 10802 25929 10804 25956
rect 10804 25929 10836 25956
rect 10874 25929 10906 25956
rect 10906 25929 10908 25956
rect 10946 25929 10974 25956
rect 10974 25929 10980 25956
rect 11018 25929 11042 25956
rect 11042 25929 11052 25956
rect 11090 25929 11110 25956
rect 11110 25929 11124 25956
rect 11162 25929 11178 25956
rect 11178 25929 11196 25956
rect 11234 25929 11246 25956
rect 11246 25929 11268 25956
rect 11306 25929 11314 25956
rect 11314 25929 11340 25956
rect 11378 25929 11382 25956
rect 11382 25929 11412 25956
rect 11450 25929 11484 25963
rect 11522 25956 11556 25963
rect 11594 25956 11628 25963
rect 11666 25956 11700 25963
rect 11738 25956 11772 25963
rect 11810 25956 11844 25963
rect 11882 25956 11916 25963
rect 11954 25956 11988 25963
rect 12026 25956 12060 25963
rect 12098 25956 12132 25963
rect 12170 25956 12204 25963
rect 12242 25956 12276 25963
rect 12314 25956 12348 25963
rect 12386 25956 12420 25963
rect 12458 25956 12492 25963
rect 12530 25956 12564 25963
rect 12602 25956 12636 25963
rect 11522 25929 11552 25956
rect 11552 25929 11556 25956
rect 11594 25929 11620 25956
rect 11620 25929 11628 25956
rect 11666 25929 11688 25956
rect 11688 25929 11700 25956
rect 11738 25929 11756 25956
rect 11756 25929 11772 25956
rect 11810 25929 11824 25956
rect 11824 25929 11844 25956
rect 11882 25929 11892 25956
rect 11892 25929 11916 25956
rect 11954 25929 11960 25956
rect 11960 25929 11988 25956
rect 12026 25929 12028 25956
rect 12028 25929 12060 25956
rect 12098 25929 12130 25956
rect 12130 25929 12132 25956
rect 12170 25929 12198 25956
rect 12198 25929 12204 25956
rect 12242 25929 12266 25956
rect 12266 25929 12276 25956
rect 12314 25929 12334 25956
rect 12334 25929 12348 25956
rect 12386 25929 12402 25956
rect 12402 25929 12420 25956
rect 12458 25929 12470 25956
rect 12470 25929 12492 25956
rect 12530 25929 12538 25956
rect 12538 25929 12564 25956
rect 12602 25929 12606 25956
rect 12606 25929 12636 25956
rect 12674 25929 12708 25963
rect 12746 25956 12780 25963
rect 12818 25956 12852 25963
rect 12890 25956 12924 25963
rect 12962 25956 12996 25963
rect 13034 25956 13068 25963
rect 13106 25956 13140 25963
rect 13178 25956 13212 25963
rect 13250 25956 13284 25963
rect 13322 25956 13356 25963
rect 13394 25956 13428 25963
rect 13466 25956 13500 25963
rect 13538 25956 13572 25963
rect 13610 25956 13644 25963
rect 13682 25956 13716 25963
rect 13754 25956 13788 25963
rect 13826 25956 13860 25963
rect 12746 25929 12776 25956
rect 12776 25929 12780 25956
rect 12818 25929 12844 25956
rect 12844 25929 12852 25956
rect 12890 25929 12912 25956
rect 12912 25929 12924 25956
rect 12962 25929 12980 25956
rect 12980 25929 12996 25956
rect 13034 25929 13048 25956
rect 13048 25929 13068 25956
rect 13106 25929 13116 25956
rect 13116 25929 13140 25956
rect 13178 25929 13184 25956
rect 13184 25929 13212 25956
rect 13250 25929 13252 25956
rect 13252 25929 13284 25956
rect 13322 25929 13354 25956
rect 13354 25929 13356 25956
rect 13394 25929 13422 25956
rect 13422 25929 13428 25956
rect 13466 25929 13490 25956
rect 13490 25929 13500 25956
rect 13538 25929 13558 25956
rect 13558 25929 13572 25956
rect 13610 25929 13626 25956
rect 13626 25929 13644 25956
rect 13682 25929 13694 25956
rect 13694 25929 13716 25956
rect 13754 25929 13762 25956
rect 13762 25929 13788 25956
rect 13826 25929 13830 25956
rect 13830 25929 13860 25956
rect 13898 25929 13932 25963
rect 13970 25956 14004 25963
rect 14042 25956 14076 25963
rect 14114 25956 14148 25963
rect 14186 25956 14220 25963
rect 14258 25956 14292 25963
rect 14330 25956 14364 25963
rect 14402 25956 14436 25963
rect 14474 25956 14508 25963
rect 14546 25956 14580 25963
rect 14618 25956 14652 25963
rect 14690 25956 14724 25963
rect 13970 25929 14000 25956
rect 14000 25929 14004 25956
rect 14042 25929 14068 25956
rect 14068 25929 14076 25956
rect 14114 25929 14136 25956
rect 14136 25929 14148 25956
rect 14186 25929 14204 25956
rect 14204 25929 14220 25956
rect 14258 25929 14272 25956
rect 14272 25929 14292 25956
rect 14330 25929 14340 25956
rect 14340 25929 14364 25956
rect 14402 25929 14408 25956
rect 14408 25929 14436 25956
rect 14474 25929 14476 25956
rect 14476 25929 14508 25956
rect 14546 25929 14578 25956
rect 14578 25929 14580 25956
rect 14618 25929 14646 25956
rect 14646 25929 14652 25956
rect 14690 25929 14714 25956
rect 14714 25929 14724 25956
rect 243 25884 277 25889
rect 316 25884 350 25889
rect 389 25884 423 25889
rect 462 25884 496 25889
rect 535 25884 569 25889
rect 608 25884 642 25889
rect 681 25884 715 25889
rect 754 25884 788 25889
rect 827 25884 861 25889
rect 900 25884 934 25889
rect 973 25884 1007 25889
rect 1046 25884 1080 25889
rect 1119 25884 1153 25889
rect 1192 25884 1226 25889
rect 1265 25884 1299 25889
rect 1338 25884 1372 25889
rect 1411 25884 1445 25889
rect 243 25855 276 25884
rect 276 25855 277 25884
rect 316 25855 345 25884
rect 345 25855 350 25884
rect 389 25855 414 25884
rect 414 25855 423 25884
rect 462 25855 483 25884
rect 483 25855 496 25884
rect 535 25855 552 25884
rect 552 25855 569 25884
rect 608 25855 621 25884
rect 621 25855 642 25884
rect 681 25855 690 25884
rect 690 25855 715 25884
rect 754 25855 759 25884
rect 759 25855 788 25884
rect 827 25855 828 25884
rect 828 25855 861 25884
rect 900 25855 931 25884
rect 931 25855 934 25884
rect 973 25855 1000 25884
rect 1000 25855 1007 25884
rect 1046 25855 1069 25884
rect 1069 25855 1080 25884
rect 1119 25855 1138 25884
rect 1138 25855 1153 25884
rect 1192 25855 1207 25884
rect 1207 25855 1226 25884
rect 1265 25855 1276 25884
rect 1276 25855 1299 25884
rect 1338 25855 1345 25884
rect 1345 25855 1372 25884
rect 1411 25855 1414 25884
rect 1414 25855 1445 25884
rect 1484 25855 1518 25889
rect 1557 25884 1591 25889
rect 1630 25884 1664 25889
rect 1703 25884 1737 25889
rect 1776 25884 1810 25889
rect 1849 25884 1883 25889
rect 1922 25884 1956 25889
rect 1995 25884 2029 25889
rect 2068 25884 2102 25889
rect 2141 25884 2175 25889
rect 2214 25884 2248 25889
rect 2287 25884 2321 25889
rect 2360 25884 2394 25889
rect 2433 25884 2467 25889
rect 2506 25884 2540 25889
rect 2579 25884 2613 25889
rect 2652 25884 2686 25889
rect 1557 25855 1587 25884
rect 1587 25855 1591 25884
rect 1630 25855 1656 25884
rect 1656 25855 1664 25884
rect 1703 25855 1725 25884
rect 1725 25855 1737 25884
rect 1776 25855 1794 25884
rect 1794 25855 1810 25884
rect 1849 25855 1863 25884
rect 1863 25855 1883 25884
rect 1922 25855 1932 25884
rect 1932 25855 1956 25884
rect 1995 25855 2001 25884
rect 2001 25855 2029 25884
rect 2068 25855 2070 25884
rect 2070 25855 2102 25884
rect 2141 25855 2173 25884
rect 2173 25855 2175 25884
rect 2214 25855 2242 25884
rect 2242 25855 2248 25884
rect 2287 25855 2311 25884
rect 2311 25855 2321 25884
rect 2360 25855 2380 25884
rect 2380 25855 2394 25884
rect 2433 25855 2449 25884
rect 2449 25855 2467 25884
rect 2506 25855 2518 25884
rect 2518 25855 2540 25884
rect 2579 25855 2587 25884
rect 2587 25855 2613 25884
rect 2652 25855 2656 25884
rect 2656 25855 2686 25884
rect 2725 25855 2759 25889
rect 2798 25884 2832 25889
rect 2871 25884 2905 25889
rect 2944 25884 2978 25889
rect 3017 25884 3051 25889
rect 3090 25884 3124 25889
rect 3163 25884 3197 25889
rect 3236 25884 3270 25889
rect 3309 25884 3343 25889
rect 3382 25884 3416 25889
rect 3455 25884 3489 25889
rect 3528 25884 3562 25889
rect 3601 25884 3635 25889
rect 3674 25884 3708 25889
rect 3746 25884 3780 25889
rect 3818 25884 3852 25889
rect 3890 25884 3924 25889
rect 3962 25884 3996 25889
rect 4034 25884 4068 25889
rect 2798 25855 2829 25884
rect 2829 25855 2832 25884
rect 2871 25855 2898 25884
rect 2898 25855 2905 25884
rect 2944 25855 2967 25884
rect 2967 25855 2978 25884
rect 3017 25855 3036 25884
rect 3036 25855 3051 25884
rect 3090 25855 3105 25884
rect 3105 25855 3124 25884
rect 3163 25855 3174 25884
rect 3174 25855 3197 25884
rect 3236 25855 3243 25884
rect 3243 25855 3270 25884
rect 3309 25855 3312 25884
rect 3312 25855 3343 25884
rect 3382 25855 3415 25884
rect 3415 25855 3416 25884
rect 3455 25855 3484 25884
rect 3484 25855 3489 25884
rect 3528 25855 3553 25884
rect 3553 25855 3562 25884
rect 3601 25855 3622 25884
rect 3622 25855 3635 25884
rect 3674 25855 3691 25884
rect 3691 25855 3708 25884
rect 3746 25855 3760 25884
rect 3760 25855 3780 25884
rect 3818 25855 3829 25884
rect 3829 25855 3852 25884
rect 3890 25855 3898 25884
rect 3898 25855 3924 25884
rect 3962 25855 3967 25884
rect 3967 25855 3996 25884
rect 4034 25855 4036 25884
rect 4036 25855 4068 25884
rect 4106 25855 4140 25889
rect 4178 25884 4212 25889
rect 4250 25884 4284 25889
rect 4322 25884 4356 25889
rect 4394 25884 4428 25889
rect 4466 25884 4500 25889
rect 4538 25884 4572 25889
rect 4610 25884 4644 25889
rect 4682 25884 4716 25889
rect 4754 25884 4788 25889
rect 4826 25884 4860 25889
rect 4898 25884 4932 25889
rect 4970 25884 5004 25889
rect 5042 25884 5076 25889
rect 5114 25884 5148 25889
rect 5186 25884 5220 25889
rect 5258 25884 5292 25889
rect 4178 25855 4208 25884
rect 4208 25855 4212 25884
rect 4250 25855 4276 25884
rect 4276 25855 4284 25884
rect 4322 25855 4344 25884
rect 4344 25855 4356 25884
rect 4394 25855 4412 25884
rect 4412 25855 4428 25884
rect 4466 25855 4480 25884
rect 4480 25855 4500 25884
rect 4538 25855 4548 25884
rect 4548 25855 4572 25884
rect 4610 25855 4616 25884
rect 4616 25855 4644 25884
rect 4682 25855 4684 25884
rect 4684 25855 4716 25884
rect 4754 25855 4786 25884
rect 4786 25855 4788 25884
rect 4826 25855 4854 25884
rect 4854 25855 4860 25884
rect 4898 25855 4922 25884
rect 4922 25855 4932 25884
rect 4970 25855 4990 25884
rect 4990 25855 5004 25884
rect 5042 25855 5058 25884
rect 5058 25855 5076 25884
rect 5114 25855 5126 25884
rect 5126 25855 5148 25884
rect 5186 25855 5194 25884
rect 5194 25855 5220 25884
rect 5258 25855 5262 25884
rect 5262 25855 5292 25884
rect 5330 25855 5364 25889
rect 5402 25884 5436 25889
rect 5474 25884 5508 25889
rect 5546 25884 5580 25889
rect 5618 25884 5652 25889
rect 5690 25884 5724 25889
rect 5762 25884 5796 25889
rect 5834 25884 5868 25889
rect 5906 25884 5940 25889
rect 5978 25884 6012 25889
rect 6050 25884 6084 25889
rect 6122 25884 6156 25889
rect 6194 25884 6228 25889
rect 6266 25884 6300 25889
rect 6338 25884 6372 25889
rect 6410 25884 6444 25889
rect 6482 25884 6516 25889
rect 5402 25855 5432 25884
rect 5432 25855 5436 25884
rect 5474 25855 5500 25884
rect 5500 25855 5508 25884
rect 5546 25855 5568 25884
rect 5568 25855 5580 25884
rect 5618 25855 5636 25884
rect 5636 25855 5652 25884
rect 5690 25855 5704 25884
rect 5704 25855 5724 25884
rect 5762 25855 5772 25884
rect 5772 25855 5796 25884
rect 5834 25855 5840 25884
rect 5840 25855 5868 25884
rect 5906 25855 5908 25884
rect 5908 25855 5940 25884
rect 5978 25855 6010 25884
rect 6010 25855 6012 25884
rect 6050 25855 6078 25884
rect 6078 25855 6084 25884
rect 6122 25855 6146 25884
rect 6146 25855 6156 25884
rect 6194 25855 6214 25884
rect 6214 25855 6228 25884
rect 6266 25855 6282 25884
rect 6282 25855 6300 25884
rect 6338 25855 6350 25884
rect 6350 25855 6372 25884
rect 6410 25855 6418 25884
rect 6418 25855 6444 25884
rect 6482 25855 6486 25884
rect 6486 25855 6516 25884
rect 6554 25855 6588 25889
rect 6626 25884 6660 25889
rect 6698 25884 6732 25889
rect 6770 25884 6804 25889
rect 6842 25884 6876 25889
rect 6914 25884 6948 25889
rect 6986 25884 7020 25889
rect 7058 25884 7092 25889
rect 7130 25884 7164 25889
rect 7202 25884 7236 25889
rect 7274 25884 7308 25889
rect 7346 25884 7380 25889
rect 7418 25884 7452 25889
rect 7490 25884 7524 25889
rect 7562 25884 7596 25889
rect 7634 25884 7668 25889
rect 7706 25884 7740 25889
rect 6626 25855 6656 25884
rect 6656 25855 6660 25884
rect 6698 25855 6724 25884
rect 6724 25855 6732 25884
rect 6770 25855 6792 25884
rect 6792 25855 6804 25884
rect 6842 25855 6860 25884
rect 6860 25855 6876 25884
rect 6914 25855 6928 25884
rect 6928 25855 6948 25884
rect 6986 25855 6996 25884
rect 6996 25855 7020 25884
rect 7058 25855 7064 25884
rect 7064 25855 7092 25884
rect 7130 25855 7132 25884
rect 7132 25855 7164 25884
rect 7202 25855 7234 25884
rect 7234 25855 7236 25884
rect 7274 25855 7302 25884
rect 7302 25855 7308 25884
rect 7346 25855 7370 25884
rect 7370 25855 7380 25884
rect 7418 25855 7438 25884
rect 7438 25855 7452 25884
rect 7490 25855 7506 25884
rect 7506 25855 7524 25884
rect 7562 25855 7574 25884
rect 7574 25855 7596 25884
rect 7634 25855 7642 25884
rect 7642 25855 7668 25884
rect 7706 25855 7710 25884
rect 7710 25855 7740 25884
rect 7778 25855 7812 25889
rect 7850 25884 7884 25889
rect 7922 25884 7956 25889
rect 7994 25884 8028 25889
rect 8066 25884 8100 25889
rect 8138 25884 8172 25889
rect 8210 25884 8244 25889
rect 8282 25884 8316 25889
rect 8354 25884 8388 25889
rect 8426 25884 8460 25889
rect 8498 25884 8532 25889
rect 8570 25884 8604 25889
rect 8642 25884 8676 25889
rect 8714 25884 8748 25889
rect 8786 25884 8820 25889
rect 8858 25884 8892 25889
rect 8930 25884 8964 25889
rect 7850 25855 7880 25884
rect 7880 25855 7884 25884
rect 7922 25855 7948 25884
rect 7948 25855 7956 25884
rect 7994 25855 8016 25884
rect 8016 25855 8028 25884
rect 8066 25855 8084 25884
rect 8084 25855 8100 25884
rect 8138 25855 8152 25884
rect 8152 25855 8172 25884
rect 8210 25855 8220 25884
rect 8220 25855 8244 25884
rect 8282 25855 8288 25884
rect 8288 25855 8316 25884
rect 8354 25855 8356 25884
rect 8356 25855 8388 25884
rect 8426 25855 8458 25884
rect 8458 25855 8460 25884
rect 8498 25855 8526 25884
rect 8526 25855 8532 25884
rect 8570 25855 8594 25884
rect 8594 25855 8604 25884
rect 8642 25855 8662 25884
rect 8662 25855 8676 25884
rect 8714 25855 8730 25884
rect 8730 25855 8748 25884
rect 8786 25855 8798 25884
rect 8798 25855 8820 25884
rect 8858 25855 8866 25884
rect 8866 25855 8892 25884
rect 8930 25855 8934 25884
rect 8934 25855 8964 25884
rect 9002 25855 9036 25889
rect 9074 25884 9108 25889
rect 9146 25884 9180 25889
rect 9218 25884 9252 25889
rect 9290 25884 9324 25889
rect 9362 25884 9396 25889
rect 9434 25884 9468 25889
rect 9506 25884 9540 25889
rect 9578 25884 9612 25889
rect 9650 25884 9684 25889
rect 9722 25884 9756 25889
rect 9794 25884 9828 25889
rect 9866 25884 9900 25889
rect 9938 25884 9972 25889
rect 10010 25884 10044 25889
rect 10082 25884 10116 25889
rect 10154 25884 10188 25889
rect 9074 25855 9104 25884
rect 9104 25855 9108 25884
rect 9146 25855 9172 25884
rect 9172 25855 9180 25884
rect 9218 25855 9240 25884
rect 9240 25855 9252 25884
rect 9290 25855 9308 25884
rect 9308 25855 9324 25884
rect 9362 25855 9376 25884
rect 9376 25855 9396 25884
rect 9434 25855 9444 25884
rect 9444 25855 9468 25884
rect 9506 25855 9512 25884
rect 9512 25855 9540 25884
rect 9578 25855 9580 25884
rect 9580 25855 9612 25884
rect 9650 25855 9682 25884
rect 9682 25855 9684 25884
rect 9722 25855 9750 25884
rect 9750 25855 9756 25884
rect 9794 25855 9818 25884
rect 9818 25855 9828 25884
rect 9866 25855 9886 25884
rect 9886 25855 9900 25884
rect 9938 25855 9954 25884
rect 9954 25855 9972 25884
rect 10010 25855 10022 25884
rect 10022 25855 10044 25884
rect 10082 25855 10090 25884
rect 10090 25855 10116 25884
rect 10154 25855 10158 25884
rect 10158 25855 10188 25884
rect 10226 25855 10260 25889
rect 10298 25884 10332 25889
rect 10370 25884 10404 25889
rect 10442 25884 10476 25889
rect 10514 25884 10548 25889
rect 10586 25884 10620 25889
rect 10658 25884 10692 25889
rect 10730 25884 10764 25889
rect 10802 25884 10836 25889
rect 10874 25884 10908 25889
rect 10946 25884 10980 25889
rect 11018 25884 11052 25889
rect 11090 25884 11124 25889
rect 11162 25884 11196 25889
rect 11234 25884 11268 25889
rect 11306 25884 11340 25889
rect 11378 25884 11412 25889
rect 10298 25855 10328 25884
rect 10328 25855 10332 25884
rect 10370 25855 10396 25884
rect 10396 25855 10404 25884
rect 10442 25855 10464 25884
rect 10464 25855 10476 25884
rect 10514 25855 10532 25884
rect 10532 25855 10548 25884
rect 10586 25855 10600 25884
rect 10600 25855 10620 25884
rect 10658 25855 10668 25884
rect 10668 25855 10692 25884
rect 10730 25855 10736 25884
rect 10736 25855 10764 25884
rect 10802 25855 10804 25884
rect 10804 25855 10836 25884
rect 10874 25855 10906 25884
rect 10906 25855 10908 25884
rect 10946 25855 10974 25884
rect 10974 25855 10980 25884
rect 11018 25855 11042 25884
rect 11042 25855 11052 25884
rect 11090 25855 11110 25884
rect 11110 25855 11124 25884
rect 11162 25855 11178 25884
rect 11178 25855 11196 25884
rect 11234 25855 11246 25884
rect 11246 25855 11268 25884
rect 11306 25855 11314 25884
rect 11314 25855 11340 25884
rect 11378 25855 11382 25884
rect 11382 25855 11412 25884
rect 11450 25855 11484 25889
rect 11522 25884 11556 25889
rect 11594 25884 11628 25889
rect 11666 25884 11700 25889
rect 11738 25884 11772 25889
rect 11810 25884 11844 25889
rect 11882 25884 11916 25889
rect 11954 25884 11988 25889
rect 12026 25884 12060 25889
rect 12098 25884 12132 25889
rect 12170 25884 12204 25889
rect 12242 25884 12276 25889
rect 12314 25884 12348 25889
rect 12386 25884 12420 25889
rect 12458 25884 12492 25889
rect 12530 25884 12564 25889
rect 12602 25884 12636 25889
rect 11522 25855 11552 25884
rect 11552 25855 11556 25884
rect 11594 25855 11620 25884
rect 11620 25855 11628 25884
rect 11666 25855 11688 25884
rect 11688 25855 11700 25884
rect 11738 25855 11756 25884
rect 11756 25855 11772 25884
rect 11810 25855 11824 25884
rect 11824 25855 11844 25884
rect 11882 25855 11892 25884
rect 11892 25855 11916 25884
rect 11954 25855 11960 25884
rect 11960 25855 11988 25884
rect 12026 25855 12028 25884
rect 12028 25855 12060 25884
rect 12098 25855 12130 25884
rect 12130 25855 12132 25884
rect 12170 25855 12198 25884
rect 12198 25855 12204 25884
rect 12242 25855 12266 25884
rect 12266 25855 12276 25884
rect 12314 25855 12334 25884
rect 12334 25855 12348 25884
rect 12386 25855 12402 25884
rect 12402 25855 12420 25884
rect 12458 25855 12470 25884
rect 12470 25855 12492 25884
rect 12530 25855 12538 25884
rect 12538 25855 12564 25884
rect 12602 25855 12606 25884
rect 12606 25855 12636 25884
rect 12674 25855 12708 25889
rect 12746 25884 12780 25889
rect 12818 25884 12852 25889
rect 12890 25884 12924 25889
rect 12962 25884 12996 25889
rect 13034 25884 13068 25889
rect 13106 25884 13140 25889
rect 13178 25884 13212 25889
rect 13250 25884 13284 25889
rect 13322 25884 13356 25889
rect 13394 25884 13428 25889
rect 13466 25884 13500 25889
rect 13538 25884 13572 25889
rect 13610 25884 13644 25889
rect 13682 25884 13716 25889
rect 13754 25884 13788 25889
rect 13826 25884 13860 25889
rect 12746 25855 12776 25884
rect 12776 25855 12780 25884
rect 12818 25855 12844 25884
rect 12844 25855 12852 25884
rect 12890 25855 12912 25884
rect 12912 25855 12924 25884
rect 12962 25855 12980 25884
rect 12980 25855 12996 25884
rect 13034 25855 13048 25884
rect 13048 25855 13068 25884
rect 13106 25855 13116 25884
rect 13116 25855 13140 25884
rect 13178 25855 13184 25884
rect 13184 25855 13212 25884
rect 13250 25855 13252 25884
rect 13252 25855 13284 25884
rect 13322 25855 13354 25884
rect 13354 25855 13356 25884
rect 13394 25855 13422 25884
rect 13422 25855 13428 25884
rect 13466 25855 13490 25884
rect 13490 25855 13500 25884
rect 13538 25855 13558 25884
rect 13558 25855 13572 25884
rect 13610 25855 13626 25884
rect 13626 25855 13644 25884
rect 13682 25855 13694 25884
rect 13694 25855 13716 25884
rect 13754 25855 13762 25884
rect 13762 25855 13788 25884
rect 13826 25855 13830 25884
rect 13830 25855 13860 25884
rect 13898 25855 13932 25889
rect 13970 25884 14004 25889
rect 14042 25884 14076 25889
rect 14114 25884 14148 25889
rect 14186 25884 14220 25889
rect 14258 25884 14292 25889
rect 14330 25884 14364 25889
rect 14402 25884 14436 25889
rect 14474 25884 14508 25889
rect 14546 25884 14580 25889
rect 14618 25884 14652 25889
rect 14690 25884 14724 25889
rect 13970 25855 14000 25884
rect 14000 25855 14004 25884
rect 14042 25855 14068 25884
rect 14068 25855 14076 25884
rect 14114 25855 14136 25884
rect 14136 25855 14148 25884
rect 14186 25855 14204 25884
rect 14204 25855 14220 25884
rect 14258 25855 14272 25884
rect 14272 25855 14292 25884
rect 14330 25855 14340 25884
rect 14340 25855 14364 25884
rect 14402 25855 14408 25884
rect 14408 25855 14436 25884
rect 14474 25855 14476 25884
rect 14476 25855 14508 25884
rect 14546 25855 14578 25884
rect 14578 25855 14580 25884
rect 14618 25855 14646 25884
rect 14646 25855 14652 25884
rect 14690 25855 14714 25884
rect 14714 25855 14724 25884
rect 243 25812 277 25815
rect 316 25812 350 25815
rect 389 25812 423 25815
rect 462 25812 496 25815
rect 535 25812 569 25815
rect 608 25812 642 25815
rect 681 25812 715 25815
rect 754 25812 788 25815
rect 827 25812 861 25815
rect 900 25812 934 25815
rect 973 25812 1007 25815
rect 1046 25812 1080 25815
rect 1119 25812 1153 25815
rect 1192 25812 1226 25815
rect 1265 25812 1299 25815
rect 1338 25812 1372 25815
rect 1411 25812 1445 25815
rect 243 25781 276 25812
rect 276 25781 277 25812
rect 316 25781 345 25812
rect 345 25781 350 25812
rect 389 25781 414 25812
rect 414 25781 423 25812
rect 462 25781 483 25812
rect 483 25781 496 25812
rect 535 25781 552 25812
rect 552 25781 569 25812
rect 608 25781 621 25812
rect 621 25781 642 25812
rect 681 25781 690 25812
rect 690 25781 715 25812
rect 754 25781 759 25812
rect 759 25781 788 25812
rect 827 25781 828 25812
rect 828 25781 861 25812
rect 900 25781 931 25812
rect 931 25781 934 25812
rect 973 25781 1000 25812
rect 1000 25781 1007 25812
rect 1046 25781 1069 25812
rect 1069 25781 1080 25812
rect 1119 25781 1138 25812
rect 1138 25781 1153 25812
rect 1192 25781 1207 25812
rect 1207 25781 1226 25812
rect 1265 25781 1276 25812
rect 1276 25781 1299 25812
rect 1338 25781 1345 25812
rect 1345 25781 1372 25812
rect 1411 25781 1414 25812
rect 1414 25781 1445 25812
rect 1484 25781 1518 25815
rect 1557 25812 1591 25815
rect 1630 25812 1664 25815
rect 1703 25812 1737 25815
rect 1776 25812 1810 25815
rect 1849 25812 1883 25815
rect 1922 25812 1956 25815
rect 1995 25812 2029 25815
rect 2068 25812 2102 25815
rect 2141 25812 2175 25815
rect 2214 25812 2248 25815
rect 2287 25812 2321 25815
rect 2360 25812 2394 25815
rect 2433 25812 2467 25815
rect 2506 25812 2540 25815
rect 2579 25812 2613 25815
rect 2652 25812 2686 25815
rect 1557 25781 1587 25812
rect 1587 25781 1591 25812
rect 1630 25781 1656 25812
rect 1656 25781 1664 25812
rect 1703 25781 1725 25812
rect 1725 25781 1737 25812
rect 1776 25781 1794 25812
rect 1794 25781 1810 25812
rect 1849 25781 1863 25812
rect 1863 25781 1883 25812
rect 1922 25781 1932 25812
rect 1932 25781 1956 25812
rect 1995 25781 2001 25812
rect 2001 25781 2029 25812
rect 2068 25781 2070 25812
rect 2070 25781 2102 25812
rect 2141 25781 2173 25812
rect 2173 25781 2175 25812
rect 2214 25781 2242 25812
rect 2242 25781 2248 25812
rect 2287 25781 2311 25812
rect 2311 25781 2321 25812
rect 2360 25781 2380 25812
rect 2380 25781 2394 25812
rect 2433 25781 2449 25812
rect 2449 25781 2467 25812
rect 2506 25781 2518 25812
rect 2518 25781 2540 25812
rect 2579 25781 2587 25812
rect 2587 25781 2613 25812
rect 2652 25781 2656 25812
rect 2656 25781 2686 25812
rect 2725 25781 2759 25815
rect 2798 25812 2832 25815
rect 2871 25812 2905 25815
rect 2944 25812 2978 25815
rect 3017 25812 3051 25815
rect 3090 25812 3124 25815
rect 3163 25812 3197 25815
rect 3236 25812 3270 25815
rect 3309 25812 3343 25815
rect 3382 25812 3416 25815
rect 3455 25812 3489 25815
rect 3528 25812 3562 25815
rect 3601 25812 3635 25815
rect 3674 25812 3708 25815
rect 3746 25812 3780 25815
rect 3818 25812 3852 25815
rect 3890 25812 3924 25815
rect 3962 25812 3996 25815
rect 4034 25812 4068 25815
rect 2798 25781 2829 25812
rect 2829 25781 2832 25812
rect 2871 25781 2898 25812
rect 2898 25781 2905 25812
rect 2944 25781 2967 25812
rect 2967 25781 2978 25812
rect 3017 25781 3036 25812
rect 3036 25781 3051 25812
rect 3090 25781 3105 25812
rect 3105 25781 3124 25812
rect 3163 25781 3174 25812
rect 3174 25781 3197 25812
rect 3236 25781 3243 25812
rect 3243 25781 3270 25812
rect 3309 25781 3312 25812
rect 3312 25781 3343 25812
rect 3382 25781 3415 25812
rect 3415 25781 3416 25812
rect 3455 25781 3484 25812
rect 3484 25781 3489 25812
rect 3528 25781 3553 25812
rect 3553 25781 3562 25812
rect 3601 25781 3622 25812
rect 3622 25781 3635 25812
rect 3674 25781 3691 25812
rect 3691 25781 3708 25812
rect 3746 25781 3760 25812
rect 3760 25781 3780 25812
rect 3818 25781 3829 25812
rect 3829 25781 3852 25812
rect 3890 25781 3898 25812
rect 3898 25781 3924 25812
rect 3962 25781 3967 25812
rect 3967 25781 3996 25812
rect 4034 25781 4036 25812
rect 4036 25781 4068 25812
rect 4106 25781 4140 25815
rect 4178 25812 4212 25815
rect 4250 25812 4284 25815
rect 4322 25812 4356 25815
rect 4394 25812 4428 25815
rect 4466 25812 4500 25815
rect 4538 25812 4572 25815
rect 4610 25812 4644 25815
rect 4682 25812 4716 25815
rect 4754 25812 4788 25815
rect 4826 25812 4860 25815
rect 4898 25812 4932 25815
rect 4970 25812 5004 25815
rect 5042 25812 5076 25815
rect 5114 25812 5148 25815
rect 5186 25812 5220 25815
rect 5258 25812 5292 25815
rect 4178 25781 4208 25812
rect 4208 25781 4212 25812
rect 4250 25781 4276 25812
rect 4276 25781 4284 25812
rect 4322 25781 4344 25812
rect 4344 25781 4356 25812
rect 4394 25781 4412 25812
rect 4412 25781 4428 25812
rect 4466 25781 4480 25812
rect 4480 25781 4500 25812
rect 4538 25781 4548 25812
rect 4548 25781 4572 25812
rect 4610 25781 4616 25812
rect 4616 25781 4644 25812
rect 4682 25781 4684 25812
rect 4684 25781 4716 25812
rect 4754 25781 4786 25812
rect 4786 25781 4788 25812
rect 4826 25781 4854 25812
rect 4854 25781 4860 25812
rect 4898 25781 4922 25812
rect 4922 25781 4932 25812
rect 4970 25781 4990 25812
rect 4990 25781 5004 25812
rect 5042 25781 5058 25812
rect 5058 25781 5076 25812
rect 5114 25781 5126 25812
rect 5126 25781 5148 25812
rect 5186 25781 5194 25812
rect 5194 25781 5220 25812
rect 5258 25781 5262 25812
rect 5262 25781 5292 25812
rect 5330 25781 5364 25815
rect 5402 25812 5436 25815
rect 5474 25812 5508 25815
rect 5546 25812 5580 25815
rect 5618 25812 5652 25815
rect 5690 25812 5724 25815
rect 5762 25812 5796 25815
rect 5834 25812 5868 25815
rect 5906 25812 5940 25815
rect 5978 25812 6012 25815
rect 6050 25812 6084 25815
rect 6122 25812 6156 25815
rect 6194 25812 6228 25815
rect 6266 25812 6300 25815
rect 6338 25812 6372 25815
rect 6410 25812 6444 25815
rect 6482 25812 6516 25815
rect 5402 25781 5432 25812
rect 5432 25781 5436 25812
rect 5474 25781 5500 25812
rect 5500 25781 5508 25812
rect 5546 25781 5568 25812
rect 5568 25781 5580 25812
rect 5618 25781 5636 25812
rect 5636 25781 5652 25812
rect 5690 25781 5704 25812
rect 5704 25781 5724 25812
rect 5762 25781 5772 25812
rect 5772 25781 5796 25812
rect 5834 25781 5840 25812
rect 5840 25781 5868 25812
rect 5906 25781 5908 25812
rect 5908 25781 5940 25812
rect 5978 25781 6010 25812
rect 6010 25781 6012 25812
rect 6050 25781 6078 25812
rect 6078 25781 6084 25812
rect 6122 25781 6146 25812
rect 6146 25781 6156 25812
rect 6194 25781 6214 25812
rect 6214 25781 6228 25812
rect 6266 25781 6282 25812
rect 6282 25781 6300 25812
rect 6338 25781 6350 25812
rect 6350 25781 6372 25812
rect 6410 25781 6418 25812
rect 6418 25781 6444 25812
rect 6482 25781 6486 25812
rect 6486 25781 6516 25812
rect 6554 25781 6588 25815
rect 6626 25812 6660 25815
rect 6698 25812 6732 25815
rect 6770 25812 6804 25815
rect 6842 25812 6876 25815
rect 6914 25812 6948 25815
rect 6986 25812 7020 25815
rect 7058 25812 7092 25815
rect 7130 25812 7164 25815
rect 7202 25812 7236 25815
rect 7274 25812 7308 25815
rect 7346 25812 7380 25815
rect 7418 25812 7452 25815
rect 7490 25812 7524 25815
rect 7562 25812 7596 25815
rect 7634 25812 7668 25815
rect 7706 25812 7740 25815
rect 6626 25781 6656 25812
rect 6656 25781 6660 25812
rect 6698 25781 6724 25812
rect 6724 25781 6732 25812
rect 6770 25781 6792 25812
rect 6792 25781 6804 25812
rect 6842 25781 6860 25812
rect 6860 25781 6876 25812
rect 6914 25781 6928 25812
rect 6928 25781 6948 25812
rect 6986 25781 6996 25812
rect 6996 25781 7020 25812
rect 7058 25781 7064 25812
rect 7064 25781 7092 25812
rect 7130 25781 7132 25812
rect 7132 25781 7164 25812
rect 7202 25781 7234 25812
rect 7234 25781 7236 25812
rect 7274 25781 7302 25812
rect 7302 25781 7308 25812
rect 7346 25781 7370 25812
rect 7370 25781 7380 25812
rect 7418 25781 7438 25812
rect 7438 25781 7452 25812
rect 7490 25781 7506 25812
rect 7506 25781 7524 25812
rect 7562 25781 7574 25812
rect 7574 25781 7596 25812
rect 7634 25781 7642 25812
rect 7642 25781 7668 25812
rect 7706 25781 7710 25812
rect 7710 25781 7740 25812
rect 7778 25781 7812 25815
rect 7850 25812 7884 25815
rect 7922 25812 7956 25815
rect 7994 25812 8028 25815
rect 8066 25812 8100 25815
rect 8138 25812 8172 25815
rect 8210 25812 8244 25815
rect 8282 25812 8316 25815
rect 8354 25812 8388 25815
rect 8426 25812 8460 25815
rect 8498 25812 8532 25815
rect 8570 25812 8604 25815
rect 8642 25812 8676 25815
rect 8714 25812 8748 25815
rect 8786 25812 8820 25815
rect 8858 25812 8892 25815
rect 8930 25812 8964 25815
rect 7850 25781 7880 25812
rect 7880 25781 7884 25812
rect 7922 25781 7948 25812
rect 7948 25781 7956 25812
rect 7994 25781 8016 25812
rect 8016 25781 8028 25812
rect 8066 25781 8084 25812
rect 8084 25781 8100 25812
rect 8138 25781 8152 25812
rect 8152 25781 8172 25812
rect 8210 25781 8220 25812
rect 8220 25781 8244 25812
rect 8282 25781 8288 25812
rect 8288 25781 8316 25812
rect 8354 25781 8356 25812
rect 8356 25781 8388 25812
rect 8426 25781 8458 25812
rect 8458 25781 8460 25812
rect 8498 25781 8526 25812
rect 8526 25781 8532 25812
rect 8570 25781 8594 25812
rect 8594 25781 8604 25812
rect 8642 25781 8662 25812
rect 8662 25781 8676 25812
rect 8714 25781 8730 25812
rect 8730 25781 8748 25812
rect 8786 25781 8798 25812
rect 8798 25781 8820 25812
rect 8858 25781 8866 25812
rect 8866 25781 8892 25812
rect 8930 25781 8934 25812
rect 8934 25781 8964 25812
rect 9002 25781 9036 25815
rect 9074 25812 9108 25815
rect 9146 25812 9180 25815
rect 9218 25812 9252 25815
rect 9290 25812 9324 25815
rect 9362 25812 9396 25815
rect 9434 25812 9468 25815
rect 9506 25812 9540 25815
rect 9578 25812 9612 25815
rect 9650 25812 9684 25815
rect 9722 25812 9756 25815
rect 9794 25812 9828 25815
rect 9866 25812 9900 25815
rect 9938 25812 9972 25815
rect 10010 25812 10044 25815
rect 10082 25812 10116 25815
rect 10154 25812 10188 25815
rect 9074 25781 9104 25812
rect 9104 25781 9108 25812
rect 9146 25781 9172 25812
rect 9172 25781 9180 25812
rect 9218 25781 9240 25812
rect 9240 25781 9252 25812
rect 9290 25781 9308 25812
rect 9308 25781 9324 25812
rect 9362 25781 9376 25812
rect 9376 25781 9396 25812
rect 9434 25781 9444 25812
rect 9444 25781 9468 25812
rect 9506 25781 9512 25812
rect 9512 25781 9540 25812
rect 9578 25781 9580 25812
rect 9580 25781 9612 25812
rect 9650 25781 9682 25812
rect 9682 25781 9684 25812
rect 9722 25781 9750 25812
rect 9750 25781 9756 25812
rect 9794 25781 9818 25812
rect 9818 25781 9828 25812
rect 9866 25781 9886 25812
rect 9886 25781 9900 25812
rect 9938 25781 9954 25812
rect 9954 25781 9972 25812
rect 10010 25781 10022 25812
rect 10022 25781 10044 25812
rect 10082 25781 10090 25812
rect 10090 25781 10116 25812
rect 10154 25781 10158 25812
rect 10158 25781 10188 25812
rect 10226 25781 10260 25815
rect 10298 25812 10332 25815
rect 10370 25812 10404 25815
rect 10442 25812 10476 25815
rect 10514 25812 10548 25815
rect 10586 25812 10620 25815
rect 10658 25812 10692 25815
rect 10730 25812 10764 25815
rect 10802 25812 10836 25815
rect 10874 25812 10908 25815
rect 10946 25812 10980 25815
rect 11018 25812 11052 25815
rect 11090 25812 11124 25815
rect 11162 25812 11196 25815
rect 11234 25812 11268 25815
rect 11306 25812 11340 25815
rect 11378 25812 11412 25815
rect 10298 25781 10328 25812
rect 10328 25781 10332 25812
rect 10370 25781 10396 25812
rect 10396 25781 10404 25812
rect 10442 25781 10464 25812
rect 10464 25781 10476 25812
rect 10514 25781 10532 25812
rect 10532 25781 10548 25812
rect 10586 25781 10600 25812
rect 10600 25781 10620 25812
rect 10658 25781 10668 25812
rect 10668 25781 10692 25812
rect 10730 25781 10736 25812
rect 10736 25781 10764 25812
rect 10802 25781 10804 25812
rect 10804 25781 10836 25812
rect 10874 25781 10906 25812
rect 10906 25781 10908 25812
rect 10946 25781 10974 25812
rect 10974 25781 10980 25812
rect 11018 25781 11042 25812
rect 11042 25781 11052 25812
rect 11090 25781 11110 25812
rect 11110 25781 11124 25812
rect 11162 25781 11178 25812
rect 11178 25781 11196 25812
rect 11234 25781 11246 25812
rect 11246 25781 11268 25812
rect 11306 25781 11314 25812
rect 11314 25781 11340 25812
rect 11378 25781 11382 25812
rect 11382 25781 11412 25812
rect 11450 25781 11484 25815
rect 11522 25812 11556 25815
rect 11594 25812 11628 25815
rect 11666 25812 11700 25815
rect 11738 25812 11772 25815
rect 11810 25812 11844 25815
rect 11882 25812 11916 25815
rect 11954 25812 11988 25815
rect 12026 25812 12060 25815
rect 12098 25812 12132 25815
rect 12170 25812 12204 25815
rect 12242 25812 12276 25815
rect 12314 25812 12348 25815
rect 12386 25812 12420 25815
rect 12458 25812 12492 25815
rect 12530 25812 12564 25815
rect 12602 25812 12636 25815
rect 11522 25781 11552 25812
rect 11552 25781 11556 25812
rect 11594 25781 11620 25812
rect 11620 25781 11628 25812
rect 11666 25781 11688 25812
rect 11688 25781 11700 25812
rect 11738 25781 11756 25812
rect 11756 25781 11772 25812
rect 11810 25781 11824 25812
rect 11824 25781 11844 25812
rect 11882 25781 11892 25812
rect 11892 25781 11916 25812
rect 11954 25781 11960 25812
rect 11960 25781 11988 25812
rect 12026 25781 12028 25812
rect 12028 25781 12060 25812
rect 12098 25781 12130 25812
rect 12130 25781 12132 25812
rect 12170 25781 12198 25812
rect 12198 25781 12204 25812
rect 12242 25781 12266 25812
rect 12266 25781 12276 25812
rect 12314 25781 12334 25812
rect 12334 25781 12348 25812
rect 12386 25781 12402 25812
rect 12402 25781 12420 25812
rect 12458 25781 12470 25812
rect 12470 25781 12492 25812
rect 12530 25781 12538 25812
rect 12538 25781 12564 25812
rect 12602 25781 12606 25812
rect 12606 25781 12636 25812
rect 12674 25781 12708 25815
rect 12746 25812 12780 25815
rect 12818 25812 12852 25815
rect 12890 25812 12924 25815
rect 12962 25812 12996 25815
rect 13034 25812 13068 25815
rect 13106 25812 13140 25815
rect 13178 25812 13212 25815
rect 13250 25812 13284 25815
rect 13322 25812 13356 25815
rect 13394 25812 13428 25815
rect 13466 25812 13500 25815
rect 13538 25812 13572 25815
rect 13610 25812 13644 25815
rect 13682 25812 13716 25815
rect 13754 25812 13788 25815
rect 13826 25812 13860 25815
rect 12746 25781 12776 25812
rect 12776 25781 12780 25812
rect 12818 25781 12844 25812
rect 12844 25781 12852 25812
rect 12890 25781 12912 25812
rect 12912 25781 12924 25812
rect 12962 25781 12980 25812
rect 12980 25781 12996 25812
rect 13034 25781 13048 25812
rect 13048 25781 13068 25812
rect 13106 25781 13116 25812
rect 13116 25781 13140 25812
rect 13178 25781 13184 25812
rect 13184 25781 13212 25812
rect 13250 25781 13252 25812
rect 13252 25781 13284 25812
rect 13322 25781 13354 25812
rect 13354 25781 13356 25812
rect 13394 25781 13422 25812
rect 13422 25781 13428 25812
rect 13466 25781 13490 25812
rect 13490 25781 13500 25812
rect 13538 25781 13558 25812
rect 13558 25781 13572 25812
rect 13610 25781 13626 25812
rect 13626 25781 13644 25812
rect 13682 25781 13694 25812
rect 13694 25781 13716 25812
rect 13754 25781 13762 25812
rect 13762 25781 13788 25812
rect 13826 25781 13830 25812
rect 13830 25781 13860 25812
rect 13898 25781 13932 25815
rect 13970 25812 14004 25815
rect 14042 25812 14076 25815
rect 14114 25812 14148 25815
rect 14186 25812 14220 25815
rect 14258 25812 14292 25815
rect 14330 25812 14364 25815
rect 14402 25812 14436 25815
rect 14474 25812 14508 25815
rect 14546 25812 14580 25815
rect 14618 25812 14652 25815
rect 14690 25812 14724 25815
rect 13970 25781 14000 25812
rect 14000 25781 14004 25812
rect 14042 25781 14068 25812
rect 14068 25781 14076 25812
rect 14114 25781 14136 25812
rect 14136 25781 14148 25812
rect 14186 25781 14204 25812
rect 14204 25781 14220 25812
rect 14258 25781 14272 25812
rect 14272 25781 14292 25812
rect 14330 25781 14340 25812
rect 14340 25781 14364 25812
rect 14402 25781 14408 25812
rect 14408 25781 14436 25812
rect 14474 25781 14476 25812
rect 14476 25781 14508 25812
rect 14546 25781 14578 25812
rect 14578 25781 14580 25812
rect 14618 25781 14646 25812
rect 14646 25781 14652 25812
rect 14690 25781 14714 25812
rect 14714 25781 14724 25812
rect 243 25740 277 25741
rect 316 25740 350 25741
rect 389 25740 423 25741
rect 462 25740 496 25741
rect 535 25740 569 25741
rect 608 25740 642 25741
rect 681 25740 715 25741
rect 754 25740 788 25741
rect 827 25740 861 25741
rect 900 25740 934 25741
rect 973 25740 1007 25741
rect 1046 25740 1080 25741
rect 1119 25740 1153 25741
rect 1192 25740 1226 25741
rect 1265 25740 1299 25741
rect 1338 25740 1372 25741
rect 1411 25740 1445 25741
rect 243 25707 276 25740
rect 276 25707 277 25740
rect 316 25707 345 25740
rect 345 25707 350 25740
rect 389 25707 414 25740
rect 414 25707 423 25740
rect 462 25707 483 25740
rect 483 25707 496 25740
rect 535 25707 552 25740
rect 552 25707 569 25740
rect 608 25707 621 25740
rect 621 25707 642 25740
rect 681 25707 690 25740
rect 690 25707 715 25740
rect 754 25707 759 25740
rect 759 25707 788 25740
rect 827 25707 828 25740
rect 828 25707 861 25740
rect 900 25707 931 25740
rect 931 25707 934 25740
rect 973 25707 1000 25740
rect 1000 25707 1007 25740
rect 1046 25707 1069 25740
rect 1069 25707 1080 25740
rect 1119 25707 1138 25740
rect 1138 25707 1153 25740
rect 1192 25707 1207 25740
rect 1207 25707 1226 25740
rect 1265 25707 1276 25740
rect 1276 25707 1299 25740
rect 1338 25707 1345 25740
rect 1345 25707 1372 25740
rect 1411 25707 1414 25740
rect 1414 25707 1445 25740
rect 1484 25707 1518 25741
rect 1557 25740 1591 25741
rect 1630 25740 1664 25741
rect 1703 25740 1737 25741
rect 1776 25740 1810 25741
rect 1849 25740 1883 25741
rect 1922 25740 1956 25741
rect 1995 25740 2029 25741
rect 2068 25740 2102 25741
rect 2141 25740 2175 25741
rect 2214 25740 2248 25741
rect 2287 25740 2321 25741
rect 2360 25740 2394 25741
rect 2433 25740 2467 25741
rect 2506 25740 2540 25741
rect 2579 25740 2613 25741
rect 2652 25740 2686 25741
rect 1557 25707 1587 25740
rect 1587 25707 1591 25740
rect 1630 25707 1656 25740
rect 1656 25707 1664 25740
rect 1703 25707 1725 25740
rect 1725 25707 1737 25740
rect 1776 25707 1794 25740
rect 1794 25707 1810 25740
rect 1849 25707 1863 25740
rect 1863 25707 1883 25740
rect 1922 25707 1932 25740
rect 1932 25707 1956 25740
rect 1995 25707 2001 25740
rect 2001 25707 2029 25740
rect 2068 25707 2070 25740
rect 2070 25707 2102 25740
rect 2141 25707 2173 25740
rect 2173 25707 2175 25740
rect 2214 25707 2242 25740
rect 2242 25707 2248 25740
rect 2287 25707 2311 25740
rect 2311 25707 2321 25740
rect 2360 25707 2380 25740
rect 2380 25707 2394 25740
rect 2433 25707 2449 25740
rect 2449 25707 2467 25740
rect 2506 25707 2518 25740
rect 2518 25707 2540 25740
rect 2579 25707 2587 25740
rect 2587 25707 2613 25740
rect 2652 25707 2656 25740
rect 2656 25707 2686 25740
rect 2725 25707 2759 25741
rect 2798 25740 2832 25741
rect 2871 25740 2905 25741
rect 2944 25740 2978 25741
rect 3017 25740 3051 25741
rect 3090 25740 3124 25741
rect 3163 25740 3197 25741
rect 3236 25740 3270 25741
rect 3309 25740 3343 25741
rect 3382 25740 3416 25741
rect 3455 25740 3489 25741
rect 3528 25740 3562 25741
rect 3601 25740 3635 25741
rect 3674 25740 3708 25741
rect 3746 25740 3780 25741
rect 3818 25740 3852 25741
rect 3890 25740 3924 25741
rect 3962 25740 3996 25741
rect 4034 25740 4068 25741
rect 2798 25707 2829 25740
rect 2829 25707 2832 25740
rect 2871 25707 2898 25740
rect 2898 25707 2905 25740
rect 2944 25707 2967 25740
rect 2967 25707 2978 25740
rect 3017 25707 3036 25740
rect 3036 25707 3051 25740
rect 3090 25707 3105 25740
rect 3105 25707 3124 25740
rect 3163 25707 3174 25740
rect 3174 25707 3197 25740
rect 3236 25707 3243 25740
rect 3243 25707 3270 25740
rect 3309 25707 3312 25740
rect 3312 25707 3343 25740
rect 3382 25707 3415 25740
rect 3415 25707 3416 25740
rect 3455 25707 3484 25740
rect 3484 25707 3489 25740
rect 3528 25707 3553 25740
rect 3553 25707 3562 25740
rect 3601 25707 3622 25740
rect 3622 25707 3635 25740
rect 3674 25707 3691 25740
rect 3691 25707 3708 25740
rect 3746 25707 3760 25740
rect 3760 25707 3780 25740
rect 3818 25707 3829 25740
rect 3829 25707 3852 25740
rect 3890 25707 3898 25740
rect 3898 25707 3924 25740
rect 3962 25707 3967 25740
rect 3967 25707 3996 25740
rect 4034 25707 4036 25740
rect 4036 25707 4068 25740
rect 4106 25707 4140 25741
rect 4178 25740 4212 25741
rect 4250 25740 4284 25741
rect 4322 25740 4356 25741
rect 4394 25740 4428 25741
rect 4466 25740 4500 25741
rect 4538 25740 4572 25741
rect 4610 25740 4644 25741
rect 4682 25740 4716 25741
rect 4754 25740 4788 25741
rect 4826 25740 4860 25741
rect 4898 25740 4932 25741
rect 4970 25740 5004 25741
rect 5042 25740 5076 25741
rect 5114 25740 5148 25741
rect 5186 25740 5220 25741
rect 5258 25740 5292 25741
rect 4178 25707 4208 25740
rect 4208 25707 4212 25740
rect 4250 25707 4276 25740
rect 4276 25707 4284 25740
rect 4322 25707 4344 25740
rect 4344 25707 4356 25740
rect 4394 25707 4412 25740
rect 4412 25707 4428 25740
rect 4466 25707 4480 25740
rect 4480 25707 4500 25740
rect 4538 25707 4548 25740
rect 4548 25707 4572 25740
rect 4610 25707 4616 25740
rect 4616 25707 4644 25740
rect 4682 25707 4684 25740
rect 4684 25707 4716 25740
rect 4754 25707 4786 25740
rect 4786 25707 4788 25740
rect 4826 25707 4854 25740
rect 4854 25707 4860 25740
rect 4898 25707 4922 25740
rect 4922 25707 4932 25740
rect 4970 25707 4990 25740
rect 4990 25707 5004 25740
rect 5042 25707 5058 25740
rect 5058 25707 5076 25740
rect 5114 25707 5126 25740
rect 5126 25707 5148 25740
rect 5186 25707 5194 25740
rect 5194 25707 5220 25740
rect 5258 25707 5262 25740
rect 5262 25707 5292 25740
rect 5330 25707 5364 25741
rect 5402 25740 5436 25741
rect 5474 25740 5508 25741
rect 5546 25740 5580 25741
rect 5618 25740 5652 25741
rect 5690 25740 5724 25741
rect 5762 25740 5796 25741
rect 5834 25740 5868 25741
rect 5906 25740 5940 25741
rect 5978 25740 6012 25741
rect 6050 25740 6084 25741
rect 6122 25740 6156 25741
rect 6194 25740 6228 25741
rect 6266 25740 6300 25741
rect 6338 25740 6372 25741
rect 6410 25740 6444 25741
rect 6482 25740 6516 25741
rect 5402 25707 5432 25740
rect 5432 25707 5436 25740
rect 5474 25707 5500 25740
rect 5500 25707 5508 25740
rect 5546 25707 5568 25740
rect 5568 25707 5580 25740
rect 5618 25707 5636 25740
rect 5636 25707 5652 25740
rect 5690 25707 5704 25740
rect 5704 25707 5724 25740
rect 5762 25707 5772 25740
rect 5772 25707 5796 25740
rect 5834 25707 5840 25740
rect 5840 25707 5868 25740
rect 5906 25707 5908 25740
rect 5908 25707 5940 25740
rect 5978 25707 6010 25740
rect 6010 25707 6012 25740
rect 6050 25707 6078 25740
rect 6078 25707 6084 25740
rect 6122 25707 6146 25740
rect 6146 25707 6156 25740
rect 6194 25707 6214 25740
rect 6214 25707 6228 25740
rect 6266 25707 6282 25740
rect 6282 25707 6300 25740
rect 6338 25707 6350 25740
rect 6350 25707 6372 25740
rect 6410 25707 6418 25740
rect 6418 25707 6444 25740
rect 6482 25707 6486 25740
rect 6486 25707 6516 25740
rect 6554 25707 6588 25741
rect 6626 25740 6660 25741
rect 6698 25740 6732 25741
rect 6770 25740 6804 25741
rect 6842 25740 6876 25741
rect 6914 25740 6948 25741
rect 6986 25740 7020 25741
rect 7058 25740 7092 25741
rect 7130 25740 7164 25741
rect 7202 25740 7236 25741
rect 7274 25740 7308 25741
rect 7346 25740 7380 25741
rect 7418 25740 7452 25741
rect 7490 25740 7524 25741
rect 7562 25740 7596 25741
rect 7634 25740 7668 25741
rect 7706 25740 7740 25741
rect 6626 25707 6656 25740
rect 6656 25707 6660 25740
rect 6698 25707 6724 25740
rect 6724 25707 6732 25740
rect 6770 25707 6792 25740
rect 6792 25707 6804 25740
rect 6842 25707 6860 25740
rect 6860 25707 6876 25740
rect 6914 25707 6928 25740
rect 6928 25707 6948 25740
rect 6986 25707 6996 25740
rect 6996 25707 7020 25740
rect 7058 25707 7064 25740
rect 7064 25707 7092 25740
rect 7130 25707 7132 25740
rect 7132 25707 7164 25740
rect 7202 25707 7234 25740
rect 7234 25707 7236 25740
rect 7274 25707 7302 25740
rect 7302 25707 7308 25740
rect 7346 25707 7370 25740
rect 7370 25707 7380 25740
rect 7418 25707 7438 25740
rect 7438 25707 7452 25740
rect 7490 25707 7506 25740
rect 7506 25707 7524 25740
rect 7562 25707 7574 25740
rect 7574 25707 7596 25740
rect 7634 25707 7642 25740
rect 7642 25707 7668 25740
rect 7706 25707 7710 25740
rect 7710 25707 7740 25740
rect 7778 25707 7812 25741
rect 7850 25740 7884 25741
rect 7922 25740 7956 25741
rect 7994 25740 8028 25741
rect 8066 25740 8100 25741
rect 8138 25740 8172 25741
rect 8210 25740 8244 25741
rect 8282 25740 8316 25741
rect 8354 25740 8388 25741
rect 8426 25740 8460 25741
rect 8498 25740 8532 25741
rect 8570 25740 8604 25741
rect 8642 25740 8676 25741
rect 8714 25740 8748 25741
rect 8786 25740 8820 25741
rect 8858 25740 8892 25741
rect 8930 25740 8964 25741
rect 7850 25707 7880 25740
rect 7880 25707 7884 25740
rect 7922 25707 7948 25740
rect 7948 25707 7956 25740
rect 7994 25707 8016 25740
rect 8016 25707 8028 25740
rect 8066 25707 8084 25740
rect 8084 25707 8100 25740
rect 8138 25707 8152 25740
rect 8152 25707 8172 25740
rect 8210 25707 8220 25740
rect 8220 25707 8244 25740
rect 8282 25707 8288 25740
rect 8288 25707 8316 25740
rect 8354 25707 8356 25740
rect 8356 25707 8388 25740
rect 8426 25707 8458 25740
rect 8458 25707 8460 25740
rect 8498 25707 8526 25740
rect 8526 25707 8532 25740
rect 8570 25707 8594 25740
rect 8594 25707 8604 25740
rect 8642 25707 8662 25740
rect 8662 25707 8676 25740
rect 8714 25707 8730 25740
rect 8730 25707 8748 25740
rect 8786 25707 8798 25740
rect 8798 25707 8820 25740
rect 8858 25707 8866 25740
rect 8866 25707 8892 25740
rect 8930 25707 8934 25740
rect 8934 25707 8964 25740
rect 9002 25707 9036 25741
rect 9074 25740 9108 25741
rect 9146 25740 9180 25741
rect 9218 25740 9252 25741
rect 9290 25740 9324 25741
rect 9362 25740 9396 25741
rect 9434 25740 9468 25741
rect 9506 25740 9540 25741
rect 9578 25740 9612 25741
rect 9650 25740 9684 25741
rect 9722 25740 9756 25741
rect 9794 25740 9828 25741
rect 9866 25740 9900 25741
rect 9938 25740 9972 25741
rect 10010 25740 10044 25741
rect 10082 25740 10116 25741
rect 10154 25740 10188 25741
rect 9074 25707 9104 25740
rect 9104 25707 9108 25740
rect 9146 25707 9172 25740
rect 9172 25707 9180 25740
rect 9218 25707 9240 25740
rect 9240 25707 9252 25740
rect 9290 25707 9308 25740
rect 9308 25707 9324 25740
rect 9362 25707 9376 25740
rect 9376 25707 9396 25740
rect 9434 25707 9444 25740
rect 9444 25707 9468 25740
rect 9506 25707 9512 25740
rect 9512 25707 9540 25740
rect 9578 25707 9580 25740
rect 9580 25707 9612 25740
rect 9650 25707 9682 25740
rect 9682 25707 9684 25740
rect 9722 25707 9750 25740
rect 9750 25707 9756 25740
rect 9794 25707 9818 25740
rect 9818 25707 9828 25740
rect 9866 25707 9886 25740
rect 9886 25707 9900 25740
rect 9938 25707 9954 25740
rect 9954 25707 9972 25740
rect 10010 25707 10022 25740
rect 10022 25707 10044 25740
rect 10082 25707 10090 25740
rect 10090 25707 10116 25740
rect 10154 25707 10158 25740
rect 10158 25707 10188 25740
rect 10226 25707 10260 25741
rect 10298 25740 10332 25741
rect 10370 25740 10404 25741
rect 10442 25740 10476 25741
rect 10514 25740 10548 25741
rect 10586 25740 10620 25741
rect 10658 25740 10692 25741
rect 10730 25740 10764 25741
rect 10802 25740 10836 25741
rect 10874 25740 10908 25741
rect 10946 25740 10980 25741
rect 11018 25740 11052 25741
rect 11090 25740 11124 25741
rect 11162 25740 11196 25741
rect 11234 25740 11268 25741
rect 11306 25740 11340 25741
rect 11378 25740 11412 25741
rect 10298 25707 10328 25740
rect 10328 25707 10332 25740
rect 10370 25707 10396 25740
rect 10396 25707 10404 25740
rect 10442 25707 10464 25740
rect 10464 25707 10476 25740
rect 10514 25707 10532 25740
rect 10532 25707 10548 25740
rect 10586 25707 10600 25740
rect 10600 25707 10620 25740
rect 10658 25707 10668 25740
rect 10668 25707 10692 25740
rect 10730 25707 10736 25740
rect 10736 25707 10764 25740
rect 10802 25707 10804 25740
rect 10804 25707 10836 25740
rect 10874 25707 10906 25740
rect 10906 25707 10908 25740
rect 10946 25707 10974 25740
rect 10974 25707 10980 25740
rect 11018 25707 11042 25740
rect 11042 25707 11052 25740
rect 11090 25707 11110 25740
rect 11110 25707 11124 25740
rect 11162 25707 11178 25740
rect 11178 25707 11196 25740
rect 11234 25707 11246 25740
rect 11246 25707 11268 25740
rect 11306 25707 11314 25740
rect 11314 25707 11340 25740
rect 11378 25707 11382 25740
rect 11382 25707 11412 25740
rect 11450 25707 11484 25741
rect 11522 25740 11556 25741
rect 11594 25740 11628 25741
rect 11666 25740 11700 25741
rect 11738 25740 11772 25741
rect 11810 25740 11844 25741
rect 11882 25740 11916 25741
rect 11954 25740 11988 25741
rect 12026 25740 12060 25741
rect 12098 25740 12132 25741
rect 12170 25740 12204 25741
rect 12242 25740 12276 25741
rect 12314 25740 12348 25741
rect 12386 25740 12420 25741
rect 12458 25740 12492 25741
rect 12530 25740 12564 25741
rect 12602 25740 12636 25741
rect 11522 25707 11552 25740
rect 11552 25707 11556 25740
rect 11594 25707 11620 25740
rect 11620 25707 11628 25740
rect 11666 25707 11688 25740
rect 11688 25707 11700 25740
rect 11738 25707 11756 25740
rect 11756 25707 11772 25740
rect 11810 25707 11824 25740
rect 11824 25707 11844 25740
rect 11882 25707 11892 25740
rect 11892 25707 11916 25740
rect 11954 25707 11960 25740
rect 11960 25707 11988 25740
rect 12026 25707 12028 25740
rect 12028 25707 12060 25740
rect 12098 25707 12130 25740
rect 12130 25707 12132 25740
rect 12170 25707 12198 25740
rect 12198 25707 12204 25740
rect 12242 25707 12266 25740
rect 12266 25707 12276 25740
rect 12314 25707 12334 25740
rect 12334 25707 12348 25740
rect 12386 25707 12402 25740
rect 12402 25707 12420 25740
rect 12458 25707 12470 25740
rect 12470 25707 12492 25740
rect 12530 25707 12538 25740
rect 12538 25707 12564 25740
rect 12602 25707 12606 25740
rect 12606 25707 12636 25740
rect 12674 25707 12708 25741
rect 12746 25740 12780 25741
rect 12818 25740 12852 25741
rect 12890 25740 12924 25741
rect 12962 25740 12996 25741
rect 13034 25740 13068 25741
rect 13106 25740 13140 25741
rect 13178 25740 13212 25741
rect 13250 25740 13284 25741
rect 13322 25740 13356 25741
rect 13394 25740 13428 25741
rect 13466 25740 13500 25741
rect 13538 25740 13572 25741
rect 13610 25740 13644 25741
rect 13682 25740 13716 25741
rect 13754 25740 13788 25741
rect 13826 25740 13860 25741
rect 12746 25707 12776 25740
rect 12776 25707 12780 25740
rect 12818 25707 12844 25740
rect 12844 25707 12852 25740
rect 12890 25707 12912 25740
rect 12912 25707 12924 25740
rect 12962 25707 12980 25740
rect 12980 25707 12996 25740
rect 13034 25707 13048 25740
rect 13048 25707 13068 25740
rect 13106 25707 13116 25740
rect 13116 25707 13140 25740
rect 13178 25707 13184 25740
rect 13184 25707 13212 25740
rect 13250 25707 13252 25740
rect 13252 25707 13284 25740
rect 13322 25707 13354 25740
rect 13354 25707 13356 25740
rect 13394 25707 13422 25740
rect 13422 25707 13428 25740
rect 13466 25707 13490 25740
rect 13490 25707 13500 25740
rect 13538 25707 13558 25740
rect 13558 25707 13572 25740
rect 13610 25707 13626 25740
rect 13626 25707 13644 25740
rect 13682 25707 13694 25740
rect 13694 25707 13716 25740
rect 13754 25707 13762 25740
rect 13762 25707 13788 25740
rect 13826 25707 13830 25740
rect 13830 25707 13860 25740
rect 13898 25707 13932 25741
rect 13970 25740 14004 25741
rect 14042 25740 14076 25741
rect 14114 25740 14148 25741
rect 14186 25740 14220 25741
rect 14258 25740 14292 25741
rect 14330 25740 14364 25741
rect 14402 25740 14436 25741
rect 14474 25740 14508 25741
rect 14546 25740 14580 25741
rect 14618 25740 14652 25741
rect 14690 25740 14724 25741
rect 13970 25707 14000 25740
rect 14000 25707 14004 25740
rect 14042 25707 14068 25740
rect 14068 25707 14076 25740
rect 14114 25707 14136 25740
rect 14136 25707 14148 25740
rect 14186 25707 14204 25740
rect 14204 25707 14220 25740
rect 14258 25707 14272 25740
rect 14272 25707 14292 25740
rect 14330 25707 14340 25740
rect 14340 25707 14364 25740
rect 14402 25707 14408 25740
rect 14408 25707 14436 25740
rect 14474 25707 14476 25740
rect 14476 25707 14508 25740
rect 14546 25707 14578 25740
rect 14578 25707 14580 25740
rect 14618 25707 14646 25740
rect 14646 25707 14652 25740
rect 14690 25707 14714 25740
rect 14714 25707 14724 25740
rect 243 25634 276 25667
rect 276 25634 277 25667
rect 316 25634 345 25667
rect 345 25634 350 25667
rect 389 25634 414 25667
rect 414 25634 423 25667
rect 462 25634 483 25667
rect 483 25634 496 25667
rect 535 25634 552 25667
rect 552 25634 569 25667
rect 608 25634 621 25667
rect 621 25634 642 25667
rect 681 25634 690 25667
rect 690 25634 715 25667
rect 754 25634 759 25667
rect 759 25634 788 25667
rect 827 25634 828 25667
rect 828 25634 861 25667
rect 900 25634 931 25667
rect 931 25634 934 25667
rect 973 25634 1000 25667
rect 1000 25634 1007 25667
rect 1046 25634 1069 25667
rect 1069 25634 1080 25667
rect 1119 25634 1138 25667
rect 1138 25634 1153 25667
rect 1192 25634 1207 25667
rect 1207 25634 1226 25667
rect 1265 25634 1276 25667
rect 1276 25634 1299 25667
rect 1338 25634 1345 25667
rect 1345 25634 1372 25667
rect 1411 25634 1414 25667
rect 1414 25634 1445 25667
rect 243 25633 277 25634
rect 316 25633 350 25634
rect 389 25633 423 25634
rect 462 25633 496 25634
rect 535 25633 569 25634
rect 608 25633 642 25634
rect 681 25633 715 25634
rect 754 25633 788 25634
rect 827 25633 861 25634
rect 900 25633 934 25634
rect 973 25633 1007 25634
rect 1046 25633 1080 25634
rect 1119 25633 1153 25634
rect 1192 25633 1226 25634
rect 1265 25633 1299 25634
rect 1338 25633 1372 25634
rect 1411 25633 1445 25634
rect 1484 25633 1518 25667
rect 1557 25634 1587 25667
rect 1587 25634 1591 25667
rect 1630 25634 1656 25667
rect 1656 25634 1664 25667
rect 1703 25634 1725 25667
rect 1725 25634 1737 25667
rect 1776 25634 1794 25667
rect 1794 25634 1810 25667
rect 1849 25634 1863 25667
rect 1863 25634 1883 25667
rect 1922 25634 1932 25667
rect 1932 25634 1956 25667
rect 1995 25634 2001 25667
rect 2001 25634 2029 25667
rect 2068 25634 2070 25667
rect 2070 25634 2102 25667
rect 2141 25634 2173 25667
rect 2173 25634 2175 25667
rect 2214 25634 2242 25667
rect 2242 25634 2248 25667
rect 2287 25634 2311 25667
rect 2311 25634 2321 25667
rect 2360 25634 2380 25667
rect 2380 25634 2394 25667
rect 2433 25634 2449 25667
rect 2449 25634 2467 25667
rect 2506 25634 2518 25667
rect 2518 25634 2540 25667
rect 2579 25634 2587 25667
rect 2587 25634 2613 25667
rect 2652 25634 2656 25667
rect 2656 25634 2686 25667
rect 1557 25633 1591 25634
rect 1630 25633 1664 25634
rect 1703 25633 1737 25634
rect 1776 25633 1810 25634
rect 1849 25633 1883 25634
rect 1922 25633 1956 25634
rect 1995 25633 2029 25634
rect 2068 25633 2102 25634
rect 2141 25633 2175 25634
rect 2214 25633 2248 25634
rect 2287 25633 2321 25634
rect 2360 25633 2394 25634
rect 2433 25633 2467 25634
rect 2506 25633 2540 25634
rect 2579 25633 2613 25634
rect 2652 25633 2686 25634
rect 2725 25633 2759 25667
rect 2798 25634 2829 25667
rect 2829 25634 2832 25667
rect 2871 25634 2898 25667
rect 2898 25634 2905 25667
rect 2944 25634 2967 25667
rect 2967 25634 2978 25667
rect 3017 25634 3036 25667
rect 3036 25634 3051 25667
rect 3090 25634 3105 25667
rect 3105 25634 3124 25667
rect 3163 25634 3174 25667
rect 3174 25634 3197 25667
rect 3236 25634 3243 25667
rect 3243 25634 3270 25667
rect 3309 25634 3312 25667
rect 3312 25634 3343 25667
rect 3382 25634 3415 25667
rect 3415 25634 3416 25667
rect 3455 25634 3484 25667
rect 3484 25634 3489 25667
rect 3528 25634 3553 25667
rect 3553 25634 3562 25667
rect 3601 25634 3622 25667
rect 3622 25634 3635 25667
rect 3674 25634 3691 25667
rect 3691 25634 3708 25667
rect 3746 25634 3760 25667
rect 3760 25634 3780 25667
rect 3818 25634 3829 25667
rect 3829 25634 3852 25667
rect 3890 25634 3898 25667
rect 3898 25634 3924 25667
rect 3962 25634 3967 25667
rect 3967 25634 3996 25667
rect 4034 25634 4036 25667
rect 4036 25634 4068 25667
rect 2798 25633 2832 25634
rect 2871 25633 2905 25634
rect 2944 25633 2978 25634
rect 3017 25633 3051 25634
rect 3090 25633 3124 25634
rect 3163 25633 3197 25634
rect 3236 25633 3270 25634
rect 3309 25633 3343 25634
rect 3382 25633 3416 25634
rect 3455 25633 3489 25634
rect 3528 25633 3562 25634
rect 3601 25633 3635 25634
rect 3674 25633 3708 25634
rect 3746 25633 3780 25634
rect 3818 25633 3852 25634
rect 3890 25633 3924 25634
rect 3962 25633 3996 25634
rect 4034 25633 4068 25634
rect 4106 25633 4140 25667
rect 4178 25634 4208 25667
rect 4208 25634 4212 25667
rect 4250 25634 4276 25667
rect 4276 25634 4284 25667
rect 4322 25634 4344 25667
rect 4344 25634 4356 25667
rect 4394 25634 4412 25667
rect 4412 25634 4428 25667
rect 4466 25634 4480 25667
rect 4480 25634 4500 25667
rect 4538 25634 4548 25667
rect 4548 25634 4572 25667
rect 4610 25634 4616 25667
rect 4616 25634 4644 25667
rect 4682 25634 4684 25667
rect 4684 25634 4716 25667
rect 4754 25634 4786 25667
rect 4786 25634 4788 25667
rect 4826 25634 4854 25667
rect 4854 25634 4860 25667
rect 4898 25634 4922 25667
rect 4922 25634 4932 25667
rect 4970 25634 4990 25667
rect 4990 25634 5004 25667
rect 5042 25634 5058 25667
rect 5058 25634 5076 25667
rect 5114 25634 5126 25667
rect 5126 25634 5148 25667
rect 5186 25634 5194 25667
rect 5194 25634 5220 25667
rect 5258 25634 5262 25667
rect 5262 25634 5292 25667
rect 4178 25633 4212 25634
rect 4250 25633 4284 25634
rect 4322 25633 4356 25634
rect 4394 25633 4428 25634
rect 4466 25633 4500 25634
rect 4538 25633 4572 25634
rect 4610 25633 4644 25634
rect 4682 25633 4716 25634
rect 4754 25633 4788 25634
rect 4826 25633 4860 25634
rect 4898 25633 4932 25634
rect 4970 25633 5004 25634
rect 5042 25633 5076 25634
rect 5114 25633 5148 25634
rect 5186 25633 5220 25634
rect 5258 25633 5292 25634
rect 5330 25633 5364 25667
rect 5402 25634 5432 25667
rect 5432 25634 5436 25667
rect 5474 25634 5500 25667
rect 5500 25634 5508 25667
rect 5546 25634 5568 25667
rect 5568 25634 5580 25667
rect 5618 25634 5636 25667
rect 5636 25634 5652 25667
rect 5690 25634 5704 25667
rect 5704 25634 5724 25667
rect 5762 25634 5772 25667
rect 5772 25634 5796 25667
rect 5834 25634 5840 25667
rect 5840 25634 5868 25667
rect 5906 25634 5908 25667
rect 5908 25634 5940 25667
rect 5978 25634 6010 25667
rect 6010 25634 6012 25667
rect 6050 25634 6078 25667
rect 6078 25634 6084 25667
rect 6122 25634 6146 25667
rect 6146 25634 6156 25667
rect 6194 25634 6214 25667
rect 6214 25634 6228 25667
rect 6266 25634 6282 25667
rect 6282 25634 6300 25667
rect 6338 25634 6350 25667
rect 6350 25634 6372 25667
rect 6410 25634 6418 25667
rect 6418 25634 6444 25667
rect 6482 25634 6486 25667
rect 6486 25634 6516 25667
rect 5402 25633 5436 25634
rect 5474 25633 5508 25634
rect 5546 25633 5580 25634
rect 5618 25633 5652 25634
rect 5690 25633 5724 25634
rect 5762 25633 5796 25634
rect 5834 25633 5868 25634
rect 5906 25633 5940 25634
rect 5978 25633 6012 25634
rect 6050 25633 6084 25634
rect 6122 25633 6156 25634
rect 6194 25633 6228 25634
rect 6266 25633 6300 25634
rect 6338 25633 6372 25634
rect 6410 25633 6444 25634
rect 6482 25633 6516 25634
rect 6554 25633 6588 25667
rect 6626 25634 6656 25667
rect 6656 25634 6660 25667
rect 6698 25634 6724 25667
rect 6724 25634 6732 25667
rect 6770 25634 6792 25667
rect 6792 25634 6804 25667
rect 6842 25634 6860 25667
rect 6860 25634 6876 25667
rect 6914 25634 6928 25667
rect 6928 25634 6948 25667
rect 6986 25634 6996 25667
rect 6996 25634 7020 25667
rect 7058 25634 7064 25667
rect 7064 25634 7092 25667
rect 7130 25634 7132 25667
rect 7132 25634 7164 25667
rect 7202 25634 7234 25667
rect 7234 25634 7236 25667
rect 7274 25634 7302 25667
rect 7302 25634 7308 25667
rect 7346 25634 7370 25667
rect 7370 25634 7380 25667
rect 7418 25634 7438 25667
rect 7438 25634 7452 25667
rect 7490 25634 7506 25667
rect 7506 25634 7524 25667
rect 7562 25634 7574 25667
rect 7574 25634 7596 25667
rect 7634 25634 7642 25667
rect 7642 25634 7668 25667
rect 7706 25634 7710 25667
rect 7710 25634 7740 25667
rect 6626 25633 6660 25634
rect 6698 25633 6732 25634
rect 6770 25633 6804 25634
rect 6842 25633 6876 25634
rect 6914 25633 6948 25634
rect 6986 25633 7020 25634
rect 7058 25633 7092 25634
rect 7130 25633 7164 25634
rect 7202 25633 7236 25634
rect 7274 25633 7308 25634
rect 7346 25633 7380 25634
rect 7418 25633 7452 25634
rect 7490 25633 7524 25634
rect 7562 25633 7596 25634
rect 7634 25633 7668 25634
rect 7706 25633 7740 25634
rect 7778 25633 7812 25667
rect 7850 25634 7880 25667
rect 7880 25634 7884 25667
rect 7922 25634 7948 25667
rect 7948 25634 7956 25667
rect 7994 25634 8016 25667
rect 8016 25634 8028 25667
rect 8066 25634 8084 25667
rect 8084 25634 8100 25667
rect 8138 25634 8152 25667
rect 8152 25634 8172 25667
rect 8210 25634 8220 25667
rect 8220 25634 8244 25667
rect 8282 25634 8288 25667
rect 8288 25634 8316 25667
rect 8354 25634 8356 25667
rect 8356 25634 8388 25667
rect 8426 25634 8458 25667
rect 8458 25634 8460 25667
rect 8498 25634 8526 25667
rect 8526 25634 8532 25667
rect 8570 25634 8594 25667
rect 8594 25634 8604 25667
rect 8642 25634 8662 25667
rect 8662 25634 8676 25667
rect 8714 25634 8730 25667
rect 8730 25634 8748 25667
rect 8786 25634 8798 25667
rect 8798 25634 8820 25667
rect 8858 25634 8866 25667
rect 8866 25634 8892 25667
rect 8930 25634 8934 25667
rect 8934 25634 8964 25667
rect 7850 25633 7884 25634
rect 7922 25633 7956 25634
rect 7994 25633 8028 25634
rect 8066 25633 8100 25634
rect 8138 25633 8172 25634
rect 8210 25633 8244 25634
rect 8282 25633 8316 25634
rect 8354 25633 8388 25634
rect 8426 25633 8460 25634
rect 8498 25633 8532 25634
rect 8570 25633 8604 25634
rect 8642 25633 8676 25634
rect 8714 25633 8748 25634
rect 8786 25633 8820 25634
rect 8858 25633 8892 25634
rect 8930 25633 8964 25634
rect 9002 25633 9036 25667
rect 9074 25634 9104 25667
rect 9104 25634 9108 25667
rect 9146 25634 9172 25667
rect 9172 25634 9180 25667
rect 9218 25634 9240 25667
rect 9240 25634 9252 25667
rect 9290 25634 9308 25667
rect 9308 25634 9324 25667
rect 9362 25634 9376 25667
rect 9376 25634 9396 25667
rect 9434 25634 9444 25667
rect 9444 25634 9468 25667
rect 9506 25634 9512 25667
rect 9512 25634 9540 25667
rect 9578 25634 9580 25667
rect 9580 25634 9612 25667
rect 9650 25634 9682 25667
rect 9682 25634 9684 25667
rect 9722 25634 9750 25667
rect 9750 25634 9756 25667
rect 9794 25634 9818 25667
rect 9818 25634 9828 25667
rect 9866 25634 9886 25667
rect 9886 25634 9900 25667
rect 9938 25634 9954 25667
rect 9954 25634 9972 25667
rect 10010 25634 10022 25667
rect 10022 25634 10044 25667
rect 10082 25634 10090 25667
rect 10090 25634 10116 25667
rect 10154 25634 10158 25667
rect 10158 25634 10188 25667
rect 9074 25633 9108 25634
rect 9146 25633 9180 25634
rect 9218 25633 9252 25634
rect 9290 25633 9324 25634
rect 9362 25633 9396 25634
rect 9434 25633 9468 25634
rect 9506 25633 9540 25634
rect 9578 25633 9612 25634
rect 9650 25633 9684 25634
rect 9722 25633 9756 25634
rect 9794 25633 9828 25634
rect 9866 25633 9900 25634
rect 9938 25633 9972 25634
rect 10010 25633 10044 25634
rect 10082 25633 10116 25634
rect 10154 25633 10188 25634
rect 10226 25633 10260 25667
rect 10298 25634 10328 25667
rect 10328 25634 10332 25667
rect 10370 25634 10396 25667
rect 10396 25634 10404 25667
rect 10442 25634 10464 25667
rect 10464 25634 10476 25667
rect 10514 25634 10532 25667
rect 10532 25634 10548 25667
rect 10586 25634 10600 25667
rect 10600 25634 10620 25667
rect 10658 25634 10668 25667
rect 10668 25634 10692 25667
rect 10730 25634 10736 25667
rect 10736 25634 10764 25667
rect 10802 25634 10804 25667
rect 10804 25634 10836 25667
rect 10874 25634 10906 25667
rect 10906 25634 10908 25667
rect 10946 25634 10974 25667
rect 10974 25634 10980 25667
rect 11018 25634 11042 25667
rect 11042 25634 11052 25667
rect 11090 25634 11110 25667
rect 11110 25634 11124 25667
rect 11162 25634 11178 25667
rect 11178 25634 11196 25667
rect 11234 25634 11246 25667
rect 11246 25634 11268 25667
rect 11306 25634 11314 25667
rect 11314 25634 11340 25667
rect 11378 25634 11382 25667
rect 11382 25634 11412 25667
rect 10298 25633 10332 25634
rect 10370 25633 10404 25634
rect 10442 25633 10476 25634
rect 10514 25633 10548 25634
rect 10586 25633 10620 25634
rect 10658 25633 10692 25634
rect 10730 25633 10764 25634
rect 10802 25633 10836 25634
rect 10874 25633 10908 25634
rect 10946 25633 10980 25634
rect 11018 25633 11052 25634
rect 11090 25633 11124 25634
rect 11162 25633 11196 25634
rect 11234 25633 11268 25634
rect 11306 25633 11340 25634
rect 11378 25633 11412 25634
rect 11450 25633 11484 25667
rect 11522 25634 11552 25667
rect 11552 25634 11556 25667
rect 11594 25634 11620 25667
rect 11620 25634 11628 25667
rect 11666 25634 11688 25667
rect 11688 25634 11700 25667
rect 11738 25634 11756 25667
rect 11756 25634 11772 25667
rect 11810 25634 11824 25667
rect 11824 25634 11844 25667
rect 11882 25634 11892 25667
rect 11892 25634 11916 25667
rect 11954 25634 11960 25667
rect 11960 25634 11988 25667
rect 12026 25634 12028 25667
rect 12028 25634 12060 25667
rect 12098 25634 12130 25667
rect 12130 25634 12132 25667
rect 12170 25634 12198 25667
rect 12198 25634 12204 25667
rect 12242 25634 12266 25667
rect 12266 25634 12276 25667
rect 12314 25634 12334 25667
rect 12334 25634 12348 25667
rect 12386 25634 12402 25667
rect 12402 25634 12420 25667
rect 12458 25634 12470 25667
rect 12470 25634 12492 25667
rect 12530 25634 12538 25667
rect 12538 25634 12564 25667
rect 12602 25634 12606 25667
rect 12606 25634 12636 25667
rect 11522 25633 11556 25634
rect 11594 25633 11628 25634
rect 11666 25633 11700 25634
rect 11738 25633 11772 25634
rect 11810 25633 11844 25634
rect 11882 25633 11916 25634
rect 11954 25633 11988 25634
rect 12026 25633 12060 25634
rect 12098 25633 12132 25634
rect 12170 25633 12204 25634
rect 12242 25633 12276 25634
rect 12314 25633 12348 25634
rect 12386 25633 12420 25634
rect 12458 25633 12492 25634
rect 12530 25633 12564 25634
rect 12602 25633 12636 25634
rect 12674 25633 12708 25667
rect 12746 25634 12776 25667
rect 12776 25634 12780 25667
rect 12818 25634 12844 25667
rect 12844 25634 12852 25667
rect 12890 25634 12912 25667
rect 12912 25634 12924 25667
rect 12962 25634 12980 25667
rect 12980 25634 12996 25667
rect 13034 25634 13048 25667
rect 13048 25634 13068 25667
rect 13106 25634 13116 25667
rect 13116 25634 13140 25667
rect 13178 25634 13184 25667
rect 13184 25634 13212 25667
rect 13250 25634 13252 25667
rect 13252 25634 13284 25667
rect 13322 25634 13354 25667
rect 13354 25634 13356 25667
rect 13394 25634 13422 25667
rect 13422 25634 13428 25667
rect 13466 25634 13490 25667
rect 13490 25634 13500 25667
rect 13538 25634 13558 25667
rect 13558 25634 13572 25667
rect 13610 25634 13626 25667
rect 13626 25634 13644 25667
rect 13682 25634 13694 25667
rect 13694 25634 13716 25667
rect 13754 25634 13762 25667
rect 13762 25634 13788 25667
rect 13826 25634 13830 25667
rect 13830 25634 13860 25667
rect 12746 25633 12780 25634
rect 12818 25633 12852 25634
rect 12890 25633 12924 25634
rect 12962 25633 12996 25634
rect 13034 25633 13068 25634
rect 13106 25633 13140 25634
rect 13178 25633 13212 25634
rect 13250 25633 13284 25634
rect 13322 25633 13356 25634
rect 13394 25633 13428 25634
rect 13466 25633 13500 25634
rect 13538 25633 13572 25634
rect 13610 25633 13644 25634
rect 13682 25633 13716 25634
rect 13754 25633 13788 25634
rect 13826 25633 13860 25634
rect 13898 25633 13932 25667
rect 13970 25634 14000 25667
rect 14000 25634 14004 25667
rect 14042 25634 14068 25667
rect 14068 25634 14076 25667
rect 14114 25634 14136 25667
rect 14136 25634 14148 25667
rect 14186 25634 14204 25667
rect 14204 25634 14220 25667
rect 14258 25634 14272 25667
rect 14272 25634 14292 25667
rect 14330 25634 14340 25667
rect 14340 25634 14364 25667
rect 14402 25634 14408 25667
rect 14408 25634 14436 25667
rect 14474 25634 14476 25667
rect 14476 25634 14508 25667
rect 14546 25634 14578 25667
rect 14578 25634 14580 25667
rect 14618 25634 14646 25667
rect 14646 25634 14652 25667
rect 14690 25634 14714 25667
rect 14714 25634 14724 25667
rect 13970 25633 14004 25634
rect 14042 25633 14076 25634
rect 14114 25633 14148 25634
rect 14186 25633 14220 25634
rect 14258 25633 14292 25634
rect 14330 25633 14364 25634
rect 14402 25633 14436 25634
rect 14474 25633 14508 25634
rect 14546 25633 14580 25634
rect 14618 25633 14652 25634
rect 14690 25633 14724 25634
rect 88 25007 122 25041
rect 161 25034 195 25041
rect 234 25034 268 25041
rect 307 25034 341 25041
rect 380 25034 414 25041
rect 453 25034 487 25041
rect 526 25034 560 25041
rect 599 25034 633 25041
rect 672 25034 706 25041
rect 745 25034 779 25041
rect 818 25034 852 25041
rect 891 25034 925 25041
rect 964 25034 998 25041
rect 1037 25034 1071 25041
rect 1110 25034 1144 25041
rect 1183 25034 1217 25041
rect 1256 25034 1290 25041
rect 1329 25034 1363 25041
rect 1402 25034 1436 25041
rect 1475 25034 1509 25041
rect 1548 25034 1582 25041
rect 1621 25034 1655 25041
rect 1694 25034 1728 25041
rect 1767 25034 1801 25041
rect 1840 25034 1874 25041
rect 1913 25034 1947 25041
rect 1986 25034 2020 25041
rect 2059 25034 2093 25041
rect 2132 25034 2166 25041
rect 2205 25034 2239 25041
rect 161 25007 193 25034
rect 193 25007 195 25034
rect 234 25007 262 25034
rect 262 25007 268 25034
rect 307 25007 331 25034
rect 331 25007 341 25034
rect 380 25007 400 25034
rect 400 25007 414 25034
rect 453 25007 469 25034
rect 469 25007 487 25034
rect 526 25007 538 25034
rect 538 25007 560 25034
rect 599 25007 607 25034
rect 607 25007 633 25034
rect 672 25007 676 25034
rect 676 25007 706 25034
rect 745 25007 779 25034
rect 818 25007 848 25034
rect 848 25007 852 25034
rect 891 25007 917 25034
rect 917 25007 925 25034
rect 964 25007 986 25034
rect 986 25007 998 25034
rect 1037 25007 1054 25034
rect 1054 25007 1071 25034
rect 1110 25007 1122 25034
rect 1122 25007 1144 25034
rect 1183 25007 1190 25034
rect 1190 25007 1217 25034
rect 1256 25007 1258 25034
rect 1258 25007 1290 25034
rect 1329 25007 1360 25034
rect 1360 25007 1363 25034
rect 1402 25007 1428 25034
rect 1428 25007 1436 25034
rect 1475 25007 1496 25034
rect 1496 25007 1509 25034
rect 1548 25007 1564 25034
rect 1564 25007 1582 25034
rect 1621 25007 1632 25034
rect 1632 25007 1655 25034
rect 1694 25007 1700 25034
rect 1700 25007 1728 25034
rect 1767 25007 1768 25034
rect 1768 25007 1801 25034
rect 1840 25007 1870 25034
rect 1870 25007 1874 25034
rect 1913 25007 1938 25034
rect 1938 25007 1947 25034
rect 1986 25007 2006 25034
rect 2006 25007 2020 25034
rect 2059 25007 2074 25034
rect 2074 25007 2093 25034
rect 2132 25007 2142 25034
rect 2142 25007 2166 25034
rect 2205 25007 2210 25034
rect 2210 25007 2239 25034
rect 2278 25007 2312 25041
rect 2351 25034 2385 25041
rect 2424 25034 2458 25041
rect 2497 25034 2531 25041
rect 2570 25034 2604 25041
rect 2643 25034 2677 25041
rect 2716 25034 2750 25041
rect 2789 25034 2823 25041
rect 2862 25034 2896 25041
rect 2935 25034 2969 25041
rect 3008 25034 3042 25041
rect 3081 25034 3115 25041
rect 3154 25034 3188 25041
rect 3227 25034 3261 25041
rect 3300 25034 3334 25041
rect 3373 25034 3407 25041
rect 3446 25034 3480 25041
rect 3519 25034 3553 25041
rect 3592 25034 3626 25041
rect 3665 25034 3699 25041
rect 3738 25034 3772 25041
rect 3811 25034 3845 25041
rect 3884 25034 3918 25041
rect 3957 25034 3991 25041
rect 4030 25034 4064 25041
rect 4103 25034 4137 25041
rect 4176 25034 4210 25041
rect 4249 25034 4283 25041
rect 4322 25034 4356 25041
rect 4395 25034 4429 25041
rect 4468 25034 14870 25041
rect 2351 25007 2380 25034
rect 2380 25007 2385 25034
rect 2424 25007 2448 25034
rect 2448 25007 2458 25034
rect 2497 25007 2516 25034
rect 2516 25007 2531 25034
rect 2570 25007 2584 25034
rect 2584 25007 2604 25034
rect 2643 25007 2652 25034
rect 2652 25007 2677 25034
rect 2716 25007 2720 25034
rect 2720 25007 2750 25034
rect 2789 25007 2822 25034
rect 2822 25007 2823 25034
rect 2862 25007 2890 25034
rect 2890 25007 2896 25034
rect 2935 25007 2958 25034
rect 2958 25007 2969 25034
rect 3008 25007 3026 25034
rect 3026 25007 3042 25034
rect 3081 25007 3094 25034
rect 3094 25007 3115 25034
rect 3154 25007 3162 25034
rect 3162 25007 3188 25034
rect 3227 25007 3230 25034
rect 3230 25007 3261 25034
rect 3300 25007 3332 25034
rect 3332 25007 3334 25034
rect 3373 25007 3400 25034
rect 3400 25007 3407 25034
rect 3446 25007 3468 25034
rect 3468 25007 3480 25034
rect 3519 25007 3536 25034
rect 3536 25007 3553 25034
rect 3592 25007 3604 25034
rect 3604 25007 3626 25034
rect 3665 25007 3672 25034
rect 3672 25007 3699 25034
rect 3738 25007 3740 25034
rect 3740 25007 3772 25034
rect 3811 25007 3842 25034
rect 3842 25007 3845 25034
rect 3884 25007 3910 25034
rect 3910 25007 3918 25034
rect 3957 25007 3978 25034
rect 3978 25007 3991 25034
rect 4030 25007 4046 25034
rect 4046 25007 4064 25034
rect 4103 25007 4114 25034
rect 4114 25007 4137 25034
rect 4176 25007 4182 25034
rect 4182 25007 4210 25034
rect 4249 25007 4250 25034
rect 4250 25007 4283 25034
rect 4322 25007 4352 25034
rect 4352 25007 4356 25034
rect 4395 25007 4420 25034
rect 4420 25007 4429 25034
rect 4468 25000 4488 25034
rect 4488 25000 4522 25034
rect 4522 25000 4556 25034
rect 4556 25000 4590 25034
rect 4590 25000 4624 25034
rect 4624 25000 4658 25034
rect 4658 25000 4692 25034
rect 4692 25000 4726 25034
rect 4726 25000 4760 25034
rect 4760 25000 4794 25034
rect 4794 25000 4828 25034
rect 4828 25000 4862 25034
rect 4862 25000 4896 25034
rect 4896 25000 4930 25034
rect 4930 25000 4964 25034
rect 4964 25000 4998 25034
rect 4998 25000 5032 25034
rect 5032 25000 5066 25034
rect 5066 25000 5100 25034
rect 5100 25000 5134 25034
rect 5134 25000 5168 25034
rect 5168 25000 5202 25034
rect 5202 25000 5236 25034
rect 5236 25000 5270 25034
rect 5270 25000 5304 25034
rect 5304 25000 5338 25034
rect 5338 25000 5372 25034
rect 5372 25000 5406 25034
rect 5406 25000 5440 25034
rect 5440 25000 5474 25034
rect 5474 25000 5508 25034
rect 5508 25000 5542 25034
rect 5542 25000 5576 25034
rect 5576 25000 5610 25034
rect 5610 25000 5644 25034
rect 5644 25000 5678 25034
rect 5678 25000 5712 25034
rect 5712 25000 5746 25034
rect 5746 25000 5780 25034
rect 5780 25000 5814 25034
rect 5814 25000 5848 25034
rect 5848 25000 5882 25034
rect 5882 25000 5916 25034
rect 5916 25000 5950 25034
rect 5950 25000 5984 25034
rect 5984 25000 6018 25034
rect 6018 25000 6052 25034
rect 6052 25000 6086 25034
rect 6086 25000 6120 25034
rect 6120 25000 6154 25034
rect 6154 25000 6188 25034
rect 6188 25000 6222 25034
rect 6222 25000 6256 25034
rect 6256 25000 6290 25034
rect 6290 25000 6324 25034
rect 6324 25000 6358 25034
rect 6358 25000 6392 25034
rect 6392 25000 6426 25034
rect 6426 25000 6460 25034
rect 6460 25000 6494 25034
rect 6494 25000 6528 25034
rect 6528 25000 6562 25034
rect 6562 25000 6596 25034
rect 6596 25000 6630 25034
rect 6630 25000 6664 25034
rect 6664 25000 6698 25034
rect 6698 25000 6732 25034
rect 6732 25000 6766 25034
rect 6766 25000 6800 25034
rect 6800 25000 6834 25034
rect 6834 25000 6868 25034
rect 6868 25000 6902 25034
rect 6902 25000 6936 25034
rect 6936 25000 6970 25034
rect 6970 25000 7004 25034
rect 7004 25000 7038 25034
rect 7038 25000 7072 25034
rect 7072 25000 7106 25034
rect 7106 25000 7140 25034
rect 7140 25000 7174 25034
rect 7174 25000 7208 25034
rect 7208 25000 7242 25034
rect 7242 25000 7276 25034
rect 7276 25000 7310 25034
rect 7310 25000 7344 25034
rect 7344 25000 7378 25034
rect 7378 25000 7412 25034
rect 7412 25000 7446 25034
rect 7446 25000 7480 25034
rect 7480 25000 7514 25034
rect 7514 25000 7548 25034
rect 7548 25000 7582 25034
rect 7582 25000 7616 25034
rect 7616 25000 7650 25034
rect 7650 25000 7684 25034
rect 7684 25000 7718 25034
rect 7718 25000 7752 25034
rect 7752 25000 7786 25034
rect 7786 25000 7820 25034
rect 7820 25000 7854 25034
rect 7854 25000 7888 25034
rect 7888 25000 7922 25034
rect 7922 25000 7956 25034
rect 7956 25000 7990 25034
rect 7990 25000 8024 25034
rect 8024 25000 8058 25034
rect 8058 25000 8092 25034
rect 8092 25000 8126 25034
rect 8126 25000 8160 25034
rect 8160 25000 8194 25034
rect 8194 25000 8228 25034
rect 8228 25000 8262 25034
rect 8262 25000 8296 25034
rect 8296 25000 8330 25034
rect 8330 25000 8364 25034
rect 8364 25000 8398 25034
rect 8398 25000 8432 25034
rect 8432 25000 8466 25034
rect 8466 25000 8500 25034
rect 8500 25000 8534 25034
rect 8534 25000 8568 25034
rect 8568 25000 8602 25034
rect 8602 25000 8636 25034
rect 8636 25000 8670 25034
rect 8670 25000 8704 25034
rect 8704 25000 8738 25034
rect 8738 25000 8772 25034
rect 8772 25000 8806 25034
rect 8806 25000 8840 25034
rect 8840 25000 8874 25034
rect 8874 25000 8908 25034
rect 8908 25000 8942 25034
rect 8942 25000 8976 25034
rect 8976 25000 9010 25034
rect 9010 25000 9044 25034
rect 9044 25000 9078 25034
rect 9078 25000 9112 25034
rect 9112 25000 9146 25034
rect 9146 25000 9180 25034
rect 9180 25000 9214 25034
rect 9214 25000 9248 25034
rect 9248 25000 9282 25034
rect 9282 25000 9316 25034
rect 9316 25000 9350 25034
rect 9350 25000 9384 25034
rect 9384 25000 9418 25034
rect 9418 25000 9452 25034
rect 9452 25000 9486 25034
rect 9486 25000 9520 25034
rect 9520 25000 9554 25034
rect 9554 25000 9588 25034
rect 9588 25000 9622 25034
rect 9622 25000 9656 25034
rect 9656 25000 9690 25034
rect 9690 25000 9724 25034
rect 9724 25000 9758 25034
rect 9758 25000 9792 25034
rect 9792 25000 9826 25034
rect 9826 25000 9860 25034
rect 9860 25000 9894 25034
rect 9894 25000 9928 25034
rect 9928 25000 9962 25034
rect 9962 25000 9996 25034
rect 9996 25000 10030 25034
rect 10030 25000 10064 25034
rect 10064 25000 10098 25034
rect 10098 25000 10132 25034
rect 10132 25000 10166 25034
rect 10166 25000 10200 25034
rect 10200 25000 10234 25034
rect 10234 25000 10268 25034
rect 10268 25000 10302 25034
rect 10302 25000 10336 25034
rect 10336 25000 10370 25034
rect 10370 25000 10404 25034
rect 10404 25000 10438 25034
rect 10438 25000 10472 25034
rect 10472 25000 10506 25034
rect 10506 25000 10540 25034
rect 10540 25000 10574 25034
rect 10574 25000 10608 25034
rect 10608 25000 10642 25034
rect 10642 25000 10676 25034
rect 10676 25000 10710 25034
rect 10710 25000 10744 25034
rect 10744 25000 10778 25034
rect 10778 25000 10812 25034
rect 10812 25000 10846 25034
rect 10846 25000 10880 25034
rect 10880 25000 10914 25034
rect 10914 25000 10948 25034
rect 10948 25000 10982 25034
rect 10982 25000 11016 25034
rect 11016 25000 11050 25034
rect 11050 25000 11084 25034
rect 11084 25000 11118 25034
rect 11118 25000 11152 25034
rect 11152 25000 11186 25034
rect 11186 25000 11220 25034
rect 11220 25000 11254 25034
rect 11254 25000 11288 25034
rect 11288 25000 11322 25034
rect 11322 25000 11356 25034
rect 11356 25000 11390 25034
rect 11390 25000 11424 25034
rect 11424 25000 11458 25034
rect 11458 25000 11492 25034
rect 11492 25000 11526 25034
rect 11526 25000 11560 25034
rect 11560 25000 11594 25034
rect 11594 25000 11628 25034
rect 11628 25000 11662 25034
rect 11662 25000 11696 25034
rect 11696 25000 11730 25034
rect 11730 25000 11764 25034
rect 11764 25000 11798 25034
rect 11798 25000 11832 25034
rect 11832 25000 11866 25034
rect 11866 25000 11900 25034
rect 11900 25000 11934 25034
rect 11934 25000 11968 25034
rect 11968 25000 12002 25034
rect 12002 25000 12036 25034
rect 12036 25000 12070 25034
rect 12070 25000 12104 25034
rect 12104 25000 12138 25034
rect 12138 25000 12172 25034
rect 12172 25000 12206 25034
rect 12206 25000 12240 25034
rect 12240 25000 12274 25034
rect 12274 25000 12308 25034
rect 12308 25000 12342 25034
rect 12342 25000 12376 25034
rect 12376 25000 12410 25034
rect 12410 25000 12444 25034
rect 12444 25000 12478 25034
rect 12478 25000 12512 25034
rect 12512 25000 12546 25034
rect 12546 25000 12580 25034
rect 12580 25000 12614 25034
rect 12614 25000 12648 25034
rect 12648 25000 12682 25034
rect 12682 25000 12716 25034
rect 12716 25000 12750 25034
rect 12750 25000 12784 25034
rect 12784 25000 12818 25034
rect 12818 25000 12852 25034
rect 12852 25000 12886 25034
rect 12886 25000 12920 25034
rect 12920 25000 12954 25034
rect 12954 25000 12988 25034
rect 12988 25000 13022 25034
rect 13022 25000 13056 25034
rect 13056 25000 13090 25034
rect 13090 25000 13124 25034
rect 13124 25000 13158 25034
rect 13158 25000 13192 25034
rect 13192 25000 13226 25034
rect 13226 25000 13260 25034
rect 13260 25000 13294 25034
rect 13294 25000 13328 25034
rect 13328 25000 13362 25034
rect 13362 25000 13396 25034
rect 13396 25000 13430 25034
rect 13430 25000 13464 25034
rect 13464 25000 13498 25034
rect 13498 25000 13532 25034
rect 13532 25000 13566 25034
rect 13566 25000 13600 25034
rect 13600 25000 13634 25034
rect 13634 25000 13668 25034
rect 13668 25000 13702 25034
rect 13702 25000 13736 25034
rect 13736 25000 13770 25034
rect 13770 25000 13804 25034
rect 13804 25000 13838 25034
rect 13838 25000 13872 25034
rect 13872 25000 13906 25034
rect 13906 25000 13940 25034
rect 13940 25000 13974 25034
rect 13974 25000 14008 25034
rect 14008 25000 14042 25034
rect 14042 25000 14076 25034
rect 14076 25000 14110 25034
rect 14110 25000 14144 25034
rect 14144 25000 14178 25034
rect 14178 25000 14212 25034
rect 14212 25000 14246 25034
rect 14246 25000 14280 25034
rect 14280 25000 14314 25034
rect 14314 25000 14348 25034
rect 14348 25000 14382 25034
rect 14382 25000 14416 25034
rect 14416 25000 14450 25034
rect 14450 25000 14484 25034
rect 14484 25000 14518 25034
rect 14518 25000 14552 25034
rect 14552 25000 14586 25034
rect 14586 25000 14620 25034
rect 14620 25000 14654 25034
rect 14654 25000 14688 25034
rect 14688 25000 14722 25034
rect 14722 25000 14756 25034
rect 14756 25000 14790 25034
rect 14790 25000 14824 25034
rect 14824 25000 14858 25034
rect 14858 25000 14870 25034
rect 88 24935 122 24969
rect 161 24962 195 24969
rect 234 24962 268 24969
rect 307 24962 341 24969
rect 380 24962 414 24969
rect 453 24962 487 24969
rect 526 24962 560 24969
rect 599 24962 633 24969
rect 672 24962 706 24969
rect 745 24962 779 24969
rect 818 24962 852 24969
rect 891 24962 925 24969
rect 964 24962 998 24969
rect 1037 24962 1071 24969
rect 1110 24962 1144 24969
rect 1183 24962 1217 24969
rect 1256 24962 1290 24969
rect 1329 24962 1363 24969
rect 1402 24962 1436 24969
rect 1475 24962 1509 24969
rect 1548 24962 1582 24969
rect 1621 24962 1655 24969
rect 1694 24962 1728 24969
rect 1767 24962 1801 24969
rect 1840 24962 1874 24969
rect 1913 24962 1947 24969
rect 1986 24962 2020 24969
rect 2059 24962 2093 24969
rect 2132 24962 2166 24969
rect 2205 24962 2239 24969
rect 161 24935 193 24962
rect 193 24935 195 24962
rect 234 24935 262 24962
rect 262 24935 268 24962
rect 307 24935 331 24962
rect 331 24935 341 24962
rect 380 24935 400 24962
rect 400 24935 414 24962
rect 453 24935 469 24962
rect 469 24935 487 24962
rect 526 24935 538 24962
rect 538 24935 560 24962
rect 599 24935 607 24962
rect 607 24935 633 24962
rect 672 24935 676 24962
rect 676 24935 706 24962
rect 745 24935 779 24962
rect 818 24935 848 24962
rect 848 24935 852 24962
rect 891 24935 917 24962
rect 917 24935 925 24962
rect 964 24935 986 24962
rect 986 24935 998 24962
rect 1037 24935 1054 24962
rect 1054 24935 1071 24962
rect 1110 24935 1122 24962
rect 1122 24935 1144 24962
rect 1183 24935 1190 24962
rect 1190 24935 1217 24962
rect 1256 24935 1258 24962
rect 1258 24935 1290 24962
rect 1329 24935 1360 24962
rect 1360 24935 1363 24962
rect 1402 24935 1428 24962
rect 1428 24935 1436 24962
rect 1475 24935 1496 24962
rect 1496 24935 1509 24962
rect 1548 24935 1564 24962
rect 1564 24935 1582 24962
rect 1621 24935 1632 24962
rect 1632 24935 1655 24962
rect 1694 24935 1700 24962
rect 1700 24935 1728 24962
rect 1767 24935 1768 24962
rect 1768 24935 1801 24962
rect 1840 24935 1870 24962
rect 1870 24935 1874 24962
rect 1913 24935 1938 24962
rect 1938 24935 1947 24962
rect 1986 24935 2006 24962
rect 2006 24935 2020 24962
rect 2059 24935 2074 24962
rect 2074 24935 2093 24962
rect 2132 24935 2142 24962
rect 2142 24935 2166 24962
rect 2205 24935 2210 24962
rect 2210 24935 2239 24962
rect 2278 24935 2312 24969
rect 2351 24962 2385 24969
rect 2424 24962 2458 24969
rect 2497 24962 2531 24969
rect 2570 24962 2604 24969
rect 2643 24962 2677 24969
rect 2716 24962 2750 24969
rect 2789 24962 2823 24969
rect 2862 24962 2896 24969
rect 2935 24962 2969 24969
rect 3008 24962 3042 24969
rect 3081 24962 3115 24969
rect 3154 24962 3188 24969
rect 3227 24962 3261 24969
rect 3300 24962 3334 24969
rect 3373 24962 3407 24969
rect 3446 24962 3480 24969
rect 3519 24962 3553 24969
rect 3592 24962 3626 24969
rect 3665 24962 3699 24969
rect 3738 24962 3772 24969
rect 3811 24962 3845 24969
rect 3884 24962 3918 24969
rect 3957 24962 3991 24969
rect 4030 24962 4064 24969
rect 4103 24962 4137 24969
rect 4176 24962 4210 24969
rect 4249 24962 4283 24969
rect 4322 24962 4356 24969
rect 4395 24962 4429 24969
rect 4468 24962 14870 25000
rect 2351 24935 2380 24962
rect 2380 24935 2385 24962
rect 2424 24935 2448 24962
rect 2448 24935 2458 24962
rect 2497 24935 2516 24962
rect 2516 24935 2531 24962
rect 2570 24935 2584 24962
rect 2584 24935 2604 24962
rect 2643 24935 2652 24962
rect 2652 24935 2677 24962
rect 2716 24935 2720 24962
rect 2720 24935 2750 24962
rect 2789 24935 2822 24962
rect 2822 24935 2823 24962
rect 2862 24935 2890 24962
rect 2890 24935 2896 24962
rect 2935 24935 2958 24962
rect 2958 24935 2969 24962
rect 3008 24935 3026 24962
rect 3026 24935 3042 24962
rect 3081 24935 3094 24962
rect 3094 24935 3115 24962
rect 3154 24935 3162 24962
rect 3162 24935 3188 24962
rect 3227 24935 3230 24962
rect 3230 24935 3261 24962
rect 3300 24935 3332 24962
rect 3332 24935 3334 24962
rect 3373 24935 3400 24962
rect 3400 24935 3407 24962
rect 3446 24935 3468 24962
rect 3468 24935 3480 24962
rect 3519 24935 3536 24962
rect 3536 24935 3553 24962
rect 3592 24935 3604 24962
rect 3604 24935 3626 24962
rect 3665 24935 3672 24962
rect 3672 24935 3699 24962
rect 3738 24935 3740 24962
rect 3740 24935 3772 24962
rect 3811 24935 3842 24962
rect 3842 24935 3845 24962
rect 3884 24935 3910 24962
rect 3910 24935 3918 24962
rect 3957 24935 3978 24962
rect 3978 24935 3991 24962
rect 4030 24935 4046 24962
rect 4046 24935 4064 24962
rect 4103 24935 4114 24962
rect 4114 24935 4137 24962
rect 4176 24935 4182 24962
rect 4182 24935 4210 24962
rect 4249 24935 4250 24962
rect 4250 24935 4283 24962
rect 4322 24935 4352 24962
rect 4352 24935 4356 24962
rect 4395 24935 4420 24962
rect 4420 24935 4429 24962
rect 4468 24928 4488 24962
rect 4488 24928 4522 24962
rect 4522 24928 4556 24962
rect 4556 24928 4590 24962
rect 4590 24928 4624 24962
rect 4624 24928 4658 24962
rect 4658 24928 4692 24962
rect 4692 24928 4726 24962
rect 4726 24928 4760 24962
rect 4760 24928 4794 24962
rect 4794 24928 4828 24962
rect 4828 24928 4862 24962
rect 4862 24928 4896 24962
rect 4896 24928 4930 24962
rect 4930 24928 4964 24962
rect 4964 24928 4998 24962
rect 4998 24928 5032 24962
rect 5032 24928 5066 24962
rect 5066 24928 5100 24962
rect 5100 24928 5134 24962
rect 5134 24928 5168 24962
rect 5168 24928 5202 24962
rect 5202 24928 5236 24962
rect 5236 24928 5270 24962
rect 5270 24928 5304 24962
rect 5304 24928 5338 24962
rect 5338 24928 5372 24962
rect 5372 24928 5406 24962
rect 5406 24928 5440 24962
rect 5440 24928 5474 24962
rect 5474 24928 5508 24962
rect 5508 24928 5542 24962
rect 5542 24928 5576 24962
rect 5576 24928 5610 24962
rect 5610 24928 5644 24962
rect 5644 24928 5678 24962
rect 5678 24928 5712 24962
rect 5712 24928 5746 24962
rect 5746 24928 5780 24962
rect 5780 24928 5814 24962
rect 5814 24928 5848 24962
rect 5848 24928 5882 24962
rect 5882 24928 5916 24962
rect 5916 24928 5950 24962
rect 5950 24928 5984 24962
rect 5984 24928 6018 24962
rect 6018 24928 6052 24962
rect 6052 24928 6086 24962
rect 6086 24928 6120 24962
rect 6120 24928 6154 24962
rect 6154 24928 6188 24962
rect 6188 24928 6222 24962
rect 6222 24928 6256 24962
rect 6256 24928 6290 24962
rect 6290 24928 6324 24962
rect 6324 24928 6358 24962
rect 6358 24928 6392 24962
rect 6392 24928 6426 24962
rect 6426 24928 6460 24962
rect 6460 24928 6494 24962
rect 6494 24928 6528 24962
rect 6528 24928 6562 24962
rect 6562 24928 6596 24962
rect 6596 24928 6630 24962
rect 6630 24928 6664 24962
rect 6664 24928 6698 24962
rect 6698 24928 6732 24962
rect 6732 24928 6766 24962
rect 6766 24928 6800 24962
rect 6800 24928 6834 24962
rect 6834 24928 6868 24962
rect 6868 24928 6902 24962
rect 6902 24928 6936 24962
rect 6936 24928 6970 24962
rect 6970 24928 7004 24962
rect 7004 24928 7038 24962
rect 7038 24928 7072 24962
rect 7072 24928 7106 24962
rect 7106 24928 7140 24962
rect 7140 24928 7174 24962
rect 7174 24928 7208 24962
rect 7208 24928 7242 24962
rect 7242 24928 7276 24962
rect 7276 24928 7310 24962
rect 7310 24928 7344 24962
rect 7344 24928 7378 24962
rect 7378 24928 7412 24962
rect 7412 24928 7446 24962
rect 7446 24928 7480 24962
rect 7480 24928 7514 24962
rect 7514 24928 7548 24962
rect 7548 24928 7582 24962
rect 7582 24928 7616 24962
rect 7616 24928 7650 24962
rect 7650 24928 7684 24962
rect 7684 24928 7718 24962
rect 7718 24928 7752 24962
rect 7752 24928 7786 24962
rect 7786 24928 7820 24962
rect 7820 24928 7854 24962
rect 7854 24928 7888 24962
rect 7888 24928 7922 24962
rect 7922 24928 7956 24962
rect 7956 24928 7990 24962
rect 7990 24928 8024 24962
rect 8024 24928 8058 24962
rect 8058 24928 8092 24962
rect 8092 24928 8126 24962
rect 8126 24928 8160 24962
rect 8160 24928 8194 24962
rect 8194 24928 8228 24962
rect 8228 24928 8262 24962
rect 8262 24928 8296 24962
rect 8296 24928 8330 24962
rect 8330 24928 8364 24962
rect 8364 24928 8398 24962
rect 8398 24928 8432 24962
rect 8432 24928 8466 24962
rect 8466 24928 8500 24962
rect 8500 24928 8534 24962
rect 8534 24928 8568 24962
rect 8568 24928 8602 24962
rect 8602 24928 8636 24962
rect 8636 24928 8670 24962
rect 8670 24928 8704 24962
rect 8704 24928 8738 24962
rect 8738 24928 8772 24962
rect 8772 24928 8806 24962
rect 8806 24928 8840 24962
rect 8840 24928 8874 24962
rect 8874 24928 8908 24962
rect 8908 24928 8942 24962
rect 8942 24928 8976 24962
rect 8976 24928 9010 24962
rect 9010 24928 9044 24962
rect 9044 24928 9078 24962
rect 9078 24928 9112 24962
rect 9112 24928 9146 24962
rect 9146 24928 9180 24962
rect 9180 24928 9214 24962
rect 9214 24928 9248 24962
rect 9248 24928 9282 24962
rect 9282 24928 9316 24962
rect 9316 24928 9350 24962
rect 9350 24928 9384 24962
rect 9384 24928 9418 24962
rect 9418 24928 9452 24962
rect 9452 24928 9486 24962
rect 9486 24928 9520 24962
rect 9520 24928 9554 24962
rect 9554 24928 9588 24962
rect 9588 24928 9622 24962
rect 9622 24928 9656 24962
rect 9656 24928 9690 24962
rect 9690 24928 9724 24962
rect 9724 24928 9758 24962
rect 9758 24928 9792 24962
rect 9792 24928 9826 24962
rect 9826 24928 9860 24962
rect 9860 24928 9894 24962
rect 9894 24928 9928 24962
rect 9928 24928 9962 24962
rect 9962 24928 9996 24962
rect 9996 24928 10030 24962
rect 10030 24928 10064 24962
rect 10064 24928 10098 24962
rect 10098 24928 10132 24962
rect 10132 24928 10166 24962
rect 10166 24928 10200 24962
rect 10200 24928 10234 24962
rect 10234 24928 10268 24962
rect 10268 24928 10302 24962
rect 10302 24928 10336 24962
rect 10336 24928 10370 24962
rect 10370 24928 10404 24962
rect 10404 24928 10438 24962
rect 10438 24928 10472 24962
rect 10472 24928 10506 24962
rect 10506 24928 10540 24962
rect 10540 24928 10574 24962
rect 10574 24928 10608 24962
rect 10608 24928 10642 24962
rect 10642 24928 10676 24962
rect 10676 24928 10710 24962
rect 10710 24928 10744 24962
rect 10744 24928 10778 24962
rect 10778 24928 10812 24962
rect 10812 24928 10846 24962
rect 10846 24928 10880 24962
rect 10880 24928 10914 24962
rect 10914 24928 10948 24962
rect 10948 24928 10982 24962
rect 10982 24928 11016 24962
rect 11016 24928 11050 24962
rect 11050 24928 11084 24962
rect 11084 24928 11118 24962
rect 11118 24928 11152 24962
rect 11152 24928 11186 24962
rect 11186 24928 11220 24962
rect 11220 24928 11254 24962
rect 11254 24928 11288 24962
rect 11288 24928 11322 24962
rect 11322 24928 11356 24962
rect 11356 24928 11390 24962
rect 11390 24928 11424 24962
rect 11424 24928 11458 24962
rect 11458 24928 11492 24962
rect 11492 24928 11526 24962
rect 11526 24928 11560 24962
rect 11560 24928 11594 24962
rect 11594 24928 11628 24962
rect 11628 24928 11662 24962
rect 11662 24928 11696 24962
rect 11696 24928 11730 24962
rect 11730 24928 11764 24962
rect 11764 24928 11798 24962
rect 11798 24928 11832 24962
rect 11832 24928 11866 24962
rect 11866 24928 11900 24962
rect 11900 24928 11934 24962
rect 11934 24928 11968 24962
rect 11968 24928 12002 24962
rect 12002 24928 12036 24962
rect 12036 24928 12070 24962
rect 12070 24928 12104 24962
rect 12104 24928 12138 24962
rect 12138 24928 12172 24962
rect 12172 24928 12206 24962
rect 12206 24928 12240 24962
rect 12240 24928 12274 24962
rect 12274 24928 12308 24962
rect 12308 24928 12342 24962
rect 12342 24928 12376 24962
rect 12376 24928 12410 24962
rect 12410 24928 12444 24962
rect 12444 24928 12478 24962
rect 12478 24928 12512 24962
rect 12512 24928 12546 24962
rect 12546 24928 12580 24962
rect 12580 24928 12614 24962
rect 12614 24928 12648 24962
rect 12648 24928 12682 24962
rect 12682 24928 12716 24962
rect 12716 24928 12750 24962
rect 12750 24928 12784 24962
rect 12784 24928 12818 24962
rect 12818 24928 12852 24962
rect 12852 24928 12886 24962
rect 12886 24928 12920 24962
rect 12920 24928 12954 24962
rect 12954 24928 12988 24962
rect 12988 24928 13022 24962
rect 13022 24928 13056 24962
rect 13056 24928 13090 24962
rect 13090 24928 13124 24962
rect 13124 24928 13158 24962
rect 13158 24928 13192 24962
rect 13192 24928 13226 24962
rect 13226 24928 13260 24962
rect 13260 24928 13294 24962
rect 13294 24928 13328 24962
rect 13328 24928 13362 24962
rect 13362 24928 13396 24962
rect 13396 24928 13430 24962
rect 13430 24928 13464 24962
rect 13464 24928 13498 24962
rect 13498 24928 13532 24962
rect 13532 24928 13566 24962
rect 13566 24928 13600 24962
rect 13600 24928 13634 24962
rect 13634 24928 13668 24962
rect 13668 24928 13702 24962
rect 13702 24928 13736 24962
rect 13736 24928 13770 24962
rect 13770 24928 13804 24962
rect 13804 24928 13838 24962
rect 13838 24928 13872 24962
rect 13872 24928 13906 24962
rect 13906 24928 13940 24962
rect 13940 24928 13974 24962
rect 13974 24928 14008 24962
rect 14008 24928 14042 24962
rect 14042 24928 14076 24962
rect 14076 24928 14110 24962
rect 14110 24928 14144 24962
rect 14144 24928 14178 24962
rect 14178 24928 14212 24962
rect 14212 24928 14246 24962
rect 14246 24928 14280 24962
rect 14280 24928 14314 24962
rect 14314 24928 14348 24962
rect 14348 24928 14382 24962
rect 14382 24928 14416 24962
rect 14416 24928 14450 24962
rect 14450 24928 14484 24962
rect 14484 24928 14518 24962
rect 14518 24928 14552 24962
rect 14552 24928 14586 24962
rect 14586 24928 14620 24962
rect 14620 24928 14654 24962
rect 14654 24928 14688 24962
rect 14688 24928 14722 24962
rect 14722 24928 14756 24962
rect 14756 24928 14790 24962
rect 14790 24928 14824 24962
rect 14824 24928 14858 24962
rect 14858 24928 14870 24962
rect 88 24863 122 24897
rect 161 24890 195 24897
rect 234 24890 268 24897
rect 307 24890 341 24897
rect 380 24890 414 24897
rect 453 24890 487 24897
rect 526 24890 560 24897
rect 599 24890 633 24897
rect 672 24890 706 24897
rect 745 24890 779 24897
rect 818 24890 852 24897
rect 891 24890 925 24897
rect 964 24890 998 24897
rect 1037 24890 1071 24897
rect 1110 24890 1144 24897
rect 1183 24890 1217 24897
rect 1256 24890 1290 24897
rect 1329 24890 1363 24897
rect 1402 24890 1436 24897
rect 1475 24890 1509 24897
rect 1548 24890 1582 24897
rect 1621 24890 1655 24897
rect 1694 24890 1728 24897
rect 1767 24890 1801 24897
rect 1840 24890 1874 24897
rect 1913 24890 1947 24897
rect 1986 24890 2020 24897
rect 2059 24890 2093 24897
rect 2132 24890 2166 24897
rect 2205 24890 2239 24897
rect 161 24863 193 24890
rect 193 24863 195 24890
rect 234 24863 262 24890
rect 262 24863 268 24890
rect 307 24863 331 24890
rect 331 24863 341 24890
rect 380 24863 400 24890
rect 400 24863 414 24890
rect 453 24863 469 24890
rect 469 24863 487 24890
rect 526 24863 538 24890
rect 538 24863 560 24890
rect 599 24863 607 24890
rect 607 24863 633 24890
rect 672 24863 676 24890
rect 676 24863 706 24890
rect 745 24863 779 24890
rect 818 24863 848 24890
rect 848 24863 852 24890
rect 891 24863 917 24890
rect 917 24863 925 24890
rect 964 24863 986 24890
rect 986 24863 998 24890
rect 1037 24863 1054 24890
rect 1054 24863 1071 24890
rect 1110 24863 1122 24890
rect 1122 24863 1144 24890
rect 1183 24863 1190 24890
rect 1190 24863 1217 24890
rect 1256 24863 1258 24890
rect 1258 24863 1290 24890
rect 1329 24863 1360 24890
rect 1360 24863 1363 24890
rect 1402 24863 1428 24890
rect 1428 24863 1436 24890
rect 1475 24863 1496 24890
rect 1496 24863 1509 24890
rect 1548 24863 1564 24890
rect 1564 24863 1582 24890
rect 1621 24863 1632 24890
rect 1632 24863 1655 24890
rect 1694 24863 1700 24890
rect 1700 24863 1728 24890
rect 1767 24863 1768 24890
rect 1768 24863 1801 24890
rect 1840 24863 1870 24890
rect 1870 24863 1874 24890
rect 1913 24863 1938 24890
rect 1938 24863 1947 24890
rect 1986 24863 2006 24890
rect 2006 24863 2020 24890
rect 2059 24863 2074 24890
rect 2074 24863 2093 24890
rect 2132 24863 2142 24890
rect 2142 24863 2166 24890
rect 2205 24863 2210 24890
rect 2210 24863 2239 24890
rect 2278 24863 2312 24897
rect 2351 24890 2385 24897
rect 2424 24890 2458 24897
rect 2497 24890 2531 24897
rect 2570 24890 2604 24897
rect 2643 24890 2677 24897
rect 2716 24890 2750 24897
rect 2789 24890 2823 24897
rect 2862 24890 2896 24897
rect 2935 24890 2969 24897
rect 3008 24890 3042 24897
rect 3081 24890 3115 24897
rect 3154 24890 3188 24897
rect 3227 24890 3261 24897
rect 3300 24890 3334 24897
rect 3373 24890 3407 24897
rect 3446 24890 3480 24897
rect 3519 24890 3553 24897
rect 3592 24890 3626 24897
rect 3665 24890 3699 24897
rect 3738 24890 3772 24897
rect 3811 24890 3845 24897
rect 3884 24890 3918 24897
rect 3957 24890 3991 24897
rect 4030 24890 4064 24897
rect 4103 24890 4137 24897
rect 4176 24890 4210 24897
rect 4249 24890 4283 24897
rect 4322 24890 4356 24897
rect 4395 24890 4429 24897
rect 4468 24890 14870 24928
rect 2351 24863 2380 24890
rect 2380 24863 2385 24890
rect 2424 24863 2448 24890
rect 2448 24863 2458 24890
rect 2497 24863 2516 24890
rect 2516 24863 2531 24890
rect 2570 24863 2584 24890
rect 2584 24863 2604 24890
rect 2643 24863 2652 24890
rect 2652 24863 2677 24890
rect 2716 24863 2720 24890
rect 2720 24863 2750 24890
rect 2789 24863 2822 24890
rect 2822 24863 2823 24890
rect 2862 24863 2890 24890
rect 2890 24863 2896 24890
rect 2935 24863 2958 24890
rect 2958 24863 2969 24890
rect 3008 24863 3026 24890
rect 3026 24863 3042 24890
rect 3081 24863 3094 24890
rect 3094 24863 3115 24890
rect 3154 24863 3162 24890
rect 3162 24863 3188 24890
rect 3227 24863 3230 24890
rect 3230 24863 3261 24890
rect 3300 24863 3332 24890
rect 3332 24863 3334 24890
rect 3373 24863 3400 24890
rect 3400 24863 3407 24890
rect 3446 24863 3468 24890
rect 3468 24863 3480 24890
rect 3519 24863 3536 24890
rect 3536 24863 3553 24890
rect 3592 24863 3604 24890
rect 3604 24863 3626 24890
rect 3665 24863 3672 24890
rect 3672 24863 3699 24890
rect 3738 24863 3740 24890
rect 3740 24863 3772 24890
rect 3811 24863 3842 24890
rect 3842 24863 3845 24890
rect 3884 24863 3910 24890
rect 3910 24863 3918 24890
rect 3957 24863 3978 24890
rect 3978 24863 3991 24890
rect 4030 24863 4046 24890
rect 4046 24863 4064 24890
rect 4103 24863 4114 24890
rect 4114 24863 4137 24890
rect 4176 24863 4182 24890
rect 4182 24863 4210 24890
rect 4249 24863 4250 24890
rect 4250 24863 4283 24890
rect 4322 24863 4352 24890
rect 4352 24863 4356 24890
rect 4395 24863 4420 24890
rect 4420 24863 4429 24890
rect 4468 24856 4488 24890
rect 4488 24856 4522 24890
rect 4522 24856 4556 24890
rect 4556 24856 4590 24890
rect 4590 24856 4624 24890
rect 4624 24856 4658 24890
rect 4658 24856 4692 24890
rect 4692 24856 4726 24890
rect 4726 24856 4760 24890
rect 4760 24856 4794 24890
rect 4794 24856 4828 24890
rect 4828 24856 4862 24890
rect 4862 24856 4896 24890
rect 4896 24856 4930 24890
rect 4930 24856 4964 24890
rect 4964 24856 4998 24890
rect 4998 24856 5032 24890
rect 5032 24856 5066 24890
rect 5066 24856 5100 24890
rect 5100 24856 5134 24890
rect 5134 24856 5168 24890
rect 5168 24856 5202 24890
rect 5202 24856 5236 24890
rect 5236 24856 5270 24890
rect 5270 24856 5304 24890
rect 5304 24856 5338 24890
rect 5338 24856 5372 24890
rect 5372 24856 5406 24890
rect 5406 24856 5440 24890
rect 5440 24856 5474 24890
rect 5474 24856 5508 24890
rect 5508 24856 5542 24890
rect 5542 24856 5576 24890
rect 5576 24856 5610 24890
rect 5610 24856 5644 24890
rect 5644 24856 5678 24890
rect 5678 24856 5712 24890
rect 5712 24856 5746 24890
rect 5746 24856 5780 24890
rect 5780 24856 5814 24890
rect 5814 24856 5848 24890
rect 5848 24856 5882 24890
rect 5882 24856 5916 24890
rect 5916 24856 5950 24890
rect 5950 24856 5984 24890
rect 5984 24856 6018 24890
rect 6018 24856 6052 24890
rect 6052 24856 6086 24890
rect 6086 24856 6120 24890
rect 6120 24856 6154 24890
rect 6154 24856 6188 24890
rect 6188 24856 6222 24890
rect 6222 24856 6256 24890
rect 6256 24856 6290 24890
rect 6290 24856 6324 24890
rect 6324 24856 6358 24890
rect 6358 24856 6392 24890
rect 6392 24856 6426 24890
rect 6426 24856 6460 24890
rect 6460 24856 6494 24890
rect 6494 24856 6528 24890
rect 6528 24856 6562 24890
rect 6562 24856 6596 24890
rect 6596 24856 6630 24890
rect 6630 24856 6664 24890
rect 6664 24856 6698 24890
rect 6698 24856 6732 24890
rect 6732 24856 6766 24890
rect 6766 24856 6800 24890
rect 6800 24856 6834 24890
rect 6834 24856 6868 24890
rect 6868 24856 6902 24890
rect 6902 24856 6936 24890
rect 6936 24856 6970 24890
rect 6970 24856 7004 24890
rect 7004 24856 7038 24890
rect 7038 24856 7072 24890
rect 7072 24856 7106 24890
rect 7106 24856 7140 24890
rect 7140 24856 7174 24890
rect 7174 24856 7208 24890
rect 7208 24856 7242 24890
rect 7242 24856 7276 24890
rect 7276 24856 7310 24890
rect 7310 24856 7344 24890
rect 7344 24856 7378 24890
rect 7378 24856 7412 24890
rect 7412 24856 7446 24890
rect 7446 24856 7480 24890
rect 7480 24856 7514 24890
rect 7514 24856 7548 24890
rect 7548 24856 7582 24890
rect 7582 24856 7616 24890
rect 7616 24856 7650 24890
rect 7650 24856 7684 24890
rect 7684 24856 7718 24890
rect 7718 24856 7752 24890
rect 7752 24856 7786 24890
rect 7786 24856 7820 24890
rect 7820 24856 7854 24890
rect 7854 24856 7888 24890
rect 7888 24856 7922 24890
rect 7922 24856 7956 24890
rect 7956 24856 7990 24890
rect 7990 24856 8024 24890
rect 8024 24856 8058 24890
rect 8058 24856 8092 24890
rect 8092 24856 8126 24890
rect 8126 24856 8160 24890
rect 8160 24856 8194 24890
rect 8194 24856 8228 24890
rect 8228 24856 8262 24890
rect 8262 24856 8296 24890
rect 8296 24856 8330 24890
rect 8330 24856 8364 24890
rect 8364 24856 8398 24890
rect 8398 24856 8432 24890
rect 8432 24856 8466 24890
rect 8466 24856 8500 24890
rect 8500 24856 8534 24890
rect 8534 24856 8568 24890
rect 8568 24856 8602 24890
rect 8602 24856 8636 24890
rect 8636 24856 8670 24890
rect 8670 24856 8704 24890
rect 8704 24856 8738 24890
rect 8738 24856 8772 24890
rect 8772 24856 8806 24890
rect 8806 24856 8840 24890
rect 8840 24856 8874 24890
rect 8874 24856 8908 24890
rect 8908 24856 8942 24890
rect 8942 24856 8976 24890
rect 8976 24856 9010 24890
rect 9010 24856 9044 24890
rect 9044 24856 9078 24890
rect 9078 24856 9112 24890
rect 9112 24856 9146 24890
rect 9146 24856 9180 24890
rect 9180 24856 9214 24890
rect 9214 24856 9248 24890
rect 9248 24856 9282 24890
rect 9282 24856 9316 24890
rect 9316 24856 9350 24890
rect 9350 24856 9384 24890
rect 9384 24856 9418 24890
rect 9418 24856 9452 24890
rect 9452 24856 9486 24890
rect 9486 24856 9520 24890
rect 9520 24856 9554 24890
rect 9554 24856 9588 24890
rect 9588 24856 9622 24890
rect 9622 24856 9656 24890
rect 9656 24856 9690 24890
rect 9690 24856 9724 24890
rect 9724 24856 9758 24890
rect 9758 24856 9792 24890
rect 9792 24856 9826 24890
rect 9826 24856 9860 24890
rect 9860 24856 9894 24890
rect 9894 24856 9928 24890
rect 9928 24856 9962 24890
rect 9962 24856 9996 24890
rect 9996 24856 10030 24890
rect 10030 24856 10064 24890
rect 10064 24856 10098 24890
rect 10098 24856 10132 24890
rect 10132 24856 10166 24890
rect 10166 24856 10200 24890
rect 10200 24856 10234 24890
rect 10234 24856 10268 24890
rect 10268 24856 10302 24890
rect 10302 24856 10336 24890
rect 10336 24856 10370 24890
rect 10370 24856 10404 24890
rect 10404 24856 10438 24890
rect 10438 24856 10472 24890
rect 10472 24856 10506 24890
rect 10506 24856 10540 24890
rect 10540 24856 10574 24890
rect 10574 24856 10608 24890
rect 10608 24856 10642 24890
rect 10642 24856 10676 24890
rect 10676 24856 10710 24890
rect 10710 24856 10744 24890
rect 10744 24856 10778 24890
rect 10778 24856 10812 24890
rect 10812 24856 10846 24890
rect 10846 24856 10880 24890
rect 10880 24856 10914 24890
rect 10914 24856 10948 24890
rect 10948 24856 10982 24890
rect 10982 24856 11016 24890
rect 11016 24856 11050 24890
rect 11050 24856 11084 24890
rect 11084 24856 11118 24890
rect 11118 24856 11152 24890
rect 11152 24856 11186 24890
rect 11186 24856 11220 24890
rect 11220 24856 11254 24890
rect 11254 24856 11288 24890
rect 11288 24856 11322 24890
rect 11322 24856 11356 24890
rect 11356 24856 11390 24890
rect 11390 24856 11424 24890
rect 11424 24856 11458 24890
rect 11458 24856 11492 24890
rect 11492 24856 11526 24890
rect 11526 24856 11560 24890
rect 11560 24856 11594 24890
rect 11594 24856 11628 24890
rect 11628 24856 11662 24890
rect 11662 24856 11696 24890
rect 11696 24856 11730 24890
rect 11730 24856 11764 24890
rect 11764 24856 11798 24890
rect 11798 24856 11832 24890
rect 11832 24856 11866 24890
rect 11866 24856 11900 24890
rect 11900 24856 11934 24890
rect 11934 24856 11968 24890
rect 11968 24856 12002 24890
rect 12002 24856 12036 24890
rect 12036 24856 12070 24890
rect 12070 24856 12104 24890
rect 12104 24856 12138 24890
rect 12138 24856 12172 24890
rect 12172 24856 12206 24890
rect 12206 24856 12240 24890
rect 12240 24856 12274 24890
rect 12274 24856 12308 24890
rect 12308 24856 12342 24890
rect 12342 24856 12376 24890
rect 12376 24856 12410 24890
rect 12410 24856 12444 24890
rect 12444 24856 12478 24890
rect 12478 24856 12512 24890
rect 12512 24856 12546 24890
rect 12546 24856 12580 24890
rect 12580 24856 12614 24890
rect 12614 24856 12648 24890
rect 12648 24856 12682 24890
rect 12682 24856 12716 24890
rect 12716 24856 12750 24890
rect 12750 24856 12784 24890
rect 12784 24856 12818 24890
rect 12818 24856 12852 24890
rect 12852 24856 12886 24890
rect 12886 24856 12920 24890
rect 12920 24856 12954 24890
rect 12954 24856 12988 24890
rect 12988 24856 13022 24890
rect 13022 24856 13056 24890
rect 13056 24856 13090 24890
rect 13090 24856 13124 24890
rect 13124 24856 13158 24890
rect 13158 24856 13192 24890
rect 13192 24856 13226 24890
rect 13226 24856 13260 24890
rect 13260 24856 13294 24890
rect 13294 24856 13328 24890
rect 13328 24856 13362 24890
rect 13362 24856 13396 24890
rect 13396 24856 13430 24890
rect 13430 24856 13464 24890
rect 13464 24856 13498 24890
rect 13498 24856 13532 24890
rect 13532 24856 13566 24890
rect 13566 24856 13600 24890
rect 13600 24856 13634 24890
rect 13634 24856 13668 24890
rect 13668 24856 13702 24890
rect 13702 24856 13736 24890
rect 13736 24856 13770 24890
rect 13770 24856 13804 24890
rect 13804 24856 13838 24890
rect 13838 24856 13872 24890
rect 13872 24856 13906 24890
rect 13906 24856 13940 24890
rect 13940 24856 13974 24890
rect 13974 24856 14008 24890
rect 14008 24856 14042 24890
rect 14042 24856 14076 24890
rect 14076 24856 14110 24890
rect 14110 24856 14144 24890
rect 14144 24856 14178 24890
rect 14178 24856 14212 24890
rect 14212 24856 14246 24890
rect 14246 24856 14280 24890
rect 14280 24856 14314 24890
rect 14314 24856 14348 24890
rect 14348 24856 14382 24890
rect 14382 24856 14416 24890
rect 14416 24856 14450 24890
rect 14450 24856 14484 24890
rect 14484 24856 14518 24890
rect 14518 24856 14552 24890
rect 14552 24856 14586 24890
rect 14586 24856 14620 24890
rect 14620 24856 14654 24890
rect 14654 24856 14688 24890
rect 14688 24856 14722 24890
rect 14722 24856 14756 24890
rect 14756 24856 14790 24890
rect 14790 24856 14824 24890
rect 14824 24856 14858 24890
rect 14858 24856 14870 24890
rect 88 24791 122 24825
rect 161 24818 195 24825
rect 234 24818 268 24825
rect 307 24818 341 24825
rect 380 24818 414 24825
rect 453 24818 487 24825
rect 526 24818 560 24825
rect 599 24818 633 24825
rect 672 24818 706 24825
rect 745 24818 779 24825
rect 818 24818 852 24825
rect 891 24818 925 24825
rect 964 24818 998 24825
rect 1037 24818 1071 24825
rect 1110 24818 1144 24825
rect 1183 24818 1217 24825
rect 1256 24818 1290 24825
rect 1329 24818 1363 24825
rect 1402 24818 1436 24825
rect 1475 24818 1509 24825
rect 1548 24818 1582 24825
rect 1621 24818 1655 24825
rect 1694 24818 1728 24825
rect 1767 24818 1801 24825
rect 1840 24818 1874 24825
rect 1913 24818 1947 24825
rect 1986 24818 2020 24825
rect 2059 24818 2093 24825
rect 2132 24818 2166 24825
rect 2205 24818 2239 24825
rect 161 24791 193 24818
rect 193 24791 195 24818
rect 234 24791 262 24818
rect 262 24791 268 24818
rect 307 24791 331 24818
rect 331 24791 341 24818
rect 380 24791 400 24818
rect 400 24791 414 24818
rect 453 24791 469 24818
rect 469 24791 487 24818
rect 526 24791 538 24818
rect 538 24791 560 24818
rect 599 24791 607 24818
rect 607 24791 633 24818
rect 672 24791 676 24818
rect 676 24791 706 24818
rect 745 24791 779 24818
rect 818 24791 848 24818
rect 848 24791 852 24818
rect 891 24791 917 24818
rect 917 24791 925 24818
rect 964 24791 986 24818
rect 986 24791 998 24818
rect 1037 24791 1054 24818
rect 1054 24791 1071 24818
rect 1110 24791 1122 24818
rect 1122 24791 1144 24818
rect 1183 24791 1190 24818
rect 1190 24791 1217 24818
rect 1256 24791 1258 24818
rect 1258 24791 1290 24818
rect 1329 24791 1360 24818
rect 1360 24791 1363 24818
rect 1402 24791 1428 24818
rect 1428 24791 1436 24818
rect 1475 24791 1496 24818
rect 1496 24791 1509 24818
rect 1548 24791 1564 24818
rect 1564 24791 1582 24818
rect 1621 24791 1632 24818
rect 1632 24791 1655 24818
rect 1694 24791 1700 24818
rect 1700 24791 1728 24818
rect 1767 24791 1768 24818
rect 1768 24791 1801 24818
rect 1840 24791 1870 24818
rect 1870 24791 1874 24818
rect 1913 24791 1938 24818
rect 1938 24791 1947 24818
rect 1986 24791 2006 24818
rect 2006 24791 2020 24818
rect 2059 24791 2074 24818
rect 2074 24791 2093 24818
rect 2132 24791 2142 24818
rect 2142 24791 2166 24818
rect 2205 24791 2210 24818
rect 2210 24791 2239 24818
rect 2278 24791 2312 24825
rect 2351 24818 2385 24825
rect 2424 24818 2458 24825
rect 2497 24818 2531 24825
rect 2570 24818 2604 24825
rect 2643 24818 2677 24825
rect 2716 24818 2750 24825
rect 2789 24818 2823 24825
rect 2862 24818 2896 24825
rect 2935 24818 2969 24825
rect 3008 24818 3042 24825
rect 3081 24818 3115 24825
rect 3154 24818 3188 24825
rect 3227 24818 3261 24825
rect 3300 24818 3334 24825
rect 3373 24818 3407 24825
rect 3446 24818 3480 24825
rect 3519 24818 3553 24825
rect 3592 24818 3626 24825
rect 3665 24818 3699 24825
rect 3738 24818 3772 24825
rect 3811 24818 3845 24825
rect 3884 24818 3918 24825
rect 3957 24818 3991 24825
rect 4030 24818 4064 24825
rect 4103 24818 4137 24825
rect 4176 24818 4210 24825
rect 4249 24818 4283 24825
rect 4322 24818 4356 24825
rect 4395 24818 4429 24825
rect 4468 24818 14870 24856
rect 2351 24791 2380 24818
rect 2380 24791 2385 24818
rect 2424 24791 2448 24818
rect 2448 24791 2458 24818
rect 2497 24791 2516 24818
rect 2516 24791 2531 24818
rect 2570 24791 2584 24818
rect 2584 24791 2604 24818
rect 2643 24791 2652 24818
rect 2652 24791 2677 24818
rect 2716 24791 2720 24818
rect 2720 24791 2750 24818
rect 2789 24791 2822 24818
rect 2822 24791 2823 24818
rect 2862 24791 2890 24818
rect 2890 24791 2896 24818
rect 2935 24791 2958 24818
rect 2958 24791 2969 24818
rect 3008 24791 3026 24818
rect 3026 24791 3042 24818
rect 3081 24791 3094 24818
rect 3094 24791 3115 24818
rect 3154 24791 3162 24818
rect 3162 24791 3188 24818
rect 3227 24791 3230 24818
rect 3230 24791 3261 24818
rect 3300 24791 3332 24818
rect 3332 24791 3334 24818
rect 3373 24791 3400 24818
rect 3400 24791 3407 24818
rect 3446 24791 3468 24818
rect 3468 24791 3480 24818
rect 3519 24791 3536 24818
rect 3536 24791 3553 24818
rect 3592 24791 3604 24818
rect 3604 24791 3626 24818
rect 3665 24791 3672 24818
rect 3672 24791 3699 24818
rect 3738 24791 3740 24818
rect 3740 24791 3772 24818
rect 3811 24791 3842 24818
rect 3842 24791 3845 24818
rect 3884 24791 3910 24818
rect 3910 24791 3918 24818
rect 3957 24791 3978 24818
rect 3978 24791 3991 24818
rect 4030 24791 4046 24818
rect 4046 24791 4064 24818
rect 4103 24791 4114 24818
rect 4114 24791 4137 24818
rect 4176 24791 4182 24818
rect 4182 24791 4210 24818
rect 4249 24791 4250 24818
rect 4250 24791 4283 24818
rect 4322 24791 4352 24818
rect 4352 24791 4356 24818
rect 4395 24791 4420 24818
rect 4420 24791 4429 24818
rect 4468 24784 4488 24818
rect 4488 24784 4522 24818
rect 4522 24784 4556 24818
rect 4556 24784 4590 24818
rect 4590 24784 4624 24818
rect 4624 24784 4658 24818
rect 4658 24784 4692 24818
rect 4692 24784 4726 24818
rect 4726 24784 4760 24818
rect 4760 24784 4794 24818
rect 4794 24784 4828 24818
rect 4828 24784 4862 24818
rect 4862 24784 4896 24818
rect 4896 24784 4930 24818
rect 4930 24784 4964 24818
rect 4964 24784 4998 24818
rect 4998 24784 5032 24818
rect 5032 24784 5066 24818
rect 5066 24784 5100 24818
rect 5100 24784 5134 24818
rect 5134 24784 5168 24818
rect 5168 24784 5202 24818
rect 5202 24784 5236 24818
rect 5236 24784 5270 24818
rect 5270 24784 5304 24818
rect 5304 24784 5338 24818
rect 5338 24784 5372 24818
rect 5372 24784 5406 24818
rect 5406 24784 5440 24818
rect 5440 24784 5474 24818
rect 5474 24784 5508 24818
rect 5508 24784 5542 24818
rect 5542 24784 5576 24818
rect 5576 24784 5610 24818
rect 5610 24784 5644 24818
rect 5644 24784 5678 24818
rect 5678 24784 5712 24818
rect 5712 24784 5746 24818
rect 5746 24784 5780 24818
rect 5780 24784 5814 24818
rect 5814 24784 5848 24818
rect 5848 24784 5882 24818
rect 5882 24784 5916 24818
rect 5916 24784 5950 24818
rect 5950 24784 5984 24818
rect 5984 24784 6018 24818
rect 6018 24784 6052 24818
rect 6052 24784 6086 24818
rect 6086 24784 6120 24818
rect 6120 24784 6154 24818
rect 6154 24784 6188 24818
rect 6188 24784 6222 24818
rect 6222 24784 6256 24818
rect 6256 24784 6290 24818
rect 6290 24784 6324 24818
rect 6324 24784 6358 24818
rect 6358 24784 6392 24818
rect 6392 24784 6426 24818
rect 6426 24784 6460 24818
rect 6460 24784 6494 24818
rect 6494 24784 6528 24818
rect 6528 24784 6562 24818
rect 6562 24784 6596 24818
rect 6596 24784 6630 24818
rect 6630 24784 6664 24818
rect 6664 24784 6698 24818
rect 6698 24784 6732 24818
rect 6732 24784 6766 24818
rect 6766 24784 6800 24818
rect 6800 24784 6834 24818
rect 6834 24784 6868 24818
rect 6868 24784 6902 24818
rect 6902 24784 6936 24818
rect 6936 24784 6970 24818
rect 6970 24784 7004 24818
rect 7004 24784 7038 24818
rect 7038 24784 7072 24818
rect 7072 24784 7106 24818
rect 7106 24784 7140 24818
rect 7140 24784 7174 24818
rect 7174 24784 7208 24818
rect 7208 24784 7242 24818
rect 7242 24784 7276 24818
rect 7276 24784 7310 24818
rect 7310 24784 7344 24818
rect 7344 24784 7378 24818
rect 7378 24784 7412 24818
rect 7412 24784 7446 24818
rect 7446 24784 7480 24818
rect 7480 24784 7514 24818
rect 7514 24784 7548 24818
rect 7548 24784 7582 24818
rect 7582 24784 7616 24818
rect 7616 24784 7650 24818
rect 7650 24784 7684 24818
rect 7684 24784 7718 24818
rect 7718 24784 7752 24818
rect 7752 24784 7786 24818
rect 7786 24784 7820 24818
rect 7820 24784 7854 24818
rect 7854 24784 7888 24818
rect 7888 24784 7922 24818
rect 7922 24784 7956 24818
rect 7956 24784 7990 24818
rect 7990 24784 8024 24818
rect 8024 24784 8058 24818
rect 8058 24784 8092 24818
rect 8092 24784 8126 24818
rect 8126 24784 8160 24818
rect 8160 24784 8194 24818
rect 8194 24784 8228 24818
rect 8228 24784 8262 24818
rect 8262 24784 8296 24818
rect 8296 24784 8330 24818
rect 8330 24784 8364 24818
rect 8364 24784 8398 24818
rect 8398 24784 8432 24818
rect 8432 24784 8466 24818
rect 8466 24784 8500 24818
rect 8500 24784 8534 24818
rect 8534 24784 8568 24818
rect 8568 24784 8602 24818
rect 8602 24784 8636 24818
rect 8636 24784 8670 24818
rect 8670 24784 8704 24818
rect 8704 24784 8738 24818
rect 8738 24784 8772 24818
rect 8772 24784 8806 24818
rect 8806 24784 8840 24818
rect 8840 24784 8874 24818
rect 8874 24784 8908 24818
rect 8908 24784 8942 24818
rect 8942 24784 8976 24818
rect 8976 24784 9010 24818
rect 9010 24784 9044 24818
rect 9044 24784 9078 24818
rect 9078 24784 9112 24818
rect 9112 24784 9146 24818
rect 9146 24784 9180 24818
rect 9180 24784 9214 24818
rect 9214 24784 9248 24818
rect 9248 24784 9282 24818
rect 9282 24784 9316 24818
rect 9316 24784 9350 24818
rect 9350 24784 9384 24818
rect 9384 24784 9418 24818
rect 9418 24784 9452 24818
rect 9452 24784 9486 24818
rect 9486 24784 9520 24818
rect 9520 24784 9554 24818
rect 9554 24784 9588 24818
rect 9588 24784 9622 24818
rect 9622 24784 9656 24818
rect 9656 24784 9690 24818
rect 9690 24784 9724 24818
rect 9724 24784 9758 24818
rect 9758 24784 9792 24818
rect 9792 24784 9826 24818
rect 9826 24784 9860 24818
rect 9860 24784 9894 24818
rect 9894 24784 9928 24818
rect 9928 24784 9962 24818
rect 9962 24784 9996 24818
rect 9996 24784 10030 24818
rect 10030 24784 10064 24818
rect 10064 24784 10098 24818
rect 10098 24784 10132 24818
rect 10132 24784 10166 24818
rect 10166 24784 10200 24818
rect 10200 24784 10234 24818
rect 10234 24784 10268 24818
rect 10268 24784 10302 24818
rect 10302 24784 10336 24818
rect 10336 24784 10370 24818
rect 10370 24784 10404 24818
rect 10404 24784 10438 24818
rect 10438 24784 10472 24818
rect 10472 24784 10506 24818
rect 10506 24784 10540 24818
rect 10540 24784 10574 24818
rect 10574 24784 10608 24818
rect 10608 24784 10642 24818
rect 10642 24784 10676 24818
rect 10676 24784 10710 24818
rect 10710 24784 10744 24818
rect 10744 24784 10778 24818
rect 10778 24784 10812 24818
rect 10812 24784 10846 24818
rect 10846 24784 10880 24818
rect 10880 24784 10914 24818
rect 10914 24784 10948 24818
rect 10948 24784 10982 24818
rect 10982 24784 11016 24818
rect 11016 24784 11050 24818
rect 11050 24784 11084 24818
rect 11084 24784 11118 24818
rect 11118 24784 11152 24818
rect 11152 24784 11186 24818
rect 11186 24784 11220 24818
rect 11220 24784 11254 24818
rect 11254 24784 11288 24818
rect 11288 24784 11322 24818
rect 11322 24784 11356 24818
rect 11356 24784 11390 24818
rect 11390 24784 11424 24818
rect 11424 24784 11458 24818
rect 11458 24784 11492 24818
rect 11492 24784 11526 24818
rect 11526 24784 11560 24818
rect 11560 24784 11594 24818
rect 11594 24784 11628 24818
rect 11628 24784 11662 24818
rect 11662 24784 11696 24818
rect 11696 24784 11730 24818
rect 11730 24784 11764 24818
rect 11764 24784 11798 24818
rect 11798 24784 11832 24818
rect 11832 24784 11866 24818
rect 11866 24784 11900 24818
rect 11900 24784 11934 24818
rect 11934 24784 11968 24818
rect 11968 24784 12002 24818
rect 12002 24784 12036 24818
rect 12036 24784 12070 24818
rect 12070 24784 12104 24818
rect 12104 24784 12138 24818
rect 12138 24784 12172 24818
rect 12172 24784 12206 24818
rect 12206 24784 12240 24818
rect 12240 24784 12274 24818
rect 12274 24784 12308 24818
rect 12308 24784 12342 24818
rect 12342 24784 12376 24818
rect 12376 24784 12410 24818
rect 12410 24784 12444 24818
rect 12444 24784 12478 24818
rect 12478 24784 12512 24818
rect 12512 24784 12546 24818
rect 12546 24784 12580 24818
rect 12580 24784 12614 24818
rect 12614 24784 12648 24818
rect 12648 24784 12682 24818
rect 12682 24784 12716 24818
rect 12716 24784 12750 24818
rect 12750 24784 12784 24818
rect 12784 24784 12818 24818
rect 12818 24784 12852 24818
rect 12852 24784 12886 24818
rect 12886 24784 12920 24818
rect 12920 24784 12954 24818
rect 12954 24784 12988 24818
rect 12988 24784 13022 24818
rect 13022 24784 13056 24818
rect 13056 24784 13090 24818
rect 13090 24784 13124 24818
rect 13124 24784 13158 24818
rect 13158 24784 13192 24818
rect 13192 24784 13226 24818
rect 13226 24784 13260 24818
rect 13260 24784 13294 24818
rect 13294 24784 13328 24818
rect 13328 24784 13362 24818
rect 13362 24784 13396 24818
rect 13396 24784 13430 24818
rect 13430 24784 13464 24818
rect 13464 24784 13498 24818
rect 13498 24784 13532 24818
rect 13532 24784 13566 24818
rect 13566 24784 13600 24818
rect 13600 24784 13634 24818
rect 13634 24784 13668 24818
rect 13668 24784 13702 24818
rect 13702 24784 13736 24818
rect 13736 24784 13770 24818
rect 13770 24784 13804 24818
rect 13804 24784 13838 24818
rect 13838 24784 13872 24818
rect 13872 24784 13906 24818
rect 13906 24784 13940 24818
rect 13940 24784 13974 24818
rect 13974 24784 14008 24818
rect 14008 24784 14042 24818
rect 14042 24784 14076 24818
rect 14076 24784 14110 24818
rect 14110 24784 14144 24818
rect 14144 24784 14178 24818
rect 14178 24784 14212 24818
rect 14212 24784 14246 24818
rect 14246 24784 14280 24818
rect 14280 24784 14314 24818
rect 14314 24784 14348 24818
rect 14348 24784 14382 24818
rect 14382 24784 14416 24818
rect 14416 24784 14450 24818
rect 14450 24784 14484 24818
rect 14484 24784 14518 24818
rect 14518 24784 14552 24818
rect 14552 24784 14586 24818
rect 14586 24784 14620 24818
rect 14620 24784 14654 24818
rect 14654 24784 14688 24818
rect 14688 24784 14722 24818
rect 14722 24784 14756 24818
rect 14756 24784 14790 24818
rect 14790 24784 14824 24818
rect 14824 24784 14858 24818
rect 14858 24784 14870 24818
rect 88 24719 122 24753
rect 161 24746 195 24753
rect 234 24746 268 24753
rect 307 24746 341 24753
rect 380 24746 414 24753
rect 453 24746 487 24753
rect 526 24746 560 24753
rect 599 24746 633 24753
rect 672 24746 706 24753
rect 745 24746 779 24753
rect 818 24746 852 24753
rect 891 24746 925 24753
rect 964 24746 998 24753
rect 1037 24746 1071 24753
rect 1110 24746 1144 24753
rect 1183 24746 1217 24753
rect 1256 24746 1290 24753
rect 1329 24746 1363 24753
rect 1402 24746 1436 24753
rect 1475 24746 1509 24753
rect 1548 24746 1582 24753
rect 1621 24746 1655 24753
rect 1694 24746 1728 24753
rect 1767 24746 1801 24753
rect 1840 24746 1874 24753
rect 1913 24746 1947 24753
rect 1986 24746 2020 24753
rect 2059 24746 2093 24753
rect 2132 24746 2166 24753
rect 2205 24746 2239 24753
rect 161 24719 193 24746
rect 193 24719 195 24746
rect 234 24719 262 24746
rect 262 24719 268 24746
rect 307 24719 331 24746
rect 331 24719 341 24746
rect 380 24719 400 24746
rect 400 24719 414 24746
rect 453 24719 469 24746
rect 469 24719 487 24746
rect 526 24719 538 24746
rect 538 24719 560 24746
rect 599 24719 607 24746
rect 607 24719 633 24746
rect 672 24719 676 24746
rect 676 24719 706 24746
rect 745 24719 779 24746
rect 818 24719 848 24746
rect 848 24719 852 24746
rect 891 24719 917 24746
rect 917 24719 925 24746
rect 964 24719 986 24746
rect 986 24719 998 24746
rect 1037 24719 1054 24746
rect 1054 24719 1071 24746
rect 1110 24719 1122 24746
rect 1122 24719 1144 24746
rect 1183 24719 1190 24746
rect 1190 24719 1217 24746
rect 1256 24719 1258 24746
rect 1258 24719 1290 24746
rect 1329 24719 1360 24746
rect 1360 24719 1363 24746
rect 1402 24719 1428 24746
rect 1428 24719 1436 24746
rect 1475 24719 1496 24746
rect 1496 24719 1509 24746
rect 1548 24719 1564 24746
rect 1564 24719 1582 24746
rect 1621 24719 1632 24746
rect 1632 24719 1655 24746
rect 1694 24719 1700 24746
rect 1700 24719 1728 24746
rect 1767 24719 1768 24746
rect 1768 24719 1801 24746
rect 1840 24719 1870 24746
rect 1870 24719 1874 24746
rect 1913 24719 1938 24746
rect 1938 24719 1947 24746
rect 1986 24719 2006 24746
rect 2006 24719 2020 24746
rect 2059 24719 2074 24746
rect 2074 24719 2093 24746
rect 2132 24719 2142 24746
rect 2142 24719 2166 24746
rect 2205 24719 2210 24746
rect 2210 24719 2239 24746
rect 2278 24719 2312 24753
rect 2351 24746 2385 24753
rect 2424 24746 2458 24753
rect 2497 24746 2531 24753
rect 2570 24746 2604 24753
rect 2643 24746 2677 24753
rect 2716 24746 2750 24753
rect 2789 24746 2823 24753
rect 2862 24746 2896 24753
rect 2935 24746 2969 24753
rect 3008 24746 3042 24753
rect 3081 24746 3115 24753
rect 3154 24746 3188 24753
rect 3227 24746 3261 24753
rect 3300 24746 3334 24753
rect 3373 24746 3407 24753
rect 3446 24746 3480 24753
rect 3519 24746 3553 24753
rect 3592 24746 3626 24753
rect 3665 24746 3699 24753
rect 3738 24746 3772 24753
rect 3811 24746 3845 24753
rect 3884 24746 3918 24753
rect 3957 24746 3991 24753
rect 4030 24746 4064 24753
rect 4103 24746 4137 24753
rect 4176 24746 4210 24753
rect 4249 24746 4283 24753
rect 4322 24746 4356 24753
rect 4395 24746 4429 24753
rect 4468 24746 14870 24784
rect 2351 24719 2380 24746
rect 2380 24719 2385 24746
rect 2424 24719 2448 24746
rect 2448 24719 2458 24746
rect 2497 24719 2516 24746
rect 2516 24719 2531 24746
rect 2570 24719 2584 24746
rect 2584 24719 2604 24746
rect 2643 24719 2652 24746
rect 2652 24719 2677 24746
rect 2716 24719 2720 24746
rect 2720 24719 2750 24746
rect 2789 24719 2822 24746
rect 2822 24719 2823 24746
rect 2862 24719 2890 24746
rect 2890 24719 2896 24746
rect 2935 24719 2958 24746
rect 2958 24719 2969 24746
rect 3008 24719 3026 24746
rect 3026 24719 3042 24746
rect 3081 24719 3094 24746
rect 3094 24719 3115 24746
rect 3154 24719 3162 24746
rect 3162 24719 3188 24746
rect 3227 24719 3230 24746
rect 3230 24719 3261 24746
rect 3300 24719 3332 24746
rect 3332 24719 3334 24746
rect 3373 24719 3400 24746
rect 3400 24719 3407 24746
rect 3446 24719 3468 24746
rect 3468 24719 3480 24746
rect 3519 24719 3536 24746
rect 3536 24719 3553 24746
rect 3592 24719 3604 24746
rect 3604 24719 3626 24746
rect 3665 24719 3672 24746
rect 3672 24719 3699 24746
rect 3738 24719 3740 24746
rect 3740 24719 3772 24746
rect 3811 24719 3842 24746
rect 3842 24719 3845 24746
rect 3884 24719 3910 24746
rect 3910 24719 3918 24746
rect 3957 24719 3978 24746
rect 3978 24719 3991 24746
rect 4030 24719 4046 24746
rect 4046 24719 4064 24746
rect 4103 24719 4114 24746
rect 4114 24719 4137 24746
rect 4176 24719 4182 24746
rect 4182 24719 4210 24746
rect 4249 24719 4250 24746
rect 4250 24719 4283 24746
rect 4322 24719 4352 24746
rect 4352 24719 4356 24746
rect 4395 24719 4420 24746
rect 4420 24719 4429 24746
rect 4468 24719 4488 24746
rect 4488 24719 4522 24746
rect 4522 24719 4556 24746
rect 4556 24719 4590 24746
rect 4590 24719 4624 24746
rect 4624 24719 4658 24746
rect 4658 24719 4692 24746
rect 4692 24719 4726 24746
rect 4726 24719 4760 24746
rect 4760 24719 4794 24746
rect 4794 24719 4828 24746
rect 4828 24719 4862 24746
rect 4862 24719 4896 24746
rect 4896 24719 4930 24746
rect 4930 24719 4964 24746
rect 4964 24719 4998 24746
rect 4998 24719 5032 24746
rect 5032 24719 5066 24746
rect 5066 24719 5100 24746
rect 5100 24719 5134 24746
rect 5134 24719 5168 24746
rect 5168 24719 5202 24746
rect 5202 24719 5236 24746
rect 5236 24719 5270 24746
rect 5270 24719 5304 24746
rect 5304 24719 5338 24746
rect 5338 24719 5372 24746
rect 5372 24719 5406 24746
rect 5406 24719 5440 24746
rect 5440 24719 5474 24746
rect 5474 24719 5508 24746
rect 5508 24719 5542 24746
rect 5542 24719 5576 24746
rect 5576 24719 5610 24746
rect 5610 24719 5644 24746
rect 5644 24719 5678 24746
rect 5678 24719 5712 24746
rect 5712 24719 5746 24746
rect 5746 24719 5780 24746
rect 5780 24719 5814 24746
rect 5814 24719 5848 24746
rect 5848 24719 5882 24746
rect 5882 24719 5916 24746
rect 5916 24719 5950 24746
rect 5950 24719 5984 24746
rect 5984 24719 6018 24746
rect 6018 24719 6052 24746
rect 6052 24719 6086 24746
rect 6086 24719 6120 24746
rect 6120 24719 6154 24746
rect 6154 24719 6188 24746
rect 6188 24719 6222 24746
rect 6222 24719 6256 24746
rect 6256 24719 6290 24746
rect 6290 24719 6324 24746
rect 6324 24719 6358 24746
rect 6358 24719 6392 24746
rect 6392 24719 6426 24746
rect 6426 24719 6460 24746
rect 6460 24719 6494 24746
rect 6494 24719 6528 24746
rect 6528 24719 6562 24746
rect 6562 24719 6596 24746
rect 6596 24719 6630 24746
rect 6630 24719 6664 24746
rect 6664 24719 6698 24746
rect 6698 24719 6732 24746
rect 6732 24719 6766 24746
rect 6766 24719 6800 24746
rect 6800 24719 6834 24746
rect 6834 24719 6868 24746
rect 6868 24719 6902 24746
rect 6902 24719 6936 24746
rect 6936 24719 6970 24746
rect 6970 24719 7004 24746
rect 7004 24719 7038 24746
rect 7038 24719 7072 24746
rect 7072 24719 7106 24746
rect 7106 24719 7140 24746
rect 7140 24719 7174 24746
rect 7174 24719 7208 24746
rect 7208 24719 7242 24746
rect 7242 24719 7276 24746
rect 7276 24719 7310 24746
rect 7310 24719 7344 24746
rect 7344 24719 7378 24746
rect 7378 24719 7412 24746
rect 7412 24719 7446 24746
rect 7446 24719 7480 24746
rect 7480 24719 7514 24746
rect 7514 24719 7548 24746
rect 7548 24719 7582 24746
rect 7582 24719 7616 24746
rect 7616 24719 7650 24746
rect 7650 24719 7684 24746
rect 7684 24719 7718 24746
rect 7718 24719 7752 24746
rect 7752 24719 7786 24746
rect 7786 24719 7820 24746
rect 7820 24719 7854 24746
rect 7854 24719 7888 24746
rect 7888 24719 7922 24746
rect 7922 24719 7956 24746
rect 7956 24719 7990 24746
rect 7990 24719 8024 24746
rect 8024 24719 8058 24746
rect 8058 24719 8092 24746
rect 8092 24719 8126 24746
rect 8126 24719 8160 24746
rect 8160 24719 8194 24746
rect 8194 24719 8228 24746
rect 8228 24719 8262 24746
rect 8262 24719 8296 24746
rect 8296 24719 8330 24746
rect 8330 24719 8364 24746
rect 8364 24719 8398 24746
rect 8398 24719 8432 24746
rect 8432 24719 8466 24746
rect 8466 24719 8500 24746
rect 8500 24719 8534 24746
rect 8534 24719 8568 24746
rect 8568 24719 8602 24746
rect 8602 24719 8636 24746
rect 8636 24719 8670 24746
rect 8670 24719 8704 24746
rect 8704 24719 8738 24746
rect 8738 24719 8772 24746
rect 8772 24719 8806 24746
rect 8806 24719 8840 24746
rect 8840 24719 8874 24746
rect 8874 24719 8908 24746
rect 8908 24719 8942 24746
rect 8942 24719 8976 24746
rect 8976 24719 9010 24746
rect 9010 24719 9044 24746
rect 9044 24719 9078 24746
rect 9078 24719 9112 24746
rect 9112 24719 9146 24746
rect 9146 24719 9180 24746
rect 9180 24719 9214 24746
rect 9214 24719 9248 24746
rect 9248 24719 9282 24746
rect 9282 24719 9316 24746
rect 9316 24719 9350 24746
rect 9350 24719 9384 24746
rect 9384 24719 9418 24746
rect 9418 24719 9452 24746
rect 9452 24719 9486 24746
rect 9486 24719 9520 24746
rect 9520 24719 9554 24746
rect 9554 24719 9588 24746
rect 9588 24719 9622 24746
rect 9622 24719 9656 24746
rect 9656 24719 9690 24746
rect 9690 24719 9724 24746
rect 9724 24719 9758 24746
rect 9758 24719 9792 24746
rect 9792 24719 9826 24746
rect 9826 24719 9860 24746
rect 9860 24719 9894 24746
rect 9894 24719 9928 24746
rect 9928 24719 9962 24746
rect 9962 24719 9996 24746
rect 9996 24719 10030 24746
rect 10030 24719 10064 24746
rect 10064 24719 10098 24746
rect 10098 24719 10132 24746
rect 10132 24719 10166 24746
rect 10166 24719 10200 24746
rect 10200 24719 10234 24746
rect 10234 24719 10268 24746
rect 10268 24719 10302 24746
rect 10302 24719 10336 24746
rect 10336 24719 10370 24746
rect 10370 24719 10404 24746
rect 10404 24719 10438 24746
rect 10438 24719 10472 24746
rect 10472 24719 10506 24746
rect 10506 24719 10540 24746
rect 10540 24719 10574 24746
rect 10574 24719 10608 24746
rect 10608 24719 10642 24746
rect 10642 24719 10676 24746
rect 10676 24719 10710 24746
rect 10710 24719 10744 24746
rect 10744 24719 10778 24746
rect 10778 24719 10812 24746
rect 10812 24719 10846 24746
rect 10846 24719 10880 24746
rect 10880 24719 10914 24746
rect 10914 24719 10948 24746
rect 10948 24719 10982 24746
rect 10982 24719 11016 24746
rect 11016 24719 11050 24746
rect 11050 24719 11084 24746
rect 11084 24719 11118 24746
rect 11118 24719 11152 24746
rect 11152 24719 11186 24746
rect 11186 24719 11220 24746
rect 11220 24719 11254 24746
rect 11254 24719 11288 24746
rect 11288 24719 11322 24746
rect 11322 24719 11356 24746
rect 11356 24719 11390 24746
rect 11390 24719 11424 24746
rect 11424 24719 11458 24746
rect 11458 24719 11492 24746
rect 11492 24719 11526 24746
rect 11526 24719 11560 24746
rect 11560 24719 11594 24746
rect 11594 24719 11628 24746
rect 11628 24719 11662 24746
rect 11662 24719 11696 24746
rect 11696 24719 11730 24746
rect 11730 24719 11764 24746
rect 11764 24719 11798 24746
rect 11798 24719 11832 24746
rect 11832 24719 11866 24746
rect 11866 24719 11900 24746
rect 11900 24719 11934 24746
rect 11934 24719 11968 24746
rect 11968 24719 12002 24746
rect 12002 24719 12036 24746
rect 12036 24719 12070 24746
rect 12070 24719 12104 24746
rect 12104 24719 12138 24746
rect 12138 24719 12172 24746
rect 12172 24719 12206 24746
rect 12206 24719 12240 24746
rect 12240 24719 12274 24746
rect 12274 24719 12308 24746
rect 12308 24719 12342 24746
rect 12342 24719 12376 24746
rect 12376 24719 12410 24746
rect 12410 24719 12444 24746
rect 12444 24719 12478 24746
rect 12478 24719 12512 24746
rect 12512 24719 12546 24746
rect 12546 24719 12580 24746
rect 12580 24719 12614 24746
rect 12614 24719 12648 24746
rect 12648 24719 12682 24746
rect 12682 24719 12716 24746
rect 12716 24719 12750 24746
rect 12750 24719 12784 24746
rect 12784 24719 12818 24746
rect 12818 24719 12852 24746
rect 12852 24719 12886 24746
rect 12886 24719 12920 24746
rect 12920 24719 12954 24746
rect 12954 24719 12988 24746
rect 12988 24719 13022 24746
rect 13022 24719 13056 24746
rect 13056 24719 13090 24746
rect 13090 24719 13124 24746
rect 13124 24719 13158 24746
rect 13158 24719 13192 24746
rect 13192 24719 13226 24746
rect 13226 24719 13260 24746
rect 13260 24719 13294 24746
rect 13294 24719 13328 24746
rect 13328 24719 13362 24746
rect 13362 24719 13396 24746
rect 13396 24719 13430 24746
rect 13430 24719 13464 24746
rect 13464 24719 13498 24746
rect 13498 24719 13532 24746
rect 13532 24719 13566 24746
rect 13566 24719 13600 24746
rect 13600 24719 13634 24746
rect 13634 24719 13668 24746
rect 13668 24719 13702 24746
rect 13702 24719 13736 24746
rect 13736 24719 13770 24746
rect 13770 24719 13804 24746
rect 13804 24719 13838 24746
rect 13838 24719 13872 24746
rect 13872 24719 13906 24746
rect 13906 24719 13940 24746
rect 13940 24719 13974 24746
rect 13974 24719 14008 24746
rect 14008 24719 14042 24746
rect 14042 24719 14076 24746
rect 14076 24719 14110 24746
rect 14110 24719 14144 24746
rect 14144 24719 14178 24746
rect 14178 24719 14212 24746
rect 14212 24719 14246 24746
rect 14246 24719 14280 24746
rect 14280 24719 14314 24746
rect 14314 24719 14348 24746
rect 14348 24719 14382 24746
rect 14382 24719 14416 24746
rect 14416 24719 14450 24746
rect 14450 24719 14484 24746
rect 14484 24719 14518 24746
rect 14518 24719 14552 24746
rect 14552 24719 14586 24746
rect 14586 24719 14620 24746
rect 14620 24719 14654 24746
rect 14654 24719 14688 24746
rect 14688 24719 14722 24746
rect 14722 24719 14756 24746
rect 14756 24719 14790 24746
rect 14790 24719 14824 24746
rect 14824 24719 14858 24746
rect 14858 24719 14870 24746
rect 70 19825 77 19858
rect 77 19825 104 19858
rect 143 19825 146 19858
rect 146 19825 177 19858
rect 216 19825 249 19858
rect 249 19825 250 19858
rect 289 19825 318 19858
rect 318 19825 323 19858
rect 362 19825 387 19858
rect 387 19825 396 19858
rect 435 19825 456 19858
rect 456 19825 469 19858
rect 508 19825 525 19858
rect 525 19825 542 19858
rect 581 19825 594 19858
rect 594 19825 615 19858
rect 654 19825 663 19858
rect 663 19825 688 19858
rect 727 19825 732 19858
rect 732 19825 761 19858
rect 800 19825 801 19858
rect 801 19825 834 19858
rect 873 19825 905 19858
rect 905 19825 907 19858
rect 946 19825 974 19858
rect 974 19825 980 19858
rect 1019 19825 1043 19858
rect 1043 19825 1053 19858
rect 1092 19825 1112 19858
rect 1112 19825 1126 19858
rect 1165 19825 1181 19858
rect 1181 19825 1199 19858
rect 1238 19825 1250 19858
rect 1250 19825 1272 19858
rect 1311 19825 1319 19858
rect 1319 19825 1345 19858
rect 1384 19825 1388 19858
rect 1388 19825 1418 19858
rect 1457 19825 1491 19858
rect 1530 19825 1560 19858
rect 1560 19825 1564 19858
rect 1603 19825 1629 19858
rect 1629 19825 1637 19858
rect 1676 19825 1698 19858
rect 1698 19825 1710 19858
rect 1749 19825 1767 19858
rect 1767 19825 1783 19858
rect 1822 19825 1836 19858
rect 1836 19825 1856 19858
rect 1895 19825 1905 19858
rect 1905 19825 1929 19858
rect 1968 19825 1974 19858
rect 1974 19825 2002 19858
rect 2041 19825 2043 19858
rect 2043 19825 2075 19858
rect 2114 19825 2147 19858
rect 2147 19825 2148 19858
rect 2187 19825 2216 19858
rect 2216 19825 2221 19858
rect 2260 19825 2285 19858
rect 2285 19825 2294 19858
rect 2333 19825 2354 19858
rect 2354 19825 2367 19858
rect 2406 19825 2423 19858
rect 2423 19825 2440 19858
rect 2479 19825 2492 19858
rect 2492 19825 2513 19858
rect 2552 19825 2561 19858
rect 2561 19825 2586 19858
rect 2625 19825 2630 19858
rect 2630 19825 2659 19858
rect 2698 19825 2699 19858
rect 2699 19825 2732 19858
rect 2771 19825 2802 19858
rect 2802 19825 2805 19858
rect 2844 19825 2871 19858
rect 2871 19825 2878 19858
rect 2917 19825 2940 19858
rect 2940 19825 2951 19858
rect 2990 19825 3009 19858
rect 3009 19825 3024 19858
rect 3063 19825 3078 19858
rect 3078 19825 3097 19858
rect 3136 19825 3147 19858
rect 3147 19825 3170 19858
rect 70 19824 104 19825
rect 143 19824 177 19825
rect 216 19824 250 19825
rect 289 19824 323 19825
rect 362 19824 396 19825
rect 435 19824 469 19825
rect 508 19824 542 19825
rect 581 19824 615 19825
rect 654 19824 688 19825
rect 727 19824 761 19825
rect 800 19824 834 19825
rect 873 19824 907 19825
rect 946 19824 980 19825
rect 1019 19824 1053 19825
rect 1092 19824 1126 19825
rect 1165 19824 1199 19825
rect 1238 19824 1272 19825
rect 1311 19824 1345 19825
rect 1384 19824 1418 19825
rect 1457 19824 1491 19825
rect 1530 19824 1564 19825
rect 1603 19824 1637 19825
rect 1676 19824 1710 19825
rect 1749 19824 1783 19825
rect 1822 19824 1856 19825
rect 1895 19824 1929 19825
rect 1968 19824 2002 19825
rect 2041 19824 2075 19825
rect 2114 19824 2148 19825
rect 2187 19824 2221 19825
rect 2260 19824 2294 19825
rect 2333 19824 2367 19825
rect 2406 19824 2440 19825
rect 2479 19824 2513 19825
rect 2552 19824 2586 19825
rect 2625 19824 2659 19825
rect 2698 19824 2732 19825
rect 2771 19824 2805 19825
rect 2844 19824 2878 19825
rect 2917 19824 2951 19825
rect 2990 19824 3024 19825
rect 3063 19824 3097 19825
rect 3136 19824 3170 19825
rect 3209 19824 3243 19858
rect 3282 19824 3316 19858
rect 3354 19824 3388 19858
rect 3426 19824 3460 19858
rect 3498 19824 3532 19858
rect 3570 19824 3604 19858
rect 3642 19824 3676 19858
rect 3714 19824 3748 19858
rect 3786 19824 3820 19858
rect 3858 19824 3892 19858
rect 3930 19824 3964 19858
rect 4002 19824 4036 19858
rect 4074 19824 4108 19858
rect 4146 19824 4180 19858
rect 4218 19824 4252 19858
rect 4290 19824 4324 19858
rect 4362 19824 4396 19858
rect 4434 19824 4468 19858
rect 4506 19824 4540 19858
rect 4578 19824 4612 19858
rect 4650 19824 4684 19858
rect 4722 19824 4756 19858
rect 4794 19824 4828 19858
rect 4866 19824 4900 19858
rect 4938 19824 4972 19858
rect 5010 19824 5044 19858
rect 5082 19824 5116 19858
rect 5154 19824 5188 19858
rect 5226 19824 5260 19858
rect 5298 19824 5332 19858
rect 5370 19824 5404 19858
rect 5442 19824 5476 19858
rect 5514 19824 5548 19858
rect 5586 19824 5620 19858
rect 5658 19824 5692 19858
rect 5730 19824 5764 19858
rect 5802 19824 5836 19858
rect 5874 19824 5908 19858
rect 5946 19824 5980 19858
rect 6018 19824 6052 19858
rect 6090 19824 6124 19858
rect 6162 19824 6196 19858
rect 6234 19824 6268 19858
rect 6306 19824 6340 19858
rect 6378 19824 6412 19858
rect 6450 19824 6484 19858
rect 6522 19824 6556 19858
rect 6594 19824 6628 19858
rect 6666 19824 6700 19858
rect 6738 19824 6772 19858
rect 6810 19824 6844 19858
rect 6882 19824 6916 19858
rect 6954 19824 6988 19858
rect 7026 19824 7060 19858
rect 7098 19824 7132 19858
rect 7170 19824 7204 19858
rect 7242 19824 7276 19858
rect 7314 19824 7348 19858
rect 7386 19824 7420 19858
rect 7458 19824 7492 19858
rect 7530 19824 7564 19858
rect 7602 19824 7636 19858
rect 7674 19824 7708 19858
rect 7746 19824 7780 19858
rect 7818 19824 7852 19858
rect 7890 19824 7924 19858
rect 7962 19824 7996 19858
rect 8034 19824 8068 19858
rect 8106 19824 8140 19858
rect 8178 19824 8212 19858
rect 8250 19824 8284 19858
rect 8322 19824 8356 19858
rect 8394 19824 8428 19858
rect 8466 19824 8500 19858
rect 8538 19824 8572 19858
rect 8610 19824 8644 19858
rect 8682 19824 8716 19858
rect 8754 19824 8788 19858
rect 8826 19824 8860 19858
rect 8898 19824 8932 19858
rect 8970 19824 9004 19858
rect 9042 19824 9076 19858
rect 9114 19824 9148 19858
rect 9186 19824 9220 19858
rect 9258 19824 9292 19858
rect 9330 19824 9364 19858
rect 9402 19824 9436 19858
rect 9474 19824 9508 19858
rect 9546 19824 9580 19858
rect 9618 19824 9652 19858
rect 9690 19824 9724 19858
rect 9762 19824 9796 19858
rect 9834 19824 9868 19858
rect 9906 19824 9940 19858
rect 9978 19824 10012 19858
rect 10050 19824 10084 19858
rect 10122 19824 10156 19858
rect 10194 19824 10228 19858
rect 10266 19824 10300 19858
rect 10338 19824 10372 19858
rect 10410 19824 10444 19858
rect 10482 19824 10516 19858
rect 10554 19824 10588 19858
rect 10626 19824 10660 19858
rect 10698 19824 10732 19858
rect 10770 19824 10804 19858
rect 10842 19824 10876 19858
rect 10914 19824 10948 19858
rect 10986 19824 11020 19858
rect 11058 19824 11092 19858
rect 11130 19824 11164 19858
rect 11202 19824 11236 19858
rect 11274 19824 11308 19858
rect 11346 19824 11380 19858
rect 11418 19824 11452 19858
rect 11490 19824 11524 19858
rect 11562 19824 11596 19858
rect 11634 19824 11668 19858
rect 11706 19824 11740 19858
rect 11778 19824 11812 19858
rect 11850 19824 11884 19858
rect 11922 19824 11956 19858
rect 11994 19824 12028 19858
rect 12066 19824 12100 19858
rect 12138 19824 12172 19858
rect 12210 19824 12244 19858
rect 12282 19824 12316 19858
rect 12354 19824 12388 19858
rect 12426 19824 12460 19858
rect 12498 19824 12532 19858
rect 12570 19824 12604 19858
rect 12642 19824 12676 19858
rect 12714 19824 12748 19858
rect 12786 19824 12820 19858
rect 12858 19824 12892 19858
rect 12930 19824 12964 19858
rect 13002 19824 13036 19858
rect 13074 19824 13108 19858
rect 13146 19824 13180 19858
rect 13218 19824 13252 19858
rect 13290 19824 13324 19858
rect 13362 19824 13396 19858
rect 13434 19824 13468 19858
rect 13506 19824 13540 19858
rect 13578 19824 13612 19858
rect 13650 19824 13684 19858
rect 13722 19824 13756 19858
rect 13794 19824 13828 19858
rect 13866 19824 13900 19858
rect 13938 19824 13972 19858
rect 14010 19824 14044 19858
rect 14082 19824 14116 19858
rect 14154 19824 14188 19858
rect 14226 19824 14260 19858
rect 14298 19824 14332 19858
rect 14370 19824 14404 19858
rect 14442 19824 14476 19858
rect 14514 19831 14548 19858
rect 14586 19831 14620 19858
rect 14658 19831 14692 19858
rect 14514 19824 14518 19831
rect 14518 19824 14548 19831
rect 14586 19824 14601 19831
rect 14601 19824 14620 19831
rect 14658 19824 14684 19831
rect 14684 19824 14692 19831
rect 14730 19831 14764 19858
rect 14802 19831 14836 19858
rect 14730 19824 14733 19831
rect 14733 19824 14764 19831
rect 14802 19824 14816 19831
rect 14816 19824 14836 19831
rect 14874 19824 14908 19858
rect 70 19757 77 19772
rect 77 19757 104 19772
rect 143 19757 146 19772
rect 146 19757 177 19772
rect 216 19757 249 19772
rect 249 19757 250 19772
rect 289 19757 318 19772
rect 318 19757 323 19772
rect 362 19757 387 19772
rect 387 19757 396 19772
rect 435 19757 456 19772
rect 456 19757 469 19772
rect 508 19757 525 19772
rect 525 19757 542 19772
rect 581 19757 594 19772
rect 594 19757 615 19772
rect 654 19757 663 19772
rect 663 19757 688 19772
rect 727 19757 732 19772
rect 732 19757 761 19772
rect 800 19757 801 19772
rect 801 19757 834 19772
rect 873 19757 905 19772
rect 905 19757 907 19772
rect 946 19757 974 19772
rect 974 19757 980 19772
rect 1019 19757 1043 19772
rect 1043 19757 1053 19772
rect 1092 19757 1112 19772
rect 1112 19757 1126 19772
rect 1165 19757 1181 19772
rect 1181 19757 1199 19772
rect 1238 19757 1250 19772
rect 1250 19757 1272 19772
rect 1311 19757 1319 19772
rect 1319 19757 1345 19772
rect 1384 19757 1388 19772
rect 1388 19757 1418 19772
rect 1457 19757 1491 19772
rect 1530 19757 1560 19772
rect 1560 19757 1564 19772
rect 1603 19757 1629 19772
rect 1629 19757 1637 19772
rect 1676 19757 1698 19772
rect 1698 19757 1710 19772
rect 1749 19757 1767 19772
rect 1767 19757 1783 19772
rect 1822 19757 1836 19772
rect 1836 19757 1856 19772
rect 1895 19757 1905 19772
rect 1905 19757 1929 19772
rect 1968 19757 1974 19772
rect 1974 19757 2002 19772
rect 2041 19757 2043 19772
rect 2043 19757 2075 19772
rect 2114 19757 2147 19772
rect 2147 19757 2148 19772
rect 2187 19757 2216 19772
rect 2216 19757 2221 19772
rect 2260 19757 2285 19772
rect 2285 19757 2294 19772
rect 2333 19757 2354 19772
rect 2354 19757 2367 19772
rect 2406 19757 2423 19772
rect 2423 19757 2440 19772
rect 2479 19757 2492 19772
rect 2492 19757 2513 19772
rect 2552 19757 2561 19772
rect 2561 19757 2586 19772
rect 2625 19757 2630 19772
rect 2630 19757 2659 19772
rect 2698 19757 2699 19772
rect 2699 19757 2732 19772
rect 2771 19757 2802 19772
rect 2802 19757 2805 19772
rect 2844 19757 2871 19772
rect 2871 19757 2878 19772
rect 2917 19757 2940 19772
rect 2940 19757 2951 19772
rect 2990 19757 3009 19772
rect 3009 19757 3024 19772
rect 3063 19757 3078 19772
rect 3078 19757 3097 19772
rect 3136 19757 3147 19772
rect 3147 19757 3170 19772
rect 70 19738 104 19757
rect 143 19738 177 19757
rect 216 19738 250 19757
rect 289 19738 323 19757
rect 362 19738 396 19757
rect 435 19738 469 19757
rect 508 19738 542 19757
rect 581 19738 615 19757
rect 654 19738 688 19757
rect 727 19738 761 19757
rect 800 19738 834 19757
rect 873 19738 907 19757
rect 946 19738 980 19757
rect 1019 19738 1053 19757
rect 1092 19738 1126 19757
rect 1165 19738 1199 19757
rect 1238 19738 1272 19757
rect 1311 19738 1345 19757
rect 1384 19738 1418 19757
rect 1457 19738 1491 19757
rect 1530 19738 1564 19757
rect 1603 19738 1637 19757
rect 1676 19738 1710 19757
rect 1749 19738 1783 19757
rect 1822 19738 1856 19757
rect 1895 19738 1929 19757
rect 1968 19738 2002 19757
rect 2041 19738 2075 19757
rect 2114 19738 2148 19757
rect 2187 19738 2221 19757
rect 2260 19738 2294 19757
rect 2333 19738 2367 19757
rect 2406 19738 2440 19757
rect 2479 19738 2513 19757
rect 2552 19738 2586 19757
rect 2625 19738 2659 19757
rect 2698 19738 2732 19757
rect 2771 19738 2805 19757
rect 2844 19738 2878 19757
rect 2917 19738 2951 19757
rect 2990 19738 3024 19757
rect 3063 19738 3097 19757
rect 3136 19738 3170 19757
rect 3209 19738 3243 19772
rect 3282 19738 3316 19772
rect 3354 19738 3388 19772
rect 3426 19738 3460 19772
rect 3498 19738 3532 19772
rect 3570 19738 3604 19772
rect 3642 19738 3676 19772
rect 3714 19738 3748 19772
rect 3786 19738 3820 19772
rect 3858 19738 3892 19772
rect 3930 19738 3964 19772
rect 4002 19738 4036 19772
rect 4074 19738 4108 19772
rect 4146 19738 4180 19772
rect 4218 19738 4252 19772
rect 4290 19738 4324 19772
rect 4362 19738 4396 19772
rect 4434 19738 4468 19772
rect 4506 19738 4540 19772
rect 4578 19738 4612 19772
rect 4650 19738 4684 19772
rect 4722 19738 4756 19772
rect 4794 19738 4828 19772
rect 4866 19738 4900 19772
rect 4938 19738 4972 19772
rect 5010 19738 5044 19772
rect 5082 19738 5116 19772
rect 5154 19738 5188 19772
rect 5226 19738 5260 19772
rect 5298 19738 5332 19772
rect 5370 19738 5404 19772
rect 5442 19738 5476 19772
rect 5514 19738 5548 19772
rect 5586 19738 5620 19772
rect 5658 19738 5692 19772
rect 5730 19738 5764 19772
rect 5802 19738 5836 19772
rect 5874 19738 5908 19772
rect 5946 19738 5980 19772
rect 6018 19738 6052 19772
rect 6090 19738 6124 19772
rect 6162 19738 6196 19772
rect 6234 19738 6268 19772
rect 6306 19738 6340 19772
rect 6378 19738 6412 19772
rect 6450 19738 6484 19772
rect 6522 19738 6556 19772
rect 6594 19738 6628 19772
rect 6666 19738 6700 19772
rect 6738 19738 6772 19772
rect 6810 19738 6844 19772
rect 6882 19738 6916 19772
rect 6954 19738 6988 19772
rect 7026 19738 7060 19772
rect 7098 19738 7132 19772
rect 7170 19738 7204 19772
rect 7242 19738 7276 19772
rect 7314 19738 7348 19772
rect 7386 19738 7420 19772
rect 7458 19738 7492 19772
rect 7530 19738 7564 19772
rect 7602 19738 7636 19772
rect 7674 19738 7708 19772
rect 7746 19738 7780 19772
rect 7818 19738 7852 19772
rect 7890 19738 7924 19772
rect 7962 19738 7996 19772
rect 8034 19738 8068 19772
rect 8106 19738 8140 19772
rect 8178 19738 8212 19772
rect 8250 19738 8284 19772
rect 8322 19738 8356 19772
rect 8394 19738 8428 19772
rect 8466 19738 8500 19772
rect 8538 19738 8572 19772
rect 8610 19738 8644 19772
rect 8682 19738 8716 19772
rect 8754 19738 8788 19772
rect 8826 19738 8860 19772
rect 8898 19738 8932 19772
rect 8970 19738 9004 19772
rect 9042 19738 9076 19772
rect 9114 19738 9148 19772
rect 9186 19738 9220 19772
rect 9258 19738 9292 19772
rect 9330 19738 9364 19772
rect 9402 19738 9436 19772
rect 9474 19738 9508 19772
rect 9546 19738 9580 19772
rect 9618 19738 9652 19772
rect 9690 19738 9724 19772
rect 9762 19738 9796 19772
rect 9834 19738 9868 19772
rect 9906 19738 9940 19772
rect 9978 19738 10012 19772
rect 10050 19738 10084 19772
rect 10122 19738 10156 19772
rect 10194 19738 10228 19772
rect 10266 19738 10300 19772
rect 10338 19738 10372 19772
rect 10410 19738 10444 19772
rect 10482 19738 10516 19772
rect 10554 19738 10588 19772
rect 10626 19738 10660 19772
rect 10698 19738 10732 19772
rect 10770 19738 10804 19772
rect 10842 19738 10876 19772
rect 10914 19738 10948 19772
rect 10986 19738 11020 19772
rect 11058 19738 11092 19772
rect 11130 19738 11164 19772
rect 11202 19738 11236 19772
rect 11274 19738 11308 19772
rect 11346 19738 11380 19772
rect 11418 19738 11452 19772
rect 11490 19738 11524 19772
rect 11562 19738 11596 19772
rect 11634 19738 11668 19772
rect 11706 19738 11740 19772
rect 11778 19738 11812 19772
rect 11850 19738 11884 19772
rect 11922 19738 11956 19772
rect 11994 19738 12028 19772
rect 12066 19738 12100 19772
rect 12138 19738 12172 19772
rect 12210 19738 12244 19772
rect 12282 19738 12316 19772
rect 12354 19738 12388 19772
rect 12426 19738 12460 19772
rect 12498 19738 12532 19772
rect 12570 19738 12604 19772
rect 12642 19738 12676 19772
rect 12714 19738 12748 19772
rect 12786 19738 12820 19772
rect 12858 19738 12892 19772
rect 12930 19738 12964 19772
rect 13002 19738 13036 19772
rect 13074 19738 13108 19772
rect 13146 19738 13180 19772
rect 13218 19738 13252 19772
rect 13290 19738 13324 19772
rect 13362 19738 13396 19772
rect 13434 19738 13468 19772
rect 13506 19738 13540 19772
rect 13578 19738 13612 19772
rect 13650 19738 13684 19772
rect 13722 19738 13756 19772
rect 13794 19738 13828 19772
rect 13866 19738 13900 19772
rect 13938 19738 13972 19772
rect 14010 19738 14044 19772
rect 14082 19738 14116 19772
rect 14154 19738 14188 19772
rect 14226 19738 14260 19772
rect 14298 19738 14332 19772
rect 14370 19738 14404 19772
rect 14442 19738 14476 19772
rect 14514 19761 14548 19772
rect 14586 19761 14620 19772
rect 14658 19761 14692 19772
rect 14514 19738 14518 19761
rect 14518 19738 14548 19761
rect 14586 19738 14601 19761
rect 14601 19738 14620 19761
rect 14658 19738 14684 19761
rect 14684 19738 14692 19761
rect 14730 19761 14764 19772
rect 14802 19761 14836 19772
rect 14730 19738 14733 19761
rect 14733 19738 14764 19761
rect 14802 19738 14816 19761
rect 14816 19738 14836 19761
rect 14874 19738 14908 19772
rect 70 19655 104 19686
rect 143 19655 177 19686
rect 216 19655 250 19686
rect 289 19655 323 19686
rect 362 19655 396 19686
rect 435 19655 469 19686
rect 508 19655 542 19686
rect 581 19655 615 19686
rect 654 19655 688 19686
rect 727 19655 761 19686
rect 800 19655 834 19686
rect 873 19655 907 19686
rect 946 19655 980 19686
rect 1019 19655 1053 19686
rect 1092 19655 1126 19686
rect 1165 19655 1199 19686
rect 1238 19655 1272 19686
rect 1311 19655 1345 19686
rect 1384 19655 1418 19686
rect 1457 19655 1491 19686
rect 1530 19655 1564 19686
rect 1603 19655 1637 19686
rect 1676 19655 1710 19686
rect 1749 19655 1783 19686
rect 1822 19655 1856 19686
rect 1895 19655 1929 19686
rect 1968 19655 2002 19686
rect 2041 19655 2075 19686
rect 2114 19655 2148 19686
rect 2187 19655 2221 19686
rect 2260 19655 2294 19686
rect 2333 19655 2367 19686
rect 2406 19655 2440 19686
rect 2479 19655 2513 19686
rect 2552 19655 2586 19686
rect 2625 19655 2659 19686
rect 2698 19655 2732 19686
rect 2771 19655 2805 19686
rect 2844 19655 2878 19686
rect 2917 19655 2951 19686
rect 2990 19655 3024 19686
rect 3063 19655 3097 19686
rect 3136 19655 3170 19686
rect 70 19652 77 19655
rect 77 19652 104 19655
rect 143 19652 146 19655
rect 146 19652 177 19655
rect 216 19652 249 19655
rect 249 19652 250 19655
rect 289 19652 318 19655
rect 318 19652 323 19655
rect 362 19652 387 19655
rect 387 19652 396 19655
rect 435 19652 456 19655
rect 456 19652 469 19655
rect 508 19652 525 19655
rect 525 19652 542 19655
rect 581 19652 594 19655
rect 594 19652 615 19655
rect 654 19652 663 19655
rect 663 19652 688 19655
rect 727 19652 732 19655
rect 732 19652 761 19655
rect 800 19652 801 19655
rect 801 19652 834 19655
rect 873 19652 905 19655
rect 905 19652 907 19655
rect 946 19652 974 19655
rect 974 19652 980 19655
rect 1019 19652 1043 19655
rect 1043 19652 1053 19655
rect 1092 19652 1112 19655
rect 1112 19652 1126 19655
rect 1165 19652 1181 19655
rect 1181 19652 1199 19655
rect 1238 19652 1250 19655
rect 1250 19652 1272 19655
rect 1311 19652 1319 19655
rect 1319 19652 1345 19655
rect 1384 19652 1388 19655
rect 1388 19652 1418 19655
rect 1457 19652 1491 19655
rect 1530 19652 1560 19655
rect 1560 19652 1564 19655
rect 1603 19652 1629 19655
rect 1629 19652 1637 19655
rect 1676 19652 1698 19655
rect 1698 19652 1710 19655
rect 1749 19652 1767 19655
rect 1767 19652 1783 19655
rect 1822 19652 1836 19655
rect 1836 19652 1856 19655
rect 1895 19652 1905 19655
rect 1905 19652 1929 19655
rect 1968 19652 1974 19655
rect 1974 19652 2002 19655
rect 2041 19652 2043 19655
rect 2043 19652 2075 19655
rect 2114 19652 2147 19655
rect 2147 19652 2148 19655
rect 2187 19652 2216 19655
rect 2216 19652 2221 19655
rect 2260 19652 2285 19655
rect 2285 19652 2294 19655
rect 2333 19652 2354 19655
rect 2354 19652 2367 19655
rect 2406 19652 2423 19655
rect 2423 19652 2440 19655
rect 2479 19652 2492 19655
rect 2492 19652 2513 19655
rect 2552 19652 2561 19655
rect 2561 19652 2586 19655
rect 2625 19652 2630 19655
rect 2630 19652 2659 19655
rect 2698 19652 2699 19655
rect 2699 19652 2732 19655
rect 2771 19652 2802 19655
rect 2802 19652 2805 19655
rect 2844 19652 2871 19655
rect 2871 19652 2878 19655
rect 2917 19652 2940 19655
rect 2940 19652 2951 19655
rect 2990 19652 3009 19655
rect 3009 19652 3024 19655
rect 3063 19652 3078 19655
rect 3078 19652 3097 19655
rect 3136 19652 3147 19655
rect 3147 19652 3170 19655
rect 3209 19652 3243 19686
rect 3282 19652 3316 19686
rect 3354 19652 3388 19686
rect 3426 19652 3460 19686
rect 3498 19652 3532 19686
rect 3570 19652 3604 19686
rect 3642 19652 3676 19686
rect 3714 19652 3748 19686
rect 3786 19652 3820 19686
rect 3858 19652 3892 19686
rect 3930 19652 3964 19686
rect 4002 19652 4036 19686
rect 4074 19652 4108 19686
rect 4146 19652 4180 19686
rect 4218 19652 4252 19686
rect 4290 19652 4324 19686
rect 4362 19652 4396 19686
rect 4434 19652 4468 19686
rect 4506 19652 4540 19686
rect 4578 19652 4612 19686
rect 4650 19652 4684 19686
rect 4722 19652 4756 19686
rect 4794 19652 4828 19686
rect 4866 19652 4900 19686
rect 4938 19652 4972 19686
rect 5010 19652 5044 19686
rect 5082 19652 5116 19686
rect 5154 19652 5188 19686
rect 5226 19652 5260 19686
rect 5298 19652 5332 19686
rect 5370 19652 5404 19686
rect 5442 19652 5476 19686
rect 5514 19652 5548 19686
rect 5586 19652 5620 19686
rect 5658 19652 5692 19686
rect 5730 19652 5764 19686
rect 5802 19652 5836 19686
rect 5874 19652 5908 19686
rect 5946 19652 5980 19686
rect 6018 19652 6052 19686
rect 6090 19652 6124 19686
rect 6162 19652 6196 19686
rect 6234 19652 6268 19686
rect 6306 19652 6340 19686
rect 6378 19652 6412 19686
rect 6450 19652 6484 19686
rect 6522 19652 6556 19686
rect 6594 19652 6628 19686
rect 6666 19652 6700 19686
rect 6738 19652 6772 19686
rect 6810 19652 6844 19686
rect 6882 19652 6916 19686
rect 6954 19652 6988 19686
rect 7026 19652 7060 19686
rect 7098 19652 7132 19686
rect 7170 19652 7204 19686
rect 7242 19652 7276 19686
rect 7314 19652 7348 19686
rect 7386 19652 7420 19686
rect 7458 19652 7492 19686
rect 7530 19652 7564 19686
rect 7602 19652 7636 19686
rect 7674 19652 7708 19686
rect 7746 19652 7780 19686
rect 7818 19652 7852 19686
rect 7890 19652 7924 19686
rect 7962 19652 7996 19686
rect 8034 19652 8068 19686
rect 8106 19652 8140 19686
rect 8178 19652 8212 19686
rect 8250 19652 8284 19686
rect 8322 19652 8356 19686
rect 8394 19652 8428 19686
rect 8466 19652 8500 19686
rect 8538 19652 8572 19686
rect 8610 19652 8644 19686
rect 8682 19652 8716 19686
rect 8754 19652 8788 19686
rect 8826 19652 8860 19686
rect 8898 19652 8932 19686
rect 8970 19652 9004 19686
rect 9042 19652 9076 19686
rect 9114 19652 9148 19686
rect 9186 19652 9220 19686
rect 9258 19652 9292 19686
rect 9330 19652 9364 19686
rect 9402 19652 9436 19686
rect 9474 19652 9508 19686
rect 9546 19652 9580 19686
rect 9618 19652 9652 19686
rect 9690 19652 9724 19686
rect 9762 19652 9796 19686
rect 9834 19652 9868 19686
rect 9906 19652 9940 19686
rect 9978 19652 10012 19686
rect 10050 19652 10084 19686
rect 10122 19652 10156 19686
rect 10194 19652 10228 19686
rect 10266 19652 10300 19686
rect 10338 19652 10372 19686
rect 10410 19652 10444 19686
rect 10482 19652 10516 19686
rect 10554 19652 10588 19686
rect 10626 19652 10660 19686
rect 10698 19652 10732 19686
rect 10770 19652 10804 19686
rect 10842 19652 10876 19686
rect 10914 19652 10948 19686
rect 10986 19652 11020 19686
rect 11058 19652 11092 19686
rect 11130 19652 11164 19686
rect 11202 19652 11236 19686
rect 11274 19652 11308 19686
rect 11346 19652 11380 19686
rect 11418 19652 11452 19686
rect 11490 19652 11524 19686
rect 11562 19652 11596 19686
rect 11634 19652 11668 19686
rect 11706 19652 11740 19686
rect 11778 19652 11812 19686
rect 11850 19652 11884 19686
rect 11922 19652 11956 19686
rect 11994 19652 12028 19686
rect 12066 19652 12100 19686
rect 12138 19652 12172 19686
rect 12210 19652 12244 19686
rect 12282 19652 12316 19686
rect 12354 19652 12388 19686
rect 12426 19652 12460 19686
rect 12498 19652 12532 19686
rect 12570 19652 12604 19686
rect 12642 19652 12676 19686
rect 12714 19652 12748 19686
rect 12786 19652 12820 19686
rect 12858 19652 12892 19686
rect 12930 19652 12964 19686
rect 13002 19652 13036 19686
rect 13074 19652 13108 19686
rect 13146 19652 13180 19686
rect 13218 19652 13252 19686
rect 13290 19652 13324 19686
rect 13362 19652 13396 19686
rect 13434 19652 13468 19686
rect 13506 19652 13540 19686
rect 13578 19652 13612 19686
rect 13650 19652 13684 19686
rect 13722 19652 13756 19686
rect 13794 19652 13828 19686
rect 13866 19652 13900 19686
rect 13938 19652 13972 19686
rect 14010 19652 14044 19686
rect 14082 19652 14116 19686
rect 14154 19652 14188 19686
rect 14226 19652 14260 19686
rect 14298 19652 14332 19686
rect 14370 19652 14404 19686
rect 14442 19652 14476 19686
rect 14514 19657 14518 19686
rect 14518 19657 14548 19686
rect 14586 19657 14601 19686
rect 14601 19657 14620 19686
rect 14658 19657 14684 19686
rect 14684 19657 14692 19686
rect 14514 19652 14548 19657
rect 14586 19652 14620 19657
rect 14658 19652 14692 19657
rect 14730 19657 14733 19686
rect 14733 19657 14764 19686
rect 14802 19657 14816 19686
rect 14816 19657 14836 19686
rect 14730 19652 14764 19657
rect 14802 19652 14836 19657
rect 14874 19652 14908 19686
rect 70 19585 104 19600
rect 143 19585 177 19600
rect 216 19585 250 19600
rect 289 19585 323 19600
rect 362 19585 396 19600
rect 435 19585 469 19600
rect 508 19585 542 19600
rect 581 19585 615 19600
rect 654 19585 688 19600
rect 727 19585 761 19600
rect 800 19585 834 19600
rect 873 19585 907 19600
rect 946 19585 980 19600
rect 1019 19585 1053 19600
rect 1092 19585 1126 19600
rect 1165 19585 1199 19600
rect 1238 19585 1272 19600
rect 1311 19585 1345 19600
rect 1384 19585 1418 19600
rect 1457 19585 1491 19600
rect 1530 19585 1564 19600
rect 1603 19585 1637 19600
rect 1676 19585 1710 19600
rect 1749 19585 1783 19600
rect 1822 19585 1856 19600
rect 1895 19585 1929 19600
rect 1968 19585 2002 19600
rect 2041 19585 2075 19600
rect 2114 19585 2148 19600
rect 2187 19585 2221 19600
rect 2260 19585 2294 19600
rect 2333 19585 2367 19600
rect 2406 19585 2440 19600
rect 2479 19585 2513 19600
rect 2552 19585 2586 19600
rect 2625 19585 2659 19600
rect 2698 19585 2732 19600
rect 2771 19585 2805 19600
rect 2844 19585 2878 19600
rect 2917 19585 2951 19600
rect 2990 19585 3024 19600
rect 3063 19585 3097 19600
rect 3136 19585 3170 19600
rect 3209 19585 3243 19600
rect 3282 19585 3316 19600
rect 70 19566 77 19585
rect 77 19566 104 19585
rect 143 19566 146 19585
rect 146 19566 177 19585
rect 216 19566 249 19585
rect 249 19566 250 19585
rect 289 19566 318 19585
rect 318 19566 323 19585
rect 362 19566 387 19585
rect 387 19566 396 19585
rect 435 19566 456 19585
rect 456 19566 469 19585
rect 508 19566 525 19585
rect 525 19566 542 19585
rect 581 19566 594 19585
rect 594 19566 615 19585
rect 654 19566 663 19585
rect 663 19566 688 19585
rect 727 19566 732 19585
rect 732 19566 761 19585
rect 800 19566 801 19585
rect 801 19566 834 19585
rect 873 19566 905 19585
rect 905 19566 907 19585
rect 946 19566 974 19585
rect 974 19566 980 19585
rect 1019 19566 1043 19585
rect 1043 19566 1053 19585
rect 1092 19566 1112 19585
rect 1112 19566 1126 19585
rect 1165 19566 1181 19585
rect 1181 19566 1199 19585
rect 1238 19566 1250 19585
rect 1250 19566 1272 19585
rect 1311 19566 1319 19585
rect 1319 19566 1345 19585
rect 1384 19566 1388 19585
rect 1388 19566 1418 19585
rect 1457 19566 1491 19585
rect 1530 19566 1560 19585
rect 1560 19566 1564 19585
rect 1603 19566 1629 19585
rect 1629 19566 1637 19585
rect 1676 19566 1698 19585
rect 1698 19566 1710 19585
rect 1749 19566 1767 19585
rect 1767 19566 1783 19585
rect 1822 19566 1836 19585
rect 1836 19566 1856 19585
rect 1895 19566 1905 19585
rect 1905 19566 1929 19585
rect 1968 19566 1974 19585
rect 1974 19566 2002 19585
rect 2041 19566 2043 19585
rect 2043 19566 2075 19585
rect 2114 19566 2147 19585
rect 2147 19566 2148 19585
rect 2187 19566 2216 19585
rect 2216 19566 2221 19585
rect 2260 19566 2285 19585
rect 2285 19566 2294 19585
rect 2333 19566 2354 19585
rect 2354 19566 2367 19585
rect 2406 19566 2423 19585
rect 2423 19566 2440 19585
rect 2479 19566 2492 19585
rect 2492 19566 2513 19585
rect 2552 19566 2561 19585
rect 2561 19566 2586 19585
rect 2625 19566 2630 19585
rect 2630 19566 2659 19585
rect 2698 19566 2699 19585
rect 2699 19566 2732 19585
rect 2771 19566 2802 19585
rect 2802 19566 2805 19585
rect 2844 19566 2871 19585
rect 2871 19566 2878 19585
rect 2917 19566 2940 19585
rect 2940 19566 2951 19585
rect 2990 19566 3009 19585
rect 3009 19566 3024 19585
rect 3063 19566 3078 19585
rect 3078 19566 3097 19585
rect 3136 19566 3147 19585
rect 3147 19566 3170 19585
rect 3209 19566 3216 19585
rect 3216 19566 3243 19585
rect 3282 19566 3285 19585
rect 3285 19566 3316 19585
rect 3354 19566 3388 19600
rect 3426 19585 3460 19600
rect 3498 19585 3532 19600
rect 3570 19585 3604 19600
rect 3642 19585 3676 19600
rect 3714 19585 3748 19600
rect 3786 19585 3820 19600
rect 3858 19585 3892 19600
rect 3930 19585 3964 19600
rect 4002 19585 4036 19600
rect 4074 19585 4108 19600
rect 4146 19585 4180 19600
rect 4218 19585 4252 19600
rect 4290 19585 4324 19600
rect 4362 19585 4396 19600
rect 4434 19585 4468 19600
rect 4506 19585 4540 19600
rect 4578 19585 4612 19600
rect 4650 19585 4684 19600
rect 4722 19585 4756 19600
rect 4794 19585 4828 19600
rect 4866 19585 4900 19600
rect 4938 19585 4972 19600
rect 5010 19585 5044 19600
rect 5082 19585 5116 19600
rect 5154 19585 5188 19600
rect 5226 19585 5260 19600
rect 5298 19585 5332 19600
rect 5370 19585 5404 19600
rect 5442 19585 5476 19600
rect 5514 19585 5548 19600
rect 5586 19585 5620 19600
rect 5658 19585 5692 19600
rect 5730 19585 5764 19600
rect 5802 19585 5836 19600
rect 5874 19585 5908 19600
rect 5946 19585 5980 19600
rect 6018 19585 6052 19600
rect 6090 19585 6124 19600
rect 6162 19585 6196 19600
rect 6234 19585 6268 19600
rect 6306 19585 6340 19600
rect 6378 19585 6412 19600
rect 6450 19585 6484 19600
rect 6522 19585 6556 19600
rect 6594 19585 6628 19600
rect 6666 19585 6700 19600
rect 6738 19585 6772 19600
rect 6810 19585 6844 19600
rect 6882 19585 6916 19600
rect 6954 19585 6988 19600
rect 7026 19585 7060 19600
rect 7098 19585 7132 19600
rect 7170 19585 7204 19600
rect 7242 19585 7276 19600
rect 7314 19585 7348 19600
rect 7386 19585 7420 19600
rect 7458 19585 7492 19600
rect 7530 19585 7564 19600
rect 7602 19585 7636 19600
rect 7674 19585 7708 19600
rect 7746 19585 7780 19600
rect 7818 19585 7852 19600
rect 7890 19585 7924 19600
rect 7962 19585 7996 19600
rect 8034 19585 8068 19600
rect 8106 19585 8140 19600
rect 8178 19585 8212 19600
rect 8250 19585 8284 19600
rect 8322 19585 8356 19600
rect 8394 19585 8428 19600
rect 8466 19585 8500 19600
rect 8538 19585 8572 19600
rect 8610 19585 8644 19600
rect 8682 19585 8716 19600
rect 8754 19585 8788 19600
rect 8826 19585 8860 19600
rect 8898 19585 8932 19600
rect 8970 19585 9004 19600
rect 9042 19585 9076 19600
rect 9114 19585 9148 19600
rect 9186 19585 9220 19600
rect 9258 19585 9292 19600
rect 9330 19585 9364 19600
rect 9402 19585 9436 19600
rect 9474 19585 9508 19600
rect 9546 19585 9580 19600
rect 9618 19585 9652 19600
rect 9690 19585 9724 19600
rect 9762 19585 9796 19600
rect 9834 19585 9868 19600
rect 9906 19585 9940 19600
rect 9978 19585 10012 19600
rect 10050 19585 10084 19600
rect 10122 19585 10156 19600
rect 10194 19585 10228 19600
rect 10266 19585 10300 19600
rect 10338 19585 10372 19600
rect 10410 19585 10444 19600
rect 10482 19585 10516 19600
rect 10554 19585 10588 19600
rect 10626 19585 10660 19600
rect 10698 19585 10732 19600
rect 10770 19585 10804 19600
rect 10842 19585 10876 19600
rect 10914 19585 10948 19600
rect 10986 19585 11020 19600
rect 11058 19585 11092 19600
rect 11130 19585 11164 19600
rect 11202 19585 11236 19600
rect 11274 19585 11308 19600
rect 11346 19585 11380 19600
rect 11418 19585 11452 19600
rect 11490 19585 11524 19600
rect 11562 19585 11596 19600
rect 11634 19585 11668 19600
rect 11706 19585 11740 19600
rect 3426 19566 3458 19585
rect 3458 19566 3460 19585
rect 3498 19566 3527 19585
rect 3527 19566 3532 19585
rect 3570 19566 3596 19585
rect 3596 19566 3604 19585
rect 3642 19566 3665 19585
rect 3665 19566 3676 19585
rect 3714 19566 3733 19585
rect 3733 19566 3748 19585
rect 3786 19566 3801 19585
rect 3801 19566 3820 19585
rect 3858 19566 3869 19585
rect 3869 19566 3892 19585
rect 3930 19566 3937 19585
rect 3937 19566 3964 19585
rect 4002 19566 4005 19585
rect 4005 19566 4036 19585
rect 4074 19566 4107 19585
rect 4107 19566 4108 19585
rect 4146 19566 4175 19585
rect 4175 19566 4180 19585
rect 4218 19566 4243 19585
rect 4243 19566 4252 19585
rect 4290 19566 4311 19585
rect 4311 19566 4324 19585
rect 4362 19566 4379 19585
rect 4379 19566 4396 19585
rect 4434 19566 4447 19585
rect 4447 19566 4468 19585
rect 4506 19566 4515 19585
rect 4515 19566 4540 19585
rect 4578 19566 4583 19585
rect 4583 19566 4612 19585
rect 4650 19566 4651 19585
rect 4651 19566 4684 19585
rect 4722 19566 4753 19585
rect 4753 19566 4756 19585
rect 4794 19566 4821 19585
rect 4821 19566 4828 19585
rect 4866 19566 4889 19585
rect 4889 19566 4900 19585
rect 4938 19566 4957 19585
rect 4957 19566 4972 19585
rect 5010 19566 5025 19585
rect 5025 19566 5044 19585
rect 5082 19566 5093 19585
rect 5093 19566 5116 19585
rect 5154 19566 5161 19585
rect 5161 19566 5188 19585
rect 5226 19566 5229 19585
rect 5229 19566 5260 19585
rect 5298 19566 5331 19585
rect 5331 19566 5332 19585
rect 5370 19566 5399 19585
rect 5399 19566 5404 19585
rect 5442 19566 5467 19585
rect 5467 19566 5476 19585
rect 5514 19566 5535 19585
rect 5535 19566 5548 19585
rect 5586 19566 5603 19585
rect 5603 19566 5620 19585
rect 5658 19566 5671 19585
rect 5671 19566 5692 19585
rect 5730 19566 5739 19585
rect 5739 19566 5764 19585
rect 5802 19566 5807 19585
rect 5807 19566 5836 19585
rect 5874 19566 5875 19585
rect 5875 19566 5908 19585
rect 5946 19566 5977 19585
rect 5977 19566 5980 19585
rect 6018 19566 6045 19585
rect 6045 19566 6052 19585
rect 6090 19566 6113 19585
rect 6113 19566 6124 19585
rect 6162 19566 6181 19585
rect 6181 19566 6196 19585
rect 6234 19566 6249 19585
rect 6249 19566 6268 19585
rect 6306 19566 6317 19585
rect 6317 19566 6340 19585
rect 6378 19566 6385 19585
rect 6385 19566 6412 19585
rect 6450 19566 6453 19585
rect 6453 19566 6484 19585
rect 6522 19566 6555 19585
rect 6555 19566 6556 19585
rect 6594 19566 6623 19585
rect 6623 19566 6628 19585
rect 6666 19566 6691 19585
rect 6691 19566 6700 19585
rect 6738 19566 6759 19585
rect 6759 19566 6772 19585
rect 6810 19566 6827 19585
rect 6827 19566 6844 19585
rect 6882 19566 6895 19585
rect 6895 19566 6916 19585
rect 6954 19566 6963 19585
rect 6963 19566 6988 19585
rect 7026 19566 7031 19585
rect 7031 19566 7060 19585
rect 7098 19566 7099 19585
rect 7099 19566 7132 19585
rect 7170 19566 7201 19585
rect 7201 19566 7204 19585
rect 7242 19566 7269 19585
rect 7269 19566 7276 19585
rect 7314 19566 7337 19585
rect 7337 19566 7348 19585
rect 7386 19566 7405 19585
rect 7405 19566 7420 19585
rect 7458 19566 7473 19585
rect 7473 19566 7492 19585
rect 7530 19566 7541 19585
rect 7541 19566 7564 19585
rect 7602 19566 7609 19585
rect 7609 19566 7636 19585
rect 7674 19566 7677 19585
rect 7677 19566 7708 19585
rect 7746 19566 7779 19585
rect 7779 19566 7780 19585
rect 7818 19566 7847 19585
rect 7847 19566 7852 19585
rect 7890 19566 7915 19585
rect 7915 19566 7924 19585
rect 7962 19566 7983 19585
rect 7983 19566 7996 19585
rect 8034 19566 8051 19585
rect 8051 19566 8068 19585
rect 8106 19566 8119 19585
rect 8119 19566 8140 19585
rect 8178 19566 8187 19585
rect 8187 19566 8212 19585
rect 8250 19566 8255 19585
rect 8255 19566 8284 19585
rect 8322 19566 8323 19585
rect 8323 19566 8356 19585
rect 8394 19566 8425 19585
rect 8425 19566 8428 19585
rect 8466 19566 8493 19585
rect 8493 19566 8500 19585
rect 8538 19566 8561 19585
rect 8561 19566 8572 19585
rect 8610 19566 8629 19585
rect 8629 19566 8644 19585
rect 8682 19566 8697 19585
rect 8697 19566 8716 19585
rect 8754 19566 8765 19585
rect 8765 19566 8788 19585
rect 8826 19566 8833 19585
rect 8833 19566 8860 19585
rect 8898 19566 8901 19585
rect 8901 19566 8932 19585
rect 8970 19566 9003 19585
rect 9003 19566 9004 19585
rect 9042 19566 9071 19585
rect 9071 19566 9076 19585
rect 9114 19566 9139 19585
rect 9139 19566 9148 19585
rect 9186 19566 9207 19585
rect 9207 19566 9220 19585
rect 9258 19566 9275 19585
rect 9275 19566 9292 19585
rect 9330 19566 9343 19585
rect 9343 19566 9364 19585
rect 9402 19566 9411 19585
rect 9411 19566 9436 19585
rect 9474 19566 9479 19585
rect 9479 19566 9508 19585
rect 9546 19566 9547 19585
rect 9547 19566 9580 19585
rect 9618 19566 9649 19585
rect 9649 19566 9652 19585
rect 9690 19566 9717 19585
rect 9717 19566 9724 19585
rect 9762 19566 9785 19585
rect 9785 19566 9796 19585
rect 9834 19566 9853 19585
rect 9853 19566 9868 19585
rect 9906 19566 9921 19585
rect 9921 19566 9940 19585
rect 9978 19566 9989 19585
rect 9989 19566 10012 19585
rect 10050 19566 10057 19585
rect 10057 19566 10084 19585
rect 10122 19566 10125 19585
rect 10125 19566 10156 19585
rect 10194 19566 10227 19585
rect 10227 19566 10228 19585
rect 10266 19566 10295 19585
rect 10295 19566 10300 19585
rect 10338 19566 10363 19585
rect 10363 19566 10372 19585
rect 10410 19566 10431 19585
rect 10431 19566 10444 19585
rect 10482 19566 10499 19585
rect 10499 19566 10516 19585
rect 10554 19566 10567 19585
rect 10567 19566 10588 19585
rect 10626 19566 10635 19585
rect 10635 19566 10660 19585
rect 10698 19566 10703 19585
rect 10703 19566 10732 19585
rect 10770 19566 10771 19585
rect 10771 19566 10804 19585
rect 10842 19566 10873 19585
rect 10873 19566 10876 19585
rect 10914 19566 10941 19585
rect 10941 19566 10948 19585
rect 10986 19566 11009 19585
rect 11009 19566 11020 19585
rect 11058 19566 11077 19585
rect 11077 19566 11092 19585
rect 11130 19566 11145 19585
rect 11145 19566 11164 19585
rect 11202 19566 11213 19585
rect 11213 19566 11236 19585
rect 11274 19566 11281 19585
rect 11281 19566 11308 19585
rect 11346 19566 11349 19585
rect 11349 19566 11380 19585
rect 11418 19566 11451 19585
rect 11451 19566 11452 19585
rect 11490 19566 11519 19585
rect 11519 19566 11524 19585
rect 11562 19566 11587 19585
rect 11587 19566 11596 19585
rect 11634 19566 11655 19585
rect 11655 19566 11668 19585
rect 11706 19566 11723 19585
rect 11723 19566 11740 19585
rect 11778 19566 11812 19600
rect 11850 19566 11884 19600
rect 11922 19566 11956 19600
rect 11994 19566 12028 19600
rect 12066 19566 12100 19600
rect 12138 19566 12172 19600
rect 12210 19566 12244 19600
rect 12282 19566 12316 19600
rect 12354 19566 12388 19600
rect 12426 19566 12460 19600
rect 12498 19566 12532 19600
rect 12570 19566 12604 19600
rect 12642 19566 12676 19600
rect 12714 19566 12748 19600
rect 12786 19566 12820 19600
rect 12858 19566 12892 19600
rect 12930 19566 12964 19600
rect 13002 19566 13036 19600
rect 13074 19566 13108 19600
rect 13146 19566 13180 19600
rect 13218 19566 13252 19600
rect 13290 19566 13324 19600
rect 13362 19566 13396 19600
rect 13434 19566 13468 19600
rect 13506 19566 13540 19600
rect 13578 19566 13612 19600
rect 13650 19566 13684 19600
rect 13722 19566 13756 19600
rect 13794 19566 13828 19600
rect 13866 19566 13900 19600
rect 13938 19566 13972 19600
rect 14010 19566 14044 19600
rect 14082 19566 14116 19600
rect 14154 19566 14188 19600
rect 14226 19566 14260 19600
rect 14298 19566 14332 19600
rect 14370 19566 14404 19600
rect 14442 19566 14476 19600
rect 14514 19587 14518 19600
rect 14518 19587 14548 19600
rect 14586 19587 14601 19600
rect 14601 19587 14620 19600
rect 14658 19587 14684 19600
rect 14684 19587 14692 19600
rect 14514 19566 14548 19587
rect 14586 19566 14620 19587
rect 14658 19566 14692 19587
rect 14730 19587 14733 19600
rect 14733 19587 14764 19600
rect 14802 19587 14816 19600
rect 14816 19587 14836 19600
rect 14730 19566 14764 19587
rect 14802 19566 14836 19587
rect 14874 19566 14908 19600
rect 209 18379 243 18382
rect 282 18379 316 18382
rect 355 18379 389 18382
rect 428 18379 462 18382
rect 501 18379 535 18382
rect 574 18379 608 18382
rect 647 18379 681 18382
rect 720 18379 754 18382
rect 793 18379 827 18382
rect 866 18379 900 18382
rect 939 18379 973 18382
rect 1012 18379 1046 18382
rect 1085 18379 1119 18382
rect 1158 18379 1192 18382
rect 1231 18379 1265 18382
rect 1304 18379 1338 18382
rect 1377 18379 1411 18382
rect 1450 18379 1484 18382
rect 1523 18379 1557 18382
rect 1596 18379 1630 18382
rect 1669 18379 1703 18382
rect 1742 18379 1776 18382
rect 1815 18379 1849 18382
rect 1888 18379 1922 18382
rect 1961 18379 1995 18382
rect 2034 18379 2068 18382
rect 2107 18379 2141 18382
rect 2180 18379 2214 18382
rect 2253 18379 2287 18382
rect 2326 18379 2360 18382
rect 2399 18379 2433 18382
rect 2472 18379 2506 18382
rect 2545 18379 2579 18382
rect 2618 18379 2652 18382
rect 2691 18379 2725 18382
rect 2764 18379 2798 18382
rect 2837 18379 2871 18382
rect 2910 18379 2944 18382
rect 2983 18379 3017 18382
rect 3056 18379 3090 18382
rect 3129 18379 3163 18382
rect 3202 18379 3236 18382
rect 3275 18379 3309 18382
rect 3348 18379 3382 18382
rect 3421 18379 3455 18382
rect 3494 18379 3528 18382
rect 3566 18379 3600 18382
rect 3638 18379 3672 18382
rect 3710 18379 3744 18382
rect 3782 18379 3816 18382
rect 3854 18379 3888 18382
rect 3926 18379 3960 18382
rect 3998 18379 4032 18382
rect 4070 18379 4104 18382
rect 4142 18379 4176 18382
rect 4214 18379 4248 18382
rect 4286 18379 4320 18382
rect 4358 18379 4392 18382
rect 4430 18379 4464 18382
rect 4502 18379 4536 18382
rect 4574 18379 4608 18382
rect 4646 18379 4680 18382
rect 4718 18379 4752 18382
rect 4790 18379 4824 18382
rect 4862 18379 4896 18382
rect 4934 18379 4968 18382
rect 5006 18379 5040 18382
rect 5078 18379 5112 18382
rect 5150 18379 5184 18382
rect 5222 18379 5256 18382
rect 5294 18379 5328 18382
rect 5366 18379 5400 18382
rect 5438 18379 5472 18382
rect 5510 18379 5544 18382
rect 5582 18379 5616 18382
rect 5654 18379 5688 18382
rect 5726 18379 5760 18382
rect 5798 18379 5832 18382
rect 5870 18379 5904 18382
rect 5942 18379 5976 18382
rect 6014 18379 6048 18382
rect 6086 18379 6120 18382
rect 6158 18379 6192 18382
rect 6230 18379 6264 18382
rect 6302 18379 6336 18382
rect 6374 18379 6408 18382
rect 6446 18379 6480 18382
rect 6518 18379 6552 18382
rect 6590 18379 6624 18382
rect 6662 18379 6696 18382
rect 6734 18379 6768 18382
rect 6806 18379 6840 18382
rect 6878 18379 6912 18382
rect 6950 18379 6984 18382
rect 7022 18379 7056 18382
rect 7094 18379 7128 18382
rect 7166 18379 7200 18382
rect 7238 18379 7272 18382
rect 7310 18379 7344 18382
rect 7382 18379 7416 18382
rect 7454 18379 7488 18382
rect 7526 18379 7560 18382
rect 7598 18379 7632 18382
rect 7670 18379 7704 18382
rect 7742 18379 7776 18382
rect 7814 18379 7848 18382
rect 7886 18379 7920 18382
rect 7958 18379 7992 18382
rect 8030 18379 8064 18382
rect 8102 18379 8136 18382
rect 8174 18379 8208 18382
rect 8246 18379 8280 18382
rect 8318 18379 8352 18382
rect 8390 18379 8424 18382
rect 8462 18379 8496 18382
rect 8534 18379 8568 18382
rect 8606 18379 8640 18382
rect 8678 18379 8712 18382
rect 8750 18379 8784 18382
rect 8822 18379 8856 18382
rect 8894 18379 8928 18382
rect 8966 18379 9000 18382
rect 9038 18379 9072 18382
rect 9110 18379 9144 18382
rect 9182 18379 9216 18382
rect 9254 18379 9288 18382
rect 9326 18379 9360 18382
rect 9398 18379 9432 18382
rect 9470 18379 9504 18382
rect 9542 18379 9576 18382
rect 9614 18379 9648 18382
rect 9686 18379 9720 18382
rect 9758 18379 9792 18382
rect 9830 18379 9864 18382
rect 9902 18379 9936 18382
rect 9974 18379 10008 18382
rect 10046 18379 10080 18382
rect 10118 18379 10152 18382
rect 10190 18379 10224 18382
rect 10262 18379 10296 18382
rect 10334 18379 10368 18382
rect 10406 18379 10440 18382
rect 10478 18379 10512 18382
rect 10550 18379 10584 18382
rect 10622 18379 10656 18382
rect 10694 18379 10728 18382
rect 10766 18379 10800 18382
rect 10838 18379 10872 18382
rect 10910 18379 10944 18382
rect 10982 18379 11016 18382
rect 11054 18379 11088 18382
rect 11126 18379 11160 18382
rect 11198 18379 11232 18382
rect 11270 18379 11304 18382
rect 11342 18379 11376 18382
rect 11414 18379 11448 18382
rect 11486 18379 11520 18382
rect 11558 18379 11592 18382
rect 11630 18379 11664 18382
rect 11702 18379 11736 18382
rect 11774 18379 11808 18382
rect 11846 18379 11880 18382
rect 11918 18379 11952 18382
rect 11990 18379 12024 18382
rect 12062 18379 12096 18382
rect 12134 18379 12168 18382
rect 12206 18379 12240 18382
rect 12278 18379 12312 18382
rect 12350 18379 12384 18382
rect 12422 18379 12456 18382
rect 12494 18379 12528 18382
rect 12566 18379 12600 18382
rect 12638 18379 12672 18382
rect 12710 18379 12744 18382
rect 12782 18379 12816 18382
rect 12854 18379 12888 18382
rect 12926 18379 12960 18382
rect 12998 18379 13032 18382
rect 13070 18379 13104 18382
rect 13142 18379 13176 18382
rect 13214 18379 13248 18382
rect 13286 18379 13320 18382
rect 13358 18379 13392 18382
rect 13430 18379 13464 18382
rect 13502 18379 13536 18382
rect 13574 18379 13608 18382
rect 13646 18379 13680 18382
rect 13718 18379 13752 18382
rect 13790 18379 13824 18382
rect 13862 18379 13896 18382
rect 13934 18379 13968 18382
rect 14006 18379 14040 18382
rect 14078 18379 14112 18382
rect 14150 18379 14184 18382
rect 14222 18379 14256 18382
rect 14294 18379 14328 18382
rect 14366 18379 14400 18382
rect 14438 18379 14472 18382
rect 14510 18379 14544 18382
rect 14582 18379 14616 18382
rect 14654 18379 14688 18382
rect 14726 18379 14760 18382
rect 209 18348 221 18379
rect 221 18348 243 18379
rect 282 18348 290 18379
rect 290 18348 316 18379
rect 355 18348 359 18379
rect 359 18348 389 18379
rect 428 18348 461 18379
rect 461 18348 462 18379
rect 501 18348 529 18379
rect 529 18348 535 18379
rect 574 18348 597 18379
rect 597 18348 608 18379
rect 647 18348 665 18379
rect 665 18348 681 18379
rect 720 18348 733 18379
rect 733 18348 754 18379
rect 793 18348 801 18379
rect 801 18348 827 18379
rect 866 18348 869 18379
rect 869 18348 900 18379
rect 939 18348 971 18379
rect 971 18348 973 18379
rect 1012 18348 1039 18379
rect 1039 18348 1046 18379
rect 1085 18348 1107 18379
rect 1107 18348 1119 18379
rect 1158 18348 1175 18379
rect 1175 18348 1192 18379
rect 1231 18348 1243 18379
rect 1243 18348 1265 18379
rect 1304 18348 1311 18379
rect 1311 18348 1338 18379
rect 1377 18348 1379 18379
rect 1379 18348 1411 18379
rect 1450 18348 1481 18379
rect 1481 18348 1484 18379
rect 1523 18348 1549 18379
rect 1549 18348 1557 18379
rect 1596 18348 1617 18379
rect 1617 18348 1630 18379
rect 1669 18348 1685 18379
rect 1685 18348 1703 18379
rect 1742 18348 1753 18379
rect 1753 18348 1776 18379
rect 1815 18348 1821 18379
rect 1821 18348 1849 18379
rect 1888 18348 1889 18379
rect 1889 18348 1922 18379
rect 1961 18348 1991 18379
rect 1991 18348 1995 18379
rect 2034 18348 2059 18379
rect 2059 18348 2068 18379
rect 2107 18348 2127 18379
rect 2127 18348 2141 18379
rect 2180 18348 2195 18379
rect 2195 18348 2214 18379
rect 2253 18348 2263 18379
rect 2263 18348 2287 18379
rect 2326 18348 2331 18379
rect 2331 18348 2360 18379
rect 2399 18348 2433 18379
rect 2472 18348 2501 18379
rect 2501 18348 2506 18379
rect 2545 18348 2569 18379
rect 2569 18348 2579 18379
rect 2618 18348 2637 18379
rect 2637 18348 2652 18379
rect 2691 18348 2705 18379
rect 2705 18348 2725 18379
rect 2764 18348 2773 18379
rect 2773 18348 2798 18379
rect 2837 18348 2841 18379
rect 2841 18348 2871 18379
rect 2910 18348 2943 18379
rect 2943 18348 2944 18379
rect 2983 18348 3011 18379
rect 3011 18348 3017 18379
rect 3056 18348 3079 18379
rect 3079 18348 3090 18379
rect 3129 18348 3147 18379
rect 3147 18348 3163 18379
rect 3202 18348 3215 18379
rect 3215 18348 3236 18379
rect 3275 18348 3283 18379
rect 3283 18348 3309 18379
rect 3348 18348 3351 18379
rect 3351 18348 3382 18379
rect 3421 18348 3453 18379
rect 3453 18348 3455 18379
rect 3494 18348 3521 18379
rect 3521 18348 3528 18379
rect 3566 18348 3589 18379
rect 3589 18348 3600 18379
rect 3638 18348 3657 18379
rect 3657 18348 3672 18379
rect 3710 18348 3725 18379
rect 3725 18348 3744 18379
rect 3782 18348 3793 18379
rect 3793 18348 3816 18379
rect 3854 18348 3861 18379
rect 3861 18348 3888 18379
rect 3926 18348 3929 18379
rect 3929 18348 3960 18379
rect 3998 18348 4031 18379
rect 4031 18348 4032 18379
rect 4070 18348 4099 18379
rect 4099 18348 4104 18379
rect 4142 18348 4167 18379
rect 4167 18348 4176 18379
rect 4214 18348 4235 18379
rect 4235 18348 4248 18379
rect 4286 18348 4303 18379
rect 4303 18348 4320 18379
rect 4358 18348 4371 18379
rect 4371 18348 4392 18379
rect 4430 18348 4439 18379
rect 4439 18348 4464 18379
rect 4502 18348 4507 18379
rect 4507 18348 4536 18379
rect 4574 18348 4575 18379
rect 4575 18348 4608 18379
rect 4646 18348 4677 18379
rect 4677 18348 4680 18379
rect 4718 18348 4745 18379
rect 4745 18348 4752 18379
rect 4790 18348 4813 18379
rect 4813 18348 4824 18379
rect 4862 18348 4881 18379
rect 4881 18348 4896 18379
rect 4934 18348 4949 18379
rect 4949 18348 4968 18379
rect 5006 18348 5017 18379
rect 5017 18348 5040 18379
rect 5078 18348 5085 18379
rect 5085 18348 5112 18379
rect 5150 18348 5153 18379
rect 5153 18348 5184 18379
rect 5222 18348 5255 18379
rect 5255 18348 5256 18379
rect 5294 18348 5323 18379
rect 5323 18348 5328 18379
rect 5366 18348 5391 18379
rect 5391 18348 5400 18379
rect 5438 18348 5459 18379
rect 5459 18348 5472 18379
rect 5510 18348 5527 18379
rect 5527 18348 5544 18379
rect 5582 18348 5595 18379
rect 5595 18348 5616 18379
rect 5654 18348 5663 18379
rect 5663 18348 5688 18379
rect 5726 18348 5731 18379
rect 5731 18348 5760 18379
rect 5798 18348 5799 18379
rect 5799 18348 5832 18379
rect 5870 18348 5901 18379
rect 5901 18348 5904 18379
rect 5942 18348 5969 18379
rect 5969 18348 5976 18379
rect 6014 18348 6037 18379
rect 6037 18348 6048 18379
rect 6086 18348 6105 18379
rect 6105 18348 6120 18379
rect 6158 18348 6173 18379
rect 6173 18348 6192 18379
rect 6230 18348 6241 18379
rect 6241 18348 6264 18379
rect 6302 18348 6309 18379
rect 6309 18348 6336 18379
rect 6374 18348 6377 18379
rect 6377 18348 6408 18379
rect 6446 18348 6479 18379
rect 6479 18348 6480 18379
rect 6518 18348 6547 18379
rect 6547 18348 6552 18379
rect 6590 18348 6615 18379
rect 6615 18348 6624 18379
rect 6662 18348 6683 18379
rect 6683 18348 6696 18379
rect 6734 18348 6751 18379
rect 6751 18348 6768 18379
rect 6806 18348 6819 18379
rect 6819 18348 6840 18379
rect 6878 18348 6887 18379
rect 6887 18348 6912 18379
rect 6950 18348 6955 18379
rect 6955 18348 6984 18379
rect 7022 18348 7023 18379
rect 7023 18348 7056 18379
rect 7094 18348 7125 18379
rect 7125 18348 7128 18379
rect 7166 18348 7193 18379
rect 7193 18348 7200 18379
rect 7238 18348 7261 18379
rect 7261 18348 7272 18379
rect 7310 18348 7329 18379
rect 7329 18348 7344 18379
rect 7382 18348 7397 18379
rect 7397 18348 7416 18379
rect 7454 18348 7465 18379
rect 7465 18348 7488 18379
rect 7526 18348 7533 18379
rect 7533 18348 7560 18379
rect 7598 18348 7601 18379
rect 7601 18348 7632 18379
rect 7670 18348 7703 18379
rect 7703 18348 7704 18379
rect 7742 18348 7771 18379
rect 7771 18348 7776 18379
rect 7814 18348 7839 18379
rect 7839 18348 7848 18379
rect 7886 18348 7907 18379
rect 7907 18348 7920 18379
rect 7958 18348 7975 18379
rect 7975 18348 7992 18379
rect 8030 18348 8043 18379
rect 8043 18348 8064 18379
rect 8102 18348 8111 18379
rect 8111 18348 8136 18379
rect 8174 18348 8179 18379
rect 8179 18348 8208 18379
rect 8246 18348 8247 18379
rect 8247 18348 8280 18379
rect 8318 18348 8349 18379
rect 8349 18348 8352 18379
rect 8390 18348 8417 18379
rect 8417 18348 8424 18379
rect 8462 18348 8485 18379
rect 8485 18348 8496 18379
rect 8534 18348 8553 18379
rect 8553 18348 8568 18379
rect 8606 18348 8621 18379
rect 8621 18348 8640 18379
rect 8678 18348 8689 18379
rect 8689 18348 8712 18379
rect 8750 18348 8757 18379
rect 8757 18348 8784 18379
rect 8822 18348 8825 18379
rect 8825 18348 8856 18379
rect 8894 18348 8927 18379
rect 8927 18348 8928 18379
rect 8966 18348 8995 18379
rect 8995 18348 9000 18379
rect 9038 18348 9063 18379
rect 9063 18348 9072 18379
rect 9110 18348 9131 18379
rect 9131 18348 9144 18379
rect 9182 18348 9199 18379
rect 9199 18348 9216 18379
rect 9254 18348 9267 18379
rect 9267 18348 9288 18379
rect 9326 18348 9335 18379
rect 9335 18348 9360 18379
rect 9398 18348 9403 18379
rect 9403 18348 9432 18379
rect 9470 18348 9471 18379
rect 9471 18348 9504 18379
rect 9542 18348 9573 18379
rect 9573 18348 9576 18379
rect 9614 18348 9641 18379
rect 9641 18348 9648 18379
rect 9686 18348 9709 18379
rect 9709 18348 9720 18379
rect 9758 18348 9777 18379
rect 9777 18348 9792 18379
rect 9830 18348 9845 18379
rect 9845 18348 9864 18379
rect 9902 18348 9913 18379
rect 9913 18348 9936 18379
rect 9974 18348 9981 18379
rect 9981 18348 10008 18379
rect 10046 18348 10049 18379
rect 10049 18348 10080 18379
rect 10118 18348 10151 18379
rect 10151 18348 10152 18379
rect 10190 18348 10219 18379
rect 10219 18348 10224 18379
rect 10262 18348 10287 18379
rect 10287 18348 10296 18379
rect 10334 18348 10355 18379
rect 10355 18348 10368 18379
rect 10406 18348 10423 18379
rect 10423 18348 10440 18379
rect 10478 18348 10491 18379
rect 10491 18348 10512 18379
rect 10550 18348 10559 18379
rect 10559 18348 10584 18379
rect 10622 18348 10627 18379
rect 10627 18348 10656 18379
rect 10694 18348 10695 18379
rect 10695 18348 10728 18379
rect 10766 18348 10797 18379
rect 10797 18348 10800 18379
rect 10838 18348 10865 18379
rect 10865 18348 10872 18379
rect 10910 18348 10933 18379
rect 10933 18348 10944 18379
rect 10982 18348 11001 18379
rect 11001 18348 11016 18379
rect 11054 18348 11069 18379
rect 11069 18348 11088 18379
rect 11126 18348 11137 18379
rect 11137 18348 11160 18379
rect 11198 18348 11205 18379
rect 11205 18348 11232 18379
rect 11270 18348 11273 18379
rect 11273 18348 11304 18379
rect 11342 18348 11375 18379
rect 11375 18348 11376 18379
rect 11414 18348 11443 18379
rect 11443 18348 11448 18379
rect 11486 18348 11511 18379
rect 11511 18348 11520 18379
rect 11558 18348 11579 18379
rect 11579 18348 11592 18379
rect 11630 18348 11647 18379
rect 11647 18348 11664 18379
rect 11702 18348 11715 18379
rect 11715 18348 11736 18379
rect 11774 18348 11783 18379
rect 11783 18348 11808 18379
rect 11846 18348 11851 18379
rect 11851 18348 11880 18379
rect 11918 18348 11919 18379
rect 11919 18348 11952 18379
rect 11990 18348 12021 18379
rect 12021 18348 12024 18379
rect 12062 18348 12089 18379
rect 12089 18348 12096 18379
rect 12134 18348 12157 18379
rect 12157 18348 12168 18379
rect 12206 18348 12225 18379
rect 12225 18348 12240 18379
rect 12278 18348 12293 18379
rect 12293 18348 12312 18379
rect 12350 18348 12361 18379
rect 12361 18348 12384 18379
rect 12422 18348 12429 18379
rect 12429 18348 12456 18379
rect 12494 18348 12497 18379
rect 12497 18348 12528 18379
rect 12566 18348 12599 18379
rect 12599 18348 12600 18379
rect 12638 18348 12667 18379
rect 12667 18348 12672 18379
rect 12710 18348 12735 18379
rect 12735 18348 12744 18379
rect 12782 18348 12803 18379
rect 12803 18348 12816 18379
rect 12854 18348 12871 18379
rect 12871 18348 12888 18379
rect 12926 18348 12939 18379
rect 12939 18348 12960 18379
rect 12998 18348 13007 18379
rect 13007 18348 13032 18379
rect 13070 18348 13075 18379
rect 13075 18348 13104 18379
rect 13142 18348 13143 18379
rect 13143 18348 13176 18379
rect 13214 18348 13245 18379
rect 13245 18348 13248 18379
rect 13286 18348 13313 18379
rect 13313 18348 13320 18379
rect 13358 18348 13381 18379
rect 13381 18348 13392 18379
rect 13430 18348 13449 18379
rect 13449 18348 13464 18379
rect 13502 18348 13517 18379
rect 13517 18348 13536 18379
rect 13574 18348 13585 18379
rect 13585 18348 13608 18379
rect 13646 18348 13653 18379
rect 13653 18348 13680 18379
rect 13718 18348 13721 18379
rect 13721 18348 13752 18379
rect 13790 18348 13823 18379
rect 13823 18348 13824 18379
rect 13862 18348 13891 18379
rect 13891 18348 13896 18379
rect 13934 18348 13959 18379
rect 13959 18348 13968 18379
rect 14006 18348 14027 18379
rect 14027 18348 14040 18379
rect 14078 18348 14095 18379
rect 14095 18348 14112 18379
rect 14150 18348 14163 18379
rect 14163 18348 14184 18379
rect 14222 18348 14231 18379
rect 14231 18348 14256 18379
rect 14294 18348 14299 18379
rect 14299 18348 14328 18379
rect 14366 18348 14367 18379
rect 14367 18348 14400 18379
rect 14438 18348 14469 18379
rect 14469 18348 14472 18379
rect 14510 18348 14537 18379
rect 14537 18348 14544 18379
rect 14582 18348 14605 18379
rect 14605 18348 14616 18379
rect 14654 18348 14673 18379
rect 14673 18348 14688 18379
rect 14726 18348 14741 18379
rect 14741 18348 14760 18379
rect 209 18275 221 18306
rect 221 18275 243 18306
rect 282 18275 290 18306
rect 290 18275 316 18306
rect 355 18275 359 18306
rect 359 18275 389 18306
rect 428 18275 461 18306
rect 461 18275 462 18306
rect 501 18275 529 18306
rect 529 18275 535 18306
rect 574 18275 597 18306
rect 597 18275 608 18306
rect 647 18275 665 18306
rect 665 18275 681 18306
rect 720 18275 733 18306
rect 733 18275 754 18306
rect 793 18275 801 18306
rect 801 18275 827 18306
rect 866 18275 869 18306
rect 869 18275 900 18306
rect 939 18275 971 18306
rect 971 18275 973 18306
rect 1012 18275 1039 18306
rect 1039 18275 1046 18306
rect 1085 18275 1107 18306
rect 1107 18275 1119 18306
rect 1158 18275 1175 18306
rect 1175 18275 1192 18306
rect 1231 18275 1243 18306
rect 1243 18275 1265 18306
rect 1304 18275 1311 18306
rect 1311 18275 1338 18306
rect 1377 18275 1379 18306
rect 1379 18275 1411 18306
rect 1450 18275 1481 18306
rect 1481 18275 1484 18306
rect 1523 18275 1549 18306
rect 1549 18275 1557 18306
rect 1596 18275 1617 18306
rect 1617 18275 1630 18306
rect 1669 18275 1685 18306
rect 1685 18275 1703 18306
rect 1742 18275 1753 18306
rect 1753 18275 1776 18306
rect 1815 18275 1821 18306
rect 1821 18275 1849 18306
rect 1888 18275 1889 18306
rect 1889 18275 1922 18306
rect 1961 18275 1991 18306
rect 1991 18275 1995 18306
rect 2034 18275 2059 18306
rect 2059 18275 2068 18306
rect 2107 18275 2127 18306
rect 2127 18275 2141 18306
rect 2180 18275 2195 18306
rect 2195 18275 2214 18306
rect 2253 18275 2263 18306
rect 2263 18275 2287 18306
rect 2326 18275 2331 18306
rect 2331 18275 2360 18306
rect 2399 18275 2433 18306
rect 2472 18275 2501 18306
rect 2501 18275 2506 18306
rect 2545 18275 2569 18306
rect 2569 18275 2579 18306
rect 2618 18275 2637 18306
rect 2637 18275 2652 18306
rect 2691 18275 2705 18306
rect 2705 18275 2725 18306
rect 2764 18275 2773 18306
rect 2773 18275 2798 18306
rect 2837 18275 2841 18306
rect 2841 18275 2871 18306
rect 2910 18275 2943 18306
rect 2943 18275 2944 18306
rect 2983 18275 3011 18306
rect 3011 18275 3017 18306
rect 3056 18275 3079 18306
rect 3079 18275 3090 18306
rect 3129 18275 3147 18306
rect 3147 18275 3163 18306
rect 3202 18275 3215 18306
rect 3215 18275 3236 18306
rect 3275 18275 3283 18306
rect 3283 18275 3309 18306
rect 3348 18275 3351 18306
rect 3351 18275 3382 18306
rect 3421 18275 3453 18306
rect 3453 18275 3455 18306
rect 3494 18275 3521 18306
rect 3521 18275 3528 18306
rect 3566 18275 3589 18306
rect 3589 18275 3600 18306
rect 3638 18275 3657 18306
rect 3657 18275 3672 18306
rect 3710 18275 3725 18306
rect 3725 18275 3744 18306
rect 3782 18275 3793 18306
rect 3793 18275 3816 18306
rect 3854 18275 3861 18306
rect 3861 18275 3888 18306
rect 3926 18275 3929 18306
rect 3929 18275 3960 18306
rect 3998 18275 4031 18306
rect 4031 18275 4032 18306
rect 4070 18275 4099 18306
rect 4099 18275 4104 18306
rect 4142 18275 4167 18306
rect 4167 18275 4176 18306
rect 4214 18275 4235 18306
rect 4235 18275 4248 18306
rect 4286 18275 4303 18306
rect 4303 18275 4320 18306
rect 4358 18275 4371 18306
rect 4371 18275 4392 18306
rect 4430 18275 4439 18306
rect 4439 18275 4464 18306
rect 4502 18275 4507 18306
rect 4507 18275 4536 18306
rect 4574 18275 4575 18306
rect 4575 18275 4608 18306
rect 4646 18275 4677 18306
rect 4677 18275 4680 18306
rect 4718 18275 4745 18306
rect 4745 18275 4752 18306
rect 4790 18275 4813 18306
rect 4813 18275 4824 18306
rect 4862 18275 4881 18306
rect 4881 18275 4896 18306
rect 4934 18275 4949 18306
rect 4949 18275 4968 18306
rect 5006 18275 5017 18306
rect 5017 18275 5040 18306
rect 5078 18275 5085 18306
rect 5085 18275 5112 18306
rect 5150 18275 5153 18306
rect 5153 18275 5184 18306
rect 5222 18275 5255 18306
rect 5255 18275 5256 18306
rect 5294 18275 5323 18306
rect 5323 18275 5328 18306
rect 5366 18275 5391 18306
rect 5391 18275 5400 18306
rect 5438 18275 5459 18306
rect 5459 18275 5472 18306
rect 5510 18275 5527 18306
rect 5527 18275 5544 18306
rect 5582 18275 5595 18306
rect 5595 18275 5616 18306
rect 5654 18275 5663 18306
rect 5663 18275 5688 18306
rect 5726 18275 5731 18306
rect 5731 18275 5760 18306
rect 5798 18275 5799 18306
rect 5799 18275 5832 18306
rect 5870 18275 5901 18306
rect 5901 18275 5904 18306
rect 5942 18275 5969 18306
rect 5969 18275 5976 18306
rect 6014 18275 6037 18306
rect 6037 18275 6048 18306
rect 6086 18275 6105 18306
rect 6105 18275 6120 18306
rect 6158 18275 6173 18306
rect 6173 18275 6192 18306
rect 6230 18275 6241 18306
rect 6241 18275 6264 18306
rect 6302 18275 6309 18306
rect 6309 18275 6336 18306
rect 6374 18275 6377 18306
rect 6377 18275 6408 18306
rect 6446 18275 6479 18306
rect 6479 18275 6480 18306
rect 6518 18275 6547 18306
rect 6547 18275 6552 18306
rect 6590 18275 6615 18306
rect 6615 18275 6624 18306
rect 6662 18275 6683 18306
rect 6683 18275 6696 18306
rect 6734 18275 6751 18306
rect 6751 18275 6768 18306
rect 6806 18275 6819 18306
rect 6819 18275 6840 18306
rect 6878 18275 6887 18306
rect 6887 18275 6912 18306
rect 6950 18275 6955 18306
rect 6955 18275 6984 18306
rect 7022 18275 7023 18306
rect 7023 18275 7056 18306
rect 7094 18275 7125 18306
rect 7125 18275 7128 18306
rect 7166 18275 7193 18306
rect 7193 18275 7200 18306
rect 7238 18275 7261 18306
rect 7261 18275 7272 18306
rect 7310 18275 7329 18306
rect 7329 18275 7344 18306
rect 7382 18275 7397 18306
rect 7397 18275 7416 18306
rect 7454 18275 7465 18306
rect 7465 18275 7488 18306
rect 7526 18275 7533 18306
rect 7533 18275 7560 18306
rect 7598 18275 7601 18306
rect 7601 18275 7632 18306
rect 7670 18275 7703 18306
rect 7703 18275 7704 18306
rect 7742 18275 7771 18306
rect 7771 18275 7776 18306
rect 7814 18275 7839 18306
rect 7839 18275 7848 18306
rect 7886 18275 7907 18306
rect 7907 18275 7920 18306
rect 7958 18275 7975 18306
rect 7975 18275 7992 18306
rect 8030 18275 8043 18306
rect 8043 18275 8064 18306
rect 8102 18275 8111 18306
rect 8111 18275 8136 18306
rect 8174 18275 8179 18306
rect 8179 18275 8208 18306
rect 8246 18275 8247 18306
rect 8247 18275 8280 18306
rect 8318 18275 8349 18306
rect 8349 18275 8352 18306
rect 8390 18275 8417 18306
rect 8417 18275 8424 18306
rect 8462 18275 8485 18306
rect 8485 18275 8496 18306
rect 8534 18275 8553 18306
rect 8553 18275 8568 18306
rect 8606 18275 8621 18306
rect 8621 18275 8640 18306
rect 8678 18275 8689 18306
rect 8689 18275 8712 18306
rect 8750 18275 8757 18306
rect 8757 18275 8784 18306
rect 8822 18275 8825 18306
rect 8825 18275 8856 18306
rect 8894 18275 8927 18306
rect 8927 18275 8928 18306
rect 8966 18275 8995 18306
rect 8995 18275 9000 18306
rect 9038 18275 9063 18306
rect 9063 18275 9072 18306
rect 9110 18275 9131 18306
rect 9131 18275 9144 18306
rect 9182 18275 9199 18306
rect 9199 18275 9216 18306
rect 9254 18275 9267 18306
rect 9267 18275 9288 18306
rect 9326 18275 9335 18306
rect 9335 18275 9360 18306
rect 9398 18275 9403 18306
rect 9403 18275 9432 18306
rect 9470 18275 9471 18306
rect 9471 18275 9504 18306
rect 9542 18275 9573 18306
rect 9573 18275 9576 18306
rect 9614 18275 9641 18306
rect 9641 18275 9648 18306
rect 9686 18275 9709 18306
rect 9709 18275 9720 18306
rect 9758 18275 9777 18306
rect 9777 18275 9792 18306
rect 9830 18275 9845 18306
rect 9845 18275 9864 18306
rect 9902 18275 9913 18306
rect 9913 18275 9936 18306
rect 9974 18275 9981 18306
rect 9981 18275 10008 18306
rect 10046 18275 10049 18306
rect 10049 18275 10080 18306
rect 10118 18275 10151 18306
rect 10151 18275 10152 18306
rect 10190 18275 10219 18306
rect 10219 18275 10224 18306
rect 10262 18275 10287 18306
rect 10287 18275 10296 18306
rect 10334 18275 10355 18306
rect 10355 18275 10368 18306
rect 10406 18275 10423 18306
rect 10423 18275 10440 18306
rect 10478 18275 10491 18306
rect 10491 18275 10512 18306
rect 10550 18275 10559 18306
rect 10559 18275 10584 18306
rect 10622 18275 10627 18306
rect 10627 18275 10656 18306
rect 10694 18275 10695 18306
rect 10695 18275 10728 18306
rect 10766 18275 10797 18306
rect 10797 18275 10800 18306
rect 10838 18275 10865 18306
rect 10865 18275 10872 18306
rect 10910 18275 10933 18306
rect 10933 18275 10944 18306
rect 10982 18275 11001 18306
rect 11001 18275 11016 18306
rect 11054 18275 11069 18306
rect 11069 18275 11088 18306
rect 11126 18275 11137 18306
rect 11137 18275 11160 18306
rect 11198 18275 11205 18306
rect 11205 18275 11232 18306
rect 11270 18275 11273 18306
rect 11273 18275 11304 18306
rect 11342 18275 11375 18306
rect 11375 18275 11376 18306
rect 11414 18275 11443 18306
rect 11443 18275 11448 18306
rect 11486 18275 11511 18306
rect 11511 18275 11520 18306
rect 11558 18275 11579 18306
rect 11579 18275 11592 18306
rect 11630 18275 11647 18306
rect 11647 18275 11664 18306
rect 11702 18275 11715 18306
rect 11715 18275 11736 18306
rect 11774 18275 11783 18306
rect 11783 18275 11808 18306
rect 11846 18275 11851 18306
rect 11851 18275 11880 18306
rect 11918 18275 11919 18306
rect 11919 18275 11952 18306
rect 11990 18275 12021 18306
rect 12021 18275 12024 18306
rect 12062 18275 12089 18306
rect 12089 18275 12096 18306
rect 12134 18275 12157 18306
rect 12157 18275 12168 18306
rect 12206 18275 12225 18306
rect 12225 18275 12240 18306
rect 12278 18275 12293 18306
rect 12293 18275 12312 18306
rect 12350 18275 12361 18306
rect 12361 18275 12384 18306
rect 12422 18275 12429 18306
rect 12429 18275 12456 18306
rect 12494 18275 12497 18306
rect 12497 18275 12528 18306
rect 12566 18275 12599 18306
rect 12599 18275 12600 18306
rect 12638 18275 12667 18306
rect 12667 18275 12672 18306
rect 12710 18275 12735 18306
rect 12735 18275 12744 18306
rect 12782 18275 12803 18306
rect 12803 18275 12816 18306
rect 12854 18275 12871 18306
rect 12871 18275 12888 18306
rect 12926 18275 12939 18306
rect 12939 18275 12960 18306
rect 12998 18275 13007 18306
rect 13007 18275 13032 18306
rect 13070 18275 13075 18306
rect 13075 18275 13104 18306
rect 13142 18275 13143 18306
rect 13143 18275 13176 18306
rect 13214 18275 13245 18306
rect 13245 18275 13248 18306
rect 13286 18275 13313 18306
rect 13313 18275 13320 18306
rect 13358 18275 13381 18306
rect 13381 18275 13392 18306
rect 13430 18275 13449 18306
rect 13449 18275 13464 18306
rect 13502 18275 13517 18306
rect 13517 18275 13536 18306
rect 13574 18275 13585 18306
rect 13585 18275 13608 18306
rect 13646 18275 13653 18306
rect 13653 18275 13680 18306
rect 13718 18275 13721 18306
rect 13721 18275 13752 18306
rect 13790 18275 13823 18306
rect 13823 18275 13824 18306
rect 13862 18275 13891 18306
rect 13891 18275 13896 18306
rect 13934 18275 13959 18306
rect 13959 18275 13968 18306
rect 14006 18275 14027 18306
rect 14027 18275 14040 18306
rect 14078 18275 14095 18306
rect 14095 18275 14112 18306
rect 14150 18275 14163 18306
rect 14163 18275 14184 18306
rect 14222 18275 14231 18306
rect 14231 18275 14256 18306
rect 14294 18275 14299 18306
rect 14299 18275 14328 18306
rect 14366 18275 14367 18306
rect 14367 18275 14400 18306
rect 14438 18275 14469 18306
rect 14469 18275 14472 18306
rect 14510 18275 14537 18306
rect 14537 18275 14544 18306
rect 14582 18275 14605 18306
rect 14605 18275 14616 18306
rect 14654 18275 14673 18306
rect 14673 18275 14688 18306
rect 14726 18275 14741 18306
rect 14741 18275 14760 18306
rect 209 18272 243 18275
rect 282 18272 316 18275
rect 355 18272 389 18275
rect 428 18272 462 18275
rect 501 18272 535 18275
rect 574 18272 608 18275
rect 647 18272 681 18275
rect 720 18272 754 18275
rect 793 18272 827 18275
rect 866 18272 900 18275
rect 939 18272 973 18275
rect 1012 18272 1046 18275
rect 1085 18272 1119 18275
rect 1158 18272 1192 18275
rect 1231 18272 1265 18275
rect 1304 18272 1338 18275
rect 1377 18272 1411 18275
rect 1450 18272 1484 18275
rect 1523 18272 1557 18275
rect 1596 18272 1630 18275
rect 1669 18272 1703 18275
rect 1742 18272 1776 18275
rect 1815 18272 1849 18275
rect 1888 18272 1922 18275
rect 1961 18272 1995 18275
rect 2034 18272 2068 18275
rect 2107 18272 2141 18275
rect 2180 18272 2214 18275
rect 2253 18272 2287 18275
rect 2326 18272 2360 18275
rect 2399 18272 2433 18275
rect 2472 18272 2506 18275
rect 2545 18272 2579 18275
rect 2618 18272 2652 18275
rect 2691 18272 2725 18275
rect 2764 18272 2798 18275
rect 2837 18272 2871 18275
rect 2910 18272 2944 18275
rect 2983 18272 3017 18275
rect 3056 18272 3090 18275
rect 3129 18272 3163 18275
rect 3202 18272 3236 18275
rect 3275 18272 3309 18275
rect 3348 18272 3382 18275
rect 3421 18272 3455 18275
rect 3494 18272 3528 18275
rect 3566 18272 3600 18275
rect 3638 18272 3672 18275
rect 3710 18272 3744 18275
rect 3782 18272 3816 18275
rect 3854 18272 3888 18275
rect 3926 18272 3960 18275
rect 3998 18272 4032 18275
rect 4070 18272 4104 18275
rect 4142 18272 4176 18275
rect 4214 18272 4248 18275
rect 4286 18272 4320 18275
rect 4358 18272 4392 18275
rect 4430 18272 4464 18275
rect 4502 18272 4536 18275
rect 4574 18272 4608 18275
rect 4646 18272 4680 18275
rect 4718 18272 4752 18275
rect 4790 18272 4824 18275
rect 4862 18272 4896 18275
rect 4934 18272 4968 18275
rect 5006 18272 5040 18275
rect 5078 18272 5112 18275
rect 5150 18272 5184 18275
rect 5222 18272 5256 18275
rect 5294 18272 5328 18275
rect 5366 18272 5400 18275
rect 5438 18272 5472 18275
rect 5510 18272 5544 18275
rect 5582 18272 5616 18275
rect 5654 18272 5688 18275
rect 5726 18272 5760 18275
rect 5798 18272 5832 18275
rect 5870 18272 5904 18275
rect 5942 18272 5976 18275
rect 6014 18272 6048 18275
rect 6086 18272 6120 18275
rect 6158 18272 6192 18275
rect 6230 18272 6264 18275
rect 6302 18272 6336 18275
rect 6374 18272 6408 18275
rect 6446 18272 6480 18275
rect 6518 18272 6552 18275
rect 6590 18272 6624 18275
rect 6662 18272 6696 18275
rect 6734 18272 6768 18275
rect 6806 18272 6840 18275
rect 6878 18272 6912 18275
rect 6950 18272 6984 18275
rect 7022 18272 7056 18275
rect 7094 18272 7128 18275
rect 7166 18272 7200 18275
rect 7238 18272 7272 18275
rect 7310 18272 7344 18275
rect 7382 18272 7416 18275
rect 7454 18272 7488 18275
rect 7526 18272 7560 18275
rect 7598 18272 7632 18275
rect 7670 18272 7704 18275
rect 7742 18272 7776 18275
rect 7814 18272 7848 18275
rect 7886 18272 7920 18275
rect 7958 18272 7992 18275
rect 8030 18272 8064 18275
rect 8102 18272 8136 18275
rect 8174 18272 8208 18275
rect 8246 18272 8280 18275
rect 8318 18272 8352 18275
rect 8390 18272 8424 18275
rect 8462 18272 8496 18275
rect 8534 18272 8568 18275
rect 8606 18272 8640 18275
rect 8678 18272 8712 18275
rect 8750 18272 8784 18275
rect 8822 18272 8856 18275
rect 8894 18272 8928 18275
rect 8966 18272 9000 18275
rect 9038 18272 9072 18275
rect 9110 18272 9144 18275
rect 9182 18272 9216 18275
rect 9254 18272 9288 18275
rect 9326 18272 9360 18275
rect 9398 18272 9432 18275
rect 9470 18272 9504 18275
rect 9542 18272 9576 18275
rect 9614 18272 9648 18275
rect 9686 18272 9720 18275
rect 9758 18272 9792 18275
rect 9830 18272 9864 18275
rect 9902 18272 9936 18275
rect 9974 18272 10008 18275
rect 10046 18272 10080 18275
rect 10118 18272 10152 18275
rect 10190 18272 10224 18275
rect 10262 18272 10296 18275
rect 10334 18272 10368 18275
rect 10406 18272 10440 18275
rect 10478 18272 10512 18275
rect 10550 18272 10584 18275
rect 10622 18272 10656 18275
rect 10694 18272 10728 18275
rect 10766 18272 10800 18275
rect 10838 18272 10872 18275
rect 10910 18272 10944 18275
rect 10982 18272 11016 18275
rect 11054 18272 11088 18275
rect 11126 18272 11160 18275
rect 11198 18272 11232 18275
rect 11270 18272 11304 18275
rect 11342 18272 11376 18275
rect 11414 18272 11448 18275
rect 11486 18272 11520 18275
rect 11558 18272 11592 18275
rect 11630 18272 11664 18275
rect 11702 18272 11736 18275
rect 11774 18272 11808 18275
rect 11846 18272 11880 18275
rect 11918 18272 11952 18275
rect 11990 18272 12024 18275
rect 12062 18272 12096 18275
rect 12134 18272 12168 18275
rect 12206 18272 12240 18275
rect 12278 18272 12312 18275
rect 12350 18272 12384 18275
rect 12422 18272 12456 18275
rect 12494 18272 12528 18275
rect 12566 18272 12600 18275
rect 12638 18272 12672 18275
rect 12710 18272 12744 18275
rect 12782 18272 12816 18275
rect 12854 18272 12888 18275
rect 12926 18272 12960 18275
rect 12998 18272 13032 18275
rect 13070 18272 13104 18275
rect 13142 18272 13176 18275
rect 13214 18272 13248 18275
rect 13286 18272 13320 18275
rect 13358 18272 13392 18275
rect 13430 18272 13464 18275
rect 13502 18272 13536 18275
rect 13574 18272 13608 18275
rect 13646 18272 13680 18275
rect 13718 18272 13752 18275
rect 13790 18272 13824 18275
rect 13862 18272 13896 18275
rect 13934 18272 13968 18275
rect 14006 18272 14040 18275
rect 14078 18272 14112 18275
rect 14150 18272 14184 18275
rect 14222 18272 14256 18275
rect 14294 18272 14328 18275
rect 14366 18272 14400 18275
rect 14438 18272 14472 18275
rect 14510 18272 14544 18275
rect 14582 18272 14616 18275
rect 14654 18272 14688 18275
rect 14726 18272 14760 18275
rect 209 18205 221 18230
rect 221 18205 243 18230
rect 282 18205 290 18230
rect 290 18205 316 18230
rect 355 18205 359 18230
rect 359 18205 389 18230
rect 428 18205 461 18230
rect 461 18205 462 18230
rect 501 18205 529 18230
rect 529 18205 535 18230
rect 574 18205 597 18230
rect 597 18205 608 18230
rect 647 18205 665 18230
rect 665 18205 681 18230
rect 720 18205 733 18230
rect 733 18205 754 18230
rect 793 18205 801 18230
rect 801 18205 827 18230
rect 866 18205 869 18230
rect 869 18205 900 18230
rect 939 18205 971 18230
rect 971 18205 973 18230
rect 1012 18205 1039 18230
rect 1039 18205 1046 18230
rect 1085 18205 1107 18230
rect 1107 18205 1119 18230
rect 1158 18205 1175 18230
rect 1175 18205 1192 18230
rect 1231 18205 1243 18230
rect 1243 18205 1265 18230
rect 1304 18205 1311 18230
rect 1311 18205 1338 18230
rect 1377 18205 1379 18230
rect 1379 18205 1411 18230
rect 1450 18205 1481 18230
rect 1481 18205 1484 18230
rect 1523 18205 1549 18230
rect 1549 18205 1557 18230
rect 1596 18205 1617 18230
rect 1617 18205 1630 18230
rect 1669 18205 1685 18230
rect 1685 18205 1703 18230
rect 1742 18205 1753 18230
rect 1753 18205 1776 18230
rect 1815 18205 1821 18230
rect 1821 18205 1849 18230
rect 1888 18205 1889 18230
rect 1889 18205 1922 18230
rect 1961 18205 1991 18230
rect 1991 18205 1995 18230
rect 2034 18205 2059 18230
rect 2059 18205 2068 18230
rect 2107 18205 2127 18230
rect 2127 18205 2141 18230
rect 2180 18205 2195 18230
rect 2195 18205 2214 18230
rect 2253 18205 2263 18230
rect 2263 18205 2287 18230
rect 2326 18205 2331 18230
rect 2331 18205 2360 18230
rect 2399 18205 2433 18230
rect 2472 18205 2501 18230
rect 2501 18205 2506 18230
rect 2545 18205 2569 18230
rect 2569 18205 2579 18230
rect 2618 18205 2637 18230
rect 2637 18205 2652 18230
rect 2691 18205 2705 18230
rect 2705 18205 2725 18230
rect 2764 18205 2773 18230
rect 2773 18205 2798 18230
rect 2837 18205 2841 18230
rect 2841 18205 2871 18230
rect 2910 18205 2943 18230
rect 2943 18205 2944 18230
rect 2983 18205 3011 18230
rect 3011 18205 3017 18230
rect 3056 18205 3079 18230
rect 3079 18205 3090 18230
rect 3129 18205 3147 18230
rect 3147 18205 3163 18230
rect 3202 18205 3215 18230
rect 3215 18205 3236 18230
rect 3275 18205 3283 18230
rect 3283 18205 3309 18230
rect 3348 18205 3351 18230
rect 3351 18205 3382 18230
rect 3421 18205 3453 18230
rect 3453 18205 3455 18230
rect 3494 18205 3521 18230
rect 3521 18205 3528 18230
rect 3566 18205 3589 18230
rect 3589 18205 3600 18230
rect 3638 18205 3657 18230
rect 3657 18205 3672 18230
rect 3710 18205 3725 18230
rect 3725 18205 3744 18230
rect 3782 18205 3793 18230
rect 3793 18205 3816 18230
rect 3854 18205 3861 18230
rect 3861 18205 3888 18230
rect 3926 18205 3929 18230
rect 3929 18205 3960 18230
rect 3998 18205 4031 18230
rect 4031 18205 4032 18230
rect 4070 18205 4099 18230
rect 4099 18205 4104 18230
rect 4142 18205 4167 18230
rect 4167 18205 4176 18230
rect 4214 18205 4235 18230
rect 4235 18205 4248 18230
rect 4286 18205 4303 18230
rect 4303 18205 4320 18230
rect 4358 18205 4371 18230
rect 4371 18205 4392 18230
rect 4430 18205 4439 18230
rect 4439 18205 4464 18230
rect 4502 18205 4507 18230
rect 4507 18205 4536 18230
rect 4574 18205 4575 18230
rect 4575 18205 4608 18230
rect 4646 18205 4677 18230
rect 4677 18205 4680 18230
rect 4718 18205 4745 18230
rect 4745 18205 4752 18230
rect 4790 18205 4813 18230
rect 4813 18205 4824 18230
rect 4862 18205 4881 18230
rect 4881 18205 4896 18230
rect 4934 18205 4949 18230
rect 4949 18205 4968 18230
rect 5006 18205 5017 18230
rect 5017 18205 5040 18230
rect 5078 18205 5085 18230
rect 5085 18205 5112 18230
rect 5150 18205 5153 18230
rect 5153 18205 5184 18230
rect 5222 18205 5255 18230
rect 5255 18205 5256 18230
rect 5294 18205 5323 18230
rect 5323 18205 5328 18230
rect 5366 18205 5391 18230
rect 5391 18205 5400 18230
rect 5438 18205 5459 18230
rect 5459 18205 5472 18230
rect 5510 18205 5527 18230
rect 5527 18205 5544 18230
rect 5582 18205 5595 18230
rect 5595 18205 5616 18230
rect 5654 18205 5663 18230
rect 5663 18205 5688 18230
rect 5726 18205 5731 18230
rect 5731 18205 5760 18230
rect 5798 18205 5799 18230
rect 5799 18205 5832 18230
rect 5870 18205 5901 18230
rect 5901 18205 5904 18230
rect 5942 18205 5969 18230
rect 5969 18205 5976 18230
rect 6014 18205 6037 18230
rect 6037 18205 6048 18230
rect 6086 18205 6105 18230
rect 6105 18205 6120 18230
rect 6158 18205 6173 18230
rect 6173 18205 6192 18230
rect 6230 18205 6241 18230
rect 6241 18205 6264 18230
rect 6302 18205 6309 18230
rect 6309 18205 6336 18230
rect 6374 18205 6377 18230
rect 6377 18205 6408 18230
rect 6446 18205 6479 18230
rect 6479 18205 6480 18230
rect 6518 18205 6547 18230
rect 6547 18205 6552 18230
rect 6590 18205 6615 18230
rect 6615 18205 6624 18230
rect 6662 18205 6683 18230
rect 6683 18205 6696 18230
rect 6734 18205 6751 18230
rect 6751 18205 6768 18230
rect 6806 18205 6819 18230
rect 6819 18205 6840 18230
rect 6878 18205 6887 18230
rect 6887 18205 6912 18230
rect 6950 18205 6955 18230
rect 6955 18205 6984 18230
rect 7022 18205 7023 18230
rect 7023 18205 7056 18230
rect 7094 18205 7125 18230
rect 7125 18205 7128 18230
rect 7166 18205 7193 18230
rect 7193 18205 7200 18230
rect 7238 18205 7261 18230
rect 7261 18205 7272 18230
rect 7310 18205 7329 18230
rect 7329 18205 7344 18230
rect 7382 18205 7397 18230
rect 7397 18205 7416 18230
rect 7454 18205 7465 18230
rect 7465 18205 7488 18230
rect 7526 18205 7533 18230
rect 7533 18205 7560 18230
rect 7598 18205 7601 18230
rect 7601 18205 7632 18230
rect 7670 18205 7703 18230
rect 7703 18205 7704 18230
rect 7742 18205 7771 18230
rect 7771 18205 7776 18230
rect 7814 18205 7839 18230
rect 7839 18205 7848 18230
rect 7886 18205 7907 18230
rect 7907 18205 7920 18230
rect 7958 18205 7975 18230
rect 7975 18205 7992 18230
rect 8030 18205 8043 18230
rect 8043 18205 8064 18230
rect 8102 18205 8111 18230
rect 8111 18205 8136 18230
rect 8174 18205 8179 18230
rect 8179 18205 8208 18230
rect 8246 18205 8247 18230
rect 8247 18205 8280 18230
rect 8318 18205 8349 18230
rect 8349 18205 8352 18230
rect 8390 18205 8417 18230
rect 8417 18205 8424 18230
rect 8462 18205 8485 18230
rect 8485 18205 8496 18230
rect 8534 18205 8553 18230
rect 8553 18205 8568 18230
rect 8606 18205 8621 18230
rect 8621 18205 8640 18230
rect 8678 18205 8689 18230
rect 8689 18205 8712 18230
rect 8750 18205 8757 18230
rect 8757 18205 8784 18230
rect 8822 18205 8825 18230
rect 8825 18205 8856 18230
rect 8894 18205 8927 18230
rect 8927 18205 8928 18230
rect 8966 18205 8995 18230
rect 8995 18205 9000 18230
rect 9038 18205 9063 18230
rect 9063 18205 9072 18230
rect 9110 18205 9131 18230
rect 9131 18205 9144 18230
rect 9182 18205 9199 18230
rect 9199 18205 9216 18230
rect 9254 18205 9267 18230
rect 9267 18205 9288 18230
rect 9326 18205 9335 18230
rect 9335 18205 9360 18230
rect 9398 18205 9403 18230
rect 9403 18205 9432 18230
rect 9470 18205 9471 18230
rect 9471 18205 9504 18230
rect 9542 18205 9573 18230
rect 9573 18205 9576 18230
rect 9614 18205 9641 18230
rect 9641 18205 9648 18230
rect 9686 18205 9709 18230
rect 9709 18205 9720 18230
rect 9758 18205 9777 18230
rect 9777 18205 9792 18230
rect 9830 18205 9845 18230
rect 9845 18205 9864 18230
rect 9902 18205 9913 18230
rect 9913 18205 9936 18230
rect 9974 18205 9981 18230
rect 9981 18205 10008 18230
rect 10046 18205 10049 18230
rect 10049 18205 10080 18230
rect 10118 18205 10151 18230
rect 10151 18205 10152 18230
rect 10190 18205 10219 18230
rect 10219 18205 10224 18230
rect 10262 18205 10287 18230
rect 10287 18205 10296 18230
rect 10334 18205 10355 18230
rect 10355 18205 10368 18230
rect 10406 18205 10423 18230
rect 10423 18205 10440 18230
rect 10478 18205 10491 18230
rect 10491 18205 10512 18230
rect 10550 18205 10559 18230
rect 10559 18205 10584 18230
rect 10622 18205 10627 18230
rect 10627 18205 10656 18230
rect 10694 18205 10695 18230
rect 10695 18205 10728 18230
rect 10766 18205 10797 18230
rect 10797 18205 10800 18230
rect 10838 18205 10865 18230
rect 10865 18205 10872 18230
rect 10910 18205 10933 18230
rect 10933 18205 10944 18230
rect 10982 18205 11001 18230
rect 11001 18205 11016 18230
rect 11054 18205 11069 18230
rect 11069 18205 11088 18230
rect 11126 18205 11137 18230
rect 11137 18205 11160 18230
rect 11198 18205 11205 18230
rect 11205 18205 11232 18230
rect 11270 18205 11273 18230
rect 11273 18205 11304 18230
rect 11342 18205 11375 18230
rect 11375 18205 11376 18230
rect 11414 18205 11443 18230
rect 11443 18205 11448 18230
rect 11486 18205 11511 18230
rect 11511 18205 11520 18230
rect 11558 18205 11579 18230
rect 11579 18205 11592 18230
rect 11630 18205 11647 18230
rect 11647 18205 11664 18230
rect 11702 18205 11715 18230
rect 11715 18205 11736 18230
rect 11774 18205 11783 18230
rect 11783 18205 11808 18230
rect 11846 18205 11851 18230
rect 11851 18205 11880 18230
rect 11918 18205 11919 18230
rect 11919 18205 11952 18230
rect 11990 18205 12021 18230
rect 12021 18205 12024 18230
rect 12062 18205 12089 18230
rect 12089 18205 12096 18230
rect 12134 18205 12157 18230
rect 12157 18205 12168 18230
rect 12206 18205 12225 18230
rect 12225 18205 12240 18230
rect 12278 18205 12293 18230
rect 12293 18205 12312 18230
rect 12350 18205 12361 18230
rect 12361 18205 12384 18230
rect 12422 18205 12429 18230
rect 12429 18205 12456 18230
rect 12494 18205 12497 18230
rect 12497 18205 12528 18230
rect 12566 18205 12599 18230
rect 12599 18205 12600 18230
rect 12638 18205 12667 18230
rect 12667 18205 12672 18230
rect 12710 18205 12735 18230
rect 12735 18205 12744 18230
rect 12782 18205 12803 18230
rect 12803 18205 12816 18230
rect 12854 18205 12871 18230
rect 12871 18205 12888 18230
rect 12926 18205 12939 18230
rect 12939 18205 12960 18230
rect 12998 18205 13007 18230
rect 13007 18205 13032 18230
rect 13070 18205 13075 18230
rect 13075 18205 13104 18230
rect 13142 18205 13143 18230
rect 13143 18205 13176 18230
rect 13214 18205 13245 18230
rect 13245 18205 13248 18230
rect 13286 18205 13313 18230
rect 13313 18205 13320 18230
rect 13358 18205 13381 18230
rect 13381 18205 13392 18230
rect 13430 18205 13449 18230
rect 13449 18205 13464 18230
rect 13502 18205 13517 18230
rect 13517 18205 13536 18230
rect 13574 18205 13585 18230
rect 13585 18205 13608 18230
rect 13646 18205 13653 18230
rect 13653 18205 13680 18230
rect 13718 18205 13721 18230
rect 13721 18205 13752 18230
rect 13790 18205 13823 18230
rect 13823 18205 13824 18230
rect 13862 18205 13891 18230
rect 13891 18205 13896 18230
rect 13934 18205 13959 18230
rect 13959 18205 13968 18230
rect 14006 18205 14027 18230
rect 14027 18205 14040 18230
rect 14078 18205 14095 18230
rect 14095 18205 14112 18230
rect 14150 18205 14163 18230
rect 14163 18205 14184 18230
rect 14222 18205 14231 18230
rect 14231 18205 14256 18230
rect 14294 18205 14299 18230
rect 14299 18205 14328 18230
rect 14366 18205 14367 18230
rect 14367 18205 14400 18230
rect 14438 18205 14469 18230
rect 14469 18205 14472 18230
rect 14510 18205 14537 18230
rect 14537 18205 14544 18230
rect 14582 18205 14605 18230
rect 14605 18205 14616 18230
rect 14654 18205 14673 18230
rect 14673 18205 14688 18230
rect 14726 18205 14741 18230
rect 14741 18205 14760 18230
rect 209 18196 243 18205
rect 282 18196 316 18205
rect 355 18196 389 18205
rect 428 18196 462 18205
rect 501 18196 535 18205
rect 574 18196 608 18205
rect 647 18196 681 18205
rect 720 18196 754 18205
rect 793 18196 827 18205
rect 866 18196 900 18205
rect 939 18196 973 18205
rect 1012 18196 1046 18205
rect 1085 18196 1119 18205
rect 1158 18196 1192 18205
rect 1231 18196 1265 18205
rect 1304 18196 1338 18205
rect 1377 18196 1411 18205
rect 1450 18196 1484 18205
rect 1523 18196 1557 18205
rect 1596 18196 1630 18205
rect 1669 18196 1703 18205
rect 1742 18196 1776 18205
rect 1815 18196 1849 18205
rect 1888 18196 1922 18205
rect 1961 18196 1995 18205
rect 2034 18196 2068 18205
rect 2107 18196 2141 18205
rect 2180 18196 2214 18205
rect 2253 18196 2287 18205
rect 2326 18196 2360 18205
rect 2399 18196 2433 18205
rect 2472 18196 2506 18205
rect 2545 18196 2579 18205
rect 2618 18196 2652 18205
rect 2691 18196 2725 18205
rect 2764 18196 2798 18205
rect 2837 18196 2871 18205
rect 2910 18196 2944 18205
rect 2983 18196 3017 18205
rect 3056 18196 3090 18205
rect 3129 18196 3163 18205
rect 3202 18196 3236 18205
rect 3275 18196 3309 18205
rect 3348 18196 3382 18205
rect 3421 18196 3455 18205
rect 3494 18196 3528 18205
rect 3566 18196 3600 18205
rect 3638 18196 3672 18205
rect 3710 18196 3744 18205
rect 3782 18196 3816 18205
rect 3854 18196 3888 18205
rect 3926 18196 3960 18205
rect 3998 18196 4032 18205
rect 4070 18196 4104 18205
rect 4142 18196 4176 18205
rect 4214 18196 4248 18205
rect 4286 18196 4320 18205
rect 4358 18196 4392 18205
rect 4430 18196 4464 18205
rect 4502 18196 4536 18205
rect 4574 18196 4608 18205
rect 4646 18196 4680 18205
rect 4718 18196 4752 18205
rect 4790 18196 4824 18205
rect 4862 18196 4896 18205
rect 4934 18196 4968 18205
rect 5006 18196 5040 18205
rect 5078 18196 5112 18205
rect 5150 18196 5184 18205
rect 5222 18196 5256 18205
rect 5294 18196 5328 18205
rect 5366 18196 5400 18205
rect 5438 18196 5472 18205
rect 5510 18196 5544 18205
rect 5582 18196 5616 18205
rect 5654 18196 5688 18205
rect 5726 18196 5760 18205
rect 5798 18196 5832 18205
rect 5870 18196 5904 18205
rect 5942 18196 5976 18205
rect 6014 18196 6048 18205
rect 6086 18196 6120 18205
rect 6158 18196 6192 18205
rect 6230 18196 6264 18205
rect 6302 18196 6336 18205
rect 6374 18196 6408 18205
rect 6446 18196 6480 18205
rect 6518 18196 6552 18205
rect 6590 18196 6624 18205
rect 6662 18196 6696 18205
rect 6734 18196 6768 18205
rect 6806 18196 6840 18205
rect 6878 18196 6912 18205
rect 6950 18196 6984 18205
rect 7022 18196 7056 18205
rect 7094 18196 7128 18205
rect 7166 18196 7200 18205
rect 7238 18196 7272 18205
rect 7310 18196 7344 18205
rect 7382 18196 7416 18205
rect 7454 18196 7488 18205
rect 7526 18196 7560 18205
rect 7598 18196 7632 18205
rect 7670 18196 7704 18205
rect 7742 18196 7776 18205
rect 7814 18196 7848 18205
rect 7886 18196 7920 18205
rect 7958 18196 7992 18205
rect 8030 18196 8064 18205
rect 8102 18196 8136 18205
rect 8174 18196 8208 18205
rect 8246 18196 8280 18205
rect 8318 18196 8352 18205
rect 8390 18196 8424 18205
rect 8462 18196 8496 18205
rect 8534 18196 8568 18205
rect 8606 18196 8640 18205
rect 8678 18196 8712 18205
rect 8750 18196 8784 18205
rect 8822 18196 8856 18205
rect 8894 18196 8928 18205
rect 8966 18196 9000 18205
rect 9038 18196 9072 18205
rect 9110 18196 9144 18205
rect 9182 18196 9216 18205
rect 9254 18196 9288 18205
rect 9326 18196 9360 18205
rect 9398 18196 9432 18205
rect 9470 18196 9504 18205
rect 9542 18196 9576 18205
rect 9614 18196 9648 18205
rect 9686 18196 9720 18205
rect 9758 18196 9792 18205
rect 9830 18196 9864 18205
rect 9902 18196 9936 18205
rect 9974 18196 10008 18205
rect 10046 18196 10080 18205
rect 10118 18196 10152 18205
rect 10190 18196 10224 18205
rect 10262 18196 10296 18205
rect 10334 18196 10368 18205
rect 10406 18196 10440 18205
rect 10478 18196 10512 18205
rect 10550 18196 10584 18205
rect 10622 18196 10656 18205
rect 10694 18196 10728 18205
rect 10766 18196 10800 18205
rect 10838 18196 10872 18205
rect 10910 18196 10944 18205
rect 10982 18196 11016 18205
rect 11054 18196 11088 18205
rect 11126 18196 11160 18205
rect 11198 18196 11232 18205
rect 11270 18196 11304 18205
rect 11342 18196 11376 18205
rect 11414 18196 11448 18205
rect 11486 18196 11520 18205
rect 11558 18196 11592 18205
rect 11630 18196 11664 18205
rect 11702 18196 11736 18205
rect 11774 18196 11808 18205
rect 11846 18196 11880 18205
rect 11918 18196 11952 18205
rect 11990 18196 12024 18205
rect 12062 18196 12096 18205
rect 12134 18196 12168 18205
rect 12206 18196 12240 18205
rect 12278 18196 12312 18205
rect 12350 18196 12384 18205
rect 12422 18196 12456 18205
rect 12494 18196 12528 18205
rect 12566 18196 12600 18205
rect 12638 18196 12672 18205
rect 12710 18196 12744 18205
rect 12782 18196 12816 18205
rect 12854 18196 12888 18205
rect 12926 18196 12960 18205
rect 12998 18196 13032 18205
rect 13070 18196 13104 18205
rect 13142 18196 13176 18205
rect 13214 18196 13248 18205
rect 13286 18196 13320 18205
rect 13358 18196 13392 18205
rect 13430 18196 13464 18205
rect 13502 18196 13536 18205
rect 13574 18196 13608 18205
rect 13646 18196 13680 18205
rect 13718 18196 13752 18205
rect 13790 18196 13824 18205
rect 13862 18196 13896 18205
rect 13934 18196 13968 18205
rect 14006 18196 14040 18205
rect 14078 18196 14112 18205
rect 14150 18196 14184 18205
rect 14222 18196 14256 18205
rect 14294 18196 14328 18205
rect 14366 18196 14400 18205
rect 14438 18196 14472 18205
rect 14510 18196 14544 18205
rect 14582 18196 14616 18205
rect 14654 18196 14688 18205
rect 14726 18196 14760 18205
rect 209 18135 221 18154
rect 221 18135 243 18154
rect 282 18135 290 18154
rect 290 18135 316 18154
rect 355 18135 359 18154
rect 359 18135 389 18154
rect 428 18135 461 18154
rect 461 18135 462 18154
rect 501 18135 529 18154
rect 529 18135 535 18154
rect 574 18135 597 18154
rect 597 18135 608 18154
rect 647 18135 665 18154
rect 665 18135 681 18154
rect 720 18135 733 18154
rect 733 18135 754 18154
rect 793 18135 801 18154
rect 801 18135 827 18154
rect 866 18135 869 18154
rect 869 18135 900 18154
rect 939 18135 971 18154
rect 971 18135 973 18154
rect 1012 18135 1039 18154
rect 1039 18135 1046 18154
rect 1085 18135 1107 18154
rect 1107 18135 1119 18154
rect 1158 18135 1175 18154
rect 1175 18135 1192 18154
rect 1231 18135 1243 18154
rect 1243 18135 1265 18154
rect 1304 18135 1311 18154
rect 1311 18135 1338 18154
rect 1377 18135 1379 18154
rect 1379 18135 1411 18154
rect 1450 18135 1481 18154
rect 1481 18135 1484 18154
rect 1523 18135 1549 18154
rect 1549 18135 1557 18154
rect 1596 18135 1617 18154
rect 1617 18135 1630 18154
rect 1669 18135 1685 18154
rect 1685 18135 1703 18154
rect 1742 18135 1753 18154
rect 1753 18135 1776 18154
rect 1815 18135 1821 18154
rect 1821 18135 1849 18154
rect 1888 18135 1889 18154
rect 1889 18135 1922 18154
rect 1961 18135 1991 18154
rect 1991 18135 1995 18154
rect 2034 18135 2059 18154
rect 2059 18135 2068 18154
rect 2107 18135 2127 18154
rect 2127 18135 2141 18154
rect 2180 18135 2195 18154
rect 2195 18135 2214 18154
rect 2253 18135 2263 18154
rect 2263 18135 2287 18154
rect 2326 18135 2331 18154
rect 2331 18135 2360 18154
rect 2399 18135 2433 18154
rect 2472 18135 2501 18154
rect 2501 18135 2506 18154
rect 2545 18135 2569 18154
rect 2569 18135 2579 18154
rect 2618 18135 2637 18154
rect 2637 18135 2652 18154
rect 2691 18135 2705 18154
rect 2705 18135 2725 18154
rect 2764 18135 2773 18154
rect 2773 18135 2798 18154
rect 2837 18135 2841 18154
rect 2841 18135 2871 18154
rect 2910 18135 2943 18154
rect 2943 18135 2944 18154
rect 2983 18135 3011 18154
rect 3011 18135 3017 18154
rect 3056 18135 3079 18154
rect 3079 18135 3090 18154
rect 3129 18135 3147 18154
rect 3147 18135 3163 18154
rect 3202 18135 3215 18154
rect 3215 18135 3236 18154
rect 3275 18135 3283 18154
rect 3283 18135 3309 18154
rect 3348 18135 3351 18154
rect 3351 18135 3382 18154
rect 3421 18135 3453 18154
rect 3453 18135 3455 18154
rect 3494 18135 3521 18154
rect 3521 18135 3528 18154
rect 3566 18135 3589 18154
rect 3589 18135 3600 18154
rect 3638 18135 3657 18154
rect 3657 18135 3672 18154
rect 3710 18135 3725 18154
rect 3725 18135 3744 18154
rect 3782 18135 3793 18154
rect 3793 18135 3816 18154
rect 3854 18135 3861 18154
rect 3861 18135 3888 18154
rect 3926 18135 3929 18154
rect 3929 18135 3960 18154
rect 3998 18135 4031 18154
rect 4031 18135 4032 18154
rect 4070 18135 4099 18154
rect 4099 18135 4104 18154
rect 4142 18135 4167 18154
rect 4167 18135 4176 18154
rect 4214 18135 4235 18154
rect 4235 18135 4248 18154
rect 4286 18135 4303 18154
rect 4303 18135 4320 18154
rect 4358 18135 4371 18154
rect 4371 18135 4392 18154
rect 4430 18135 4439 18154
rect 4439 18135 4464 18154
rect 4502 18135 4507 18154
rect 4507 18135 4536 18154
rect 4574 18135 4575 18154
rect 4575 18135 4608 18154
rect 4646 18135 4677 18154
rect 4677 18135 4680 18154
rect 4718 18135 4745 18154
rect 4745 18135 4752 18154
rect 4790 18135 4813 18154
rect 4813 18135 4824 18154
rect 4862 18135 4881 18154
rect 4881 18135 4896 18154
rect 4934 18135 4949 18154
rect 4949 18135 4968 18154
rect 5006 18135 5017 18154
rect 5017 18135 5040 18154
rect 5078 18135 5085 18154
rect 5085 18135 5112 18154
rect 5150 18135 5153 18154
rect 5153 18135 5184 18154
rect 5222 18135 5255 18154
rect 5255 18135 5256 18154
rect 5294 18135 5323 18154
rect 5323 18135 5328 18154
rect 5366 18135 5391 18154
rect 5391 18135 5400 18154
rect 5438 18135 5459 18154
rect 5459 18135 5472 18154
rect 5510 18135 5527 18154
rect 5527 18135 5544 18154
rect 5582 18135 5595 18154
rect 5595 18135 5616 18154
rect 5654 18135 5663 18154
rect 5663 18135 5688 18154
rect 5726 18135 5731 18154
rect 5731 18135 5760 18154
rect 5798 18135 5799 18154
rect 5799 18135 5832 18154
rect 5870 18135 5901 18154
rect 5901 18135 5904 18154
rect 5942 18135 5969 18154
rect 5969 18135 5976 18154
rect 6014 18135 6037 18154
rect 6037 18135 6048 18154
rect 6086 18135 6105 18154
rect 6105 18135 6120 18154
rect 6158 18135 6173 18154
rect 6173 18135 6192 18154
rect 6230 18135 6241 18154
rect 6241 18135 6264 18154
rect 6302 18135 6309 18154
rect 6309 18135 6336 18154
rect 6374 18135 6377 18154
rect 6377 18135 6408 18154
rect 6446 18135 6479 18154
rect 6479 18135 6480 18154
rect 6518 18135 6547 18154
rect 6547 18135 6552 18154
rect 6590 18135 6615 18154
rect 6615 18135 6624 18154
rect 6662 18135 6683 18154
rect 6683 18135 6696 18154
rect 6734 18135 6751 18154
rect 6751 18135 6768 18154
rect 6806 18135 6819 18154
rect 6819 18135 6840 18154
rect 6878 18135 6887 18154
rect 6887 18135 6912 18154
rect 6950 18135 6955 18154
rect 6955 18135 6984 18154
rect 7022 18135 7023 18154
rect 7023 18135 7056 18154
rect 7094 18135 7125 18154
rect 7125 18135 7128 18154
rect 7166 18135 7193 18154
rect 7193 18135 7200 18154
rect 7238 18135 7261 18154
rect 7261 18135 7272 18154
rect 7310 18135 7329 18154
rect 7329 18135 7344 18154
rect 7382 18135 7397 18154
rect 7397 18135 7416 18154
rect 7454 18135 7465 18154
rect 7465 18135 7488 18154
rect 7526 18135 7533 18154
rect 7533 18135 7560 18154
rect 7598 18135 7601 18154
rect 7601 18135 7632 18154
rect 7670 18135 7703 18154
rect 7703 18135 7704 18154
rect 7742 18135 7771 18154
rect 7771 18135 7776 18154
rect 7814 18135 7839 18154
rect 7839 18135 7848 18154
rect 7886 18135 7907 18154
rect 7907 18135 7920 18154
rect 7958 18135 7975 18154
rect 7975 18135 7992 18154
rect 8030 18135 8043 18154
rect 8043 18135 8064 18154
rect 8102 18135 8111 18154
rect 8111 18135 8136 18154
rect 8174 18135 8179 18154
rect 8179 18135 8208 18154
rect 8246 18135 8247 18154
rect 8247 18135 8280 18154
rect 8318 18135 8349 18154
rect 8349 18135 8352 18154
rect 8390 18135 8417 18154
rect 8417 18135 8424 18154
rect 8462 18135 8485 18154
rect 8485 18135 8496 18154
rect 8534 18135 8553 18154
rect 8553 18135 8568 18154
rect 8606 18135 8621 18154
rect 8621 18135 8640 18154
rect 8678 18135 8689 18154
rect 8689 18135 8712 18154
rect 8750 18135 8757 18154
rect 8757 18135 8784 18154
rect 8822 18135 8825 18154
rect 8825 18135 8856 18154
rect 8894 18135 8927 18154
rect 8927 18135 8928 18154
rect 8966 18135 8995 18154
rect 8995 18135 9000 18154
rect 9038 18135 9063 18154
rect 9063 18135 9072 18154
rect 9110 18135 9131 18154
rect 9131 18135 9144 18154
rect 9182 18135 9199 18154
rect 9199 18135 9216 18154
rect 9254 18135 9267 18154
rect 9267 18135 9288 18154
rect 9326 18135 9335 18154
rect 9335 18135 9360 18154
rect 9398 18135 9403 18154
rect 9403 18135 9432 18154
rect 9470 18135 9471 18154
rect 9471 18135 9504 18154
rect 9542 18135 9573 18154
rect 9573 18135 9576 18154
rect 9614 18135 9641 18154
rect 9641 18135 9648 18154
rect 9686 18135 9709 18154
rect 9709 18135 9720 18154
rect 9758 18135 9777 18154
rect 9777 18135 9792 18154
rect 9830 18135 9845 18154
rect 9845 18135 9864 18154
rect 9902 18135 9913 18154
rect 9913 18135 9936 18154
rect 9974 18135 9981 18154
rect 9981 18135 10008 18154
rect 10046 18135 10049 18154
rect 10049 18135 10080 18154
rect 10118 18135 10151 18154
rect 10151 18135 10152 18154
rect 10190 18135 10219 18154
rect 10219 18135 10224 18154
rect 10262 18135 10287 18154
rect 10287 18135 10296 18154
rect 10334 18135 10355 18154
rect 10355 18135 10368 18154
rect 10406 18135 10423 18154
rect 10423 18135 10440 18154
rect 10478 18135 10491 18154
rect 10491 18135 10512 18154
rect 10550 18135 10559 18154
rect 10559 18135 10584 18154
rect 10622 18135 10627 18154
rect 10627 18135 10656 18154
rect 10694 18135 10695 18154
rect 10695 18135 10728 18154
rect 10766 18135 10797 18154
rect 10797 18135 10800 18154
rect 10838 18135 10865 18154
rect 10865 18135 10872 18154
rect 10910 18135 10933 18154
rect 10933 18135 10944 18154
rect 10982 18135 11001 18154
rect 11001 18135 11016 18154
rect 11054 18135 11069 18154
rect 11069 18135 11088 18154
rect 11126 18135 11137 18154
rect 11137 18135 11160 18154
rect 11198 18135 11205 18154
rect 11205 18135 11232 18154
rect 11270 18135 11273 18154
rect 11273 18135 11304 18154
rect 11342 18135 11375 18154
rect 11375 18135 11376 18154
rect 11414 18135 11443 18154
rect 11443 18135 11448 18154
rect 11486 18135 11511 18154
rect 11511 18135 11520 18154
rect 11558 18135 11579 18154
rect 11579 18135 11592 18154
rect 11630 18135 11647 18154
rect 11647 18135 11664 18154
rect 11702 18135 11715 18154
rect 11715 18135 11736 18154
rect 11774 18135 11783 18154
rect 11783 18135 11808 18154
rect 11846 18135 11851 18154
rect 11851 18135 11880 18154
rect 11918 18135 11919 18154
rect 11919 18135 11952 18154
rect 11990 18135 12021 18154
rect 12021 18135 12024 18154
rect 12062 18135 12089 18154
rect 12089 18135 12096 18154
rect 12134 18135 12157 18154
rect 12157 18135 12168 18154
rect 12206 18135 12225 18154
rect 12225 18135 12240 18154
rect 12278 18135 12293 18154
rect 12293 18135 12312 18154
rect 12350 18135 12361 18154
rect 12361 18135 12384 18154
rect 12422 18135 12429 18154
rect 12429 18135 12456 18154
rect 12494 18135 12497 18154
rect 12497 18135 12528 18154
rect 12566 18135 12599 18154
rect 12599 18135 12600 18154
rect 12638 18135 12667 18154
rect 12667 18135 12672 18154
rect 12710 18135 12735 18154
rect 12735 18135 12744 18154
rect 12782 18135 12803 18154
rect 12803 18135 12816 18154
rect 12854 18135 12871 18154
rect 12871 18135 12888 18154
rect 12926 18135 12939 18154
rect 12939 18135 12960 18154
rect 12998 18135 13007 18154
rect 13007 18135 13032 18154
rect 13070 18135 13075 18154
rect 13075 18135 13104 18154
rect 13142 18135 13143 18154
rect 13143 18135 13176 18154
rect 13214 18135 13245 18154
rect 13245 18135 13248 18154
rect 13286 18135 13313 18154
rect 13313 18135 13320 18154
rect 13358 18135 13381 18154
rect 13381 18135 13392 18154
rect 13430 18135 13449 18154
rect 13449 18135 13464 18154
rect 13502 18135 13517 18154
rect 13517 18135 13536 18154
rect 13574 18135 13585 18154
rect 13585 18135 13608 18154
rect 13646 18135 13653 18154
rect 13653 18135 13680 18154
rect 13718 18135 13721 18154
rect 13721 18135 13752 18154
rect 13790 18135 13823 18154
rect 13823 18135 13824 18154
rect 13862 18135 13891 18154
rect 13891 18135 13896 18154
rect 13934 18135 13959 18154
rect 13959 18135 13968 18154
rect 14006 18135 14027 18154
rect 14027 18135 14040 18154
rect 14078 18135 14095 18154
rect 14095 18135 14112 18154
rect 14150 18135 14163 18154
rect 14163 18135 14184 18154
rect 14222 18135 14231 18154
rect 14231 18135 14256 18154
rect 14294 18135 14299 18154
rect 14299 18135 14328 18154
rect 14366 18135 14367 18154
rect 14367 18135 14400 18154
rect 14438 18135 14469 18154
rect 14469 18135 14472 18154
rect 14510 18135 14537 18154
rect 14537 18135 14544 18154
rect 14582 18135 14605 18154
rect 14605 18135 14616 18154
rect 14654 18135 14673 18154
rect 14673 18135 14688 18154
rect 14726 18135 14741 18154
rect 14741 18135 14760 18154
rect 209 18120 243 18135
rect 282 18120 316 18135
rect 355 18120 389 18135
rect 428 18120 462 18135
rect 501 18120 535 18135
rect 574 18120 608 18135
rect 647 18120 681 18135
rect 720 18120 754 18135
rect 793 18120 827 18135
rect 866 18120 900 18135
rect 939 18120 973 18135
rect 1012 18120 1046 18135
rect 1085 18120 1119 18135
rect 1158 18120 1192 18135
rect 1231 18120 1265 18135
rect 1304 18120 1338 18135
rect 1377 18120 1411 18135
rect 1450 18120 1484 18135
rect 1523 18120 1557 18135
rect 1596 18120 1630 18135
rect 1669 18120 1703 18135
rect 1742 18120 1776 18135
rect 1815 18120 1849 18135
rect 1888 18120 1922 18135
rect 1961 18120 1995 18135
rect 2034 18120 2068 18135
rect 2107 18120 2141 18135
rect 2180 18120 2214 18135
rect 2253 18120 2287 18135
rect 2326 18120 2360 18135
rect 2399 18120 2433 18135
rect 2472 18120 2506 18135
rect 2545 18120 2579 18135
rect 2618 18120 2652 18135
rect 2691 18120 2725 18135
rect 2764 18120 2798 18135
rect 2837 18120 2871 18135
rect 2910 18120 2944 18135
rect 2983 18120 3017 18135
rect 3056 18120 3090 18135
rect 3129 18120 3163 18135
rect 3202 18120 3236 18135
rect 3275 18120 3309 18135
rect 3348 18120 3382 18135
rect 3421 18120 3455 18135
rect 3494 18120 3528 18135
rect 3566 18120 3600 18135
rect 3638 18120 3672 18135
rect 3710 18120 3744 18135
rect 3782 18120 3816 18135
rect 3854 18120 3888 18135
rect 3926 18120 3960 18135
rect 3998 18120 4032 18135
rect 4070 18120 4104 18135
rect 4142 18120 4176 18135
rect 4214 18120 4248 18135
rect 4286 18120 4320 18135
rect 4358 18120 4392 18135
rect 4430 18120 4464 18135
rect 4502 18120 4536 18135
rect 4574 18120 4608 18135
rect 4646 18120 4680 18135
rect 4718 18120 4752 18135
rect 4790 18120 4824 18135
rect 4862 18120 4896 18135
rect 4934 18120 4968 18135
rect 5006 18120 5040 18135
rect 5078 18120 5112 18135
rect 5150 18120 5184 18135
rect 5222 18120 5256 18135
rect 5294 18120 5328 18135
rect 5366 18120 5400 18135
rect 5438 18120 5472 18135
rect 5510 18120 5544 18135
rect 5582 18120 5616 18135
rect 5654 18120 5688 18135
rect 5726 18120 5760 18135
rect 5798 18120 5832 18135
rect 5870 18120 5904 18135
rect 5942 18120 5976 18135
rect 6014 18120 6048 18135
rect 6086 18120 6120 18135
rect 6158 18120 6192 18135
rect 6230 18120 6264 18135
rect 6302 18120 6336 18135
rect 6374 18120 6408 18135
rect 6446 18120 6480 18135
rect 6518 18120 6552 18135
rect 6590 18120 6624 18135
rect 6662 18120 6696 18135
rect 6734 18120 6768 18135
rect 6806 18120 6840 18135
rect 6878 18120 6912 18135
rect 6950 18120 6984 18135
rect 7022 18120 7056 18135
rect 7094 18120 7128 18135
rect 7166 18120 7200 18135
rect 7238 18120 7272 18135
rect 7310 18120 7344 18135
rect 7382 18120 7416 18135
rect 7454 18120 7488 18135
rect 7526 18120 7560 18135
rect 7598 18120 7632 18135
rect 7670 18120 7704 18135
rect 7742 18120 7776 18135
rect 7814 18120 7848 18135
rect 7886 18120 7920 18135
rect 7958 18120 7992 18135
rect 8030 18120 8064 18135
rect 8102 18120 8136 18135
rect 8174 18120 8208 18135
rect 8246 18120 8280 18135
rect 8318 18120 8352 18135
rect 8390 18120 8424 18135
rect 8462 18120 8496 18135
rect 8534 18120 8568 18135
rect 8606 18120 8640 18135
rect 8678 18120 8712 18135
rect 8750 18120 8784 18135
rect 8822 18120 8856 18135
rect 8894 18120 8928 18135
rect 8966 18120 9000 18135
rect 9038 18120 9072 18135
rect 9110 18120 9144 18135
rect 9182 18120 9216 18135
rect 9254 18120 9288 18135
rect 9326 18120 9360 18135
rect 9398 18120 9432 18135
rect 9470 18120 9504 18135
rect 9542 18120 9576 18135
rect 9614 18120 9648 18135
rect 9686 18120 9720 18135
rect 9758 18120 9792 18135
rect 9830 18120 9864 18135
rect 9902 18120 9936 18135
rect 9974 18120 10008 18135
rect 10046 18120 10080 18135
rect 10118 18120 10152 18135
rect 10190 18120 10224 18135
rect 10262 18120 10296 18135
rect 10334 18120 10368 18135
rect 10406 18120 10440 18135
rect 10478 18120 10512 18135
rect 10550 18120 10584 18135
rect 10622 18120 10656 18135
rect 10694 18120 10728 18135
rect 10766 18120 10800 18135
rect 10838 18120 10872 18135
rect 10910 18120 10944 18135
rect 10982 18120 11016 18135
rect 11054 18120 11088 18135
rect 11126 18120 11160 18135
rect 11198 18120 11232 18135
rect 11270 18120 11304 18135
rect 11342 18120 11376 18135
rect 11414 18120 11448 18135
rect 11486 18120 11520 18135
rect 11558 18120 11592 18135
rect 11630 18120 11664 18135
rect 11702 18120 11736 18135
rect 11774 18120 11808 18135
rect 11846 18120 11880 18135
rect 11918 18120 11952 18135
rect 11990 18120 12024 18135
rect 12062 18120 12096 18135
rect 12134 18120 12168 18135
rect 12206 18120 12240 18135
rect 12278 18120 12312 18135
rect 12350 18120 12384 18135
rect 12422 18120 12456 18135
rect 12494 18120 12528 18135
rect 12566 18120 12600 18135
rect 12638 18120 12672 18135
rect 12710 18120 12744 18135
rect 12782 18120 12816 18135
rect 12854 18120 12888 18135
rect 12926 18120 12960 18135
rect 12998 18120 13032 18135
rect 13070 18120 13104 18135
rect 13142 18120 13176 18135
rect 13214 18120 13248 18135
rect 13286 18120 13320 18135
rect 13358 18120 13392 18135
rect 13430 18120 13464 18135
rect 13502 18120 13536 18135
rect 13574 18120 13608 18135
rect 13646 18120 13680 18135
rect 13718 18120 13752 18135
rect 13790 18120 13824 18135
rect 13862 18120 13896 18135
rect 13934 18120 13968 18135
rect 14006 18120 14040 18135
rect 14078 18120 14112 18135
rect 14150 18120 14184 18135
rect 14222 18120 14256 18135
rect 14294 18120 14328 18135
rect 14366 18120 14400 18135
rect 14438 18120 14472 18135
rect 14510 18120 14544 18135
rect 14582 18120 14616 18135
rect 14654 18120 14688 18135
rect 14726 18120 14760 18135
rect 209 18065 221 18078
rect 221 18065 243 18078
rect 282 18065 290 18078
rect 290 18065 316 18078
rect 355 18065 359 18078
rect 359 18065 389 18078
rect 428 18065 461 18078
rect 461 18065 462 18078
rect 501 18065 529 18078
rect 529 18065 535 18078
rect 574 18065 597 18078
rect 597 18065 608 18078
rect 647 18065 665 18078
rect 665 18065 681 18078
rect 720 18065 733 18078
rect 733 18065 754 18078
rect 793 18065 801 18078
rect 801 18065 827 18078
rect 866 18065 869 18078
rect 869 18065 900 18078
rect 939 18065 971 18078
rect 971 18065 973 18078
rect 1012 18065 1039 18078
rect 1039 18065 1046 18078
rect 1085 18065 1107 18078
rect 1107 18065 1119 18078
rect 1158 18065 1175 18078
rect 1175 18065 1192 18078
rect 1231 18065 1243 18078
rect 1243 18065 1265 18078
rect 1304 18065 1311 18078
rect 1311 18065 1338 18078
rect 1377 18065 1379 18078
rect 1379 18065 1411 18078
rect 1450 18065 1481 18078
rect 1481 18065 1484 18078
rect 1523 18065 1549 18078
rect 1549 18065 1557 18078
rect 1596 18065 1617 18078
rect 1617 18065 1630 18078
rect 1669 18065 1685 18078
rect 1685 18065 1703 18078
rect 1742 18065 1753 18078
rect 1753 18065 1776 18078
rect 1815 18065 1821 18078
rect 1821 18065 1849 18078
rect 1888 18065 1889 18078
rect 1889 18065 1922 18078
rect 1961 18065 1991 18078
rect 1991 18065 1995 18078
rect 2034 18065 2059 18078
rect 2059 18065 2068 18078
rect 2107 18065 2127 18078
rect 2127 18065 2141 18078
rect 2180 18065 2195 18078
rect 2195 18065 2214 18078
rect 2253 18065 2263 18078
rect 2263 18065 2287 18078
rect 2326 18065 2331 18078
rect 2331 18065 2360 18078
rect 2399 18065 2433 18078
rect 2472 18065 2501 18078
rect 2501 18065 2506 18078
rect 2545 18065 2569 18078
rect 2569 18065 2579 18078
rect 2618 18065 2637 18078
rect 2637 18065 2652 18078
rect 2691 18065 2705 18078
rect 2705 18065 2725 18078
rect 2764 18065 2773 18078
rect 2773 18065 2798 18078
rect 2837 18065 2841 18078
rect 2841 18065 2871 18078
rect 2910 18065 2943 18078
rect 2943 18065 2944 18078
rect 2983 18065 3011 18078
rect 3011 18065 3017 18078
rect 3056 18065 3079 18078
rect 3079 18065 3090 18078
rect 3129 18065 3147 18078
rect 3147 18065 3163 18078
rect 3202 18065 3215 18078
rect 3215 18065 3236 18078
rect 3275 18065 3283 18078
rect 3283 18065 3309 18078
rect 3348 18065 3351 18078
rect 3351 18065 3382 18078
rect 3421 18065 3453 18078
rect 3453 18065 3455 18078
rect 3494 18065 3521 18078
rect 3521 18065 3528 18078
rect 3566 18065 3589 18078
rect 3589 18065 3600 18078
rect 3638 18065 3657 18078
rect 3657 18065 3672 18078
rect 3710 18065 3725 18078
rect 3725 18065 3744 18078
rect 3782 18065 3793 18078
rect 3793 18065 3816 18078
rect 3854 18065 3861 18078
rect 3861 18065 3888 18078
rect 3926 18065 3929 18078
rect 3929 18065 3960 18078
rect 3998 18065 4031 18078
rect 4031 18065 4032 18078
rect 4070 18065 4099 18078
rect 4099 18065 4104 18078
rect 4142 18065 4167 18078
rect 4167 18065 4176 18078
rect 4214 18065 4235 18078
rect 4235 18065 4248 18078
rect 4286 18065 4303 18078
rect 4303 18065 4320 18078
rect 4358 18065 4371 18078
rect 4371 18065 4392 18078
rect 4430 18065 4439 18078
rect 4439 18065 4464 18078
rect 4502 18065 4507 18078
rect 4507 18065 4536 18078
rect 4574 18065 4575 18078
rect 4575 18065 4608 18078
rect 4646 18065 4677 18078
rect 4677 18065 4680 18078
rect 4718 18065 4745 18078
rect 4745 18065 4752 18078
rect 4790 18065 4813 18078
rect 4813 18065 4824 18078
rect 4862 18065 4881 18078
rect 4881 18065 4896 18078
rect 4934 18065 4949 18078
rect 4949 18065 4968 18078
rect 5006 18065 5017 18078
rect 5017 18065 5040 18078
rect 5078 18065 5085 18078
rect 5085 18065 5112 18078
rect 5150 18065 5153 18078
rect 5153 18065 5184 18078
rect 5222 18065 5255 18078
rect 5255 18065 5256 18078
rect 5294 18065 5323 18078
rect 5323 18065 5328 18078
rect 5366 18065 5391 18078
rect 5391 18065 5400 18078
rect 5438 18065 5459 18078
rect 5459 18065 5472 18078
rect 5510 18065 5527 18078
rect 5527 18065 5544 18078
rect 5582 18065 5595 18078
rect 5595 18065 5616 18078
rect 5654 18065 5663 18078
rect 5663 18065 5688 18078
rect 5726 18065 5731 18078
rect 5731 18065 5760 18078
rect 5798 18065 5799 18078
rect 5799 18065 5832 18078
rect 5870 18065 5901 18078
rect 5901 18065 5904 18078
rect 5942 18065 5969 18078
rect 5969 18065 5976 18078
rect 6014 18065 6037 18078
rect 6037 18065 6048 18078
rect 6086 18065 6105 18078
rect 6105 18065 6120 18078
rect 6158 18065 6173 18078
rect 6173 18065 6192 18078
rect 6230 18065 6241 18078
rect 6241 18065 6264 18078
rect 6302 18065 6309 18078
rect 6309 18065 6336 18078
rect 6374 18065 6377 18078
rect 6377 18065 6408 18078
rect 6446 18065 6479 18078
rect 6479 18065 6480 18078
rect 6518 18065 6547 18078
rect 6547 18065 6552 18078
rect 6590 18065 6615 18078
rect 6615 18065 6624 18078
rect 6662 18065 6683 18078
rect 6683 18065 6696 18078
rect 6734 18065 6751 18078
rect 6751 18065 6768 18078
rect 6806 18065 6819 18078
rect 6819 18065 6840 18078
rect 6878 18065 6887 18078
rect 6887 18065 6912 18078
rect 6950 18065 6955 18078
rect 6955 18065 6984 18078
rect 7022 18065 7023 18078
rect 7023 18065 7056 18078
rect 7094 18065 7125 18078
rect 7125 18065 7128 18078
rect 7166 18065 7193 18078
rect 7193 18065 7200 18078
rect 7238 18065 7261 18078
rect 7261 18065 7272 18078
rect 7310 18065 7329 18078
rect 7329 18065 7344 18078
rect 7382 18065 7397 18078
rect 7397 18065 7416 18078
rect 7454 18065 7465 18078
rect 7465 18065 7488 18078
rect 7526 18065 7533 18078
rect 7533 18065 7560 18078
rect 7598 18065 7601 18078
rect 7601 18065 7632 18078
rect 7670 18065 7703 18078
rect 7703 18065 7704 18078
rect 7742 18065 7771 18078
rect 7771 18065 7776 18078
rect 7814 18065 7839 18078
rect 7839 18065 7848 18078
rect 7886 18065 7907 18078
rect 7907 18065 7920 18078
rect 7958 18065 7975 18078
rect 7975 18065 7992 18078
rect 8030 18065 8043 18078
rect 8043 18065 8064 18078
rect 8102 18065 8111 18078
rect 8111 18065 8136 18078
rect 8174 18065 8179 18078
rect 8179 18065 8208 18078
rect 8246 18065 8247 18078
rect 8247 18065 8280 18078
rect 8318 18065 8349 18078
rect 8349 18065 8352 18078
rect 8390 18065 8417 18078
rect 8417 18065 8424 18078
rect 8462 18065 8485 18078
rect 8485 18065 8496 18078
rect 8534 18065 8553 18078
rect 8553 18065 8568 18078
rect 8606 18065 8621 18078
rect 8621 18065 8640 18078
rect 8678 18065 8689 18078
rect 8689 18065 8712 18078
rect 8750 18065 8757 18078
rect 8757 18065 8784 18078
rect 8822 18065 8825 18078
rect 8825 18065 8856 18078
rect 8894 18065 8927 18078
rect 8927 18065 8928 18078
rect 8966 18065 8995 18078
rect 8995 18065 9000 18078
rect 9038 18065 9063 18078
rect 9063 18065 9072 18078
rect 9110 18065 9131 18078
rect 9131 18065 9144 18078
rect 9182 18065 9199 18078
rect 9199 18065 9216 18078
rect 9254 18065 9267 18078
rect 9267 18065 9288 18078
rect 9326 18065 9335 18078
rect 9335 18065 9360 18078
rect 9398 18065 9403 18078
rect 9403 18065 9432 18078
rect 9470 18065 9471 18078
rect 9471 18065 9504 18078
rect 9542 18065 9573 18078
rect 9573 18065 9576 18078
rect 9614 18065 9641 18078
rect 9641 18065 9648 18078
rect 9686 18065 9709 18078
rect 9709 18065 9720 18078
rect 9758 18065 9777 18078
rect 9777 18065 9792 18078
rect 9830 18065 9845 18078
rect 9845 18065 9864 18078
rect 9902 18065 9913 18078
rect 9913 18065 9936 18078
rect 9974 18065 9981 18078
rect 9981 18065 10008 18078
rect 10046 18065 10049 18078
rect 10049 18065 10080 18078
rect 10118 18065 10151 18078
rect 10151 18065 10152 18078
rect 10190 18065 10219 18078
rect 10219 18065 10224 18078
rect 10262 18065 10287 18078
rect 10287 18065 10296 18078
rect 10334 18065 10355 18078
rect 10355 18065 10368 18078
rect 10406 18065 10423 18078
rect 10423 18065 10440 18078
rect 10478 18065 10491 18078
rect 10491 18065 10512 18078
rect 10550 18065 10559 18078
rect 10559 18065 10584 18078
rect 10622 18065 10627 18078
rect 10627 18065 10656 18078
rect 10694 18065 10695 18078
rect 10695 18065 10728 18078
rect 10766 18065 10797 18078
rect 10797 18065 10800 18078
rect 10838 18065 10865 18078
rect 10865 18065 10872 18078
rect 10910 18065 10933 18078
rect 10933 18065 10944 18078
rect 10982 18065 11001 18078
rect 11001 18065 11016 18078
rect 11054 18065 11069 18078
rect 11069 18065 11088 18078
rect 11126 18065 11137 18078
rect 11137 18065 11160 18078
rect 11198 18065 11205 18078
rect 11205 18065 11232 18078
rect 11270 18065 11273 18078
rect 11273 18065 11304 18078
rect 11342 18065 11375 18078
rect 11375 18065 11376 18078
rect 11414 18065 11443 18078
rect 11443 18065 11448 18078
rect 11486 18065 11511 18078
rect 11511 18065 11520 18078
rect 11558 18065 11579 18078
rect 11579 18065 11592 18078
rect 11630 18065 11647 18078
rect 11647 18065 11664 18078
rect 11702 18065 11715 18078
rect 11715 18065 11736 18078
rect 11774 18065 11783 18078
rect 11783 18065 11808 18078
rect 11846 18065 11851 18078
rect 11851 18065 11880 18078
rect 11918 18065 11919 18078
rect 11919 18065 11952 18078
rect 11990 18065 12021 18078
rect 12021 18065 12024 18078
rect 12062 18065 12089 18078
rect 12089 18065 12096 18078
rect 12134 18065 12157 18078
rect 12157 18065 12168 18078
rect 12206 18065 12225 18078
rect 12225 18065 12240 18078
rect 12278 18065 12293 18078
rect 12293 18065 12312 18078
rect 12350 18065 12361 18078
rect 12361 18065 12384 18078
rect 12422 18065 12429 18078
rect 12429 18065 12456 18078
rect 12494 18065 12497 18078
rect 12497 18065 12528 18078
rect 12566 18065 12599 18078
rect 12599 18065 12600 18078
rect 12638 18065 12667 18078
rect 12667 18065 12672 18078
rect 12710 18065 12735 18078
rect 12735 18065 12744 18078
rect 12782 18065 12803 18078
rect 12803 18065 12816 18078
rect 12854 18065 12871 18078
rect 12871 18065 12888 18078
rect 12926 18065 12939 18078
rect 12939 18065 12960 18078
rect 12998 18065 13007 18078
rect 13007 18065 13032 18078
rect 13070 18065 13075 18078
rect 13075 18065 13104 18078
rect 13142 18065 13143 18078
rect 13143 18065 13176 18078
rect 13214 18065 13245 18078
rect 13245 18065 13248 18078
rect 13286 18065 13313 18078
rect 13313 18065 13320 18078
rect 13358 18065 13381 18078
rect 13381 18065 13392 18078
rect 13430 18065 13449 18078
rect 13449 18065 13464 18078
rect 13502 18065 13517 18078
rect 13517 18065 13536 18078
rect 13574 18065 13585 18078
rect 13585 18065 13608 18078
rect 13646 18065 13653 18078
rect 13653 18065 13680 18078
rect 13718 18065 13721 18078
rect 13721 18065 13752 18078
rect 13790 18065 13823 18078
rect 13823 18065 13824 18078
rect 13862 18065 13891 18078
rect 13891 18065 13896 18078
rect 13934 18065 13959 18078
rect 13959 18065 13968 18078
rect 14006 18065 14027 18078
rect 14027 18065 14040 18078
rect 14078 18065 14095 18078
rect 14095 18065 14112 18078
rect 14150 18065 14163 18078
rect 14163 18065 14184 18078
rect 14222 18065 14231 18078
rect 14231 18065 14256 18078
rect 14294 18065 14299 18078
rect 14299 18065 14328 18078
rect 14366 18065 14367 18078
rect 14367 18065 14400 18078
rect 14438 18065 14469 18078
rect 14469 18065 14472 18078
rect 14510 18065 14537 18078
rect 14537 18065 14544 18078
rect 14582 18065 14605 18078
rect 14605 18065 14616 18078
rect 14654 18065 14673 18078
rect 14673 18065 14688 18078
rect 14726 18065 14741 18078
rect 14741 18065 14760 18078
rect 209 18044 243 18065
rect 282 18044 316 18065
rect 355 18044 389 18065
rect 428 18044 462 18065
rect 501 18044 535 18065
rect 574 18044 608 18065
rect 647 18044 681 18065
rect 720 18044 754 18065
rect 793 18044 827 18065
rect 866 18044 900 18065
rect 939 18044 973 18065
rect 1012 18044 1046 18065
rect 1085 18044 1119 18065
rect 1158 18044 1192 18065
rect 1231 18044 1265 18065
rect 1304 18044 1338 18065
rect 1377 18044 1411 18065
rect 1450 18044 1484 18065
rect 1523 18044 1557 18065
rect 1596 18044 1630 18065
rect 1669 18044 1703 18065
rect 1742 18044 1776 18065
rect 1815 18044 1849 18065
rect 1888 18044 1922 18065
rect 1961 18044 1995 18065
rect 2034 18044 2068 18065
rect 2107 18044 2141 18065
rect 2180 18044 2214 18065
rect 2253 18044 2287 18065
rect 2326 18044 2360 18065
rect 2399 18044 2433 18065
rect 2472 18044 2506 18065
rect 2545 18044 2579 18065
rect 2618 18044 2652 18065
rect 2691 18044 2725 18065
rect 2764 18044 2798 18065
rect 2837 18044 2871 18065
rect 2910 18044 2944 18065
rect 2983 18044 3017 18065
rect 3056 18044 3090 18065
rect 3129 18044 3163 18065
rect 3202 18044 3236 18065
rect 3275 18044 3309 18065
rect 3348 18044 3382 18065
rect 3421 18044 3455 18065
rect 3494 18044 3528 18065
rect 3566 18044 3600 18065
rect 3638 18044 3672 18065
rect 3710 18044 3744 18065
rect 3782 18044 3816 18065
rect 3854 18044 3888 18065
rect 3926 18044 3960 18065
rect 3998 18044 4032 18065
rect 4070 18044 4104 18065
rect 4142 18044 4176 18065
rect 4214 18044 4248 18065
rect 4286 18044 4320 18065
rect 4358 18044 4392 18065
rect 4430 18044 4464 18065
rect 4502 18044 4536 18065
rect 4574 18044 4608 18065
rect 4646 18044 4680 18065
rect 4718 18044 4752 18065
rect 4790 18044 4824 18065
rect 4862 18044 4896 18065
rect 4934 18044 4968 18065
rect 5006 18044 5040 18065
rect 5078 18044 5112 18065
rect 5150 18044 5184 18065
rect 5222 18044 5256 18065
rect 5294 18044 5328 18065
rect 5366 18044 5400 18065
rect 5438 18044 5472 18065
rect 5510 18044 5544 18065
rect 5582 18044 5616 18065
rect 5654 18044 5688 18065
rect 5726 18044 5760 18065
rect 5798 18044 5832 18065
rect 5870 18044 5904 18065
rect 5942 18044 5976 18065
rect 6014 18044 6048 18065
rect 6086 18044 6120 18065
rect 6158 18044 6192 18065
rect 6230 18044 6264 18065
rect 6302 18044 6336 18065
rect 6374 18044 6408 18065
rect 6446 18044 6480 18065
rect 6518 18044 6552 18065
rect 6590 18044 6624 18065
rect 6662 18044 6696 18065
rect 6734 18044 6768 18065
rect 6806 18044 6840 18065
rect 6878 18044 6912 18065
rect 6950 18044 6984 18065
rect 7022 18044 7056 18065
rect 7094 18044 7128 18065
rect 7166 18044 7200 18065
rect 7238 18044 7272 18065
rect 7310 18044 7344 18065
rect 7382 18044 7416 18065
rect 7454 18044 7488 18065
rect 7526 18044 7560 18065
rect 7598 18044 7632 18065
rect 7670 18044 7704 18065
rect 7742 18044 7776 18065
rect 7814 18044 7848 18065
rect 7886 18044 7920 18065
rect 7958 18044 7992 18065
rect 8030 18044 8064 18065
rect 8102 18044 8136 18065
rect 8174 18044 8208 18065
rect 8246 18044 8280 18065
rect 8318 18044 8352 18065
rect 8390 18044 8424 18065
rect 8462 18044 8496 18065
rect 8534 18044 8568 18065
rect 8606 18044 8640 18065
rect 8678 18044 8712 18065
rect 8750 18044 8784 18065
rect 8822 18044 8856 18065
rect 8894 18044 8928 18065
rect 8966 18044 9000 18065
rect 9038 18044 9072 18065
rect 9110 18044 9144 18065
rect 9182 18044 9216 18065
rect 9254 18044 9288 18065
rect 9326 18044 9360 18065
rect 9398 18044 9432 18065
rect 9470 18044 9504 18065
rect 9542 18044 9576 18065
rect 9614 18044 9648 18065
rect 9686 18044 9720 18065
rect 9758 18044 9792 18065
rect 9830 18044 9864 18065
rect 9902 18044 9936 18065
rect 9974 18044 10008 18065
rect 10046 18044 10080 18065
rect 10118 18044 10152 18065
rect 10190 18044 10224 18065
rect 10262 18044 10296 18065
rect 10334 18044 10368 18065
rect 10406 18044 10440 18065
rect 10478 18044 10512 18065
rect 10550 18044 10584 18065
rect 10622 18044 10656 18065
rect 10694 18044 10728 18065
rect 10766 18044 10800 18065
rect 10838 18044 10872 18065
rect 10910 18044 10944 18065
rect 10982 18044 11016 18065
rect 11054 18044 11088 18065
rect 11126 18044 11160 18065
rect 11198 18044 11232 18065
rect 11270 18044 11304 18065
rect 11342 18044 11376 18065
rect 11414 18044 11448 18065
rect 11486 18044 11520 18065
rect 11558 18044 11592 18065
rect 11630 18044 11664 18065
rect 11702 18044 11736 18065
rect 11774 18044 11808 18065
rect 11846 18044 11880 18065
rect 11918 18044 11952 18065
rect 11990 18044 12024 18065
rect 12062 18044 12096 18065
rect 12134 18044 12168 18065
rect 12206 18044 12240 18065
rect 12278 18044 12312 18065
rect 12350 18044 12384 18065
rect 12422 18044 12456 18065
rect 12494 18044 12528 18065
rect 12566 18044 12600 18065
rect 12638 18044 12672 18065
rect 12710 18044 12744 18065
rect 12782 18044 12816 18065
rect 12854 18044 12888 18065
rect 12926 18044 12960 18065
rect 12998 18044 13032 18065
rect 13070 18044 13104 18065
rect 13142 18044 13176 18065
rect 13214 18044 13248 18065
rect 13286 18044 13320 18065
rect 13358 18044 13392 18065
rect 13430 18044 13464 18065
rect 13502 18044 13536 18065
rect 13574 18044 13608 18065
rect 13646 18044 13680 18065
rect 13718 18044 13752 18065
rect 13790 18044 13824 18065
rect 13862 18044 13896 18065
rect 13934 18044 13968 18065
rect 14006 18044 14040 18065
rect 14078 18044 14112 18065
rect 14150 18044 14184 18065
rect 14222 18044 14256 18065
rect 14294 18044 14328 18065
rect 14366 18044 14400 18065
rect 14438 18044 14472 18065
rect 14510 18044 14544 18065
rect 14582 18044 14616 18065
rect 14654 18044 14688 18065
rect 14726 18044 14760 18065
rect 209 17995 221 18002
rect 221 17995 243 18002
rect 282 17995 290 18002
rect 290 17995 316 18002
rect 355 17995 359 18002
rect 359 17995 389 18002
rect 428 17995 461 18002
rect 461 17995 462 18002
rect 501 17995 529 18002
rect 529 17995 535 18002
rect 574 17995 597 18002
rect 597 17995 608 18002
rect 647 17995 665 18002
rect 665 17995 681 18002
rect 720 17995 733 18002
rect 733 17995 754 18002
rect 793 17995 801 18002
rect 801 17995 827 18002
rect 866 17995 869 18002
rect 869 17995 900 18002
rect 939 17995 971 18002
rect 971 17995 973 18002
rect 1012 17995 1039 18002
rect 1039 17995 1046 18002
rect 1085 17995 1107 18002
rect 1107 17995 1119 18002
rect 1158 17995 1175 18002
rect 1175 17995 1192 18002
rect 1231 17995 1243 18002
rect 1243 17995 1265 18002
rect 1304 17995 1311 18002
rect 1311 17995 1338 18002
rect 1377 17995 1379 18002
rect 1379 17995 1411 18002
rect 1450 17995 1481 18002
rect 1481 17995 1484 18002
rect 1523 17995 1549 18002
rect 1549 17995 1557 18002
rect 1596 17995 1617 18002
rect 1617 17995 1630 18002
rect 1669 17995 1685 18002
rect 1685 17995 1703 18002
rect 1742 17995 1753 18002
rect 1753 17995 1776 18002
rect 1815 17995 1821 18002
rect 1821 17995 1849 18002
rect 1888 17995 1889 18002
rect 1889 17995 1922 18002
rect 1961 17995 1991 18002
rect 1991 17995 1995 18002
rect 2034 17995 2059 18002
rect 2059 17995 2068 18002
rect 2107 17995 2127 18002
rect 2127 17995 2141 18002
rect 2180 17995 2195 18002
rect 2195 17995 2214 18002
rect 2253 17995 2263 18002
rect 2263 17995 2287 18002
rect 2326 17995 2331 18002
rect 2331 17995 2360 18002
rect 2399 17995 2433 18002
rect 2472 17995 2501 18002
rect 2501 17995 2506 18002
rect 2545 17995 2569 18002
rect 2569 17995 2579 18002
rect 2618 17995 2637 18002
rect 2637 17995 2652 18002
rect 2691 17995 2705 18002
rect 2705 17995 2725 18002
rect 2764 17995 2773 18002
rect 2773 17995 2798 18002
rect 2837 17995 2841 18002
rect 2841 17995 2871 18002
rect 2910 17995 2943 18002
rect 2943 17995 2944 18002
rect 2983 17995 3011 18002
rect 3011 17995 3017 18002
rect 3056 17995 3079 18002
rect 3079 17995 3090 18002
rect 3129 17995 3147 18002
rect 3147 17995 3163 18002
rect 3202 17995 3215 18002
rect 3215 17995 3236 18002
rect 3275 17995 3283 18002
rect 3283 17995 3309 18002
rect 3348 17995 3351 18002
rect 3351 17995 3382 18002
rect 3421 17995 3453 18002
rect 3453 17995 3455 18002
rect 3494 17995 3521 18002
rect 3521 17995 3528 18002
rect 3566 17995 3589 18002
rect 3589 17995 3600 18002
rect 3638 17995 3657 18002
rect 3657 17995 3672 18002
rect 3710 17995 3725 18002
rect 3725 17995 3744 18002
rect 3782 17995 3793 18002
rect 3793 17995 3816 18002
rect 3854 17995 3861 18002
rect 3861 17995 3888 18002
rect 3926 17995 3929 18002
rect 3929 17995 3960 18002
rect 3998 17995 4031 18002
rect 4031 17995 4032 18002
rect 4070 17995 4099 18002
rect 4099 17995 4104 18002
rect 4142 17995 4167 18002
rect 4167 17995 4176 18002
rect 4214 17995 4235 18002
rect 4235 17995 4248 18002
rect 4286 17995 4303 18002
rect 4303 17995 4320 18002
rect 4358 17995 4371 18002
rect 4371 17995 4392 18002
rect 4430 17995 4439 18002
rect 4439 17995 4464 18002
rect 4502 17995 4507 18002
rect 4507 17995 4536 18002
rect 4574 17995 4575 18002
rect 4575 17995 4608 18002
rect 4646 17995 4677 18002
rect 4677 17995 4680 18002
rect 4718 17995 4745 18002
rect 4745 17995 4752 18002
rect 4790 17995 4813 18002
rect 4813 17995 4824 18002
rect 4862 17995 4881 18002
rect 4881 17995 4896 18002
rect 4934 17995 4949 18002
rect 4949 17995 4968 18002
rect 5006 17995 5017 18002
rect 5017 17995 5040 18002
rect 5078 17995 5085 18002
rect 5085 17995 5112 18002
rect 5150 17995 5153 18002
rect 5153 17995 5184 18002
rect 5222 17995 5255 18002
rect 5255 17995 5256 18002
rect 5294 17995 5323 18002
rect 5323 17995 5328 18002
rect 5366 17995 5391 18002
rect 5391 17995 5400 18002
rect 5438 17995 5459 18002
rect 5459 17995 5472 18002
rect 5510 17995 5527 18002
rect 5527 17995 5544 18002
rect 5582 17995 5595 18002
rect 5595 17995 5616 18002
rect 5654 17995 5663 18002
rect 5663 17995 5688 18002
rect 5726 17995 5731 18002
rect 5731 17995 5760 18002
rect 5798 17995 5799 18002
rect 5799 17995 5832 18002
rect 5870 17995 5901 18002
rect 5901 17995 5904 18002
rect 5942 17995 5969 18002
rect 5969 17995 5976 18002
rect 6014 17995 6037 18002
rect 6037 17995 6048 18002
rect 6086 17995 6105 18002
rect 6105 17995 6120 18002
rect 6158 17995 6173 18002
rect 6173 17995 6192 18002
rect 6230 17995 6241 18002
rect 6241 17995 6264 18002
rect 6302 17995 6309 18002
rect 6309 17995 6336 18002
rect 6374 17995 6377 18002
rect 6377 17995 6408 18002
rect 6446 17995 6479 18002
rect 6479 17995 6480 18002
rect 6518 17995 6547 18002
rect 6547 17995 6552 18002
rect 6590 17995 6615 18002
rect 6615 17995 6624 18002
rect 6662 17995 6683 18002
rect 6683 17995 6696 18002
rect 6734 17995 6751 18002
rect 6751 17995 6768 18002
rect 6806 17995 6819 18002
rect 6819 17995 6840 18002
rect 6878 17995 6887 18002
rect 6887 17995 6912 18002
rect 6950 17995 6955 18002
rect 6955 17995 6984 18002
rect 7022 17995 7023 18002
rect 7023 17995 7056 18002
rect 7094 17995 7125 18002
rect 7125 17995 7128 18002
rect 7166 17995 7193 18002
rect 7193 17995 7200 18002
rect 7238 17995 7261 18002
rect 7261 17995 7272 18002
rect 7310 17995 7329 18002
rect 7329 17995 7344 18002
rect 7382 17995 7397 18002
rect 7397 17995 7416 18002
rect 7454 17995 7465 18002
rect 7465 17995 7488 18002
rect 7526 17995 7533 18002
rect 7533 17995 7560 18002
rect 7598 17995 7601 18002
rect 7601 17995 7632 18002
rect 7670 17995 7703 18002
rect 7703 17995 7704 18002
rect 7742 17995 7771 18002
rect 7771 17995 7776 18002
rect 7814 17995 7839 18002
rect 7839 17995 7848 18002
rect 7886 17995 7907 18002
rect 7907 17995 7920 18002
rect 7958 17995 7975 18002
rect 7975 17995 7992 18002
rect 8030 17995 8043 18002
rect 8043 17995 8064 18002
rect 8102 17995 8111 18002
rect 8111 17995 8136 18002
rect 8174 17995 8179 18002
rect 8179 17995 8208 18002
rect 8246 17995 8247 18002
rect 8247 17995 8280 18002
rect 8318 17995 8349 18002
rect 8349 17995 8352 18002
rect 8390 17995 8417 18002
rect 8417 17995 8424 18002
rect 8462 17995 8485 18002
rect 8485 17995 8496 18002
rect 8534 17995 8553 18002
rect 8553 17995 8568 18002
rect 8606 17995 8621 18002
rect 8621 17995 8640 18002
rect 8678 17995 8689 18002
rect 8689 17995 8712 18002
rect 8750 17995 8757 18002
rect 8757 17995 8784 18002
rect 8822 17995 8825 18002
rect 8825 17995 8856 18002
rect 8894 17995 8927 18002
rect 8927 17995 8928 18002
rect 8966 17995 8995 18002
rect 8995 17995 9000 18002
rect 9038 17995 9063 18002
rect 9063 17995 9072 18002
rect 9110 17995 9131 18002
rect 9131 17995 9144 18002
rect 9182 17995 9199 18002
rect 9199 17995 9216 18002
rect 9254 17995 9267 18002
rect 9267 17995 9288 18002
rect 9326 17995 9335 18002
rect 9335 17995 9360 18002
rect 9398 17995 9403 18002
rect 9403 17995 9432 18002
rect 9470 17995 9471 18002
rect 9471 17995 9504 18002
rect 9542 17995 9573 18002
rect 9573 17995 9576 18002
rect 9614 17995 9641 18002
rect 9641 17995 9648 18002
rect 9686 17995 9709 18002
rect 9709 17995 9720 18002
rect 9758 17995 9777 18002
rect 9777 17995 9792 18002
rect 9830 17995 9845 18002
rect 9845 17995 9864 18002
rect 9902 17995 9913 18002
rect 9913 17995 9936 18002
rect 9974 17995 9981 18002
rect 9981 17995 10008 18002
rect 10046 17995 10049 18002
rect 10049 17995 10080 18002
rect 10118 17995 10151 18002
rect 10151 17995 10152 18002
rect 10190 17995 10219 18002
rect 10219 17995 10224 18002
rect 10262 17995 10287 18002
rect 10287 17995 10296 18002
rect 10334 17995 10355 18002
rect 10355 17995 10368 18002
rect 10406 17995 10423 18002
rect 10423 17995 10440 18002
rect 10478 17995 10491 18002
rect 10491 17995 10512 18002
rect 10550 17995 10559 18002
rect 10559 17995 10584 18002
rect 10622 17995 10627 18002
rect 10627 17995 10656 18002
rect 10694 17995 10695 18002
rect 10695 17995 10728 18002
rect 10766 17995 10797 18002
rect 10797 17995 10800 18002
rect 10838 17995 10865 18002
rect 10865 17995 10872 18002
rect 10910 17995 10933 18002
rect 10933 17995 10944 18002
rect 10982 17995 11001 18002
rect 11001 17995 11016 18002
rect 11054 17995 11069 18002
rect 11069 17995 11088 18002
rect 11126 17995 11137 18002
rect 11137 17995 11160 18002
rect 11198 17995 11205 18002
rect 11205 17995 11232 18002
rect 11270 17995 11273 18002
rect 11273 17995 11304 18002
rect 11342 17995 11375 18002
rect 11375 17995 11376 18002
rect 11414 17995 11443 18002
rect 11443 17995 11448 18002
rect 11486 17995 11511 18002
rect 11511 17995 11520 18002
rect 11558 17995 11579 18002
rect 11579 17995 11592 18002
rect 11630 17995 11647 18002
rect 11647 17995 11664 18002
rect 11702 17995 11715 18002
rect 11715 17995 11736 18002
rect 11774 17995 11783 18002
rect 11783 17995 11808 18002
rect 11846 17995 11851 18002
rect 11851 17995 11880 18002
rect 11918 17995 11919 18002
rect 11919 17995 11952 18002
rect 11990 17995 12021 18002
rect 12021 17995 12024 18002
rect 12062 17995 12089 18002
rect 12089 17995 12096 18002
rect 12134 17995 12157 18002
rect 12157 17995 12168 18002
rect 12206 17995 12225 18002
rect 12225 17995 12240 18002
rect 12278 17995 12293 18002
rect 12293 17995 12312 18002
rect 12350 17995 12361 18002
rect 12361 17995 12384 18002
rect 12422 17995 12429 18002
rect 12429 17995 12456 18002
rect 12494 17995 12497 18002
rect 12497 17995 12528 18002
rect 12566 17995 12599 18002
rect 12599 17995 12600 18002
rect 12638 17995 12667 18002
rect 12667 17995 12672 18002
rect 12710 17995 12735 18002
rect 12735 17995 12744 18002
rect 12782 17995 12803 18002
rect 12803 17995 12816 18002
rect 12854 17995 12871 18002
rect 12871 17995 12888 18002
rect 12926 17995 12939 18002
rect 12939 17995 12960 18002
rect 12998 17995 13007 18002
rect 13007 17995 13032 18002
rect 13070 17995 13075 18002
rect 13075 17995 13104 18002
rect 13142 17995 13143 18002
rect 13143 17995 13176 18002
rect 13214 17995 13245 18002
rect 13245 17995 13248 18002
rect 13286 17995 13313 18002
rect 13313 17995 13320 18002
rect 13358 17995 13381 18002
rect 13381 17995 13392 18002
rect 13430 17995 13449 18002
rect 13449 17995 13464 18002
rect 13502 17995 13517 18002
rect 13517 17995 13536 18002
rect 13574 17995 13585 18002
rect 13585 17995 13608 18002
rect 13646 17995 13653 18002
rect 13653 17995 13680 18002
rect 13718 17995 13721 18002
rect 13721 17995 13752 18002
rect 13790 17995 13823 18002
rect 13823 17995 13824 18002
rect 13862 17995 13891 18002
rect 13891 17995 13896 18002
rect 13934 17995 13959 18002
rect 13959 17995 13968 18002
rect 14006 17995 14027 18002
rect 14027 17995 14040 18002
rect 14078 17995 14095 18002
rect 14095 17995 14112 18002
rect 14150 17995 14163 18002
rect 14163 17995 14184 18002
rect 14222 17995 14231 18002
rect 14231 17995 14256 18002
rect 14294 17995 14299 18002
rect 14299 17995 14328 18002
rect 14366 17995 14367 18002
rect 14367 17995 14400 18002
rect 14438 17995 14469 18002
rect 14469 17995 14472 18002
rect 14510 17995 14537 18002
rect 14537 17995 14544 18002
rect 14582 17995 14605 18002
rect 14605 17995 14616 18002
rect 14654 17995 14673 18002
rect 14673 17995 14688 18002
rect 14726 17995 14741 18002
rect 14741 17995 14760 18002
rect 209 17968 243 17995
rect 282 17968 316 17995
rect 355 17968 389 17995
rect 428 17968 462 17995
rect 501 17968 535 17995
rect 574 17968 608 17995
rect 647 17968 681 17995
rect 720 17968 754 17995
rect 793 17968 827 17995
rect 866 17968 900 17995
rect 939 17968 973 17995
rect 1012 17968 1046 17995
rect 1085 17968 1119 17995
rect 1158 17968 1192 17995
rect 1231 17968 1265 17995
rect 1304 17968 1338 17995
rect 1377 17968 1411 17995
rect 1450 17968 1484 17995
rect 1523 17968 1557 17995
rect 1596 17968 1630 17995
rect 1669 17968 1703 17995
rect 1742 17968 1776 17995
rect 1815 17968 1849 17995
rect 1888 17968 1922 17995
rect 1961 17968 1995 17995
rect 2034 17968 2068 17995
rect 2107 17968 2141 17995
rect 2180 17968 2214 17995
rect 2253 17968 2287 17995
rect 2326 17968 2360 17995
rect 2399 17968 2433 17995
rect 2472 17968 2506 17995
rect 2545 17968 2579 17995
rect 2618 17968 2652 17995
rect 2691 17968 2725 17995
rect 2764 17968 2798 17995
rect 2837 17968 2871 17995
rect 2910 17968 2944 17995
rect 2983 17968 3017 17995
rect 3056 17968 3090 17995
rect 3129 17968 3163 17995
rect 3202 17968 3236 17995
rect 3275 17968 3309 17995
rect 3348 17968 3382 17995
rect 3421 17968 3455 17995
rect 3494 17968 3528 17995
rect 3566 17968 3600 17995
rect 3638 17968 3672 17995
rect 3710 17968 3744 17995
rect 3782 17968 3816 17995
rect 3854 17968 3888 17995
rect 3926 17968 3960 17995
rect 3998 17968 4032 17995
rect 4070 17968 4104 17995
rect 4142 17968 4176 17995
rect 4214 17968 4248 17995
rect 4286 17968 4320 17995
rect 4358 17968 4392 17995
rect 4430 17968 4464 17995
rect 4502 17968 4536 17995
rect 4574 17968 4608 17995
rect 4646 17968 4680 17995
rect 4718 17968 4752 17995
rect 4790 17968 4824 17995
rect 4862 17968 4896 17995
rect 4934 17968 4968 17995
rect 5006 17968 5040 17995
rect 5078 17968 5112 17995
rect 5150 17968 5184 17995
rect 5222 17968 5256 17995
rect 5294 17968 5328 17995
rect 5366 17968 5400 17995
rect 5438 17968 5472 17995
rect 5510 17968 5544 17995
rect 5582 17968 5616 17995
rect 5654 17968 5688 17995
rect 5726 17968 5760 17995
rect 5798 17968 5832 17995
rect 5870 17968 5904 17995
rect 5942 17968 5976 17995
rect 6014 17968 6048 17995
rect 6086 17968 6120 17995
rect 6158 17968 6192 17995
rect 6230 17968 6264 17995
rect 6302 17968 6336 17995
rect 6374 17968 6408 17995
rect 6446 17968 6480 17995
rect 6518 17968 6552 17995
rect 6590 17968 6624 17995
rect 6662 17968 6696 17995
rect 6734 17968 6768 17995
rect 6806 17968 6840 17995
rect 6878 17968 6912 17995
rect 6950 17968 6984 17995
rect 7022 17968 7056 17995
rect 7094 17968 7128 17995
rect 7166 17968 7200 17995
rect 7238 17968 7272 17995
rect 7310 17968 7344 17995
rect 7382 17968 7416 17995
rect 7454 17968 7488 17995
rect 7526 17968 7560 17995
rect 7598 17968 7632 17995
rect 7670 17968 7704 17995
rect 7742 17968 7776 17995
rect 7814 17968 7848 17995
rect 7886 17968 7920 17995
rect 7958 17968 7992 17995
rect 8030 17968 8064 17995
rect 8102 17968 8136 17995
rect 8174 17968 8208 17995
rect 8246 17968 8280 17995
rect 8318 17968 8352 17995
rect 8390 17968 8424 17995
rect 8462 17968 8496 17995
rect 8534 17968 8568 17995
rect 8606 17968 8640 17995
rect 8678 17968 8712 17995
rect 8750 17968 8784 17995
rect 8822 17968 8856 17995
rect 8894 17968 8928 17995
rect 8966 17968 9000 17995
rect 9038 17968 9072 17995
rect 9110 17968 9144 17995
rect 9182 17968 9216 17995
rect 9254 17968 9288 17995
rect 9326 17968 9360 17995
rect 9398 17968 9432 17995
rect 9470 17968 9504 17995
rect 9542 17968 9576 17995
rect 9614 17968 9648 17995
rect 9686 17968 9720 17995
rect 9758 17968 9792 17995
rect 9830 17968 9864 17995
rect 9902 17968 9936 17995
rect 9974 17968 10008 17995
rect 10046 17968 10080 17995
rect 10118 17968 10152 17995
rect 10190 17968 10224 17995
rect 10262 17968 10296 17995
rect 10334 17968 10368 17995
rect 10406 17968 10440 17995
rect 10478 17968 10512 17995
rect 10550 17968 10584 17995
rect 10622 17968 10656 17995
rect 10694 17968 10728 17995
rect 10766 17968 10800 17995
rect 10838 17968 10872 17995
rect 10910 17968 10944 17995
rect 10982 17968 11016 17995
rect 11054 17968 11088 17995
rect 11126 17968 11160 17995
rect 11198 17968 11232 17995
rect 11270 17968 11304 17995
rect 11342 17968 11376 17995
rect 11414 17968 11448 17995
rect 11486 17968 11520 17995
rect 11558 17968 11592 17995
rect 11630 17968 11664 17995
rect 11702 17968 11736 17995
rect 11774 17968 11808 17995
rect 11846 17968 11880 17995
rect 11918 17968 11952 17995
rect 11990 17968 12024 17995
rect 12062 17968 12096 17995
rect 12134 17968 12168 17995
rect 12206 17968 12240 17995
rect 12278 17968 12312 17995
rect 12350 17968 12384 17995
rect 12422 17968 12456 17995
rect 12494 17968 12528 17995
rect 12566 17968 12600 17995
rect 12638 17968 12672 17995
rect 12710 17968 12744 17995
rect 12782 17968 12816 17995
rect 12854 17968 12888 17995
rect 12926 17968 12960 17995
rect 12998 17968 13032 17995
rect 13070 17968 13104 17995
rect 13142 17968 13176 17995
rect 13214 17968 13248 17995
rect 13286 17968 13320 17995
rect 13358 17968 13392 17995
rect 13430 17968 13464 17995
rect 13502 17968 13536 17995
rect 13574 17968 13608 17995
rect 13646 17968 13680 17995
rect 13718 17968 13752 17995
rect 13790 17968 13824 17995
rect 13862 17968 13896 17995
rect 13934 17968 13968 17995
rect 14006 17968 14040 17995
rect 14078 17968 14112 17995
rect 14150 17968 14184 17995
rect 14222 17968 14256 17995
rect 14294 17968 14328 17995
rect 14366 17968 14400 17995
rect 14438 17968 14472 17995
rect 14510 17968 14544 17995
rect 14582 17968 14616 17995
rect 14654 17968 14688 17995
rect 14726 17968 14760 17995
rect 209 17925 221 17926
rect 221 17925 243 17926
rect 282 17925 290 17926
rect 290 17925 316 17926
rect 355 17925 359 17926
rect 359 17925 389 17926
rect 428 17925 461 17926
rect 461 17925 462 17926
rect 501 17925 529 17926
rect 529 17925 535 17926
rect 574 17925 597 17926
rect 597 17925 608 17926
rect 647 17925 665 17926
rect 665 17925 681 17926
rect 720 17925 733 17926
rect 733 17925 754 17926
rect 793 17925 801 17926
rect 801 17925 827 17926
rect 866 17925 869 17926
rect 869 17925 900 17926
rect 939 17925 971 17926
rect 971 17925 973 17926
rect 1012 17925 1039 17926
rect 1039 17925 1046 17926
rect 1085 17925 1107 17926
rect 1107 17925 1119 17926
rect 1158 17925 1175 17926
rect 1175 17925 1192 17926
rect 1231 17925 1243 17926
rect 1243 17925 1265 17926
rect 1304 17925 1311 17926
rect 1311 17925 1338 17926
rect 1377 17925 1379 17926
rect 1379 17925 1411 17926
rect 1450 17925 1481 17926
rect 1481 17925 1484 17926
rect 1523 17925 1549 17926
rect 1549 17925 1557 17926
rect 1596 17925 1617 17926
rect 1617 17925 1630 17926
rect 1669 17925 1685 17926
rect 1685 17925 1703 17926
rect 1742 17925 1753 17926
rect 1753 17925 1776 17926
rect 1815 17925 1821 17926
rect 1821 17925 1849 17926
rect 1888 17925 1889 17926
rect 1889 17925 1922 17926
rect 1961 17925 1991 17926
rect 1991 17925 1995 17926
rect 2034 17925 2059 17926
rect 2059 17925 2068 17926
rect 2107 17925 2127 17926
rect 2127 17925 2141 17926
rect 2180 17925 2195 17926
rect 2195 17925 2214 17926
rect 2253 17925 2263 17926
rect 2263 17925 2287 17926
rect 2326 17925 2331 17926
rect 2331 17925 2360 17926
rect 2399 17925 2433 17926
rect 2472 17925 2501 17926
rect 2501 17925 2506 17926
rect 2545 17925 2569 17926
rect 2569 17925 2579 17926
rect 2618 17925 2637 17926
rect 2637 17925 2652 17926
rect 2691 17925 2705 17926
rect 2705 17925 2725 17926
rect 2764 17925 2773 17926
rect 2773 17925 2798 17926
rect 2837 17925 2841 17926
rect 2841 17925 2871 17926
rect 2910 17925 2943 17926
rect 2943 17925 2944 17926
rect 2983 17925 3011 17926
rect 3011 17925 3017 17926
rect 3056 17925 3079 17926
rect 3079 17925 3090 17926
rect 3129 17925 3147 17926
rect 3147 17925 3163 17926
rect 3202 17925 3215 17926
rect 3215 17925 3236 17926
rect 3275 17925 3283 17926
rect 3283 17925 3309 17926
rect 3348 17925 3351 17926
rect 3351 17925 3382 17926
rect 3421 17925 3453 17926
rect 3453 17925 3455 17926
rect 3494 17925 3521 17926
rect 3521 17925 3528 17926
rect 3566 17925 3589 17926
rect 3589 17925 3600 17926
rect 3638 17925 3657 17926
rect 3657 17925 3672 17926
rect 3710 17925 3725 17926
rect 3725 17925 3744 17926
rect 3782 17925 3793 17926
rect 3793 17925 3816 17926
rect 3854 17925 3861 17926
rect 3861 17925 3888 17926
rect 3926 17925 3929 17926
rect 3929 17925 3960 17926
rect 3998 17925 4031 17926
rect 4031 17925 4032 17926
rect 4070 17925 4099 17926
rect 4099 17925 4104 17926
rect 4142 17925 4167 17926
rect 4167 17925 4176 17926
rect 4214 17925 4235 17926
rect 4235 17925 4248 17926
rect 4286 17925 4303 17926
rect 4303 17925 4320 17926
rect 4358 17925 4371 17926
rect 4371 17925 4392 17926
rect 4430 17925 4439 17926
rect 4439 17925 4464 17926
rect 4502 17925 4507 17926
rect 4507 17925 4536 17926
rect 4574 17925 4575 17926
rect 4575 17925 4608 17926
rect 4646 17925 4677 17926
rect 4677 17925 4680 17926
rect 4718 17925 4745 17926
rect 4745 17925 4752 17926
rect 4790 17925 4813 17926
rect 4813 17925 4824 17926
rect 4862 17925 4881 17926
rect 4881 17925 4896 17926
rect 4934 17925 4949 17926
rect 4949 17925 4968 17926
rect 5006 17925 5017 17926
rect 5017 17925 5040 17926
rect 5078 17925 5085 17926
rect 5085 17925 5112 17926
rect 5150 17925 5153 17926
rect 5153 17925 5184 17926
rect 5222 17925 5255 17926
rect 5255 17925 5256 17926
rect 5294 17925 5323 17926
rect 5323 17925 5328 17926
rect 5366 17925 5391 17926
rect 5391 17925 5400 17926
rect 5438 17925 5459 17926
rect 5459 17925 5472 17926
rect 5510 17925 5527 17926
rect 5527 17925 5544 17926
rect 5582 17925 5595 17926
rect 5595 17925 5616 17926
rect 5654 17925 5663 17926
rect 5663 17925 5688 17926
rect 5726 17925 5731 17926
rect 5731 17925 5760 17926
rect 5798 17925 5799 17926
rect 5799 17925 5832 17926
rect 5870 17925 5901 17926
rect 5901 17925 5904 17926
rect 5942 17925 5969 17926
rect 5969 17925 5976 17926
rect 6014 17925 6037 17926
rect 6037 17925 6048 17926
rect 6086 17925 6105 17926
rect 6105 17925 6120 17926
rect 6158 17925 6173 17926
rect 6173 17925 6192 17926
rect 6230 17925 6241 17926
rect 6241 17925 6264 17926
rect 6302 17925 6309 17926
rect 6309 17925 6336 17926
rect 6374 17925 6377 17926
rect 6377 17925 6408 17926
rect 6446 17925 6479 17926
rect 6479 17925 6480 17926
rect 6518 17925 6547 17926
rect 6547 17925 6552 17926
rect 6590 17925 6615 17926
rect 6615 17925 6624 17926
rect 6662 17925 6683 17926
rect 6683 17925 6696 17926
rect 6734 17925 6751 17926
rect 6751 17925 6768 17926
rect 6806 17925 6819 17926
rect 6819 17925 6840 17926
rect 6878 17925 6887 17926
rect 6887 17925 6912 17926
rect 6950 17925 6955 17926
rect 6955 17925 6984 17926
rect 7022 17925 7023 17926
rect 7023 17925 7056 17926
rect 7094 17925 7125 17926
rect 7125 17925 7128 17926
rect 7166 17925 7193 17926
rect 7193 17925 7200 17926
rect 7238 17925 7261 17926
rect 7261 17925 7272 17926
rect 7310 17925 7329 17926
rect 7329 17925 7344 17926
rect 7382 17925 7397 17926
rect 7397 17925 7416 17926
rect 7454 17925 7465 17926
rect 7465 17925 7488 17926
rect 7526 17925 7533 17926
rect 7533 17925 7560 17926
rect 7598 17925 7601 17926
rect 7601 17925 7632 17926
rect 7670 17925 7703 17926
rect 7703 17925 7704 17926
rect 7742 17925 7771 17926
rect 7771 17925 7776 17926
rect 7814 17925 7839 17926
rect 7839 17925 7848 17926
rect 7886 17925 7907 17926
rect 7907 17925 7920 17926
rect 7958 17925 7975 17926
rect 7975 17925 7992 17926
rect 8030 17925 8043 17926
rect 8043 17925 8064 17926
rect 8102 17925 8111 17926
rect 8111 17925 8136 17926
rect 8174 17925 8179 17926
rect 8179 17925 8208 17926
rect 8246 17925 8247 17926
rect 8247 17925 8280 17926
rect 8318 17925 8349 17926
rect 8349 17925 8352 17926
rect 8390 17925 8417 17926
rect 8417 17925 8424 17926
rect 8462 17925 8485 17926
rect 8485 17925 8496 17926
rect 8534 17925 8553 17926
rect 8553 17925 8568 17926
rect 8606 17925 8621 17926
rect 8621 17925 8640 17926
rect 8678 17925 8689 17926
rect 8689 17925 8712 17926
rect 8750 17925 8757 17926
rect 8757 17925 8784 17926
rect 8822 17925 8825 17926
rect 8825 17925 8856 17926
rect 8894 17925 8927 17926
rect 8927 17925 8928 17926
rect 8966 17925 8995 17926
rect 8995 17925 9000 17926
rect 9038 17925 9063 17926
rect 9063 17925 9072 17926
rect 9110 17925 9131 17926
rect 9131 17925 9144 17926
rect 9182 17925 9199 17926
rect 9199 17925 9216 17926
rect 9254 17925 9267 17926
rect 9267 17925 9288 17926
rect 9326 17925 9335 17926
rect 9335 17925 9360 17926
rect 9398 17925 9403 17926
rect 9403 17925 9432 17926
rect 9470 17925 9471 17926
rect 9471 17925 9504 17926
rect 9542 17925 9573 17926
rect 9573 17925 9576 17926
rect 9614 17925 9641 17926
rect 9641 17925 9648 17926
rect 9686 17925 9709 17926
rect 9709 17925 9720 17926
rect 9758 17925 9777 17926
rect 9777 17925 9792 17926
rect 9830 17925 9845 17926
rect 9845 17925 9864 17926
rect 9902 17925 9913 17926
rect 9913 17925 9936 17926
rect 9974 17925 9981 17926
rect 9981 17925 10008 17926
rect 10046 17925 10049 17926
rect 10049 17925 10080 17926
rect 10118 17925 10151 17926
rect 10151 17925 10152 17926
rect 10190 17925 10219 17926
rect 10219 17925 10224 17926
rect 10262 17925 10287 17926
rect 10287 17925 10296 17926
rect 10334 17925 10355 17926
rect 10355 17925 10368 17926
rect 10406 17925 10423 17926
rect 10423 17925 10440 17926
rect 10478 17925 10491 17926
rect 10491 17925 10512 17926
rect 10550 17925 10559 17926
rect 10559 17925 10584 17926
rect 10622 17925 10627 17926
rect 10627 17925 10656 17926
rect 10694 17925 10695 17926
rect 10695 17925 10728 17926
rect 10766 17925 10797 17926
rect 10797 17925 10800 17926
rect 10838 17925 10865 17926
rect 10865 17925 10872 17926
rect 10910 17925 10933 17926
rect 10933 17925 10944 17926
rect 10982 17925 11001 17926
rect 11001 17925 11016 17926
rect 11054 17925 11069 17926
rect 11069 17925 11088 17926
rect 11126 17925 11137 17926
rect 11137 17925 11160 17926
rect 11198 17925 11205 17926
rect 11205 17925 11232 17926
rect 11270 17925 11273 17926
rect 11273 17925 11304 17926
rect 11342 17925 11375 17926
rect 11375 17925 11376 17926
rect 11414 17925 11443 17926
rect 11443 17925 11448 17926
rect 11486 17925 11511 17926
rect 11511 17925 11520 17926
rect 11558 17925 11579 17926
rect 11579 17925 11592 17926
rect 11630 17925 11647 17926
rect 11647 17925 11664 17926
rect 11702 17925 11715 17926
rect 11715 17925 11736 17926
rect 11774 17925 11783 17926
rect 11783 17925 11808 17926
rect 11846 17925 11851 17926
rect 11851 17925 11880 17926
rect 11918 17925 11919 17926
rect 11919 17925 11952 17926
rect 11990 17925 12021 17926
rect 12021 17925 12024 17926
rect 12062 17925 12089 17926
rect 12089 17925 12096 17926
rect 12134 17925 12157 17926
rect 12157 17925 12168 17926
rect 12206 17925 12225 17926
rect 12225 17925 12240 17926
rect 12278 17925 12293 17926
rect 12293 17925 12312 17926
rect 12350 17925 12361 17926
rect 12361 17925 12384 17926
rect 12422 17925 12429 17926
rect 12429 17925 12456 17926
rect 12494 17925 12497 17926
rect 12497 17925 12528 17926
rect 12566 17925 12599 17926
rect 12599 17925 12600 17926
rect 12638 17925 12667 17926
rect 12667 17925 12672 17926
rect 12710 17925 12735 17926
rect 12735 17925 12744 17926
rect 12782 17925 12803 17926
rect 12803 17925 12816 17926
rect 12854 17925 12871 17926
rect 12871 17925 12888 17926
rect 12926 17925 12939 17926
rect 12939 17925 12960 17926
rect 12998 17925 13007 17926
rect 13007 17925 13032 17926
rect 13070 17925 13075 17926
rect 13075 17925 13104 17926
rect 13142 17925 13143 17926
rect 13143 17925 13176 17926
rect 13214 17925 13245 17926
rect 13245 17925 13248 17926
rect 13286 17925 13313 17926
rect 13313 17925 13320 17926
rect 13358 17925 13381 17926
rect 13381 17925 13392 17926
rect 13430 17925 13449 17926
rect 13449 17925 13464 17926
rect 13502 17925 13517 17926
rect 13517 17925 13536 17926
rect 13574 17925 13585 17926
rect 13585 17925 13608 17926
rect 13646 17925 13653 17926
rect 13653 17925 13680 17926
rect 13718 17925 13721 17926
rect 13721 17925 13752 17926
rect 13790 17925 13823 17926
rect 13823 17925 13824 17926
rect 13862 17925 13891 17926
rect 13891 17925 13896 17926
rect 13934 17925 13959 17926
rect 13959 17925 13968 17926
rect 14006 17925 14027 17926
rect 14027 17925 14040 17926
rect 14078 17925 14095 17926
rect 14095 17925 14112 17926
rect 14150 17925 14163 17926
rect 14163 17925 14184 17926
rect 14222 17925 14231 17926
rect 14231 17925 14256 17926
rect 14294 17925 14299 17926
rect 14299 17925 14328 17926
rect 14366 17925 14367 17926
rect 14367 17925 14400 17926
rect 14438 17925 14469 17926
rect 14469 17925 14472 17926
rect 14510 17925 14537 17926
rect 14537 17925 14544 17926
rect 14582 17925 14605 17926
rect 14605 17925 14616 17926
rect 14654 17925 14673 17926
rect 14673 17925 14688 17926
rect 14726 17925 14741 17926
rect 14741 17925 14760 17926
rect 209 17892 243 17925
rect 282 17892 316 17925
rect 355 17892 389 17925
rect 428 17892 462 17925
rect 501 17892 535 17925
rect 574 17892 608 17925
rect 647 17892 681 17925
rect 720 17892 754 17925
rect 793 17892 827 17925
rect 866 17892 900 17925
rect 939 17892 973 17925
rect 1012 17892 1046 17925
rect 1085 17892 1119 17925
rect 1158 17892 1192 17925
rect 1231 17892 1265 17925
rect 1304 17892 1338 17925
rect 1377 17892 1411 17925
rect 1450 17892 1484 17925
rect 1523 17892 1557 17925
rect 1596 17892 1630 17925
rect 1669 17892 1703 17925
rect 1742 17892 1776 17925
rect 1815 17892 1849 17925
rect 1888 17892 1922 17925
rect 1961 17892 1995 17925
rect 2034 17892 2068 17925
rect 2107 17892 2141 17925
rect 2180 17892 2214 17925
rect 2253 17892 2287 17925
rect 2326 17892 2360 17925
rect 2399 17892 2433 17925
rect 2472 17892 2506 17925
rect 2545 17892 2579 17925
rect 2618 17892 2652 17925
rect 2691 17892 2725 17925
rect 2764 17892 2798 17925
rect 2837 17892 2871 17925
rect 2910 17892 2944 17925
rect 2983 17892 3017 17925
rect 3056 17892 3090 17925
rect 3129 17892 3163 17925
rect 3202 17892 3236 17925
rect 3275 17892 3309 17925
rect 3348 17892 3382 17925
rect 3421 17892 3455 17925
rect 3494 17892 3528 17925
rect 3566 17892 3600 17925
rect 3638 17892 3672 17925
rect 3710 17892 3744 17925
rect 3782 17892 3816 17925
rect 3854 17892 3888 17925
rect 3926 17892 3960 17925
rect 3998 17892 4032 17925
rect 4070 17892 4104 17925
rect 4142 17892 4176 17925
rect 4214 17892 4248 17925
rect 4286 17892 4320 17925
rect 4358 17892 4392 17925
rect 4430 17892 4464 17925
rect 4502 17892 4536 17925
rect 4574 17892 4608 17925
rect 4646 17892 4680 17925
rect 4718 17892 4752 17925
rect 4790 17892 4824 17925
rect 4862 17892 4896 17925
rect 4934 17892 4968 17925
rect 5006 17892 5040 17925
rect 5078 17892 5112 17925
rect 5150 17892 5184 17925
rect 5222 17892 5256 17925
rect 5294 17892 5328 17925
rect 5366 17892 5400 17925
rect 5438 17892 5472 17925
rect 5510 17892 5544 17925
rect 5582 17892 5616 17925
rect 5654 17892 5688 17925
rect 5726 17892 5760 17925
rect 5798 17892 5832 17925
rect 5870 17892 5904 17925
rect 5942 17892 5976 17925
rect 6014 17892 6048 17925
rect 6086 17892 6120 17925
rect 6158 17892 6192 17925
rect 6230 17892 6264 17925
rect 6302 17892 6336 17925
rect 6374 17892 6408 17925
rect 6446 17892 6480 17925
rect 6518 17892 6552 17925
rect 6590 17892 6624 17925
rect 6662 17892 6696 17925
rect 6734 17892 6768 17925
rect 6806 17892 6840 17925
rect 6878 17892 6912 17925
rect 6950 17892 6984 17925
rect 7022 17892 7056 17925
rect 7094 17892 7128 17925
rect 7166 17892 7200 17925
rect 7238 17892 7272 17925
rect 7310 17892 7344 17925
rect 7382 17892 7416 17925
rect 7454 17892 7488 17925
rect 7526 17892 7560 17925
rect 7598 17892 7632 17925
rect 7670 17892 7704 17925
rect 7742 17892 7776 17925
rect 7814 17892 7848 17925
rect 7886 17892 7920 17925
rect 7958 17892 7992 17925
rect 8030 17892 8064 17925
rect 8102 17892 8136 17925
rect 8174 17892 8208 17925
rect 8246 17892 8280 17925
rect 8318 17892 8352 17925
rect 8390 17892 8424 17925
rect 8462 17892 8496 17925
rect 8534 17892 8568 17925
rect 8606 17892 8640 17925
rect 8678 17892 8712 17925
rect 8750 17892 8784 17925
rect 8822 17892 8856 17925
rect 8894 17892 8928 17925
rect 8966 17892 9000 17925
rect 9038 17892 9072 17925
rect 9110 17892 9144 17925
rect 9182 17892 9216 17925
rect 9254 17892 9288 17925
rect 9326 17892 9360 17925
rect 9398 17892 9432 17925
rect 9470 17892 9504 17925
rect 9542 17892 9576 17925
rect 9614 17892 9648 17925
rect 9686 17892 9720 17925
rect 9758 17892 9792 17925
rect 9830 17892 9864 17925
rect 9902 17892 9936 17925
rect 9974 17892 10008 17925
rect 10046 17892 10080 17925
rect 10118 17892 10152 17925
rect 10190 17892 10224 17925
rect 10262 17892 10296 17925
rect 10334 17892 10368 17925
rect 10406 17892 10440 17925
rect 10478 17892 10512 17925
rect 10550 17892 10584 17925
rect 10622 17892 10656 17925
rect 10694 17892 10728 17925
rect 10766 17892 10800 17925
rect 10838 17892 10872 17925
rect 10910 17892 10944 17925
rect 10982 17892 11016 17925
rect 11054 17892 11088 17925
rect 11126 17892 11160 17925
rect 11198 17892 11232 17925
rect 11270 17892 11304 17925
rect 11342 17892 11376 17925
rect 11414 17892 11448 17925
rect 11486 17892 11520 17925
rect 11558 17892 11592 17925
rect 11630 17892 11664 17925
rect 11702 17892 11736 17925
rect 11774 17892 11808 17925
rect 11846 17892 11880 17925
rect 11918 17892 11952 17925
rect 11990 17892 12024 17925
rect 12062 17892 12096 17925
rect 12134 17892 12168 17925
rect 12206 17892 12240 17925
rect 12278 17892 12312 17925
rect 12350 17892 12384 17925
rect 12422 17892 12456 17925
rect 12494 17892 12528 17925
rect 12566 17892 12600 17925
rect 12638 17892 12672 17925
rect 12710 17892 12744 17925
rect 12782 17892 12816 17925
rect 12854 17892 12888 17925
rect 12926 17892 12960 17925
rect 12998 17892 13032 17925
rect 13070 17892 13104 17925
rect 13142 17892 13176 17925
rect 13214 17892 13248 17925
rect 13286 17892 13320 17925
rect 13358 17892 13392 17925
rect 13430 17892 13464 17925
rect 13502 17892 13536 17925
rect 13574 17892 13608 17925
rect 13646 17892 13680 17925
rect 13718 17892 13752 17925
rect 13790 17892 13824 17925
rect 13862 17892 13896 17925
rect 13934 17892 13968 17925
rect 14006 17892 14040 17925
rect 14078 17892 14112 17925
rect 14150 17892 14184 17925
rect 14222 17892 14256 17925
rect 14294 17892 14328 17925
rect 14366 17892 14400 17925
rect 14438 17892 14472 17925
rect 14510 17892 14544 17925
rect 14582 17892 14616 17925
rect 14654 17892 14688 17925
rect 14726 17892 14760 17925
<< metal1 >>
rect 14279 35712 14285 35764
rect 14337 35712 14349 35764
rect 14401 35712 14407 35764
rect 14279 35632 14285 35684
rect 14337 35632 14349 35684
rect 14401 35632 14407 35684
rect 14279 35552 14285 35604
rect 14337 35552 14349 35604
rect 14401 35552 14407 35604
rect 575 28632 1189 28633
rect 575 28580 581 28632
rect 633 28580 650 28632
rect 702 28580 719 28632
rect 771 28580 788 28632
rect 840 28580 857 28632
rect 909 28580 926 28632
rect 978 28580 995 28632
rect 1047 28580 1063 28632
rect 1115 28580 1131 28632
rect 1183 28580 1189 28632
rect 575 28558 1189 28580
rect 575 28506 581 28558
rect 633 28506 650 28558
rect 702 28506 719 28558
rect 771 28506 788 28558
rect 840 28506 857 28558
rect 909 28506 926 28558
rect 978 28506 995 28558
rect 1047 28506 1063 28558
rect 1115 28506 1131 28558
rect 1183 28506 1189 28558
rect 575 28484 1189 28506
rect 575 28432 581 28484
rect 633 28432 650 28484
rect 702 28432 719 28484
rect 771 28432 788 28484
rect 840 28432 857 28484
rect 909 28432 926 28484
rect 978 28432 995 28484
rect 1047 28432 1063 28484
rect 1115 28432 1131 28484
rect 1183 28432 1189 28484
rect 3472 28581 3478 28633
rect 3530 28581 3546 28633
rect 3598 28581 3614 28633
rect 3666 28581 3682 28633
rect 3734 28581 3750 28633
rect 3802 28581 3818 28633
rect 3870 28581 3886 28633
rect 3938 28581 3954 28633
rect 4006 28581 4021 28633
rect 4073 28581 4088 28633
rect 4140 28581 4155 28633
rect 4207 28581 4222 28633
rect 4274 28581 4289 28633
rect 4341 28581 4356 28633
rect 4408 28581 4423 28633
rect 4475 28581 4490 28633
rect 4542 28581 4557 28633
rect 4609 28581 4615 28633
rect 3472 28559 4615 28581
rect 3472 28507 3478 28559
rect 3530 28507 3546 28559
rect 3598 28507 3614 28559
rect 3666 28507 3682 28559
rect 3734 28507 3750 28559
rect 3802 28507 3818 28559
rect 3870 28507 3886 28559
rect 3938 28507 3954 28559
rect 4006 28507 4021 28559
rect 4073 28507 4088 28559
rect 4140 28507 4155 28559
rect 4207 28507 4222 28559
rect 4274 28507 4289 28559
rect 4341 28507 4356 28559
rect 4408 28507 4423 28559
rect 4475 28507 4490 28559
rect 4542 28507 4557 28559
rect 4609 28507 4615 28559
rect 3472 28485 4615 28507
rect 3472 28433 3478 28485
rect 3530 28433 3546 28485
rect 3598 28433 3614 28485
rect 3666 28433 3682 28485
rect 3734 28433 3750 28485
rect 3802 28433 3818 28485
rect 3870 28433 3886 28485
rect 3938 28433 3954 28485
rect 4006 28433 4021 28485
rect 4073 28433 4088 28485
rect 4140 28433 4155 28485
rect 4207 28433 4222 28485
rect 4274 28433 4289 28485
rect 4341 28433 4356 28485
rect 4408 28433 4423 28485
rect 4475 28433 4490 28485
rect 4542 28433 4557 28485
rect 4609 28433 4615 28485
rect 5455 28581 5461 28633
rect 5513 28581 5528 28633
rect 5580 28581 5595 28633
rect 5647 28581 5662 28633
rect 5714 28581 5729 28633
rect 5781 28581 5796 28633
rect 5848 28581 5863 28633
rect 5915 28581 5930 28633
rect 5982 28581 5997 28633
rect 6049 28581 6064 28633
rect 6116 28581 6132 28633
rect 6184 28581 6200 28633
rect 6252 28581 6268 28633
rect 6320 28581 6336 28633
rect 6388 28581 6404 28633
rect 6456 28581 6472 28633
rect 6524 28581 6540 28633
rect 6592 28581 6598 28633
rect 5455 28559 6598 28581
rect 5455 28507 5461 28559
rect 5513 28507 5528 28559
rect 5580 28507 5595 28559
rect 5647 28507 5662 28559
rect 5714 28507 5729 28559
rect 5781 28507 5796 28559
rect 5848 28507 5863 28559
rect 5915 28507 5930 28559
rect 5982 28507 5997 28559
rect 6049 28507 6064 28559
rect 6116 28507 6132 28559
rect 6184 28507 6200 28559
rect 6252 28507 6268 28559
rect 6320 28507 6336 28559
rect 6388 28507 6404 28559
rect 6456 28507 6472 28559
rect 6524 28507 6540 28559
rect 6592 28507 6598 28559
rect 5455 28485 6598 28507
rect 5455 28433 5461 28485
rect 5513 28433 5528 28485
rect 5580 28433 5595 28485
rect 5647 28433 5662 28485
rect 5714 28433 5729 28485
rect 5781 28433 5796 28485
rect 5848 28433 5863 28485
rect 5915 28433 5930 28485
rect 5982 28433 5997 28485
rect 6049 28433 6064 28485
rect 6116 28433 6132 28485
rect 6184 28433 6200 28485
rect 6252 28433 6268 28485
rect 6320 28433 6336 28485
rect 6388 28433 6404 28485
rect 6456 28433 6472 28485
rect 6524 28433 6540 28485
rect 6592 28433 6598 28485
rect 7439 28581 7445 28633
rect 7497 28581 7512 28633
rect 7564 28581 7579 28633
rect 7631 28581 7646 28633
rect 7698 28581 7713 28633
rect 7765 28581 7780 28633
rect 7832 28581 7847 28633
rect 7899 28581 7914 28633
rect 7966 28581 7981 28633
rect 8033 28581 8048 28633
rect 8100 28581 8116 28633
rect 8168 28581 8184 28633
rect 8236 28581 8252 28633
rect 8304 28581 8320 28633
rect 8372 28581 8388 28633
rect 8440 28581 8456 28633
rect 8508 28581 8524 28633
rect 8576 28581 8582 28633
rect 7439 28559 8582 28581
rect 7439 28507 7445 28559
rect 7497 28507 7512 28559
rect 7564 28507 7579 28559
rect 7631 28507 7646 28559
rect 7698 28507 7713 28559
rect 7765 28507 7780 28559
rect 7832 28507 7847 28559
rect 7899 28507 7914 28559
rect 7966 28507 7981 28559
rect 8033 28507 8048 28559
rect 8100 28507 8116 28559
rect 8168 28507 8184 28559
rect 8236 28507 8252 28559
rect 8304 28507 8320 28559
rect 8372 28507 8388 28559
rect 8440 28507 8456 28559
rect 8508 28507 8524 28559
rect 8576 28507 8582 28559
rect 7439 28485 8582 28507
rect 7439 28433 7445 28485
rect 7497 28433 7512 28485
rect 7564 28433 7579 28485
rect 7631 28433 7646 28485
rect 7698 28433 7713 28485
rect 7765 28433 7780 28485
rect 7832 28433 7847 28485
rect 7899 28433 7914 28485
rect 7966 28433 7981 28485
rect 8033 28433 8048 28485
rect 8100 28433 8116 28485
rect 8168 28433 8184 28485
rect 8236 28433 8252 28485
rect 8304 28433 8320 28485
rect 8372 28433 8388 28485
rect 8440 28433 8456 28485
rect 8508 28433 8524 28485
rect 8576 28433 8582 28485
rect 9423 28581 9429 28633
rect 9481 28581 9517 28633
rect 9569 28581 9575 28633
rect 9423 28559 9575 28581
rect 9423 28507 9429 28559
rect 9481 28507 9517 28559
rect 9569 28507 9575 28559
rect 9423 28485 9575 28507
rect 9423 28433 9429 28485
rect 9481 28433 9517 28485
rect 9569 28433 9575 28485
rect 14281 28627 14639 28633
rect 14281 28575 14282 28627
rect 14334 28575 14358 28627
rect 14410 28575 14434 28627
rect 14486 28575 14510 28627
rect 14562 28575 14586 28627
rect 14638 28575 14639 28627
rect 14281 28562 14639 28575
rect 14281 28510 14282 28562
rect 14334 28510 14358 28562
rect 14410 28510 14434 28562
rect 14486 28510 14510 28562
rect 14562 28510 14586 28562
rect 14638 28510 14639 28562
rect 14281 28497 14639 28510
rect 14281 28445 14282 28497
rect 14334 28445 14358 28497
rect 14410 28445 14434 28497
rect 14486 28445 14510 28497
rect 14562 28445 14586 28497
rect 14638 28445 14639 28497
rect 575 28431 1189 28432
rect 14281 28432 14639 28445
tri 14048 28198 14281 28431 ne
rect 14281 28380 14282 28432
rect 14334 28380 14358 28432
rect 14410 28380 14434 28432
rect 14486 28380 14510 28432
rect 14562 28380 14586 28432
rect 14638 28431 14639 28432
rect 14638 28380 15029 28431
rect 14281 28367 15029 28380
rect 14281 28315 14282 28367
rect 14334 28315 14358 28367
rect 14410 28315 14434 28367
rect 14486 28315 14510 28367
rect 14562 28315 14586 28367
rect 14638 28315 15029 28367
rect 14281 28302 15029 28315
rect 14281 28250 14282 28302
rect 14334 28250 14358 28302
rect 14410 28250 14434 28302
rect 14486 28250 14510 28302
rect 14562 28250 14586 28302
rect 14638 28250 15029 28302
rect 14281 28237 15029 28250
rect 14281 28185 14282 28237
rect 14334 28185 14358 28237
rect 14410 28185 14434 28237
rect 14486 28185 14510 28237
rect 14562 28185 14586 28237
rect 14638 28185 15029 28237
rect 14281 28171 15029 28185
rect 100 28124 13929 28129
rect 100 28122 1303 28124
rect 1355 28122 1371 28124
rect 1423 28122 1439 28124
rect 1491 28122 1507 28124
rect 1559 28122 1575 28124
rect 100 28088 112 28122
rect 146 28088 185 28122
rect 219 28088 258 28122
rect 292 28088 331 28122
rect 365 28088 404 28122
rect 438 28088 477 28122
rect 511 28088 550 28122
rect 584 28088 623 28122
rect 657 28088 696 28122
rect 730 28088 769 28122
rect 803 28088 842 28122
rect 876 28088 915 28122
rect 949 28088 988 28122
rect 1022 28088 1061 28122
rect 1095 28088 1134 28122
rect 1168 28088 1207 28122
rect 1241 28088 1280 28122
rect 1423 28088 1426 28122
rect 1491 28088 1499 28122
rect 1559 28088 1571 28122
rect 100 28072 1303 28088
rect 1355 28072 1371 28088
rect 1423 28072 1439 28088
rect 1491 28072 1507 28088
rect 1559 28072 1575 28088
rect 1627 28072 1643 28124
rect 1695 28072 1711 28124
rect 1763 28072 1779 28124
rect 1831 28072 1847 28124
rect 1899 28072 1914 28124
rect 1966 28072 1981 28124
rect 2033 28122 12157 28124
rect 2037 28088 2075 28122
rect 2109 28088 2147 28122
rect 2181 28088 2219 28122
rect 2253 28088 2291 28122
rect 2325 28088 2363 28122
rect 2397 28088 2435 28122
rect 2469 28088 2507 28122
rect 2541 28088 2579 28122
rect 2613 28088 2651 28122
rect 2685 28088 2723 28122
rect 2757 28088 2795 28122
rect 2829 28088 2867 28122
rect 2901 28088 2939 28122
rect 2973 28088 3011 28122
rect 3045 28088 3083 28122
rect 3117 28088 3155 28122
rect 3189 28088 3227 28122
rect 3261 28088 3299 28122
rect 3333 28088 3371 28122
rect 3405 28088 3443 28122
rect 3477 28088 3515 28122
rect 3549 28088 3587 28122
rect 3621 28088 3659 28122
rect 3693 28088 3731 28122
rect 3765 28088 3803 28122
rect 3837 28088 3875 28122
rect 3909 28088 3947 28122
rect 3981 28088 4019 28122
rect 4053 28088 4091 28122
rect 4125 28088 4163 28122
rect 4197 28088 4235 28122
rect 4269 28088 4307 28122
rect 4341 28088 4379 28122
rect 4413 28088 4451 28122
rect 4485 28088 4523 28122
rect 4557 28088 4595 28122
rect 4629 28088 4667 28122
rect 4701 28088 4739 28122
rect 4773 28088 4811 28122
rect 4845 28088 4883 28122
rect 4917 28088 4955 28122
rect 4989 28088 5027 28122
rect 5061 28088 5099 28122
rect 5133 28088 5171 28122
rect 5205 28088 5243 28122
rect 5277 28088 5315 28122
rect 5349 28088 5387 28122
rect 5421 28088 5459 28122
rect 5493 28088 5531 28122
rect 5565 28088 5603 28122
rect 5637 28088 5675 28122
rect 5709 28088 5747 28122
rect 5781 28088 5819 28122
rect 5853 28088 5891 28122
rect 5925 28088 5963 28122
rect 5997 28088 6035 28122
rect 6069 28088 6107 28122
rect 6141 28088 6179 28122
rect 6213 28088 6251 28122
rect 6285 28088 6323 28122
rect 6357 28088 6395 28122
rect 6429 28088 6467 28122
rect 6501 28088 6539 28122
rect 6573 28088 6611 28122
rect 6645 28088 6683 28122
rect 6717 28088 6755 28122
rect 6789 28088 6827 28122
rect 6861 28088 6899 28122
rect 6933 28088 6971 28122
rect 7005 28088 7043 28122
rect 7077 28088 7115 28122
rect 7149 28088 7187 28122
rect 7221 28088 7259 28122
rect 7293 28088 7331 28122
rect 7365 28088 7403 28122
rect 7437 28088 7475 28122
rect 7509 28088 7547 28122
rect 7581 28088 7619 28122
rect 7653 28088 7691 28122
rect 7725 28088 7763 28122
rect 7797 28088 7835 28122
rect 7869 28088 7907 28122
rect 7941 28088 7979 28122
rect 8013 28088 8051 28122
rect 8085 28088 8123 28122
rect 8157 28088 8195 28122
rect 8229 28088 8267 28122
rect 8301 28088 8339 28122
rect 8373 28088 8411 28122
rect 8445 28088 8483 28122
rect 8517 28088 8555 28122
rect 8589 28088 8627 28122
rect 8661 28088 8699 28122
rect 8733 28088 8771 28122
rect 8805 28088 8843 28122
rect 8877 28088 8915 28122
rect 8949 28088 8987 28122
rect 9021 28088 9059 28122
rect 9093 28088 9131 28122
rect 9165 28088 9203 28122
rect 9237 28088 9275 28122
rect 9309 28088 9347 28122
rect 9381 28088 9419 28122
rect 9453 28088 9491 28122
rect 9525 28088 9563 28122
rect 9597 28088 9635 28122
rect 9669 28088 9707 28122
rect 9741 28088 9779 28122
rect 9813 28088 9851 28122
rect 9885 28088 9923 28122
rect 9957 28088 9995 28122
rect 10029 28088 10067 28122
rect 10101 28088 10139 28122
rect 10173 28088 10211 28122
rect 10245 28088 10283 28122
rect 10317 28088 10355 28122
rect 10389 28088 10427 28122
rect 10461 28088 10499 28122
rect 10533 28088 10571 28122
rect 10605 28088 10643 28122
rect 10677 28088 10715 28122
rect 10749 28088 10787 28122
rect 10821 28088 10859 28122
rect 10893 28088 10931 28122
rect 10965 28088 11003 28122
rect 11037 28088 11075 28122
rect 11109 28088 11147 28122
rect 11181 28088 11219 28122
rect 11253 28088 11291 28122
rect 11325 28088 11363 28122
rect 11397 28088 11435 28122
rect 11469 28088 11507 28122
rect 11541 28088 11579 28122
rect 11613 28088 11651 28122
rect 11685 28088 11723 28122
rect 11757 28088 11795 28122
rect 11829 28088 11867 28122
rect 11901 28088 11939 28122
rect 11973 28088 12011 28122
rect 12045 28088 12083 28122
rect 12117 28088 12155 28122
rect 2033 28072 12157 28088
rect 12209 28072 12225 28124
rect 12277 28072 12293 28124
rect 12345 28072 12361 28124
rect 12413 28072 12429 28124
rect 12481 28072 12497 28124
rect 12549 28072 12565 28124
rect 12617 28122 12633 28124
rect 12685 28122 12701 28124
rect 12753 28122 12768 28124
rect 12820 28122 12835 28124
rect 12887 28122 13929 28124
rect 12621 28088 12633 28122
rect 12693 28088 12701 28122
rect 12765 28088 12768 28122
rect 12909 28088 12947 28122
rect 12981 28088 13019 28122
rect 13053 28088 13091 28122
rect 13125 28088 13163 28122
rect 13197 28088 13235 28122
rect 13269 28088 13307 28122
rect 13341 28088 13379 28122
rect 13413 28088 13451 28122
rect 13485 28088 13523 28122
rect 13557 28088 13595 28122
rect 13629 28088 13667 28122
rect 13701 28088 13739 28122
rect 13773 28088 13811 28122
rect 13845 28088 13883 28122
rect 13917 28088 13929 28122
rect 12617 28072 12633 28088
rect 12685 28072 12701 28088
rect 12753 28072 12768 28088
rect 12820 28072 12835 28088
rect 12887 28072 13929 28088
rect 100 28058 13929 28072
rect 100 28040 1303 28058
rect 1355 28040 1371 28058
rect 1423 28040 1439 28058
rect 1491 28040 1507 28058
rect 1559 28040 1575 28058
rect 100 28006 112 28040
rect 146 28006 185 28040
rect 219 28006 258 28040
rect 292 28006 331 28040
rect 365 28006 404 28040
rect 438 28006 477 28040
rect 511 28006 550 28040
rect 584 28006 623 28040
rect 657 28006 696 28040
rect 730 28006 769 28040
rect 803 28006 842 28040
rect 876 28006 915 28040
rect 949 28006 988 28040
rect 1022 28006 1061 28040
rect 1095 28006 1134 28040
rect 1168 28006 1207 28040
rect 1241 28006 1280 28040
rect 1423 28006 1426 28040
rect 1491 28006 1499 28040
rect 1559 28006 1571 28040
rect 1627 28006 1643 28058
rect 1695 28006 1711 28058
rect 1763 28006 1779 28058
rect 1831 28006 1847 28058
rect 1899 28006 1914 28058
rect 1966 28006 1981 28058
rect 2033 28040 12157 28058
rect 2037 28006 2075 28040
rect 2109 28006 2147 28040
rect 2181 28006 2219 28040
rect 2253 28006 2291 28040
rect 2325 28006 2363 28040
rect 2397 28006 2435 28040
rect 2469 28006 2507 28040
rect 2541 28006 2579 28040
rect 2613 28006 2651 28040
rect 2685 28006 2723 28040
rect 2757 28006 2795 28040
rect 2829 28006 2867 28040
rect 2901 28006 2939 28040
rect 2973 28006 3011 28040
rect 3045 28006 3083 28040
rect 3117 28006 3155 28040
rect 3189 28006 3227 28040
rect 3261 28006 3299 28040
rect 3333 28006 3371 28040
rect 3405 28006 3443 28040
rect 3477 28006 3515 28040
rect 3549 28006 3587 28040
rect 3621 28006 3659 28040
rect 3693 28006 3731 28040
rect 3765 28006 3803 28040
rect 3837 28006 3875 28040
rect 3909 28006 3947 28040
rect 3981 28006 4019 28040
rect 4053 28006 4091 28040
rect 4125 28006 4163 28040
rect 4197 28006 4235 28040
rect 4269 28006 4307 28040
rect 4341 28006 4379 28040
rect 4413 28006 4451 28040
rect 4485 28006 4523 28040
rect 4557 28006 4595 28040
rect 4629 28006 4667 28040
rect 4701 28006 4739 28040
rect 4773 28006 4811 28040
rect 4845 28006 4883 28040
rect 4917 28006 4955 28040
rect 4989 28006 5027 28040
rect 5061 28006 5099 28040
rect 5133 28006 5171 28040
rect 5205 28006 5243 28040
rect 5277 28006 5315 28040
rect 5349 28006 5387 28040
rect 5421 28006 5459 28040
rect 5493 28006 5531 28040
rect 5565 28006 5603 28040
rect 5637 28006 5675 28040
rect 5709 28006 5747 28040
rect 5781 28006 5819 28040
rect 5853 28006 5891 28040
rect 5925 28006 5963 28040
rect 5997 28006 6035 28040
rect 6069 28006 6107 28040
rect 6141 28006 6179 28040
rect 6213 28006 6251 28040
rect 6285 28006 6323 28040
rect 6357 28006 6395 28040
rect 6429 28006 6467 28040
rect 6501 28006 6539 28040
rect 6573 28006 6611 28040
rect 6645 28006 6683 28040
rect 6717 28006 6755 28040
rect 6789 28006 6827 28040
rect 6861 28006 6899 28040
rect 6933 28006 6971 28040
rect 7005 28006 7043 28040
rect 7077 28006 7115 28040
rect 7149 28006 7187 28040
rect 7221 28006 7259 28040
rect 7293 28006 7331 28040
rect 7365 28006 7403 28040
rect 7437 28006 7475 28040
rect 7509 28006 7547 28040
rect 7581 28006 7619 28040
rect 7653 28006 7691 28040
rect 7725 28006 7763 28040
rect 7797 28006 7835 28040
rect 7869 28006 7907 28040
rect 7941 28006 7979 28040
rect 8013 28006 8051 28040
rect 8085 28006 8123 28040
rect 8157 28006 8195 28040
rect 8229 28006 8267 28040
rect 8301 28006 8339 28040
rect 8373 28006 8411 28040
rect 8445 28006 8483 28040
rect 8517 28006 8555 28040
rect 8589 28006 8627 28040
rect 8661 28006 8699 28040
rect 8733 28006 8771 28040
rect 8805 28006 8843 28040
rect 8877 28006 8915 28040
rect 8949 28006 8987 28040
rect 9021 28006 9059 28040
rect 9093 28006 9131 28040
rect 9165 28006 9203 28040
rect 9237 28006 9275 28040
rect 9309 28006 9347 28040
rect 9381 28006 9419 28040
rect 9453 28006 9491 28040
rect 9525 28006 9563 28040
rect 9597 28006 9635 28040
rect 9669 28006 9707 28040
rect 9741 28006 9779 28040
rect 9813 28006 9851 28040
rect 9885 28006 9923 28040
rect 9957 28006 9995 28040
rect 10029 28006 10067 28040
rect 10101 28006 10139 28040
rect 10173 28006 10211 28040
rect 10245 28006 10283 28040
rect 10317 28006 10355 28040
rect 10389 28006 10427 28040
rect 10461 28006 10499 28040
rect 10533 28006 10571 28040
rect 10605 28006 10643 28040
rect 10677 28006 10715 28040
rect 10749 28006 10787 28040
rect 10821 28006 10859 28040
rect 10893 28006 10931 28040
rect 10965 28006 11003 28040
rect 11037 28006 11075 28040
rect 11109 28006 11147 28040
rect 11181 28006 11219 28040
rect 11253 28006 11291 28040
rect 11325 28006 11363 28040
rect 11397 28006 11435 28040
rect 11469 28006 11507 28040
rect 11541 28006 11579 28040
rect 11613 28006 11651 28040
rect 11685 28006 11723 28040
rect 11757 28006 11795 28040
rect 11829 28006 11867 28040
rect 11901 28006 11939 28040
rect 11973 28006 12011 28040
rect 12045 28006 12083 28040
rect 12117 28006 12155 28040
rect 12209 28006 12225 28058
rect 12277 28006 12293 28058
rect 12345 28006 12361 28058
rect 12413 28006 12429 28058
rect 12481 28006 12497 28058
rect 12549 28006 12565 28058
rect 12617 28040 12633 28058
rect 12685 28040 12701 28058
rect 12753 28040 12768 28058
rect 12820 28040 12835 28058
rect 12887 28040 13929 28058
rect 12621 28006 12633 28040
rect 12693 28006 12701 28040
rect 12765 28006 12768 28040
rect 12909 28006 12947 28040
rect 12981 28006 13019 28040
rect 13053 28006 13091 28040
rect 13125 28006 13163 28040
rect 13197 28006 13235 28040
rect 13269 28006 13307 28040
rect 13341 28006 13379 28040
rect 13413 28006 13451 28040
rect 13485 28006 13523 28040
rect 13557 28006 13595 28040
rect 13629 28006 13667 28040
rect 13701 28006 13739 28040
rect 13773 28006 13811 28040
rect 13845 28006 13883 28040
rect 13917 28006 13929 28040
rect 100 27992 13929 28006
rect 100 27958 1303 27992
rect 1355 27958 1371 27992
rect 1423 27958 1439 27992
rect 1491 27958 1507 27992
rect 1559 27958 1575 27992
rect 100 27924 112 27958
rect 146 27924 185 27958
rect 219 27924 258 27958
rect 292 27924 331 27958
rect 365 27924 404 27958
rect 438 27924 477 27958
rect 511 27924 550 27958
rect 584 27924 623 27958
rect 657 27924 696 27958
rect 730 27924 769 27958
rect 803 27924 842 27958
rect 876 27924 915 27958
rect 949 27924 988 27958
rect 1022 27924 1061 27958
rect 1095 27924 1134 27958
rect 1168 27924 1207 27958
rect 1241 27924 1280 27958
rect 1423 27940 1426 27958
rect 1491 27940 1499 27958
rect 1559 27940 1571 27958
rect 1627 27940 1643 27992
rect 1695 27940 1711 27992
rect 1763 27940 1779 27992
rect 1831 27940 1847 27992
rect 1899 27940 1914 27992
rect 1966 27940 1981 27992
rect 2033 27958 12157 27992
rect 1314 27926 1353 27940
rect 1387 27926 1426 27940
rect 1460 27926 1499 27940
rect 1533 27926 1571 27940
rect 1605 27926 1643 27940
rect 1677 27926 1715 27940
rect 1749 27926 1787 27940
rect 1821 27926 1859 27940
rect 1893 27926 1931 27940
rect 1965 27926 2003 27940
rect 1423 27924 1426 27926
rect 1491 27924 1499 27926
rect 1559 27924 1571 27926
rect 100 27876 1303 27924
rect 1355 27876 1371 27924
rect 1423 27876 1439 27924
rect 1491 27876 1507 27924
rect 1559 27876 1575 27924
rect 100 27842 112 27876
rect 146 27842 185 27876
rect 219 27842 258 27876
rect 292 27842 331 27876
rect 365 27842 404 27876
rect 438 27842 477 27876
rect 511 27842 550 27876
rect 584 27842 623 27876
rect 657 27842 696 27876
rect 730 27842 769 27876
rect 803 27842 842 27876
rect 876 27842 915 27876
rect 949 27842 988 27876
rect 1022 27842 1061 27876
rect 1095 27842 1134 27876
rect 1168 27842 1207 27876
rect 1241 27842 1280 27876
rect 1423 27874 1426 27876
rect 1491 27874 1499 27876
rect 1559 27874 1571 27876
rect 1627 27874 1643 27926
rect 1695 27874 1711 27926
rect 1763 27874 1779 27926
rect 1831 27874 1847 27926
rect 1899 27874 1914 27926
rect 1966 27874 1981 27926
rect 2037 27924 2075 27958
rect 2109 27924 2147 27958
rect 2181 27924 2219 27958
rect 2253 27924 2291 27958
rect 2325 27924 2363 27958
rect 2397 27924 2435 27958
rect 2469 27924 2507 27958
rect 2541 27924 2579 27958
rect 2613 27924 2651 27958
rect 2685 27924 2723 27958
rect 2757 27924 2795 27958
rect 2829 27924 2867 27958
rect 2901 27924 2939 27958
rect 2973 27924 3011 27958
rect 3045 27924 3083 27958
rect 3117 27924 3155 27958
rect 3189 27924 3227 27958
rect 3261 27924 3299 27958
rect 3333 27924 3371 27958
rect 3405 27924 3443 27958
rect 3477 27924 3515 27958
rect 3549 27924 3587 27958
rect 3621 27924 3659 27958
rect 3693 27924 3731 27958
rect 3765 27924 3803 27958
rect 3837 27924 3875 27958
rect 3909 27924 3947 27958
rect 3981 27924 4019 27958
rect 4053 27924 4091 27958
rect 4125 27924 4163 27958
rect 4197 27924 4235 27958
rect 4269 27924 4307 27958
rect 4341 27924 4379 27958
rect 4413 27924 4451 27958
rect 4485 27924 4523 27958
rect 4557 27924 4595 27958
rect 4629 27924 4667 27958
rect 4701 27924 4739 27958
rect 4773 27924 4811 27958
rect 4845 27924 4883 27958
rect 4917 27924 4955 27958
rect 4989 27924 5027 27958
rect 5061 27924 5099 27958
rect 5133 27924 5171 27958
rect 5205 27924 5243 27958
rect 5277 27924 5315 27958
rect 5349 27924 5387 27958
rect 5421 27924 5459 27958
rect 5493 27924 5531 27958
rect 5565 27924 5603 27958
rect 5637 27924 5675 27958
rect 5709 27924 5747 27958
rect 5781 27924 5819 27958
rect 5853 27924 5891 27958
rect 5925 27924 5963 27958
rect 5997 27924 6035 27958
rect 6069 27924 6107 27958
rect 6141 27924 6179 27958
rect 6213 27924 6251 27958
rect 6285 27924 6323 27958
rect 6357 27924 6395 27958
rect 6429 27924 6467 27958
rect 6501 27924 6539 27958
rect 6573 27924 6611 27958
rect 6645 27924 6683 27958
rect 6717 27924 6755 27958
rect 6789 27924 6827 27958
rect 6861 27924 6899 27958
rect 6933 27924 6971 27958
rect 7005 27924 7043 27958
rect 7077 27924 7115 27958
rect 7149 27924 7187 27958
rect 7221 27924 7259 27958
rect 7293 27924 7331 27958
rect 7365 27924 7403 27958
rect 7437 27924 7475 27958
rect 7509 27924 7547 27958
rect 7581 27924 7619 27958
rect 7653 27924 7691 27958
rect 7725 27924 7763 27958
rect 7797 27924 7835 27958
rect 7869 27924 7907 27958
rect 7941 27924 7979 27958
rect 8013 27924 8051 27958
rect 8085 27924 8123 27958
rect 8157 27924 8195 27958
rect 8229 27924 8267 27958
rect 8301 27924 8339 27958
rect 8373 27924 8411 27958
rect 8445 27924 8483 27958
rect 8517 27924 8555 27958
rect 8589 27924 8627 27958
rect 8661 27924 8699 27958
rect 8733 27924 8771 27958
rect 8805 27924 8843 27958
rect 8877 27924 8915 27958
rect 8949 27924 8987 27958
rect 9021 27924 9059 27958
rect 9093 27924 9131 27958
rect 9165 27924 9203 27958
rect 9237 27924 9275 27958
rect 9309 27924 9347 27958
rect 9381 27924 9419 27958
rect 9453 27924 9491 27958
rect 9525 27924 9563 27958
rect 9597 27924 9635 27958
rect 9669 27924 9707 27958
rect 9741 27924 9779 27958
rect 9813 27924 9851 27958
rect 9885 27924 9923 27958
rect 9957 27924 9995 27958
rect 10029 27924 10067 27958
rect 10101 27924 10139 27958
rect 10173 27924 10211 27958
rect 10245 27924 10283 27958
rect 10317 27924 10355 27958
rect 10389 27924 10427 27958
rect 10461 27924 10499 27958
rect 10533 27924 10571 27958
rect 10605 27924 10643 27958
rect 10677 27924 10715 27958
rect 10749 27924 10787 27958
rect 10821 27924 10859 27958
rect 10893 27924 10931 27958
rect 10965 27924 11003 27958
rect 11037 27924 11075 27958
rect 11109 27924 11147 27958
rect 11181 27924 11219 27958
rect 11253 27924 11291 27958
rect 11325 27924 11363 27958
rect 11397 27924 11435 27958
rect 11469 27924 11507 27958
rect 11541 27924 11579 27958
rect 11613 27924 11651 27958
rect 11685 27924 11723 27958
rect 11757 27924 11795 27958
rect 11829 27924 11867 27958
rect 11901 27924 11939 27958
rect 11973 27924 12011 27958
rect 12045 27924 12083 27958
rect 12117 27924 12155 27958
rect 12209 27940 12225 27992
rect 12277 27940 12293 27992
rect 12345 27940 12361 27992
rect 12413 27940 12429 27992
rect 12481 27940 12497 27992
rect 12549 27940 12565 27992
rect 12617 27958 12633 27992
rect 12685 27958 12701 27992
rect 12753 27958 12768 27992
rect 12820 27958 12835 27992
rect 12887 27958 13929 27992
rect 12621 27940 12633 27958
rect 12693 27940 12701 27958
rect 12765 27940 12768 27958
rect 12189 27926 12227 27940
rect 12261 27926 12299 27940
rect 12333 27926 12371 27940
rect 12405 27926 12443 27940
rect 12477 27926 12515 27940
rect 12549 27926 12587 27940
rect 12621 27926 12659 27940
rect 12693 27926 12731 27940
rect 12765 27926 12803 27940
rect 12837 27926 12875 27940
rect 2033 27876 12157 27924
rect 1314 27860 1353 27874
rect 1387 27860 1426 27874
rect 1460 27860 1499 27874
rect 1533 27860 1571 27874
rect 1605 27860 1643 27874
rect 1677 27860 1715 27874
rect 1749 27860 1787 27874
rect 1821 27860 1859 27874
rect 1893 27860 1931 27874
rect 1965 27860 2003 27874
rect 1423 27842 1426 27860
rect 1491 27842 1499 27860
rect 1559 27842 1571 27860
rect 100 27808 1303 27842
rect 1355 27808 1371 27842
rect 1423 27808 1439 27842
rect 1491 27808 1507 27842
rect 1559 27808 1575 27842
rect 1627 27808 1643 27860
rect 1695 27808 1711 27860
rect 1763 27808 1779 27860
rect 1831 27808 1847 27860
rect 1899 27808 1914 27860
rect 1966 27808 1981 27860
rect 2037 27842 2075 27876
rect 2109 27842 2147 27876
rect 2181 27842 2219 27876
rect 2253 27842 2291 27876
rect 2325 27842 2363 27876
rect 2397 27842 2435 27876
rect 2469 27842 2507 27876
rect 2541 27842 2579 27876
rect 2613 27842 2651 27876
rect 2685 27842 2723 27876
rect 2757 27842 2795 27876
rect 2829 27842 2867 27876
rect 2901 27842 2939 27876
rect 2973 27842 3011 27876
rect 3045 27842 3083 27876
rect 3117 27842 3155 27876
rect 3189 27842 3227 27876
rect 3261 27842 3299 27876
rect 3333 27842 3371 27876
rect 3405 27842 3443 27876
rect 3477 27842 3515 27876
rect 3549 27842 3587 27876
rect 3621 27842 3659 27876
rect 3693 27842 3731 27876
rect 3765 27842 3803 27876
rect 3837 27842 3875 27876
rect 3909 27842 3947 27876
rect 3981 27842 4019 27876
rect 4053 27842 4091 27876
rect 4125 27842 4163 27876
rect 4197 27842 4235 27876
rect 4269 27842 4307 27876
rect 4341 27842 4379 27876
rect 4413 27842 4451 27876
rect 4485 27842 4523 27876
rect 4557 27842 4595 27876
rect 4629 27842 4667 27876
rect 4701 27842 4739 27876
rect 4773 27842 4811 27876
rect 4845 27842 4883 27876
rect 4917 27842 4955 27876
rect 4989 27842 5027 27876
rect 5061 27842 5099 27876
rect 5133 27842 5171 27876
rect 5205 27842 5243 27876
rect 5277 27842 5315 27876
rect 5349 27842 5387 27876
rect 5421 27842 5459 27876
rect 5493 27842 5531 27876
rect 5565 27842 5603 27876
rect 5637 27842 5675 27876
rect 5709 27842 5747 27876
rect 5781 27842 5819 27876
rect 5853 27842 5891 27876
rect 5925 27842 5963 27876
rect 5997 27842 6035 27876
rect 6069 27842 6107 27876
rect 6141 27842 6179 27876
rect 6213 27842 6251 27876
rect 6285 27842 6323 27876
rect 6357 27842 6395 27876
rect 6429 27842 6467 27876
rect 6501 27842 6539 27876
rect 6573 27842 6611 27876
rect 6645 27842 6683 27876
rect 6717 27842 6755 27876
rect 6789 27842 6827 27876
rect 6861 27842 6899 27876
rect 6933 27842 6971 27876
rect 7005 27842 7043 27876
rect 7077 27842 7115 27876
rect 7149 27842 7187 27876
rect 7221 27842 7259 27876
rect 7293 27842 7331 27876
rect 7365 27842 7403 27876
rect 7437 27842 7475 27876
rect 7509 27842 7547 27876
rect 7581 27842 7619 27876
rect 7653 27842 7691 27876
rect 7725 27842 7763 27876
rect 7797 27842 7835 27876
rect 7869 27842 7907 27876
rect 7941 27842 7979 27876
rect 8013 27842 8051 27876
rect 8085 27842 8123 27876
rect 8157 27842 8195 27876
rect 8229 27842 8267 27876
rect 8301 27842 8339 27876
rect 8373 27842 8411 27876
rect 8445 27842 8483 27876
rect 8517 27842 8555 27876
rect 8589 27842 8627 27876
rect 8661 27842 8699 27876
rect 8733 27842 8771 27876
rect 8805 27842 8843 27876
rect 8877 27842 8915 27876
rect 8949 27842 8987 27876
rect 9021 27842 9059 27876
rect 9093 27842 9131 27876
rect 9165 27842 9203 27876
rect 9237 27842 9275 27876
rect 9309 27842 9347 27876
rect 9381 27842 9419 27876
rect 9453 27842 9491 27876
rect 9525 27842 9563 27876
rect 9597 27842 9635 27876
rect 9669 27842 9707 27876
rect 9741 27842 9779 27876
rect 9813 27842 9851 27876
rect 9885 27842 9923 27876
rect 9957 27842 9995 27876
rect 10029 27842 10067 27876
rect 10101 27842 10139 27876
rect 10173 27842 10211 27876
rect 10245 27842 10283 27876
rect 10317 27842 10355 27876
rect 10389 27842 10427 27876
rect 10461 27842 10499 27876
rect 10533 27842 10571 27876
rect 10605 27842 10643 27876
rect 10677 27842 10715 27876
rect 10749 27842 10787 27876
rect 10821 27842 10859 27876
rect 10893 27842 10931 27876
rect 10965 27842 11003 27876
rect 11037 27842 11075 27876
rect 11109 27842 11147 27876
rect 11181 27842 11219 27876
rect 11253 27842 11291 27876
rect 11325 27842 11363 27876
rect 11397 27842 11435 27876
rect 11469 27842 11507 27876
rect 11541 27842 11579 27876
rect 11613 27842 11651 27876
rect 11685 27842 11723 27876
rect 11757 27842 11795 27876
rect 11829 27842 11867 27876
rect 11901 27842 11939 27876
rect 11973 27842 12011 27876
rect 12045 27842 12083 27876
rect 12117 27842 12155 27876
rect 12209 27874 12225 27926
rect 12277 27874 12293 27926
rect 12345 27874 12361 27926
rect 12413 27874 12429 27926
rect 12481 27874 12497 27926
rect 12549 27874 12565 27926
rect 12621 27924 12633 27926
rect 12693 27924 12701 27926
rect 12765 27924 12768 27926
rect 12909 27924 12947 27958
rect 12981 27924 13019 27958
rect 13053 27924 13091 27958
rect 13125 27924 13163 27958
rect 13197 27924 13235 27958
rect 13269 27924 13307 27958
rect 13341 27924 13379 27958
rect 13413 27924 13451 27958
rect 13485 27924 13523 27958
rect 13557 27924 13595 27958
rect 13629 27924 13667 27958
rect 13701 27924 13739 27958
rect 13773 27924 13811 27958
rect 13845 27924 13883 27958
rect 13917 27924 13929 27958
rect 12617 27876 12633 27924
rect 12685 27876 12701 27924
rect 12753 27876 12768 27924
rect 12820 27876 12835 27924
rect 12887 27876 13929 27924
rect 12621 27874 12633 27876
rect 12693 27874 12701 27876
rect 12765 27874 12768 27876
rect 12189 27860 12227 27874
rect 12261 27860 12299 27874
rect 12333 27860 12371 27874
rect 12405 27860 12443 27874
rect 12477 27860 12515 27874
rect 12549 27860 12587 27874
rect 12621 27860 12659 27874
rect 12693 27860 12731 27874
rect 12765 27860 12803 27874
rect 12837 27860 12875 27874
rect 2033 27808 12157 27842
rect 12209 27808 12225 27860
rect 12277 27808 12293 27860
rect 12345 27808 12361 27860
rect 12413 27808 12429 27860
rect 12481 27808 12497 27860
rect 12549 27808 12565 27860
rect 12621 27842 12633 27860
rect 12693 27842 12701 27860
rect 12765 27842 12768 27860
rect 12909 27842 12947 27876
rect 12981 27842 13019 27876
rect 13053 27842 13091 27876
rect 13125 27842 13163 27876
rect 13197 27842 13235 27876
rect 13269 27842 13307 27876
rect 13341 27842 13379 27876
rect 13413 27842 13451 27876
rect 13485 27842 13523 27876
rect 13557 27842 13595 27876
rect 13629 27842 13667 27876
rect 13701 27842 13739 27876
rect 13773 27842 13811 27876
rect 13845 27842 13883 27876
rect 13917 27842 13929 27876
rect 12617 27808 12633 27842
rect 12685 27808 12701 27842
rect 12753 27808 12768 27842
rect 12820 27808 12835 27842
rect 12887 27808 13929 27842
rect 100 27794 13929 27808
rect 100 27760 112 27794
rect 146 27760 185 27794
rect 219 27760 258 27794
rect 292 27760 331 27794
rect 365 27760 404 27794
rect 438 27760 477 27794
rect 511 27760 550 27794
rect 584 27760 623 27794
rect 657 27760 696 27794
rect 730 27760 769 27794
rect 803 27760 842 27794
rect 876 27760 915 27794
rect 949 27760 988 27794
rect 1022 27760 1061 27794
rect 1095 27760 1134 27794
rect 1168 27760 1207 27794
rect 1241 27760 1280 27794
rect 1423 27760 1426 27794
rect 1491 27760 1499 27794
rect 1559 27760 1571 27794
rect 100 27742 1303 27760
rect 1355 27742 1371 27760
rect 1423 27742 1439 27760
rect 1491 27742 1507 27760
rect 1559 27742 1575 27760
rect 1627 27742 1643 27794
rect 1695 27742 1711 27794
rect 1763 27742 1779 27794
rect 1831 27742 1847 27794
rect 1899 27742 1914 27794
rect 1966 27742 1981 27794
rect 2037 27760 2075 27794
rect 2109 27760 2147 27794
rect 2181 27760 2219 27794
rect 2253 27760 2291 27794
rect 2325 27760 2363 27794
rect 2397 27760 2435 27794
rect 2469 27760 2507 27794
rect 2541 27760 2579 27794
rect 2613 27760 2651 27794
rect 2685 27760 2723 27794
rect 2757 27760 2795 27794
rect 2829 27760 2867 27794
rect 2901 27760 2939 27794
rect 2973 27760 3011 27794
rect 3045 27760 3083 27794
rect 3117 27760 3155 27794
rect 3189 27760 3227 27794
rect 3261 27760 3299 27794
rect 3333 27760 3371 27794
rect 3405 27760 3443 27794
rect 3477 27760 3515 27794
rect 3549 27760 3587 27794
rect 3621 27760 3659 27794
rect 3693 27760 3731 27794
rect 3765 27760 3803 27794
rect 3837 27760 3875 27794
rect 3909 27760 3947 27794
rect 3981 27760 4019 27794
rect 4053 27760 4091 27794
rect 4125 27760 4163 27794
rect 4197 27760 4235 27794
rect 4269 27760 4307 27794
rect 4341 27760 4379 27794
rect 4413 27760 4451 27794
rect 4485 27760 4523 27794
rect 4557 27760 4595 27794
rect 4629 27760 4667 27794
rect 4701 27760 4739 27794
rect 4773 27760 4811 27794
rect 4845 27760 4883 27794
rect 4917 27760 4955 27794
rect 4989 27760 5027 27794
rect 5061 27760 5099 27794
rect 5133 27760 5171 27794
rect 5205 27760 5243 27794
rect 5277 27760 5315 27794
rect 5349 27760 5387 27794
rect 5421 27760 5459 27794
rect 5493 27760 5531 27794
rect 5565 27760 5603 27794
rect 5637 27760 5675 27794
rect 5709 27760 5747 27794
rect 5781 27760 5819 27794
rect 5853 27760 5891 27794
rect 5925 27760 5963 27794
rect 5997 27760 6035 27794
rect 6069 27760 6107 27794
rect 6141 27760 6179 27794
rect 6213 27760 6251 27794
rect 6285 27760 6323 27794
rect 6357 27760 6395 27794
rect 6429 27760 6467 27794
rect 6501 27760 6539 27794
rect 6573 27760 6611 27794
rect 6645 27760 6683 27794
rect 6717 27760 6755 27794
rect 6789 27760 6827 27794
rect 6861 27760 6899 27794
rect 6933 27760 6971 27794
rect 7005 27760 7043 27794
rect 7077 27760 7115 27794
rect 7149 27760 7187 27794
rect 7221 27760 7259 27794
rect 7293 27760 7331 27794
rect 7365 27760 7403 27794
rect 7437 27760 7475 27794
rect 7509 27760 7547 27794
rect 7581 27760 7619 27794
rect 7653 27760 7691 27794
rect 7725 27760 7763 27794
rect 7797 27760 7835 27794
rect 7869 27760 7907 27794
rect 7941 27760 7979 27794
rect 8013 27760 8051 27794
rect 8085 27760 8123 27794
rect 8157 27760 8195 27794
rect 8229 27760 8267 27794
rect 8301 27760 8339 27794
rect 8373 27760 8411 27794
rect 8445 27760 8483 27794
rect 8517 27760 8555 27794
rect 8589 27760 8627 27794
rect 8661 27760 8699 27794
rect 8733 27760 8771 27794
rect 8805 27760 8843 27794
rect 8877 27760 8915 27794
rect 8949 27760 8987 27794
rect 9021 27760 9059 27794
rect 9093 27760 9131 27794
rect 9165 27760 9203 27794
rect 9237 27760 9275 27794
rect 9309 27760 9347 27794
rect 9381 27760 9419 27794
rect 9453 27760 9491 27794
rect 9525 27760 9563 27794
rect 9597 27760 9635 27794
rect 9669 27760 9707 27794
rect 9741 27760 9779 27794
rect 9813 27760 9851 27794
rect 9885 27760 9923 27794
rect 9957 27760 9995 27794
rect 10029 27760 10067 27794
rect 10101 27760 10139 27794
rect 10173 27760 10211 27794
rect 10245 27760 10283 27794
rect 10317 27760 10355 27794
rect 10389 27760 10427 27794
rect 10461 27760 10499 27794
rect 10533 27760 10571 27794
rect 10605 27760 10643 27794
rect 10677 27760 10715 27794
rect 10749 27760 10787 27794
rect 10821 27760 10859 27794
rect 10893 27760 10931 27794
rect 10965 27760 11003 27794
rect 11037 27760 11075 27794
rect 11109 27760 11147 27794
rect 11181 27760 11219 27794
rect 11253 27760 11291 27794
rect 11325 27760 11363 27794
rect 11397 27760 11435 27794
rect 11469 27760 11507 27794
rect 11541 27760 11579 27794
rect 11613 27760 11651 27794
rect 11685 27760 11723 27794
rect 11757 27760 11795 27794
rect 11829 27760 11867 27794
rect 11901 27760 11939 27794
rect 11973 27760 12011 27794
rect 12045 27760 12083 27794
rect 12117 27760 12155 27794
rect 2033 27742 12157 27760
rect 12209 27742 12225 27794
rect 12277 27742 12293 27794
rect 12345 27742 12361 27794
rect 12413 27742 12429 27794
rect 12481 27742 12497 27794
rect 12549 27742 12565 27794
rect 12621 27760 12633 27794
rect 12693 27760 12701 27794
rect 12765 27760 12768 27794
rect 12909 27760 12947 27794
rect 12981 27760 13019 27794
rect 13053 27760 13091 27794
rect 13125 27760 13163 27794
rect 13197 27760 13235 27794
rect 13269 27760 13307 27794
rect 13341 27760 13379 27794
rect 13413 27760 13451 27794
rect 13485 27760 13523 27794
rect 13557 27760 13595 27794
rect 13629 27760 13667 27794
rect 13701 27760 13739 27794
rect 13773 27760 13811 27794
rect 13845 27760 13883 27794
rect 13917 27760 13929 27794
rect 12617 27742 12633 27760
rect 12685 27742 12701 27760
rect 12753 27742 12768 27760
rect 12820 27742 12835 27760
rect 12887 27742 13929 27760
rect 100 27728 13929 27742
rect 100 27712 1303 27728
rect 1355 27712 1371 27728
rect 1423 27712 1439 27728
rect 1491 27712 1507 27728
rect 1559 27712 1575 27728
rect 100 27678 112 27712
rect 146 27678 185 27712
rect 219 27678 258 27712
rect 292 27678 331 27712
rect 365 27678 404 27712
rect 438 27678 477 27712
rect 511 27678 550 27712
rect 584 27678 623 27712
rect 657 27678 696 27712
rect 730 27678 769 27712
rect 803 27678 842 27712
rect 876 27678 915 27712
rect 949 27678 988 27712
rect 1022 27678 1061 27712
rect 1095 27678 1134 27712
rect 1168 27678 1207 27712
rect 1241 27678 1280 27712
rect 1423 27678 1426 27712
rect 1491 27678 1499 27712
rect 1559 27678 1571 27712
rect 100 27676 1303 27678
rect 1355 27676 1371 27678
rect 1423 27676 1439 27678
rect 1491 27676 1507 27678
rect 1559 27676 1575 27678
rect 1627 27676 1643 27728
rect 1695 27676 1711 27728
rect 1763 27676 1779 27728
rect 1831 27676 1847 27728
rect 1899 27676 1914 27728
rect 1966 27676 1981 27728
rect 2033 27712 12157 27728
rect 2037 27678 2075 27712
rect 2109 27678 2147 27712
rect 2181 27678 2219 27712
rect 2253 27678 2291 27712
rect 2325 27678 2363 27712
rect 2397 27678 2435 27712
rect 2469 27678 2507 27712
rect 2541 27678 2579 27712
rect 2613 27678 2651 27712
rect 2685 27678 2723 27712
rect 2757 27678 2795 27712
rect 2829 27678 2867 27712
rect 2901 27678 2939 27712
rect 2973 27678 3011 27712
rect 3045 27678 3083 27712
rect 3117 27678 3155 27712
rect 3189 27678 3227 27712
rect 3261 27678 3299 27712
rect 3333 27678 3371 27712
rect 3405 27678 3443 27712
rect 3477 27678 3515 27712
rect 3549 27678 3587 27712
rect 3621 27678 3659 27712
rect 3693 27678 3731 27712
rect 3765 27678 3803 27712
rect 3837 27678 3875 27712
rect 3909 27678 3947 27712
rect 3981 27678 4019 27712
rect 4053 27678 4091 27712
rect 4125 27678 4163 27712
rect 4197 27678 4235 27712
rect 4269 27678 4307 27712
rect 4341 27678 4379 27712
rect 4413 27678 4451 27712
rect 4485 27678 4523 27712
rect 4557 27678 4595 27712
rect 4629 27678 4667 27712
rect 4701 27678 4739 27712
rect 4773 27678 4811 27712
rect 4845 27678 4883 27712
rect 4917 27678 4955 27712
rect 4989 27678 5027 27712
rect 5061 27678 5099 27712
rect 5133 27678 5171 27712
rect 5205 27678 5243 27712
rect 5277 27678 5315 27712
rect 5349 27678 5387 27712
rect 5421 27678 5459 27712
rect 5493 27678 5531 27712
rect 5565 27678 5603 27712
rect 5637 27678 5675 27712
rect 5709 27678 5747 27712
rect 5781 27678 5819 27712
rect 5853 27678 5891 27712
rect 5925 27678 5963 27712
rect 5997 27678 6035 27712
rect 6069 27678 6107 27712
rect 6141 27678 6179 27712
rect 6213 27678 6251 27712
rect 6285 27678 6323 27712
rect 6357 27678 6395 27712
rect 6429 27678 6467 27712
rect 6501 27678 6539 27712
rect 6573 27678 6611 27712
rect 6645 27678 6683 27712
rect 6717 27678 6755 27712
rect 6789 27678 6827 27712
rect 6861 27678 6899 27712
rect 6933 27678 6971 27712
rect 7005 27678 7043 27712
rect 7077 27678 7115 27712
rect 7149 27678 7187 27712
rect 7221 27678 7259 27712
rect 7293 27678 7331 27712
rect 7365 27678 7403 27712
rect 7437 27678 7475 27712
rect 7509 27678 7547 27712
rect 7581 27678 7619 27712
rect 7653 27678 7691 27712
rect 7725 27678 7763 27712
rect 7797 27678 7835 27712
rect 7869 27678 7907 27712
rect 7941 27678 7979 27712
rect 8013 27678 8051 27712
rect 8085 27678 8123 27712
rect 8157 27678 8195 27712
rect 8229 27678 8267 27712
rect 8301 27678 8339 27712
rect 8373 27678 8411 27712
rect 8445 27678 8483 27712
rect 8517 27678 8555 27712
rect 8589 27678 8627 27712
rect 8661 27678 8699 27712
rect 8733 27678 8771 27712
rect 8805 27678 8843 27712
rect 8877 27678 8915 27712
rect 8949 27678 8987 27712
rect 9021 27678 9059 27712
rect 9093 27678 9131 27712
rect 9165 27678 9203 27712
rect 9237 27678 9275 27712
rect 9309 27678 9347 27712
rect 9381 27678 9419 27712
rect 9453 27678 9491 27712
rect 9525 27678 9563 27712
rect 9597 27678 9635 27712
rect 9669 27678 9707 27712
rect 9741 27678 9779 27712
rect 9813 27678 9851 27712
rect 9885 27678 9923 27712
rect 9957 27678 9995 27712
rect 10029 27678 10067 27712
rect 10101 27678 10139 27712
rect 10173 27678 10211 27712
rect 10245 27678 10283 27712
rect 10317 27678 10355 27712
rect 10389 27678 10427 27712
rect 10461 27678 10499 27712
rect 10533 27678 10571 27712
rect 10605 27678 10643 27712
rect 10677 27678 10715 27712
rect 10749 27678 10787 27712
rect 10821 27678 10859 27712
rect 10893 27678 10931 27712
rect 10965 27678 11003 27712
rect 11037 27678 11075 27712
rect 11109 27678 11147 27712
rect 11181 27678 11219 27712
rect 11253 27678 11291 27712
rect 11325 27678 11363 27712
rect 11397 27678 11435 27712
rect 11469 27678 11507 27712
rect 11541 27678 11579 27712
rect 11613 27678 11651 27712
rect 11685 27678 11723 27712
rect 11757 27678 11795 27712
rect 11829 27678 11867 27712
rect 11901 27678 11939 27712
rect 11973 27678 12011 27712
rect 12045 27678 12083 27712
rect 12117 27678 12155 27712
rect 2033 27676 12157 27678
rect 12209 27676 12225 27728
rect 12277 27676 12293 27728
rect 12345 27676 12361 27728
rect 12413 27676 12429 27728
rect 12481 27676 12497 27728
rect 12549 27676 12565 27728
rect 12617 27712 12633 27728
rect 12685 27712 12701 27728
rect 12753 27712 12768 27728
rect 12820 27712 12835 27728
rect 12887 27712 13929 27728
rect 12621 27678 12633 27712
rect 12693 27678 12701 27712
rect 12765 27678 12768 27712
rect 12909 27678 12947 27712
rect 12981 27678 13019 27712
rect 13053 27678 13091 27712
rect 13125 27678 13163 27712
rect 13197 27678 13235 27712
rect 13269 27678 13307 27712
rect 13341 27678 13379 27712
rect 13413 27678 13451 27712
rect 13485 27678 13523 27712
rect 13557 27678 13595 27712
rect 13629 27678 13667 27712
rect 13701 27678 13739 27712
rect 13773 27678 13811 27712
rect 13845 27678 13883 27712
rect 13917 27678 13929 27712
rect 12617 27676 12633 27678
rect 12685 27676 12701 27678
rect 12753 27676 12768 27678
rect 12820 27676 12835 27678
rect 12887 27676 13929 27678
rect 100 27671 13929 27676
rect 14281 28119 14282 28171
rect 14334 28119 14358 28171
rect 14410 28119 14434 28171
rect 14486 28119 14510 28171
rect 14562 28119 14586 28171
rect 14638 28119 15029 28171
rect 14281 28105 15029 28119
rect 14281 28053 14282 28105
rect 14334 28053 14358 28105
rect 14410 28053 14434 28105
rect 14486 28053 14510 28105
rect 14562 28053 14586 28105
rect 14638 28053 15029 28105
rect 14281 28039 15029 28053
rect 14281 27987 14282 28039
rect 14334 27987 14358 28039
rect 14410 27987 14434 28039
rect 14486 27987 14510 28039
rect 14562 27987 14586 28039
rect 14638 27987 15029 28039
rect 14281 27973 15029 27987
rect 14281 27921 14282 27973
rect 14334 27921 14358 27973
rect 14410 27921 14434 27973
rect 14486 27921 14510 27973
rect 14562 27921 14586 27973
rect 14638 27921 15029 27973
rect 14281 27907 15029 27921
rect 14281 27855 14282 27907
rect 14334 27855 14358 27907
rect 14410 27855 14434 27907
rect 14486 27855 14510 27907
rect 14562 27855 14586 27907
rect 14638 27855 15029 27907
rect 14281 27841 15029 27855
rect 14281 27789 14282 27841
rect 14334 27789 14358 27841
rect 14410 27789 14434 27841
rect 14486 27789 14510 27841
rect 14562 27789 14586 27841
rect 14638 27789 15029 27841
rect 14281 27775 15029 27789
rect 14281 27723 14282 27775
rect 14334 27723 14358 27775
rect 14410 27723 14434 27775
rect 14486 27723 14510 27775
rect 14562 27723 14586 27775
rect 14638 27723 15029 27775
rect 14281 27709 15029 27723
rect 14281 27657 14282 27709
rect 14334 27657 14358 27709
rect 14410 27657 14434 27709
rect 14486 27657 14510 27709
rect 14562 27657 14586 27709
rect 14638 27657 15029 27709
tri 14000 27370 14281 27651 se
rect 14281 27643 15029 27657
rect 14281 27591 14282 27643
rect 14334 27591 14358 27643
rect 14410 27591 14434 27643
rect 14486 27591 14510 27643
rect 14562 27591 14586 27643
rect 14638 27591 15029 27643
rect 14281 27577 15029 27591
rect 14281 27525 14282 27577
rect 14334 27525 14358 27577
rect 14410 27525 14434 27577
rect 14486 27525 14510 27577
rect 14562 27525 14586 27577
rect 14638 27525 15029 27577
rect 14281 27511 15029 27525
rect 14281 27459 14282 27511
rect 14334 27459 14358 27511
rect 14410 27459 14434 27511
rect 14486 27459 14510 27511
rect 14562 27459 14586 27511
rect 14638 27459 15029 27511
rect 14281 27445 15029 27459
rect 14281 27393 14282 27445
rect 14334 27393 14358 27445
rect 14410 27393 14434 27445
rect 14486 27393 14510 27445
rect 14562 27393 14586 27445
rect 14638 27393 15029 27445
rect 14281 27379 15029 27393
rect 14281 27370 14282 27379
rect 0 27369 14282 27370
rect 0 27362 3478 27369
rect 3530 27362 3546 27369
rect 3598 27362 3614 27369
rect 0 27355 827 27362
rect 0 27321 163 27355
rect 197 27321 237 27355
rect 271 27321 311 27355
rect 345 27321 385 27355
rect 419 27321 459 27355
rect 493 27321 533 27355
rect 567 27321 606 27355
rect 640 27321 679 27355
rect 713 27321 752 27355
rect 786 27328 827 27355
rect 861 27328 899 27362
rect 933 27328 971 27362
rect 1005 27328 1043 27362
rect 1077 27328 1115 27362
rect 1149 27328 1187 27362
rect 1221 27328 1259 27362
rect 1293 27328 1331 27362
rect 1365 27328 1403 27362
rect 1437 27328 1475 27362
rect 1509 27328 1547 27362
rect 1581 27328 1619 27362
rect 1653 27328 1691 27362
rect 1725 27328 1764 27362
rect 1798 27328 1837 27362
rect 1871 27328 1910 27362
rect 1944 27328 1983 27362
rect 2017 27328 2056 27362
rect 2090 27355 3392 27362
rect 2090 27328 2142 27355
rect 786 27321 2142 27328
rect 2176 27321 2221 27355
rect 2255 27321 2300 27355
rect 2334 27321 2379 27355
rect 2413 27321 2458 27355
rect 2492 27321 2536 27355
rect 2570 27321 2614 27355
rect 2648 27321 2692 27355
rect 2726 27321 2770 27355
rect 2804 27321 2848 27355
rect 2882 27321 2926 27355
rect 2960 27328 3392 27355
rect 3426 27328 3465 27362
rect 3530 27328 3538 27362
rect 3598 27328 3611 27362
rect 2960 27321 3478 27328
rect 0 27317 3478 27321
rect 3530 27317 3546 27328
rect 3598 27317 3614 27328
rect 3666 27317 3682 27369
rect 3734 27317 3750 27369
rect 3802 27317 3818 27369
rect 3870 27317 3886 27369
rect 3938 27317 3954 27369
rect 4006 27362 4021 27369
rect 4073 27362 4088 27369
rect 4140 27362 4155 27369
rect 4207 27362 4222 27369
rect 4274 27362 4289 27369
rect 4341 27362 4356 27369
rect 4408 27362 4423 27369
rect 4475 27362 4490 27369
rect 4542 27362 4557 27369
rect 4609 27362 5461 27369
rect 5513 27362 5529 27369
rect 5581 27362 5597 27369
rect 5649 27362 5665 27369
rect 5717 27362 5733 27369
rect 5785 27362 5801 27369
rect 5853 27362 5869 27369
rect 5921 27362 5937 27369
rect 5989 27362 6004 27369
rect 6056 27362 6071 27369
rect 4010 27328 4021 27362
rect 4083 27328 4088 27362
rect 4408 27328 4410 27362
rect 4475 27328 4482 27362
rect 4542 27328 4554 27362
rect 4609 27328 4626 27362
rect 4660 27328 4698 27362
rect 4732 27328 4770 27362
rect 4804 27328 4842 27362
rect 4876 27328 4914 27362
rect 4948 27328 4986 27362
rect 5020 27328 5058 27362
rect 5092 27328 5130 27362
rect 5164 27328 5202 27362
rect 5236 27328 5274 27362
rect 5308 27328 5346 27362
rect 5380 27328 5418 27362
rect 5452 27328 5461 27362
rect 5524 27328 5529 27362
rect 5596 27328 5597 27362
rect 5921 27328 5922 27362
rect 5989 27328 5994 27362
rect 6056 27328 6066 27362
rect 4006 27317 4021 27328
rect 4073 27317 4088 27328
rect 4140 27317 4155 27328
rect 4207 27317 4222 27328
rect 4274 27317 4289 27328
rect 4341 27317 4356 27328
rect 4408 27317 4423 27328
rect 4475 27317 4490 27328
rect 4542 27317 4557 27328
rect 4609 27317 5461 27328
rect 5513 27317 5529 27328
rect 5581 27317 5597 27328
rect 5649 27317 5665 27328
rect 5717 27317 5733 27328
rect 5785 27317 5801 27328
rect 5853 27317 5869 27328
rect 5921 27317 5937 27328
rect 5989 27317 6004 27328
rect 6056 27317 6071 27328
rect 6123 27317 6138 27369
rect 6190 27317 6205 27369
rect 6257 27317 6272 27369
rect 6324 27317 6339 27369
rect 6391 27317 6406 27369
rect 6458 27362 6473 27369
rect 6525 27362 6540 27369
rect 6592 27362 7445 27369
rect 7497 27362 7513 27369
rect 7565 27362 7581 27369
rect 6460 27328 6473 27362
rect 6532 27328 6540 27362
rect 6604 27328 6642 27362
rect 6676 27328 6714 27362
rect 6748 27328 6786 27362
rect 6820 27328 6858 27362
rect 6892 27328 6930 27362
rect 6964 27328 7002 27362
rect 7036 27328 7074 27362
rect 7108 27328 7146 27362
rect 7180 27328 7218 27362
rect 7252 27328 7290 27362
rect 7324 27328 7362 27362
rect 7396 27328 7434 27362
rect 7497 27328 7506 27362
rect 7565 27328 7578 27362
rect 6458 27317 6473 27328
rect 6525 27317 6540 27328
rect 6592 27317 7445 27328
rect 7497 27317 7513 27328
rect 7565 27317 7581 27328
rect 7633 27317 7649 27369
rect 7701 27317 7717 27369
rect 7769 27317 7785 27369
rect 7837 27317 7853 27369
rect 7905 27317 7921 27369
rect 7973 27317 7988 27369
rect 8040 27362 8055 27369
rect 8107 27362 8122 27369
rect 8174 27362 8189 27369
rect 8241 27362 8256 27369
rect 8308 27362 8323 27369
rect 8375 27362 8390 27369
rect 8442 27362 8457 27369
rect 8509 27362 8524 27369
rect 8576 27364 14282 27369
rect 8576 27362 9423 27364
rect 9475 27362 9523 27364
rect 9575 27362 14282 27364
rect 14334 27362 14358 27379
rect 14410 27362 14434 27379
rect 14486 27362 14510 27379
rect 14562 27362 14586 27379
rect 14638 27362 15029 27379
rect 8044 27328 8055 27362
rect 8116 27328 8122 27362
rect 8188 27328 8189 27362
rect 8509 27328 8514 27362
rect 8576 27328 8586 27362
rect 8620 27328 8658 27362
rect 8692 27328 8730 27362
rect 8764 27328 8802 27362
rect 8836 27328 8874 27362
rect 8908 27328 8946 27362
rect 8980 27328 9018 27362
rect 9052 27328 9090 27362
rect 9124 27328 9162 27362
rect 9196 27328 9234 27362
rect 9268 27328 9306 27362
rect 9340 27328 9378 27362
rect 9412 27328 9423 27362
rect 9484 27328 9522 27362
rect 9575 27328 9594 27362
rect 9628 27328 9666 27362
rect 9700 27328 9738 27362
rect 9772 27328 9810 27362
rect 9844 27328 9882 27362
rect 9916 27328 9954 27362
rect 9988 27328 10026 27362
rect 10060 27328 10098 27362
rect 10132 27328 10170 27362
rect 10204 27328 10242 27362
rect 10276 27328 10314 27362
rect 10348 27328 10386 27362
rect 10420 27328 10458 27362
rect 10492 27328 10530 27362
rect 10564 27328 10602 27362
rect 10636 27328 10674 27362
rect 10708 27328 10746 27362
rect 10780 27328 10818 27362
rect 10852 27328 10890 27362
rect 10924 27328 10962 27362
rect 10996 27328 11034 27362
rect 11068 27328 11106 27362
rect 11140 27328 11178 27362
rect 11212 27328 11250 27362
rect 11284 27328 11322 27362
rect 11356 27328 11394 27362
rect 11428 27328 11466 27362
rect 11500 27328 11538 27362
rect 11572 27328 11610 27362
rect 11644 27328 11682 27362
rect 11716 27328 11754 27362
rect 11788 27328 11826 27362
rect 11860 27328 11898 27362
rect 11932 27328 11970 27362
rect 12004 27328 12042 27362
rect 12076 27328 12114 27362
rect 12148 27328 12186 27362
rect 12220 27328 12258 27362
rect 12292 27328 12330 27362
rect 12364 27328 12402 27362
rect 12436 27328 12474 27362
rect 12508 27328 12546 27362
rect 12580 27328 12618 27362
rect 12652 27328 12690 27362
rect 12724 27328 12762 27362
rect 12796 27328 12834 27362
rect 12868 27328 12906 27362
rect 12940 27328 12978 27362
rect 13012 27328 13050 27362
rect 13084 27328 13122 27362
rect 13156 27328 13194 27362
rect 13228 27328 13266 27362
rect 13300 27328 13338 27362
rect 13372 27328 13410 27362
rect 13444 27328 13482 27362
rect 13516 27328 13554 27362
rect 13588 27328 13626 27362
rect 13660 27328 13698 27362
rect 13732 27328 13770 27362
rect 13804 27328 13842 27362
rect 13876 27328 13914 27362
rect 13948 27328 13986 27362
rect 14020 27328 14058 27362
rect 14092 27328 14130 27362
rect 14164 27328 14202 27362
rect 14236 27328 14274 27362
rect 14334 27328 14346 27362
rect 14410 27328 14418 27362
rect 14486 27328 14490 27362
rect 14668 27328 14706 27362
rect 14740 27328 14778 27362
rect 14812 27328 14850 27362
rect 14884 27328 15029 27362
rect 8040 27317 8055 27328
rect 8107 27317 8122 27328
rect 8174 27317 8189 27328
rect 8241 27317 8256 27328
rect 8308 27317 8323 27328
rect 8375 27317 8390 27328
rect 8442 27317 8457 27328
rect 8509 27317 8524 27328
rect 8576 27317 9423 27328
rect 0 27315 9423 27317
rect 0 27301 2158 27315
tri 643 27238 706 27301 ne
rect 706 27238 2158 27301
tri 2158 27238 2235 27315 nw
tri 3259 27238 3336 27315 ne
rect 3336 27312 9423 27315
rect 9475 27312 9523 27328
rect 9575 27327 14282 27328
rect 14334 27327 14358 27328
rect 14410 27327 14434 27328
rect 14486 27327 14510 27328
rect 14562 27327 14586 27328
rect 14638 27327 15029 27328
rect 9575 27313 15029 27327
rect 9575 27312 14282 27313
rect 3336 27268 14282 27312
rect 3336 27243 9423 27268
rect 3336 27238 3478 27243
rect 3530 27238 3546 27243
rect 3598 27238 3614 27243
tri 706 27204 740 27238 ne
rect 740 27204 827 27238
rect 861 27204 899 27238
rect 933 27204 971 27238
rect 1005 27204 1043 27238
rect 1077 27204 1115 27238
rect 1149 27204 1187 27238
rect 1221 27204 1259 27238
rect 1293 27204 1331 27238
rect 1365 27204 1403 27238
rect 1437 27204 1475 27238
rect 1509 27204 1547 27238
rect 1581 27204 1619 27238
rect 1653 27204 1691 27238
rect 1725 27204 1764 27238
rect 1798 27204 1837 27238
rect 1871 27204 1910 27238
rect 1944 27204 1983 27238
rect 2017 27204 2056 27238
rect 2090 27204 2124 27238
tri 2124 27204 2158 27238 nw
tri 3336 27204 3370 27238 ne
rect 3370 27204 3392 27238
rect 3426 27204 3465 27238
rect 3530 27204 3538 27238
rect 3598 27204 3611 27238
tri 740 27198 746 27204 ne
rect 746 27198 2118 27204
tri 2118 27198 2124 27204 nw
tri 3370 27198 3376 27204 ne
rect 3376 27198 3478 27204
tri 746 27189 755 27198 ne
rect 755 27189 2109 27198
tri 2109 27189 2118 27198 nw
tri 3376 27189 3385 27198 ne
rect 3385 27191 3478 27198
rect 3530 27191 3546 27204
rect 3598 27191 3614 27204
rect 3666 27191 3682 27243
rect 3734 27191 3750 27243
rect 3802 27191 3818 27243
rect 3870 27191 3886 27243
rect 3938 27191 3954 27243
rect 4006 27238 4021 27243
rect 4073 27238 4088 27243
rect 4140 27238 4155 27243
rect 4207 27238 4222 27243
rect 4274 27238 4289 27243
rect 4341 27238 4356 27243
rect 4408 27238 4423 27243
rect 4475 27238 4490 27243
rect 4542 27238 4557 27243
rect 4609 27238 5461 27243
rect 5513 27238 5529 27243
rect 5581 27238 5597 27243
rect 5649 27238 5665 27243
rect 5717 27238 5733 27243
rect 5785 27238 5801 27243
rect 5853 27238 5869 27243
rect 5921 27238 5937 27243
rect 5989 27238 6004 27243
rect 6056 27238 6071 27243
rect 4010 27204 4021 27238
rect 4083 27204 4088 27238
rect 4408 27204 4410 27238
rect 4475 27204 4482 27238
rect 4542 27204 4554 27238
rect 4609 27204 4626 27238
rect 4660 27204 4698 27238
rect 4732 27204 4770 27238
rect 4804 27204 4842 27238
rect 4876 27204 4914 27238
rect 4948 27204 4986 27238
rect 5020 27204 5058 27238
rect 5092 27204 5130 27238
rect 5164 27204 5202 27238
rect 5236 27204 5274 27238
rect 5308 27204 5346 27238
rect 5380 27204 5418 27238
rect 5452 27204 5461 27238
rect 5524 27204 5529 27238
rect 5596 27204 5597 27238
rect 5921 27204 5922 27238
rect 5989 27204 5994 27238
rect 6056 27204 6066 27238
rect 4006 27191 4021 27204
rect 4073 27191 4088 27204
rect 4140 27191 4155 27204
rect 4207 27191 4222 27204
rect 4274 27191 4289 27204
rect 4341 27191 4356 27204
rect 4408 27191 4423 27204
rect 4475 27191 4490 27204
rect 4542 27191 4557 27204
rect 4609 27191 5461 27204
rect 5513 27191 5529 27204
rect 5581 27191 5597 27204
rect 5649 27191 5665 27204
rect 5717 27191 5733 27204
rect 5785 27191 5801 27204
rect 5853 27191 5869 27204
rect 5921 27191 5937 27204
rect 5989 27191 6004 27204
rect 6056 27191 6071 27204
rect 6123 27191 6138 27243
rect 6190 27191 6205 27243
rect 6257 27191 6272 27243
rect 6324 27191 6339 27243
rect 6391 27191 6406 27243
rect 6458 27238 6473 27243
rect 6525 27238 6540 27243
rect 6592 27238 7445 27243
rect 7497 27238 7513 27243
rect 7565 27238 7581 27243
rect 6460 27204 6473 27238
rect 6532 27204 6540 27238
rect 6604 27204 6642 27238
rect 6676 27204 6714 27238
rect 6748 27204 6786 27238
rect 6820 27204 6858 27238
rect 6892 27204 6930 27238
rect 6964 27204 7002 27238
rect 7036 27204 7074 27238
rect 7108 27204 7146 27238
rect 7180 27204 7218 27238
rect 7252 27204 7290 27238
rect 7324 27204 7362 27238
rect 7396 27204 7434 27238
rect 7497 27204 7506 27238
rect 7565 27204 7578 27238
rect 6458 27191 6473 27204
rect 6525 27191 6540 27204
rect 6592 27191 7445 27204
rect 7497 27191 7513 27204
rect 7565 27191 7581 27204
rect 7633 27191 7649 27243
rect 7701 27191 7717 27243
rect 7769 27191 7785 27243
rect 7837 27191 7853 27243
rect 7905 27191 7921 27243
rect 7973 27191 7988 27243
rect 8040 27238 8055 27243
rect 8107 27238 8122 27243
rect 8174 27238 8189 27243
rect 8241 27238 8256 27243
rect 8308 27238 8323 27243
rect 8375 27238 8390 27243
rect 8442 27238 8457 27243
rect 8509 27238 8524 27243
rect 8576 27238 9423 27243
rect 9475 27238 9523 27268
rect 9575 27261 14282 27268
rect 14334 27261 14358 27313
rect 14410 27261 14434 27313
rect 14486 27261 14510 27313
rect 14562 27261 14586 27313
rect 14638 27261 15029 27313
rect 9575 27247 15029 27261
rect 9575 27238 14282 27247
rect 14334 27238 14358 27247
rect 14410 27238 14434 27247
rect 14486 27238 14510 27247
rect 14562 27238 14586 27247
rect 14638 27238 15029 27247
rect 8044 27204 8055 27238
rect 8116 27204 8122 27238
rect 8188 27204 8189 27238
rect 8509 27204 8514 27238
rect 8576 27204 8586 27238
rect 8620 27204 8658 27238
rect 8692 27204 8730 27238
rect 8764 27204 8802 27238
rect 8836 27204 8874 27238
rect 8908 27204 8946 27238
rect 8980 27204 9018 27238
rect 9052 27204 9090 27238
rect 9124 27204 9162 27238
rect 9196 27204 9234 27238
rect 9268 27204 9306 27238
rect 9340 27204 9378 27238
rect 9412 27216 9423 27238
rect 9412 27204 9450 27216
rect 9484 27204 9522 27238
rect 9575 27216 9594 27238
rect 9556 27204 9594 27216
rect 9628 27204 9666 27238
rect 9700 27204 9738 27238
rect 9772 27204 9810 27238
rect 9844 27204 9882 27238
rect 9916 27204 9954 27238
rect 9988 27204 10026 27238
rect 10060 27204 10098 27238
rect 10132 27204 10170 27238
rect 10204 27204 10242 27238
rect 10276 27204 10314 27238
rect 10348 27204 10386 27238
rect 10420 27204 10458 27238
rect 10492 27204 10530 27238
rect 10564 27204 10602 27238
rect 10636 27204 10674 27238
rect 10708 27204 10746 27238
rect 10780 27204 10818 27238
rect 10852 27204 10890 27238
rect 10924 27204 10962 27238
rect 10996 27204 11034 27238
rect 11068 27204 11106 27238
rect 11140 27204 11178 27238
rect 11212 27204 11250 27238
rect 11284 27204 11322 27238
rect 11356 27204 11394 27238
rect 11428 27204 11466 27238
rect 11500 27204 11538 27238
rect 11572 27204 11610 27238
rect 11644 27204 11682 27238
rect 11716 27204 11754 27238
rect 11788 27204 11826 27238
rect 11860 27204 11898 27238
rect 11932 27204 11970 27238
rect 12004 27204 12042 27238
rect 12076 27204 12114 27238
rect 12148 27204 12186 27238
rect 12220 27204 12258 27238
rect 12292 27204 12330 27238
rect 12364 27204 12402 27238
rect 12436 27204 12474 27238
rect 12508 27204 12546 27238
rect 12580 27204 12618 27238
rect 12652 27204 12690 27238
rect 12724 27204 12762 27238
rect 12796 27204 12834 27238
rect 12868 27204 12906 27238
rect 12940 27204 12978 27238
rect 13012 27204 13050 27238
rect 13084 27204 13122 27238
rect 13156 27204 13194 27238
rect 13228 27204 13266 27238
rect 13300 27204 13338 27238
rect 13372 27204 13410 27238
rect 13444 27204 13482 27238
rect 13516 27204 13554 27238
rect 13588 27204 13626 27238
rect 13660 27204 13698 27238
rect 13732 27204 13770 27238
rect 13804 27204 13842 27238
rect 13876 27204 13914 27238
rect 13948 27204 13986 27238
rect 14020 27204 14058 27238
rect 14092 27204 14130 27238
rect 14164 27204 14202 27238
rect 14236 27204 14274 27238
rect 14334 27204 14346 27238
rect 14410 27204 14418 27238
rect 14486 27204 14490 27238
rect 14668 27204 14706 27238
rect 14740 27204 14778 27238
rect 14812 27204 14850 27238
rect 14884 27204 15029 27238
rect 8040 27191 8055 27204
rect 8107 27191 8122 27204
rect 8174 27191 8189 27204
rect 8241 27191 8256 27204
rect 8308 27191 8323 27204
rect 8375 27191 8390 27204
rect 8442 27191 8457 27204
rect 8509 27191 8524 27204
rect 8576 27195 14282 27204
rect 14334 27195 14358 27204
rect 14410 27195 14434 27204
rect 14486 27195 14510 27204
rect 14562 27195 14586 27204
rect 14638 27195 15029 27204
rect 8576 27191 15029 27195
rect 3385 27189 15029 27191
rect 2359 26948 2365 27000
rect 2417 26948 2440 27000
rect 2492 26948 2515 27000
rect 2567 26948 2589 27000
rect 2641 26948 2663 27000
rect 2715 26948 2721 27000
rect 2359 26878 2721 26948
rect 2359 26826 2365 26878
rect 2417 26826 2440 26878
rect 2492 26826 2515 26878
rect 2567 26826 2589 26878
rect 2641 26826 2663 26878
rect 2715 26826 2721 26878
rect 231 26185 14736 26193
rect 231 26151 243 26185
rect 277 26151 316 26185
rect 350 26151 389 26185
rect 423 26151 462 26185
rect 496 26151 535 26185
rect 569 26151 608 26185
rect 642 26151 681 26185
rect 715 26151 754 26185
rect 788 26151 827 26185
rect 861 26151 900 26185
rect 934 26151 973 26185
rect 1007 26151 1046 26185
rect 1080 26151 1119 26185
rect 1153 26151 1192 26185
rect 1226 26151 1265 26185
rect 1299 26151 1338 26185
rect 1372 26151 1411 26185
rect 1445 26151 1484 26185
rect 1518 26151 1557 26185
rect 1591 26151 1630 26185
rect 1664 26151 1703 26185
rect 1737 26151 1776 26185
rect 1810 26151 1849 26185
rect 1883 26151 1922 26185
rect 1956 26151 1995 26185
rect 2029 26151 2068 26185
rect 2102 26151 2141 26185
rect 2175 26151 2214 26185
rect 2248 26151 2287 26185
rect 2321 26151 2360 26185
rect 2394 26151 2433 26185
rect 2467 26181 2506 26185
rect 2540 26181 2579 26185
rect 2613 26181 2652 26185
rect 2467 26151 2480 26181
rect 2540 26151 2550 26181
rect 2613 26151 2620 26181
rect 2686 26151 2725 26185
rect 2759 26151 2798 26185
rect 2832 26151 2871 26185
rect 2905 26151 2944 26185
rect 2978 26151 3017 26185
rect 3051 26151 3090 26185
rect 3124 26151 3163 26185
rect 3197 26151 3236 26185
rect 3270 26151 3309 26185
rect 3343 26151 3382 26185
rect 3416 26151 3455 26185
rect 3489 26181 3528 26185
rect 3562 26181 3601 26185
rect 3635 26181 3674 26185
rect 3524 26151 3528 26181
rect 3594 26151 3601 26181
rect 3664 26151 3674 26181
rect 3708 26151 3746 26185
rect 3780 26151 3818 26185
rect 3852 26151 3890 26185
rect 3924 26151 3962 26185
rect 3996 26151 4034 26185
rect 4068 26151 4106 26185
rect 4140 26151 4178 26185
rect 4212 26151 4250 26185
rect 4284 26151 4322 26185
rect 4356 26151 4394 26185
rect 4428 26181 4466 26185
rect 4500 26181 4538 26185
rect 4572 26181 4610 26185
rect 4644 26181 4682 26185
rect 4428 26151 4464 26181
rect 231 26129 2480 26151
rect 2532 26129 2550 26151
rect 2602 26129 2620 26151
rect 2672 26129 3472 26151
rect 3524 26129 3542 26151
rect 3594 26129 3612 26151
rect 3664 26129 4464 26151
rect 4516 26129 4534 26181
rect 4586 26129 4604 26181
rect 4656 26151 4682 26181
rect 4716 26151 4754 26185
rect 4788 26151 4826 26185
rect 4860 26151 4898 26185
rect 4932 26151 4970 26185
rect 5004 26151 5042 26185
rect 5076 26151 5114 26185
rect 5148 26151 5186 26185
rect 5220 26151 5258 26185
rect 5292 26151 5330 26185
rect 5364 26151 5402 26185
rect 5436 26181 5474 26185
rect 5508 26181 5546 26185
rect 5580 26181 5618 26185
rect 5436 26151 5456 26181
rect 4656 26129 5456 26151
rect 5508 26129 5526 26181
rect 5580 26151 5596 26181
rect 5652 26151 5690 26185
rect 5724 26151 5762 26185
rect 5796 26151 5834 26185
rect 5868 26151 5906 26185
rect 5940 26151 5978 26185
rect 6012 26151 6050 26185
rect 6084 26151 6122 26185
rect 6156 26151 6194 26185
rect 6228 26151 6266 26185
rect 6300 26151 6338 26185
rect 6372 26151 6410 26185
rect 6444 26181 6482 26185
rect 6516 26181 6554 26185
rect 6588 26181 6626 26185
rect 6444 26151 6448 26181
rect 6516 26151 6518 26181
rect 6660 26151 6698 26185
rect 6732 26151 6770 26185
rect 6804 26151 6842 26185
rect 6876 26151 6914 26185
rect 6948 26151 6986 26185
rect 7020 26151 7058 26185
rect 7092 26151 7130 26185
rect 7164 26151 7202 26185
rect 7236 26151 7274 26185
rect 7308 26151 7346 26185
rect 7380 26151 7418 26185
rect 7452 26181 7490 26185
rect 7524 26181 7562 26185
rect 7596 26181 7634 26185
rect 7632 26151 7634 26181
rect 7668 26151 7706 26185
rect 7740 26151 7778 26185
rect 7812 26151 7850 26185
rect 7884 26151 7922 26185
rect 7956 26151 7994 26185
rect 8028 26151 8066 26185
rect 8100 26151 8138 26185
rect 8172 26151 8210 26185
rect 8244 26151 8282 26185
rect 8316 26151 8354 26185
rect 8388 26151 8426 26185
rect 8460 26181 8498 26185
rect 8532 26181 8570 26185
rect 8604 26181 8642 26185
rect 8484 26151 8498 26181
rect 8554 26151 8570 26181
rect 8624 26151 8642 26181
rect 8676 26151 8714 26185
rect 8748 26151 8786 26185
rect 8820 26151 8858 26185
rect 8892 26151 8930 26185
rect 8964 26151 9002 26185
rect 9036 26151 9074 26185
rect 9108 26151 9146 26185
rect 9180 26151 9218 26185
rect 9252 26151 9290 26185
rect 9324 26151 9362 26185
rect 9396 26181 9434 26185
rect 9468 26181 9506 26185
rect 9540 26181 9578 26185
rect 9612 26181 9650 26185
rect 9396 26151 9424 26181
rect 5578 26129 5596 26151
rect 5648 26129 6448 26151
rect 6500 26129 6518 26151
rect 6570 26129 6588 26151
rect 6640 26129 7440 26151
rect 7492 26129 7510 26151
rect 7562 26129 7580 26151
rect 7632 26129 8432 26151
rect 8484 26129 8502 26151
rect 8554 26129 8572 26151
rect 8624 26129 9424 26151
rect 9476 26129 9494 26181
rect 9546 26129 9564 26181
rect 9616 26151 9650 26181
rect 9684 26151 9722 26185
rect 9756 26151 9794 26185
rect 9828 26151 9866 26185
rect 9900 26151 9938 26185
rect 9972 26151 10010 26185
rect 10044 26151 10082 26185
rect 10116 26151 10154 26185
rect 10188 26151 10226 26185
rect 10260 26151 10298 26185
rect 10332 26151 10370 26185
rect 10404 26151 10442 26185
rect 10476 26151 10514 26185
rect 10548 26151 10586 26185
rect 10620 26151 10658 26185
rect 10692 26151 10730 26185
rect 10764 26151 10802 26185
rect 10836 26151 10874 26185
rect 10908 26151 10946 26185
rect 10980 26151 11018 26185
rect 11052 26151 11090 26185
rect 11124 26151 11162 26185
rect 11196 26151 11234 26185
rect 11268 26151 11306 26185
rect 11340 26151 11378 26185
rect 11412 26151 11450 26185
rect 11484 26151 11522 26185
rect 11556 26151 11594 26185
rect 11628 26151 11666 26185
rect 11700 26151 11738 26185
rect 11772 26151 11810 26185
rect 11844 26151 11882 26185
rect 11916 26151 11954 26185
rect 11988 26151 12026 26185
rect 12060 26151 12098 26185
rect 12132 26151 12170 26185
rect 12204 26151 12242 26185
rect 12276 26151 12314 26185
rect 12348 26151 12386 26185
rect 12420 26151 12458 26185
rect 12492 26151 12530 26185
rect 12564 26151 12602 26185
rect 12636 26151 12674 26185
rect 12708 26151 12746 26185
rect 12780 26151 12818 26185
rect 12852 26151 12890 26185
rect 12924 26151 12962 26185
rect 12996 26151 13034 26185
rect 13068 26151 13106 26185
rect 13140 26151 13178 26185
rect 13212 26151 13250 26185
rect 13284 26151 13322 26185
rect 13356 26151 13394 26185
rect 13428 26151 13466 26185
rect 13500 26151 13538 26185
rect 13572 26151 13610 26185
rect 13644 26151 13682 26185
rect 13716 26151 13754 26185
rect 13788 26151 13826 26185
rect 13860 26151 13898 26185
rect 13932 26151 13970 26185
rect 14004 26151 14042 26185
rect 14076 26151 14114 26185
rect 14148 26151 14186 26185
rect 14220 26151 14258 26185
rect 14292 26151 14330 26185
rect 14364 26151 14402 26185
rect 14436 26151 14474 26185
rect 14508 26151 14546 26185
rect 14580 26151 14618 26185
rect 14652 26151 14690 26185
rect 14724 26151 14736 26185
rect 9616 26129 14736 26151
rect 231 26111 14736 26129
rect 231 26077 243 26111
rect 277 26077 316 26111
rect 350 26077 389 26111
rect 423 26077 462 26111
rect 496 26077 535 26111
rect 569 26077 608 26111
rect 642 26077 681 26111
rect 715 26077 754 26111
rect 788 26077 827 26111
rect 861 26077 900 26111
rect 934 26077 973 26111
rect 1007 26077 1046 26111
rect 1080 26077 1119 26111
rect 1153 26077 1192 26111
rect 1226 26077 1265 26111
rect 1299 26077 1338 26111
rect 1372 26077 1411 26111
rect 1445 26077 1484 26111
rect 1518 26077 1557 26111
rect 1591 26077 1630 26111
rect 1664 26077 1703 26111
rect 1737 26077 1776 26111
rect 1810 26077 1849 26111
rect 1883 26077 1922 26111
rect 1956 26077 1995 26111
rect 2029 26077 2068 26111
rect 2102 26077 2141 26111
rect 2175 26077 2214 26111
rect 2248 26077 2287 26111
rect 2321 26077 2360 26111
rect 2394 26077 2433 26111
rect 2467 26077 2480 26111
rect 2540 26077 2550 26111
rect 2613 26077 2620 26111
rect 2686 26077 2725 26111
rect 2759 26077 2798 26111
rect 2832 26077 2871 26111
rect 2905 26077 2944 26111
rect 2978 26077 3017 26111
rect 3051 26077 3090 26111
rect 3124 26077 3163 26111
rect 3197 26077 3236 26111
rect 3270 26077 3309 26111
rect 3343 26077 3382 26111
rect 3416 26077 3455 26111
rect 3524 26077 3528 26111
rect 3594 26077 3601 26111
rect 3664 26077 3674 26111
rect 3708 26077 3746 26111
rect 3780 26077 3818 26111
rect 3852 26077 3890 26111
rect 3924 26077 3962 26111
rect 3996 26077 4034 26111
rect 4068 26077 4106 26111
rect 4140 26077 4178 26111
rect 4212 26077 4250 26111
rect 4284 26077 4322 26111
rect 4356 26077 4394 26111
rect 4428 26077 4464 26111
rect 231 26059 2480 26077
rect 2532 26059 2550 26077
rect 2602 26059 2620 26077
rect 2672 26059 3472 26077
rect 3524 26059 3542 26077
rect 3594 26059 3612 26077
rect 3664 26059 4464 26077
rect 4516 26059 4534 26111
rect 4586 26059 4604 26111
rect 4656 26077 4682 26111
rect 4716 26077 4754 26111
rect 4788 26077 4826 26111
rect 4860 26077 4898 26111
rect 4932 26077 4970 26111
rect 5004 26077 5042 26111
rect 5076 26077 5114 26111
rect 5148 26077 5186 26111
rect 5220 26077 5258 26111
rect 5292 26077 5330 26111
rect 5364 26077 5402 26111
rect 5436 26077 5456 26111
rect 4656 26059 5456 26077
rect 5508 26059 5526 26111
rect 5580 26077 5596 26111
rect 5652 26077 5690 26111
rect 5724 26077 5762 26111
rect 5796 26077 5834 26111
rect 5868 26077 5906 26111
rect 5940 26077 5978 26111
rect 6012 26077 6050 26111
rect 6084 26077 6122 26111
rect 6156 26077 6194 26111
rect 6228 26077 6266 26111
rect 6300 26077 6338 26111
rect 6372 26077 6410 26111
rect 6444 26077 6448 26111
rect 6516 26077 6518 26111
rect 6660 26077 6698 26111
rect 6732 26077 6770 26111
rect 6804 26077 6842 26111
rect 6876 26077 6914 26111
rect 6948 26077 6986 26111
rect 7020 26077 7058 26111
rect 7092 26077 7130 26111
rect 7164 26077 7202 26111
rect 7236 26077 7274 26111
rect 7308 26077 7346 26111
rect 7380 26077 7418 26111
rect 7632 26077 7634 26111
rect 7668 26077 7706 26111
rect 7740 26077 7778 26111
rect 7812 26077 7850 26111
rect 7884 26077 7922 26111
rect 7956 26077 7994 26111
rect 8028 26077 8066 26111
rect 8100 26077 8138 26111
rect 8172 26077 8210 26111
rect 8244 26077 8282 26111
rect 8316 26077 8354 26111
rect 8388 26077 8426 26111
rect 8484 26077 8498 26111
rect 8554 26077 8570 26111
rect 8624 26077 8642 26111
rect 8676 26077 8714 26111
rect 8748 26077 8786 26111
rect 8820 26077 8858 26111
rect 8892 26077 8930 26111
rect 8964 26077 9002 26111
rect 9036 26077 9074 26111
rect 9108 26077 9146 26111
rect 9180 26077 9218 26111
rect 9252 26077 9290 26111
rect 9324 26077 9362 26111
rect 9396 26077 9424 26111
rect 5578 26059 5596 26077
rect 5648 26059 6448 26077
rect 6500 26059 6518 26077
rect 6570 26059 6588 26077
rect 6640 26059 7440 26077
rect 7492 26059 7510 26077
rect 7562 26059 7580 26077
rect 7632 26059 8432 26077
rect 8484 26059 8502 26077
rect 8554 26059 8572 26077
rect 8624 26059 9424 26077
rect 9476 26059 9494 26111
rect 9546 26059 9564 26111
rect 9616 26077 9650 26111
rect 9684 26077 9722 26111
rect 9756 26077 9794 26111
rect 9828 26077 9866 26111
rect 9900 26077 9938 26111
rect 9972 26077 10010 26111
rect 10044 26077 10082 26111
rect 10116 26077 10154 26111
rect 10188 26077 10226 26111
rect 10260 26077 10298 26111
rect 10332 26077 10370 26111
rect 10404 26077 10442 26111
rect 10476 26077 10514 26111
rect 10548 26077 10586 26111
rect 10620 26077 10658 26111
rect 10692 26077 10730 26111
rect 10764 26077 10802 26111
rect 10836 26077 10874 26111
rect 10908 26077 10946 26111
rect 10980 26077 11018 26111
rect 11052 26077 11090 26111
rect 11124 26077 11162 26111
rect 11196 26077 11234 26111
rect 11268 26077 11306 26111
rect 11340 26077 11378 26111
rect 11412 26077 11450 26111
rect 11484 26077 11522 26111
rect 11556 26077 11594 26111
rect 11628 26077 11666 26111
rect 11700 26077 11738 26111
rect 11772 26077 11810 26111
rect 11844 26077 11882 26111
rect 11916 26077 11954 26111
rect 11988 26077 12026 26111
rect 12060 26077 12098 26111
rect 12132 26077 12170 26111
rect 12204 26077 12242 26111
rect 12276 26077 12314 26111
rect 12348 26077 12386 26111
rect 12420 26077 12458 26111
rect 12492 26077 12530 26111
rect 12564 26077 12602 26111
rect 12636 26077 12674 26111
rect 12708 26077 12746 26111
rect 12780 26077 12818 26111
rect 12852 26077 12890 26111
rect 12924 26077 12962 26111
rect 12996 26077 13034 26111
rect 13068 26077 13106 26111
rect 13140 26077 13178 26111
rect 13212 26077 13250 26111
rect 13284 26077 13322 26111
rect 13356 26077 13394 26111
rect 13428 26077 13466 26111
rect 13500 26077 13538 26111
rect 13572 26077 13610 26111
rect 13644 26077 13682 26111
rect 13716 26077 13754 26111
rect 13788 26077 13826 26111
rect 13860 26077 13898 26111
rect 13932 26077 13970 26111
rect 14004 26077 14042 26111
rect 14076 26077 14114 26111
rect 14148 26077 14186 26111
rect 14220 26077 14258 26111
rect 14292 26077 14330 26111
rect 14364 26077 14402 26111
rect 14436 26077 14474 26111
rect 14508 26077 14546 26111
rect 14580 26077 14618 26111
rect 14652 26077 14690 26111
rect 14724 26077 14736 26111
rect 9616 26059 14736 26077
rect 231 26041 14736 26059
rect 231 26037 2480 26041
rect 2532 26037 2550 26041
rect 2602 26037 2620 26041
rect 2672 26037 3472 26041
rect 3524 26037 3542 26041
rect 3594 26037 3612 26041
rect 3664 26037 4464 26041
rect 231 26003 243 26037
rect 277 26003 316 26037
rect 350 26003 389 26037
rect 423 26003 462 26037
rect 496 26003 535 26037
rect 569 26003 608 26037
rect 642 26003 681 26037
rect 715 26003 754 26037
rect 788 26003 827 26037
rect 861 26003 900 26037
rect 934 26003 973 26037
rect 1007 26003 1046 26037
rect 1080 26003 1119 26037
rect 1153 26003 1192 26037
rect 1226 26003 1265 26037
rect 1299 26003 1338 26037
rect 1372 26003 1411 26037
rect 1445 26003 1484 26037
rect 1518 26003 1557 26037
rect 1591 26003 1630 26037
rect 1664 26003 1703 26037
rect 1737 26003 1776 26037
rect 1810 26003 1849 26037
rect 1883 26003 1922 26037
rect 1956 26003 1995 26037
rect 2029 26003 2068 26037
rect 2102 26003 2141 26037
rect 2175 26003 2214 26037
rect 2248 26003 2287 26037
rect 2321 26003 2360 26037
rect 2394 26003 2433 26037
rect 2467 26003 2480 26037
rect 2540 26003 2550 26037
rect 2613 26003 2620 26037
rect 2686 26003 2725 26037
rect 2759 26003 2798 26037
rect 2832 26003 2871 26037
rect 2905 26003 2944 26037
rect 2978 26003 3017 26037
rect 3051 26003 3090 26037
rect 3124 26003 3163 26037
rect 3197 26003 3236 26037
rect 3270 26003 3309 26037
rect 3343 26003 3382 26037
rect 3416 26003 3455 26037
rect 3524 26003 3528 26037
rect 3594 26003 3601 26037
rect 3664 26003 3674 26037
rect 3708 26003 3746 26037
rect 3780 26003 3818 26037
rect 3852 26003 3890 26037
rect 3924 26003 3962 26037
rect 3996 26003 4034 26037
rect 4068 26003 4106 26037
rect 4140 26003 4178 26037
rect 4212 26003 4250 26037
rect 4284 26003 4322 26037
rect 4356 26003 4394 26037
rect 4428 26003 4464 26037
rect 231 25989 2480 26003
rect 2532 25989 2550 26003
rect 2602 25989 2620 26003
rect 2672 25989 3472 26003
rect 3524 25989 3542 26003
rect 3594 25989 3612 26003
rect 3664 25989 4464 26003
rect 4516 25989 4534 26041
rect 4586 25989 4604 26041
rect 4656 26037 5456 26041
rect 4656 26003 4682 26037
rect 4716 26003 4754 26037
rect 4788 26003 4826 26037
rect 4860 26003 4898 26037
rect 4932 26003 4970 26037
rect 5004 26003 5042 26037
rect 5076 26003 5114 26037
rect 5148 26003 5186 26037
rect 5220 26003 5258 26037
rect 5292 26003 5330 26037
rect 5364 26003 5402 26037
rect 5436 26003 5456 26037
rect 4656 25989 5456 26003
rect 5508 25989 5526 26041
rect 5578 26037 5596 26041
rect 5648 26037 6448 26041
rect 6500 26037 6518 26041
rect 6570 26037 6588 26041
rect 6640 26037 7440 26041
rect 7492 26037 7510 26041
rect 7562 26037 7580 26041
rect 7632 26037 8432 26041
rect 8484 26037 8502 26041
rect 8554 26037 8572 26041
rect 8624 26037 9424 26041
rect 5580 26003 5596 26037
rect 5652 26003 5690 26037
rect 5724 26003 5762 26037
rect 5796 26003 5834 26037
rect 5868 26003 5906 26037
rect 5940 26003 5978 26037
rect 6012 26003 6050 26037
rect 6084 26003 6122 26037
rect 6156 26003 6194 26037
rect 6228 26003 6266 26037
rect 6300 26003 6338 26037
rect 6372 26003 6410 26037
rect 6444 26003 6448 26037
rect 6516 26003 6518 26037
rect 6660 26003 6698 26037
rect 6732 26003 6770 26037
rect 6804 26003 6842 26037
rect 6876 26003 6914 26037
rect 6948 26003 6986 26037
rect 7020 26003 7058 26037
rect 7092 26003 7130 26037
rect 7164 26003 7202 26037
rect 7236 26003 7274 26037
rect 7308 26003 7346 26037
rect 7380 26003 7418 26037
rect 7632 26003 7634 26037
rect 7668 26003 7706 26037
rect 7740 26003 7778 26037
rect 7812 26003 7850 26037
rect 7884 26003 7922 26037
rect 7956 26003 7994 26037
rect 8028 26003 8066 26037
rect 8100 26003 8138 26037
rect 8172 26003 8210 26037
rect 8244 26003 8282 26037
rect 8316 26003 8354 26037
rect 8388 26003 8426 26037
rect 8484 26003 8498 26037
rect 8554 26003 8570 26037
rect 8624 26003 8642 26037
rect 8676 26003 8714 26037
rect 8748 26003 8786 26037
rect 8820 26003 8858 26037
rect 8892 26003 8930 26037
rect 8964 26003 9002 26037
rect 9036 26003 9074 26037
rect 9108 26003 9146 26037
rect 9180 26003 9218 26037
rect 9252 26003 9290 26037
rect 9324 26003 9362 26037
rect 9396 26003 9424 26037
rect 5578 25989 5596 26003
rect 5648 25989 6448 26003
rect 6500 25989 6518 26003
rect 6570 25989 6588 26003
rect 6640 25989 7440 26003
rect 7492 25989 7510 26003
rect 7562 25989 7580 26003
rect 7632 25989 8432 26003
rect 8484 25989 8502 26003
rect 8554 25989 8572 26003
rect 8624 25989 9424 26003
rect 9476 25989 9494 26041
rect 9546 25989 9564 26041
rect 9616 26037 14736 26041
rect 9616 26003 9650 26037
rect 9684 26003 9722 26037
rect 9756 26003 9794 26037
rect 9828 26003 9866 26037
rect 9900 26003 9938 26037
rect 9972 26003 10010 26037
rect 10044 26003 10082 26037
rect 10116 26003 10154 26037
rect 10188 26003 10226 26037
rect 10260 26003 10298 26037
rect 10332 26003 10370 26037
rect 10404 26003 10442 26037
rect 10476 26003 10514 26037
rect 10548 26003 10586 26037
rect 10620 26003 10658 26037
rect 10692 26003 10730 26037
rect 10764 26003 10802 26037
rect 10836 26003 10874 26037
rect 10908 26003 10946 26037
rect 10980 26003 11018 26037
rect 11052 26003 11090 26037
rect 11124 26003 11162 26037
rect 11196 26003 11234 26037
rect 11268 26003 11306 26037
rect 11340 26003 11378 26037
rect 11412 26003 11450 26037
rect 11484 26003 11522 26037
rect 11556 26003 11594 26037
rect 11628 26003 11666 26037
rect 11700 26003 11738 26037
rect 11772 26003 11810 26037
rect 11844 26003 11882 26037
rect 11916 26003 11954 26037
rect 11988 26003 12026 26037
rect 12060 26003 12098 26037
rect 12132 26003 12170 26037
rect 12204 26003 12242 26037
rect 12276 26003 12314 26037
rect 12348 26003 12386 26037
rect 12420 26003 12458 26037
rect 12492 26003 12530 26037
rect 12564 26003 12602 26037
rect 12636 26003 12674 26037
rect 12708 26003 12746 26037
rect 12780 26003 12818 26037
rect 12852 26003 12890 26037
rect 12924 26003 12962 26037
rect 12996 26003 13034 26037
rect 13068 26003 13106 26037
rect 13140 26003 13178 26037
rect 13212 26003 13250 26037
rect 13284 26003 13322 26037
rect 13356 26003 13394 26037
rect 13428 26003 13466 26037
rect 13500 26003 13538 26037
rect 13572 26003 13610 26037
rect 13644 26003 13682 26037
rect 13716 26003 13754 26037
rect 13788 26003 13826 26037
rect 13860 26003 13898 26037
rect 13932 26003 13970 26037
rect 14004 26003 14042 26037
rect 14076 26003 14114 26037
rect 14148 26003 14186 26037
rect 14220 26003 14258 26037
rect 14292 26003 14330 26037
rect 14364 26003 14402 26037
rect 14436 26003 14474 26037
rect 14508 26003 14546 26037
rect 14580 26003 14618 26037
rect 14652 26003 14690 26037
rect 14724 26003 14736 26037
rect 9616 25989 14736 26003
rect 231 25971 14736 25989
rect 231 25963 2480 25971
rect 2532 25963 2550 25971
rect 2602 25963 2620 25971
rect 2672 25963 3472 25971
rect 3524 25963 3542 25971
rect 3594 25963 3612 25971
rect 3664 25963 4464 25971
rect 231 25929 243 25963
rect 277 25929 316 25963
rect 350 25929 389 25963
rect 423 25929 462 25963
rect 496 25929 535 25963
rect 569 25929 608 25963
rect 642 25929 681 25963
rect 715 25929 754 25963
rect 788 25929 827 25963
rect 861 25929 900 25963
rect 934 25929 973 25963
rect 1007 25929 1046 25963
rect 1080 25929 1119 25963
rect 1153 25929 1192 25963
rect 1226 25929 1265 25963
rect 1299 25929 1338 25963
rect 1372 25929 1411 25963
rect 1445 25929 1484 25963
rect 1518 25929 1557 25963
rect 1591 25929 1630 25963
rect 1664 25929 1703 25963
rect 1737 25929 1776 25963
rect 1810 25929 1849 25963
rect 1883 25929 1922 25963
rect 1956 25929 1995 25963
rect 2029 25929 2068 25963
rect 2102 25929 2141 25963
rect 2175 25929 2214 25963
rect 2248 25929 2287 25963
rect 2321 25929 2360 25963
rect 2394 25929 2433 25963
rect 2467 25929 2480 25963
rect 2540 25929 2550 25963
rect 2613 25929 2620 25963
rect 2686 25929 2725 25963
rect 2759 25929 2798 25963
rect 2832 25929 2871 25963
rect 2905 25929 2944 25963
rect 2978 25929 3017 25963
rect 3051 25929 3090 25963
rect 3124 25929 3163 25963
rect 3197 25929 3236 25963
rect 3270 25929 3309 25963
rect 3343 25929 3382 25963
rect 3416 25929 3455 25963
rect 3524 25929 3528 25963
rect 3594 25929 3601 25963
rect 3664 25929 3674 25963
rect 3708 25929 3746 25963
rect 3780 25929 3818 25963
rect 3852 25929 3890 25963
rect 3924 25929 3962 25963
rect 3996 25929 4034 25963
rect 4068 25929 4106 25963
rect 4140 25929 4178 25963
rect 4212 25929 4250 25963
rect 4284 25929 4322 25963
rect 4356 25929 4394 25963
rect 4428 25929 4464 25963
rect 231 25919 2480 25929
rect 2532 25919 2550 25929
rect 2602 25919 2620 25929
rect 2672 25919 3472 25929
rect 3524 25919 3542 25929
rect 3594 25919 3612 25929
rect 3664 25919 4464 25929
rect 4516 25919 4534 25971
rect 4586 25919 4604 25971
rect 4656 25963 5456 25971
rect 4656 25929 4682 25963
rect 4716 25929 4754 25963
rect 4788 25929 4826 25963
rect 4860 25929 4898 25963
rect 4932 25929 4970 25963
rect 5004 25929 5042 25963
rect 5076 25929 5114 25963
rect 5148 25929 5186 25963
rect 5220 25929 5258 25963
rect 5292 25929 5330 25963
rect 5364 25929 5402 25963
rect 5436 25929 5456 25963
rect 4656 25919 5456 25929
rect 5508 25919 5526 25971
rect 5578 25963 5596 25971
rect 5648 25963 6448 25971
rect 6500 25963 6518 25971
rect 6570 25963 6588 25971
rect 6640 25963 7440 25971
rect 7492 25963 7510 25971
rect 7562 25963 7580 25971
rect 7632 25963 8432 25971
rect 8484 25963 8502 25971
rect 8554 25963 8572 25971
rect 8624 25963 9424 25971
rect 5580 25929 5596 25963
rect 5652 25929 5690 25963
rect 5724 25929 5762 25963
rect 5796 25929 5834 25963
rect 5868 25929 5906 25963
rect 5940 25929 5978 25963
rect 6012 25929 6050 25963
rect 6084 25929 6122 25963
rect 6156 25929 6194 25963
rect 6228 25929 6266 25963
rect 6300 25929 6338 25963
rect 6372 25929 6410 25963
rect 6444 25929 6448 25963
rect 6516 25929 6518 25963
rect 6660 25929 6698 25963
rect 6732 25929 6770 25963
rect 6804 25929 6842 25963
rect 6876 25929 6914 25963
rect 6948 25929 6986 25963
rect 7020 25929 7058 25963
rect 7092 25929 7130 25963
rect 7164 25929 7202 25963
rect 7236 25929 7274 25963
rect 7308 25929 7346 25963
rect 7380 25929 7418 25963
rect 7632 25929 7634 25963
rect 7668 25929 7706 25963
rect 7740 25929 7778 25963
rect 7812 25929 7850 25963
rect 7884 25929 7922 25963
rect 7956 25929 7994 25963
rect 8028 25929 8066 25963
rect 8100 25929 8138 25963
rect 8172 25929 8210 25963
rect 8244 25929 8282 25963
rect 8316 25929 8354 25963
rect 8388 25929 8426 25963
rect 8484 25929 8498 25963
rect 8554 25929 8570 25963
rect 8624 25929 8642 25963
rect 8676 25929 8714 25963
rect 8748 25929 8786 25963
rect 8820 25929 8858 25963
rect 8892 25929 8930 25963
rect 8964 25929 9002 25963
rect 9036 25929 9074 25963
rect 9108 25929 9146 25963
rect 9180 25929 9218 25963
rect 9252 25929 9290 25963
rect 9324 25929 9362 25963
rect 9396 25929 9424 25963
rect 5578 25919 5596 25929
rect 5648 25919 6448 25929
rect 6500 25919 6518 25929
rect 6570 25919 6588 25929
rect 6640 25919 7440 25929
rect 7492 25919 7510 25929
rect 7562 25919 7580 25929
rect 7632 25919 8432 25929
rect 8484 25919 8502 25929
rect 8554 25919 8572 25929
rect 8624 25919 9424 25929
rect 9476 25919 9494 25971
rect 9546 25919 9564 25971
rect 9616 25963 14736 25971
rect 9616 25929 9650 25963
rect 9684 25929 9722 25963
rect 9756 25929 9794 25963
rect 9828 25929 9866 25963
rect 9900 25929 9938 25963
rect 9972 25929 10010 25963
rect 10044 25929 10082 25963
rect 10116 25929 10154 25963
rect 10188 25929 10226 25963
rect 10260 25929 10298 25963
rect 10332 25929 10370 25963
rect 10404 25929 10442 25963
rect 10476 25929 10514 25963
rect 10548 25929 10586 25963
rect 10620 25929 10658 25963
rect 10692 25929 10730 25963
rect 10764 25929 10802 25963
rect 10836 25929 10874 25963
rect 10908 25929 10946 25963
rect 10980 25929 11018 25963
rect 11052 25929 11090 25963
rect 11124 25929 11162 25963
rect 11196 25929 11234 25963
rect 11268 25929 11306 25963
rect 11340 25929 11378 25963
rect 11412 25929 11450 25963
rect 11484 25929 11522 25963
rect 11556 25929 11594 25963
rect 11628 25929 11666 25963
rect 11700 25929 11738 25963
rect 11772 25929 11810 25963
rect 11844 25929 11882 25963
rect 11916 25929 11954 25963
rect 11988 25929 12026 25963
rect 12060 25929 12098 25963
rect 12132 25929 12170 25963
rect 12204 25929 12242 25963
rect 12276 25929 12314 25963
rect 12348 25929 12386 25963
rect 12420 25929 12458 25963
rect 12492 25929 12530 25963
rect 12564 25929 12602 25963
rect 12636 25929 12674 25963
rect 12708 25929 12746 25963
rect 12780 25929 12818 25963
rect 12852 25929 12890 25963
rect 12924 25929 12962 25963
rect 12996 25929 13034 25963
rect 13068 25929 13106 25963
rect 13140 25929 13178 25963
rect 13212 25929 13250 25963
rect 13284 25929 13322 25963
rect 13356 25929 13394 25963
rect 13428 25929 13466 25963
rect 13500 25929 13538 25963
rect 13572 25929 13610 25963
rect 13644 25929 13682 25963
rect 13716 25929 13754 25963
rect 13788 25929 13826 25963
rect 13860 25929 13898 25963
rect 13932 25929 13970 25963
rect 14004 25929 14042 25963
rect 14076 25929 14114 25963
rect 14148 25929 14186 25963
rect 14220 25929 14258 25963
rect 14292 25929 14330 25963
rect 14364 25929 14402 25963
rect 14436 25929 14474 25963
rect 14508 25929 14546 25963
rect 14580 25929 14618 25963
rect 14652 25929 14690 25963
rect 14724 25929 14736 25963
rect 9616 25919 14736 25929
rect 231 25901 14736 25919
rect 231 25889 2480 25901
rect 2532 25889 2550 25901
rect 2602 25889 2620 25901
rect 2672 25889 3472 25901
rect 3524 25889 3542 25901
rect 3594 25889 3612 25901
rect 3664 25889 4464 25901
rect 231 25855 243 25889
rect 277 25855 316 25889
rect 350 25855 389 25889
rect 423 25855 462 25889
rect 496 25855 535 25889
rect 569 25855 608 25889
rect 642 25855 681 25889
rect 715 25855 754 25889
rect 788 25855 827 25889
rect 861 25855 900 25889
rect 934 25855 973 25889
rect 1007 25855 1046 25889
rect 1080 25855 1119 25889
rect 1153 25855 1192 25889
rect 1226 25855 1265 25889
rect 1299 25855 1338 25889
rect 1372 25855 1411 25889
rect 1445 25855 1484 25889
rect 1518 25855 1557 25889
rect 1591 25855 1630 25889
rect 1664 25855 1703 25889
rect 1737 25855 1776 25889
rect 1810 25855 1849 25889
rect 1883 25855 1922 25889
rect 1956 25855 1995 25889
rect 2029 25855 2068 25889
rect 2102 25855 2141 25889
rect 2175 25855 2214 25889
rect 2248 25855 2287 25889
rect 2321 25855 2360 25889
rect 2394 25855 2433 25889
rect 2467 25855 2480 25889
rect 2540 25855 2550 25889
rect 2613 25855 2620 25889
rect 2686 25855 2725 25889
rect 2759 25855 2798 25889
rect 2832 25855 2871 25889
rect 2905 25855 2944 25889
rect 2978 25855 3017 25889
rect 3051 25855 3090 25889
rect 3124 25855 3163 25889
rect 3197 25855 3236 25889
rect 3270 25855 3309 25889
rect 3343 25855 3382 25889
rect 3416 25855 3455 25889
rect 3524 25855 3528 25889
rect 3594 25855 3601 25889
rect 3664 25855 3674 25889
rect 3708 25855 3746 25889
rect 3780 25855 3818 25889
rect 3852 25855 3890 25889
rect 3924 25855 3962 25889
rect 3996 25855 4034 25889
rect 4068 25855 4106 25889
rect 4140 25855 4178 25889
rect 4212 25855 4250 25889
rect 4284 25855 4322 25889
rect 4356 25855 4394 25889
rect 4428 25855 4464 25889
rect 231 25849 2480 25855
rect 2532 25849 2550 25855
rect 2602 25849 2620 25855
rect 2672 25849 3472 25855
rect 3524 25849 3542 25855
rect 3594 25849 3612 25855
rect 3664 25849 4464 25855
rect 4516 25849 4534 25901
rect 4586 25849 4604 25901
rect 4656 25889 5456 25901
rect 4656 25855 4682 25889
rect 4716 25855 4754 25889
rect 4788 25855 4826 25889
rect 4860 25855 4898 25889
rect 4932 25855 4970 25889
rect 5004 25855 5042 25889
rect 5076 25855 5114 25889
rect 5148 25855 5186 25889
rect 5220 25855 5258 25889
rect 5292 25855 5330 25889
rect 5364 25855 5402 25889
rect 5436 25855 5456 25889
rect 4656 25849 5456 25855
rect 5508 25849 5526 25901
rect 5578 25889 5596 25901
rect 5648 25889 6448 25901
rect 6500 25889 6518 25901
rect 6570 25889 6588 25901
rect 6640 25889 7440 25901
rect 7492 25889 7510 25901
rect 7562 25889 7580 25901
rect 7632 25889 8432 25901
rect 8484 25889 8502 25901
rect 8554 25889 8572 25901
rect 8624 25889 9424 25901
rect 5580 25855 5596 25889
rect 5652 25855 5690 25889
rect 5724 25855 5762 25889
rect 5796 25855 5834 25889
rect 5868 25855 5906 25889
rect 5940 25855 5978 25889
rect 6012 25855 6050 25889
rect 6084 25855 6122 25889
rect 6156 25855 6194 25889
rect 6228 25855 6266 25889
rect 6300 25855 6338 25889
rect 6372 25855 6410 25889
rect 6444 25855 6448 25889
rect 6516 25855 6518 25889
rect 6660 25855 6698 25889
rect 6732 25855 6770 25889
rect 6804 25855 6842 25889
rect 6876 25855 6914 25889
rect 6948 25855 6986 25889
rect 7020 25855 7058 25889
rect 7092 25855 7130 25889
rect 7164 25855 7202 25889
rect 7236 25855 7274 25889
rect 7308 25855 7346 25889
rect 7380 25855 7418 25889
rect 7632 25855 7634 25889
rect 7668 25855 7706 25889
rect 7740 25855 7778 25889
rect 7812 25855 7850 25889
rect 7884 25855 7922 25889
rect 7956 25855 7994 25889
rect 8028 25855 8066 25889
rect 8100 25855 8138 25889
rect 8172 25855 8210 25889
rect 8244 25855 8282 25889
rect 8316 25855 8354 25889
rect 8388 25855 8426 25889
rect 8484 25855 8498 25889
rect 8554 25855 8570 25889
rect 8624 25855 8642 25889
rect 8676 25855 8714 25889
rect 8748 25855 8786 25889
rect 8820 25855 8858 25889
rect 8892 25855 8930 25889
rect 8964 25855 9002 25889
rect 9036 25855 9074 25889
rect 9108 25855 9146 25889
rect 9180 25855 9218 25889
rect 9252 25855 9290 25889
rect 9324 25855 9362 25889
rect 9396 25855 9424 25889
rect 5578 25849 5596 25855
rect 5648 25849 6448 25855
rect 6500 25849 6518 25855
rect 6570 25849 6588 25855
rect 6640 25849 7440 25855
rect 7492 25849 7510 25855
rect 7562 25849 7580 25855
rect 7632 25849 8432 25855
rect 8484 25849 8502 25855
rect 8554 25849 8572 25855
rect 8624 25849 9424 25855
rect 9476 25849 9494 25901
rect 9546 25849 9564 25901
rect 9616 25889 14736 25901
rect 9616 25855 9650 25889
rect 9684 25855 9722 25889
rect 9756 25855 9794 25889
rect 9828 25855 9866 25889
rect 9900 25855 9938 25889
rect 9972 25855 10010 25889
rect 10044 25855 10082 25889
rect 10116 25855 10154 25889
rect 10188 25855 10226 25889
rect 10260 25855 10298 25889
rect 10332 25855 10370 25889
rect 10404 25855 10442 25889
rect 10476 25855 10514 25889
rect 10548 25855 10586 25889
rect 10620 25855 10658 25889
rect 10692 25855 10730 25889
rect 10764 25855 10802 25889
rect 10836 25855 10874 25889
rect 10908 25855 10946 25889
rect 10980 25855 11018 25889
rect 11052 25855 11090 25889
rect 11124 25855 11162 25889
rect 11196 25855 11234 25889
rect 11268 25855 11306 25889
rect 11340 25855 11378 25889
rect 11412 25855 11450 25889
rect 11484 25855 11522 25889
rect 11556 25855 11594 25889
rect 11628 25855 11666 25889
rect 11700 25855 11738 25889
rect 11772 25855 11810 25889
rect 11844 25855 11882 25889
rect 11916 25855 11954 25889
rect 11988 25855 12026 25889
rect 12060 25855 12098 25889
rect 12132 25855 12170 25889
rect 12204 25855 12242 25889
rect 12276 25855 12314 25889
rect 12348 25855 12386 25889
rect 12420 25855 12458 25889
rect 12492 25855 12530 25889
rect 12564 25855 12602 25889
rect 12636 25855 12674 25889
rect 12708 25855 12746 25889
rect 12780 25855 12818 25889
rect 12852 25855 12890 25889
rect 12924 25855 12962 25889
rect 12996 25855 13034 25889
rect 13068 25855 13106 25889
rect 13140 25855 13178 25889
rect 13212 25855 13250 25889
rect 13284 25855 13322 25889
rect 13356 25855 13394 25889
rect 13428 25855 13466 25889
rect 13500 25855 13538 25889
rect 13572 25855 13610 25889
rect 13644 25855 13682 25889
rect 13716 25855 13754 25889
rect 13788 25855 13826 25889
rect 13860 25855 13898 25889
rect 13932 25855 13970 25889
rect 14004 25855 14042 25889
rect 14076 25855 14114 25889
rect 14148 25855 14186 25889
rect 14220 25855 14258 25889
rect 14292 25855 14330 25889
rect 14364 25855 14402 25889
rect 14436 25855 14474 25889
rect 14508 25855 14546 25889
rect 14580 25855 14618 25889
rect 14652 25855 14690 25889
rect 14724 25855 14736 25889
rect 9616 25849 14736 25855
rect 231 25831 14736 25849
rect 231 25815 2480 25831
rect 2532 25815 2550 25831
rect 2602 25815 2620 25831
rect 2672 25815 3472 25831
rect 3524 25815 3542 25831
rect 3594 25815 3612 25831
rect 3664 25815 4464 25831
rect 231 25781 243 25815
rect 277 25781 316 25815
rect 350 25781 389 25815
rect 423 25781 462 25815
rect 496 25781 535 25815
rect 569 25781 608 25815
rect 642 25781 681 25815
rect 715 25781 754 25815
rect 788 25781 827 25815
rect 861 25781 900 25815
rect 934 25781 973 25815
rect 1007 25781 1046 25815
rect 1080 25781 1119 25815
rect 1153 25781 1192 25815
rect 1226 25781 1265 25815
rect 1299 25781 1338 25815
rect 1372 25781 1411 25815
rect 1445 25781 1484 25815
rect 1518 25781 1557 25815
rect 1591 25781 1630 25815
rect 1664 25781 1703 25815
rect 1737 25781 1776 25815
rect 1810 25781 1849 25815
rect 1883 25781 1922 25815
rect 1956 25781 1995 25815
rect 2029 25781 2068 25815
rect 2102 25781 2141 25815
rect 2175 25781 2214 25815
rect 2248 25781 2287 25815
rect 2321 25781 2360 25815
rect 2394 25781 2433 25815
rect 2467 25781 2480 25815
rect 2540 25781 2550 25815
rect 2613 25781 2620 25815
rect 2686 25781 2725 25815
rect 2759 25781 2798 25815
rect 2832 25781 2871 25815
rect 2905 25781 2944 25815
rect 2978 25781 3017 25815
rect 3051 25781 3090 25815
rect 3124 25781 3163 25815
rect 3197 25781 3236 25815
rect 3270 25781 3309 25815
rect 3343 25781 3382 25815
rect 3416 25781 3455 25815
rect 3524 25781 3528 25815
rect 3594 25781 3601 25815
rect 3664 25781 3674 25815
rect 3708 25781 3746 25815
rect 3780 25781 3818 25815
rect 3852 25781 3890 25815
rect 3924 25781 3962 25815
rect 3996 25781 4034 25815
rect 4068 25781 4106 25815
rect 4140 25781 4178 25815
rect 4212 25781 4250 25815
rect 4284 25781 4322 25815
rect 4356 25781 4394 25815
rect 4428 25781 4464 25815
rect 231 25779 2480 25781
rect 2532 25779 2550 25781
rect 2602 25779 2620 25781
rect 2672 25779 3472 25781
rect 3524 25779 3542 25781
rect 3594 25779 3612 25781
rect 3664 25779 4464 25781
rect 4516 25779 4534 25831
rect 4586 25779 4604 25831
rect 4656 25815 5456 25831
rect 4656 25781 4682 25815
rect 4716 25781 4754 25815
rect 4788 25781 4826 25815
rect 4860 25781 4898 25815
rect 4932 25781 4970 25815
rect 5004 25781 5042 25815
rect 5076 25781 5114 25815
rect 5148 25781 5186 25815
rect 5220 25781 5258 25815
rect 5292 25781 5330 25815
rect 5364 25781 5402 25815
rect 5436 25781 5456 25815
rect 4656 25779 5456 25781
rect 5508 25779 5526 25831
rect 5578 25815 5596 25831
rect 5648 25815 6448 25831
rect 6500 25815 6518 25831
rect 6570 25815 6588 25831
rect 6640 25815 7440 25831
rect 7492 25815 7510 25831
rect 7562 25815 7580 25831
rect 7632 25815 8432 25831
rect 8484 25815 8502 25831
rect 8554 25815 8572 25831
rect 8624 25815 9424 25831
rect 5580 25781 5596 25815
rect 5652 25781 5690 25815
rect 5724 25781 5762 25815
rect 5796 25781 5834 25815
rect 5868 25781 5906 25815
rect 5940 25781 5978 25815
rect 6012 25781 6050 25815
rect 6084 25781 6122 25815
rect 6156 25781 6194 25815
rect 6228 25781 6266 25815
rect 6300 25781 6338 25815
rect 6372 25781 6410 25815
rect 6444 25781 6448 25815
rect 6516 25781 6518 25815
rect 6660 25781 6698 25815
rect 6732 25781 6770 25815
rect 6804 25781 6842 25815
rect 6876 25781 6914 25815
rect 6948 25781 6986 25815
rect 7020 25781 7058 25815
rect 7092 25781 7130 25815
rect 7164 25781 7202 25815
rect 7236 25781 7274 25815
rect 7308 25781 7346 25815
rect 7380 25781 7418 25815
rect 7632 25781 7634 25815
rect 7668 25781 7706 25815
rect 7740 25781 7778 25815
rect 7812 25781 7850 25815
rect 7884 25781 7922 25815
rect 7956 25781 7994 25815
rect 8028 25781 8066 25815
rect 8100 25781 8138 25815
rect 8172 25781 8210 25815
rect 8244 25781 8282 25815
rect 8316 25781 8354 25815
rect 8388 25781 8426 25815
rect 8484 25781 8498 25815
rect 8554 25781 8570 25815
rect 8624 25781 8642 25815
rect 8676 25781 8714 25815
rect 8748 25781 8786 25815
rect 8820 25781 8858 25815
rect 8892 25781 8930 25815
rect 8964 25781 9002 25815
rect 9036 25781 9074 25815
rect 9108 25781 9146 25815
rect 9180 25781 9218 25815
rect 9252 25781 9290 25815
rect 9324 25781 9362 25815
rect 9396 25781 9424 25815
rect 5578 25779 5596 25781
rect 5648 25779 6448 25781
rect 6500 25779 6518 25781
rect 6570 25779 6588 25781
rect 6640 25779 7440 25781
rect 7492 25779 7510 25781
rect 7562 25779 7580 25781
rect 7632 25779 8432 25781
rect 8484 25779 8502 25781
rect 8554 25779 8572 25781
rect 8624 25779 9424 25781
rect 9476 25779 9494 25831
rect 9546 25779 9564 25831
rect 9616 25815 14736 25831
rect 9616 25781 9650 25815
rect 9684 25781 9722 25815
rect 9756 25781 9794 25815
rect 9828 25781 9866 25815
rect 9900 25781 9938 25815
rect 9972 25781 10010 25815
rect 10044 25781 10082 25815
rect 10116 25781 10154 25815
rect 10188 25781 10226 25815
rect 10260 25781 10298 25815
rect 10332 25781 10370 25815
rect 10404 25781 10442 25815
rect 10476 25781 10514 25815
rect 10548 25781 10586 25815
rect 10620 25781 10658 25815
rect 10692 25781 10730 25815
rect 10764 25781 10802 25815
rect 10836 25781 10874 25815
rect 10908 25781 10946 25815
rect 10980 25781 11018 25815
rect 11052 25781 11090 25815
rect 11124 25781 11162 25815
rect 11196 25781 11234 25815
rect 11268 25781 11306 25815
rect 11340 25781 11378 25815
rect 11412 25781 11450 25815
rect 11484 25781 11522 25815
rect 11556 25781 11594 25815
rect 11628 25781 11666 25815
rect 11700 25781 11738 25815
rect 11772 25781 11810 25815
rect 11844 25781 11882 25815
rect 11916 25781 11954 25815
rect 11988 25781 12026 25815
rect 12060 25781 12098 25815
rect 12132 25781 12170 25815
rect 12204 25781 12242 25815
rect 12276 25781 12314 25815
rect 12348 25781 12386 25815
rect 12420 25781 12458 25815
rect 12492 25781 12530 25815
rect 12564 25781 12602 25815
rect 12636 25781 12674 25815
rect 12708 25781 12746 25815
rect 12780 25781 12818 25815
rect 12852 25781 12890 25815
rect 12924 25781 12962 25815
rect 12996 25781 13034 25815
rect 13068 25781 13106 25815
rect 13140 25781 13178 25815
rect 13212 25781 13250 25815
rect 13284 25781 13322 25815
rect 13356 25781 13394 25815
rect 13428 25781 13466 25815
rect 13500 25781 13538 25815
rect 13572 25781 13610 25815
rect 13644 25781 13682 25815
rect 13716 25781 13754 25815
rect 13788 25781 13826 25815
rect 13860 25781 13898 25815
rect 13932 25781 13970 25815
rect 14004 25781 14042 25815
rect 14076 25781 14114 25815
rect 14148 25781 14186 25815
rect 14220 25781 14258 25815
rect 14292 25781 14330 25815
rect 14364 25781 14402 25815
rect 14436 25781 14474 25815
rect 14508 25781 14546 25815
rect 14580 25781 14618 25815
rect 14652 25781 14690 25815
rect 14724 25781 14736 25815
rect 9616 25779 14736 25781
rect 231 25760 14736 25779
rect 231 25741 2480 25760
rect 2532 25741 2550 25760
rect 2602 25741 2620 25760
rect 2672 25741 3472 25760
rect 3524 25741 3542 25760
rect 3594 25741 3612 25760
rect 3664 25741 4464 25760
rect 231 25707 243 25741
rect 277 25707 316 25741
rect 350 25707 389 25741
rect 423 25707 462 25741
rect 496 25707 535 25741
rect 569 25707 608 25741
rect 642 25707 681 25741
rect 715 25707 754 25741
rect 788 25707 827 25741
rect 861 25707 900 25741
rect 934 25707 973 25741
rect 1007 25707 1046 25741
rect 1080 25707 1119 25741
rect 1153 25707 1192 25741
rect 1226 25707 1265 25741
rect 1299 25707 1338 25741
rect 1372 25707 1411 25741
rect 1445 25707 1484 25741
rect 1518 25707 1557 25741
rect 1591 25707 1630 25741
rect 1664 25707 1703 25741
rect 1737 25707 1776 25741
rect 1810 25707 1849 25741
rect 1883 25707 1922 25741
rect 1956 25707 1995 25741
rect 2029 25707 2068 25741
rect 2102 25707 2141 25741
rect 2175 25707 2214 25741
rect 2248 25707 2287 25741
rect 2321 25707 2360 25741
rect 2394 25707 2433 25741
rect 2467 25708 2480 25741
rect 2540 25708 2550 25741
rect 2613 25708 2620 25741
rect 2467 25707 2506 25708
rect 2540 25707 2579 25708
rect 2613 25707 2652 25708
rect 2686 25707 2725 25741
rect 2759 25707 2798 25741
rect 2832 25707 2871 25741
rect 2905 25707 2944 25741
rect 2978 25707 3017 25741
rect 3051 25707 3090 25741
rect 3124 25707 3163 25741
rect 3197 25707 3236 25741
rect 3270 25707 3309 25741
rect 3343 25707 3382 25741
rect 3416 25707 3455 25741
rect 3524 25708 3528 25741
rect 3594 25708 3601 25741
rect 3664 25708 3674 25741
rect 3489 25707 3528 25708
rect 3562 25707 3601 25708
rect 3635 25707 3674 25708
rect 3708 25707 3746 25741
rect 3780 25707 3818 25741
rect 3852 25707 3890 25741
rect 3924 25707 3962 25741
rect 3996 25707 4034 25741
rect 4068 25707 4106 25741
rect 4140 25707 4178 25741
rect 4212 25707 4250 25741
rect 4284 25707 4322 25741
rect 4356 25707 4394 25741
rect 4428 25708 4464 25741
rect 4516 25708 4534 25760
rect 4586 25708 4604 25760
rect 4656 25741 5456 25760
rect 4656 25708 4682 25741
rect 4428 25707 4466 25708
rect 4500 25707 4538 25708
rect 4572 25707 4610 25708
rect 4644 25707 4682 25708
rect 4716 25707 4754 25741
rect 4788 25707 4826 25741
rect 4860 25707 4898 25741
rect 4932 25707 4970 25741
rect 5004 25707 5042 25741
rect 5076 25707 5114 25741
rect 5148 25707 5186 25741
rect 5220 25707 5258 25741
rect 5292 25707 5330 25741
rect 5364 25707 5402 25741
rect 5436 25708 5456 25741
rect 5508 25708 5526 25760
rect 5578 25741 5596 25760
rect 5648 25741 6448 25760
rect 6500 25741 6518 25760
rect 6570 25741 6588 25760
rect 6640 25741 7440 25760
rect 7492 25741 7510 25760
rect 7562 25741 7580 25760
rect 7632 25741 8432 25760
rect 8484 25741 8502 25760
rect 8554 25741 8572 25760
rect 8624 25741 9424 25760
rect 5580 25708 5596 25741
rect 5436 25707 5474 25708
rect 5508 25707 5546 25708
rect 5580 25707 5618 25708
rect 5652 25707 5690 25741
rect 5724 25707 5762 25741
rect 5796 25707 5834 25741
rect 5868 25707 5906 25741
rect 5940 25707 5978 25741
rect 6012 25707 6050 25741
rect 6084 25707 6122 25741
rect 6156 25707 6194 25741
rect 6228 25707 6266 25741
rect 6300 25707 6338 25741
rect 6372 25707 6410 25741
rect 6444 25708 6448 25741
rect 6516 25708 6518 25741
rect 6444 25707 6482 25708
rect 6516 25707 6554 25708
rect 6588 25707 6626 25708
rect 6660 25707 6698 25741
rect 6732 25707 6770 25741
rect 6804 25707 6842 25741
rect 6876 25707 6914 25741
rect 6948 25707 6986 25741
rect 7020 25707 7058 25741
rect 7092 25707 7130 25741
rect 7164 25707 7202 25741
rect 7236 25707 7274 25741
rect 7308 25707 7346 25741
rect 7380 25707 7418 25741
rect 7632 25708 7634 25741
rect 7452 25707 7490 25708
rect 7524 25707 7562 25708
rect 7596 25707 7634 25708
rect 7668 25707 7706 25741
rect 7740 25707 7778 25741
rect 7812 25707 7850 25741
rect 7884 25707 7922 25741
rect 7956 25707 7994 25741
rect 8028 25707 8066 25741
rect 8100 25707 8138 25741
rect 8172 25707 8210 25741
rect 8244 25707 8282 25741
rect 8316 25707 8354 25741
rect 8388 25707 8426 25741
rect 8484 25708 8498 25741
rect 8554 25708 8570 25741
rect 8624 25708 8642 25741
rect 8460 25707 8498 25708
rect 8532 25707 8570 25708
rect 8604 25707 8642 25708
rect 8676 25707 8714 25741
rect 8748 25707 8786 25741
rect 8820 25707 8858 25741
rect 8892 25707 8930 25741
rect 8964 25707 9002 25741
rect 9036 25707 9074 25741
rect 9108 25707 9146 25741
rect 9180 25707 9218 25741
rect 9252 25707 9290 25741
rect 9324 25707 9362 25741
rect 9396 25708 9424 25741
rect 9476 25708 9494 25760
rect 9546 25708 9564 25760
rect 9616 25741 14736 25760
rect 9616 25708 9650 25741
rect 9396 25707 9434 25708
rect 9468 25707 9506 25708
rect 9540 25707 9578 25708
rect 9612 25707 9650 25708
rect 9684 25707 9722 25741
rect 9756 25707 9794 25741
rect 9828 25707 9866 25741
rect 9900 25707 9938 25741
rect 9972 25707 10010 25741
rect 10044 25707 10082 25741
rect 10116 25707 10154 25741
rect 10188 25707 10226 25741
rect 10260 25707 10298 25741
rect 10332 25707 10370 25741
rect 10404 25707 10442 25741
rect 10476 25707 10514 25741
rect 10548 25707 10586 25741
rect 10620 25707 10658 25741
rect 10692 25707 10730 25741
rect 10764 25707 10802 25741
rect 10836 25707 10874 25741
rect 10908 25707 10946 25741
rect 10980 25707 11018 25741
rect 11052 25707 11090 25741
rect 11124 25707 11162 25741
rect 11196 25707 11234 25741
rect 11268 25707 11306 25741
rect 11340 25707 11378 25741
rect 11412 25707 11450 25741
rect 11484 25707 11522 25741
rect 11556 25707 11594 25741
rect 11628 25707 11666 25741
rect 11700 25707 11738 25741
rect 11772 25707 11810 25741
rect 11844 25707 11882 25741
rect 11916 25707 11954 25741
rect 11988 25707 12026 25741
rect 12060 25707 12098 25741
rect 12132 25707 12170 25741
rect 12204 25707 12242 25741
rect 12276 25707 12314 25741
rect 12348 25707 12386 25741
rect 12420 25707 12458 25741
rect 12492 25707 12530 25741
rect 12564 25707 12602 25741
rect 12636 25707 12674 25741
rect 12708 25707 12746 25741
rect 12780 25707 12818 25741
rect 12852 25707 12890 25741
rect 12924 25707 12962 25741
rect 12996 25707 13034 25741
rect 13068 25707 13106 25741
rect 13140 25707 13178 25741
rect 13212 25707 13250 25741
rect 13284 25707 13322 25741
rect 13356 25707 13394 25741
rect 13428 25707 13466 25741
rect 13500 25707 13538 25741
rect 13572 25707 13610 25741
rect 13644 25707 13682 25741
rect 13716 25707 13754 25741
rect 13788 25707 13826 25741
rect 13860 25707 13898 25741
rect 13932 25707 13970 25741
rect 14004 25707 14042 25741
rect 14076 25707 14114 25741
rect 14148 25707 14186 25741
rect 14220 25707 14258 25741
rect 14292 25707 14330 25741
rect 14364 25707 14402 25741
rect 14436 25707 14474 25741
rect 14508 25707 14546 25741
rect 14580 25707 14618 25741
rect 14652 25707 14690 25741
rect 14724 25707 14736 25741
rect 231 25689 14736 25707
rect 231 25667 2480 25689
rect 2532 25667 2550 25689
rect 2602 25667 2620 25689
rect 2672 25667 3472 25689
rect 3524 25667 3542 25689
rect 3594 25667 3612 25689
rect 3664 25667 4464 25689
rect 231 25633 243 25667
rect 277 25633 316 25667
rect 350 25633 389 25667
rect 423 25633 462 25667
rect 496 25633 535 25667
rect 569 25633 608 25667
rect 642 25633 681 25667
rect 715 25633 754 25667
rect 788 25633 827 25667
rect 861 25633 900 25667
rect 934 25633 973 25667
rect 1007 25633 1046 25667
rect 1080 25633 1119 25667
rect 1153 25633 1192 25667
rect 1226 25633 1265 25667
rect 1299 25633 1338 25667
rect 1372 25633 1411 25667
rect 1445 25633 1484 25667
rect 1518 25633 1557 25667
rect 1591 25633 1630 25667
rect 1664 25633 1703 25667
rect 1737 25633 1776 25667
rect 1810 25633 1849 25667
rect 1883 25633 1922 25667
rect 1956 25633 1995 25667
rect 2029 25633 2068 25667
rect 2102 25633 2141 25667
rect 2175 25633 2214 25667
rect 2248 25633 2287 25667
rect 2321 25633 2360 25667
rect 2394 25633 2433 25667
rect 2467 25637 2480 25667
rect 2540 25637 2550 25667
rect 2613 25637 2620 25667
rect 2467 25633 2506 25637
rect 2540 25633 2579 25637
rect 2613 25633 2652 25637
rect 2686 25633 2725 25667
rect 2759 25633 2798 25667
rect 2832 25633 2871 25667
rect 2905 25633 2944 25667
rect 2978 25633 3017 25667
rect 3051 25633 3090 25667
rect 3124 25633 3163 25667
rect 3197 25633 3236 25667
rect 3270 25633 3309 25667
rect 3343 25633 3382 25667
rect 3416 25633 3455 25667
rect 3524 25637 3528 25667
rect 3594 25637 3601 25667
rect 3664 25637 3674 25667
rect 3489 25633 3528 25637
rect 3562 25633 3601 25637
rect 3635 25633 3674 25637
rect 3708 25633 3746 25667
rect 3780 25633 3818 25667
rect 3852 25633 3890 25667
rect 3924 25633 3962 25667
rect 3996 25633 4034 25667
rect 4068 25633 4106 25667
rect 4140 25633 4178 25667
rect 4212 25633 4250 25667
rect 4284 25633 4322 25667
rect 4356 25633 4394 25667
rect 4428 25637 4464 25667
rect 4516 25637 4534 25689
rect 4586 25637 4604 25689
rect 4656 25667 5456 25689
rect 4656 25637 4682 25667
rect 4428 25633 4466 25637
rect 4500 25633 4538 25637
rect 4572 25633 4610 25637
rect 4644 25633 4682 25637
rect 4716 25633 4754 25667
rect 4788 25633 4826 25667
rect 4860 25633 4898 25667
rect 4932 25633 4970 25667
rect 5004 25633 5042 25667
rect 5076 25633 5114 25667
rect 5148 25633 5186 25667
rect 5220 25633 5258 25667
rect 5292 25633 5330 25667
rect 5364 25633 5402 25667
rect 5436 25637 5456 25667
rect 5508 25637 5526 25689
rect 5578 25667 5596 25689
rect 5648 25667 6448 25689
rect 6500 25667 6518 25689
rect 6570 25667 6588 25689
rect 6640 25667 7440 25689
rect 7492 25667 7510 25689
rect 7562 25667 7580 25689
rect 7632 25667 8432 25689
rect 8484 25667 8502 25689
rect 8554 25667 8572 25689
rect 8624 25667 9424 25689
rect 5580 25637 5596 25667
rect 5436 25633 5474 25637
rect 5508 25633 5546 25637
rect 5580 25633 5618 25637
rect 5652 25633 5690 25667
rect 5724 25633 5762 25667
rect 5796 25633 5834 25667
rect 5868 25633 5906 25667
rect 5940 25633 5978 25667
rect 6012 25633 6050 25667
rect 6084 25633 6122 25667
rect 6156 25633 6194 25667
rect 6228 25633 6266 25667
rect 6300 25633 6338 25667
rect 6372 25633 6410 25667
rect 6444 25637 6448 25667
rect 6516 25637 6518 25667
rect 6444 25633 6482 25637
rect 6516 25633 6554 25637
rect 6588 25633 6626 25637
rect 6660 25633 6698 25667
rect 6732 25633 6770 25667
rect 6804 25633 6842 25667
rect 6876 25633 6914 25667
rect 6948 25633 6986 25667
rect 7020 25633 7058 25667
rect 7092 25633 7130 25667
rect 7164 25633 7202 25667
rect 7236 25633 7274 25667
rect 7308 25633 7346 25667
rect 7380 25633 7418 25667
rect 7632 25637 7634 25667
rect 7452 25633 7490 25637
rect 7524 25633 7562 25637
rect 7596 25633 7634 25637
rect 7668 25633 7706 25667
rect 7740 25633 7778 25667
rect 7812 25633 7850 25667
rect 7884 25633 7922 25667
rect 7956 25633 7994 25667
rect 8028 25633 8066 25667
rect 8100 25633 8138 25667
rect 8172 25633 8210 25667
rect 8244 25633 8282 25667
rect 8316 25633 8354 25667
rect 8388 25633 8426 25667
rect 8484 25637 8498 25667
rect 8554 25637 8570 25667
rect 8624 25637 8642 25667
rect 8460 25633 8498 25637
rect 8532 25633 8570 25637
rect 8604 25633 8642 25637
rect 8676 25633 8714 25667
rect 8748 25633 8786 25667
rect 8820 25633 8858 25667
rect 8892 25633 8930 25667
rect 8964 25633 9002 25667
rect 9036 25633 9074 25667
rect 9108 25633 9146 25667
rect 9180 25633 9218 25667
rect 9252 25633 9290 25667
rect 9324 25633 9362 25667
rect 9396 25637 9424 25667
rect 9476 25637 9494 25689
rect 9546 25637 9564 25689
rect 9616 25667 14736 25689
rect 9616 25637 9650 25667
rect 9396 25633 9434 25637
rect 9468 25633 9506 25637
rect 9540 25633 9578 25637
rect 9612 25633 9650 25637
rect 9684 25633 9722 25667
rect 9756 25633 9794 25667
rect 9828 25633 9866 25667
rect 9900 25633 9938 25667
rect 9972 25633 10010 25667
rect 10044 25633 10082 25667
rect 10116 25633 10154 25667
rect 10188 25633 10226 25667
rect 10260 25633 10298 25667
rect 10332 25633 10370 25667
rect 10404 25633 10442 25667
rect 10476 25633 10514 25667
rect 10548 25633 10586 25667
rect 10620 25633 10658 25667
rect 10692 25633 10730 25667
rect 10764 25633 10802 25667
rect 10836 25633 10874 25667
rect 10908 25633 10946 25667
rect 10980 25633 11018 25667
rect 11052 25633 11090 25667
rect 11124 25633 11162 25667
rect 11196 25633 11234 25667
rect 11268 25633 11306 25667
rect 11340 25633 11378 25667
rect 11412 25633 11450 25667
rect 11484 25633 11522 25667
rect 11556 25633 11594 25667
rect 11628 25633 11666 25667
rect 11700 25633 11738 25667
rect 11772 25633 11810 25667
rect 11844 25633 11882 25667
rect 11916 25633 11954 25667
rect 11988 25633 12026 25667
rect 12060 25633 12098 25667
rect 12132 25633 12170 25667
rect 12204 25633 12242 25667
rect 12276 25633 12314 25667
rect 12348 25633 12386 25667
rect 12420 25633 12458 25667
rect 12492 25633 12530 25667
rect 12564 25633 12602 25667
rect 12636 25633 12674 25667
rect 12708 25633 12746 25667
rect 12780 25633 12818 25667
rect 12852 25633 12890 25667
rect 12924 25633 12962 25667
rect 12996 25633 13034 25667
rect 13068 25633 13106 25667
rect 13140 25633 13178 25667
rect 13212 25633 13250 25667
rect 13284 25633 13322 25667
rect 13356 25633 13394 25667
rect 13428 25633 13466 25667
rect 13500 25633 13538 25667
rect 13572 25633 13610 25667
rect 13644 25633 13682 25667
rect 13716 25633 13754 25667
rect 13788 25633 13826 25667
rect 13860 25633 13898 25667
rect 13932 25633 13970 25667
rect 14004 25633 14042 25667
rect 14076 25633 14114 25667
rect 14148 25633 14186 25667
rect 14220 25633 14258 25667
rect 14292 25633 14330 25667
rect 14364 25633 14402 25667
rect 14436 25633 14474 25667
rect 14508 25633 14546 25667
rect 14580 25633 14618 25667
rect 14652 25633 14690 25667
rect 14724 25633 14736 25667
rect 231 25625 14736 25633
rect -29 25041 15029 25052
rect -29 25007 88 25041
rect 122 25007 161 25041
rect 195 25007 234 25041
rect 268 25007 307 25041
rect 341 25007 380 25041
rect 414 25007 453 25041
rect 487 25007 526 25041
rect 560 25007 599 25041
rect 633 25007 672 25041
rect 706 25007 745 25041
rect 779 25007 818 25041
rect 852 25007 891 25041
rect 925 25007 964 25041
rect 998 25007 1037 25041
rect 1071 25007 1110 25041
rect 1144 25007 1183 25041
rect 1217 25007 1256 25041
rect 1290 25037 1329 25041
rect 1363 25037 1402 25041
rect 1436 25037 1475 25041
rect 1509 25037 1548 25041
rect 1582 25037 1621 25041
rect 1655 25037 1694 25041
rect 1728 25037 1767 25041
rect 1801 25037 1840 25041
rect 1874 25037 1913 25041
rect 1947 25037 1986 25041
rect 2020 25037 2059 25041
rect 1290 25007 1303 25037
rect 1363 25007 1371 25037
rect 1436 25007 1439 25037
rect 1763 25007 1767 25037
rect 1831 25007 1840 25037
rect 1899 25007 1913 25037
rect -29 24985 1303 25007
rect 1355 24985 1371 25007
rect 1423 24985 1439 25007
rect 1491 24985 1507 25007
rect 1559 24985 1575 25007
rect 1627 24985 1643 25007
rect 1695 24985 1711 25007
rect 1763 24985 1779 25007
rect 1831 24985 1847 25007
rect 1899 24985 1914 25007
rect 1966 24985 1981 25037
rect 2033 25007 2059 25037
rect 2093 25007 2132 25041
rect 2166 25007 2205 25041
rect 2239 25007 2278 25041
rect 2312 25007 2351 25041
rect 2385 25007 2424 25041
rect 2458 25007 2497 25041
rect 2531 25007 2570 25041
rect 2604 25007 2643 25041
rect 2677 25007 2716 25041
rect 2750 25007 2789 25041
rect 2823 25007 2862 25041
rect 2896 25007 2935 25041
rect 2969 25007 3008 25041
rect 3042 25007 3081 25041
rect 3115 25007 3154 25041
rect 3188 25007 3227 25041
rect 3261 25007 3300 25041
rect 3334 25007 3373 25041
rect 3407 25007 3446 25041
rect 3480 25007 3519 25041
rect 3553 25007 3592 25041
rect 3626 25007 3665 25041
rect 3699 25007 3738 25041
rect 3772 25007 3811 25041
rect 3845 25007 3884 25041
rect 3918 25007 3957 25041
rect 3991 25007 4030 25041
rect 4064 25007 4103 25041
rect 4137 25007 4176 25041
rect 4210 25007 4249 25041
rect 4283 25007 4322 25041
rect 4356 25007 4395 25041
rect 4429 25007 4468 25041
rect 2033 24985 4468 25007
rect -29 24969 4468 24985
rect -29 24935 88 24969
rect 122 24935 161 24969
rect 195 24935 234 24969
rect 268 24935 307 24969
rect 341 24935 380 24969
rect 414 24935 453 24969
rect 487 24935 526 24969
rect 560 24935 599 24969
rect 633 24935 672 24969
rect 706 24935 745 24969
rect 779 24935 818 24969
rect 852 24935 891 24969
rect 925 24935 964 24969
rect 998 24935 1037 24969
rect 1071 24935 1110 24969
rect 1144 24935 1183 24969
rect 1217 24935 1256 24969
rect 1290 24967 1329 24969
rect 1363 24967 1402 24969
rect 1436 24967 1475 24969
rect 1509 24967 1548 24969
rect 1582 24967 1621 24969
rect 1655 24967 1694 24969
rect 1728 24967 1767 24969
rect 1801 24967 1840 24969
rect 1874 24967 1913 24969
rect 1947 24967 1986 24969
rect 2020 24967 2059 24969
rect 1290 24935 1303 24967
rect 1363 24935 1371 24967
rect 1436 24935 1439 24967
rect 1763 24935 1767 24967
rect 1831 24935 1840 24967
rect 1899 24935 1913 24967
rect -29 24915 1303 24935
rect 1355 24915 1371 24935
rect 1423 24915 1439 24935
rect 1491 24915 1507 24935
rect 1559 24915 1575 24935
rect 1627 24915 1643 24935
rect 1695 24915 1711 24935
rect 1763 24915 1779 24935
rect 1831 24915 1847 24935
rect 1899 24915 1914 24935
rect 1966 24915 1981 24967
rect 2033 24935 2059 24967
rect 2093 24935 2132 24969
rect 2166 24935 2205 24969
rect 2239 24935 2278 24969
rect 2312 24935 2351 24969
rect 2385 24935 2424 24969
rect 2458 24935 2497 24969
rect 2531 24935 2570 24969
rect 2604 24935 2643 24969
rect 2677 24935 2716 24969
rect 2750 24935 2789 24969
rect 2823 24935 2862 24969
rect 2896 24935 2935 24969
rect 2969 24935 3008 24969
rect 3042 24935 3081 24969
rect 3115 24935 3154 24969
rect 3188 24935 3227 24969
rect 3261 24935 3300 24969
rect 3334 24935 3373 24969
rect 3407 24935 3446 24969
rect 3480 24935 3519 24969
rect 3553 24935 3592 24969
rect 3626 24935 3665 24969
rect 3699 24935 3738 24969
rect 3772 24935 3811 24969
rect 3845 24935 3884 24969
rect 3918 24935 3957 24969
rect 3991 24935 4030 24969
rect 4064 24935 4103 24969
rect 4137 24935 4176 24969
rect 4210 24935 4249 24969
rect 4283 24935 4322 24969
rect 4356 24935 4395 24969
rect 4429 24935 4468 24969
rect 2033 24915 4468 24935
rect -29 24897 4468 24915
rect -29 24863 88 24897
rect 122 24863 161 24897
rect 195 24863 234 24897
rect 268 24863 307 24897
rect 341 24863 380 24897
rect 414 24863 453 24897
rect 487 24863 526 24897
rect 560 24863 599 24897
rect 633 24863 672 24897
rect 706 24863 745 24897
rect 779 24863 818 24897
rect 852 24863 891 24897
rect 925 24863 964 24897
rect 998 24863 1037 24897
rect 1071 24863 1110 24897
rect 1144 24863 1183 24897
rect 1217 24863 1256 24897
rect 1290 24863 1303 24897
rect 1363 24863 1371 24897
rect 1436 24863 1439 24897
rect 1763 24863 1767 24897
rect 1831 24863 1840 24897
rect 1899 24863 1913 24897
rect -29 24845 1303 24863
rect 1355 24845 1371 24863
rect 1423 24845 1439 24863
rect 1491 24845 1507 24863
rect 1559 24845 1575 24863
rect 1627 24845 1643 24863
rect 1695 24845 1711 24863
rect 1763 24845 1779 24863
rect 1831 24845 1847 24863
rect 1899 24845 1914 24863
rect 1966 24845 1981 24897
rect 2033 24863 2059 24897
rect 2093 24863 2132 24897
rect 2166 24863 2205 24897
rect 2239 24863 2278 24897
rect 2312 24863 2351 24897
rect 2385 24863 2424 24897
rect 2458 24863 2497 24897
rect 2531 24863 2570 24897
rect 2604 24863 2643 24897
rect 2677 24863 2716 24897
rect 2750 24863 2789 24897
rect 2823 24863 2862 24897
rect 2896 24863 2935 24897
rect 2969 24863 3008 24897
rect 3042 24863 3081 24897
rect 3115 24863 3154 24897
rect 3188 24863 3227 24897
rect 3261 24863 3300 24897
rect 3334 24863 3373 24897
rect 3407 24863 3446 24897
rect 3480 24863 3519 24897
rect 3553 24863 3592 24897
rect 3626 24863 3665 24897
rect 3699 24863 3738 24897
rect 3772 24863 3811 24897
rect 3845 24863 3884 24897
rect 3918 24863 3957 24897
rect 3991 24863 4030 24897
rect 4064 24863 4103 24897
rect 4137 24863 4176 24897
rect 4210 24863 4249 24897
rect 4283 24863 4322 24897
rect 4356 24863 4395 24897
rect 4429 24863 4468 24897
rect 2033 24845 4468 24863
rect -29 24827 4468 24845
rect -29 24825 1303 24827
rect 1355 24825 1371 24827
rect 1423 24825 1439 24827
rect 1491 24825 1507 24827
rect 1559 24825 1575 24827
rect 1627 24825 1643 24827
rect 1695 24825 1711 24827
rect 1763 24825 1779 24827
rect 1831 24825 1847 24827
rect 1899 24825 1914 24827
rect -29 24791 88 24825
rect 122 24791 161 24825
rect 195 24791 234 24825
rect 268 24791 307 24825
rect 341 24791 380 24825
rect 414 24791 453 24825
rect 487 24791 526 24825
rect 560 24791 599 24825
rect 633 24791 672 24825
rect 706 24791 745 24825
rect 779 24791 818 24825
rect 852 24791 891 24825
rect 925 24791 964 24825
rect 998 24791 1037 24825
rect 1071 24791 1110 24825
rect 1144 24791 1183 24825
rect 1217 24791 1256 24825
rect 1290 24791 1303 24825
rect 1363 24791 1371 24825
rect 1436 24791 1439 24825
rect 1763 24791 1767 24825
rect 1831 24791 1840 24825
rect 1899 24791 1913 24825
rect -29 24775 1303 24791
rect 1355 24775 1371 24791
rect 1423 24775 1439 24791
rect 1491 24775 1507 24791
rect 1559 24775 1575 24791
rect 1627 24775 1643 24791
rect 1695 24775 1711 24791
rect 1763 24775 1779 24791
rect 1831 24775 1847 24791
rect 1899 24775 1914 24791
rect 1966 24775 1981 24827
rect 2033 24825 4468 24827
rect 2033 24791 2059 24825
rect 2093 24791 2132 24825
rect 2166 24791 2205 24825
rect 2239 24791 2278 24825
rect 2312 24791 2351 24825
rect 2385 24791 2424 24825
rect 2458 24791 2497 24825
rect 2531 24791 2570 24825
rect 2604 24791 2643 24825
rect 2677 24791 2716 24825
rect 2750 24791 2789 24825
rect 2823 24791 2862 24825
rect 2896 24791 2935 24825
rect 2969 24791 3008 24825
rect 3042 24791 3081 24825
rect 3115 24791 3154 24825
rect 3188 24791 3227 24825
rect 3261 24791 3300 24825
rect 3334 24791 3373 24825
rect 3407 24791 3446 24825
rect 3480 24791 3519 24825
rect 3553 24791 3592 24825
rect 3626 24791 3665 24825
rect 3699 24791 3738 24825
rect 3772 24791 3811 24825
rect 3845 24791 3884 24825
rect 3918 24791 3957 24825
rect 3991 24791 4030 24825
rect 4064 24791 4103 24825
rect 4137 24791 4176 24825
rect 4210 24791 4249 24825
rect 4283 24791 4322 24825
rect 4356 24791 4395 24825
rect 4429 24791 4468 24825
rect 2033 24775 4468 24791
rect -29 24757 4468 24775
rect -29 24753 1303 24757
rect 1355 24753 1371 24757
rect 1423 24753 1439 24757
rect 1491 24753 1507 24757
rect 1559 24753 1575 24757
rect 1627 24753 1643 24757
rect 1695 24753 1711 24757
rect 1763 24753 1779 24757
rect 1831 24753 1847 24757
rect 1899 24753 1914 24757
rect -29 24719 88 24753
rect 122 24719 161 24753
rect 195 24719 234 24753
rect 268 24719 307 24753
rect 341 24719 380 24753
rect 414 24719 453 24753
rect 487 24719 526 24753
rect 560 24719 599 24753
rect 633 24719 672 24753
rect 706 24719 745 24753
rect 779 24719 818 24753
rect 852 24719 891 24753
rect 925 24719 964 24753
rect 998 24719 1037 24753
rect 1071 24719 1110 24753
rect 1144 24719 1183 24753
rect 1217 24719 1256 24753
rect 1290 24719 1303 24753
rect 1363 24719 1371 24753
rect 1436 24719 1439 24753
rect 1763 24719 1767 24753
rect 1831 24719 1840 24753
rect 1899 24719 1913 24753
rect -29 24705 1303 24719
rect 1355 24705 1371 24719
rect 1423 24705 1439 24719
rect 1491 24705 1507 24719
rect 1559 24705 1575 24719
rect 1627 24705 1643 24719
rect 1695 24705 1711 24719
rect 1763 24705 1779 24719
rect 1831 24705 1847 24719
rect 1899 24705 1914 24719
rect 1966 24705 1981 24757
rect 2033 24753 4468 24757
rect 2033 24719 2059 24753
rect 2093 24719 2132 24753
rect 2166 24719 2205 24753
rect 2239 24719 2278 24753
rect 2312 24719 2351 24753
rect 2385 24719 2424 24753
rect 2458 24719 2497 24753
rect 2531 24719 2570 24753
rect 2604 24719 2643 24753
rect 2677 24719 2716 24753
rect 2750 24719 2789 24753
rect 2823 24719 2862 24753
rect 2896 24719 2935 24753
rect 2969 24719 3008 24753
rect 3042 24719 3081 24753
rect 3115 24719 3154 24753
rect 3188 24719 3227 24753
rect 3261 24719 3300 24753
rect 3334 24719 3373 24753
rect 3407 24719 3446 24753
rect 3480 24719 3519 24753
rect 3553 24719 3592 24753
rect 3626 24719 3665 24753
rect 3699 24719 3738 24753
rect 3772 24719 3811 24753
rect 3845 24719 3884 24753
rect 3918 24719 3957 24753
rect 3991 24719 4030 24753
rect 4064 24719 4103 24753
rect 4137 24719 4176 24753
rect 4210 24719 4249 24753
rect 4283 24719 4322 24753
rect 4356 24719 4395 24753
rect 4429 24719 4468 24753
rect 14870 24719 15029 25041
rect 2033 24705 12157 24719
rect 12209 24705 12225 24719
rect 12277 24705 12293 24719
rect 12345 24705 12361 24719
rect 12413 24705 12429 24719
rect 12481 24705 12497 24719
rect 12549 24705 12565 24719
rect 12617 24705 12633 24719
rect 12685 24705 12701 24719
rect 12753 24705 12768 24719
rect 12820 24705 12835 24719
rect 12887 24705 15029 24719
rect -29 24687 15029 24705
rect -29 24683 1303 24687
rect 1297 24635 1303 24683
rect 1355 24635 1371 24687
rect 1423 24635 1439 24687
rect 1491 24635 1507 24687
rect 1559 24635 1575 24687
rect 1627 24635 1643 24687
rect 1695 24635 1711 24687
rect 1763 24635 1779 24687
rect 1831 24635 1847 24687
rect 1899 24635 1914 24687
rect 1966 24635 1981 24687
rect 2033 24683 12157 24687
rect 2033 24635 2039 24683
rect 1297 24617 2039 24635
rect 1297 24565 1303 24617
rect 1355 24565 1371 24617
rect 1423 24565 1439 24617
rect 1491 24565 1507 24617
rect 1559 24565 1575 24617
rect 1627 24565 1643 24617
rect 1695 24565 1711 24617
rect 1763 24565 1779 24617
rect 1831 24565 1847 24617
rect 1899 24565 1914 24617
rect 1966 24565 1981 24617
rect 2033 24565 2039 24617
rect 1297 24547 2039 24565
rect 1297 24495 1303 24547
rect 1355 24495 1371 24547
rect 1423 24495 1439 24547
rect 1491 24495 1507 24547
rect 1559 24495 1575 24547
rect 1627 24495 1643 24547
rect 1695 24495 1711 24547
rect 1763 24495 1779 24547
rect 1831 24495 1847 24547
rect 1899 24495 1914 24547
rect 1966 24495 1981 24547
rect 2033 24495 2039 24547
rect 1297 24493 2039 24495
rect 12151 24635 12157 24683
rect 12209 24635 12225 24687
rect 12277 24635 12293 24687
rect 12345 24635 12361 24687
rect 12413 24635 12429 24687
rect 12481 24635 12497 24687
rect 12549 24635 12565 24687
rect 12617 24635 12633 24687
rect 12685 24635 12701 24687
rect 12753 24635 12768 24687
rect 12820 24635 12835 24687
rect 12887 24683 15029 24687
rect 12887 24635 12893 24683
rect 12151 24617 12893 24635
rect 12151 24565 12157 24617
rect 12209 24565 12225 24617
rect 12277 24565 12293 24617
rect 12345 24565 12361 24617
rect 12413 24565 12429 24617
rect 12481 24565 12497 24617
rect 12549 24565 12565 24617
rect 12617 24565 12633 24617
rect 12685 24565 12701 24617
rect 12753 24565 12768 24617
rect 12820 24565 12835 24617
rect 12887 24565 12893 24617
rect 12151 24547 12893 24565
rect 12151 24495 12157 24547
rect 12209 24495 12225 24547
rect 12277 24495 12293 24547
rect 12345 24495 12361 24547
rect 12413 24495 12429 24547
rect 12481 24495 12497 24547
rect 12549 24495 12565 24547
rect 12617 24495 12633 24547
rect 12685 24495 12701 24547
rect 12753 24495 12768 24547
rect 12820 24495 12835 24547
rect 12887 24495 12893 24547
rect 12151 24493 12893 24495
rect 14754 21413 14940 21419
rect 14754 21361 14755 21413
rect 14807 21361 14821 21413
rect 14873 21361 14887 21413
rect 14939 21361 14940 21413
rect 14754 21348 14940 21361
rect 14754 21296 14755 21348
rect 14807 21296 14821 21348
rect 14873 21296 14887 21348
rect 14939 21296 14940 21348
rect 14754 21282 14940 21296
rect 14754 21230 14755 21282
rect 14807 21230 14821 21282
rect 14873 21230 14887 21282
rect 14939 21230 14940 21282
rect 14754 21216 14940 21230
rect 14754 21164 14755 21216
rect 14807 21164 14821 21216
rect 14873 21164 14887 21216
rect 14939 21164 14940 21216
rect 14754 21150 14940 21164
rect 14754 21098 14755 21150
rect 14807 21098 14821 21150
rect 14873 21098 14887 21150
rect 14939 21098 14940 21150
rect 14754 21084 14940 21098
rect 14754 21032 14755 21084
rect 14807 21032 14821 21084
rect 14873 21032 14887 21084
rect 14939 21032 14940 21084
rect 14754 21018 14940 21032
rect 14754 20966 14755 21018
rect 14807 20966 14821 21018
rect 14873 20966 14887 21018
rect 14939 20966 14940 21018
rect 14754 20952 14940 20966
rect 14754 20900 14755 20952
rect 14807 20900 14821 20952
rect 14873 20900 14887 20952
rect 14939 20900 14940 20952
rect 14754 20886 14940 20900
rect 14754 20834 14755 20886
rect 14807 20834 14821 20886
rect 14873 20834 14887 20886
rect 14939 20834 14940 20886
rect 14754 20820 14940 20834
rect 14754 20768 14755 20820
rect 14807 20768 14821 20820
rect 14873 20768 14887 20820
rect 14939 20768 14940 20820
rect 14754 20754 14940 20768
rect 14754 20702 14755 20754
rect 14807 20702 14821 20754
rect 14873 20702 14887 20754
rect 14939 20702 14940 20754
rect 14754 20688 14940 20702
rect 14754 20636 14755 20688
rect 14807 20636 14821 20688
rect 14873 20636 14887 20688
rect 14939 20636 14940 20688
rect 14754 20622 14940 20636
rect 14754 20570 14755 20622
rect 14807 20570 14821 20622
rect 14873 20570 14887 20622
rect 14939 20570 14940 20622
rect 14754 20556 14940 20570
rect 14754 20504 14755 20556
rect 14807 20504 14821 20556
rect 14873 20504 14887 20556
rect 14939 20504 14940 20556
rect 14754 20490 14940 20504
rect 14754 20438 14755 20490
rect 14807 20438 14821 20490
rect 14873 20438 14887 20490
rect 14939 20438 14940 20490
rect 14754 20424 14940 20438
rect 14754 20372 14755 20424
rect 14807 20372 14821 20424
rect 14873 20372 14887 20424
rect 14939 20372 14940 20424
rect 14754 20358 14940 20372
rect 14754 20306 14755 20358
rect 14807 20306 14821 20358
rect 14873 20306 14887 20358
rect 14939 20306 14940 20358
rect 14754 20292 14940 20306
rect 14754 20240 14755 20292
rect 14807 20240 14821 20292
rect 14873 20240 14887 20292
rect 14939 20240 14940 20292
rect 14754 20226 14940 20240
rect 14754 20174 14755 20226
rect 14807 20174 14821 20226
rect 14873 20174 14887 20226
rect 14939 20174 14940 20226
rect 14754 20160 14940 20174
rect 14754 20108 14755 20160
rect 14807 20108 14821 20160
rect 14873 20108 14887 20160
rect 14939 20108 14940 20160
rect 14754 20094 14940 20108
rect 14754 20042 14755 20094
rect 14807 20042 14821 20094
rect 14873 20042 14887 20094
rect 14939 20042 14940 20094
rect 14754 20028 14940 20042
rect 14754 19976 14755 20028
rect 14807 19976 14821 20028
rect 14873 19976 14887 20028
rect 14939 19976 14940 20028
rect 195 19964 1266 19967
rect 195 19912 201 19964
rect 253 19912 269 19964
rect 321 19912 337 19964
rect 389 19912 404 19964
rect 456 19912 471 19964
rect 523 19912 538 19964
rect 590 19912 605 19964
rect 657 19912 672 19964
rect 724 19912 739 19964
rect 791 19912 806 19964
rect 858 19912 873 19964
rect 925 19912 940 19964
rect 992 19912 1007 19964
rect 1059 19912 1074 19964
rect 1126 19912 1141 19964
rect 1193 19912 1208 19964
rect 1260 19912 1266 19964
rect 195 19896 1266 19912
rect 195 19884 201 19896
rect -29 19858 201 19884
rect -29 19824 70 19858
rect 104 19824 143 19858
rect 177 19844 201 19858
rect 253 19844 269 19896
rect 321 19858 337 19896
rect 389 19858 404 19896
rect 456 19858 471 19896
rect 523 19858 538 19896
rect 590 19858 605 19896
rect 657 19858 672 19896
rect 724 19858 739 19896
rect 791 19858 806 19896
rect 323 19844 337 19858
rect 396 19844 404 19858
rect 469 19844 471 19858
rect 724 19844 727 19858
rect 791 19844 800 19858
rect 858 19844 873 19896
rect 925 19844 940 19896
rect 992 19844 1007 19896
rect 1059 19844 1074 19896
rect 1126 19844 1141 19896
rect 1193 19858 1208 19896
rect 1260 19884 1266 19896
rect 8194 19964 9265 19967
rect 8194 19912 8200 19964
rect 8252 19912 8268 19964
rect 8320 19912 8336 19964
rect 8388 19912 8403 19964
rect 8455 19912 8470 19964
rect 8522 19912 8537 19964
rect 8589 19912 8604 19964
rect 8656 19912 8671 19964
rect 8723 19912 8738 19964
rect 8790 19912 8805 19964
rect 8857 19912 8872 19964
rect 8924 19912 8939 19964
rect 8991 19912 9006 19964
rect 9058 19912 9073 19964
rect 9125 19912 9140 19964
rect 9192 19912 9207 19964
rect 9259 19912 9265 19964
rect 8194 19896 9265 19912
rect 8194 19884 8200 19896
rect 1260 19858 8200 19884
rect 8252 19858 8268 19896
rect 8320 19858 8336 19896
rect 8388 19858 8403 19896
rect 8455 19858 8470 19896
rect 1199 19844 1208 19858
rect 177 19828 216 19844
rect 250 19828 289 19844
rect 323 19828 362 19844
rect 396 19828 435 19844
rect 469 19828 508 19844
rect 542 19828 581 19844
rect 615 19828 654 19844
rect 688 19828 727 19844
rect 761 19828 800 19844
rect 834 19828 873 19844
rect 907 19828 946 19844
rect 980 19828 1019 19844
rect 1053 19828 1092 19844
rect 1126 19828 1165 19844
rect 1199 19828 1238 19844
rect 177 19824 201 19828
rect -29 19776 201 19824
rect 253 19776 269 19828
rect 323 19824 337 19828
rect 396 19824 404 19828
rect 469 19824 471 19828
rect 724 19824 727 19828
rect 791 19824 800 19828
rect 321 19776 337 19824
rect 389 19776 404 19824
rect 456 19776 471 19824
rect 523 19776 538 19824
rect 590 19776 605 19824
rect 657 19776 672 19824
rect 724 19776 739 19824
rect 791 19776 806 19824
rect 858 19776 873 19828
rect 925 19776 940 19828
rect 992 19776 1007 19828
rect 1059 19776 1074 19828
rect 1126 19776 1141 19828
rect 1199 19824 1208 19828
rect 1272 19824 1311 19858
rect 1345 19824 1384 19858
rect 1418 19824 1457 19858
rect 1491 19824 1530 19858
rect 1564 19824 1603 19858
rect 1637 19824 1676 19858
rect 1710 19824 1749 19858
rect 1783 19824 1822 19858
rect 1856 19824 1895 19858
rect 1929 19824 1968 19858
rect 2002 19824 2041 19858
rect 2075 19824 2114 19858
rect 2148 19824 2187 19858
rect 2221 19824 2260 19858
rect 2294 19824 2333 19858
rect 2367 19824 2406 19858
rect 2440 19824 2479 19858
rect 2513 19824 2552 19858
rect 2586 19824 2625 19858
rect 2659 19824 2698 19858
rect 2732 19824 2771 19858
rect 2805 19824 2844 19858
rect 2878 19824 2917 19858
rect 2951 19824 2990 19858
rect 3024 19824 3063 19858
rect 3097 19824 3136 19858
rect 3170 19824 3209 19858
rect 3243 19824 3282 19858
rect 3316 19824 3354 19858
rect 3388 19824 3426 19858
rect 3460 19824 3498 19858
rect 3532 19824 3570 19858
rect 3604 19824 3642 19858
rect 3676 19824 3714 19858
rect 3748 19824 3786 19858
rect 3820 19824 3858 19858
rect 3892 19824 3930 19858
rect 3964 19824 4002 19858
rect 4036 19824 4074 19858
rect 4108 19824 4146 19858
rect 4180 19824 4218 19858
rect 4252 19824 4290 19858
rect 4324 19824 4362 19858
rect 4396 19824 4434 19858
rect 4468 19824 4506 19858
rect 4540 19824 4578 19858
rect 4612 19824 4650 19858
rect 4684 19824 4722 19858
rect 4756 19824 4794 19858
rect 4828 19824 4866 19858
rect 4900 19824 4938 19858
rect 4972 19824 5010 19858
rect 5044 19824 5082 19858
rect 5116 19824 5154 19858
rect 5188 19824 5226 19858
rect 5260 19824 5298 19858
rect 5332 19824 5370 19858
rect 5404 19824 5442 19858
rect 5476 19824 5514 19858
rect 5548 19824 5586 19858
rect 5620 19824 5658 19858
rect 5692 19824 5730 19858
rect 5764 19824 5802 19858
rect 5836 19824 5874 19858
rect 5908 19824 5946 19858
rect 5980 19824 6018 19858
rect 6052 19824 6090 19858
rect 6124 19824 6162 19858
rect 6196 19824 6234 19858
rect 6268 19824 6306 19858
rect 6340 19824 6378 19858
rect 6412 19824 6450 19858
rect 6484 19824 6522 19858
rect 6556 19824 6594 19858
rect 6628 19824 6666 19858
rect 6700 19824 6738 19858
rect 6772 19824 6810 19858
rect 6844 19824 6882 19858
rect 6916 19824 6954 19858
rect 6988 19824 7026 19858
rect 7060 19824 7098 19858
rect 7132 19824 7170 19858
rect 7204 19824 7242 19858
rect 7276 19824 7314 19858
rect 7348 19824 7386 19858
rect 7420 19824 7458 19858
rect 7492 19824 7530 19858
rect 7564 19824 7602 19858
rect 7636 19824 7674 19858
rect 7708 19824 7746 19858
rect 7780 19824 7818 19858
rect 7852 19824 7890 19858
rect 7924 19824 7962 19858
rect 7996 19824 8034 19858
rect 8068 19824 8106 19858
rect 8140 19824 8178 19858
rect 8320 19844 8322 19858
rect 8388 19844 8394 19858
rect 8455 19844 8466 19858
rect 8522 19844 8537 19896
rect 8589 19844 8604 19896
rect 8656 19844 8671 19896
rect 8723 19844 8738 19896
rect 8790 19844 8805 19896
rect 8857 19858 8872 19896
rect 8924 19858 8939 19896
rect 8991 19858 9006 19896
rect 9058 19858 9073 19896
rect 9125 19858 9140 19896
rect 9192 19858 9207 19896
rect 9259 19884 9265 19896
rect 14754 19962 14940 19976
rect 14754 19910 14755 19962
rect 14807 19910 14821 19962
rect 14873 19910 14887 19962
rect 14939 19910 14940 19962
rect 14754 19896 14940 19910
rect 14754 19884 14755 19896
rect 9259 19858 14755 19884
rect 14807 19858 14821 19896
rect 14873 19858 14887 19896
rect 14939 19884 14940 19896
rect 14939 19864 15029 19884
rect 8860 19844 8872 19858
rect 8932 19844 8939 19858
rect 9004 19844 9006 19858
rect 8212 19828 8250 19844
rect 8284 19828 8322 19844
rect 8356 19828 8394 19844
rect 8428 19828 8466 19844
rect 8500 19828 8538 19844
rect 8572 19828 8610 19844
rect 8644 19828 8682 19844
rect 8716 19828 8754 19844
rect 8788 19828 8826 19844
rect 8860 19828 8898 19844
rect 8932 19828 8970 19844
rect 9004 19828 9042 19844
rect 9076 19828 9114 19844
rect 9148 19828 9186 19844
rect 9220 19828 9258 19844
rect 8320 19824 8322 19828
rect 8388 19824 8394 19828
rect 8455 19824 8466 19828
rect 1193 19776 1208 19824
rect 1260 19776 8200 19824
rect 8252 19776 8268 19824
rect 8320 19776 8336 19824
rect 8388 19776 8403 19824
rect 8455 19776 8470 19824
rect 8522 19776 8537 19828
rect 8589 19776 8604 19828
rect 8656 19776 8671 19828
rect 8723 19776 8738 19828
rect 8790 19776 8805 19828
rect 8860 19824 8872 19828
rect 8932 19824 8939 19828
rect 9004 19824 9006 19828
rect 9292 19824 9330 19858
rect 9364 19824 9402 19858
rect 9436 19824 9474 19858
rect 9508 19824 9546 19858
rect 9580 19824 9618 19858
rect 9652 19824 9690 19858
rect 9724 19824 9762 19858
rect 9796 19824 9834 19858
rect 9868 19824 9906 19858
rect 9940 19824 9978 19858
rect 10012 19824 10050 19858
rect 10084 19824 10122 19858
rect 10156 19824 10194 19858
rect 10228 19824 10266 19858
rect 10300 19824 10338 19858
rect 10372 19824 10410 19858
rect 10444 19824 10482 19858
rect 10516 19824 10554 19858
rect 10588 19824 10626 19858
rect 10660 19824 10698 19858
rect 10732 19824 10770 19858
rect 10804 19824 10842 19858
rect 10876 19824 10914 19858
rect 10948 19824 10986 19858
rect 11020 19824 11058 19858
rect 11092 19824 11130 19858
rect 11164 19824 11202 19858
rect 11236 19824 11274 19858
rect 11308 19824 11346 19858
rect 11380 19824 11418 19858
rect 11452 19824 11490 19858
rect 11524 19824 11562 19858
rect 11596 19824 11634 19858
rect 11668 19824 11706 19858
rect 11740 19824 11778 19858
rect 11812 19824 11850 19858
rect 11884 19824 11922 19858
rect 11956 19824 11994 19858
rect 12028 19824 12066 19858
rect 12100 19824 12138 19858
rect 12172 19824 12210 19858
rect 12244 19824 12282 19858
rect 12316 19824 12354 19858
rect 12388 19824 12426 19858
rect 12460 19824 12498 19858
rect 12532 19824 12570 19858
rect 12604 19824 12642 19858
rect 12676 19824 12714 19858
rect 12748 19824 12786 19858
rect 12820 19824 12858 19858
rect 12892 19824 12930 19858
rect 12964 19824 13002 19858
rect 13036 19824 13074 19858
rect 13108 19824 13146 19858
rect 13180 19824 13218 19858
rect 13252 19824 13290 19858
rect 13324 19824 13362 19858
rect 13396 19824 13434 19858
rect 13468 19824 13506 19858
rect 13540 19824 13578 19858
rect 13612 19824 13650 19858
rect 13684 19824 13722 19858
rect 13756 19824 13794 19858
rect 13828 19824 13866 19858
rect 13900 19824 13938 19858
rect 13972 19824 14010 19858
rect 14044 19824 14082 19858
rect 14116 19824 14154 19858
rect 14188 19824 14226 19858
rect 14260 19824 14298 19858
rect 14332 19824 14370 19858
rect 14404 19824 14442 19858
rect 14476 19824 14514 19858
rect 14548 19824 14586 19858
rect 14620 19824 14658 19858
rect 14692 19824 14730 19858
rect 14873 19844 14874 19858
rect 14939 19844 14971 19864
rect 14764 19830 14802 19844
rect 14836 19830 14874 19844
rect 14908 19830 14971 19844
tri 14971 19835 15000 19864 nw
rect 14873 19824 14874 19830
rect 8857 19776 8872 19824
rect 8924 19776 8939 19824
rect 8991 19776 9006 19824
rect 9058 19776 9073 19824
rect 9125 19776 9140 19824
rect 9192 19776 9207 19824
rect 9259 19778 14755 19824
rect 14807 19778 14821 19824
rect 14873 19778 14887 19824
rect 14939 19778 14971 19830
rect 9259 19776 14971 19778
rect -29 19772 14971 19776
rect -29 19738 70 19772
rect 104 19738 143 19772
rect 177 19760 216 19772
rect 250 19760 289 19772
rect 323 19760 362 19772
rect 396 19760 435 19772
rect 469 19760 508 19772
rect 542 19760 581 19772
rect 615 19760 654 19772
rect 688 19760 727 19772
rect 761 19760 800 19772
rect 834 19760 873 19772
rect 907 19760 946 19772
rect 980 19760 1019 19772
rect 1053 19760 1092 19772
rect 1126 19760 1165 19772
rect 1199 19760 1238 19772
rect 177 19738 201 19760
rect -29 19708 201 19738
rect 253 19708 269 19760
rect 323 19738 337 19760
rect 396 19738 404 19760
rect 469 19738 471 19760
rect 724 19738 727 19760
rect 791 19738 800 19760
rect 321 19708 337 19738
rect 389 19708 404 19738
rect 456 19708 471 19738
rect 523 19708 538 19738
rect 590 19708 605 19738
rect 657 19708 672 19738
rect 724 19708 739 19738
rect 791 19708 806 19738
rect 858 19708 873 19760
rect 925 19708 940 19760
rect 992 19708 1007 19760
rect 1059 19708 1074 19760
rect 1126 19708 1141 19760
rect 1199 19738 1208 19760
rect 1272 19738 1311 19772
rect 1345 19738 1384 19772
rect 1418 19738 1457 19772
rect 1491 19738 1530 19772
rect 1564 19738 1603 19772
rect 1637 19738 1676 19772
rect 1710 19738 1749 19772
rect 1783 19738 1822 19772
rect 1856 19738 1895 19772
rect 1929 19738 1968 19772
rect 2002 19738 2041 19772
rect 2075 19738 2114 19772
rect 2148 19738 2187 19772
rect 2221 19738 2260 19772
rect 2294 19738 2333 19772
rect 2367 19738 2406 19772
rect 2440 19738 2479 19772
rect 2513 19738 2552 19772
rect 2586 19738 2625 19772
rect 2659 19738 2698 19772
rect 2732 19738 2771 19772
rect 2805 19738 2844 19772
rect 2878 19738 2917 19772
rect 2951 19738 2990 19772
rect 3024 19738 3063 19772
rect 3097 19738 3136 19772
rect 3170 19738 3209 19772
rect 3243 19738 3282 19772
rect 3316 19738 3354 19772
rect 3388 19738 3426 19772
rect 3460 19738 3498 19772
rect 3532 19738 3570 19772
rect 3604 19738 3642 19772
rect 3676 19738 3714 19772
rect 3748 19738 3786 19772
rect 3820 19738 3858 19772
rect 3892 19738 3930 19772
rect 3964 19738 4002 19772
rect 4036 19738 4074 19772
rect 4108 19738 4146 19772
rect 4180 19738 4218 19772
rect 4252 19738 4290 19772
rect 4324 19738 4362 19772
rect 4396 19738 4434 19772
rect 4468 19738 4506 19772
rect 4540 19738 4578 19772
rect 4612 19738 4650 19772
rect 4684 19738 4722 19772
rect 4756 19738 4794 19772
rect 4828 19738 4866 19772
rect 4900 19738 4938 19772
rect 4972 19738 5010 19772
rect 5044 19738 5082 19772
rect 5116 19738 5154 19772
rect 5188 19738 5226 19772
rect 5260 19738 5298 19772
rect 5332 19738 5370 19772
rect 5404 19738 5442 19772
rect 5476 19738 5514 19772
rect 5548 19738 5586 19772
rect 5620 19738 5658 19772
rect 5692 19738 5730 19772
rect 5764 19738 5802 19772
rect 5836 19738 5874 19772
rect 5908 19738 5946 19772
rect 5980 19738 6018 19772
rect 6052 19738 6090 19772
rect 6124 19738 6162 19772
rect 6196 19738 6234 19772
rect 6268 19738 6306 19772
rect 6340 19738 6378 19772
rect 6412 19738 6450 19772
rect 6484 19738 6522 19772
rect 6556 19738 6594 19772
rect 6628 19738 6666 19772
rect 6700 19738 6738 19772
rect 6772 19738 6810 19772
rect 6844 19738 6882 19772
rect 6916 19738 6954 19772
rect 6988 19738 7026 19772
rect 7060 19738 7098 19772
rect 7132 19738 7170 19772
rect 7204 19738 7242 19772
rect 7276 19738 7314 19772
rect 7348 19738 7386 19772
rect 7420 19738 7458 19772
rect 7492 19738 7530 19772
rect 7564 19738 7602 19772
rect 7636 19738 7674 19772
rect 7708 19738 7746 19772
rect 7780 19738 7818 19772
rect 7852 19738 7890 19772
rect 7924 19738 7962 19772
rect 7996 19738 8034 19772
rect 8068 19738 8106 19772
rect 8140 19738 8178 19772
rect 8212 19760 8250 19772
rect 8284 19760 8322 19772
rect 8356 19760 8394 19772
rect 8428 19760 8466 19772
rect 8500 19760 8538 19772
rect 8572 19760 8610 19772
rect 8644 19760 8682 19772
rect 8716 19760 8754 19772
rect 8788 19760 8826 19772
rect 8860 19760 8898 19772
rect 8932 19760 8970 19772
rect 9004 19760 9042 19772
rect 9076 19760 9114 19772
rect 9148 19760 9186 19772
rect 9220 19760 9258 19772
rect 8320 19738 8322 19760
rect 8388 19738 8394 19760
rect 8455 19738 8466 19760
rect 1193 19708 1208 19738
rect 1260 19708 8200 19738
rect 8252 19708 8268 19738
rect 8320 19708 8336 19738
rect 8388 19708 8403 19738
rect 8455 19708 8470 19738
rect 8522 19708 8537 19760
rect 8589 19708 8604 19760
rect 8656 19708 8671 19760
rect 8723 19708 8738 19760
rect 8790 19708 8805 19760
rect 8860 19738 8872 19760
rect 8932 19738 8939 19760
rect 9004 19738 9006 19760
rect 9292 19738 9330 19772
rect 9364 19738 9402 19772
rect 9436 19738 9474 19772
rect 9508 19738 9546 19772
rect 9580 19738 9618 19772
rect 9652 19738 9690 19772
rect 9724 19738 9762 19772
rect 9796 19738 9834 19772
rect 9868 19738 9906 19772
rect 9940 19738 9978 19772
rect 10012 19738 10050 19772
rect 10084 19738 10122 19772
rect 10156 19738 10194 19772
rect 10228 19738 10266 19772
rect 10300 19738 10338 19772
rect 10372 19738 10410 19772
rect 10444 19738 10482 19772
rect 10516 19738 10554 19772
rect 10588 19738 10626 19772
rect 10660 19738 10698 19772
rect 10732 19738 10770 19772
rect 10804 19738 10842 19772
rect 10876 19738 10914 19772
rect 10948 19738 10986 19772
rect 11020 19738 11058 19772
rect 11092 19738 11130 19772
rect 11164 19738 11202 19772
rect 11236 19738 11274 19772
rect 11308 19738 11346 19772
rect 11380 19738 11418 19772
rect 11452 19738 11490 19772
rect 11524 19738 11562 19772
rect 11596 19738 11634 19772
rect 11668 19738 11706 19772
rect 11740 19738 11778 19772
rect 11812 19738 11850 19772
rect 11884 19738 11922 19772
rect 11956 19738 11994 19772
rect 12028 19738 12066 19772
rect 12100 19738 12138 19772
rect 12172 19738 12210 19772
rect 12244 19738 12282 19772
rect 12316 19738 12354 19772
rect 12388 19738 12426 19772
rect 12460 19738 12498 19772
rect 12532 19738 12570 19772
rect 12604 19738 12642 19772
rect 12676 19738 12714 19772
rect 12748 19738 12786 19772
rect 12820 19738 12858 19772
rect 12892 19738 12930 19772
rect 12964 19738 13002 19772
rect 13036 19738 13074 19772
rect 13108 19738 13146 19772
rect 13180 19738 13218 19772
rect 13252 19738 13290 19772
rect 13324 19738 13362 19772
rect 13396 19738 13434 19772
rect 13468 19738 13506 19772
rect 13540 19738 13578 19772
rect 13612 19738 13650 19772
rect 13684 19738 13722 19772
rect 13756 19738 13794 19772
rect 13828 19738 13866 19772
rect 13900 19738 13938 19772
rect 13972 19738 14010 19772
rect 14044 19738 14082 19772
rect 14116 19738 14154 19772
rect 14188 19738 14226 19772
rect 14260 19738 14298 19772
rect 14332 19738 14370 19772
rect 14404 19738 14442 19772
rect 14476 19738 14514 19772
rect 14548 19738 14586 19772
rect 14620 19738 14658 19772
rect 14692 19738 14730 19772
rect 14764 19764 14802 19772
rect 14836 19764 14874 19772
rect 14908 19764 14971 19772
rect 14873 19738 14874 19764
rect 8857 19708 8872 19738
rect 8924 19708 8939 19738
rect 8991 19708 9006 19738
rect 9058 19708 9073 19738
rect 9125 19708 9140 19738
rect 9192 19708 9207 19738
rect 9259 19712 14755 19738
rect 14807 19712 14821 19738
rect 14873 19712 14887 19738
rect 14939 19712 14971 19764
rect 9259 19708 14971 19712
rect -29 19698 14971 19708
rect -29 19692 14755 19698
rect -29 19686 201 19692
rect -29 19652 70 19686
rect 104 19652 143 19686
rect 177 19652 201 19686
rect -29 19640 201 19652
rect 253 19640 269 19692
rect 321 19686 337 19692
rect 389 19686 404 19692
rect 456 19686 471 19692
rect 523 19686 538 19692
rect 590 19686 605 19692
rect 657 19686 672 19692
rect 724 19686 739 19692
rect 791 19686 806 19692
rect 323 19652 337 19686
rect 396 19652 404 19686
rect 469 19652 471 19686
rect 724 19652 727 19686
rect 791 19652 800 19686
rect 321 19640 337 19652
rect 389 19640 404 19652
rect 456 19640 471 19652
rect 523 19640 538 19652
rect 590 19640 605 19652
rect 657 19640 672 19652
rect 724 19640 739 19652
rect 791 19640 806 19652
rect 858 19640 873 19692
rect 925 19640 940 19692
rect 992 19640 1007 19692
rect 1059 19640 1074 19692
rect 1126 19640 1141 19692
rect 1193 19686 1208 19692
rect 1260 19686 8200 19692
rect 8252 19686 8268 19692
rect 8320 19686 8336 19692
rect 8388 19686 8403 19692
rect 8455 19686 8470 19692
rect 1199 19652 1208 19686
rect 1272 19652 1311 19686
rect 1345 19652 1384 19686
rect 1418 19652 1457 19686
rect 1491 19652 1530 19686
rect 1564 19652 1603 19686
rect 1637 19652 1676 19686
rect 1710 19652 1749 19686
rect 1783 19652 1822 19686
rect 1856 19652 1895 19686
rect 1929 19652 1968 19686
rect 2002 19652 2041 19686
rect 2075 19652 2114 19686
rect 2148 19652 2187 19686
rect 2221 19652 2260 19686
rect 2294 19652 2333 19686
rect 2367 19652 2406 19686
rect 2440 19652 2479 19686
rect 2513 19652 2552 19686
rect 2586 19652 2625 19686
rect 2659 19652 2698 19686
rect 2732 19652 2771 19686
rect 2805 19652 2844 19686
rect 2878 19652 2917 19686
rect 2951 19652 2990 19686
rect 3024 19652 3063 19686
rect 3097 19652 3136 19686
rect 3170 19652 3209 19686
rect 3243 19652 3282 19686
rect 3316 19652 3354 19686
rect 3388 19652 3426 19686
rect 3460 19652 3498 19686
rect 3532 19652 3570 19686
rect 3604 19652 3642 19686
rect 3676 19652 3714 19686
rect 3748 19652 3786 19686
rect 3820 19652 3858 19686
rect 3892 19652 3930 19686
rect 3964 19652 4002 19686
rect 4036 19652 4074 19686
rect 4108 19652 4146 19686
rect 4180 19652 4218 19686
rect 4252 19652 4290 19686
rect 4324 19652 4362 19686
rect 4396 19652 4434 19686
rect 4468 19652 4506 19686
rect 4540 19652 4578 19686
rect 4612 19652 4650 19686
rect 4684 19652 4722 19686
rect 4756 19652 4794 19686
rect 4828 19652 4866 19686
rect 4900 19652 4938 19686
rect 4972 19652 5010 19686
rect 5044 19652 5082 19686
rect 5116 19652 5154 19686
rect 5188 19652 5226 19686
rect 5260 19652 5298 19686
rect 5332 19652 5370 19686
rect 5404 19652 5442 19686
rect 5476 19652 5514 19686
rect 5548 19652 5586 19686
rect 5620 19652 5658 19686
rect 5692 19652 5730 19686
rect 5764 19652 5802 19686
rect 5836 19652 5874 19686
rect 5908 19652 5946 19686
rect 5980 19652 6018 19686
rect 6052 19652 6090 19686
rect 6124 19652 6162 19686
rect 6196 19652 6234 19686
rect 6268 19652 6306 19686
rect 6340 19652 6378 19686
rect 6412 19652 6450 19686
rect 6484 19652 6522 19686
rect 6556 19652 6594 19686
rect 6628 19652 6666 19686
rect 6700 19652 6738 19686
rect 6772 19652 6810 19686
rect 6844 19652 6882 19686
rect 6916 19652 6954 19686
rect 6988 19652 7026 19686
rect 7060 19652 7098 19686
rect 7132 19652 7170 19686
rect 7204 19652 7242 19686
rect 7276 19652 7314 19686
rect 7348 19652 7386 19686
rect 7420 19652 7458 19686
rect 7492 19652 7530 19686
rect 7564 19652 7602 19686
rect 7636 19652 7674 19686
rect 7708 19652 7746 19686
rect 7780 19652 7818 19686
rect 7852 19652 7890 19686
rect 7924 19652 7962 19686
rect 7996 19652 8034 19686
rect 8068 19652 8106 19686
rect 8140 19652 8178 19686
rect 8320 19652 8322 19686
rect 8388 19652 8394 19686
rect 8455 19652 8466 19686
rect 1193 19640 1208 19652
rect 1260 19640 8200 19652
rect 8252 19640 8268 19652
rect 8320 19640 8336 19652
rect 8388 19640 8403 19652
rect 8455 19640 8470 19652
rect 8522 19640 8537 19692
rect 8589 19640 8604 19692
rect 8656 19640 8671 19692
rect 8723 19640 8738 19692
rect 8790 19640 8805 19692
rect 8857 19686 8872 19692
rect 8924 19686 8939 19692
rect 8991 19686 9006 19692
rect 9058 19686 9073 19692
rect 9125 19686 9140 19692
rect 9192 19686 9207 19692
rect 9259 19686 14755 19692
rect 14807 19686 14821 19698
rect 14873 19686 14887 19698
rect 8860 19652 8872 19686
rect 8932 19652 8939 19686
rect 9004 19652 9006 19686
rect 9292 19652 9330 19686
rect 9364 19652 9402 19686
rect 9436 19652 9474 19686
rect 9508 19652 9546 19686
rect 9580 19652 9618 19686
rect 9652 19652 9690 19686
rect 9724 19652 9762 19686
rect 9796 19652 9834 19686
rect 9868 19652 9906 19686
rect 9940 19652 9978 19686
rect 10012 19652 10050 19686
rect 10084 19652 10122 19686
rect 10156 19652 10194 19686
rect 10228 19652 10266 19686
rect 10300 19652 10338 19686
rect 10372 19652 10410 19686
rect 10444 19652 10482 19686
rect 10516 19652 10554 19686
rect 10588 19652 10626 19686
rect 10660 19652 10698 19686
rect 10732 19652 10770 19686
rect 10804 19652 10842 19686
rect 10876 19652 10914 19686
rect 10948 19652 10986 19686
rect 11020 19652 11058 19686
rect 11092 19652 11130 19686
rect 11164 19652 11202 19686
rect 11236 19652 11274 19686
rect 11308 19652 11346 19686
rect 11380 19652 11418 19686
rect 11452 19652 11490 19686
rect 11524 19652 11562 19686
rect 11596 19652 11634 19686
rect 11668 19652 11706 19686
rect 11740 19652 11778 19686
rect 11812 19652 11850 19686
rect 11884 19652 11922 19686
rect 11956 19652 11994 19686
rect 12028 19652 12066 19686
rect 12100 19652 12138 19686
rect 12172 19652 12210 19686
rect 12244 19652 12282 19686
rect 12316 19652 12354 19686
rect 12388 19652 12426 19686
rect 12460 19652 12498 19686
rect 12532 19652 12570 19686
rect 12604 19652 12642 19686
rect 12676 19652 12714 19686
rect 12748 19652 12786 19686
rect 12820 19652 12858 19686
rect 12892 19652 12930 19686
rect 12964 19652 13002 19686
rect 13036 19652 13074 19686
rect 13108 19652 13146 19686
rect 13180 19652 13218 19686
rect 13252 19652 13290 19686
rect 13324 19652 13362 19686
rect 13396 19652 13434 19686
rect 13468 19652 13506 19686
rect 13540 19652 13578 19686
rect 13612 19652 13650 19686
rect 13684 19652 13722 19686
rect 13756 19652 13794 19686
rect 13828 19652 13866 19686
rect 13900 19652 13938 19686
rect 13972 19652 14010 19686
rect 14044 19652 14082 19686
rect 14116 19652 14154 19686
rect 14188 19652 14226 19686
rect 14260 19652 14298 19686
rect 14332 19652 14370 19686
rect 14404 19652 14442 19686
rect 14476 19652 14514 19686
rect 14548 19652 14586 19686
rect 14620 19652 14658 19686
rect 14692 19652 14730 19686
rect 14873 19652 14874 19686
rect 8857 19640 8872 19652
rect 8924 19640 8939 19652
rect 8991 19640 9006 19652
rect 9058 19640 9073 19652
rect 9125 19640 9140 19652
rect 9192 19640 9207 19652
rect 9259 19646 14755 19652
rect 14807 19646 14821 19652
rect 14873 19646 14887 19652
rect 14939 19646 14971 19698
rect 9259 19640 14971 19646
rect -29 19632 14971 19640
rect -29 19624 14755 19632
rect -29 19600 201 19624
rect -29 19566 70 19600
rect 104 19566 143 19600
rect 177 19572 201 19600
rect 253 19572 269 19624
rect 321 19600 337 19624
rect 389 19600 404 19624
rect 456 19600 471 19624
rect 523 19600 538 19624
rect 590 19600 605 19624
rect 657 19600 672 19624
rect 724 19600 739 19624
rect 791 19600 806 19624
rect 323 19572 337 19600
rect 396 19572 404 19600
rect 469 19572 471 19600
rect 724 19572 727 19600
rect 791 19572 800 19600
rect 858 19572 873 19624
rect 925 19572 940 19624
rect 992 19572 1007 19624
rect 1059 19572 1074 19624
rect 1126 19572 1141 19624
rect 1193 19600 1208 19624
rect 1260 19600 8200 19624
rect 8252 19600 8268 19624
rect 8320 19600 8336 19624
rect 8388 19600 8403 19624
rect 8455 19600 8470 19624
rect 1199 19572 1208 19600
rect 177 19566 216 19572
rect 250 19566 289 19572
rect 323 19566 362 19572
rect 396 19566 435 19572
rect 469 19566 508 19572
rect 542 19566 581 19572
rect 615 19566 654 19572
rect 688 19566 727 19572
rect 761 19566 800 19572
rect 834 19566 873 19572
rect 907 19566 946 19572
rect 980 19566 1019 19572
rect 1053 19566 1092 19572
rect 1126 19566 1165 19572
rect 1199 19566 1238 19572
rect 1272 19566 1311 19600
rect 1345 19566 1384 19600
rect 1418 19566 1457 19600
rect 1491 19566 1530 19600
rect 1564 19566 1603 19600
rect 1637 19566 1676 19600
rect 1710 19566 1749 19600
rect 1783 19566 1822 19600
rect 1856 19566 1895 19600
rect 1929 19566 1968 19600
rect 2002 19566 2041 19600
rect 2075 19566 2114 19600
rect 2148 19566 2187 19600
rect 2221 19566 2260 19600
rect 2294 19566 2333 19600
rect 2367 19566 2406 19600
rect 2440 19566 2479 19600
rect 2513 19566 2552 19600
rect 2586 19566 2625 19600
rect 2659 19566 2698 19600
rect 2732 19566 2771 19600
rect 2805 19566 2844 19600
rect 2878 19566 2917 19600
rect 2951 19566 2990 19600
rect 3024 19566 3063 19600
rect 3097 19566 3136 19600
rect 3170 19566 3209 19600
rect 3243 19566 3282 19600
rect 3316 19566 3354 19600
rect 3388 19566 3426 19600
rect 3460 19566 3498 19600
rect 3532 19566 3570 19600
rect 3604 19566 3642 19600
rect 3676 19566 3714 19600
rect 3748 19566 3786 19600
rect 3820 19566 3858 19600
rect 3892 19566 3930 19600
rect 3964 19566 4002 19600
rect 4036 19566 4074 19600
rect 4108 19566 4146 19600
rect 4180 19566 4218 19600
rect 4252 19566 4290 19600
rect 4324 19566 4362 19600
rect 4396 19566 4434 19600
rect 4468 19566 4506 19600
rect 4540 19566 4578 19600
rect 4612 19566 4650 19600
rect 4684 19566 4722 19600
rect 4756 19566 4794 19600
rect 4828 19566 4866 19600
rect 4900 19566 4938 19600
rect 4972 19566 5010 19600
rect 5044 19566 5082 19600
rect 5116 19566 5154 19600
rect 5188 19566 5226 19600
rect 5260 19566 5298 19600
rect 5332 19566 5370 19600
rect 5404 19566 5442 19600
rect 5476 19566 5514 19600
rect 5548 19566 5586 19600
rect 5620 19566 5658 19600
rect 5692 19566 5730 19600
rect 5764 19566 5802 19600
rect 5836 19566 5874 19600
rect 5908 19566 5946 19600
rect 5980 19566 6018 19600
rect 6052 19566 6090 19600
rect 6124 19566 6162 19600
rect 6196 19566 6234 19600
rect 6268 19566 6306 19600
rect 6340 19566 6378 19600
rect 6412 19566 6450 19600
rect 6484 19566 6522 19600
rect 6556 19566 6594 19600
rect 6628 19566 6666 19600
rect 6700 19566 6738 19600
rect 6772 19566 6810 19600
rect 6844 19566 6882 19600
rect 6916 19566 6954 19600
rect 6988 19566 7026 19600
rect 7060 19566 7098 19600
rect 7132 19566 7170 19600
rect 7204 19566 7242 19600
rect 7276 19566 7314 19600
rect 7348 19566 7386 19600
rect 7420 19566 7458 19600
rect 7492 19566 7530 19600
rect 7564 19566 7602 19600
rect 7636 19566 7674 19600
rect 7708 19566 7746 19600
rect 7780 19566 7818 19600
rect 7852 19566 7890 19600
rect 7924 19566 7962 19600
rect 7996 19566 8034 19600
rect 8068 19566 8106 19600
rect 8140 19566 8178 19600
rect 8320 19572 8322 19600
rect 8388 19572 8394 19600
rect 8455 19572 8466 19600
rect 8522 19572 8537 19624
rect 8589 19572 8604 19624
rect 8656 19572 8671 19624
rect 8723 19572 8738 19624
rect 8790 19572 8805 19624
rect 8857 19600 8872 19624
rect 8924 19600 8939 19624
rect 8991 19600 9006 19624
rect 9058 19600 9073 19624
rect 9125 19600 9140 19624
rect 9192 19600 9207 19624
rect 9259 19600 14755 19624
rect 14807 19600 14821 19632
rect 14873 19600 14887 19632
rect 8860 19572 8872 19600
rect 8932 19572 8939 19600
rect 9004 19572 9006 19600
rect 8212 19566 8250 19572
rect 8284 19566 8322 19572
rect 8356 19566 8394 19572
rect 8428 19566 8466 19572
rect 8500 19566 8538 19572
rect 8572 19566 8610 19572
rect 8644 19566 8682 19572
rect 8716 19566 8754 19572
rect 8788 19566 8826 19572
rect 8860 19566 8898 19572
rect 8932 19566 8970 19572
rect 9004 19566 9042 19572
rect 9076 19566 9114 19572
rect 9148 19566 9186 19572
rect 9220 19566 9258 19572
rect 9292 19566 9330 19600
rect 9364 19566 9402 19600
rect 9436 19566 9474 19600
rect 9508 19566 9546 19600
rect 9580 19566 9618 19600
rect 9652 19566 9690 19600
rect 9724 19566 9762 19600
rect 9796 19566 9834 19600
rect 9868 19566 9906 19600
rect 9940 19566 9978 19600
rect 10012 19566 10050 19600
rect 10084 19566 10122 19600
rect 10156 19566 10194 19600
rect 10228 19566 10266 19600
rect 10300 19566 10338 19600
rect 10372 19566 10410 19600
rect 10444 19566 10482 19600
rect 10516 19566 10554 19600
rect 10588 19566 10626 19600
rect 10660 19566 10698 19600
rect 10732 19566 10770 19600
rect 10804 19566 10842 19600
rect 10876 19566 10914 19600
rect 10948 19566 10986 19600
rect 11020 19566 11058 19600
rect 11092 19566 11130 19600
rect 11164 19566 11202 19600
rect 11236 19566 11274 19600
rect 11308 19566 11346 19600
rect 11380 19566 11418 19600
rect 11452 19566 11490 19600
rect 11524 19566 11562 19600
rect 11596 19566 11634 19600
rect 11668 19566 11706 19600
rect 11740 19566 11778 19600
rect 11812 19566 11850 19600
rect 11884 19566 11922 19600
rect 11956 19566 11994 19600
rect 12028 19566 12066 19600
rect 12100 19566 12138 19600
rect 12172 19566 12210 19600
rect 12244 19566 12282 19600
rect 12316 19566 12354 19600
rect 12388 19566 12426 19600
rect 12460 19566 12498 19600
rect 12532 19566 12570 19600
rect 12604 19566 12642 19600
rect 12676 19566 12714 19600
rect 12748 19566 12786 19600
rect 12820 19566 12858 19600
rect 12892 19566 12930 19600
rect 12964 19566 13002 19600
rect 13036 19566 13074 19600
rect 13108 19566 13146 19600
rect 13180 19566 13218 19600
rect 13252 19566 13290 19600
rect 13324 19566 13362 19600
rect 13396 19566 13434 19600
rect 13468 19566 13506 19600
rect 13540 19566 13578 19600
rect 13612 19566 13650 19600
rect 13684 19566 13722 19600
rect 13756 19566 13794 19600
rect 13828 19566 13866 19600
rect 13900 19566 13938 19600
rect 13972 19566 14010 19600
rect 14044 19566 14082 19600
rect 14116 19566 14154 19600
rect 14188 19566 14226 19600
rect 14260 19566 14298 19600
rect 14332 19566 14370 19600
rect 14404 19566 14442 19600
rect 14476 19566 14514 19600
rect 14548 19566 14586 19600
rect 14620 19566 14658 19600
rect 14692 19566 14730 19600
rect 14873 19580 14874 19600
rect 14939 19580 14971 19632
rect 14764 19566 14802 19580
rect 14836 19566 14874 19580
rect 14908 19566 14971 19580
rect -29 19560 14971 19566
rect 12610 18765 12616 18817
rect 12668 18765 12682 18817
rect 12734 18765 12740 18817
rect 12610 18685 12616 18737
rect 12668 18685 12682 18737
rect 12734 18685 12740 18737
rect 195 18387 14772 18393
rect 195 18335 201 18387
rect 253 18335 269 18387
rect 321 18335 337 18387
rect 389 18335 404 18387
rect 456 18382 471 18387
rect 523 18382 538 18387
rect 590 18382 605 18387
rect 657 18382 672 18387
rect 724 18382 739 18387
rect 791 18382 806 18387
rect 858 18382 873 18387
rect 925 18382 940 18387
rect 462 18348 471 18382
rect 535 18348 538 18382
rect 791 18348 793 18382
rect 858 18348 866 18382
rect 925 18348 939 18382
rect 456 18335 471 18348
rect 523 18335 538 18348
rect 590 18335 605 18348
rect 657 18335 672 18348
rect 724 18335 739 18348
rect 791 18335 806 18348
rect 858 18335 873 18348
rect 925 18335 940 18348
rect 992 18335 1007 18387
rect 1059 18335 1074 18387
rect 1126 18335 1141 18387
rect 1193 18335 1208 18387
rect 1260 18382 14772 18387
rect 1265 18348 1304 18382
rect 1338 18348 1377 18382
rect 1411 18348 1450 18382
rect 1484 18348 1523 18382
rect 1557 18348 1596 18382
rect 1630 18348 1669 18382
rect 1703 18348 1742 18382
rect 1776 18348 1815 18382
rect 1849 18348 1888 18382
rect 1922 18348 1961 18382
rect 1995 18348 2034 18382
rect 2068 18348 2107 18382
rect 2141 18348 2180 18382
rect 2214 18348 2253 18382
rect 2287 18348 2326 18382
rect 2360 18348 2399 18382
rect 2433 18348 2472 18382
rect 2506 18348 2545 18382
rect 2579 18348 2618 18382
rect 2652 18348 2691 18382
rect 2725 18348 2764 18382
rect 2798 18348 2837 18382
rect 2871 18348 2910 18382
rect 2944 18348 2983 18382
rect 3017 18348 3056 18382
rect 3090 18348 3129 18382
rect 3163 18348 3202 18382
rect 3236 18348 3275 18382
rect 3309 18348 3348 18382
rect 3382 18348 3421 18382
rect 3455 18348 3494 18382
rect 3528 18348 3566 18382
rect 3600 18348 3638 18382
rect 3672 18348 3710 18382
rect 3744 18348 3782 18382
rect 3816 18348 3854 18382
rect 3888 18348 3926 18382
rect 3960 18348 3998 18382
rect 4032 18348 4070 18382
rect 4104 18348 4142 18382
rect 4176 18348 4214 18382
rect 4248 18348 4286 18382
rect 4320 18348 4358 18382
rect 4392 18348 4430 18382
rect 4464 18348 4502 18382
rect 4536 18348 4574 18382
rect 4608 18348 4646 18382
rect 4680 18348 4718 18382
rect 4752 18348 4790 18382
rect 4824 18348 4862 18382
rect 4896 18348 4934 18382
rect 4968 18348 5006 18382
rect 5040 18348 5078 18382
rect 5112 18348 5150 18382
rect 5184 18348 5222 18382
rect 5256 18348 5294 18382
rect 5328 18348 5366 18382
rect 5400 18348 5438 18382
rect 5472 18348 5510 18382
rect 5544 18348 5582 18382
rect 5616 18348 5654 18382
rect 5688 18348 5726 18382
rect 5760 18348 5798 18382
rect 5832 18348 5870 18382
rect 5904 18348 5942 18382
rect 5976 18348 6014 18382
rect 6048 18348 6086 18382
rect 6120 18348 6158 18382
rect 6192 18348 6230 18382
rect 6264 18348 6302 18382
rect 6336 18348 6374 18382
rect 6408 18348 6446 18382
rect 6480 18348 6518 18382
rect 6552 18348 6590 18382
rect 6624 18348 6662 18382
rect 6696 18348 6734 18382
rect 6768 18348 6806 18382
rect 6840 18348 6878 18382
rect 6912 18348 6950 18382
rect 6984 18348 7022 18382
rect 7056 18348 7094 18382
rect 7128 18348 7166 18382
rect 7200 18348 7238 18382
rect 7272 18348 7310 18382
rect 7344 18348 7382 18382
rect 7416 18348 7454 18382
rect 7488 18348 7526 18382
rect 7560 18348 7598 18382
rect 7632 18348 7670 18382
rect 7704 18348 7742 18382
rect 7776 18348 7814 18382
rect 7848 18348 7886 18382
rect 7920 18348 7958 18382
rect 7992 18348 8030 18382
rect 8064 18348 8102 18382
rect 8136 18348 8174 18382
rect 8208 18348 8246 18382
rect 8280 18348 8318 18382
rect 8352 18348 8390 18382
rect 8424 18348 8462 18382
rect 8496 18348 8534 18382
rect 8568 18348 8606 18382
rect 8640 18348 8678 18382
rect 8712 18348 8750 18382
rect 8784 18348 8822 18382
rect 8856 18348 8894 18382
rect 8928 18348 8966 18382
rect 9000 18348 9038 18382
rect 9072 18348 9110 18382
rect 9144 18348 9182 18382
rect 9216 18348 9254 18382
rect 9288 18348 9326 18382
rect 9360 18348 9398 18382
rect 9432 18348 9470 18382
rect 9504 18348 9542 18382
rect 9576 18348 9614 18382
rect 9648 18348 9686 18382
rect 9720 18348 9758 18382
rect 9792 18348 9830 18382
rect 9864 18348 9902 18382
rect 9936 18348 9974 18382
rect 10008 18348 10046 18382
rect 10080 18348 10118 18382
rect 10152 18348 10190 18382
rect 10224 18348 10262 18382
rect 10296 18348 10334 18382
rect 10368 18348 10406 18382
rect 10440 18348 10478 18382
rect 10512 18348 10550 18382
rect 10584 18348 10622 18382
rect 10656 18348 10694 18382
rect 10728 18348 10766 18382
rect 10800 18348 10838 18382
rect 10872 18348 10910 18382
rect 10944 18348 10982 18382
rect 11016 18348 11054 18382
rect 11088 18348 11126 18382
rect 11160 18348 11198 18382
rect 11232 18348 11270 18382
rect 11304 18348 11342 18382
rect 11376 18348 11414 18382
rect 11448 18348 11486 18382
rect 11520 18348 11558 18382
rect 11592 18348 11630 18382
rect 11664 18348 11702 18382
rect 11736 18348 11774 18382
rect 11808 18348 11846 18382
rect 11880 18348 11918 18382
rect 11952 18348 11990 18382
rect 12024 18348 12062 18382
rect 12096 18348 12134 18382
rect 12168 18348 12206 18382
rect 12240 18348 12278 18382
rect 12312 18348 12350 18382
rect 12384 18348 12422 18382
rect 12456 18348 12494 18382
rect 12528 18348 12566 18382
rect 12600 18348 12638 18382
rect 12672 18348 12710 18382
rect 12744 18348 12782 18382
rect 12816 18348 12854 18382
rect 12888 18348 12926 18382
rect 12960 18348 12998 18382
rect 13032 18348 13070 18382
rect 13104 18348 13142 18382
rect 13176 18348 13214 18382
rect 13248 18348 13286 18382
rect 13320 18348 13358 18382
rect 13392 18348 13430 18382
rect 13464 18348 13502 18382
rect 13536 18348 13574 18382
rect 13608 18348 13646 18382
rect 13680 18348 13718 18382
rect 13752 18348 13790 18382
rect 13824 18348 13862 18382
rect 13896 18348 13934 18382
rect 13968 18348 14006 18382
rect 14040 18348 14078 18382
rect 14112 18348 14150 18382
rect 14184 18348 14222 18382
rect 14256 18348 14294 18382
rect 14328 18348 14366 18382
rect 14400 18348 14438 18382
rect 14472 18348 14510 18382
rect 14544 18348 14582 18382
rect 14616 18348 14654 18382
rect 14688 18348 14726 18382
rect 14760 18348 14772 18382
rect 1260 18335 14772 18348
rect 195 18323 14772 18335
rect 195 18271 201 18323
rect 253 18271 269 18323
rect 321 18271 337 18323
rect 389 18271 404 18323
rect 456 18306 471 18323
rect 523 18306 538 18323
rect 590 18306 605 18323
rect 657 18306 672 18323
rect 724 18306 739 18323
rect 791 18306 806 18323
rect 858 18306 873 18323
rect 925 18306 940 18323
rect 462 18272 471 18306
rect 535 18272 538 18306
rect 791 18272 793 18306
rect 858 18272 866 18306
rect 925 18272 939 18306
rect 456 18271 471 18272
rect 523 18271 538 18272
rect 590 18271 605 18272
rect 657 18271 672 18272
rect 724 18271 739 18272
rect 791 18271 806 18272
rect 858 18271 873 18272
rect 925 18271 940 18272
rect 992 18271 1007 18323
rect 1059 18271 1074 18323
rect 1126 18271 1141 18323
rect 1193 18271 1208 18323
rect 1260 18306 14772 18323
rect 1265 18272 1304 18306
rect 1338 18272 1377 18306
rect 1411 18272 1450 18306
rect 1484 18272 1523 18306
rect 1557 18272 1596 18306
rect 1630 18272 1669 18306
rect 1703 18272 1742 18306
rect 1776 18272 1815 18306
rect 1849 18272 1888 18306
rect 1922 18272 1961 18306
rect 1995 18272 2034 18306
rect 2068 18272 2107 18306
rect 2141 18272 2180 18306
rect 2214 18272 2253 18306
rect 2287 18272 2326 18306
rect 2360 18272 2399 18306
rect 2433 18272 2472 18306
rect 2506 18272 2545 18306
rect 2579 18272 2618 18306
rect 2652 18272 2691 18306
rect 2725 18272 2764 18306
rect 2798 18272 2837 18306
rect 2871 18272 2910 18306
rect 2944 18272 2983 18306
rect 3017 18272 3056 18306
rect 3090 18272 3129 18306
rect 3163 18272 3202 18306
rect 3236 18272 3275 18306
rect 3309 18272 3348 18306
rect 3382 18272 3421 18306
rect 3455 18272 3494 18306
rect 3528 18272 3566 18306
rect 3600 18272 3638 18306
rect 3672 18272 3710 18306
rect 3744 18272 3782 18306
rect 3816 18272 3854 18306
rect 3888 18272 3926 18306
rect 3960 18272 3998 18306
rect 4032 18272 4070 18306
rect 4104 18272 4142 18306
rect 4176 18272 4214 18306
rect 4248 18272 4286 18306
rect 4320 18272 4358 18306
rect 4392 18272 4430 18306
rect 4464 18272 4502 18306
rect 4536 18272 4574 18306
rect 4608 18272 4646 18306
rect 4680 18272 4718 18306
rect 4752 18272 4790 18306
rect 4824 18272 4862 18306
rect 4896 18272 4934 18306
rect 4968 18272 5006 18306
rect 5040 18272 5078 18306
rect 5112 18272 5150 18306
rect 5184 18272 5222 18306
rect 5256 18272 5294 18306
rect 5328 18272 5366 18306
rect 5400 18272 5438 18306
rect 5472 18272 5510 18306
rect 5544 18272 5582 18306
rect 5616 18272 5654 18306
rect 5688 18272 5726 18306
rect 5760 18272 5798 18306
rect 5832 18272 5870 18306
rect 5904 18272 5942 18306
rect 5976 18272 6014 18306
rect 6048 18272 6086 18306
rect 6120 18272 6158 18306
rect 6192 18272 6230 18306
rect 6264 18272 6302 18306
rect 6336 18272 6374 18306
rect 6408 18272 6446 18306
rect 6480 18272 6518 18306
rect 6552 18272 6590 18306
rect 6624 18272 6662 18306
rect 6696 18272 6734 18306
rect 6768 18272 6806 18306
rect 6840 18272 6878 18306
rect 6912 18272 6950 18306
rect 6984 18272 7022 18306
rect 7056 18272 7094 18306
rect 7128 18272 7166 18306
rect 7200 18272 7238 18306
rect 7272 18272 7310 18306
rect 7344 18272 7382 18306
rect 7416 18272 7454 18306
rect 7488 18272 7526 18306
rect 7560 18272 7598 18306
rect 7632 18272 7670 18306
rect 7704 18272 7742 18306
rect 7776 18272 7814 18306
rect 7848 18272 7886 18306
rect 7920 18272 7958 18306
rect 7992 18272 8030 18306
rect 8064 18272 8102 18306
rect 8136 18272 8174 18306
rect 8208 18272 8246 18306
rect 8280 18272 8318 18306
rect 8352 18272 8390 18306
rect 8424 18272 8462 18306
rect 8496 18272 8534 18306
rect 8568 18272 8606 18306
rect 8640 18272 8678 18306
rect 8712 18272 8750 18306
rect 8784 18272 8822 18306
rect 8856 18272 8894 18306
rect 8928 18272 8966 18306
rect 9000 18272 9038 18306
rect 9072 18272 9110 18306
rect 9144 18272 9182 18306
rect 9216 18272 9254 18306
rect 9288 18272 9326 18306
rect 9360 18272 9398 18306
rect 9432 18272 9470 18306
rect 9504 18272 9542 18306
rect 9576 18272 9614 18306
rect 9648 18272 9686 18306
rect 9720 18272 9758 18306
rect 9792 18272 9830 18306
rect 9864 18272 9902 18306
rect 9936 18272 9974 18306
rect 10008 18272 10046 18306
rect 10080 18272 10118 18306
rect 10152 18272 10190 18306
rect 10224 18272 10262 18306
rect 10296 18272 10334 18306
rect 10368 18272 10406 18306
rect 10440 18272 10478 18306
rect 10512 18272 10550 18306
rect 10584 18272 10622 18306
rect 10656 18272 10694 18306
rect 10728 18272 10766 18306
rect 10800 18272 10838 18306
rect 10872 18272 10910 18306
rect 10944 18272 10982 18306
rect 11016 18272 11054 18306
rect 11088 18272 11126 18306
rect 11160 18272 11198 18306
rect 11232 18272 11270 18306
rect 11304 18272 11342 18306
rect 11376 18272 11414 18306
rect 11448 18272 11486 18306
rect 11520 18272 11558 18306
rect 11592 18272 11630 18306
rect 11664 18272 11702 18306
rect 11736 18272 11774 18306
rect 11808 18272 11846 18306
rect 11880 18272 11918 18306
rect 11952 18272 11990 18306
rect 12024 18272 12062 18306
rect 12096 18272 12134 18306
rect 12168 18272 12206 18306
rect 12240 18272 12278 18306
rect 12312 18272 12350 18306
rect 12384 18272 12422 18306
rect 12456 18272 12494 18306
rect 12528 18272 12566 18306
rect 12600 18272 12638 18306
rect 12672 18272 12710 18306
rect 12744 18272 12782 18306
rect 12816 18272 12854 18306
rect 12888 18272 12926 18306
rect 12960 18272 12998 18306
rect 13032 18272 13070 18306
rect 13104 18272 13142 18306
rect 13176 18272 13214 18306
rect 13248 18272 13286 18306
rect 13320 18272 13358 18306
rect 13392 18272 13430 18306
rect 13464 18272 13502 18306
rect 13536 18272 13574 18306
rect 13608 18272 13646 18306
rect 13680 18272 13718 18306
rect 13752 18272 13790 18306
rect 13824 18272 13862 18306
rect 13896 18272 13934 18306
rect 13968 18272 14006 18306
rect 14040 18272 14078 18306
rect 14112 18272 14150 18306
rect 14184 18272 14222 18306
rect 14256 18272 14294 18306
rect 14328 18272 14366 18306
rect 14400 18272 14438 18306
rect 14472 18272 14510 18306
rect 14544 18272 14582 18306
rect 14616 18272 14654 18306
rect 14688 18272 14726 18306
rect 14760 18272 14772 18306
rect 1260 18271 14772 18272
rect 195 18259 14772 18271
rect 195 18207 201 18259
rect 253 18207 269 18259
rect 321 18207 337 18259
rect 389 18207 404 18259
rect 456 18230 471 18259
rect 523 18230 538 18259
rect 590 18230 605 18259
rect 657 18230 672 18259
rect 724 18230 739 18259
rect 791 18230 806 18259
rect 858 18230 873 18259
rect 925 18230 940 18259
rect 462 18207 471 18230
rect 535 18207 538 18230
rect 791 18207 793 18230
rect 858 18207 866 18230
rect 925 18207 939 18230
rect 992 18207 1007 18259
rect 1059 18207 1074 18259
rect 1126 18207 1141 18259
rect 1193 18207 1208 18259
rect 1260 18230 14772 18259
rect 195 18196 209 18207
rect 243 18196 282 18207
rect 316 18196 355 18207
rect 389 18196 428 18207
rect 462 18196 501 18207
rect 535 18196 574 18207
rect 608 18196 647 18207
rect 681 18196 720 18207
rect 754 18196 793 18207
rect 827 18196 866 18207
rect 900 18196 939 18207
rect 973 18196 1012 18207
rect 1046 18196 1085 18207
rect 1119 18196 1158 18207
rect 1192 18196 1231 18207
rect 1265 18196 1304 18230
rect 1338 18196 1377 18230
rect 1411 18196 1450 18230
rect 1484 18196 1523 18230
rect 1557 18196 1596 18230
rect 1630 18196 1669 18230
rect 1703 18196 1742 18230
rect 1776 18196 1815 18230
rect 1849 18196 1888 18230
rect 1922 18196 1961 18230
rect 1995 18196 2034 18230
rect 2068 18196 2107 18230
rect 2141 18196 2180 18230
rect 2214 18196 2253 18230
rect 2287 18196 2326 18230
rect 2360 18196 2399 18230
rect 2433 18196 2472 18230
rect 2506 18196 2545 18230
rect 2579 18196 2618 18230
rect 2652 18196 2691 18230
rect 2725 18196 2764 18230
rect 2798 18196 2837 18230
rect 2871 18196 2910 18230
rect 2944 18196 2983 18230
rect 3017 18196 3056 18230
rect 3090 18196 3129 18230
rect 3163 18196 3202 18230
rect 3236 18196 3275 18230
rect 3309 18196 3348 18230
rect 3382 18196 3421 18230
rect 3455 18196 3494 18230
rect 3528 18196 3566 18230
rect 3600 18196 3638 18230
rect 3672 18196 3710 18230
rect 3744 18196 3782 18230
rect 3816 18196 3854 18230
rect 3888 18196 3926 18230
rect 3960 18196 3998 18230
rect 4032 18196 4070 18230
rect 4104 18196 4142 18230
rect 4176 18196 4214 18230
rect 4248 18196 4286 18230
rect 4320 18196 4358 18230
rect 4392 18196 4430 18230
rect 4464 18196 4502 18230
rect 4536 18196 4574 18230
rect 4608 18196 4646 18230
rect 4680 18196 4718 18230
rect 4752 18196 4790 18230
rect 4824 18196 4862 18230
rect 4896 18196 4934 18230
rect 4968 18196 5006 18230
rect 5040 18196 5078 18230
rect 5112 18196 5150 18230
rect 5184 18196 5222 18230
rect 5256 18196 5294 18230
rect 5328 18196 5366 18230
rect 5400 18196 5438 18230
rect 5472 18196 5510 18230
rect 5544 18196 5582 18230
rect 5616 18196 5654 18230
rect 5688 18196 5726 18230
rect 5760 18196 5798 18230
rect 5832 18196 5870 18230
rect 5904 18196 5942 18230
rect 5976 18196 6014 18230
rect 6048 18196 6086 18230
rect 6120 18196 6158 18230
rect 6192 18196 6230 18230
rect 6264 18196 6302 18230
rect 6336 18196 6374 18230
rect 6408 18196 6446 18230
rect 6480 18196 6518 18230
rect 6552 18196 6590 18230
rect 6624 18196 6662 18230
rect 6696 18196 6734 18230
rect 6768 18196 6806 18230
rect 6840 18196 6878 18230
rect 6912 18196 6950 18230
rect 6984 18196 7022 18230
rect 7056 18196 7094 18230
rect 7128 18196 7166 18230
rect 7200 18196 7238 18230
rect 7272 18196 7310 18230
rect 7344 18196 7382 18230
rect 7416 18196 7454 18230
rect 7488 18196 7526 18230
rect 7560 18196 7598 18230
rect 7632 18196 7670 18230
rect 7704 18196 7742 18230
rect 7776 18196 7814 18230
rect 7848 18196 7886 18230
rect 7920 18196 7958 18230
rect 7992 18196 8030 18230
rect 8064 18196 8102 18230
rect 8136 18196 8174 18230
rect 8208 18196 8246 18230
rect 8280 18196 8318 18230
rect 8352 18196 8390 18230
rect 8424 18196 8462 18230
rect 8496 18196 8534 18230
rect 8568 18196 8606 18230
rect 8640 18196 8678 18230
rect 8712 18196 8750 18230
rect 8784 18196 8822 18230
rect 8856 18196 8894 18230
rect 8928 18196 8966 18230
rect 9000 18196 9038 18230
rect 9072 18196 9110 18230
rect 9144 18196 9182 18230
rect 9216 18196 9254 18230
rect 9288 18196 9326 18230
rect 9360 18196 9398 18230
rect 9432 18196 9470 18230
rect 9504 18196 9542 18230
rect 9576 18196 9614 18230
rect 9648 18196 9686 18230
rect 9720 18196 9758 18230
rect 9792 18196 9830 18230
rect 9864 18196 9902 18230
rect 9936 18196 9974 18230
rect 10008 18196 10046 18230
rect 10080 18196 10118 18230
rect 10152 18196 10190 18230
rect 10224 18196 10262 18230
rect 10296 18196 10334 18230
rect 10368 18196 10406 18230
rect 10440 18196 10478 18230
rect 10512 18196 10550 18230
rect 10584 18196 10622 18230
rect 10656 18196 10694 18230
rect 10728 18196 10766 18230
rect 10800 18196 10838 18230
rect 10872 18196 10910 18230
rect 10944 18196 10982 18230
rect 11016 18196 11054 18230
rect 11088 18196 11126 18230
rect 11160 18196 11198 18230
rect 11232 18196 11270 18230
rect 11304 18196 11342 18230
rect 11376 18196 11414 18230
rect 11448 18196 11486 18230
rect 11520 18196 11558 18230
rect 11592 18196 11630 18230
rect 11664 18196 11702 18230
rect 11736 18196 11774 18230
rect 11808 18196 11846 18230
rect 11880 18196 11918 18230
rect 11952 18196 11990 18230
rect 12024 18196 12062 18230
rect 12096 18196 12134 18230
rect 12168 18196 12206 18230
rect 12240 18196 12278 18230
rect 12312 18196 12350 18230
rect 12384 18196 12422 18230
rect 12456 18196 12494 18230
rect 12528 18196 12566 18230
rect 12600 18196 12638 18230
rect 12672 18196 12710 18230
rect 12744 18196 12782 18230
rect 12816 18196 12854 18230
rect 12888 18196 12926 18230
rect 12960 18196 12998 18230
rect 13032 18196 13070 18230
rect 13104 18196 13142 18230
rect 13176 18196 13214 18230
rect 13248 18196 13286 18230
rect 13320 18196 13358 18230
rect 13392 18196 13430 18230
rect 13464 18196 13502 18230
rect 13536 18196 13574 18230
rect 13608 18196 13646 18230
rect 13680 18196 13718 18230
rect 13752 18196 13790 18230
rect 13824 18196 13862 18230
rect 13896 18196 13934 18230
rect 13968 18196 14006 18230
rect 14040 18196 14078 18230
rect 14112 18196 14150 18230
rect 14184 18196 14222 18230
rect 14256 18196 14294 18230
rect 14328 18196 14366 18230
rect 14400 18196 14438 18230
rect 14472 18196 14510 18230
rect 14544 18196 14582 18230
rect 14616 18196 14654 18230
rect 14688 18196 14726 18230
rect 14760 18196 14772 18230
rect 195 18195 14772 18196
rect 195 18143 201 18195
rect 253 18143 269 18195
rect 321 18143 337 18195
rect 389 18143 404 18195
rect 456 18154 471 18195
rect 523 18154 538 18195
rect 590 18154 605 18195
rect 657 18154 672 18195
rect 724 18154 739 18195
rect 791 18154 806 18195
rect 858 18154 873 18195
rect 925 18154 940 18195
rect 462 18143 471 18154
rect 535 18143 538 18154
rect 791 18143 793 18154
rect 858 18143 866 18154
rect 925 18143 939 18154
rect 992 18143 1007 18195
rect 1059 18143 1074 18195
rect 1126 18143 1141 18195
rect 1193 18143 1208 18195
rect 1260 18154 14772 18195
rect 195 18131 209 18143
rect 243 18131 282 18143
rect 316 18131 355 18143
rect 389 18131 428 18143
rect 462 18131 501 18143
rect 535 18131 574 18143
rect 608 18131 647 18143
rect 681 18131 720 18143
rect 754 18131 793 18143
rect 827 18131 866 18143
rect 900 18131 939 18143
rect 973 18131 1012 18143
rect 1046 18131 1085 18143
rect 1119 18131 1158 18143
rect 1192 18131 1231 18143
rect 195 18079 201 18131
rect 253 18079 269 18131
rect 321 18079 337 18131
rect 389 18079 404 18131
rect 462 18120 471 18131
rect 535 18120 538 18131
rect 791 18120 793 18131
rect 858 18120 866 18131
rect 925 18120 939 18131
rect 456 18079 471 18120
rect 523 18079 538 18120
rect 590 18079 605 18120
rect 657 18079 672 18120
rect 724 18079 739 18120
rect 791 18079 806 18120
rect 858 18079 873 18120
rect 925 18079 940 18120
rect 992 18079 1007 18131
rect 1059 18079 1074 18131
rect 1126 18079 1141 18131
rect 1193 18079 1208 18131
rect 1265 18120 1304 18154
rect 1338 18120 1377 18154
rect 1411 18120 1450 18154
rect 1484 18120 1523 18154
rect 1557 18120 1596 18154
rect 1630 18120 1669 18154
rect 1703 18120 1742 18154
rect 1776 18120 1815 18154
rect 1849 18120 1888 18154
rect 1922 18120 1961 18154
rect 1995 18120 2034 18154
rect 2068 18120 2107 18154
rect 2141 18120 2180 18154
rect 2214 18120 2253 18154
rect 2287 18120 2326 18154
rect 2360 18120 2399 18154
rect 2433 18120 2472 18154
rect 2506 18120 2545 18154
rect 2579 18120 2618 18154
rect 2652 18120 2691 18154
rect 2725 18120 2764 18154
rect 2798 18120 2837 18154
rect 2871 18120 2910 18154
rect 2944 18120 2983 18154
rect 3017 18120 3056 18154
rect 3090 18120 3129 18154
rect 3163 18120 3202 18154
rect 3236 18120 3275 18154
rect 3309 18120 3348 18154
rect 3382 18120 3421 18154
rect 3455 18120 3494 18154
rect 3528 18120 3566 18154
rect 3600 18120 3638 18154
rect 3672 18120 3710 18154
rect 3744 18120 3782 18154
rect 3816 18120 3854 18154
rect 3888 18120 3926 18154
rect 3960 18120 3998 18154
rect 4032 18120 4070 18154
rect 4104 18120 4142 18154
rect 4176 18120 4214 18154
rect 4248 18120 4286 18154
rect 4320 18120 4358 18154
rect 4392 18120 4430 18154
rect 4464 18120 4502 18154
rect 4536 18120 4574 18154
rect 4608 18120 4646 18154
rect 4680 18120 4718 18154
rect 4752 18120 4790 18154
rect 4824 18120 4862 18154
rect 4896 18120 4934 18154
rect 4968 18120 5006 18154
rect 5040 18120 5078 18154
rect 5112 18120 5150 18154
rect 5184 18120 5222 18154
rect 5256 18120 5294 18154
rect 5328 18120 5366 18154
rect 5400 18120 5438 18154
rect 5472 18120 5510 18154
rect 5544 18120 5582 18154
rect 5616 18120 5654 18154
rect 5688 18120 5726 18154
rect 5760 18120 5798 18154
rect 5832 18120 5870 18154
rect 5904 18120 5942 18154
rect 5976 18120 6014 18154
rect 6048 18120 6086 18154
rect 6120 18120 6158 18154
rect 6192 18120 6230 18154
rect 6264 18120 6302 18154
rect 6336 18120 6374 18154
rect 6408 18120 6446 18154
rect 6480 18120 6518 18154
rect 6552 18120 6590 18154
rect 6624 18120 6662 18154
rect 6696 18120 6734 18154
rect 6768 18120 6806 18154
rect 6840 18120 6878 18154
rect 6912 18120 6950 18154
rect 6984 18120 7022 18154
rect 7056 18120 7094 18154
rect 7128 18120 7166 18154
rect 7200 18120 7238 18154
rect 7272 18120 7310 18154
rect 7344 18120 7382 18154
rect 7416 18120 7454 18154
rect 7488 18120 7526 18154
rect 7560 18120 7598 18154
rect 7632 18120 7670 18154
rect 7704 18120 7742 18154
rect 7776 18120 7814 18154
rect 7848 18120 7886 18154
rect 7920 18120 7958 18154
rect 7992 18120 8030 18154
rect 8064 18120 8102 18154
rect 8136 18120 8174 18154
rect 8208 18120 8246 18154
rect 8280 18120 8318 18154
rect 8352 18120 8390 18154
rect 8424 18120 8462 18154
rect 8496 18120 8534 18154
rect 8568 18120 8606 18154
rect 8640 18120 8678 18154
rect 8712 18120 8750 18154
rect 8784 18120 8822 18154
rect 8856 18120 8894 18154
rect 8928 18120 8966 18154
rect 9000 18120 9038 18154
rect 9072 18120 9110 18154
rect 9144 18120 9182 18154
rect 9216 18120 9254 18154
rect 9288 18120 9326 18154
rect 9360 18120 9398 18154
rect 9432 18120 9470 18154
rect 9504 18120 9542 18154
rect 9576 18120 9614 18154
rect 9648 18120 9686 18154
rect 9720 18120 9758 18154
rect 9792 18120 9830 18154
rect 9864 18120 9902 18154
rect 9936 18120 9974 18154
rect 10008 18120 10046 18154
rect 10080 18120 10118 18154
rect 10152 18120 10190 18154
rect 10224 18120 10262 18154
rect 10296 18120 10334 18154
rect 10368 18120 10406 18154
rect 10440 18120 10478 18154
rect 10512 18120 10550 18154
rect 10584 18120 10622 18154
rect 10656 18120 10694 18154
rect 10728 18120 10766 18154
rect 10800 18120 10838 18154
rect 10872 18120 10910 18154
rect 10944 18120 10982 18154
rect 11016 18120 11054 18154
rect 11088 18120 11126 18154
rect 11160 18120 11198 18154
rect 11232 18120 11270 18154
rect 11304 18120 11342 18154
rect 11376 18120 11414 18154
rect 11448 18120 11486 18154
rect 11520 18120 11558 18154
rect 11592 18120 11630 18154
rect 11664 18120 11702 18154
rect 11736 18120 11774 18154
rect 11808 18120 11846 18154
rect 11880 18120 11918 18154
rect 11952 18120 11990 18154
rect 12024 18120 12062 18154
rect 12096 18120 12134 18154
rect 12168 18120 12206 18154
rect 12240 18120 12278 18154
rect 12312 18120 12350 18154
rect 12384 18120 12422 18154
rect 12456 18120 12494 18154
rect 12528 18120 12566 18154
rect 12600 18120 12638 18154
rect 12672 18120 12710 18154
rect 12744 18120 12782 18154
rect 12816 18120 12854 18154
rect 12888 18120 12926 18154
rect 12960 18120 12998 18154
rect 13032 18120 13070 18154
rect 13104 18120 13142 18154
rect 13176 18120 13214 18154
rect 13248 18120 13286 18154
rect 13320 18120 13358 18154
rect 13392 18120 13430 18154
rect 13464 18120 13502 18154
rect 13536 18120 13574 18154
rect 13608 18120 13646 18154
rect 13680 18120 13718 18154
rect 13752 18120 13790 18154
rect 13824 18120 13862 18154
rect 13896 18120 13934 18154
rect 13968 18120 14006 18154
rect 14040 18120 14078 18154
rect 14112 18120 14150 18154
rect 14184 18120 14222 18154
rect 14256 18120 14294 18154
rect 14328 18120 14366 18154
rect 14400 18120 14438 18154
rect 14472 18120 14510 18154
rect 14544 18120 14582 18154
rect 14616 18120 14654 18154
rect 14688 18120 14726 18154
rect 14760 18120 14772 18154
rect 1260 18079 14772 18120
rect 195 18078 14772 18079
rect 195 18067 209 18078
rect 243 18067 282 18078
rect 316 18067 355 18078
rect 389 18067 428 18078
rect 462 18067 501 18078
rect 535 18067 574 18078
rect 608 18067 647 18078
rect 681 18067 720 18078
rect 754 18067 793 18078
rect 827 18067 866 18078
rect 900 18067 939 18078
rect 973 18067 1012 18078
rect 1046 18067 1085 18078
rect 1119 18067 1158 18078
rect 1192 18067 1231 18078
rect 195 18015 201 18067
rect 253 18015 269 18067
rect 321 18015 337 18067
rect 389 18015 404 18067
rect 462 18044 471 18067
rect 535 18044 538 18067
rect 791 18044 793 18067
rect 858 18044 866 18067
rect 925 18044 939 18067
rect 456 18015 471 18044
rect 523 18015 538 18044
rect 590 18015 605 18044
rect 657 18015 672 18044
rect 724 18015 739 18044
rect 791 18015 806 18044
rect 858 18015 873 18044
rect 925 18015 940 18044
rect 992 18015 1007 18067
rect 1059 18015 1074 18067
rect 1126 18015 1141 18067
rect 1193 18015 1208 18067
rect 1265 18044 1304 18078
rect 1338 18044 1377 18078
rect 1411 18044 1450 18078
rect 1484 18044 1523 18078
rect 1557 18044 1596 18078
rect 1630 18044 1669 18078
rect 1703 18044 1742 18078
rect 1776 18044 1815 18078
rect 1849 18044 1888 18078
rect 1922 18044 1961 18078
rect 1995 18044 2034 18078
rect 2068 18044 2107 18078
rect 2141 18044 2180 18078
rect 2214 18044 2253 18078
rect 2287 18044 2326 18078
rect 2360 18044 2399 18078
rect 2433 18044 2472 18078
rect 2506 18044 2545 18078
rect 2579 18044 2618 18078
rect 2652 18044 2691 18078
rect 2725 18044 2764 18078
rect 2798 18044 2837 18078
rect 2871 18044 2910 18078
rect 2944 18044 2983 18078
rect 3017 18044 3056 18078
rect 3090 18044 3129 18078
rect 3163 18044 3202 18078
rect 3236 18044 3275 18078
rect 3309 18044 3348 18078
rect 3382 18044 3421 18078
rect 3455 18044 3494 18078
rect 3528 18044 3566 18078
rect 3600 18044 3638 18078
rect 3672 18044 3710 18078
rect 3744 18044 3782 18078
rect 3816 18044 3854 18078
rect 3888 18044 3926 18078
rect 3960 18044 3998 18078
rect 4032 18044 4070 18078
rect 4104 18044 4142 18078
rect 4176 18044 4214 18078
rect 4248 18044 4286 18078
rect 4320 18044 4358 18078
rect 4392 18044 4430 18078
rect 4464 18044 4502 18078
rect 4536 18044 4574 18078
rect 4608 18044 4646 18078
rect 4680 18044 4718 18078
rect 4752 18044 4790 18078
rect 4824 18044 4862 18078
rect 4896 18044 4934 18078
rect 4968 18044 5006 18078
rect 5040 18044 5078 18078
rect 5112 18044 5150 18078
rect 5184 18044 5222 18078
rect 5256 18044 5294 18078
rect 5328 18044 5366 18078
rect 5400 18044 5438 18078
rect 5472 18044 5510 18078
rect 5544 18044 5582 18078
rect 5616 18044 5654 18078
rect 5688 18044 5726 18078
rect 5760 18044 5798 18078
rect 5832 18044 5870 18078
rect 5904 18044 5942 18078
rect 5976 18044 6014 18078
rect 6048 18044 6086 18078
rect 6120 18044 6158 18078
rect 6192 18044 6230 18078
rect 6264 18044 6302 18078
rect 6336 18044 6374 18078
rect 6408 18044 6446 18078
rect 6480 18044 6518 18078
rect 6552 18044 6590 18078
rect 6624 18044 6662 18078
rect 6696 18044 6734 18078
rect 6768 18044 6806 18078
rect 6840 18044 6878 18078
rect 6912 18044 6950 18078
rect 6984 18044 7022 18078
rect 7056 18044 7094 18078
rect 7128 18044 7166 18078
rect 7200 18044 7238 18078
rect 7272 18044 7310 18078
rect 7344 18044 7382 18078
rect 7416 18044 7454 18078
rect 7488 18044 7526 18078
rect 7560 18044 7598 18078
rect 7632 18044 7670 18078
rect 7704 18044 7742 18078
rect 7776 18044 7814 18078
rect 7848 18044 7886 18078
rect 7920 18044 7958 18078
rect 7992 18044 8030 18078
rect 8064 18044 8102 18078
rect 8136 18044 8174 18078
rect 8208 18044 8246 18078
rect 8280 18044 8318 18078
rect 8352 18044 8390 18078
rect 8424 18044 8462 18078
rect 8496 18044 8534 18078
rect 8568 18044 8606 18078
rect 8640 18044 8678 18078
rect 8712 18044 8750 18078
rect 8784 18044 8822 18078
rect 8856 18044 8894 18078
rect 8928 18044 8966 18078
rect 9000 18044 9038 18078
rect 9072 18044 9110 18078
rect 9144 18044 9182 18078
rect 9216 18044 9254 18078
rect 9288 18044 9326 18078
rect 9360 18044 9398 18078
rect 9432 18044 9470 18078
rect 9504 18044 9542 18078
rect 9576 18044 9614 18078
rect 9648 18044 9686 18078
rect 9720 18044 9758 18078
rect 9792 18044 9830 18078
rect 9864 18044 9902 18078
rect 9936 18044 9974 18078
rect 10008 18044 10046 18078
rect 10080 18044 10118 18078
rect 10152 18044 10190 18078
rect 10224 18044 10262 18078
rect 10296 18044 10334 18078
rect 10368 18044 10406 18078
rect 10440 18044 10478 18078
rect 10512 18044 10550 18078
rect 10584 18044 10622 18078
rect 10656 18044 10694 18078
rect 10728 18044 10766 18078
rect 10800 18044 10838 18078
rect 10872 18044 10910 18078
rect 10944 18044 10982 18078
rect 11016 18044 11054 18078
rect 11088 18044 11126 18078
rect 11160 18044 11198 18078
rect 11232 18044 11270 18078
rect 11304 18044 11342 18078
rect 11376 18044 11414 18078
rect 11448 18044 11486 18078
rect 11520 18044 11558 18078
rect 11592 18044 11630 18078
rect 11664 18044 11702 18078
rect 11736 18044 11774 18078
rect 11808 18044 11846 18078
rect 11880 18044 11918 18078
rect 11952 18044 11990 18078
rect 12024 18044 12062 18078
rect 12096 18044 12134 18078
rect 12168 18044 12206 18078
rect 12240 18044 12278 18078
rect 12312 18044 12350 18078
rect 12384 18044 12422 18078
rect 12456 18044 12494 18078
rect 12528 18044 12566 18078
rect 12600 18044 12638 18078
rect 12672 18044 12710 18078
rect 12744 18044 12782 18078
rect 12816 18044 12854 18078
rect 12888 18044 12926 18078
rect 12960 18044 12998 18078
rect 13032 18044 13070 18078
rect 13104 18044 13142 18078
rect 13176 18044 13214 18078
rect 13248 18044 13286 18078
rect 13320 18044 13358 18078
rect 13392 18044 13430 18078
rect 13464 18044 13502 18078
rect 13536 18044 13574 18078
rect 13608 18044 13646 18078
rect 13680 18044 13718 18078
rect 13752 18044 13790 18078
rect 13824 18044 13862 18078
rect 13896 18044 13934 18078
rect 13968 18044 14006 18078
rect 14040 18044 14078 18078
rect 14112 18044 14150 18078
rect 14184 18044 14222 18078
rect 14256 18044 14294 18078
rect 14328 18044 14366 18078
rect 14400 18044 14438 18078
rect 14472 18044 14510 18078
rect 14544 18044 14582 18078
rect 14616 18044 14654 18078
rect 14688 18044 14726 18078
rect 14760 18044 14772 18078
rect 1260 18015 14772 18044
rect 195 18003 14772 18015
rect 195 17951 201 18003
rect 253 17951 269 18003
rect 321 17951 337 18003
rect 389 17951 404 18003
rect 456 18002 471 18003
rect 523 18002 538 18003
rect 590 18002 605 18003
rect 657 18002 672 18003
rect 724 18002 739 18003
rect 791 18002 806 18003
rect 858 18002 873 18003
rect 925 18002 940 18003
rect 462 17968 471 18002
rect 535 17968 538 18002
rect 791 17968 793 18002
rect 858 17968 866 18002
rect 925 17968 939 18002
rect 456 17951 471 17968
rect 523 17951 538 17968
rect 590 17951 605 17968
rect 657 17951 672 17968
rect 724 17951 739 17968
rect 791 17951 806 17968
rect 858 17951 873 17968
rect 925 17951 940 17968
rect 992 17951 1007 18003
rect 1059 17951 1074 18003
rect 1126 17951 1141 18003
rect 1193 17951 1208 18003
rect 1260 18002 14772 18003
rect 1265 17968 1304 18002
rect 1338 17968 1377 18002
rect 1411 17968 1450 18002
rect 1484 17968 1523 18002
rect 1557 17968 1596 18002
rect 1630 17968 1669 18002
rect 1703 17968 1742 18002
rect 1776 17968 1815 18002
rect 1849 17968 1888 18002
rect 1922 17968 1961 18002
rect 1995 17968 2034 18002
rect 2068 17968 2107 18002
rect 2141 17968 2180 18002
rect 2214 17968 2253 18002
rect 2287 17968 2326 18002
rect 2360 17968 2399 18002
rect 2433 17968 2472 18002
rect 2506 17968 2545 18002
rect 2579 17968 2618 18002
rect 2652 17968 2691 18002
rect 2725 17968 2764 18002
rect 2798 17968 2837 18002
rect 2871 17968 2910 18002
rect 2944 17968 2983 18002
rect 3017 17968 3056 18002
rect 3090 17968 3129 18002
rect 3163 17968 3202 18002
rect 3236 17968 3275 18002
rect 3309 17968 3348 18002
rect 3382 17968 3421 18002
rect 3455 17968 3494 18002
rect 3528 17968 3566 18002
rect 3600 17968 3638 18002
rect 3672 17968 3710 18002
rect 3744 17968 3782 18002
rect 3816 17968 3854 18002
rect 3888 17968 3926 18002
rect 3960 17968 3998 18002
rect 4032 17968 4070 18002
rect 4104 17968 4142 18002
rect 4176 17968 4214 18002
rect 4248 17968 4286 18002
rect 4320 17968 4358 18002
rect 4392 17968 4430 18002
rect 4464 17968 4502 18002
rect 4536 17968 4574 18002
rect 4608 17968 4646 18002
rect 4680 17968 4718 18002
rect 4752 17968 4790 18002
rect 4824 17968 4862 18002
rect 4896 17968 4934 18002
rect 4968 17968 5006 18002
rect 5040 17968 5078 18002
rect 5112 17968 5150 18002
rect 5184 17968 5222 18002
rect 5256 17968 5294 18002
rect 5328 17968 5366 18002
rect 5400 17968 5438 18002
rect 5472 17968 5510 18002
rect 5544 17968 5582 18002
rect 5616 17968 5654 18002
rect 5688 17968 5726 18002
rect 5760 17968 5798 18002
rect 5832 17968 5870 18002
rect 5904 17968 5942 18002
rect 5976 17968 6014 18002
rect 6048 17968 6086 18002
rect 6120 17968 6158 18002
rect 6192 17968 6230 18002
rect 6264 17968 6302 18002
rect 6336 17968 6374 18002
rect 6408 17968 6446 18002
rect 6480 17968 6518 18002
rect 6552 17968 6590 18002
rect 6624 17968 6662 18002
rect 6696 17968 6734 18002
rect 6768 17968 6806 18002
rect 6840 17968 6878 18002
rect 6912 17968 6950 18002
rect 6984 17968 7022 18002
rect 7056 17968 7094 18002
rect 7128 17968 7166 18002
rect 7200 17968 7238 18002
rect 7272 17968 7310 18002
rect 7344 17968 7382 18002
rect 7416 17968 7454 18002
rect 7488 17968 7526 18002
rect 7560 17968 7598 18002
rect 7632 17968 7670 18002
rect 7704 17968 7742 18002
rect 7776 17968 7814 18002
rect 7848 17968 7886 18002
rect 7920 17968 7958 18002
rect 7992 17968 8030 18002
rect 8064 17968 8102 18002
rect 8136 17968 8174 18002
rect 8208 17968 8246 18002
rect 8280 17968 8318 18002
rect 8352 17968 8390 18002
rect 8424 17968 8462 18002
rect 8496 17968 8534 18002
rect 8568 17968 8606 18002
rect 8640 17968 8678 18002
rect 8712 17968 8750 18002
rect 8784 17968 8822 18002
rect 8856 17968 8894 18002
rect 8928 17968 8966 18002
rect 9000 17968 9038 18002
rect 9072 17968 9110 18002
rect 9144 17968 9182 18002
rect 9216 17968 9254 18002
rect 9288 17968 9326 18002
rect 9360 17968 9398 18002
rect 9432 17968 9470 18002
rect 9504 17968 9542 18002
rect 9576 17968 9614 18002
rect 9648 17968 9686 18002
rect 9720 17968 9758 18002
rect 9792 17968 9830 18002
rect 9864 17968 9902 18002
rect 9936 17968 9974 18002
rect 10008 17968 10046 18002
rect 10080 17968 10118 18002
rect 10152 17968 10190 18002
rect 10224 17968 10262 18002
rect 10296 17968 10334 18002
rect 10368 17968 10406 18002
rect 10440 17968 10478 18002
rect 10512 17968 10550 18002
rect 10584 17968 10622 18002
rect 10656 17968 10694 18002
rect 10728 17968 10766 18002
rect 10800 17968 10838 18002
rect 10872 17968 10910 18002
rect 10944 17968 10982 18002
rect 11016 17968 11054 18002
rect 11088 17968 11126 18002
rect 11160 17968 11198 18002
rect 11232 17968 11270 18002
rect 11304 17968 11342 18002
rect 11376 17968 11414 18002
rect 11448 17968 11486 18002
rect 11520 17968 11558 18002
rect 11592 17968 11630 18002
rect 11664 17968 11702 18002
rect 11736 17968 11774 18002
rect 11808 17968 11846 18002
rect 11880 17968 11918 18002
rect 11952 17968 11990 18002
rect 12024 17968 12062 18002
rect 12096 17968 12134 18002
rect 12168 17968 12206 18002
rect 12240 17968 12278 18002
rect 12312 17968 12350 18002
rect 12384 17968 12422 18002
rect 12456 17968 12494 18002
rect 12528 17968 12566 18002
rect 12600 17968 12638 18002
rect 12672 17968 12710 18002
rect 12744 17968 12782 18002
rect 12816 17968 12854 18002
rect 12888 17968 12926 18002
rect 12960 17968 12998 18002
rect 13032 17968 13070 18002
rect 13104 17968 13142 18002
rect 13176 17968 13214 18002
rect 13248 17968 13286 18002
rect 13320 17968 13358 18002
rect 13392 17968 13430 18002
rect 13464 17968 13502 18002
rect 13536 17968 13574 18002
rect 13608 17968 13646 18002
rect 13680 17968 13718 18002
rect 13752 17968 13790 18002
rect 13824 17968 13862 18002
rect 13896 17968 13934 18002
rect 13968 17968 14006 18002
rect 14040 17968 14078 18002
rect 14112 17968 14150 18002
rect 14184 17968 14222 18002
rect 14256 17968 14294 18002
rect 14328 17968 14366 18002
rect 14400 17968 14438 18002
rect 14472 17968 14510 18002
rect 14544 17968 14582 18002
rect 14616 17968 14654 18002
rect 14688 17968 14726 18002
rect 14760 17968 14772 18002
rect 1260 17951 14772 17968
rect 195 17939 14772 17951
rect 195 17887 201 17939
rect 253 17887 269 17939
rect 321 17887 337 17939
rect 389 17887 404 17939
rect 456 17926 471 17939
rect 523 17926 538 17939
rect 590 17926 605 17939
rect 657 17926 672 17939
rect 724 17926 739 17939
rect 791 17926 806 17939
rect 858 17926 873 17939
rect 925 17926 940 17939
rect 462 17892 471 17926
rect 535 17892 538 17926
rect 791 17892 793 17926
rect 858 17892 866 17926
rect 925 17892 939 17926
rect 456 17887 471 17892
rect 523 17887 538 17892
rect 590 17887 605 17892
rect 657 17887 672 17892
rect 724 17887 739 17892
rect 791 17887 806 17892
rect 858 17887 873 17892
rect 925 17887 940 17892
rect 992 17887 1007 17939
rect 1059 17887 1074 17939
rect 1126 17887 1141 17939
rect 1193 17887 1208 17939
rect 1260 17926 14772 17939
rect 1265 17892 1304 17926
rect 1338 17892 1377 17926
rect 1411 17892 1450 17926
rect 1484 17892 1523 17926
rect 1557 17892 1596 17926
rect 1630 17892 1669 17926
rect 1703 17892 1742 17926
rect 1776 17892 1815 17926
rect 1849 17892 1888 17926
rect 1922 17892 1961 17926
rect 1995 17892 2034 17926
rect 2068 17892 2107 17926
rect 2141 17892 2180 17926
rect 2214 17892 2253 17926
rect 2287 17892 2326 17926
rect 2360 17892 2399 17926
rect 2433 17892 2472 17926
rect 2506 17892 2545 17926
rect 2579 17892 2618 17926
rect 2652 17892 2691 17926
rect 2725 17892 2764 17926
rect 2798 17892 2837 17926
rect 2871 17892 2910 17926
rect 2944 17892 2983 17926
rect 3017 17892 3056 17926
rect 3090 17892 3129 17926
rect 3163 17892 3202 17926
rect 3236 17892 3275 17926
rect 3309 17892 3348 17926
rect 3382 17892 3421 17926
rect 3455 17892 3494 17926
rect 3528 17892 3566 17926
rect 3600 17892 3638 17926
rect 3672 17892 3710 17926
rect 3744 17892 3782 17926
rect 3816 17892 3854 17926
rect 3888 17892 3926 17926
rect 3960 17892 3998 17926
rect 4032 17892 4070 17926
rect 4104 17892 4142 17926
rect 4176 17892 4214 17926
rect 4248 17892 4286 17926
rect 4320 17892 4358 17926
rect 4392 17892 4430 17926
rect 4464 17892 4502 17926
rect 4536 17892 4574 17926
rect 4608 17892 4646 17926
rect 4680 17892 4718 17926
rect 4752 17892 4790 17926
rect 4824 17892 4862 17926
rect 4896 17892 4934 17926
rect 4968 17892 5006 17926
rect 5040 17892 5078 17926
rect 5112 17892 5150 17926
rect 5184 17892 5222 17926
rect 5256 17892 5294 17926
rect 5328 17892 5366 17926
rect 5400 17892 5438 17926
rect 5472 17892 5510 17926
rect 5544 17892 5582 17926
rect 5616 17892 5654 17926
rect 5688 17892 5726 17926
rect 5760 17892 5798 17926
rect 5832 17892 5870 17926
rect 5904 17892 5942 17926
rect 5976 17892 6014 17926
rect 6048 17892 6086 17926
rect 6120 17892 6158 17926
rect 6192 17892 6230 17926
rect 6264 17892 6302 17926
rect 6336 17892 6374 17926
rect 6408 17892 6446 17926
rect 6480 17892 6518 17926
rect 6552 17892 6590 17926
rect 6624 17892 6662 17926
rect 6696 17892 6734 17926
rect 6768 17892 6806 17926
rect 6840 17892 6878 17926
rect 6912 17892 6950 17926
rect 6984 17892 7022 17926
rect 7056 17892 7094 17926
rect 7128 17892 7166 17926
rect 7200 17892 7238 17926
rect 7272 17892 7310 17926
rect 7344 17892 7382 17926
rect 7416 17892 7454 17926
rect 7488 17892 7526 17926
rect 7560 17892 7598 17926
rect 7632 17892 7670 17926
rect 7704 17892 7742 17926
rect 7776 17892 7814 17926
rect 7848 17892 7886 17926
rect 7920 17892 7958 17926
rect 7992 17892 8030 17926
rect 8064 17892 8102 17926
rect 8136 17892 8174 17926
rect 8208 17892 8246 17926
rect 8280 17892 8318 17926
rect 8352 17892 8390 17926
rect 8424 17892 8462 17926
rect 8496 17892 8534 17926
rect 8568 17892 8606 17926
rect 8640 17892 8678 17926
rect 8712 17892 8750 17926
rect 8784 17892 8822 17926
rect 8856 17892 8894 17926
rect 8928 17892 8966 17926
rect 9000 17892 9038 17926
rect 9072 17892 9110 17926
rect 9144 17892 9182 17926
rect 9216 17892 9254 17926
rect 9288 17892 9326 17926
rect 9360 17892 9398 17926
rect 9432 17892 9470 17926
rect 9504 17892 9542 17926
rect 9576 17892 9614 17926
rect 9648 17892 9686 17926
rect 9720 17892 9758 17926
rect 9792 17892 9830 17926
rect 9864 17892 9902 17926
rect 9936 17892 9974 17926
rect 10008 17892 10046 17926
rect 10080 17892 10118 17926
rect 10152 17892 10190 17926
rect 10224 17892 10262 17926
rect 10296 17892 10334 17926
rect 10368 17892 10406 17926
rect 10440 17892 10478 17926
rect 10512 17892 10550 17926
rect 10584 17892 10622 17926
rect 10656 17892 10694 17926
rect 10728 17892 10766 17926
rect 10800 17892 10838 17926
rect 10872 17892 10910 17926
rect 10944 17892 10982 17926
rect 11016 17892 11054 17926
rect 11088 17892 11126 17926
rect 11160 17892 11198 17926
rect 11232 17892 11270 17926
rect 11304 17892 11342 17926
rect 11376 17892 11414 17926
rect 11448 17892 11486 17926
rect 11520 17892 11558 17926
rect 11592 17892 11630 17926
rect 11664 17892 11702 17926
rect 11736 17892 11774 17926
rect 11808 17892 11846 17926
rect 11880 17892 11918 17926
rect 11952 17892 11990 17926
rect 12024 17892 12062 17926
rect 12096 17892 12134 17926
rect 12168 17892 12206 17926
rect 12240 17892 12278 17926
rect 12312 17892 12350 17926
rect 12384 17892 12422 17926
rect 12456 17892 12494 17926
rect 12528 17892 12566 17926
rect 12600 17892 12638 17926
rect 12672 17892 12710 17926
rect 12744 17892 12782 17926
rect 12816 17892 12854 17926
rect 12888 17892 12926 17926
rect 12960 17892 12998 17926
rect 13032 17892 13070 17926
rect 13104 17892 13142 17926
rect 13176 17892 13214 17926
rect 13248 17892 13286 17926
rect 13320 17892 13358 17926
rect 13392 17892 13430 17926
rect 13464 17892 13502 17926
rect 13536 17892 13574 17926
rect 13608 17892 13646 17926
rect 13680 17892 13718 17926
rect 13752 17892 13790 17926
rect 13824 17892 13862 17926
rect 13896 17892 13934 17926
rect 13968 17892 14006 17926
rect 14040 17892 14078 17926
rect 14112 17892 14150 17926
rect 14184 17892 14222 17926
rect 14256 17892 14294 17926
rect 14328 17892 14366 17926
rect 14400 17892 14438 17926
rect 14472 17892 14510 17926
rect 14544 17892 14582 17926
rect 14616 17892 14654 17926
rect 14688 17892 14726 17926
rect 14760 17892 14772 17926
rect 1260 17887 14772 17892
rect 195 17881 14772 17887
<< via1 >>
rect 14285 35712 14337 35764
rect 14349 35712 14401 35764
rect 14285 35632 14337 35684
rect 14349 35632 14401 35684
rect 14285 35552 14337 35604
rect 14349 35552 14401 35604
rect 581 28580 633 28632
rect 650 28580 702 28632
rect 719 28580 771 28632
rect 788 28580 840 28632
rect 857 28580 909 28632
rect 926 28580 978 28632
rect 995 28580 1047 28632
rect 1063 28580 1115 28632
rect 1131 28580 1183 28632
rect 581 28506 633 28558
rect 650 28506 702 28558
rect 719 28506 771 28558
rect 788 28506 840 28558
rect 857 28506 909 28558
rect 926 28506 978 28558
rect 995 28506 1047 28558
rect 1063 28506 1115 28558
rect 1131 28506 1183 28558
rect 581 28432 633 28484
rect 650 28432 702 28484
rect 719 28432 771 28484
rect 788 28432 840 28484
rect 857 28432 909 28484
rect 926 28432 978 28484
rect 995 28432 1047 28484
rect 1063 28432 1115 28484
rect 1131 28432 1183 28484
rect 3478 28581 3530 28633
rect 3546 28581 3598 28633
rect 3614 28581 3666 28633
rect 3682 28581 3734 28633
rect 3750 28581 3802 28633
rect 3818 28581 3870 28633
rect 3886 28581 3938 28633
rect 3954 28581 4006 28633
rect 4021 28581 4073 28633
rect 4088 28581 4140 28633
rect 4155 28581 4207 28633
rect 4222 28581 4274 28633
rect 4289 28581 4341 28633
rect 4356 28581 4408 28633
rect 4423 28581 4475 28633
rect 4490 28581 4542 28633
rect 4557 28581 4609 28633
rect 3478 28507 3530 28559
rect 3546 28507 3598 28559
rect 3614 28507 3666 28559
rect 3682 28507 3734 28559
rect 3750 28507 3802 28559
rect 3818 28507 3870 28559
rect 3886 28507 3938 28559
rect 3954 28507 4006 28559
rect 4021 28507 4073 28559
rect 4088 28507 4140 28559
rect 4155 28507 4207 28559
rect 4222 28507 4274 28559
rect 4289 28507 4341 28559
rect 4356 28507 4408 28559
rect 4423 28507 4475 28559
rect 4490 28507 4542 28559
rect 4557 28507 4609 28559
rect 3478 28433 3530 28485
rect 3546 28433 3598 28485
rect 3614 28433 3666 28485
rect 3682 28433 3734 28485
rect 3750 28433 3802 28485
rect 3818 28433 3870 28485
rect 3886 28433 3938 28485
rect 3954 28433 4006 28485
rect 4021 28433 4073 28485
rect 4088 28433 4140 28485
rect 4155 28433 4207 28485
rect 4222 28433 4274 28485
rect 4289 28433 4341 28485
rect 4356 28433 4408 28485
rect 4423 28433 4475 28485
rect 4490 28433 4542 28485
rect 4557 28433 4609 28485
rect 5461 28581 5513 28633
rect 5528 28581 5580 28633
rect 5595 28581 5647 28633
rect 5662 28581 5714 28633
rect 5729 28581 5781 28633
rect 5796 28581 5848 28633
rect 5863 28581 5915 28633
rect 5930 28581 5982 28633
rect 5997 28581 6049 28633
rect 6064 28581 6116 28633
rect 6132 28581 6184 28633
rect 6200 28581 6252 28633
rect 6268 28581 6320 28633
rect 6336 28581 6388 28633
rect 6404 28581 6456 28633
rect 6472 28581 6524 28633
rect 6540 28581 6592 28633
rect 5461 28507 5513 28559
rect 5528 28507 5580 28559
rect 5595 28507 5647 28559
rect 5662 28507 5714 28559
rect 5729 28507 5781 28559
rect 5796 28507 5848 28559
rect 5863 28507 5915 28559
rect 5930 28507 5982 28559
rect 5997 28507 6049 28559
rect 6064 28507 6116 28559
rect 6132 28507 6184 28559
rect 6200 28507 6252 28559
rect 6268 28507 6320 28559
rect 6336 28507 6388 28559
rect 6404 28507 6456 28559
rect 6472 28507 6524 28559
rect 6540 28507 6592 28559
rect 5461 28433 5513 28485
rect 5528 28433 5580 28485
rect 5595 28433 5647 28485
rect 5662 28433 5714 28485
rect 5729 28433 5781 28485
rect 5796 28433 5848 28485
rect 5863 28433 5915 28485
rect 5930 28433 5982 28485
rect 5997 28433 6049 28485
rect 6064 28433 6116 28485
rect 6132 28433 6184 28485
rect 6200 28433 6252 28485
rect 6268 28433 6320 28485
rect 6336 28433 6388 28485
rect 6404 28433 6456 28485
rect 6472 28433 6524 28485
rect 6540 28433 6592 28485
rect 7445 28581 7497 28633
rect 7512 28581 7564 28633
rect 7579 28581 7631 28633
rect 7646 28581 7698 28633
rect 7713 28581 7765 28633
rect 7780 28581 7832 28633
rect 7847 28581 7899 28633
rect 7914 28581 7966 28633
rect 7981 28581 8033 28633
rect 8048 28581 8100 28633
rect 8116 28581 8168 28633
rect 8184 28581 8236 28633
rect 8252 28581 8304 28633
rect 8320 28581 8372 28633
rect 8388 28581 8440 28633
rect 8456 28581 8508 28633
rect 8524 28581 8576 28633
rect 7445 28507 7497 28559
rect 7512 28507 7564 28559
rect 7579 28507 7631 28559
rect 7646 28507 7698 28559
rect 7713 28507 7765 28559
rect 7780 28507 7832 28559
rect 7847 28507 7899 28559
rect 7914 28507 7966 28559
rect 7981 28507 8033 28559
rect 8048 28507 8100 28559
rect 8116 28507 8168 28559
rect 8184 28507 8236 28559
rect 8252 28507 8304 28559
rect 8320 28507 8372 28559
rect 8388 28507 8440 28559
rect 8456 28507 8508 28559
rect 8524 28507 8576 28559
rect 7445 28433 7497 28485
rect 7512 28433 7564 28485
rect 7579 28433 7631 28485
rect 7646 28433 7698 28485
rect 7713 28433 7765 28485
rect 7780 28433 7832 28485
rect 7847 28433 7899 28485
rect 7914 28433 7966 28485
rect 7981 28433 8033 28485
rect 8048 28433 8100 28485
rect 8116 28433 8168 28485
rect 8184 28433 8236 28485
rect 8252 28433 8304 28485
rect 8320 28433 8372 28485
rect 8388 28433 8440 28485
rect 8456 28433 8508 28485
rect 8524 28433 8576 28485
rect 9429 28581 9481 28633
rect 9517 28581 9569 28633
rect 9429 28507 9481 28559
rect 9517 28507 9569 28559
rect 9429 28433 9481 28485
rect 9517 28433 9569 28485
rect 14282 28575 14334 28627
rect 14358 28575 14410 28627
rect 14434 28575 14486 28627
rect 14510 28575 14562 28627
rect 14586 28575 14638 28627
rect 14282 28510 14334 28562
rect 14358 28510 14410 28562
rect 14434 28510 14486 28562
rect 14510 28510 14562 28562
rect 14586 28510 14638 28562
rect 14282 28445 14334 28497
rect 14358 28445 14410 28497
rect 14434 28445 14486 28497
rect 14510 28445 14562 28497
rect 14586 28445 14638 28497
rect 14282 28380 14334 28432
rect 14358 28380 14410 28432
rect 14434 28380 14486 28432
rect 14510 28380 14562 28432
rect 14586 28380 14638 28432
rect 14282 28315 14334 28367
rect 14358 28315 14410 28367
rect 14434 28315 14486 28367
rect 14510 28315 14562 28367
rect 14586 28315 14638 28367
rect 14282 28250 14334 28302
rect 14358 28250 14410 28302
rect 14434 28250 14486 28302
rect 14510 28250 14562 28302
rect 14586 28250 14638 28302
rect 14282 28185 14334 28237
rect 14358 28185 14410 28237
rect 14434 28185 14486 28237
rect 14510 28185 14562 28237
rect 14586 28185 14638 28237
rect 1303 28122 1355 28124
rect 1371 28122 1423 28124
rect 1439 28122 1491 28124
rect 1507 28122 1559 28124
rect 1575 28122 1627 28124
rect 1303 28088 1314 28122
rect 1314 28088 1353 28122
rect 1353 28088 1355 28122
rect 1371 28088 1387 28122
rect 1387 28088 1423 28122
rect 1439 28088 1460 28122
rect 1460 28088 1491 28122
rect 1507 28088 1533 28122
rect 1533 28088 1559 28122
rect 1575 28088 1605 28122
rect 1605 28088 1627 28122
rect 1303 28072 1355 28088
rect 1371 28072 1423 28088
rect 1439 28072 1491 28088
rect 1507 28072 1559 28088
rect 1575 28072 1627 28088
rect 1643 28122 1695 28124
rect 1643 28088 1677 28122
rect 1677 28088 1695 28122
rect 1643 28072 1695 28088
rect 1711 28122 1763 28124
rect 1711 28088 1715 28122
rect 1715 28088 1749 28122
rect 1749 28088 1763 28122
rect 1711 28072 1763 28088
rect 1779 28122 1831 28124
rect 1779 28088 1787 28122
rect 1787 28088 1821 28122
rect 1821 28088 1831 28122
rect 1779 28072 1831 28088
rect 1847 28122 1899 28124
rect 1847 28088 1859 28122
rect 1859 28088 1893 28122
rect 1893 28088 1899 28122
rect 1847 28072 1899 28088
rect 1914 28122 1966 28124
rect 1914 28088 1931 28122
rect 1931 28088 1965 28122
rect 1965 28088 1966 28122
rect 1914 28072 1966 28088
rect 1981 28122 2033 28124
rect 12157 28122 12209 28124
rect 1981 28088 2003 28122
rect 2003 28088 2033 28122
rect 12157 28088 12189 28122
rect 12189 28088 12209 28122
rect 1981 28072 2033 28088
rect 12157 28072 12209 28088
rect 12225 28122 12277 28124
rect 12225 28088 12227 28122
rect 12227 28088 12261 28122
rect 12261 28088 12277 28122
rect 12225 28072 12277 28088
rect 12293 28122 12345 28124
rect 12293 28088 12299 28122
rect 12299 28088 12333 28122
rect 12333 28088 12345 28122
rect 12293 28072 12345 28088
rect 12361 28122 12413 28124
rect 12361 28088 12371 28122
rect 12371 28088 12405 28122
rect 12405 28088 12413 28122
rect 12361 28072 12413 28088
rect 12429 28122 12481 28124
rect 12429 28088 12443 28122
rect 12443 28088 12477 28122
rect 12477 28088 12481 28122
rect 12429 28072 12481 28088
rect 12497 28122 12549 28124
rect 12497 28088 12515 28122
rect 12515 28088 12549 28122
rect 12497 28072 12549 28088
rect 12565 28122 12617 28124
rect 12633 28122 12685 28124
rect 12701 28122 12753 28124
rect 12768 28122 12820 28124
rect 12835 28122 12887 28124
rect 12565 28088 12587 28122
rect 12587 28088 12617 28122
rect 12633 28088 12659 28122
rect 12659 28088 12685 28122
rect 12701 28088 12731 28122
rect 12731 28088 12753 28122
rect 12768 28088 12803 28122
rect 12803 28088 12820 28122
rect 12835 28088 12837 28122
rect 12837 28088 12875 28122
rect 12875 28088 12887 28122
rect 12565 28072 12617 28088
rect 12633 28072 12685 28088
rect 12701 28072 12753 28088
rect 12768 28072 12820 28088
rect 12835 28072 12887 28088
rect 1303 28040 1355 28058
rect 1371 28040 1423 28058
rect 1439 28040 1491 28058
rect 1507 28040 1559 28058
rect 1575 28040 1627 28058
rect 1303 28006 1314 28040
rect 1314 28006 1353 28040
rect 1353 28006 1355 28040
rect 1371 28006 1387 28040
rect 1387 28006 1423 28040
rect 1439 28006 1460 28040
rect 1460 28006 1491 28040
rect 1507 28006 1533 28040
rect 1533 28006 1559 28040
rect 1575 28006 1605 28040
rect 1605 28006 1627 28040
rect 1643 28040 1695 28058
rect 1643 28006 1677 28040
rect 1677 28006 1695 28040
rect 1711 28040 1763 28058
rect 1711 28006 1715 28040
rect 1715 28006 1749 28040
rect 1749 28006 1763 28040
rect 1779 28040 1831 28058
rect 1779 28006 1787 28040
rect 1787 28006 1821 28040
rect 1821 28006 1831 28040
rect 1847 28040 1899 28058
rect 1847 28006 1859 28040
rect 1859 28006 1893 28040
rect 1893 28006 1899 28040
rect 1914 28040 1966 28058
rect 1914 28006 1931 28040
rect 1931 28006 1965 28040
rect 1965 28006 1966 28040
rect 1981 28040 2033 28058
rect 12157 28040 12209 28058
rect 1981 28006 2003 28040
rect 2003 28006 2033 28040
rect 12157 28006 12189 28040
rect 12189 28006 12209 28040
rect 12225 28040 12277 28058
rect 12225 28006 12227 28040
rect 12227 28006 12261 28040
rect 12261 28006 12277 28040
rect 12293 28040 12345 28058
rect 12293 28006 12299 28040
rect 12299 28006 12333 28040
rect 12333 28006 12345 28040
rect 12361 28040 12413 28058
rect 12361 28006 12371 28040
rect 12371 28006 12405 28040
rect 12405 28006 12413 28040
rect 12429 28040 12481 28058
rect 12429 28006 12443 28040
rect 12443 28006 12477 28040
rect 12477 28006 12481 28040
rect 12497 28040 12549 28058
rect 12497 28006 12515 28040
rect 12515 28006 12549 28040
rect 12565 28040 12617 28058
rect 12633 28040 12685 28058
rect 12701 28040 12753 28058
rect 12768 28040 12820 28058
rect 12835 28040 12887 28058
rect 12565 28006 12587 28040
rect 12587 28006 12617 28040
rect 12633 28006 12659 28040
rect 12659 28006 12685 28040
rect 12701 28006 12731 28040
rect 12731 28006 12753 28040
rect 12768 28006 12803 28040
rect 12803 28006 12820 28040
rect 12835 28006 12837 28040
rect 12837 28006 12875 28040
rect 12875 28006 12887 28040
rect 1303 27958 1355 27992
rect 1371 27958 1423 27992
rect 1439 27958 1491 27992
rect 1507 27958 1559 27992
rect 1575 27958 1627 27992
rect 1303 27940 1314 27958
rect 1314 27940 1353 27958
rect 1353 27940 1355 27958
rect 1371 27940 1387 27958
rect 1387 27940 1423 27958
rect 1439 27940 1460 27958
rect 1460 27940 1491 27958
rect 1507 27940 1533 27958
rect 1533 27940 1559 27958
rect 1575 27940 1605 27958
rect 1605 27940 1627 27958
rect 1643 27958 1695 27992
rect 1643 27940 1677 27958
rect 1677 27940 1695 27958
rect 1711 27958 1763 27992
rect 1711 27940 1715 27958
rect 1715 27940 1749 27958
rect 1749 27940 1763 27958
rect 1779 27958 1831 27992
rect 1779 27940 1787 27958
rect 1787 27940 1821 27958
rect 1821 27940 1831 27958
rect 1847 27958 1899 27992
rect 1847 27940 1859 27958
rect 1859 27940 1893 27958
rect 1893 27940 1899 27958
rect 1914 27958 1966 27992
rect 1914 27940 1931 27958
rect 1931 27940 1965 27958
rect 1965 27940 1966 27958
rect 1981 27958 2033 27992
rect 12157 27958 12209 27992
rect 1981 27940 2003 27958
rect 2003 27940 2033 27958
rect 1303 27924 1314 27926
rect 1314 27924 1353 27926
rect 1353 27924 1355 27926
rect 1371 27924 1387 27926
rect 1387 27924 1423 27926
rect 1439 27924 1460 27926
rect 1460 27924 1491 27926
rect 1507 27924 1533 27926
rect 1533 27924 1559 27926
rect 1575 27924 1605 27926
rect 1605 27924 1627 27926
rect 1303 27876 1355 27924
rect 1371 27876 1423 27924
rect 1439 27876 1491 27924
rect 1507 27876 1559 27924
rect 1575 27876 1627 27924
rect 1303 27874 1314 27876
rect 1314 27874 1353 27876
rect 1353 27874 1355 27876
rect 1371 27874 1387 27876
rect 1387 27874 1423 27876
rect 1439 27874 1460 27876
rect 1460 27874 1491 27876
rect 1507 27874 1533 27876
rect 1533 27874 1559 27876
rect 1575 27874 1605 27876
rect 1605 27874 1627 27876
rect 1643 27924 1677 27926
rect 1677 27924 1695 27926
rect 1643 27876 1695 27924
rect 1643 27874 1677 27876
rect 1677 27874 1695 27876
rect 1711 27924 1715 27926
rect 1715 27924 1749 27926
rect 1749 27924 1763 27926
rect 1711 27876 1763 27924
rect 1711 27874 1715 27876
rect 1715 27874 1749 27876
rect 1749 27874 1763 27876
rect 1779 27924 1787 27926
rect 1787 27924 1821 27926
rect 1821 27924 1831 27926
rect 1779 27876 1831 27924
rect 1779 27874 1787 27876
rect 1787 27874 1821 27876
rect 1821 27874 1831 27876
rect 1847 27924 1859 27926
rect 1859 27924 1893 27926
rect 1893 27924 1899 27926
rect 1847 27876 1899 27924
rect 1847 27874 1859 27876
rect 1859 27874 1893 27876
rect 1893 27874 1899 27876
rect 1914 27924 1931 27926
rect 1931 27924 1965 27926
rect 1965 27924 1966 27926
rect 1914 27876 1966 27924
rect 1914 27874 1931 27876
rect 1931 27874 1965 27876
rect 1965 27874 1966 27876
rect 1981 27924 2003 27926
rect 2003 27924 2033 27926
rect 12157 27940 12189 27958
rect 12189 27940 12209 27958
rect 12225 27958 12277 27992
rect 12225 27940 12227 27958
rect 12227 27940 12261 27958
rect 12261 27940 12277 27958
rect 12293 27958 12345 27992
rect 12293 27940 12299 27958
rect 12299 27940 12333 27958
rect 12333 27940 12345 27958
rect 12361 27958 12413 27992
rect 12361 27940 12371 27958
rect 12371 27940 12405 27958
rect 12405 27940 12413 27958
rect 12429 27958 12481 27992
rect 12429 27940 12443 27958
rect 12443 27940 12477 27958
rect 12477 27940 12481 27958
rect 12497 27958 12549 27992
rect 12497 27940 12515 27958
rect 12515 27940 12549 27958
rect 12565 27958 12617 27992
rect 12633 27958 12685 27992
rect 12701 27958 12753 27992
rect 12768 27958 12820 27992
rect 12835 27958 12887 27992
rect 12565 27940 12587 27958
rect 12587 27940 12617 27958
rect 12633 27940 12659 27958
rect 12659 27940 12685 27958
rect 12701 27940 12731 27958
rect 12731 27940 12753 27958
rect 12768 27940 12803 27958
rect 12803 27940 12820 27958
rect 12835 27940 12837 27958
rect 12837 27940 12875 27958
rect 12875 27940 12887 27958
rect 12157 27924 12189 27926
rect 12189 27924 12209 27926
rect 1981 27876 2033 27924
rect 12157 27876 12209 27924
rect 1981 27874 2003 27876
rect 2003 27874 2033 27876
rect 1303 27842 1314 27860
rect 1314 27842 1353 27860
rect 1353 27842 1355 27860
rect 1371 27842 1387 27860
rect 1387 27842 1423 27860
rect 1439 27842 1460 27860
rect 1460 27842 1491 27860
rect 1507 27842 1533 27860
rect 1533 27842 1559 27860
rect 1575 27842 1605 27860
rect 1605 27842 1627 27860
rect 1303 27808 1355 27842
rect 1371 27808 1423 27842
rect 1439 27808 1491 27842
rect 1507 27808 1559 27842
rect 1575 27808 1627 27842
rect 1643 27842 1677 27860
rect 1677 27842 1695 27860
rect 1643 27808 1695 27842
rect 1711 27842 1715 27860
rect 1715 27842 1749 27860
rect 1749 27842 1763 27860
rect 1711 27808 1763 27842
rect 1779 27842 1787 27860
rect 1787 27842 1821 27860
rect 1821 27842 1831 27860
rect 1779 27808 1831 27842
rect 1847 27842 1859 27860
rect 1859 27842 1893 27860
rect 1893 27842 1899 27860
rect 1847 27808 1899 27842
rect 1914 27842 1931 27860
rect 1931 27842 1965 27860
rect 1965 27842 1966 27860
rect 1914 27808 1966 27842
rect 1981 27842 2003 27860
rect 2003 27842 2033 27860
rect 12157 27874 12189 27876
rect 12189 27874 12209 27876
rect 12225 27924 12227 27926
rect 12227 27924 12261 27926
rect 12261 27924 12277 27926
rect 12225 27876 12277 27924
rect 12225 27874 12227 27876
rect 12227 27874 12261 27876
rect 12261 27874 12277 27876
rect 12293 27924 12299 27926
rect 12299 27924 12333 27926
rect 12333 27924 12345 27926
rect 12293 27876 12345 27924
rect 12293 27874 12299 27876
rect 12299 27874 12333 27876
rect 12333 27874 12345 27876
rect 12361 27924 12371 27926
rect 12371 27924 12405 27926
rect 12405 27924 12413 27926
rect 12361 27876 12413 27924
rect 12361 27874 12371 27876
rect 12371 27874 12405 27876
rect 12405 27874 12413 27876
rect 12429 27924 12443 27926
rect 12443 27924 12477 27926
rect 12477 27924 12481 27926
rect 12429 27876 12481 27924
rect 12429 27874 12443 27876
rect 12443 27874 12477 27876
rect 12477 27874 12481 27876
rect 12497 27924 12515 27926
rect 12515 27924 12549 27926
rect 12497 27876 12549 27924
rect 12497 27874 12515 27876
rect 12515 27874 12549 27876
rect 12565 27924 12587 27926
rect 12587 27924 12617 27926
rect 12633 27924 12659 27926
rect 12659 27924 12685 27926
rect 12701 27924 12731 27926
rect 12731 27924 12753 27926
rect 12768 27924 12803 27926
rect 12803 27924 12820 27926
rect 12835 27924 12837 27926
rect 12837 27924 12875 27926
rect 12875 27924 12887 27926
rect 12565 27876 12617 27924
rect 12633 27876 12685 27924
rect 12701 27876 12753 27924
rect 12768 27876 12820 27924
rect 12835 27876 12887 27924
rect 12565 27874 12587 27876
rect 12587 27874 12617 27876
rect 12633 27874 12659 27876
rect 12659 27874 12685 27876
rect 12701 27874 12731 27876
rect 12731 27874 12753 27876
rect 12768 27874 12803 27876
rect 12803 27874 12820 27876
rect 12835 27874 12837 27876
rect 12837 27874 12875 27876
rect 12875 27874 12887 27876
rect 12157 27842 12189 27860
rect 12189 27842 12209 27860
rect 1981 27808 2033 27842
rect 12157 27808 12209 27842
rect 12225 27842 12227 27860
rect 12227 27842 12261 27860
rect 12261 27842 12277 27860
rect 12225 27808 12277 27842
rect 12293 27842 12299 27860
rect 12299 27842 12333 27860
rect 12333 27842 12345 27860
rect 12293 27808 12345 27842
rect 12361 27842 12371 27860
rect 12371 27842 12405 27860
rect 12405 27842 12413 27860
rect 12361 27808 12413 27842
rect 12429 27842 12443 27860
rect 12443 27842 12477 27860
rect 12477 27842 12481 27860
rect 12429 27808 12481 27842
rect 12497 27842 12515 27860
rect 12515 27842 12549 27860
rect 12497 27808 12549 27842
rect 12565 27842 12587 27860
rect 12587 27842 12617 27860
rect 12633 27842 12659 27860
rect 12659 27842 12685 27860
rect 12701 27842 12731 27860
rect 12731 27842 12753 27860
rect 12768 27842 12803 27860
rect 12803 27842 12820 27860
rect 12835 27842 12837 27860
rect 12837 27842 12875 27860
rect 12875 27842 12887 27860
rect 12565 27808 12617 27842
rect 12633 27808 12685 27842
rect 12701 27808 12753 27842
rect 12768 27808 12820 27842
rect 12835 27808 12887 27842
rect 1303 27760 1314 27794
rect 1314 27760 1353 27794
rect 1353 27760 1355 27794
rect 1371 27760 1387 27794
rect 1387 27760 1423 27794
rect 1439 27760 1460 27794
rect 1460 27760 1491 27794
rect 1507 27760 1533 27794
rect 1533 27760 1559 27794
rect 1575 27760 1605 27794
rect 1605 27760 1627 27794
rect 1303 27742 1355 27760
rect 1371 27742 1423 27760
rect 1439 27742 1491 27760
rect 1507 27742 1559 27760
rect 1575 27742 1627 27760
rect 1643 27760 1677 27794
rect 1677 27760 1695 27794
rect 1643 27742 1695 27760
rect 1711 27760 1715 27794
rect 1715 27760 1749 27794
rect 1749 27760 1763 27794
rect 1711 27742 1763 27760
rect 1779 27760 1787 27794
rect 1787 27760 1821 27794
rect 1821 27760 1831 27794
rect 1779 27742 1831 27760
rect 1847 27760 1859 27794
rect 1859 27760 1893 27794
rect 1893 27760 1899 27794
rect 1847 27742 1899 27760
rect 1914 27760 1931 27794
rect 1931 27760 1965 27794
rect 1965 27760 1966 27794
rect 1914 27742 1966 27760
rect 1981 27760 2003 27794
rect 2003 27760 2033 27794
rect 12157 27760 12189 27794
rect 12189 27760 12209 27794
rect 1981 27742 2033 27760
rect 12157 27742 12209 27760
rect 12225 27760 12227 27794
rect 12227 27760 12261 27794
rect 12261 27760 12277 27794
rect 12225 27742 12277 27760
rect 12293 27760 12299 27794
rect 12299 27760 12333 27794
rect 12333 27760 12345 27794
rect 12293 27742 12345 27760
rect 12361 27760 12371 27794
rect 12371 27760 12405 27794
rect 12405 27760 12413 27794
rect 12361 27742 12413 27760
rect 12429 27760 12443 27794
rect 12443 27760 12477 27794
rect 12477 27760 12481 27794
rect 12429 27742 12481 27760
rect 12497 27760 12515 27794
rect 12515 27760 12549 27794
rect 12497 27742 12549 27760
rect 12565 27760 12587 27794
rect 12587 27760 12617 27794
rect 12633 27760 12659 27794
rect 12659 27760 12685 27794
rect 12701 27760 12731 27794
rect 12731 27760 12753 27794
rect 12768 27760 12803 27794
rect 12803 27760 12820 27794
rect 12835 27760 12837 27794
rect 12837 27760 12875 27794
rect 12875 27760 12887 27794
rect 12565 27742 12617 27760
rect 12633 27742 12685 27760
rect 12701 27742 12753 27760
rect 12768 27742 12820 27760
rect 12835 27742 12887 27760
rect 1303 27712 1355 27728
rect 1371 27712 1423 27728
rect 1439 27712 1491 27728
rect 1507 27712 1559 27728
rect 1575 27712 1627 27728
rect 1303 27678 1314 27712
rect 1314 27678 1353 27712
rect 1353 27678 1355 27712
rect 1371 27678 1387 27712
rect 1387 27678 1423 27712
rect 1439 27678 1460 27712
rect 1460 27678 1491 27712
rect 1507 27678 1533 27712
rect 1533 27678 1559 27712
rect 1575 27678 1605 27712
rect 1605 27678 1627 27712
rect 1303 27676 1355 27678
rect 1371 27676 1423 27678
rect 1439 27676 1491 27678
rect 1507 27676 1559 27678
rect 1575 27676 1627 27678
rect 1643 27712 1695 27728
rect 1643 27678 1677 27712
rect 1677 27678 1695 27712
rect 1643 27676 1695 27678
rect 1711 27712 1763 27728
rect 1711 27678 1715 27712
rect 1715 27678 1749 27712
rect 1749 27678 1763 27712
rect 1711 27676 1763 27678
rect 1779 27712 1831 27728
rect 1779 27678 1787 27712
rect 1787 27678 1821 27712
rect 1821 27678 1831 27712
rect 1779 27676 1831 27678
rect 1847 27712 1899 27728
rect 1847 27678 1859 27712
rect 1859 27678 1893 27712
rect 1893 27678 1899 27712
rect 1847 27676 1899 27678
rect 1914 27712 1966 27728
rect 1914 27678 1931 27712
rect 1931 27678 1965 27712
rect 1965 27678 1966 27712
rect 1914 27676 1966 27678
rect 1981 27712 2033 27728
rect 12157 27712 12209 27728
rect 1981 27678 2003 27712
rect 2003 27678 2033 27712
rect 12157 27678 12189 27712
rect 12189 27678 12209 27712
rect 1981 27676 2033 27678
rect 12157 27676 12209 27678
rect 12225 27712 12277 27728
rect 12225 27678 12227 27712
rect 12227 27678 12261 27712
rect 12261 27678 12277 27712
rect 12225 27676 12277 27678
rect 12293 27712 12345 27728
rect 12293 27678 12299 27712
rect 12299 27678 12333 27712
rect 12333 27678 12345 27712
rect 12293 27676 12345 27678
rect 12361 27712 12413 27728
rect 12361 27678 12371 27712
rect 12371 27678 12405 27712
rect 12405 27678 12413 27712
rect 12361 27676 12413 27678
rect 12429 27712 12481 27728
rect 12429 27678 12443 27712
rect 12443 27678 12477 27712
rect 12477 27678 12481 27712
rect 12429 27676 12481 27678
rect 12497 27712 12549 27728
rect 12497 27678 12515 27712
rect 12515 27678 12549 27712
rect 12497 27676 12549 27678
rect 12565 27712 12617 27728
rect 12633 27712 12685 27728
rect 12701 27712 12753 27728
rect 12768 27712 12820 27728
rect 12835 27712 12887 27728
rect 12565 27678 12587 27712
rect 12587 27678 12617 27712
rect 12633 27678 12659 27712
rect 12659 27678 12685 27712
rect 12701 27678 12731 27712
rect 12731 27678 12753 27712
rect 12768 27678 12803 27712
rect 12803 27678 12820 27712
rect 12835 27678 12837 27712
rect 12837 27678 12875 27712
rect 12875 27678 12887 27712
rect 12565 27676 12617 27678
rect 12633 27676 12685 27678
rect 12701 27676 12753 27678
rect 12768 27676 12820 27678
rect 12835 27676 12887 27678
rect 14282 28119 14334 28171
rect 14358 28119 14410 28171
rect 14434 28119 14486 28171
rect 14510 28119 14562 28171
rect 14586 28119 14638 28171
rect 14282 28053 14334 28105
rect 14358 28053 14410 28105
rect 14434 28053 14486 28105
rect 14510 28053 14562 28105
rect 14586 28053 14638 28105
rect 14282 27987 14334 28039
rect 14358 27987 14410 28039
rect 14434 27987 14486 28039
rect 14510 27987 14562 28039
rect 14586 27987 14638 28039
rect 14282 27921 14334 27973
rect 14358 27921 14410 27973
rect 14434 27921 14486 27973
rect 14510 27921 14562 27973
rect 14586 27921 14638 27973
rect 14282 27855 14334 27907
rect 14358 27855 14410 27907
rect 14434 27855 14486 27907
rect 14510 27855 14562 27907
rect 14586 27855 14638 27907
rect 14282 27789 14334 27841
rect 14358 27789 14410 27841
rect 14434 27789 14486 27841
rect 14510 27789 14562 27841
rect 14586 27789 14638 27841
rect 14282 27723 14334 27775
rect 14358 27723 14410 27775
rect 14434 27723 14486 27775
rect 14510 27723 14562 27775
rect 14586 27723 14638 27775
rect 14282 27657 14334 27709
rect 14358 27657 14410 27709
rect 14434 27657 14486 27709
rect 14510 27657 14562 27709
rect 14586 27657 14638 27709
rect 14282 27591 14334 27643
rect 14358 27591 14410 27643
rect 14434 27591 14486 27643
rect 14510 27591 14562 27643
rect 14586 27591 14638 27643
rect 14282 27525 14334 27577
rect 14358 27525 14410 27577
rect 14434 27525 14486 27577
rect 14510 27525 14562 27577
rect 14586 27525 14638 27577
rect 14282 27459 14334 27511
rect 14358 27459 14410 27511
rect 14434 27459 14486 27511
rect 14510 27459 14562 27511
rect 14586 27459 14638 27511
rect 14282 27393 14334 27445
rect 14358 27393 14410 27445
rect 14434 27393 14486 27445
rect 14510 27393 14562 27445
rect 14586 27393 14638 27445
rect 3478 27362 3530 27369
rect 3546 27362 3598 27369
rect 3614 27362 3666 27369
rect 3478 27328 3499 27362
rect 3499 27328 3530 27362
rect 3546 27328 3572 27362
rect 3572 27328 3598 27362
rect 3614 27328 3645 27362
rect 3645 27328 3666 27362
rect 3478 27317 3530 27328
rect 3546 27317 3598 27328
rect 3614 27317 3666 27328
rect 3682 27362 3734 27369
rect 3682 27328 3684 27362
rect 3684 27328 3718 27362
rect 3718 27328 3734 27362
rect 3682 27317 3734 27328
rect 3750 27362 3802 27369
rect 3750 27328 3757 27362
rect 3757 27328 3791 27362
rect 3791 27328 3802 27362
rect 3750 27317 3802 27328
rect 3818 27362 3870 27369
rect 3818 27328 3830 27362
rect 3830 27328 3864 27362
rect 3864 27328 3870 27362
rect 3818 27317 3870 27328
rect 3886 27362 3938 27369
rect 3886 27328 3903 27362
rect 3903 27328 3937 27362
rect 3937 27328 3938 27362
rect 3886 27317 3938 27328
rect 3954 27362 4006 27369
rect 4021 27362 4073 27369
rect 4088 27362 4140 27369
rect 4155 27362 4207 27369
rect 4222 27362 4274 27369
rect 4289 27362 4341 27369
rect 4356 27362 4408 27369
rect 4423 27362 4475 27369
rect 4490 27362 4542 27369
rect 4557 27362 4609 27369
rect 5461 27362 5513 27369
rect 5529 27362 5581 27369
rect 5597 27362 5649 27369
rect 5665 27362 5717 27369
rect 5733 27362 5785 27369
rect 5801 27362 5853 27369
rect 5869 27362 5921 27369
rect 5937 27362 5989 27369
rect 6004 27362 6056 27369
rect 6071 27362 6123 27369
rect 3954 27328 3976 27362
rect 3976 27328 4006 27362
rect 4021 27328 4049 27362
rect 4049 27328 4073 27362
rect 4088 27328 4122 27362
rect 4122 27328 4140 27362
rect 4155 27328 4156 27362
rect 4156 27328 4194 27362
rect 4194 27328 4207 27362
rect 4222 27328 4228 27362
rect 4228 27328 4266 27362
rect 4266 27328 4274 27362
rect 4289 27328 4300 27362
rect 4300 27328 4338 27362
rect 4338 27328 4341 27362
rect 4356 27328 4372 27362
rect 4372 27328 4408 27362
rect 4423 27328 4444 27362
rect 4444 27328 4475 27362
rect 4490 27328 4516 27362
rect 4516 27328 4542 27362
rect 4557 27328 4588 27362
rect 4588 27328 4609 27362
rect 5461 27328 5490 27362
rect 5490 27328 5513 27362
rect 5529 27328 5562 27362
rect 5562 27328 5581 27362
rect 5597 27328 5634 27362
rect 5634 27328 5649 27362
rect 5665 27328 5668 27362
rect 5668 27328 5706 27362
rect 5706 27328 5717 27362
rect 5733 27328 5740 27362
rect 5740 27328 5778 27362
rect 5778 27328 5785 27362
rect 5801 27328 5812 27362
rect 5812 27328 5850 27362
rect 5850 27328 5853 27362
rect 5869 27328 5884 27362
rect 5884 27328 5921 27362
rect 5937 27328 5956 27362
rect 5956 27328 5989 27362
rect 6004 27328 6028 27362
rect 6028 27328 6056 27362
rect 6071 27328 6100 27362
rect 6100 27328 6123 27362
rect 3954 27317 4006 27328
rect 4021 27317 4073 27328
rect 4088 27317 4140 27328
rect 4155 27317 4207 27328
rect 4222 27317 4274 27328
rect 4289 27317 4341 27328
rect 4356 27317 4408 27328
rect 4423 27317 4475 27328
rect 4490 27317 4542 27328
rect 4557 27317 4609 27328
rect 5461 27317 5513 27328
rect 5529 27317 5581 27328
rect 5597 27317 5649 27328
rect 5665 27317 5717 27328
rect 5733 27317 5785 27328
rect 5801 27317 5853 27328
rect 5869 27317 5921 27328
rect 5937 27317 5989 27328
rect 6004 27317 6056 27328
rect 6071 27317 6123 27328
rect 6138 27362 6190 27369
rect 6138 27328 6172 27362
rect 6172 27328 6190 27362
rect 6138 27317 6190 27328
rect 6205 27362 6257 27369
rect 6205 27328 6210 27362
rect 6210 27328 6244 27362
rect 6244 27328 6257 27362
rect 6205 27317 6257 27328
rect 6272 27362 6324 27369
rect 6272 27328 6282 27362
rect 6282 27328 6316 27362
rect 6316 27328 6324 27362
rect 6272 27317 6324 27328
rect 6339 27362 6391 27369
rect 6339 27328 6354 27362
rect 6354 27328 6388 27362
rect 6388 27328 6391 27362
rect 6339 27317 6391 27328
rect 6406 27362 6458 27369
rect 6473 27362 6525 27369
rect 6540 27362 6592 27369
rect 7445 27362 7497 27369
rect 7513 27362 7565 27369
rect 7581 27362 7633 27369
rect 6406 27328 6426 27362
rect 6426 27328 6458 27362
rect 6473 27328 6498 27362
rect 6498 27328 6525 27362
rect 6540 27328 6570 27362
rect 6570 27328 6592 27362
rect 7445 27328 7468 27362
rect 7468 27328 7497 27362
rect 7513 27328 7540 27362
rect 7540 27328 7565 27362
rect 7581 27328 7612 27362
rect 7612 27328 7633 27362
rect 6406 27317 6458 27328
rect 6473 27317 6525 27328
rect 6540 27317 6592 27328
rect 7445 27317 7497 27328
rect 7513 27317 7565 27328
rect 7581 27317 7633 27328
rect 7649 27362 7701 27369
rect 7649 27328 7650 27362
rect 7650 27328 7684 27362
rect 7684 27328 7701 27362
rect 7649 27317 7701 27328
rect 7717 27362 7769 27369
rect 7717 27328 7722 27362
rect 7722 27328 7756 27362
rect 7756 27328 7769 27362
rect 7717 27317 7769 27328
rect 7785 27362 7837 27369
rect 7785 27328 7794 27362
rect 7794 27328 7828 27362
rect 7828 27328 7837 27362
rect 7785 27317 7837 27328
rect 7853 27362 7905 27369
rect 7853 27328 7866 27362
rect 7866 27328 7900 27362
rect 7900 27328 7905 27362
rect 7853 27317 7905 27328
rect 7921 27362 7973 27369
rect 7921 27328 7938 27362
rect 7938 27328 7972 27362
rect 7972 27328 7973 27362
rect 7921 27317 7973 27328
rect 7988 27362 8040 27369
rect 8055 27362 8107 27369
rect 8122 27362 8174 27369
rect 8189 27362 8241 27369
rect 8256 27362 8308 27369
rect 8323 27362 8375 27369
rect 8390 27362 8442 27369
rect 8457 27362 8509 27369
rect 8524 27362 8576 27369
rect 9423 27362 9475 27364
rect 9523 27362 9575 27364
rect 14282 27362 14334 27379
rect 14358 27362 14410 27379
rect 14434 27362 14486 27379
rect 14510 27362 14562 27379
rect 14586 27362 14638 27379
rect 7988 27328 8010 27362
rect 8010 27328 8040 27362
rect 8055 27328 8082 27362
rect 8082 27328 8107 27362
rect 8122 27328 8154 27362
rect 8154 27328 8174 27362
rect 8189 27328 8226 27362
rect 8226 27328 8241 27362
rect 8256 27328 8260 27362
rect 8260 27328 8298 27362
rect 8298 27328 8308 27362
rect 8323 27328 8332 27362
rect 8332 27328 8370 27362
rect 8370 27328 8375 27362
rect 8390 27328 8404 27362
rect 8404 27328 8442 27362
rect 8457 27328 8476 27362
rect 8476 27328 8509 27362
rect 8524 27328 8548 27362
rect 8548 27328 8576 27362
rect 9423 27328 9450 27362
rect 9450 27328 9475 27362
rect 9523 27328 9556 27362
rect 9556 27328 9575 27362
rect 14282 27328 14308 27362
rect 14308 27328 14334 27362
rect 14358 27328 14380 27362
rect 14380 27328 14410 27362
rect 14434 27328 14452 27362
rect 14452 27328 14486 27362
rect 14510 27328 14524 27362
rect 14524 27328 14562 27362
rect 14586 27328 14596 27362
rect 14596 27328 14634 27362
rect 14634 27328 14638 27362
rect 7988 27317 8040 27328
rect 8055 27317 8107 27328
rect 8122 27317 8174 27328
rect 8189 27317 8241 27328
rect 8256 27317 8308 27328
rect 8323 27317 8375 27328
rect 8390 27317 8442 27328
rect 8457 27317 8509 27328
rect 8524 27317 8576 27328
rect 9423 27312 9475 27328
rect 9523 27312 9575 27328
rect 14282 27327 14334 27328
rect 14358 27327 14410 27328
rect 14434 27327 14486 27328
rect 14510 27327 14562 27328
rect 14586 27327 14638 27328
rect 3478 27238 3530 27243
rect 3546 27238 3598 27243
rect 3614 27238 3666 27243
rect 3478 27204 3499 27238
rect 3499 27204 3530 27238
rect 3546 27204 3572 27238
rect 3572 27204 3598 27238
rect 3614 27204 3645 27238
rect 3645 27204 3666 27238
rect 3478 27191 3530 27204
rect 3546 27191 3598 27204
rect 3614 27191 3666 27204
rect 3682 27238 3734 27243
rect 3682 27204 3684 27238
rect 3684 27204 3718 27238
rect 3718 27204 3734 27238
rect 3682 27191 3734 27204
rect 3750 27238 3802 27243
rect 3750 27204 3757 27238
rect 3757 27204 3791 27238
rect 3791 27204 3802 27238
rect 3750 27191 3802 27204
rect 3818 27238 3870 27243
rect 3818 27204 3830 27238
rect 3830 27204 3864 27238
rect 3864 27204 3870 27238
rect 3818 27191 3870 27204
rect 3886 27238 3938 27243
rect 3886 27204 3903 27238
rect 3903 27204 3937 27238
rect 3937 27204 3938 27238
rect 3886 27191 3938 27204
rect 3954 27238 4006 27243
rect 4021 27238 4073 27243
rect 4088 27238 4140 27243
rect 4155 27238 4207 27243
rect 4222 27238 4274 27243
rect 4289 27238 4341 27243
rect 4356 27238 4408 27243
rect 4423 27238 4475 27243
rect 4490 27238 4542 27243
rect 4557 27238 4609 27243
rect 5461 27238 5513 27243
rect 5529 27238 5581 27243
rect 5597 27238 5649 27243
rect 5665 27238 5717 27243
rect 5733 27238 5785 27243
rect 5801 27238 5853 27243
rect 5869 27238 5921 27243
rect 5937 27238 5989 27243
rect 6004 27238 6056 27243
rect 6071 27238 6123 27243
rect 3954 27204 3976 27238
rect 3976 27204 4006 27238
rect 4021 27204 4049 27238
rect 4049 27204 4073 27238
rect 4088 27204 4122 27238
rect 4122 27204 4140 27238
rect 4155 27204 4156 27238
rect 4156 27204 4194 27238
rect 4194 27204 4207 27238
rect 4222 27204 4228 27238
rect 4228 27204 4266 27238
rect 4266 27204 4274 27238
rect 4289 27204 4300 27238
rect 4300 27204 4338 27238
rect 4338 27204 4341 27238
rect 4356 27204 4372 27238
rect 4372 27204 4408 27238
rect 4423 27204 4444 27238
rect 4444 27204 4475 27238
rect 4490 27204 4516 27238
rect 4516 27204 4542 27238
rect 4557 27204 4588 27238
rect 4588 27204 4609 27238
rect 5461 27204 5490 27238
rect 5490 27204 5513 27238
rect 5529 27204 5562 27238
rect 5562 27204 5581 27238
rect 5597 27204 5634 27238
rect 5634 27204 5649 27238
rect 5665 27204 5668 27238
rect 5668 27204 5706 27238
rect 5706 27204 5717 27238
rect 5733 27204 5740 27238
rect 5740 27204 5778 27238
rect 5778 27204 5785 27238
rect 5801 27204 5812 27238
rect 5812 27204 5850 27238
rect 5850 27204 5853 27238
rect 5869 27204 5884 27238
rect 5884 27204 5921 27238
rect 5937 27204 5956 27238
rect 5956 27204 5989 27238
rect 6004 27204 6028 27238
rect 6028 27204 6056 27238
rect 6071 27204 6100 27238
rect 6100 27204 6123 27238
rect 3954 27191 4006 27204
rect 4021 27191 4073 27204
rect 4088 27191 4140 27204
rect 4155 27191 4207 27204
rect 4222 27191 4274 27204
rect 4289 27191 4341 27204
rect 4356 27191 4408 27204
rect 4423 27191 4475 27204
rect 4490 27191 4542 27204
rect 4557 27191 4609 27204
rect 5461 27191 5513 27204
rect 5529 27191 5581 27204
rect 5597 27191 5649 27204
rect 5665 27191 5717 27204
rect 5733 27191 5785 27204
rect 5801 27191 5853 27204
rect 5869 27191 5921 27204
rect 5937 27191 5989 27204
rect 6004 27191 6056 27204
rect 6071 27191 6123 27204
rect 6138 27238 6190 27243
rect 6138 27204 6172 27238
rect 6172 27204 6190 27238
rect 6138 27191 6190 27204
rect 6205 27238 6257 27243
rect 6205 27204 6210 27238
rect 6210 27204 6244 27238
rect 6244 27204 6257 27238
rect 6205 27191 6257 27204
rect 6272 27238 6324 27243
rect 6272 27204 6282 27238
rect 6282 27204 6316 27238
rect 6316 27204 6324 27238
rect 6272 27191 6324 27204
rect 6339 27238 6391 27243
rect 6339 27204 6354 27238
rect 6354 27204 6388 27238
rect 6388 27204 6391 27238
rect 6339 27191 6391 27204
rect 6406 27238 6458 27243
rect 6473 27238 6525 27243
rect 6540 27238 6592 27243
rect 7445 27238 7497 27243
rect 7513 27238 7565 27243
rect 7581 27238 7633 27243
rect 6406 27204 6426 27238
rect 6426 27204 6458 27238
rect 6473 27204 6498 27238
rect 6498 27204 6525 27238
rect 6540 27204 6570 27238
rect 6570 27204 6592 27238
rect 7445 27204 7468 27238
rect 7468 27204 7497 27238
rect 7513 27204 7540 27238
rect 7540 27204 7565 27238
rect 7581 27204 7612 27238
rect 7612 27204 7633 27238
rect 6406 27191 6458 27204
rect 6473 27191 6525 27204
rect 6540 27191 6592 27204
rect 7445 27191 7497 27204
rect 7513 27191 7565 27204
rect 7581 27191 7633 27204
rect 7649 27238 7701 27243
rect 7649 27204 7650 27238
rect 7650 27204 7684 27238
rect 7684 27204 7701 27238
rect 7649 27191 7701 27204
rect 7717 27238 7769 27243
rect 7717 27204 7722 27238
rect 7722 27204 7756 27238
rect 7756 27204 7769 27238
rect 7717 27191 7769 27204
rect 7785 27238 7837 27243
rect 7785 27204 7794 27238
rect 7794 27204 7828 27238
rect 7828 27204 7837 27238
rect 7785 27191 7837 27204
rect 7853 27238 7905 27243
rect 7853 27204 7866 27238
rect 7866 27204 7900 27238
rect 7900 27204 7905 27238
rect 7853 27191 7905 27204
rect 7921 27238 7973 27243
rect 7921 27204 7938 27238
rect 7938 27204 7972 27238
rect 7972 27204 7973 27238
rect 7921 27191 7973 27204
rect 7988 27238 8040 27243
rect 8055 27238 8107 27243
rect 8122 27238 8174 27243
rect 8189 27238 8241 27243
rect 8256 27238 8308 27243
rect 8323 27238 8375 27243
rect 8390 27238 8442 27243
rect 8457 27238 8509 27243
rect 8524 27238 8576 27243
rect 9423 27238 9475 27268
rect 9523 27238 9575 27268
rect 14282 27261 14334 27313
rect 14358 27261 14410 27313
rect 14434 27261 14486 27313
rect 14510 27261 14562 27313
rect 14586 27261 14638 27313
rect 14282 27238 14334 27247
rect 14358 27238 14410 27247
rect 14434 27238 14486 27247
rect 14510 27238 14562 27247
rect 14586 27238 14638 27247
rect 7988 27204 8010 27238
rect 8010 27204 8040 27238
rect 8055 27204 8082 27238
rect 8082 27204 8107 27238
rect 8122 27204 8154 27238
rect 8154 27204 8174 27238
rect 8189 27204 8226 27238
rect 8226 27204 8241 27238
rect 8256 27204 8260 27238
rect 8260 27204 8298 27238
rect 8298 27204 8308 27238
rect 8323 27204 8332 27238
rect 8332 27204 8370 27238
rect 8370 27204 8375 27238
rect 8390 27204 8404 27238
rect 8404 27204 8442 27238
rect 8457 27204 8476 27238
rect 8476 27204 8509 27238
rect 8524 27204 8548 27238
rect 8548 27204 8576 27238
rect 9423 27216 9450 27238
rect 9450 27216 9475 27238
rect 9523 27216 9556 27238
rect 9556 27216 9575 27238
rect 14282 27204 14308 27238
rect 14308 27204 14334 27238
rect 14358 27204 14380 27238
rect 14380 27204 14410 27238
rect 14434 27204 14452 27238
rect 14452 27204 14486 27238
rect 14510 27204 14524 27238
rect 14524 27204 14562 27238
rect 14586 27204 14596 27238
rect 14596 27204 14634 27238
rect 14634 27204 14638 27238
rect 7988 27191 8040 27204
rect 8055 27191 8107 27204
rect 8122 27191 8174 27204
rect 8189 27191 8241 27204
rect 8256 27191 8308 27204
rect 8323 27191 8375 27204
rect 8390 27191 8442 27204
rect 8457 27191 8509 27204
rect 8524 27191 8576 27204
rect 14282 27195 14334 27204
rect 14358 27195 14410 27204
rect 14434 27195 14486 27204
rect 14510 27195 14562 27204
rect 14586 27195 14638 27204
rect 2365 26948 2417 27000
rect 2440 26948 2492 27000
rect 2515 26948 2567 27000
rect 2589 26948 2641 27000
rect 2663 26948 2715 27000
rect 2365 26826 2417 26878
rect 2440 26826 2492 26878
rect 2515 26826 2567 26878
rect 2589 26826 2641 26878
rect 2663 26826 2715 26878
rect 2480 26151 2506 26181
rect 2506 26151 2532 26181
rect 2550 26151 2579 26181
rect 2579 26151 2602 26181
rect 2620 26151 2652 26181
rect 2652 26151 2672 26181
rect 3472 26151 3489 26181
rect 3489 26151 3524 26181
rect 3542 26151 3562 26181
rect 3562 26151 3594 26181
rect 3612 26151 3635 26181
rect 3635 26151 3664 26181
rect 4464 26151 4466 26181
rect 4466 26151 4500 26181
rect 4500 26151 4516 26181
rect 2480 26129 2532 26151
rect 2550 26129 2602 26151
rect 2620 26129 2672 26151
rect 3472 26129 3524 26151
rect 3542 26129 3594 26151
rect 3612 26129 3664 26151
rect 4464 26129 4516 26151
rect 4534 26151 4538 26181
rect 4538 26151 4572 26181
rect 4572 26151 4586 26181
rect 4534 26129 4586 26151
rect 4604 26151 4610 26181
rect 4610 26151 4644 26181
rect 4644 26151 4656 26181
rect 5456 26151 5474 26181
rect 5474 26151 5508 26181
rect 4604 26129 4656 26151
rect 5456 26129 5508 26151
rect 5526 26151 5546 26181
rect 5546 26151 5578 26181
rect 5596 26151 5618 26181
rect 5618 26151 5648 26181
rect 6448 26151 6482 26181
rect 6482 26151 6500 26181
rect 6518 26151 6554 26181
rect 6554 26151 6570 26181
rect 6588 26151 6626 26181
rect 6626 26151 6640 26181
rect 7440 26151 7452 26181
rect 7452 26151 7490 26181
rect 7490 26151 7492 26181
rect 7510 26151 7524 26181
rect 7524 26151 7562 26181
rect 7580 26151 7596 26181
rect 7596 26151 7632 26181
rect 8432 26151 8460 26181
rect 8460 26151 8484 26181
rect 8502 26151 8532 26181
rect 8532 26151 8554 26181
rect 8572 26151 8604 26181
rect 8604 26151 8624 26181
rect 9424 26151 9434 26181
rect 9434 26151 9468 26181
rect 9468 26151 9476 26181
rect 5526 26129 5578 26151
rect 5596 26129 5648 26151
rect 6448 26129 6500 26151
rect 6518 26129 6570 26151
rect 6588 26129 6640 26151
rect 7440 26129 7492 26151
rect 7510 26129 7562 26151
rect 7580 26129 7632 26151
rect 8432 26129 8484 26151
rect 8502 26129 8554 26151
rect 8572 26129 8624 26151
rect 9424 26129 9476 26151
rect 9494 26151 9506 26181
rect 9506 26151 9540 26181
rect 9540 26151 9546 26181
rect 9494 26129 9546 26151
rect 9564 26151 9578 26181
rect 9578 26151 9612 26181
rect 9612 26151 9616 26181
rect 9564 26129 9616 26151
rect 2480 26077 2506 26111
rect 2506 26077 2532 26111
rect 2550 26077 2579 26111
rect 2579 26077 2602 26111
rect 2620 26077 2652 26111
rect 2652 26077 2672 26111
rect 3472 26077 3489 26111
rect 3489 26077 3524 26111
rect 3542 26077 3562 26111
rect 3562 26077 3594 26111
rect 3612 26077 3635 26111
rect 3635 26077 3664 26111
rect 4464 26077 4466 26111
rect 4466 26077 4500 26111
rect 4500 26077 4516 26111
rect 2480 26059 2532 26077
rect 2550 26059 2602 26077
rect 2620 26059 2672 26077
rect 3472 26059 3524 26077
rect 3542 26059 3594 26077
rect 3612 26059 3664 26077
rect 4464 26059 4516 26077
rect 4534 26077 4538 26111
rect 4538 26077 4572 26111
rect 4572 26077 4586 26111
rect 4534 26059 4586 26077
rect 4604 26077 4610 26111
rect 4610 26077 4644 26111
rect 4644 26077 4656 26111
rect 5456 26077 5474 26111
rect 5474 26077 5508 26111
rect 4604 26059 4656 26077
rect 5456 26059 5508 26077
rect 5526 26077 5546 26111
rect 5546 26077 5578 26111
rect 5596 26077 5618 26111
rect 5618 26077 5648 26111
rect 6448 26077 6482 26111
rect 6482 26077 6500 26111
rect 6518 26077 6554 26111
rect 6554 26077 6570 26111
rect 6588 26077 6626 26111
rect 6626 26077 6640 26111
rect 7440 26077 7452 26111
rect 7452 26077 7490 26111
rect 7490 26077 7492 26111
rect 7510 26077 7524 26111
rect 7524 26077 7562 26111
rect 7580 26077 7596 26111
rect 7596 26077 7632 26111
rect 8432 26077 8460 26111
rect 8460 26077 8484 26111
rect 8502 26077 8532 26111
rect 8532 26077 8554 26111
rect 8572 26077 8604 26111
rect 8604 26077 8624 26111
rect 9424 26077 9434 26111
rect 9434 26077 9468 26111
rect 9468 26077 9476 26111
rect 5526 26059 5578 26077
rect 5596 26059 5648 26077
rect 6448 26059 6500 26077
rect 6518 26059 6570 26077
rect 6588 26059 6640 26077
rect 7440 26059 7492 26077
rect 7510 26059 7562 26077
rect 7580 26059 7632 26077
rect 8432 26059 8484 26077
rect 8502 26059 8554 26077
rect 8572 26059 8624 26077
rect 9424 26059 9476 26077
rect 9494 26077 9506 26111
rect 9506 26077 9540 26111
rect 9540 26077 9546 26111
rect 9494 26059 9546 26077
rect 9564 26077 9578 26111
rect 9578 26077 9612 26111
rect 9612 26077 9616 26111
rect 9564 26059 9616 26077
rect 2480 26037 2532 26041
rect 2550 26037 2602 26041
rect 2620 26037 2672 26041
rect 3472 26037 3524 26041
rect 3542 26037 3594 26041
rect 3612 26037 3664 26041
rect 4464 26037 4516 26041
rect 2480 26003 2506 26037
rect 2506 26003 2532 26037
rect 2550 26003 2579 26037
rect 2579 26003 2602 26037
rect 2620 26003 2652 26037
rect 2652 26003 2672 26037
rect 3472 26003 3489 26037
rect 3489 26003 3524 26037
rect 3542 26003 3562 26037
rect 3562 26003 3594 26037
rect 3612 26003 3635 26037
rect 3635 26003 3664 26037
rect 4464 26003 4466 26037
rect 4466 26003 4500 26037
rect 4500 26003 4516 26037
rect 2480 25989 2532 26003
rect 2550 25989 2602 26003
rect 2620 25989 2672 26003
rect 3472 25989 3524 26003
rect 3542 25989 3594 26003
rect 3612 25989 3664 26003
rect 4464 25989 4516 26003
rect 4534 26037 4586 26041
rect 4534 26003 4538 26037
rect 4538 26003 4572 26037
rect 4572 26003 4586 26037
rect 4534 25989 4586 26003
rect 4604 26037 4656 26041
rect 5456 26037 5508 26041
rect 4604 26003 4610 26037
rect 4610 26003 4644 26037
rect 4644 26003 4656 26037
rect 5456 26003 5474 26037
rect 5474 26003 5508 26037
rect 4604 25989 4656 26003
rect 5456 25989 5508 26003
rect 5526 26037 5578 26041
rect 5596 26037 5648 26041
rect 6448 26037 6500 26041
rect 6518 26037 6570 26041
rect 6588 26037 6640 26041
rect 7440 26037 7492 26041
rect 7510 26037 7562 26041
rect 7580 26037 7632 26041
rect 8432 26037 8484 26041
rect 8502 26037 8554 26041
rect 8572 26037 8624 26041
rect 9424 26037 9476 26041
rect 5526 26003 5546 26037
rect 5546 26003 5578 26037
rect 5596 26003 5618 26037
rect 5618 26003 5648 26037
rect 6448 26003 6482 26037
rect 6482 26003 6500 26037
rect 6518 26003 6554 26037
rect 6554 26003 6570 26037
rect 6588 26003 6626 26037
rect 6626 26003 6640 26037
rect 7440 26003 7452 26037
rect 7452 26003 7490 26037
rect 7490 26003 7492 26037
rect 7510 26003 7524 26037
rect 7524 26003 7562 26037
rect 7580 26003 7596 26037
rect 7596 26003 7632 26037
rect 8432 26003 8460 26037
rect 8460 26003 8484 26037
rect 8502 26003 8532 26037
rect 8532 26003 8554 26037
rect 8572 26003 8604 26037
rect 8604 26003 8624 26037
rect 9424 26003 9434 26037
rect 9434 26003 9468 26037
rect 9468 26003 9476 26037
rect 5526 25989 5578 26003
rect 5596 25989 5648 26003
rect 6448 25989 6500 26003
rect 6518 25989 6570 26003
rect 6588 25989 6640 26003
rect 7440 25989 7492 26003
rect 7510 25989 7562 26003
rect 7580 25989 7632 26003
rect 8432 25989 8484 26003
rect 8502 25989 8554 26003
rect 8572 25989 8624 26003
rect 9424 25989 9476 26003
rect 9494 26037 9546 26041
rect 9494 26003 9506 26037
rect 9506 26003 9540 26037
rect 9540 26003 9546 26037
rect 9494 25989 9546 26003
rect 9564 26037 9616 26041
rect 9564 26003 9578 26037
rect 9578 26003 9612 26037
rect 9612 26003 9616 26037
rect 9564 25989 9616 26003
rect 2480 25963 2532 25971
rect 2550 25963 2602 25971
rect 2620 25963 2672 25971
rect 3472 25963 3524 25971
rect 3542 25963 3594 25971
rect 3612 25963 3664 25971
rect 4464 25963 4516 25971
rect 2480 25929 2506 25963
rect 2506 25929 2532 25963
rect 2550 25929 2579 25963
rect 2579 25929 2602 25963
rect 2620 25929 2652 25963
rect 2652 25929 2672 25963
rect 3472 25929 3489 25963
rect 3489 25929 3524 25963
rect 3542 25929 3562 25963
rect 3562 25929 3594 25963
rect 3612 25929 3635 25963
rect 3635 25929 3664 25963
rect 4464 25929 4466 25963
rect 4466 25929 4500 25963
rect 4500 25929 4516 25963
rect 2480 25919 2532 25929
rect 2550 25919 2602 25929
rect 2620 25919 2672 25929
rect 3472 25919 3524 25929
rect 3542 25919 3594 25929
rect 3612 25919 3664 25929
rect 4464 25919 4516 25929
rect 4534 25963 4586 25971
rect 4534 25929 4538 25963
rect 4538 25929 4572 25963
rect 4572 25929 4586 25963
rect 4534 25919 4586 25929
rect 4604 25963 4656 25971
rect 5456 25963 5508 25971
rect 4604 25929 4610 25963
rect 4610 25929 4644 25963
rect 4644 25929 4656 25963
rect 5456 25929 5474 25963
rect 5474 25929 5508 25963
rect 4604 25919 4656 25929
rect 5456 25919 5508 25929
rect 5526 25963 5578 25971
rect 5596 25963 5648 25971
rect 6448 25963 6500 25971
rect 6518 25963 6570 25971
rect 6588 25963 6640 25971
rect 7440 25963 7492 25971
rect 7510 25963 7562 25971
rect 7580 25963 7632 25971
rect 8432 25963 8484 25971
rect 8502 25963 8554 25971
rect 8572 25963 8624 25971
rect 9424 25963 9476 25971
rect 5526 25929 5546 25963
rect 5546 25929 5578 25963
rect 5596 25929 5618 25963
rect 5618 25929 5648 25963
rect 6448 25929 6482 25963
rect 6482 25929 6500 25963
rect 6518 25929 6554 25963
rect 6554 25929 6570 25963
rect 6588 25929 6626 25963
rect 6626 25929 6640 25963
rect 7440 25929 7452 25963
rect 7452 25929 7490 25963
rect 7490 25929 7492 25963
rect 7510 25929 7524 25963
rect 7524 25929 7562 25963
rect 7580 25929 7596 25963
rect 7596 25929 7632 25963
rect 8432 25929 8460 25963
rect 8460 25929 8484 25963
rect 8502 25929 8532 25963
rect 8532 25929 8554 25963
rect 8572 25929 8604 25963
rect 8604 25929 8624 25963
rect 9424 25929 9434 25963
rect 9434 25929 9468 25963
rect 9468 25929 9476 25963
rect 5526 25919 5578 25929
rect 5596 25919 5648 25929
rect 6448 25919 6500 25929
rect 6518 25919 6570 25929
rect 6588 25919 6640 25929
rect 7440 25919 7492 25929
rect 7510 25919 7562 25929
rect 7580 25919 7632 25929
rect 8432 25919 8484 25929
rect 8502 25919 8554 25929
rect 8572 25919 8624 25929
rect 9424 25919 9476 25929
rect 9494 25963 9546 25971
rect 9494 25929 9506 25963
rect 9506 25929 9540 25963
rect 9540 25929 9546 25963
rect 9494 25919 9546 25929
rect 9564 25963 9616 25971
rect 9564 25929 9578 25963
rect 9578 25929 9612 25963
rect 9612 25929 9616 25963
rect 9564 25919 9616 25929
rect 2480 25889 2532 25901
rect 2550 25889 2602 25901
rect 2620 25889 2672 25901
rect 3472 25889 3524 25901
rect 3542 25889 3594 25901
rect 3612 25889 3664 25901
rect 4464 25889 4516 25901
rect 2480 25855 2506 25889
rect 2506 25855 2532 25889
rect 2550 25855 2579 25889
rect 2579 25855 2602 25889
rect 2620 25855 2652 25889
rect 2652 25855 2672 25889
rect 3472 25855 3489 25889
rect 3489 25855 3524 25889
rect 3542 25855 3562 25889
rect 3562 25855 3594 25889
rect 3612 25855 3635 25889
rect 3635 25855 3664 25889
rect 4464 25855 4466 25889
rect 4466 25855 4500 25889
rect 4500 25855 4516 25889
rect 2480 25849 2532 25855
rect 2550 25849 2602 25855
rect 2620 25849 2672 25855
rect 3472 25849 3524 25855
rect 3542 25849 3594 25855
rect 3612 25849 3664 25855
rect 4464 25849 4516 25855
rect 4534 25889 4586 25901
rect 4534 25855 4538 25889
rect 4538 25855 4572 25889
rect 4572 25855 4586 25889
rect 4534 25849 4586 25855
rect 4604 25889 4656 25901
rect 5456 25889 5508 25901
rect 4604 25855 4610 25889
rect 4610 25855 4644 25889
rect 4644 25855 4656 25889
rect 5456 25855 5474 25889
rect 5474 25855 5508 25889
rect 4604 25849 4656 25855
rect 5456 25849 5508 25855
rect 5526 25889 5578 25901
rect 5596 25889 5648 25901
rect 6448 25889 6500 25901
rect 6518 25889 6570 25901
rect 6588 25889 6640 25901
rect 7440 25889 7492 25901
rect 7510 25889 7562 25901
rect 7580 25889 7632 25901
rect 8432 25889 8484 25901
rect 8502 25889 8554 25901
rect 8572 25889 8624 25901
rect 9424 25889 9476 25901
rect 5526 25855 5546 25889
rect 5546 25855 5578 25889
rect 5596 25855 5618 25889
rect 5618 25855 5648 25889
rect 6448 25855 6482 25889
rect 6482 25855 6500 25889
rect 6518 25855 6554 25889
rect 6554 25855 6570 25889
rect 6588 25855 6626 25889
rect 6626 25855 6640 25889
rect 7440 25855 7452 25889
rect 7452 25855 7490 25889
rect 7490 25855 7492 25889
rect 7510 25855 7524 25889
rect 7524 25855 7562 25889
rect 7580 25855 7596 25889
rect 7596 25855 7632 25889
rect 8432 25855 8460 25889
rect 8460 25855 8484 25889
rect 8502 25855 8532 25889
rect 8532 25855 8554 25889
rect 8572 25855 8604 25889
rect 8604 25855 8624 25889
rect 9424 25855 9434 25889
rect 9434 25855 9468 25889
rect 9468 25855 9476 25889
rect 5526 25849 5578 25855
rect 5596 25849 5648 25855
rect 6448 25849 6500 25855
rect 6518 25849 6570 25855
rect 6588 25849 6640 25855
rect 7440 25849 7492 25855
rect 7510 25849 7562 25855
rect 7580 25849 7632 25855
rect 8432 25849 8484 25855
rect 8502 25849 8554 25855
rect 8572 25849 8624 25855
rect 9424 25849 9476 25855
rect 9494 25889 9546 25901
rect 9494 25855 9506 25889
rect 9506 25855 9540 25889
rect 9540 25855 9546 25889
rect 9494 25849 9546 25855
rect 9564 25889 9616 25901
rect 9564 25855 9578 25889
rect 9578 25855 9612 25889
rect 9612 25855 9616 25889
rect 9564 25849 9616 25855
rect 2480 25815 2532 25831
rect 2550 25815 2602 25831
rect 2620 25815 2672 25831
rect 3472 25815 3524 25831
rect 3542 25815 3594 25831
rect 3612 25815 3664 25831
rect 4464 25815 4516 25831
rect 2480 25781 2506 25815
rect 2506 25781 2532 25815
rect 2550 25781 2579 25815
rect 2579 25781 2602 25815
rect 2620 25781 2652 25815
rect 2652 25781 2672 25815
rect 3472 25781 3489 25815
rect 3489 25781 3524 25815
rect 3542 25781 3562 25815
rect 3562 25781 3594 25815
rect 3612 25781 3635 25815
rect 3635 25781 3664 25815
rect 4464 25781 4466 25815
rect 4466 25781 4500 25815
rect 4500 25781 4516 25815
rect 2480 25779 2532 25781
rect 2550 25779 2602 25781
rect 2620 25779 2672 25781
rect 3472 25779 3524 25781
rect 3542 25779 3594 25781
rect 3612 25779 3664 25781
rect 4464 25779 4516 25781
rect 4534 25815 4586 25831
rect 4534 25781 4538 25815
rect 4538 25781 4572 25815
rect 4572 25781 4586 25815
rect 4534 25779 4586 25781
rect 4604 25815 4656 25831
rect 5456 25815 5508 25831
rect 4604 25781 4610 25815
rect 4610 25781 4644 25815
rect 4644 25781 4656 25815
rect 5456 25781 5474 25815
rect 5474 25781 5508 25815
rect 4604 25779 4656 25781
rect 5456 25779 5508 25781
rect 5526 25815 5578 25831
rect 5596 25815 5648 25831
rect 6448 25815 6500 25831
rect 6518 25815 6570 25831
rect 6588 25815 6640 25831
rect 7440 25815 7492 25831
rect 7510 25815 7562 25831
rect 7580 25815 7632 25831
rect 8432 25815 8484 25831
rect 8502 25815 8554 25831
rect 8572 25815 8624 25831
rect 9424 25815 9476 25831
rect 5526 25781 5546 25815
rect 5546 25781 5578 25815
rect 5596 25781 5618 25815
rect 5618 25781 5648 25815
rect 6448 25781 6482 25815
rect 6482 25781 6500 25815
rect 6518 25781 6554 25815
rect 6554 25781 6570 25815
rect 6588 25781 6626 25815
rect 6626 25781 6640 25815
rect 7440 25781 7452 25815
rect 7452 25781 7490 25815
rect 7490 25781 7492 25815
rect 7510 25781 7524 25815
rect 7524 25781 7562 25815
rect 7580 25781 7596 25815
rect 7596 25781 7632 25815
rect 8432 25781 8460 25815
rect 8460 25781 8484 25815
rect 8502 25781 8532 25815
rect 8532 25781 8554 25815
rect 8572 25781 8604 25815
rect 8604 25781 8624 25815
rect 9424 25781 9434 25815
rect 9434 25781 9468 25815
rect 9468 25781 9476 25815
rect 5526 25779 5578 25781
rect 5596 25779 5648 25781
rect 6448 25779 6500 25781
rect 6518 25779 6570 25781
rect 6588 25779 6640 25781
rect 7440 25779 7492 25781
rect 7510 25779 7562 25781
rect 7580 25779 7632 25781
rect 8432 25779 8484 25781
rect 8502 25779 8554 25781
rect 8572 25779 8624 25781
rect 9424 25779 9476 25781
rect 9494 25815 9546 25831
rect 9494 25781 9506 25815
rect 9506 25781 9540 25815
rect 9540 25781 9546 25815
rect 9494 25779 9546 25781
rect 9564 25815 9616 25831
rect 9564 25781 9578 25815
rect 9578 25781 9612 25815
rect 9612 25781 9616 25815
rect 9564 25779 9616 25781
rect 2480 25741 2532 25760
rect 2550 25741 2602 25760
rect 2620 25741 2672 25760
rect 3472 25741 3524 25760
rect 3542 25741 3594 25760
rect 3612 25741 3664 25760
rect 4464 25741 4516 25760
rect 2480 25708 2506 25741
rect 2506 25708 2532 25741
rect 2550 25708 2579 25741
rect 2579 25708 2602 25741
rect 2620 25708 2652 25741
rect 2652 25708 2672 25741
rect 3472 25708 3489 25741
rect 3489 25708 3524 25741
rect 3542 25708 3562 25741
rect 3562 25708 3594 25741
rect 3612 25708 3635 25741
rect 3635 25708 3664 25741
rect 4464 25708 4466 25741
rect 4466 25708 4500 25741
rect 4500 25708 4516 25741
rect 4534 25741 4586 25760
rect 4534 25708 4538 25741
rect 4538 25708 4572 25741
rect 4572 25708 4586 25741
rect 4604 25741 4656 25760
rect 5456 25741 5508 25760
rect 4604 25708 4610 25741
rect 4610 25708 4644 25741
rect 4644 25708 4656 25741
rect 5456 25708 5474 25741
rect 5474 25708 5508 25741
rect 5526 25741 5578 25760
rect 5596 25741 5648 25760
rect 6448 25741 6500 25760
rect 6518 25741 6570 25760
rect 6588 25741 6640 25760
rect 7440 25741 7492 25760
rect 7510 25741 7562 25760
rect 7580 25741 7632 25760
rect 8432 25741 8484 25760
rect 8502 25741 8554 25760
rect 8572 25741 8624 25760
rect 9424 25741 9476 25760
rect 5526 25708 5546 25741
rect 5546 25708 5578 25741
rect 5596 25708 5618 25741
rect 5618 25708 5648 25741
rect 6448 25708 6482 25741
rect 6482 25708 6500 25741
rect 6518 25708 6554 25741
rect 6554 25708 6570 25741
rect 6588 25708 6626 25741
rect 6626 25708 6640 25741
rect 7440 25708 7452 25741
rect 7452 25708 7490 25741
rect 7490 25708 7492 25741
rect 7510 25708 7524 25741
rect 7524 25708 7562 25741
rect 7580 25708 7596 25741
rect 7596 25708 7632 25741
rect 8432 25708 8460 25741
rect 8460 25708 8484 25741
rect 8502 25708 8532 25741
rect 8532 25708 8554 25741
rect 8572 25708 8604 25741
rect 8604 25708 8624 25741
rect 9424 25708 9434 25741
rect 9434 25708 9468 25741
rect 9468 25708 9476 25741
rect 9494 25741 9546 25760
rect 9494 25708 9506 25741
rect 9506 25708 9540 25741
rect 9540 25708 9546 25741
rect 9564 25741 9616 25760
rect 9564 25708 9578 25741
rect 9578 25708 9612 25741
rect 9612 25708 9616 25741
rect 2480 25667 2532 25689
rect 2550 25667 2602 25689
rect 2620 25667 2672 25689
rect 3472 25667 3524 25689
rect 3542 25667 3594 25689
rect 3612 25667 3664 25689
rect 4464 25667 4516 25689
rect 2480 25637 2506 25667
rect 2506 25637 2532 25667
rect 2550 25637 2579 25667
rect 2579 25637 2602 25667
rect 2620 25637 2652 25667
rect 2652 25637 2672 25667
rect 3472 25637 3489 25667
rect 3489 25637 3524 25667
rect 3542 25637 3562 25667
rect 3562 25637 3594 25667
rect 3612 25637 3635 25667
rect 3635 25637 3664 25667
rect 4464 25637 4466 25667
rect 4466 25637 4500 25667
rect 4500 25637 4516 25667
rect 4534 25667 4586 25689
rect 4534 25637 4538 25667
rect 4538 25637 4572 25667
rect 4572 25637 4586 25667
rect 4604 25667 4656 25689
rect 5456 25667 5508 25689
rect 4604 25637 4610 25667
rect 4610 25637 4644 25667
rect 4644 25637 4656 25667
rect 5456 25637 5474 25667
rect 5474 25637 5508 25667
rect 5526 25667 5578 25689
rect 5596 25667 5648 25689
rect 6448 25667 6500 25689
rect 6518 25667 6570 25689
rect 6588 25667 6640 25689
rect 7440 25667 7492 25689
rect 7510 25667 7562 25689
rect 7580 25667 7632 25689
rect 8432 25667 8484 25689
rect 8502 25667 8554 25689
rect 8572 25667 8624 25689
rect 9424 25667 9476 25689
rect 5526 25637 5546 25667
rect 5546 25637 5578 25667
rect 5596 25637 5618 25667
rect 5618 25637 5648 25667
rect 6448 25637 6482 25667
rect 6482 25637 6500 25667
rect 6518 25637 6554 25667
rect 6554 25637 6570 25667
rect 6588 25637 6626 25667
rect 6626 25637 6640 25667
rect 7440 25637 7452 25667
rect 7452 25637 7490 25667
rect 7490 25637 7492 25667
rect 7510 25637 7524 25667
rect 7524 25637 7562 25667
rect 7580 25637 7596 25667
rect 7596 25637 7632 25667
rect 8432 25637 8460 25667
rect 8460 25637 8484 25667
rect 8502 25637 8532 25667
rect 8532 25637 8554 25667
rect 8572 25637 8604 25667
rect 8604 25637 8624 25667
rect 9424 25637 9434 25667
rect 9434 25637 9468 25667
rect 9468 25637 9476 25667
rect 9494 25667 9546 25689
rect 9494 25637 9506 25667
rect 9506 25637 9540 25667
rect 9540 25637 9546 25667
rect 9564 25667 9616 25689
rect 9564 25637 9578 25667
rect 9578 25637 9612 25667
rect 9612 25637 9616 25667
rect 1303 25007 1329 25037
rect 1329 25007 1355 25037
rect 1371 25007 1402 25037
rect 1402 25007 1423 25037
rect 1439 25007 1475 25037
rect 1475 25007 1491 25037
rect 1507 25007 1509 25037
rect 1509 25007 1548 25037
rect 1548 25007 1559 25037
rect 1575 25007 1582 25037
rect 1582 25007 1621 25037
rect 1621 25007 1627 25037
rect 1643 25007 1655 25037
rect 1655 25007 1694 25037
rect 1694 25007 1695 25037
rect 1711 25007 1728 25037
rect 1728 25007 1763 25037
rect 1779 25007 1801 25037
rect 1801 25007 1831 25037
rect 1847 25007 1874 25037
rect 1874 25007 1899 25037
rect 1914 25007 1947 25037
rect 1947 25007 1966 25037
rect 1303 24985 1355 25007
rect 1371 24985 1423 25007
rect 1439 24985 1491 25007
rect 1507 24985 1559 25007
rect 1575 24985 1627 25007
rect 1643 24985 1695 25007
rect 1711 24985 1763 25007
rect 1779 24985 1831 25007
rect 1847 24985 1899 25007
rect 1914 24985 1966 25007
rect 1981 25007 1986 25037
rect 1986 25007 2020 25037
rect 2020 25007 2033 25037
rect 1981 24985 2033 25007
rect 12157 24985 12209 25037
rect 12225 24985 12277 25037
rect 12293 24985 12345 25037
rect 12361 24985 12413 25037
rect 12429 24985 12481 25037
rect 12497 24985 12549 25037
rect 12565 24985 12617 25037
rect 12633 24985 12685 25037
rect 12701 24985 12753 25037
rect 12768 24985 12820 25037
rect 12835 24985 12887 25037
rect 1303 24935 1329 24967
rect 1329 24935 1355 24967
rect 1371 24935 1402 24967
rect 1402 24935 1423 24967
rect 1439 24935 1475 24967
rect 1475 24935 1491 24967
rect 1507 24935 1509 24967
rect 1509 24935 1548 24967
rect 1548 24935 1559 24967
rect 1575 24935 1582 24967
rect 1582 24935 1621 24967
rect 1621 24935 1627 24967
rect 1643 24935 1655 24967
rect 1655 24935 1694 24967
rect 1694 24935 1695 24967
rect 1711 24935 1728 24967
rect 1728 24935 1763 24967
rect 1779 24935 1801 24967
rect 1801 24935 1831 24967
rect 1847 24935 1874 24967
rect 1874 24935 1899 24967
rect 1914 24935 1947 24967
rect 1947 24935 1966 24967
rect 1303 24915 1355 24935
rect 1371 24915 1423 24935
rect 1439 24915 1491 24935
rect 1507 24915 1559 24935
rect 1575 24915 1627 24935
rect 1643 24915 1695 24935
rect 1711 24915 1763 24935
rect 1779 24915 1831 24935
rect 1847 24915 1899 24935
rect 1914 24915 1966 24935
rect 1981 24935 1986 24967
rect 1986 24935 2020 24967
rect 2020 24935 2033 24967
rect 1981 24915 2033 24935
rect 12157 24915 12209 24967
rect 12225 24915 12277 24967
rect 12293 24915 12345 24967
rect 12361 24915 12413 24967
rect 12429 24915 12481 24967
rect 12497 24915 12549 24967
rect 12565 24915 12617 24967
rect 12633 24915 12685 24967
rect 12701 24915 12753 24967
rect 12768 24915 12820 24967
rect 12835 24915 12887 24967
rect 1303 24863 1329 24897
rect 1329 24863 1355 24897
rect 1371 24863 1402 24897
rect 1402 24863 1423 24897
rect 1439 24863 1475 24897
rect 1475 24863 1491 24897
rect 1507 24863 1509 24897
rect 1509 24863 1548 24897
rect 1548 24863 1559 24897
rect 1575 24863 1582 24897
rect 1582 24863 1621 24897
rect 1621 24863 1627 24897
rect 1643 24863 1655 24897
rect 1655 24863 1694 24897
rect 1694 24863 1695 24897
rect 1711 24863 1728 24897
rect 1728 24863 1763 24897
rect 1779 24863 1801 24897
rect 1801 24863 1831 24897
rect 1847 24863 1874 24897
rect 1874 24863 1899 24897
rect 1914 24863 1947 24897
rect 1947 24863 1966 24897
rect 1303 24845 1355 24863
rect 1371 24845 1423 24863
rect 1439 24845 1491 24863
rect 1507 24845 1559 24863
rect 1575 24845 1627 24863
rect 1643 24845 1695 24863
rect 1711 24845 1763 24863
rect 1779 24845 1831 24863
rect 1847 24845 1899 24863
rect 1914 24845 1966 24863
rect 1981 24863 1986 24897
rect 1986 24863 2020 24897
rect 2020 24863 2033 24897
rect 1981 24845 2033 24863
rect 12157 24845 12209 24897
rect 12225 24845 12277 24897
rect 12293 24845 12345 24897
rect 12361 24845 12413 24897
rect 12429 24845 12481 24897
rect 12497 24845 12549 24897
rect 12565 24845 12617 24897
rect 12633 24845 12685 24897
rect 12701 24845 12753 24897
rect 12768 24845 12820 24897
rect 12835 24845 12887 24897
rect 1303 24825 1355 24827
rect 1371 24825 1423 24827
rect 1439 24825 1491 24827
rect 1507 24825 1559 24827
rect 1575 24825 1627 24827
rect 1643 24825 1695 24827
rect 1711 24825 1763 24827
rect 1779 24825 1831 24827
rect 1847 24825 1899 24827
rect 1914 24825 1966 24827
rect 1303 24791 1329 24825
rect 1329 24791 1355 24825
rect 1371 24791 1402 24825
rect 1402 24791 1423 24825
rect 1439 24791 1475 24825
rect 1475 24791 1491 24825
rect 1507 24791 1509 24825
rect 1509 24791 1548 24825
rect 1548 24791 1559 24825
rect 1575 24791 1582 24825
rect 1582 24791 1621 24825
rect 1621 24791 1627 24825
rect 1643 24791 1655 24825
rect 1655 24791 1694 24825
rect 1694 24791 1695 24825
rect 1711 24791 1728 24825
rect 1728 24791 1763 24825
rect 1779 24791 1801 24825
rect 1801 24791 1831 24825
rect 1847 24791 1874 24825
rect 1874 24791 1899 24825
rect 1914 24791 1947 24825
rect 1947 24791 1966 24825
rect 1303 24775 1355 24791
rect 1371 24775 1423 24791
rect 1439 24775 1491 24791
rect 1507 24775 1559 24791
rect 1575 24775 1627 24791
rect 1643 24775 1695 24791
rect 1711 24775 1763 24791
rect 1779 24775 1831 24791
rect 1847 24775 1899 24791
rect 1914 24775 1966 24791
rect 1981 24825 2033 24827
rect 1981 24791 1986 24825
rect 1986 24791 2020 24825
rect 2020 24791 2033 24825
rect 1981 24775 2033 24791
rect 12157 24775 12209 24827
rect 12225 24775 12277 24827
rect 12293 24775 12345 24827
rect 12361 24775 12413 24827
rect 12429 24775 12481 24827
rect 12497 24775 12549 24827
rect 12565 24775 12617 24827
rect 12633 24775 12685 24827
rect 12701 24775 12753 24827
rect 12768 24775 12820 24827
rect 12835 24775 12887 24827
rect 1303 24753 1355 24757
rect 1371 24753 1423 24757
rect 1439 24753 1491 24757
rect 1507 24753 1559 24757
rect 1575 24753 1627 24757
rect 1643 24753 1695 24757
rect 1711 24753 1763 24757
rect 1779 24753 1831 24757
rect 1847 24753 1899 24757
rect 1914 24753 1966 24757
rect 1303 24719 1329 24753
rect 1329 24719 1355 24753
rect 1371 24719 1402 24753
rect 1402 24719 1423 24753
rect 1439 24719 1475 24753
rect 1475 24719 1491 24753
rect 1507 24719 1509 24753
rect 1509 24719 1548 24753
rect 1548 24719 1559 24753
rect 1575 24719 1582 24753
rect 1582 24719 1621 24753
rect 1621 24719 1627 24753
rect 1643 24719 1655 24753
rect 1655 24719 1694 24753
rect 1694 24719 1695 24753
rect 1711 24719 1728 24753
rect 1728 24719 1763 24753
rect 1779 24719 1801 24753
rect 1801 24719 1831 24753
rect 1847 24719 1874 24753
rect 1874 24719 1899 24753
rect 1914 24719 1947 24753
rect 1947 24719 1966 24753
rect 1303 24705 1355 24719
rect 1371 24705 1423 24719
rect 1439 24705 1491 24719
rect 1507 24705 1559 24719
rect 1575 24705 1627 24719
rect 1643 24705 1695 24719
rect 1711 24705 1763 24719
rect 1779 24705 1831 24719
rect 1847 24705 1899 24719
rect 1914 24705 1966 24719
rect 1981 24753 2033 24757
rect 1981 24719 1986 24753
rect 1986 24719 2020 24753
rect 2020 24719 2033 24753
rect 12157 24719 12209 24757
rect 12225 24719 12277 24757
rect 12293 24719 12345 24757
rect 12361 24719 12413 24757
rect 12429 24719 12481 24757
rect 12497 24719 12549 24757
rect 12565 24719 12617 24757
rect 12633 24719 12685 24757
rect 12701 24719 12753 24757
rect 12768 24719 12820 24757
rect 12835 24719 12887 24757
rect 1981 24705 2033 24719
rect 12157 24705 12209 24719
rect 12225 24705 12277 24719
rect 12293 24705 12345 24719
rect 12361 24705 12413 24719
rect 12429 24705 12481 24719
rect 12497 24705 12549 24719
rect 12565 24705 12617 24719
rect 12633 24705 12685 24719
rect 12701 24705 12753 24719
rect 12768 24705 12820 24719
rect 12835 24705 12887 24719
rect 1303 24635 1355 24687
rect 1371 24635 1423 24687
rect 1439 24635 1491 24687
rect 1507 24635 1559 24687
rect 1575 24635 1627 24687
rect 1643 24635 1695 24687
rect 1711 24635 1763 24687
rect 1779 24635 1831 24687
rect 1847 24635 1899 24687
rect 1914 24635 1966 24687
rect 1981 24635 2033 24687
rect 1303 24565 1355 24617
rect 1371 24565 1423 24617
rect 1439 24565 1491 24617
rect 1507 24565 1559 24617
rect 1575 24565 1627 24617
rect 1643 24565 1695 24617
rect 1711 24565 1763 24617
rect 1779 24565 1831 24617
rect 1847 24565 1899 24617
rect 1914 24565 1966 24617
rect 1981 24565 2033 24617
rect 1303 24495 1355 24547
rect 1371 24495 1423 24547
rect 1439 24495 1491 24547
rect 1507 24495 1559 24547
rect 1575 24495 1627 24547
rect 1643 24495 1695 24547
rect 1711 24495 1763 24547
rect 1779 24495 1831 24547
rect 1847 24495 1899 24547
rect 1914 24495 1966 24547
rect 1981 24495 2033 24547
rect 12157 24635 12209 24687
rect 12225 24635 12277 24687
rect 12293 24635 12345 24687
rect 12361 24635 12413 24687
rect 12429 24635 12481 24687
rect 12497 24635 12549 24687
rect 12565 24635 12617 24687
rect 12633 24635 12685 24687
rect 12701 24635 12753 24687
rect 12768 24635 12820 24687
rect 12835 24635 12887 24687
rect 12157 24565 12209 24617
rect 12225 24565 12277 24617
rect 12293 24565 12345 24617
rect 12361 24565 12413 24617
rect 12429 24565 12481 24617
rect 12497 24565 12549 24617
rect 12565 24565 12617 24617
rect 12633 24565 12685 24617
rect 12701 24565 12753 24617
rect 12768 24565 12820 24617
rect 12835 24565 12887 24617
rect 12157 24495 12209 24547
rect 12225 24495 12277 24547
rect 12293 24495 12345 24547
rect 12361 24495 12413 24547
rect 12429 24495 12481 24547
rect 12497 24495 12549 24547
rect 12565 24495 12617 24547
rect 12633 24495 12685 24547
rect 12701 24495 12753 24547
rect 12768 24495 12820 24547
rect 12835 24495 12887 24547
rect 14755 21361 14807 21413
rect 14821 21361 14873 21413
rect 14887 21361 14939 21413
rect 14755 21296 14807 21348
rect 14821 21296 14873 21348
rect 14887 21296 14939 21348
rect 14755 21230 14807 21282
rect 14821 21230 14873 21282
rect 14887 21230 14939 21282
rect 14755 21164 14807 21216
rect 14821 21164 14873 21216
rect 14887 21164 14939 21216
rect 14755 21098 14807 21150
rect 14821 21098 14873 21150
rect 14887 21098 14939 21150
rect 14755 21032 14807 21084
rect 14821 21032 14873 21084
rect 14887 21032 14939 21084
rect 14755 20966 14807 21018
rect 14821 20966 14873 21018
rect 14887 20966 14939 21018
rect 14755 20900 14807 20952
rect 14821 20900 14873 20952
rect 14887 20900 14939 20952
rect 14755 20834 14807 20886
rect 14821 20834 14873 20886
rect 14887 20834 14939 20886
rect 14755 20768 14807 20820
rect 14821 20768 14873 20820
rect 14887 20768 14939 20820
rect 14755 20702 14807 20754
rect 14821 20702 14873 20754
rect 14887 20702 14939 20754
rect 14755 20636 14807 20688
rect 14821 20636 14873 20688
rect 14887 20636 14939 20688
rect 14755 20570 14807 20622
rect 14821 20570 14873 20622
rect 14887 20570 14939 20622
rect 14755 20504 14807 20556
rect 14821 20504 14873 20556
rect 14887 20504 14939 20556
rect 14755 20438 14807 20490
rect 14821 20438 14873 20490
rect 14887 20438 14939 20490
rect 14755 20372 14807 20424
rect 14821 20372 14873 20424
rect 14887 20372 14939 20424
rect 14755 20306 14807 20358
rect 14821 20306 14873 20358
rect 14887 20306 14939 20358
rect 14755 20240 14807 20292
rect 14821 20240 14873 20292
rect 14887 20240 14939 20292
rect 14755 20174 14807 20226
rect 14821 20174 14873 20226
rect 14887 20174 14939 20226
rect 14755 20108 14807 20160
rect 14821 20108 14873 20160
rect 14887 20108 14939 20160
rect 14755 20042 14807 20094
rect 14821 20042 14873 20094
rect 14887 20042 14939 20094
rect 14755 19976 14807 20028
rect 14821 19976 14873 20028
rect 14887 19976 14939 20028
rect 201 19912 253 19964
rect 269 19912 321 19964
rect 337 19912 389 19964
rect 404 19912 456 19964
rect 471 19912 523 19964
rect 538 19912 590 19964
rect 605 19912 657 19964
rect 672 19912 724 19964
rect 739 19912 791 19964
rect 806 19912 858 19964
rect 873 19912 925 19964
rect 940 19912 992 19964
rect 1007 19912 1059 19964
rect 1074 19912 1126 19964
rect 1141 19912 1193 19964
rect 1208 19912 1260 19964
rect 201 19858 253 19896
rect 201 19844 216 19858
rect 216 19844 250 19858
rect 250 19844 253 19858
rect 269 19858 321 19896
rect 337 19858 389 19896
rect 404 19858 456 19896
rect 471 19858 523 19896
rect 538 19858 590 19896
rect 605 19858 657 19896
rect 672 19858 724 19896
rect 739 19858 791 19896
rect 806 19858 858 19896
rect 269 19844 289 19858
rect 289 19844 321 19858
rect 337 19844 362 19858
rect 362 19844 389 19858
rect 404 19844 435 19858
rect 435 19844 456 19858
rect 471 19844 508 19858
rect 508 19844 523 19858
rect 538 19844 542 19858
rect 542 19844 581 19858
rect 581 19844 590 19858
rect 605 19844 615 19858
rect 615 19844 654 19858
rect 654 19844 657 19858
rect 672 19844 688 19858
rect 688 19844 724 19858
rect 739 19844 761 19858
rect 761 19844 791 19858
rect 806 19844 834 19858
rect 834 19844 858 19858
rect 873 19858 925 19896
rect 873 19844 907 19858
rect 907 19844 925 19858
rect 940 19858 992 19896
rect 940 19844 946 19858
rect 946 19844 980 19858
rect 980 19844 992 19858
rect 1007 19858 1059 19896
rect 1007 19844 1019 19858
rect 1019 19844 1053 19858
rect 1053 19844 1059 19858
rect 1074 19858 1126 19896
rect 1074 19844 1092 19858
rect 1092 19844 1126 19858
rect 1141 19858 1193 19896
rect 1208 19858 1260 19896
rect 8200 19912 8252 19964
rect 8268 19912 8320 19964
rect 8336 19912 8388 19964
rect 8403 19912 8455 19964
rect 8470 19912 8522 19964
rect 8537 19912 8589 19964
rect 8604 19912 8656 19964
rect 8671 19912 8723 19964
rect 8738 19912 8790 19964
rect 8805 19912 8857 19964
rect 8872 19912 8924 19964
rect 8939 19912 8991 19964
rect 9006 19912 9058 19964
rect 9073 19912 9125 19964
rect 9140 19912 9192 19964
rect 9207 19912 9259 19964
rect 8200 19858 8252 19896
rect 8268 19858 8320 19896
rect 8336 19858 8388 19896
rect 8403 19858 8455 19896
rect 8470 19858 8522 19896
rect 1141 19844 1165 19858
rect 1165 19844 1193 19858
rect 1208 19844 1238 19858
rect 1238 19844 1260 19858
rect 201 19824 216 19828
rect 216 19824 250 19828
rect 250 19824 253 19828
rect 201 19776 253 19824
rect 269 19824 289 19828
rect 289 19824 321 19828
rect 337 19824 362 19828
rect 362 19824 389 19828
rect 404 19824 435 19828
rect 435 19824 456 19828
rect 471 19824 508 19828
rect 508 19824 523 19828
rect 538 19824 542 19828
rect 542 19824 581 19828
rect 581 19824 590 19828
rect 605 19824 615 19828
rect 615 19824 654 19828
rect 654 19824 657 19828
rect 672 19824 688 19828
rect 688 19824 724 19828
rect 739 19824 761 19828
rect 761 19824 791 19828
rect 806 19824 834 19828
rect 834 19824 858 19828
rect 269 19776 321 19824
rect 337 19776 389 19824
rect 404 19776 456 19824
rect 471 19776 523 19824
rect 538 19776 590 19824
rect 605 19776 657 19824
rect 672 19776 724 19824
rect 739 19776 791 19824
rect 806 19776 858 19824
rect 873 19824 907 19828
rect 907 19824 925 19828
rect 873 19776 925 19824
rect 940 19824 946 19828
rect 946 19824 980 19828
rect 980 19824 992 19828
rect 940 19776 992 19824
rect 1007 19824 1019 19828
rect 1019 19824 1053 19828
rect 1053 19824 1059 19828
rect 1007 19776 1059 19824
rect 1074 19824 1092 19828
rect 1092 19824 1126 19828
rect 1074 19776 1126 19824
rect 1141 19824 1165 19828
rect 1165 19824 1193 19828
rect 1208 19824 1238 19828
rect 1238 19824 1260 19828
rect 8200 19844 8212 19858
rect 8212 19844 8250 19858
rect 8250 19844 8252 19858
rect 8268 19844 8284 19858
rect 8284 19844 8320 19858
rect 8336 19844 8356 19858
rect 8356 19844 8388 19858
rect 8403 19844 8428 19858
rect 8428 19844 8455 19858
rect 8470 19844 8500 19858
rect 8500 19844 8522 19858
rect 8537 19858 8589 19896
rect 8537 19844 8538 19858
rect 8538 19844 8572 19858
rect 8572 19844 8589 19858
rect 8604 19858 8656 19896
rect 8604 19844 8610 19858
rect 8610 19844 8644 19858
rect 8644 19844 8656 19858
rect 8671 19858 8723 19896
rect 8671 19844 8682 19858
rect 8682 19844 8716 19858
rect 8716 19844 8723 19858
rect 8738 19858 8790 19896
rect 8738 19844 8754 19858
rect 8754 19844 8788 19858
rect 8788 19844 8790 19858
rect 8805 19858 8857 19896
rect 8872 19858 8924 19896
rect 8939 19858 8991 19896
rect 9006 19858 9058 19896
rect 9073 19858 9125 19896
rect 9140 19858 9192 19896
rect 9207 19858 9259 19896
rect 14755 19910 14807 19962
rect 14821 19910 14873 19962
rect 14887 19910 14939 19962
rect 14755 19858 14807 19896
rect 14821 19858 14873 19896
rect 14887 19858 14939 19896
rect 8805 19844 8826 19858
rect 8826 19844 8857 19858
rect 8872 19844 8898 19858
rect 8898 19844 8924 19858
rect 8939 19844 8970 19858
rect 8970 19844 8991 19858
rect 9006 19844 9042 19858
rect 9042 19844 9058 19858
rect 9073 19844 9076 19858
rect 9076 19844 9114 19858
rect 9114 19844 9125 19858
rect 9140 19844 9148 19858
rect 9148 19844 9186 19858
rect 9186 19844 9192 19858
rect 9207 19844 9220 19858
rect 9220 19844 9258 19858
rect 9258 19844 9259 19858
rect 8200 19824 8212 19828
rect 8212 19824 8250 19828
rect 8250 19824 8252 19828
rect 8268 19824 8284 19828
rect 8284 19824 8320 19828
rect 8336 19824 8356 19828
rect 8356 19824 8388 19828
rect 8403 19824 8428 19828
rect 8428 19824 8455 19828
rect 8470 19824 8500 19828
rect 8500 19824 8522 19828
rect 1141 19776 1193 19824
rect 1208 19776 1260 19824
rect 8200 19776 8252 19824
rect 8268 19776 8320 19824
rect 8336 19776 8388 19824
rect 8403 19776 8455 19824
rect 8470 19776 8522 19824
rect 8537 19824 8538 19828
rect 8538 19824 8572 19828
rect 8572 19824 8589 19828
rect 8537 19776 8589 19824
rect 8604 19824 8610 19828
rect 8610 19824 8644 19828
rect 8644 19824 8656 19828
rect 8604 19776 8656 19824
rect 8671 19824 8682 19828
rect 8682 19824 8716 19828
rect 8716 19824 8723 19828
rect 8671 19776 8723 19824
rect 8738 19824 8754 19828
rect 8754 19824 8788 19828
rect 8788 19824 8790 19828
rect 8738 19776 8790 19824
rect 8805 19824 8826 19828
rect 8826 19824 8857 19828
rect 8872 19824 8898 19828
rect 8898 19824 8924 19828
rect 8939 19824 8970 19828
rect 8970 19824 8991 19828
rect 9006 19824 9042 19828
rect 9042 19824 9058 19828
rect 9073 19824 9076 19828
rect 9076 19824 9114 19828
rect 9114 19824 9125 19828
rect 9140 19824 9148 19828
rect 9148 19824 9186 19828
rect 9186 19824 9192 19828
rect 9207 19824 9220 19828
rect 9220 19824 9258 19828
rect 9258 19824 9259 19828
rect 14755 19844 14764 19858
rect 14764 19844 14802 19858
rect 14802 19844 14807 19858
rect 14821 19844 14836 19858
rect 14836 19844 14873 19858
rect 14887 19844 14908 19858
rect 14908 19844 14939 19858
rect 14755 19824 14764 19830
rect 14764 19824 14802 19830
rect 14802 19824 14807 19830
rect 14821 19824 14836 19830
rect 14836 19824 14873 19830
rect 14887 19824 14908 19830
rect 14908 19824 14939 19830
rect 8805 19776 8857 19824
rect 8872 19776 8924 19824
rect 8939 19776 8991 19824
rect 9006 19776 9058 19824
rect 9073 19776 9125 19824
rect 9140 19776 9192 19824
rect 9207 19776 9259 19824
rect 14755 19778 14807 19824
rect 14821 19778 14873 19824
rect 14887 19778 14939 19824
rect 201 19738 216 19760
rect 216 19738 250 19760
rect 250 19738 253 19760
rect 201 19708 253 19738
rect 269 19738 289 19760
rect 289 19738 321 19760
rect 337 19738 362 19760
rect 362 19738 389 19760
rect 404 19738 435 19760
rect 435 19738 456 19760
rect 471 19738 508 19760
rect 508 19738 523 19760
rect 538 19738 542 19760
rect 542 19738 581 19760
rect 581 19738 590 19760
rect 605 19738 615 19760
rect 615 19738 654 19760
rect 654 19738 657 19760
rect 672 19738 688 19760
rect 688 19738 724 19760
rect 739 19738 761 19760
rect 761 19738 791 19760
rect 806 19738 834 19760
rect 834 19738 858 19760
rect 269 19708 321 19738
rect 337 19708 389 19738
rect 404 19708 456 19738
rect 471 19708 523 19738
rect 538 19708 590 19738
rect 605 19708 657 19738
rect 672 19708 724 19738
rect 739 19708 791 19738
rect 806 19708 858 19738
rect 873 19738 907 19760
rect 907 19738 925 19760
rect 873 19708 925 19738
rect 940 19738 946 19760
rect 946 19738 980 19760
rect 980 19738 992 19760
rect 940 19708 992 19738
rect 1007 19738 1019 19760
rect 1019 19738 1053 19760
rect 1053 19738 1059 19760
rect 1007 19708 1059 19738
rect 1074 19738 1092 19760
rect 1092 19738 1126 19760
rect 1074 19708 1126 19738
rect 1141 19738 1165 19760
rect 1165 19738 1193 19760
rect 1208 19738 1238 19760
rect 1238 19738 1260 19760
rect 8200 19738 8212 19760
rect 8212 19738 8250 19760
rect 8250 19738 8252 19760
rect 8268 19738 8284 19760
rect 8284 19738 8320 19760
rect 8336 19738 8356 19760
rect 8356 19738 8388 19760
rect 8403 19738 8428 19760
rect 8428 19738 8455 19760
rect 8470 19738 8500 19760
rect 8500 19738 8522 19760
rect 1141 19708 1193 19738
rect 1208 19708 1260 19738
rect 8200 19708 8252 19738
rect 8268 19708 8320 19738
rect 8336 19708 8388 19738
rect 8403 19708 8455 19738
rect 8470 19708 8522 19738
rect 8537 19738 8538 19760
rect 8538 19738 8572 19760
rect 8572 19738 8589 19760
rect 8537 19708 8589 19738
rect 8604 19738 8610 19760
rect 8610 19738 8644 19760
rect 8644 19738 8656 19760
rect 8604 19708 8656 19738
rect 8671 19738 8682 19760
rect 8682 19738 8716 19760
rect 8716 19738 8723 19760
rect 8671 19708 8723 19738
rect 8738 19738 8754 19760
rect 8754 19738 8788 19760
rect 8788 19738 8790 19760
rect 8738 19708 8790 19738
rect 8805 19738 8826 19760
rect 8826 19738 8857 19760
rect 8872 19738 8898 19760
rect 8898 19738 8924 19760
rect 8939 19738 8970 19760
rect 8970 19738 8991 19760
rect 9006 19738 9042 19760
rect 9042 19738 9058 19760
rect 9073 19738 9076 19760
rect 9076 19738 9114 19760
rect 9114 19738 9125 19760
rect 9140 19738 9148 19760
rect 9148 19738 9186 19760
rect 9186 19738 9192 19760
rect 9207 19738 9220 19760
rect 9220 19738 9258 19760
rect 9258 19738 9259 19760
rect 14755 19738 14764 19764
rect 14764 19738 14802 19764
rect 14802 19738 14807 19764
rect 14821 19738 14836 19764
rect 14836 19738 14873 19764
rect 14887 19738 14908 19764
rect 14908 19738 14939 19764
rect 8805 19708 8857 19738
rect 8872 19708 8924 19738
rect 8939 19708 8991 19738
rect 9006 19708 9058 19738
rect 9073 19708 9125 19738
rect 9140 19708 9192 19738
rect 9207 19708 9259 19738
rect 14755 19712 14807 19738
rect 14821 19712 14873 19738
rect 14887 19712 14939 19738
rect 201 19686 253 19692
rect 201 19652 216 19686
rect 216 19652 250 19686
rect 250 19652 253 19686
rect 201 19640 253 19652
rect 269 19686 321 19692
rect 337 19686 389 19692
rect 404 19686 456 19692
rect 471 19686 523 19692
rect 538 19686 590 19692
rect 605 19686 657 19692
rect 672 19686 724 19692
rect 739 19686 791 19692
rect 806 19686 858 19692
rect 269 19652 289 19686
rect 289 19652 321 19686
rect 337 19652 362 19686
rect 362 19652 389 19686
rect 404 19652 435 19686
rect 435 19652 456 19686
rect 471 19652 508 19686
rect 508 19652 523 19686
rect 538 19652 542 19686
rect 542 19652 581 19686
rect 581 19652 590 19686
rect 605 19652 615 19686
rect 615 19652 654 19686
rect 654 19652 657 19686
rect 672 19652 688 19686
rect 688 19652 724 19686
rect 739 19652 761 19686
rect 761 19652 791 19686
rect 806 19652 834 19686
rect 834 19652 858 19686
rect 269 19640 321 19652
rect 337 19640 389 19652
rect 404 19640 456 19652
rect 471 19640 523 19652
rect 538 19640 590 19652
rect 605 19640 657 19652
rect 672 19640 724 19652
rect 739 19640 791 19652
rect 806 19640 858 19652
rect 873 19686 925 19692
rect 873 19652 907 19686
rect 907 19652 925 19686
rect 873 19640 925 19652
rect 940 19686 992 19692
rect 940 19652 946 19686
rect 946 19652 980 19686
rect 980 19652 992 19686
rect 940 19640 992 19652
rect 1007 19686 1059 19692
rect 1007 19652 1019 19686
rect 1019 19652 1053 19686
rect 1053 19652 1059 19686
rect 1007 19640 1059 19652
rect 1074 19686 1126 19692
rect 1074 19652 1092 19686
rect 1092 19652 1126 19686
rect 1074 19640 1126 19652
rect 1141 19686 1193 19692
rect 1208 19686 1260 19692
rect 8200 19686 8252 19692
rect 8268 19686 8320 19692
rect 8336 19686 8388 19692
rect 8403 19686 8455 19692
rect 8470 19686 8522 19692
rect 1141 19652 1165 19686
rect 1165 19652 1193 19686
rect 1208 19652 1238 19686
rect 1238 19652 1260 19686
rect 8200 19652 8212 19686
rect 8212 19652 8250 19686
rect 8250 19652 8252 19686
rect 8268 19652 8284 19686
rect 8284 19652 8320 19686
rect 8336 19652 8356 19686
rect 8356 19652 8388 19686
rect 8403 19652 8428 19686
rect 8428 19652 8455 19686
rect 8470 19652 8500 19686
rect 8500 19652 8522 19686
rect 1141 19640 1193 19652
rect 1208 19640 1260 19652
rect 8200 19640 8252 19652
rect 8268 19640 8320 19652
rect 8336 19640 8388 19652
rect 8403 19640 8455 19652
rect 8470 19640 8522 19652
rect 8537 19686 8589 19692
rect 8537 19652 8538 19686
rect 8538 19652 8572 19686
rect 8572 19652 8589 19686
rect 8537 19640 8589 19652
rect 8604 19686 8656 19692
rect 8604 19652 8610 19686
rect 8610 19652 8644 19686
rect 8644 19652 8656 19686
rect 8604 19640 8656 19652
rect 8671 19686 8723 19692
rect 8671 19652 8682 19686
rect 8682 19652 8716 19686
rect 8716 19652 8723 19686
rect 8671 19640 8723 19652
rect 8738 19686 8790 19692
rect 8738 19652 8754 19686
rect 8754 19652 8788 19686
rect 8788 19652 8790 19686
rect 8738 19640 8790 19652
rect 8805 19686 8857 19692
rect 8872 19686 8924 19692
rect 8939 19686 8991 19692
rect 9006 19686 9058 19692
rect 9073 19686 9125 19692
rect 9140 19686 9192 19692
rect 9207 19686 9259 19692
rect 14755 19686 14807 19698
rect 14821 19686 14873 19698
rect 14887 19686 14939 19698
rect 8805 19652 8826 19686
rect 8826 19652 8857 19686
rect 8872 19652 8898 19686
rect 8898 19652 8924 19686
rect 8939 19652 8970 19686
rect 8970 19652 8991 19686
rect 9006 19652 9042 19686
rect 9042 19652 9058 19686
rect 9073 19652 9076 19686
rect 9076 19652 9114 19686
rect 9114 19652 9125 19686
rect 9140 19652 9148 19686
rect 9148 19652 9186 19686
rect 9186 19652 9192 19686
rect 9207 19652 9220 19686
rect 9220 19652 9258 19686
rect 9258 19652 9259 19686
rect 14755 19652 14764 19686
rect 14764 19652 14802 19686
rect 14802 19652 14807 19686
rect 14821 19652 14836 19686
rect 14836 19652 14873 19686
rect 14887 19652 14908 19686
rect 14908 19652 14939 19686
rect 8805 19640 8857 19652
rect 8872 19640 8924 19652
rect 8939 19640 8991 19652
rect 9006 19640 9058 19652
rect 9073 19640 9125 19652
rect 9140 19640 9192 19652
rect 9207 19640 9259 19652
rect 14755 19646 14807 19652
rect 14821 19646 14873 19652
rect 14887 19646 14939 19652
rect 201 19600 253 19624
rect 201 19572 216 19600
rect 216 19572 250 19600
rect 250 19572 253 19600
rect 269 19600 321 19624
rect 337 19600 389 19624
rect 404 19600 456 19624
rect 471 19600 523 19624
rect 538 19600 590 19624
rect 605 19600 657 19624
rect 672 19600 724 19624
rect 739 19600 791 19624
rect 806 19600 858 19624
rect 269 19572 289 19600
rect 289 19572 321 19600
rect 337 19572 362 19600
rect 362 19572 389 19600
rect 404 19572 435 19600
rect 435 19572 456 19600
rect 471 19572 508 19600
rect 508 19572 523 19600
rect 538 19572 542 19600
rect 542 19572 581 19600
rect 581 19572 590 19600
rect 605 19572 615 19600
rect 615 19572 654 19600
rect 654 19572 657 19600
rect 672 19572 688 19600
rect 688 19572 724 19600
rect 739 19572 761 19600
rect 761 19572 791 19600
rect 806 19572 834 19600
rect 834 19572 858 19600
rect 873 19600 925 19624
rect 873 19572 907 19600
rect 907 19572 925 19600
rect 940 19600 992 19624
rect 940 19572 946 19600
rect 946 19572 980 19600
rect 980 19572 992 19600
rect 1007 19600 1059 19624
rect 1007 19572 1019 19600
rect 1019 19572 1053 19600
rect 1053 19572 1059 19600
rect 1074 19600 1126 19624
rect 1074 19572 1092 19600
rect 1092 19572 1126 19600
rect 1141 19600 1193 19624
rect 1208 19600 1260 19624
rect 8200 19600 8252 19624
rect 8268 19600 8320 19624
rect 8336 19600 8388 19624
rect 8403 19600 8455 19624
rect 8470 19600 8522 19624
rect 1141 19572 1165 19600
rect 1165 19572 1193 19600
rect 1208 19572 1238 19600
rect 1238 19572 1260 19600
rect 8200 19572 8212 19600
rect 8212 19572 8250 19600
rect 8250 19572 8252 19600
rect 8268 19572 8284 19600
rect 8284 19572 8320 19600
rect 8336 19572 8356 19600
rect 8356 19572 8388 19600
rect 8403 19572 8428 19600
rect 8428 19572 8455 19600
rect 8470 19572 8500 19600
rect 8500 19572 8522 19600
rect 8537 19600 8589 19624
rect 8537 19572 8538 19600
rect 8538 19572 8572 19600
rect 8572 19572 8589 19600
rect 8604 19600 8656 19624
rect 8604 19572 8610 19600
rect 8610 19572 8644 19600
rect 8644 19572 8656 19600
rect 8671 19600 8723 19624
rect 8671 19572 8682 19600
rect 8682 19572 8716 19600
rect 8716 19572 8723 19600
rect 8738 19600 8790 19624
rect 8738 19572 8754 19600
rect 8754 19572 8788 19600
rect 8788 19572 8790 19600
rect 8805 19600 8857 19624
rect 8872 19600 8924 19624
rect 8939 19600 8991 19624
rect 9006 19600 9058 19624
rect 9073 19600 9125 19624
rect 9140 19600 9192 19624
rect 9207 19600 9259 19624
rect 14755 19600 14807 19632
rect 14821 19600 14873 19632
rect 14887 19600 14939 19632
rect 8805 19572 8826 19600
rect 8826 19572 8857 19600
rect 8872 19572 8898 19600
rect 8898 19572 8924 19600
rect 8939 19572 8970 19600
rect 8970 19572 8991 19600
rect 9006 19572 9042 19600
rect 9042 19572 9058 19600
rect 9073 19572 9076 19600
rect 9076 19572 9114 19600
rect 9114 19572 9125 19600
rect 9140 19572 9148 19600
rect 9148 19572 9186 19600
rect 9186 19572 9192 19600
rect 9207 19572 9220 19600
rect 9220 19572 9258 19600
rect 9258 19572 9259 19600
rect 14755 19580 14764 19600
rect 14764 19580 14802 19600
rect 14802 19580 14807 19600
rect 14821 19580 14836 19600
rect 14836 19580 14873 19600
rect 14887 19580 14908 19600
rect 14908 19580 14939 19600
rect 12616 18765 12668 18817
rect 12682 18765 12734 18817
rect 12616 18685 12668 18737
rect 12682 18685 12734 18737
rect 201 18382 253 18387
rect 201 18348 209 18382
rect 209 18348 243 18382
rect 243 18348 253 18382
rect 201 18335 253 18348
rect 269 18382 321 18387
rect 269 18348 282 18382
rect 282 18348 316 18382
rect 316 18348 321 18382
rect 269 18335 321 18348
rect 337 18382 389 18387
rect 337 18348 355 18382
rect 355 18348 389 18382
rect 337 18335 389 18348
rect 404 18382 456 18387
rect 471 18382 523 18387
rect 538 18382 590 18387
rect 605 18382 657 18387
rect 672 18382 724 18387
rect 739 18382 791 18387
rect 806 18382 858 18387
rect 873 18382 925 18387
rect 940 18382 992 18387
rect 404 18348 428 18382
rect 428 18348 456 18382
rect 471 18348 501 18382
rect 501 18348 523 18382
rect 538 18348 574 18382
rect 574 18348 590 18382
rect 605 18348 608 18382
rect 608 18348 647 18382
rect 647 18348 657 18382
rect 672 18348 681 18382
rect 681 18348 720 18382
rect 720 18348 724 18382
rect 739 18348 754 18382
rect 754 18348 791 18382
rect 806 18348 827 18382
rect 827 18348 858 18382
rect 873 18348 900 18382
rect 900 18348 925 18382
rect 940 18348 973 18382
rect 973 18348 992 18382
rect 404 18335 456 18348
rect 471 18335 523 18348
rect 538 18335 590 18348
rect 605 18335 657 18348
rect 672 18335 724 18348
rect 739 18335 791 18348
rect 806 18335 858 18348
rect 873 18335 925 18348
rect 940 18335 992 18348
rect 1007 18382 1059 18387
rect 1007 18348 1012 18382
rect 1012 18348 1046 18382
rect 1046 18348 1059 18382
rect 1007 18335 1059 18348
rect 1074 18382 1126 18387
rect 1074 18348 1085 18382
rect 1085 18348 1119 18382
rect 1119 18348 1126 18382
rect 1074 18335 1126 18348
rect 1141 18382 1193 18387
rect 1141 18348 1158 18382
rect 1158 18348 1192 18382
rect 1192 18348 1193 18382
rect 1141 18335 1193 18348
rect 1208 18382 1260 18387
rect 1208 18348 1231 18382
rect 1231 18348 1260 18382
rect 1208 18335 1260 18348
rect 201 18306 253 18323
rect 201 18272 209 18306
rect 209 18272 243 18306
rect 243 18272 253 18306
rect 201 18271 253 18272
rect 269 18306 321 18323
rect 269 18272 282 18306
rect 282 18272 316 18306
rect 316 18272 321 18306
rect 269 18271 321 18272
rect 337 18306 389 18323
rect 337 18272 355 18306
rect 355 18272 389 18306
rect 337 18271 389 18272
rect 404 18306 456 18323
rect 471 18306 523 18323
rect 538 18306 590 18323
rect 605 18306 657 18323
rect 672 18306 724 18323
rect 739 18306 791 18323
rect 806 18306 858 18323
rect 873 18306 925 18323
rect 940 18306 992 18323
rect 404 18272 428 18306
rect 428 18272 456 18306
rect 471 18272 501 18306
rect 501 18272 523 18306
rect 538 18272 574 18306
rect 574 18272 590 18306
rect 605 18272 608 18306
rect 608 18272 647 18306
rect 647 18272 657 18306
rect 672 18272 681 18306
rect 681 18272 720 18306
rect 720 18272 724 18306
rect 739 18272 754 18306
rect 754 18272 791 18306
rect 806 18272 827 18306
rect 827 18272 858 18306
rect 873 18272 900 18306
rect 900 18272 925 18306
rect 940 18272 973 18306
rect 973 18272 992 18306
rect 404 18271 456 18272
rect 471 18271 523 18272
rect 538 18271 590 18272
rect 605 18271 657 18272
rect 672 18271 724 18272
rect 739 18271 791 18272
rect 806 18271 858 18272
rect 873 18271 925 18272
rect 940 18271 992 18272
rect 1007 18306 1059 18323
rect 1007 18272 1012 18306
rect 1012 18272 1046 18306
rect 1046 18272 1059 18306
rect 1007 18271 1059 18272
rect 1074 18306 1126 18323
rect 1074 18272 1085 18306
rect 1085 18272 1119 18306
rect 1119 18272 1126 18306
rect 1074 18271 1126 18272
rect 1141 18306 1193 18323
rect 1141 18272 1158 18306
rect 1158 18272 1192 18306
rect 1192 18272 1193 18306
rect 1141 18271 1193 18272
rect 1208 18306 1260 18323
rect 1208 18272 1231 18306
rect 1231 18272 1260 18306
rect 1208 18271 1260 18272
rect 201 18230 253 18259
rect 201 18207 209 18230
rect 209 18207 243 18230
rect 243 18207 253 18230
rect 269 18230 321 18259
rect 269 18207 282 18230
rect 282 18207 316 18230
rect 316 18207 321 18230
rect 337 18230 389 18259
rect 337 18207 355 18230
rect 355 18207 389 18230
rect 404 18230 456 18259
rect 471 18230 523 18259
rect 538 18230 590 18259
rect 605 18230 657 18259
rect 672 18230 724 18259
rect 739 18230 791 18259
rect 806 18230 858 18259
rect 873 18230 925 18259
rect 940 18230 992 18259
rect 404 18207 428 18230
rect 428 18207 456 18230
rect 471 18207 501 18230
rect 501 18207 523 18230
rect 538 18207 574 18230
rect 574 18207 590 18230
rect 605 18207 608 18230
rect 608 18207 647 18230
rect 647 18207 657 18230
rect 672 18207 681 18230
rect 681 18207 720 18230
rect 720 18207 724 18230
rect 739 18207 754 18230
rect 754 18207 791 18230
rect 806 18207 827 18230
rect 827 18207 858 18230
rect 873 18207 900 18230
rect 900 18207 925 18230
rect 940 18207 973 18230
rect 973 18207 992 18230
rect 1007 18230 1059 18259
rect 1007 18207 1012 18230
rect 1012 18207 1046 18230
rect 1046 18207 1059 18230
rect 1074 18230 1126 18259
rect 1074 18207 1085 18230
rect 1085 18207 1119 18230
rect 1119 18207 1126 18230
rect 1141 18230 1193 18259
rect 1141 18207 1158 18230
rect 1158 18207 1192 18230
rect 1192 18207 1193 18230
rect 1208 18230 1260 18259
rect 1208 18207 1231 18230
rect 1231 18207 1260 18230
rect 201 18154 253 18195
rect 201 18143 209 18154
rect 209 18143 243 18154
rect 243 18143 253 18154
rect 269 18154 321 18195
rect 269 18143 282 18154
rect 282 18143 316 18154
rect 316 18143 321 18154
rect 337 18154 389 18195
rect 337 18143 355 18154
rect 355 18143 389 18154
rect 404 18154 456 18195
rect 471 18154 523 18195
rect 538 18154 590 18195
rect 605 18154 657 18195
rect 672 18154 724 18195
rect 739 18154 791 18195
rect 806 18154 858 18195
rect 873 18154 925 18195
rect 940 18154 992 18195
rect 404 18143 428 18154
rect 428 18143 456 18154
rect 471 18143 501 18154
rect 501 18143 523 18154
rect 538 18143 574 18154
rect 574 18143 590 18154
rect 605 18143 608 18154
rect 608 18143 647 18154
rect 647 18143 657 18154
rect 672 18143 681 18154
rect 681 18143 720 18154
rect 720 18143 724 18154
rect 739 18143 754 18154
rect 754 18143 791 18154
rect 806 18143 827 18154
rect 827 18143 858 18154
rect 873 18143 900 18154
rect 900 18143 925 18154
rect 940 18143 973 18154
rect 973 18143 992 18154
rect 1007 18154 1059 18195
rect 1007 18143 1012 18154
rect 1012 18143 1046 18154
rect 1046 18143 1059 18154
rect 1074 18154 1126 18195
rect 1074 18143 1085 18154
rect 1085 18143 1119 18154
rect 1119 18143 1126 18154
rect 1141 18154 1193 18195
rect 1141 18143 1158 18154
rect 1158 18143 1192 18154
rect 1192 18143 1193 18154
rect 1208 18154 1260 18195
rect 1208 18143 1231 18154
rect 1231 18143 1260 18154
rect 201 18120 209 18131
rect 209 18120 243 18131
rect 243 18120 253 18131
rect 201 18079 253 18120
rect 269 18120 282 18131
rect 282 18120 316 18131
rect 316 18120 321 18131
rect 269 18079 321 18120
rect 337 18120 355 18131
rect 355 18120 389 18131
rect 337 18079 389 18120
rect 404 18120 428 18131
rect 428 18120 456 18131
rect 471 18120 501 18131
rect 501 18120 523 18131
rect 538 18120 574 18131
rect 574 18120 590 18131
rect 605 18120 608 18131
rect 608 18120 647 18131
rect 647 18120 657 18131
rect 672 18120 681 18131
rect 681 18120 720 18131
rect 720 18120 724 18131
rect 739 18120 754 18131
rect 754 18120 791 18131
rect 806 18120 827 18131
rect 827 18120 858 18131
rect 873 18120 900 18131
rect 900 18120 925 18131
rect 940 18120 973 18131
rect 973 18120 992 18131
rect 404 18079 456 18120
rect 471 18079 523 18120
rect 538 18079 590 18120
rect 605 18079 657 18120
rect 672 18079 724 18120
rect 739 18079 791 18120
rect 806 18079 858 18120
rect 873 18079 925 18120
rect 940 18079 992 18120
rect 1007 18120 1012 18131
rect 1012 18120 1046 18131
rect 1046 18120 1059 18131
rect 1007 18079 1059 18120
rect 1074 18120 1085 18131
rect 1085 18120 1119 18131
rect 1119 18120 1126 18131
rect 1074 18079 1126 18120
rect 1141 18120 1158 18131
rect 1158 18120 1192 18131
rect 1192 18120 1193 18131
rect 1141 18079 1193 18120
rect 1208 18120 1231 18131
rect 1231 18120 1260 18131
rect 1208 18079 1260 18120
rect 201 18044 209 18067
rect 209 18044 243 18067
rect 243 18044 253 18067
rect 201 18015 253 18044
rect 269 18044 282 18067
rect 282 18044 316 18067
rect 316 18044 321 18067
rect 269 18015 321 18044
rect 337 18044 355 18067
rect 355 18044 389 18067
rect 337 18015 389 18044
rect 404 18044 428 18067
rect 428 18044 456 18067
rect 471 18044 501 18067
rect 501 18044 523 18067
rect 538 18044 574 18067
rect 574 18044 590 18067
rect 605 18044 608 18067
rect 608 18044 647 18067
rect 647 18044 657 18067
rect 672 18044 681 18067
rect 681 18044 720 18067
rect 720 18044 724 18067
rect 739 18044 754 18067
rect 754 18044 791 18067
rect 806 18044 827 18067
rect 827 18044 858 18067
rect 873 18044 900 18067
rect 900 18044 925 18067
rect 940 18044 973 18067
rect 973 18044 992 18067
rect 404 18015 456 18044
rect 471 18015 523 18044
rect 538 18015 590 18044
rect 605 18015 657 18044
rect 672 18015 724 18044
rect 739 18015 791 18044
rect 806 18015 858 18044
rect 873 18015 925 18044
rect 940 18015 992 18044
rect 1007 18044 1012 18067
rect 1012 18044 1046 18067
rect 1046 18044 1059 18067
rect 1007 18015 1059 18044
rect 1074 18044 1085 18067
rect 1085 18044 1119 18067
rect 1119 18044 1126 18067
rect 1074 18015 1126 18044
rect 1141 18044 1158 18067
rect 1158 18044 1192 18067
rect 1192 18044 1193 18067
rect 1141 18015 1193 18044
rect 1208 18044 1231 18067
rect 1231 18044 1260 18067
rect 1208 18015 1260 18044
rect 201 18002 253 18003
rect 201 17968 209 18002
rect 209 17968 243 18002
rect 243 17968 253 18002
rect 201 17951 253 17968
rect 269 18002 321 18003
rect 269 17968 282 18002
rect 282 17968 316 18002
rect 316 17968 321 18002
rect 269 17951 321 17968
rect 337 18002 389 18003
rect 337 17968 355 18002
rect 355 17968 389 18002
rect 337 17951 389 17968
rect 404 18002 456 18003
rect 471 18002 523 18003
rect 538 18002 590 18003
rect 605 18002 657 18003
rect 672 18002 724 18003
rect 739 18002 791 18003
rect 806 18002 858 18003
rect 873 18002 925 18003
rect 940 18002 992 18003
rect 404 17968 428 18002
rect 428 17968 456 18002
rect 471 17968 501 18002
rect 501 17968 523 18002
rect 538 17968 574 18002
rect 574 17968 590 18002
rect 605 17968 608 18002
rect 608 17968 647 18002
rect 647 17968 657 18002
rect 672 17968 681 18002
rect 681 17968 720 18002
rect 720 17968 724 18002
rect 739 17968 754 18002
rect 754 17968 791 18002
rect 806 17968 827 18002
rect 827 17968 858 18002
rect 873 17968 900 18002
rect 900 17968 925 18002
rect 940 17968 973 18002
rect 973 17968 992 18002
rect 404 17951 456 17968
rect 471 17951 523 17968
rect 538 17951 590 17968
rect 605 17951 657 17968
rect 672 17951 724 17968
rect 739 17951 791 17968
rect 806 17951 858 17968
rect 873 17951 925 17968
rect 940 17951 992 17968
rect 1007 18002 1059 18003
rect 1007 17968 1012 18002
rect 1012 17968 1046 18002
rect 1046 17968 1059 18002
rect 1007 17951 1059 17968
rect 1074 18002 1126 18003
rect 1074 17968 1085 18002
rect 1085 17968 1119 18002
rect 1119 17968 1126 18002
rect 1074 17951 1126 17968
rect 1141 18002 1193 18003
rect 1141 17968 1158 18002
rect 1158 17968 1192 18002
rect 1192 17968 1193 18002
rect 1141 17951 1193 17968
rect 1208 18002 1260 18003
rect 1208 17968 1231 18002
rect 1231 17968 1260 18002
rect 1208 17951 1260 17968
rect 201 17926 253 17939
rect 201 17892 209 17926
rect 209 17892 243 17926
rect 243 17892 253 17926
rect 201 17887 253 17892
rect 269 17926 321 17939
rect 269 17892 282 17926
rect 282 17892 316 17926
rect 316 17892 321 17926
rect 269 17887 321 17892
rect 337 17926 389 17939
rect 337 17892 355 17926
rect 355 17892 389 17926
rect 337 17887 389 17892
rect 404 17926 456 17939
rect 471 17926 523 17939
rect 538 17926 590 17939
rect 605 17926 657 17939
rect 672 17926 724 17939
rect 739 17926 791 17939
rect 806 17926 858 17939
rect 873 17926 925 17939
rect 940 17926 992 17939
rect 404 17892 428 17926
rect 428 17892 456 17926
rect 471 17892 501 17926
rect 501 17892 523 17926
rect 538 17892 574 17926
rect 574 17892 590 17926
rect 605 17892 608 17926
rect 608 17892 647 17926
rect 647 17892 657 17926
rect 672 17892 681 17926
rect 681 17892 720 17926
rect 720 17892 724 17926
rect 739 17892 754 17926
rect 754 17892 791 17926
rect 806 17892 827 17926
rect 827 17892 858 17926
rect 873 17892 900 17926
rect 900 17892 925 17926
rect 940 17892 973 17926
rect 973 17892 992 17926
rect 404 17887 456 17892
rect 471 17887 523 17892
rect 538 17887 590 17892
rect 605 17887 657 17892
rect 672 17887 724 17892
rect 739 17887 791 17892
rect 806 17887 858 17892
rect 873 17887 925 17892
rect 940 17887 992 17892
rect 1007 17926 1059 17939
rect 1007 17892 1012 17926
rect 1012 17892 1046 17926
rect 1046 17892 1059 17926
rect 1007 17887 1059 17892
rect 1074 17926 1126 17939
rect 1074 17892 1085 17926
rect 1085 17892 1119 17926
rect 1119 17892 1126 17926
rect 1074 17887 1126 17892
rect 1141 17926 1193 17939
rect 1141 17892 1158 17926
rect 1158 17892 1192 17926
rect 1192 17892 1193 17926
rect 1141 17887 1193 17892
rect 1208 17926 1260 17939
rect 1208 17892 1231 17926
rect 1231 17892 1260 17926
rect 1208 17887 1260 17892
<< metal2 >>
rect 14279 35712 14285 35764
rect 14337 35712 14349 35764
rect 14401 35712 14407 35764
rect 14279 35684 14407 35712
rect 14279 35632 14285 35684
rect 14337 35632 14349 35684
rect 14401 35632 14407 35684
rect 14279 35604 14407 35632
rect 14279 35552 14285 35604
rect 14337 35552 14349 35604
rect 14401 35552 14407 35604
rect 460 32764 688 32773
rect 460 32708 465 32764
rect 521 32708 623 32764
rect 679 32708 688 32764
rect 460 32683 688 32708
rect 460 32627 465 32683
rect 521 32627 623 32683
rect 679 32627 688 32683
rect 460 32601 688 32627
rect 460 32545 465 32601
rect 521 32545 623 32601
rect 679 32545 688 32601
rect 460 32519 688 32545
rect 460 32463 465 32519
rect 521 32463 623 32519
rect 679 32463 688 32519
rect 460 32437 688 32463
rect 460 32381 465 32437
rect 521 32381 623 32437
rect 679 32381 688 32437
rect 460 32355 688 32381
rect 460 32299 465 32355
rect 521 32299 623 32355
rect 679 32299 688 32355
rect 460 32273 688 32299
rect 460 32217 465 32273
rect 521 32217 623 32273
rect 679 32217 688 32273
rect 460 32191 688 32217
rect 460 32135 465 32191
rect 521 32135 623 32191
rect 679 32135 688 32191
rect 460 32109 688 32135
rect 460 32053 465 32109
rect 521 32053 623 32109
rect 679 32053 688 32109
rect 460 32027 688 32053
rect 14259 32761 14667 32770
rect 14315 32705 14347 32761
rect 14403 32705 14435 32761
rect 14491 32705 14523 32761
rect 14579 32705 14611 32761
rect 14259 32681 14667 32705
rect 14315 32625 14347 32681
rect 14403 32625 14435 32681
rect 14491 32625 14523 32681
rect 14579 32625 14611 32681
rect 14259 32601 14667 32625
rect 14315 32545 14347 32601
rect 14403 32545 14435 32601
rect 14491 32545 14523 32601
rect 14579 32545 14611 32601
rect 14259 32521 14667 32545
rect 14315 32465 14347 32521
rect 14403 32465 14435 32521
rect 14491 32465 14523 32521
rect 14579 32465 14611 32521
rect 14259 32441 14667 32465
rect 14315 32385 14347 32441
rect 14403 32385 14435 32441
rect 14491 32385 14523 32441
rect 14579 32385 14611 32441
rect 14259 32361 14667 32385
rect 14315 32305 14347 32361
rect 14403 32305 14435 32361
rect 14491 32305 14523 32361
rect 14579 32305 14611 32361
rect 14259 32281 14667 32305
rect 14315 32225 14347 32281
rect 14403 32225 14435 32281
rect 14491 32225 14523 32281
rect 14579 32225 14611 32281
rect 14259 32201 14667 32225
rect 14315 32145 14347 32201
rect 14403 32145 14435 32201
rect 14491 32145 14523 32201
rect 14579 32145 14611 32201
rect 14259 32121 14667 32145
rect 14315 32065 14347 32121
rect 14403 32065 14435 32121
rect 14491 32065 14523 32121
rect 14579 32065 14611 32121
rect 14259 32041 14667 32065
rect 521 31971 623 32027
rect 465 31945 679 31971
rect 521 31889 623 31945
rect 465 31863 679 31889
rect 521 31807 623 31863
rect 465 31781 679 31807
rect 521 31725 623 31781
rect 465 31699 679 31725
rect 521 31643 623 31699
rect 465 31617 679 31643
rect 521 31561 623 31617
rect 465 31535 679 31561
rect 521 31479 623 31535
rect 465 31453 679 31479
rect 521 31397 623 31453
rect 465 31371 679 31397
rect 521 31315 623 31371
rect 465 31289 679 31315
rect 521 31233 623 31289
rect 465 31207 679 31233
rect 521 31151 623 31207
rect 465 31125 679 31151
rect 521 31069 623 31125
rect 465 31043 679 31069
rect 521 30987 623 31043
rect 465 30961 679 30987
rect 521 30905 623 30961
rect 465 30879 679 30905
rect 521 30823 623 30879
rect 465 30797 679 30823
rect 521 30741 623 30797
rect 465 30715 679 30741
rect 521 30659 623 30715
rect 465 30633 679 30659
rect 521 30577 623 30633
rect 465 30551 679 30577
rect 521 30495 623 30551
rect 465 30469 679 30495
rect 521 30413 623 30469
rect 465 30387 679 30413
rect 521 30331 623 30387
rect 465 30305 679 30331
rect 521 30249 623 30305
rect 465 30223 679 30249
rect 521 30167 623 30223
rect 465 30141 679 30167
rect 521 30085 623 30141
rect 465 30059 679 30085
rect 521 30003 623 30059
rect 465 29977 679 30003
rect 521 29921 623 29977
rect 465 29895 679 29921
rect 521 29839 623 29895
rect 465 29813 679 29839
rect 521 29757 623 29813
rect 465 29731 679 29757
rect 521 29675 623 29731
rect 465 29649 679 29675
rect 521 29593 623 29649
rect 465 29567 679 29593
rect 521 29511 623 29567
rect 465 29485 679 29511
rect 521 29429 623 29485
rect 465 29420 679 29429
rect 862 32018 1052 32027
rect 918 31962 996 32018
rect 862 31936 1052 31962
rect 918 31880 996 31936
rect 862 31854 1052 31880
rect 918 31798 996 31854
rect 862 31772 1052 31798
rect 918 31716 996 31772
rect 862 31690 1052 31716
rect 918 31634 996 31690
rect 862 31608 1052 31634
rect 918 31552 996 31608
rect 862 31526 1052 31552
rect 918 31470 996 31526
rect 862 31444 1052 31470
rect 918 31388 996 31444
rect 862 31362 1052 31388
rect 918 31306 996 31362
rect 862 31280 1052 31306
rect 918 31224 996 31280
rect 862 31198 1052 31224
rect 918 31142 996 31198
rect 862 31116 1052 31142
rect 918 31060 996 31116
rect 862 31034 1052 31060
rect 918 30978 996 31034
rect 862 30952 1052 30978
rect 918 30896 996 30952
rect 862 30870 1052 30896
rect 918 30814 996 30870
rect 862 30788 1052 30814
rect 918 30732 996 30788
rect 862 30706 1052 30732
rect 918 30650 996 30706
rect 862 30624 1052 30650
rect 918 30568 996 30624
rect 862 30542 1052 30568
rect 918 30486 996 30542
rect 862 30460 1052 30486
rect 918 30404 996 30460
rect 862 30378 1052 30404
rect 918 30322 996 30378
rect 862 30296 1052 30322
rect 918 30240 996 30296
rect 862 30214 1052 30240
rect 918 30158 996 30214
rect 862 30132 1052 30158
rect 918 30076 996 30132
rect 862 30050 1052 30076
rect 918 29994 996 30050
rect 862 29968 1052 29994
rect 918 29912 996 29968
rect 862 29886 1052 29912
rect 918 29830 996 29886
rect 862 29804 1052 29830
rect 918 29748 996 29804
rect 862 29722 1052 29748
rect 918 29666 996 29722
rect 862 29640 1052 29666
rect 918 29584 996 29640
rect 862 29558 1052 29584
rect 918 29502 996 29558
rect 862 29476 1052 29502
rect 918 29420 996 29476
rect 1395 32018 1577 32027
rect 1451 31962 1521 32018
rect 1395 31937 1577 31962
rect 1451 31881 1521 31937
rect 1395 31856 1577 31881
rect 1451 31800 1521 31856
rect 1395 31775 1577 31800
rect 1451 31719 1521 31775
rect 1395 31694 1577 31719
rect 1451 31638 1521 31694
rect 1395 31613 1577 31638
rect 1451 31557 1521 31613
rect 1395 31532 1577 31557
rect 1451 31476 1521 31532
rect 1395 31451 1577 31476
rect 1451 31395 1521 31451
rect 1395 31370 1577 31395
rect 1451 31314 1521 31370
rect 1395 31289 1577 31314
rect 1451 31233 1521 31289
rect 1395 31207 1577 31233
rect 1451 31151 1521 31207
rect 1395 31125 1577 31151
rect 1451 31069 1521 31125
rect 1395 31043 1577 31069
rect 1451 30987 1521 31043
rect 1395 30961 1577 30987
rect 1451 30905 1521 30961
rect 1395 30879 1577 30905
rect 1451 30823 1521 30879
rect 1395 30797 1577 30823
rect 1451 30741 1521 30797
rect 1395 30715 1577 30741
rect 1451 30659 1521 30715
rect 1395 30633 1577 30659
rect 1451 30577 1521 30633
rect 1395 30551 1577 30577
rect 1451 30495 1521 30551
rect 1395 30469 1577 30495
rect 1451 30413 1521 30469
rect 1395 30387 1577 30413
rect 1451 30331 1521 30387
rect 1395 30305 1577 30331
rect 1451 30249 1521 30305
rect 1395 30223 1577 30249
rect 1451 30167 1521 30223
rect 1395 30141 1577 30167
rect 1451 30085 1521 30141
rect 1395 30059 1577 30085
rect 1451 30003 1521 30059
rect 1395 29977 1577 30003
rect 1451 29921 1521 29977
rect 1395 29895 1577 29921
rect 1451 29839 1521 29895
rect 1395 29813 1577 29839
rect 1451 29757 1521 29813
rect 1395 29731 1577 29757
rect 1451 29675 1521 29731
rect 1395 29649 1577 29675
rect 1451 29593 1521 29649
rect 1395 29567 1577 29593
rect 1451 29511 1521 29567
rect 1395 29485 1577 29511
rect 1451 29429 1521 29485
rect 1395 29420 1577 29429
rect 1891 32018 2073 32027
rect 1947 31962 2017 32018
rect 1891 31936 2073 31962
rect 1947 31880 2017 31936
rect 1891 31854 2073 31880
rect 1947 31798 2017 31854
rect 1891 31772 2073 31798
rect 1947 31716 2017 31772
rect 1891 31690 2073 31716
rect 1947 31634 2017 31690
rect 1891 31608 2073 31634
rect 1947 31552 2017 31608
rect 1891 31526 2073 31552
rect 1947 31470 2017 31526
rect 1891 31444 2073 31470
rect 1947 31388 2017 31444
rect 1891 31362 2073 31388
rect 1947 31306 2017 31362
rect 1891 31280 2073 31306
rect 1947 31224 2017 31280
rect 1891 31198 2073 31224
rect 1947 31142 2017 31198
rect 1891 31116 2073 31142
rect 1947 31060 2017 31116
rect 1891 31034 2073 31060
rect 1947 30978 2017 31034
rect 1891 30952 2073 30978
rect 1947 30896 2017 30952
rect 1891 30870 2073 30896
rect 1947 30814 2017 30870
rect 1891 30788 2073 30814
rect 1947 30732 2017 30788
rect 1891 30706 2073 30732
rect 1947 30650 2017 30706
rect 1891 30624 2073 30650
rect 1947 30568 2017 30624
rect 1891 30542 2073 30568
rect 1947 30486 2017 30542
rect 1891 30460 2073 30486
rect 1947 30404 2017 30460
rect 1891 30378 2073 30404
rect 1947 30322 2017 30378
rect 1891 30296 2073 30322
rect 1947 30240 2017 30296
rect 1891 30214 2073 30240
rect 1947 30158 2017 30214
rect 1891 30132 2073 30158
rect 1947 30076 2017 30132
rect 1891 30050 2073 30076
rect 1947 29994 2017 30050
rect 1891 29968 2073 29994
rect 1947 29912 2017 29968
rect 1891 29886 2073 29912
rect 1947 29830 2017 29886
rect 1891 29804 2073 29830
rect 1947 29748 2017 29804
rect 1891 29722 2073 29748
rect 1947 29666 2017 29722
rect 1891 29640 2073 29666
rect 1947 29584 2017 29640
rect 1891 29558 2073 29584
rect 1947 29502 2017 29558
rect 1891 29476 2073 29502
rect 1947 29420 2017 29476
rect 2387 32018 2569 32027
rect 2443 31962 2513 32018
rect 2387 31936 2569 31962
rect 2443 31880 2513 31936
rect 2387 31854 2569 31880
rect 2443 31798 2513 31854
rect 2387 31772 2569 31798
rect 2443 31716 2513 31772
rect 2387 31690 2569 31716
rect 2443 31634 2513 31690
rect 2387 31608 2569 31634
rect 2443 31552 2513 31608
rect 2387 31526 2569 31552
rect 2443 31470 2513 31526
rect 2387 31444 2569 31470
rect 2443 31388 2513 31444
rect 2387 31362 2569 31388
rect 2443 31306 2513 31362
rect 2387 31280 2569 31306
rect 2443 31224 2513 31280
rect 2387 31198 2569 31224
rect 2443 31142 2513 31198
rect 2387 31116 2569 31142
rect 2443 31060 2513 31116
rect 2387 31034 2569 31060
rect 2443 30978 2513 31034
rect 2387 30952 2569 30978
rect 2443 30896 2513 30952
rect 2387 30870 2569 30896
rect 2443 30814 2513 30870
rect 2387 30788 2569 30814
rect 2443 30732 2513 30788
rect 2387 30706 2569 30732
rect 2443 30650 2513 30706
rect 2387 30624 2569 30650
rect 2443 30568 2513 30624
rect 2387 30542 2569 30568
rect 2443 30486 2513 30542
rect 2387 30460 2569 30486
rect 2443 30404 2513 30460
rect 2387 30378 2569 30404
rect 2443 30322 2513 30378
rect 2387 30296 2569 30322
rect 2443 30240 2513 30296
rect 2387 30214 2569 30240
rect 2443 30158 2513 30214
rect 2387 30132 2569 30158
rect 2443 30076 2513 30132
rect 2387 30050 2569 30076
rect 2443 29994 2513 30050
rect 2387 29968 2569 29994
rect 2443 29912 2513 29968
rect 2387 29886 2569 29912
rect 2443 29830 2513 29886
rect 2387 29804 2569 29830
rect 2443 29748 2513 29804
rect 2387 29722 2569 29748
rect 2443 29666 2513 29722
rect 2387 29640 2569 29666
rect 2443 29584 2513 29640
rect 2387 29558 2569 29584
rect 2443 29502 2513 29558
rect 2387 29476 2569 29502
rect 2443 29420 2513 29476
rect 2883 32018 3065 32027
rect 2939 31962 3009 32018
rect 2883 31936 3065 31962
rect 2939 31880 3009 31936
rect 2883 31854 3065 31880
rect 2939 31798 3009 31854
rect 2883 31772 3065 31798
rect 2939 31716 3009 31772
rect 2883 31690 3065 31716
rect 2939 31634 3009 31690
rect 2883 31608 3065 31634
rect 2939 31552 3009 31608
rect 2883 31526 3065 31552
rect 2939 31470 3009 31526
rect 2883 31444 3065 31470
rect 2939 31388 3009 31444
rect 2883 31362 3065 31388
rect 2939 31306 3009 31362
rect 2883 31280 3065 31306
rect 2939 31224 3009 31280
rect 2883 31198 3065 31224
rect 2939 31142 3009 31198
rect 2883 31116 3065 31142
rect 2939 31060 3009 31116
rect 2883 31034 3065 31060
rect 2939 30978 3009 31034
rect 2883 30952 3065 30978
rect 2939 30896 3009 30952
rect 2883 30870 3065 30896
rect 2939 30814 3009 30870
rect 2883 30788 3065 30814
rect 2939 30732 3009 30788
rect 2883 30706 3065 30732
rect 2939 30650 3009 30706
rect 2883 30624 3065 30650
rect 2939 30568 3009 30624
rect 2883 30542 3065 30568
rect 2939 30486 3009 30542
rect 2883 30460 3065 30486
rect 2939 30404 3009 30460
rect 2883 30378 3065 30404
rect 2939 30322 3009 30378
rect 2883 30296 3065 30322
rect 2939 30240 3009 30296
rect 2883 30214 3065 30240
rect 2939 30158 3009 30214
rect 2883 30132 3065 30158
rect 2939 30076 3009 30132
rect 2883 30050 3065 30076
rect 2939 29994 3009 30050
rect 2883 29968 3065 29994
rect 2939 29912 3009 29968
rect 2883 29886 3065 29912
rect 2939 29830 3009 29886
rect 2883 29804 3065 29830
rect 2939 29748 3009 29804
rect 2883 29722 3065 29748
rect 2939 29666 3009 29722
rect 2883 29640 3065 29666
rect 2939 29584 3009 29640
rect 2883 29558 3065 29584
rect 2939 29502 3009 29558
rect 2883 29476 3065 29502
rect 2939 29420 3009 29476
rect 3379 32018 3561 32027
rect 3435 31962 3505 32018
rect 3379 31936 3561 31962
rect 3435 31880 3505 31936
rect 3379 31854 3561 31880
rect 3435 31798 3505 31854
rect 3379 31772 3561 31798
rect 3435 31716 3505 31772
rect 3379 31690 3561 31716
rect 3435 31634 3505 31690
rect 3379 31608 3561 31634
rect 3435 31552 3505 31608
rect 3379 31526 3561 31552
rect 3435 31470 3505 31526
rect 3379 31444 3561 31470
rect 3435 31388 3505 31444
rect 3379 31362 3561 31388
rect 3435 31306 3505 31362
rect 3379 31280 3561 31306
rect 3435 31224 3505 31280
rect 3379 31198 3561 31224
rect 3435 31142 3505 31198
rect 3379 31116 3561 31142
rect 3435 31060 3505 31116
rect 3379 31034 3561 31060
rect 3435 30978 3505 31034
rect 3379 30952 3561 30978
rect 3435 30896 3505 30952
rect 3379 30870 3561 30896
rect 3435 30814 3505 30870
rect 3379 30788 3561 30814
rect 3435 30732 3505 30788
rect 3379 30706 3561 30732
rect 3435 30650 3505 30706
rect 3379 30624 3561 30650
rect 3435 30568 3505 30624
rect 3379 30542 3561 30568
rect 3435 30486 3505 30542
rect 3379 30460 3561 30486
rect 3435 30404 3505 30460
rect 3379 30378 3561 30404
rect 3435 30322 3505 30378
rect 3379 30296 3561 30322
rect 3435 30240 3505 30296
rect 3379 30214 3561 30240
rect 3435 30158 3505 30214
rect 3379 30132 3561 30158
rect 3435 30076 3505 30132
rect 3379 30050 3561 30076
rect 3435 29994 3505 30050
rect 3379 29968 3561 29994
rect 3435 29912 3505 29968
rect 3379 29886 3561 29912
rect 3435 29830 3505 29886
rect 3379 29804 3561 29830
rect 3435 29748 3505 29804
rect 3379 29722 3561 29748
rect 3435 29666 3505 29722
rect 3379 29640 3561 29666
rect 3435 29584 3505 29640
rect 3379 29558 3561 29584
rect 3435 29502 3505 29558
rect 3379 29476 3561 29502
rect 3435 29420 3505 29476
rect 3875 32018 4057 32027
rect 3931 31962 4001 32018
rect 3875 31936 4057 31962
rect 3931 31880 4001 31936
rect 3875 31854 4057 31880
rect 3931 31798 4001 31854
rect 3875 31772 4057 31798
rect 3931 31716 4001 31772
rect 3875 31690 4057 31716
rect 3931 31634 4001 31690
rect 3875 31608 4057 31634
rect 3931 31552 4001 31608
rect 3875 31526 4057 31552
rect 3931 31470 4001 31526
rect 3875 31444 4057 31470
rect 3931 31388 4001 31444
rect 3875 31362 4057 31388
rect 3931 31306 4001 31362
rect 3875 31280 4057 31306
rect 3931 31224 4001 31280
rect 3875 31198 4057 31224
rect 3931 31142 4001 31198
rect 3875 31116 4057 31142
rect 3931 31060 4001 31116
rect 3875 31034 4057 31060
rect 3931 30978 4001 31034
rect 3875 30952 4057 30978
rect 3931 30896 4001 30952
rect 3875 30870 4057 30896
rect 3931 30814 4001 30870
rect 3875 30788 4057 30814
rect 3931 30732 4001 30788
rect 3875 30706 4057 30732
rect 3931 30650 4001 30706
rect 3875 30624 4057 30650
rect 3931 30568 4001 30624
rect 3875 30542 4057 30568
rect 3931 30486 4001 30542
rect 3875 30460 4057 30486
rect 3931 30404 4001 30460
rect 3875 30378 4057 30404
rect 3931 30322 4001 30378
rect 3875 30296 4057 30322
rect 3931 30240 4001 30296
rect 3875 30214 4057 30240
rect 3931 30158 4001 30214
rect 3875 30132 4057 30158
rect 3931 30076 4001 30132
rect 3875 30050 4057 30076
rect 3931 29994 4001 30050
rect 3875 29968 4057 29994
rect 3931 29912 4001 29968
rect 3875 29886 4057 29912
rect 3931 29830 4001 29886
rect 3875 29804 4057 29830
rect 3931 29748 4001 29804
rect 3875 29722 4057 29748
rect 3931 29666 4001 29722
rect 3875 29640 4057 29666
rect 3931 29584 4001 29640
rect 3875 29558 4057 29584
rect 3931 29502 4001 29558
rect 3875 29476 4057 29502
rect 3931 29420 4001 29476
rect 4371 32018 4553 32027
rect 4427 31962 4497 32018
rect 4371 31936 4553 31962
rect 4427 31880 4497 31936
rect 4371 31854 4553 31880
rect 4427 31798 4497 31854
rect 4371 31772 4553 31798
rect 4427 31716 4497 31772
rect 4371 31690 4553 31716
rect 4427 31634 4497 31690
rect 4371 31608 4553 31634
rect 4427 31552 4497 31608
rect 4371 31526 4553 31552
rect 4427 31470 4497 31526
rect 4371 31444 4553 31470
rect 4427 31388 4497 31444
rect 4371 31362 4553 31388
rect 4427 31306 4497 31362
rect 4371 31280 4553 31306
rect 4427 31224 4497 31280
rect 4371 31198 4553 31224
rect 4427 31142 4497 31198
rect 4371 31116 4553 31142
rect 4427 31060 4497 31116
rect 4371 31034 4553 31060
rect 4427 30978 4497 31034
rect 4371 30952 4553 30978
rect 4427 30896 4497 30952
rect 4371 30870 4553 30896
rect 4427 30814 4497 30870
rect 4371 30788 4553 30814
rect 4427 30732 4497 30788
rect 4371 30706 4553 30732
rect 4427 30650 4497 30706
rect 4371 30624 4553 30650
rect 4427 30568 4497 30624
rect 4371 30542 4553 30568
rect 4427 30486 4497 30542
rect 4371 30460 4553 30486
rect 4427 30404 4497 30460
rect 4371 30378 4553 30404
rect 4427 30322 4497 30378
rect 4371 30296 4553 30322
rect 4427 30240 4497 30296
rect 4371 30214 4553 30240
rect 4427 30158 4497 30214
rect 4371 30132 4553 30158
rect 4427 30076 4497 30132
rect 4371 30050 4553 30076
rect 4427 29994 4497 30050
rect 4371 29968 4553 29994
rect 4427 29912 4497 29968
rect 4371 29886 4553 29912
rect 4427 29830 4497 29886
rect 4371 29804 4553 29830
rect 4427 29748 4497 29804
rect 4371 29722 4553 29748
rect 4427 29666 4497 29722
rect 4371 29640 4553 29666
rect 4427 29584 4497 29640
rect 4371 29558 4553 29584
rect 4427 29502 4497 29558
rect 4371 29476 4553 29502
rect 4427 29420 4497 29476
rect 4867 32018 5049 32027
rect 4923 31962 4993 32018
rect 4867 31936 5049 31962
rect 4923 31880 4993 31936
rect 4867 31854 5049 31880
rect 4923 31798 4993 31854
rect 4867 31772 5049 31798
rect 4923 31716 4993 31772
rect 4867 31690 5049 31716
rect 4923 31634 4993 31690
rect 4867 31608 5049 31634
rect 4923 31552 4993 31608
rect 4867 31526 5049 31552
rect 4923 31470 4993 31526
rect 4867 31444 5049 31470
rect 4923 31388 4993 31444
rect 4867 31362 5049 31388
rect 4923 31306 4993 31362
rect 4867 31280 5049 31306
rect 4923 31224 4993 31280
rect 4867 31198 5049 31224
rect 4923 31142 4993 31198
rect 4867 31116 5049 31142
rect 4923 31060 4993 31116
rect 4867 31034 5049 31060
rect 4923 30978 4993 31034
rect 4867 30952 5049 30978
rect 4923 30896 4993 30952
rect 4867 30870 5049 30896
rect 4923 30814 4993 30870
rect 4867 30788 5049 30814
rect 4923 30732 4993 30788
rect 4867 30706 5049 30732
rect 4923 30650 4993 30706
rect 4867 30624 5049 30650
rect 4923 30568 4993 30624
rect 4867 30542 5049 30568
rect 4923 30486 4993 30542
rect 4867 30460 5049 30486
rect 4923 30404 4993 30460
rect 4867 30378 5049 30404
rect 4923 30322 4993 30378
rect 4867 30296 5049 30322
rect 4923 30240 4993 30296
rect 4867 30214 5049 30240
rect 4923 30158 4993 30214
rect 4867 30132 5049 30158
rect 4923 30076 4993 30132
rect 4867 30050 5049 30076
rect 4923 29994 4993 30050
rect 4867 29968 5049 29994
rect 4923 29912 4993 29968
rect 4867 29886 5049 29912
rect 4923 29830 4993 29886
rect 4867 29804 5049 29830
rect 4923 29748 4993 29804
rect 4867 29722 5049 29748
rect 4923 29666 4993 29722
rect 4867 29640 5049 29666
rect 4923 29584 4993 29640
rect 4867 29558 5049 29584
rect 4923 29502 4993 29558
rect 4867 29476 5049 29502
rect 4923 29420 4993 29476
rect 5363 32018 5545 32027
rect 5419 31962 5489 32018
rect 5363 31936 5545 31962
rect 5419 31880 5489 31936
rect 5363 31854 5545 31880
rect 5419 31798 5489 31854
rect 5363 31772 5545 31798
rect 5419 31716 5489 31772
rect 5363 31690 5545 31716
rect 5419 31634 5489 31690
rect 5363 31608 5545 31634
rect 5419 31552 5489 31608
rect 5363 31526 5545 31552
rect 5419 31470 5489 31526
rect 5363 31444 5545 31470
rect 5419 31388 5489 31444
rect 5363 31362 5545 31388
rect 5419 31306 5489 31362
rect 5363 31280 5545 31306
rect 5419 31224 5489 31280
rect 5363 31198 5545 31224
rect 5419 31142 5489 31198
rect 5363 31116 5545 31142
rect 5419 31060 5489 31116
rect 5363 31034 5545 31060
rect 5419 30978 5489 31034
rect 5363 30952 5545 30978
rect 5419 30896 5489 30952
rect 5363 30870 5545 30896
rect 5419 30814 5489 30870
rect 5363 30788 5545 30814
rect 5419 30732 5489 30788
rect 5363 30706 5545 30732
rect 5419 30650 5489 30706
rect 5363 30624 5545 30650
rect 5419 30568 5489 30624
rect 5363 30542 5545 30568
rect 5419 30486 5489 30542
rect 5363 30460 5545 30486
rect 5419 30404 5489 30460
rect 5363 30378 5545 30404
rect 5419 30322 5489 30378
rect 5363 30296 5545 30322
rect 5419 30240 5489 30296
rect 5363 30214 5545 30240
rect 5419 30158 5489 30214
rect 5363 30132 5545 30158
rect 5419 30076 5489 30132
rect 5363 30050 5545 30076
rect 5419 29994 5489 30050
rect 5363 29968 5545 29994
rect 5419 29912 5489 29968
rect 5363 29886 5545 29912
rect 5419 29830 5489 29886
rect 5363 29804 5545 29830
rect 5419 29748 5489 29804
rect 5363 29722 5545 29748
rect 5419 29666 5489 29722
rect 5363 29640 5545 29666
rect 5419 29584 5489 29640
rect 5363 29558 5545 29584
rect 5419 29502 5489 29558
rect 5363 29476 5545 29502
rect 5419 29420 5489 29476
rect 5859 32018 6041 32027
rect 5915 31962 5985 32018
rect 5859 31936 6041 31962
rect 5915 31880 5985 31936
rect 5859 31854 6041 31880
rect 5915 31798 5985 31854
rect 5859 31772 6041 31798
rect 5915 31716 5985 31772
rect 5859 31690 6041 31716
rect 5915 31634 5985 31690
rect 5859 31608 6041 31634
rect 5915 31552 5985 31608
rect 5859 31526 6041 31552
rect 5915 31470 5985 31526
rect 5859 31444 6041 31470
rect 5915 31388 5985 31444
rect 5859 31362 6041 31388
rect 5915 31306 5985 31362
rect 5859 31280 6041 31306
rect 5915 31224 5985 31280
rect 5859 31198 6041 31224
rect 5915 31142 5985 31198
rect 5859 31116 6041 31142
rect 5915 31060 5985 31116
rect 5859 31034 6041 31060
rect 5915 30978 5985 31034
rect 5859 30952 6041 30978
rect 5915 30896 5985 30952
rect 5859 30870 6041 30896
rect 5915 30814 5985 30870
rect 5859 30788 6041 30814
rect 5915 30732 5985 30788
rect 5859 30706 6041 30732
rect 5915 30650 5985 30706
rect 5859 30624 6041 30650
rect 5915 30568 5985 30624
rect 5859 30542 6041 30568
rect 5915 30486 5985 30542
rect 5859 30460 6041 30486
rect 5915 30404 5985 30460
rect 5859 30378 6041 30404
rect 5915 30322 5985 30378
rect 5859 30296 6041 30322
rect 5915 30240 5985 30296
rect 5859 30214 6041 30240
rect 5915 30158 5985 30214
rect 5859 30132 6041 30158
rect 5915 30076 5985 30132
rect 5859 30050 6041 30076
rect 5915 29994 5985 30050
rect 5859 29968 6041 29994
rect 5915 29912 5985 29968
rect 5859 29886 6041 29912
rect 5915 29830 5985 29886
rect 5859 29804 6041 29830
rect 5915 29748 5985 29804
rect 5859 29722 6041 29748
rect 5915 29666 5985 29722
rect 5859 29640 6041 29666
rect 5915 29584 5985 29640
rect 5859 29558 6041 29584
rect 5915 29502 5985 29558
rect 5859 29476 6041 29502
rect 5915 29420 5985 29476
rect 6355 32018 6537 32027
rect 6411 31962 6481 32018
rect 6355 31936 6537 31962
rect 6411 31880 6481 31936
rect 6355 31854 6537 31880
rect 6411 31798 6481 31854
rect 6355 31772 6537 31798
rect 6411 31716 6481 31772
rect 6355 31690 6537 31716
rect 6411 31634 6481 31690
rect 6355 31608 6537 31634
rect 6411 31552 6481 31608
rect 6355 31526 6537 31552
rect 6411 31470 6481 31526
rect 6355 31444 6537 31470
rect 6411 31388 6481 31444
rect 6355 31362 6537 31388
rect 6411 31306 6481 31362
rect 6355 31280 6537 31306
rect 6411 31224 6481 31280
rect 6355 31198 6537 31224
rect 6411 31142 6481 31198
rect 6355 31116 6537 31142
rect 6411 31060 6481 31116
rect 6355 31034 6537 31060
rect 6411 30978 6481 31034
rect 6355 30952 6537 30978
rect 6411 30896 6481 30952
rect 6355 30870 6537 30896
rect 6411 30814 6481 30870
rect 6355 30788 6537 30814
rect 6411 30732 6481 30788
rect 6355 30706 6537 30732
rect 6411 30650 6481 30706
rect 6355 30624 6537 30650
rect 6411 30568 6481 30624
rect 6355 30542 6537 30568
rect 6411 30486 6481 30542
rect 6355 30460 6537 30486
rect 6411 30404 6481 30460
rect 6355 30378 6537 30404
rect 6411 30322 6481 30378
rect 6355 30296 6537 30322
rect 6411 30240 6481 30296
rect 6355 30214 6537 30240
rect 6411 30158 6481 30214
rect 6355 30132 6537 30158
rect 6411 30076 6481 30132
rect 6355 30050 6537 30076
rect 6411 29994 6481 30050
rect 6355 29968 6537 29994
rect 6411 29912 6481 29968
rect 6355 29886 6537 29912
rect 6411 29830 6481 29886
rect 6355 29804 6537 29830
rect 6411 29748 6481 29804
rect 6355 29722 6537 29748
rect 6411 29666 6481 29722
rect 6355 29640 6537 29666
rect 6411 29584 6481 29640
rect 6355 29558 6537 29584
rect 6411 29502 6481 29558
rect 6355 29476 6537 29502
rect 6411 29420 6481 29476
rect 6851 32018 7033 32027
rect 6907 31962 6977 32018
rect 6851 31936 7033 31962
rect 6907 31880 6977 31936
rect 6851 31854 7033 31880
rect 6907 31798 6977 31854
rect 6851 31772 7033 31798
rect 6907 31716 6977 31772
rect 6851 31690 7033 31716
rect 6907 31634 6977 31690
rect 6851 31608 7033 31634
rect 6907 31552 6977 31608
rect 6851 31526 7033 31552
rect 6907 31470 6977 31526
rect 6851 31444 7033 31470
rect 6907 31388 6977 31444
rect 6851 31362 7033 31388
rect 6907 31306 6977 31362
rect 6851 31280 7033 31306
rect 6907 31224 6977 31280
rect 6851 31198 7033 31224
rect 6907 31142 6977 31198
rect 6851 31116 7033 31142
rect 6907 31060 6977 31116
rect 6851 31034 7033 31060
rect 6907 30978 6977 31034
rect 6851 30952 7033 30978
rect 6907 30896 6977 30952
rect 6851 30870 7033 30896
rect 6907 30814 6977 30870
rect 6851 30788 7033 30814
rect 6907 30732 6977 30788
rect 6851 30706 7033 30732
rect 6907 30650 6977 30706
rect 6851 30624 7033 30650
rect 6907 30568 6977 30624
rect 6851 30542 7033 30568
rect 6907 30486 6977 30542
rect 6851 30460 7033 30486
rect 6907 30404 6977 30460
rect 6851 30378 7033 30404
rect 6907 30322 6977 30378
rect 6851 30296 7033 30322
rect 6907 30240 6977 30296
rect 6851 30214 7033 30240
rect 6907 30158 6977 30214
rect 6851 30132 7033 30158
rect 6907 30076 6977 30132
rect 6851 30050 7033 30076
rect 6907 29994 6977 30050
rect 6851 29968 7033 29994
rect 6907 29912 6977 29968
rect 6851 29886 7033 29912
rect 6907 29830 6977 29886
rect 6851 29804 7033 29830
rect 6907 29748 6977 29804
rect 6851 29722 7033 29748
rect 6907 29666 6977 29722
rect 6851 29640 7033 29666
rect 6907 29584 6977 29640
rect 6851 29558 7033 29584
rect 6907 29502 6977 29558
rect 6851 29476 7033 29502
rect 6907 29420 6977 29476
rect 7347 32018 7529 32027
rect 7403 31962 7473 32018
rect 7347 31936 7529 31962
rect 7403 31880 7473 31936
rect 7347 31854 7529 31880
rect 7403 31798 7473 31854
rect 7347 31772 7529 31798
rect 7403 31716 7473 31772
rect 7347 31690 7529 31716
rect 7403 31634 7473 31690
rect 7347 31608 7529 31634
rect 7403 31552 7473 31608
rect 7347 31526 7529 31552
rect 7403 31470 7473 31526
rect 7347 31444 7529 31470
rect 7403 31388 7473 31444
rect 7347 31362 7529 31388
rect 7403 31306 7473 31362
rect 7347 31280 7529 31306
rect 7403 31224 7473 31280
rect 7347 31198 7529 31224
rect 7403 31142 7473 31198
rect 7347 31116 7529 31142
rect 7403 31060 7473 31116
rect 7347 31034 7529 31060
rect 7403 30978 7473 31034
rect 7347 30952 7529 30978
rect 7403 30896 7473 30952
rect 7347 30870 7529 30896
rect 7403 30814 7473 30870
rect 7347 30788 7529 30814
rect 7403 30732 7473 30788
rect 7347 30706 7529 30732
rect 7403 30650 7473 30706
rect 7347 30624 7529 30650
rect 7403 30568 7473 30624
rect 7347 30542 7529 30568
rect 7403 30486 7473 30542
rect 7347 30460 7529 30486
rect 7403 30404 7473 30460
rect 7347 30378 7529 30404
rect 7403 30322 7473 30378
rect 7347 30296 7529 30322
rect 7403 30240 7473 30296
rect 7347 30214 7529 30240
rect 7403 30158 7473 30214
rect 7347 30132 7529 30158
rect 7403 30076 7473 30132
rect 7347 30050 7529 30076
rect 7403 29994 7473 30050
rect 7347 29968 7529 29994
rect 7403 29912 7473 29968
rect 7347 29886 7529 29912
rect 7403 29830 7473 29886
rect 7347 29804 7529 29830
rect 7403 29748 7473 29804
rect 7347 29722 7529 29748
rect 7403 29666 7473 29722
rect 7347 29640 7529 29666
rect 7403 29584 7473 29640
rect 7347 29558 7529 29584
rect 7403 29502 7473 29558
rect 7347 29476 7529 29502
rect 7403 29420 7473 29476
rect 7843 32018 8025 32027
rect 7899 31962 7969 32018
rect 7843 31936 8025 31962
rect 7899 31880 7969 31936
rect 7843 31854 8025 31880
rect 7899 31798 7969 31854
rect 7843 31772 8025 31798
rect 7899 31716 7969 31772
rect 7843 31690 8025 31716
rect 7899 31634 7969 31690
rect 7843 31608 8025 31634
rect 7899 31552 7969 31608
rect 7843 31526 8025 31552
rect 7899 31470 7969 31526
rect 7843 31444 8025 31470
rect 7899 31388 7969 31444
rect 7843 31362 8025 31388
rect 7899 31306 7969 31362
rect 7843 31280 8025 31306
rect 7899 31224 7969 31280
rect 7843 31198 8025 31224
rect 7899 31142 7969 31198
rect 7843 31116 8025 31142
rect 7899 31060 7969 31116
rect 7843 31034 8025 31060
rect 7899 30978 7969 31034
rect 7843 30952 8025 30978
rect 7899 30896 7969 30952
rect 7843 30870 8025 30896
rect 7899 30814 7969 30870
rect 7843 30788 8025 30814
rect 7899 30732 7969 30788
rect 7843 30706 8025 30732
rect 7899 30650 7969 30706
rect 7843 30624 8025 30650
rect 7899 30568 7969 30624
rect 7843 30542 8025 30568
rect 7899 30486 7969 30542
rect 7843 30460 8025 30486
rect 7899 30404 7969 30460
rect 7843 30378 8025 30404
rect 7899 30322 7969 30378
rect 7843 30296 8025 30322
rect 7899 30240 7969 30296
rect 7843 30214 8025 30240
rect 7899 30158 7969 30214
rect 7843 30132 8025 30158
rect 7899 30076 7969 30132
rect 7843 30050 8025 30076
rect 7899 29994 7969 30050
rect 7843 29968 8025 29994
rect 7899 29912 7969 29968
rect 7843 29886 8025 29912
rect 7899 29830 7969 29886
rect 7843 29804 8025 29830
rect 7899 29748 7969 29804
rect 7843 29722 8025 29748
rect 7899 29666 7969 29722
rect 7843 29640 8025 29666
rect 7899 29584 7969 29640
rect 7843 29558 8025 29584
rect 7899 29502 7969 29558
rect 7843 29476 8025 29502
rect 7899 29420 7969 29476
rect 8339 32018 8521 32027
rect 8395 31962 8465 32018
rect 8339 31936 8521 31962
rect 8395 31880 8465 31936
rect 8339 31854 8521 31880
rect 8395 31798 8465 31854
rect 8339 31772 8521 31798
rect 8395 31716 8465 31772
rect 8339 31690 8521 31716
rect 8395 31634 8465 31690
rect 8339 31608 8521 31634
rect 8395 31552 8465 31608
rect 8339 31526 8521 31552
rect 8395 31470 8465 31526
rect 8339 31444 8521 31470
rect 8395 31388 8465 31444
rect 8339 31362 8521 31388
rect 8395 31306 8465 31362
rect 8339 31280 8521 31306
rect 8395 31224 8465 31280
rect 8339 31198 8521 31224
rect 8395 31142 8465 31198
rect 8339 31116 8521 31142
rect 8395 31060 8465 31116
rect 8339 31034 8521 31060
rect 8395 30978 8465 31034
rect 8339 30952 8521 30978
rect 8395 30896 8465 30952
rect 8339 30870 8521 30896
rect 8395 30814 8465 30870
rect 8339 30788 8521 30814
rect 8395 30732 8465 30788
rect 8339 30706 8521 30732
rect 8395 30650 8465 30706
rect 8339 30624 8521 30650
rect 8395 30568 8465 30624
rect 8339 30542 8521 30568
rect 8395 30486 8465 30542
rect 8339 30460 8521 30486
rect 8395 30404 8465 30460
rect 8339 30378 8521 30404
rect 8395 30322 8465 30378
rect 8339 30296 8521 30322
rect 8395 30240 8465 30296
rect 8339 30214 8521 30240
rect 8395 30158 8465 30214
rect 8339 30132 8521 30158
rect 8395 30076 8465 30132
rect 8339 30050 8521 30076
rect 8395 29994 8465 30050
rect 8339 29968 8521 29994
rect 8395 29912 8465 29968
rect 8339 29886 8521 29912
rect 8395 29830 8465 29886
rect 8339 29804 8521 29830
rect 8395 29748 8465 29804
rect 8339 29722 8521 29748
rect 8395 29666 8465 29722
rect 8339 29640 8521 29666
rect 8395 29584 8465 29640
rect 8339 29558 8521 29584
rect 8395 29502 8465 29558
rect 8339 29476 8521 29502
rect 8395 29420 8465 29476
rect 8835 32018 9017 32027
rect 8891 31962 8961 32018
rect 8835 31936 9017 31962
rect 8891 31880 8961 31936
rect 8835 31854 9017 31880
rect 8891 31798 8961 31854
rect 8835 31772 9017 31798
rect 8891 31716 8961 31772
rect 8835 31690 9017 31716
rect 8891 31634 8961 31690
rect 8835 31608 9017 31634
rect 8891 31552 8961 31608
rect 8835 31526 9017 31552
rect 8891 31470 8961 31526
rect 8835 31444 9017 31470
rect 8891 31388 8961 31444
rect 8835 31362 9017 31388
rect 8891 31306 8961 31362
rect 8835 31280 9017 31306
rect 8891 31224 8961 31280
rect 8835 31198 9017 31224
rect 8891 31142 8961 31198
rect 8835 31116 9017 31142
rect 8891 31060 8961 31116
rect 8835 31034 9017 31060
rect 8891 30978 8961 31034
rect 8835 30952 9017 30978
rect 8891 30896 8961 30952
rect 8835 30870 9017 30896
rect 8891 30814 8961 30870
rect 8835 30788 9017 30814
rect 8891 30732 8961 30788
rect 8835 30706 9017 30732
rect 8891 30650 8961 30706
rect 8835 30624 9017 30650
rect 8891 30568 8961 30624
rect 8835 30542 9017 30568
rect 8891 30486 8961 30542
rect 8835 30460 9017 30486
rect 8891 30404 8961 30460
rect 8835 30378 9017 30404
rect 8891 30322 8961 30378
rect 8835 30296 9017 30322
rect 8891 30240 8961 30296
rect 8835 30214 9017 30240
rect 8891 30158 8961 30214
rect 8835 30132 9017 30158
rect 8891 30076 8961 30132
rect 8835 30050 9017 30076
rect 8891 29994 8961 30050
rect 8835 29968 9017 29994
rect 8891 29912 8961 29968
rect 8835 29886 9017 29912
rect 8891 29830 8961 29886
rect 8835 29804 9017 29830
rect 8891 29748 8961 29804
rect 8835 29722 9017 29748
rect 8891 29666 8961 29722
rect 8835 29640 9017 29666
rect 8891 29584 8961 29640
rect 8835 29558 9017 29584
rect 8891 29502 8961 29558
rect 8835 29476 9017 29502
rect 8891 29420 8961 29476
rect 9331 32018 9513 32027
rect 9387 31962 9457 32018
rect 9331 31936 9513 31962
rect 9387 31880 9457 31936
rect 9331 31854 9513 31880
rect 9387 31798 9457 31854
rect 9331 31772 9513 31798
rect 9387 31716 9457 31772
rect 9331 31690 9513 31716
rect 9387 31634 9457 31690
rect 9331 31608 9513 31634
rect 9387 31552 9457 31608
rect 9331 31526 9513 31552
rect 9387 31470 9457 31526
rect 9331 31444 9513 31470
rect 9387 31388 9457 31444
rect 9331 31362 9513 31388
rect 9387 31306 9457 31362
rect 9331 31280 9513 31306
rect 9387 31224 9457 31280
rect 9331 31198 9513 31224
rect 9387 31142 9457 31198
rect 9331 31116 9513 31142
rect 9387 31060 9457 31116
rect 9331 31034 9513 31060
rect 9387 30978 9457 31034
rect 9331 30952 9513 30978
rect 9387 30896 9457 30952
rect 9331 30870 9513 30896
rect 9387 30814 9457 30870
rect 9331 30788 9513 30814
rect 9387 30732 9457 30788
rect 9331 30706 9513 30732
rect 9387 30650 9457 30706
rect 9331 30624 9513 30650
rect 9387 30568 9457 30624
rect 9331 30542 9513 30568
rect 9387 30486 9457 30542
rect 9331 30460 9513 30486
rect 9387 30404 9457 30460
rect 9331 30378 9513 30404
rect 9387 30322 9457 30378
rect 9331 30296 9513 30322
rect 9387 30240 9457 30296
rect 9331 30214 9513 30240
rect 9387 30158 9457 30214
rect 9331 30132 9513 30158
rect 9387 30076 9457 30132
rect 9331 30050 9513 30076
rect 9387 29994 9457 30050
rect 9331 29968 9513 29994
rect 9387 29912 9457 29968
rect 9331 29886 9513 29912
rect 9387 29830 9457 29886
rect 9331 29804 9513 29830
rect 9387 29748 9457 29804
rect 9331 29722 9513 29748
rect 9387 29666 9457 29722
rect 9331 29640 9513 29666
rect 9387 29584 9457 29640
rect 9331 29558 9513 29584
rect 9387 29502 9457 29558
rect 9331 29476 9513 29502
rect 9387 29420 9457 29476
rect 9827 32018 10009 32027
rect 9883 31962 9953 32018
rect 9827 31936 10009 31962
rect 9883 31880 9953 31936
rect 9827 31854 10009 31880
rect 9883 31798 9953 31854
rect 9827 31772 10009 31798
rect 9883 31716 9953 31772
rect 9827 31690 10009 31716
rect 9883 31634 9953 31690
rect 9827 31608 10009 31634
rect 9883 31552 9953 31608
rect 9827 31526 10009 31552
rect 9883 31470 9953 31526
rect 9827 31444 10009 31470
rect 9883 31388 9953 31444
rect 9827 31362 10009 31388
rect 9883 31306 9953 31362
rect 9827 31280 10009 31306
rect 9883 31224 9953 31280
rect 9827 31198 10009 31224
rect 9883 31142 9953 31198
rect 9827 31116 10009 31142
rect 9883 31060 9953 31116
rect 9827 31034 10009 31060
rect 9883 30978 9953 31034
rect 9827 30952 10009 30978
rect 9883 30896 9953 30952
rect 9827 30870 10009 30896
rect 9883 30814 9953 30870
rect 9827 30788 10009 30814
rect 9883 30732 9953 30788
rect 9827 30706 10009 30732
rect 9883 30650 9953 30706
rect 9827 30624 10009 30650
rect 9883 30568 9953 30624
rect 9827 30542 10009 30568
rect 9883 30486 9953 30542
rect 9827 30460 10009 30486
rect 9883 30404 9953 30460
rect 9827 30378 10009 30404
rect 9883 30322 9953 30378
rect 9827 30296 10009 30322
rect 9883 30240 9953 30296
rect 9827 30214 10009 30240
rect 9883 30158 9953 30214
rect 9827 30132 10009 30158
rect 9883 30076 9953 30132
rect 9827 30050 10009 30076
rect 9883 29994 9953 30050
rect 9827 29968 10009 29994
rect 9883 29912 9953 29968
rect 9827 29886 10009 29912
rect 9883 29830 9953 29886
rect 9827 29804 10009 29830
rect 9883 29748 9953 29804
rect 9827 29722 10009 29748
rect 9883 29666 9953 29722
rect 9827 29640 10009 29666
rect 9883 29584 9953 29640
rect 9827 29558 10009 29584
rect 9883 29502 9953 29558
rect 9827 29476 10009 29502
rect 9883 29420 9953 29476
rect 10323 32018 10505 32027
rect 10379 31962 10449 32018
rect 10323 31936 10505 31962
rect 10379 31880 10449 31936
rect 10323 31854 10505 31880
rect 10379 31798 10449 31854
rect 10323 31772 10505 31798
rect 10379 31716 10449 31772
rect 10323 31690 10505 31716
rect 10379 31634 10449 31690
rect 10323 31608 10505 31634
rect 10379 31552 10449 31608
rect 10323 31526 10505 31552
rect 10379 31470 10449 31526
rect 10323 31444 10505 31470
rect 10379 31388 10449 31444
rect 10323 31362 10505 31388
rect 10379 31306 10449 31362
rect 10323 31280 10505 31306
rect 10379 31224 10449 31280
rect 10323 31198 10505 31224
rect 10379 31142 10449 31198
rect 10323 31116 10505 31142
rect 10379 31060 10449 31116
rect 10323 31034 10505 31060
rect 10379 30978 10449 31034
rect 10323 30952 10505 30978
rect 10379 30896 10449 30952
rect 10323 30870 10505 30896
rect 10379 30814 10449 30870
rect 10323 30788 10505 30814
rect 10379 30732 10449 30788
rect 10323 30706 10505 30732
rect 10379 30650 10449 30706
rect 10323 30624 10505 30650
rect 10379 30568 10449 30624
rect 10323 30542 10505 30568
rect 10379 30486 10449 30542
rect 10323 30460 10505 30486
rect 10379 30404 10449 30460
rect 10323 30378 10505 30404
rect 10379 30322 10449 30378
rect 10323 30296 10505 30322
rect 10379 30240 10449 30296
rect 10323 30214 10505 30240
rect 10379 30158 10449 30214
rect 10323 30132 10505 30158
rect 10379 30076 10449 30132
rect 10323 30050 10505 30076
rect 10379 29994 10449 30050
rect 10323 29968 10505 29994
rect 10379 29912 10449 29968
rect 10323 29886 10505 29912
rect 10379 29830 10449 29886
rect 10323 29804 10505 29830
rect 10379 29748 10449 29804
rect 10323 29722 10505 29748
rect 10379 29666 10449 29722
rect 10323 29640 10505 29666
rect 10379 29584 10449 29640
rect 10323 29558 10505 29584
rect 10379 29502 10449 29558
rect 10323 29476 10505 29502
rect 10379 29420 10449 29476
rect 10819 32018 11001 32027
rect 10875 31962 10945 32018
rect 10819 31936 11001 31962
rect 10875 31880 10945 31936
rect 10819 31854 11001 31880
rect 10875 31798 10945 31854
rect 10819 31772 11001 31798
rect 10875 31716 10945 31772
rect 10819 31690 11001 31716
rect 10875 31634 10945 31690
rect 10819 31608 11001 31634
rect 10875 31552 10945 31608
rect 10819 31526 11001 31552
rect 10875 31470 10945 31526
rect 10819 31444 11001 31470
rect 10875 31388 10945 31444
rect 10819 31362 11001 31388
rect 10875 31306 10945 31362
rect 10819 31280 11001 31306
rect 10875 31224 10945 31280
rect 10819 31198 11001 31224
rect 10875 31142 10945 31198
rect 10819 31116 11001 31142
rect 10875 31060 10945 31116
rect 10819 31034 11001 31060
rect 10875 30978 10945 31034
rect 10819 30952 11001 30978
rect 10875 30896 10945 30952
rect 10819 30870 11001 30896
rect 10875 30814 10945 30870
rect 10819 30788 11001 30814
rect 10875 30732 10945 30788
rect 10819 30706 11001 30732
rect 10875 30650 10945 30706
rect 10819 30624 11001 30650
rect 10875 30568 10945 30624
rect 10819 30542 11001 30568
rect 10875 30486 10945 30542
rect 10819 30460 11001 30486
rect 10875 30404 10945 30460
rect 10819 30378 11001 30404
rect 10875 30322 10945 30378
rect 10819 30296 11001 30322
rect 10875 30240 10945 30296
rect 10819 30214 11001 30240
rect 10875 30158 10945 30214
rect 10819 30132 11001 30158
rect 10875 30076 10945 30132
rect 10819 30050 11001 30076
rect 10875 29994 10945 30050
rect 10819 29968 11001 29994
rect 10875 29912 10945 29968
rect 10819 29886 11001 29912
rect 10875 29830 10945 29886
rect 10819 29804 11001 29830
rect 10875 29748 10945 29804
rect 10819 29722 11001 29748
rect 10875 29666 10945 29722
rect 10819 29640 11001 29666
rect 10875 29584 10945 29640
rect 10819 29558 11001 29584
rect 10875 29502 10945 29558
rect 10819 29476 11001 29502
rect 10875 29420 10945 29476
rect 11315 32018 11497 32027
rect 11371 31962 11441 32018
rect 11315 31936 11497 31962
rect 11371 31880 11441 31936
rect 11315 31854 11497 31880
rect 11371 31798 11441 31854
rect 11315 31772 11497 31798
rect 11371 31716 11441 31772
rect 11315 31690 11497 31716
rect 11371 31634 11441 31690
rect 11315 31608 11497 31634
rect 11371 31552 11441 31608
rect 11315 31526 11497 31552
rect 11371 31470 11441 31526
rect 11315 31444 11497 31470
rect 11371 31388 11441 31444
rect 11315 31362 11497 31388
rect 11371 31306 11441 31362
rect 11315 31280 11497 31306
rect 11371 31224 11441 31280
rect 11315 31198 11497 31224
rect 11371 31142 11441 31198
rect 11315 31116 11497 31142
rect 11371 31060 11441 31116
rect 11315 31034 11497 31060
rect 11371 30978 11441 31034
rect 11315 30952 11497 30978
rect 11371 30896 11441 30952
rect 11315 30870 11497 30896
rect 11371 30814 11441 30870
rect 11315 30788 11497 30814
rect 11371 30732 11441 30788
rect 11315 30706 11497 30732
rect 11371 30650 11441 30706
rect 11315 30624 11497 30650
rect 11371 30568 11441 30624
rect 11315 30542 11497 30568
rect 11371 30486 11441 30542
rect 11315 30460 11497 30486
rect 11371 30404 11441 30460
rect 11315 30378 11497 30404
rect 11371 30322 11441 30378
rect 11315 30296 11497 30322
rect 11371 30240 11441 30296
rect 11315 30214 11497 30240
rect 11371 30158 11441 30214
rect 11315 30132 11497 30158
rect 11371 30076 11441 30132
rect 11315 30050 11497 30076
rect 11371 29994 11441 30050
rect 11315 29968 11497 29994
rect 11371 29912 11441 29968
rect 11315 29886 11497 29912
rect 11371 29830 11441 29886
rect 11315 29804 11497 29830
rect 11371 29748 11441 29804
rect 11315 29722 11497 29748
rect 11371 29666 11441 29722
rect 11315 29640 11497 29666
rect 11371 29584 11441 29640
rect 11315 29558 11497 29584
rect 11371 29502 11441 29558
rect 11315 29476 11497 29502
rect 11371 29420 11441 29476
rect 11811 32018 11993 32027
rect 11867 31962 11937 32018
rect 11811 31936 11993 31962
rect 11867 31880 11937 31936
rect 11811 31854 11993 31880
rect 11867 31798 11937 31854
rect 11811 31772 11993 31798
rect 11867 31716 11937 31772
rect 11811 31690 11993 31716
rect 11867 31634 11937 31690
rect 11811 31608 11993 31634
rect 11867 31552 11937 31608
rect 11811 31526 11993 31552
rect 11867 31470 11937 31526
rect 11811 31444 11993 31470
rect 11867 31388 11937 31444
rect 11811 31362 11993 31388
rect 11867 31306 11937 31362
rect 11811 31280 11993 31306
rect 11867 31224 11937 31280
rect 11811 31198 11993 31224
rect 11867 31142 11937 31198
rect 11811 31116 11993 31142
rect 11867 31060 11937 31116
rect 11811 31034 11993 31060
rect 11867 30978 11937 31034
rect 11811 30952 11993 30978
rect 11867 30896 11937 30952
rect 11811 30870 11993 30896
rect 11867 30814 11937 30870
rect 11811 30788 11993 30814
rect 11867 30732 11937 30788
rect 11811 30706 11993 30732
rect 11867 30650 11937 30706
rect 11811 30624 11993 30650
rect 11867 30568 11937 30624
rect 11811 30542 11993 30568
rect 11867 30486 11937 30542
rect 11811 30460 11993 30486
rect 11867 30404 11937 30460
rect 11811 30378 11993 30404
rect 11867 30322 11937 30378
rect 11811 30296 11993 30322
rect 11867 30240 11937 30296
rect 11811 30214 11993 30240
rect 11867 30158 11937 30214
rect 11811 30132 11993 30158
rect 11867 30076 11937 30132
rect 11811 30050 11993 30076
rect 11867 29994 11937 30050
rect 11811 29968 11993 29994
rect 11867 29912 11937 29968
rect 11811 29886 11993 29912
rect 11867 29830 11937 29886
rect 11811 29804 11993 29830
rect 11867 29748 11937 29804
rect 11811 29722 11993 29748
rect 11867 29666 11937 29722
rect 11811 29640 11993 29666
rect 11867 29584 11937 29640
rect 11811 29558 11993 29584
rect 11867 29502 11937 29558
rect 11811 29476 11993 29502
rect 11867 29420 11937 29476
rect 12307 32018 12489 32027
rect 12363 31962 12433 32018
rect 12307 31936 12489 31962
rect 12363 31880 12433 31936
rect 12307 31854 12489 31880
rect 12363 31798 12433 31854
rect 12307 31772 12489 31798
rect 12363 31716 12433 31772
rect 12307 31690 12489 31716
rect 12363 31634 12433 31690
rect 12307 31608 12489 31634
rect 12363 31552 12433 31608
rect 12307 31526 12489 31552
rect 12363 31470 12433 31526
rect 12307 31444 12489 31470
rect 12363 31388 12433 31444
rect 12307 31362 12489 31388
rect 12363 31306 12433 31362
rect 12307 31280 12489 31306
rect 12363 31224 12433 31280
rect 12307 31198 12489 31224
rect 12363 31142 12433 31198
rect 12307 31116 12489 31142
rect 12363 31060 12433 31116
rect 12307 31034 12489 31060
rect 12363 30978 12433 31034
rect 12307 30952 12489 30978
rect 12363 30896 12433 30952
rect 12307 30870 12489 30896
rect 12363 30814 12433 30870
rect 12307 30788 12489 30814
rect 12363 30732 12433 30788
rect 12307 30706 12489 30732
rect 12363 30650 12433 30706
rect 12307 30624 12489 30650
rect 12363 30568 12433 30624
rect 12307 30542 12489 30568
rect 12363 30486 12433 30542
rect 12307 30460 12489 30486
rect 12363 30404 12433 30460
rect 12307 30378 12489 30404
rect 12363 30322 12433 30378
rect 12307 30296 12489 30322
rect 12363 30240 12433 30296
rect 12307 30214 12489 30240
rect 12363 30158 12433 30214
rect 12307 30132 12489 30158
rect 12363 30076 12433 30132
rect 12307 30050 12489 30076
rect 12363 29994 12433 30050
rect 12307 29968 12489 29994
rect 12363 29912 12433 29968
rect 12307 29886 12489 29912
rect 12363 29830 12433 29886
rect 12307 29804 12489 29830
rect 12363 29748 12433 29804
rect 12307 29722 12489 29748
rect 12363 29666 12433 29722
rect 12307 29640 12489 29666
rect 12363 29584 12433 29640
rect 12307 29558 12489 29584
rect 12363 29502 12433 29558
rect 12307 29476 12489 29502
rect 12363 29420 12433 29476
rect 12803 32018 12985 32027
rect 12859 31962 12929 32018
rect 12803 31936 12985 31962
rect 12859 31880 12929 31936
rect 12803 31854 12985 31880
rect 12859 31798 12929 31854
rect 12803 31772 12985 31798
rect 12859 31716 12929 31772
rect 12803 31690 12985 31716
rect 12859 31634 12929 31690
rect 12803 31608 12985 31634
rect 12859 31552 12929 31608
rect 12803 31526 12985 31552
rect 12859 31470 12929 31526
rect 12803 31444 12985 31470
rect 12859 31388 12929 31444
rect 12803 31362 12985 31388
rect 12859 31306 12929 31362
rect 12803 31280 12985 31306
rect 12859 31224 12929 31280
rect 12803 31198 12985 31224
rect 12859 31142 12929 31198
rect 12803 31116 12985 31142
rect 12859 31060 12929 31116
rect 12803 31034 12985 31060
rect 12859 30978 12929 31034
rect 12803 30952 12985 30978
rect 12859 30896 12929 30952
rect 12803 30870 12985 30896
rect 12859 30814 12929 30870
rect 12803 30788 12985 30814
rect 12859 30732 12929 30788
rect 12803 30706 12985 30732
rect 12859 30650 12929 30706
rect 12803 30624 12985 30650
rect 12859 30568 12929 30624
rect 12803 30542 12985 30568
rect 12859 30486 12929 30542
rect 12803 30460 12985 30486
rect 12859 30404 12929 30460
rect 12803 30378 12985 30404
rect 12859 30322 12929 30378
rect 12803 30296 12985 30322
rect 12859 30240 12929 30296
rect 12803 30214 12985 30240
rect 12859 30158 12929 30214
rect 12803 30132 12985 30158
rect 12859 30076 12929 30132
rect 12803 30050 12985 30076
rect 12859 29994 12929 30050
rect 12803 29968 12985 29994
rect 12859 29912 12929 29968
rect 12803 29886 12985 29912
rect 12859 29830 12929 29886
rect 12803 29804 12985 29830
rect 12859 29748 12929 29804
rect 12803 29722 12985 29748
rect 12859 29666 12929 29722
rect 12803 29640 12985 29666
rect 12859 29584 12929 29640
rect 12803 29558 12985 29584
rect 12859 29502 12929 29558
rect 12803 29476 12985 29502
rect 12859 29420 12929 29476
rect 13299 32018 13481 32027
rect 13355 31962 13425 32018
rect 13299 31936 13481 31962
rect 13355 31880 13425 31936
rect 13299 31854 13481 31880
rect 13355 31798 13425 31854
rect 13299 31772 13481 31798
rect 13355 31716 13425 31772
rect 13299 31690 13481 31716
rect 13355 31634 13425 31690
rect 13299 31608 13481 31634
rect 13355 31552 13425 31608
rect 13299 31526 13481 31552
rect 13355 31470 13425 31526
rect 13299 31444 13481 31470
rect 13355 31388 13425 31444
rect 13299 31362 13481 31388
rect 13355 31306 13425 31362
rect 13299 31280 13481 31306
rect 13355 31224 13425 31280
rect 13299 31198 13481 31224
rect 13355 31142 13425 31198
rect 13299 31116 13481 31142
rect 13355 31060 13425 31116
rect 13299 31034 13481 31060
rect 13355 30978 13425 31034
rect 13299 30952 13481 30978
rect 13355 30896 13425 30952
rect 13299 30870 13481 30896
rect 13355 30814 13425 30870
rect 13299 30788 13481 30814
rect 13355 30732 13425 30788
rect 13299 30706 13481 30732
rect 13355 30650 13425 30706
rect 13299 30624 13481 30650
rect 13355 30568 13425 30624
rect 13299 30542 13481 30568
rect 13355 30486 13425 30542
rect 13299 30460 13481 30486
rect 13355 30404 13425 30460
rect 13299 30378 13481 30404
rect 13355 30322 13425 30378
rect 13299 30296 13481 30322
rect 13355 30240 13425 30296
rect 13299 30214 13481 30240
rect 13355 30158 13425 30214
rect 13299 30132 13481 30158
rect 13355 30076 13425 30132
rect 13299 30050 13481 30076
rect 13355 29994 13425 30050
rect 13299 29968 13481 29994
rect 13355 29912 13425 29968
rect 13299 29886 13481 29912
rect 13355 29830 13425 29886
rect 13299 29804 13481 29830
rect 13355 29748 13425 29804
rect 13299 29722 13481 29748
rect 13355 29666 13425 29722
rect 13299 29640 13481 29666
rect 13355 29584 13425 29640
rect 13299 29558 13481 29584
rect 13355 29502 13425 29558
rect 13299 29476 13481 29502
rect 13355 29420 13425 29476
rect 13795 32018 13977 32027
rect 13851 31962 13921 32018
rect 13795 31936 13977 31962
rect 13851 31880 13921 31936
rect 13795 31854 13977 31880
rect 13851 31798 13921 31854
rect 13795 31772 13977 31798
rect 13851 31716 13921 31772
rect 13795 31690 13977 31716
rect 13851 31634 13921 31690
rect 13795 31608 13977 31634
rect 13851 31552 13921 31608
rect 13795 31526 13977 31552
rect 13851 31470 13921 31526
rect 13795 31444 13977 31470
rect 13851 31388 13921 31444
rect 13795 31362 13977 31388
rect 13851 31306 13921 31362
rect 13795 31280 13977 31306
rect 13851 31224 13921 31280
rect 13795 31198 13977 31224
rect 13851 31142 13921 31198
rect 13795 31116 13977 31142
rect 13851 31060 13921 31116
rect 13795 31034 13977 31060
rect 13851 30978 13921 31034
rect 13795 30952 13977 30978
rect 13851 30896 13921 30952
rect 13795 30870 13977 30896
rect 13851 30814 13921 30870
rect 13795 30788 13977 30814
rect 13851 30732 13921 30788
rect 13795 30706 13977 30732
rect 13851 30650 13921 30706
rect 13795 30624 13977 30650
rect 13851 30568 13921 30624
rect 13795 30542 13977 30568
rect 13851 30486 13921 30542
rect 13795 30460 13977 30486
rect 13851 30404 13921 30460
rect 13795 30378 13977 30404
rect 13851 30322 13921 30378
rect 13795 30296 13977 30322
rect 13851 30240 13921 30296
rect 13795 30214 13977 30240
rect 13851 30158 13921 30214
rect 13795 30132 13977 30158
rect 13851 30076 13921 30132
rect 13795 30050 13977 30076
rect 13851 29994 13921 30050
rect 13795 29968 13977 29994
rect 13851 29912 13921 29968
rect 13795 29886 13977 29912
rect 13851 29830 13921 29886
rect 13795 29804 13977 29830
rect 13851 29748 13921 29804
rect 13795 29722 13977 29748
rect 13851 29666 13921 29722
rect 13795 29640 13977 29666
rect 13851 29584 13921 29640
rect 13795 29558 13977 29584
rect 13851 29502 13921 29558
rect 13795 29476 13977 29502
rect 13851 29420 13921 29476
rect 14315 31985 14347 32041
rect 14403 31985 14435 32041
rect 14491 31985 14523 32041
rect 14579 31985 14611 32041
rect 14259 31961 14667 31985
rect 14315 31905 14347 31961
rect 14403 31905 14435 31961
rect 14491 31905 14523 31961
rect 14579 31905 14611 31961
rect 14259 31881 14667 31905
rect 14315 31825 14347 31881
rect 14403 31825 14435 31881
rect 14491 31825 14523 31881
rect 14579 31825 14611 31881
rect 14259 31801 14667 31825
rect 14315 31745 14347 31801
rect 14403 31745 14435 31801
rect 14491 31745 14523 31801
rect 14579 31745 14611 31801
rect 14259 31721 14667 31745
rect 14315 31665 14347 31721
rect 14403 31665 14435 31721
rect 14491 31665 14523 31721
rect 14579 31665 14611 31721
rect 14259 31641 14667 31665
rect 14315 31585 14347 31641
rect 14403 31585 14435 31641
rect 14491 31585 14523 31641
rect 14579 31585 14611 31641
rect 14259 31561 14667 31585
rect 14315 31505 14347 31561
rect 14403 31505 14435 31561
rect 14491 31505 14523 31561
rect 14579 31505 14611 31561
rect 14259 31481 14667 31505
rect 14315 31425 14347 31481
rect 14403 31425 14435 31481
rect 14491 31425 14523 31481
rect 14579 31425 14611 31481
rect 14259 31400 14667 31425
rect 14315 31344 14347 31400
rect 14403 31344 14435 31400
rect 14491 31344 14523 31400
rect 14579 31344 14611 31400
rect 14259 31319 14667 31344
rect 14315 31263 14347 31319
rect 14403 31263 14435 31319
rect 14491 31263 14523 31319
rect 14579 31263 14611 31319
rect 14259 31238 14667 31263
rect 14315 31182 14347 31238
rect 14403 31182 14435 31238
rect 14491 31182 14523 31238
rect 14579 31182 14611 31238
rect 14259 31157 14667 31182
rect 14315 31101 14347 31157
rect 14403 31101 14435 31157
rect 14491 31101 14523 31157
rect 14579 31101 14611 31157
rect 14259 31076 14667 31101
rect 14315 31020 14347 31076
rect 14403 31020 14435 31076
rect 14491 31020 14523 31076
rect 14579 31020 14611 31076
rect 14259 30995 14667 31020
rect 14315 30939 14347 30995
rect 14403 30939 14435 30995
rect 14491 30939 14523 30995
rect 14579 30939 14611 30995
rect 14259 30914 14667 30939
rect 14315 30858 14347 30914
rect 14403 30858 14435 30914
rect 14491 30858 14523 30914
rect 14579 30858 14611 30914
rect 14259 30833 14667 30858
rect 14315 30777 14347 30833
rect 14403 30777 14435 30833
rect 14491 30777 14523 30833
rect 14579 30777 14611 30833
rect 14259 30752 14667 30777
rect 14315 30696 14347 30752
rect 14403 30696 14435 30752
rect 14491 30696 14523 30752
rect 14579 30696 14611 30752
rect 14259 30671 14667 30696
rect 14315 30615 14347 30671
rect 14403 30615 14435 30671
rect 14491 30615 14523 30671
rect 14579 30615 14611 30671
rect 14259 30590 14667 30615
rect 14315 30534 14347 30590
rect 14403 30534 14435 30590
rect 14491 30534 14523 30590
rect 14579 30534 14611 30590
rect 14259 30509 14667 30534
rect 14315 30453 14347 30509
rect 14403 30453 14435 30509
rect 14491 30453 14523 30509
rect 14579 30453 14611 30509
rect 14259 30428 14667 30453
rect 14315 30372 14347 30428
rect 14403 30372 14435 30428
rect 14491 30372 14523 30428
rect 14579 30372 14611 30428
rect 14259 30347 14667 30372
rect 14315 30291 14347 30347
rect 14403 30291 14435 30347
rect 14491 30291 14523 30347
rect 14579 30291 14611 30347
rect 14259 30266 14667 30291
rect 14315 30210 14347 30266
rect 14403 30210 14435 30266
rect 14491 30210 14523 30266
rect 14579 30210 14611 30266
rect 14259 30185 14667 30210
rect 14315 30129 14347 30185
rect 14403 30129 14435 30185
rect 14491 30129 14523 30185
rect 14579 30129 14611 30185
rect 14259 30104 14667 30129
rect 14315 30048 14347 30104
rect 14403 30048 14435 30104
rect 14491 30048 14523 30104
rect 14579 30048 14611 30104
rect 14259 30023 14667 30048
rect 14315 29967 14347 30023
rect 14403 29967 14435 30023
rect 14491 29967 14523 30023
rect 14579 29967 14611 30023
rect 14259 29942 14667 29967
rect 14315 29886 14347 29942
rect 14403 29886 14435 29942
rect 14491 29886 14523 29942
rect 14579 29886 14611 29942
rect 14259 29861 14667 29886
rect 14315 29805 14347 29861
rect 14403 29805 14435 29861
rect 14491 29805 14523 29861
rect 14579 29805 14611 29861
rect 14259 29780 14667 29805
rect 14315 29724 14347 29780
rect 14403 29724 14435 29780
rect 14491 29724 14523 29780
rect 14579 29724 14611 29780
rect 14259 29699 14667 29724
rect 14315 29643 14347 29699
rect 14403 29643 14435 29699
rect 14491 29643 14523 29699
rect 14579 29643 14611 29699
rect 14259 29618 14667 29643
rect 14315 29562 14347 29618
rect 14403 29562 14435 29618
rect 14491 29562 14523 29618
rect 14579 29562 14611 29618
rect 14259 29537 14667 29562
rect 14315 29481 14347 29537
rect 14403 29481 14435 29537
rect 14491 29481 14523 29537
rect 14579 29481 14611 29537
rect 14259 29456 14667 29481
rect 862 29411 1052 29420
rect 1890 29411 2080 29420
rect 2386 29411 2576 29420
rect 2882 29411 3072 29420
rect 3378 29411 3568 29420
rect 3874 29411 4064 29420
rect 4370 29411 4560 29420
rect 4866 29411 5056 29420
rect 5362 29411 5552 29420
rect 5858 29411 6048 29420
rect 6354 29411 6544 29420
rect 6850 29411 7040 29420
rect 7346 29411 7536 29420
rect 7842 29411 8032 29420
rect 8338 29411 8528 29420
rect 8834 29411 9024 29420
rect 9330 29411 9520 29420
rect 9826 29411 10016 29420
rect 10322 29411 10512 29420
rect 10818 29411 11008 29420
rect 11314 29411 11504 29420
rect 11810 29411 12000 29420
rect 12306 29411 12496 29420
rect 12802 29411 12992 29420
rect 13298 29411 13488 29420
rect 13794 29411 13984 29420
rect 14315 29400 14347 29456
rect 14403 29400 14435 29456
rect 14491 29400 14523 29456
rect 14579 29400 14611 29456
rect 14259 29375 14667 29400
rect 14315 29319 14347 29375
rect 14403 29319 14435 29375
rect 14491 29319 14523 29375
rect 14579 29319 14611 29375
rect 14259 29294 14667 29319
rect 14315 29238 14347 29294
rect 14403 29238 14435 29294
rect 14491 29238 14523 29294
rect 14579 29238 14611 29294
rect 14259 29213 14667 29238
rect 14315 29157 14347 29213
rect 14403 29157 14435 29213
rect 14491 29157 14523 29213
rect 14579 29157 14611 29213
rect 14259 29132 14667 29157
rect 14315 29076 14347 29132
rect 14403 29076 14435 29132
rect 14491 29076 14523 29132
rect 14579 29076 14611 29132
rect 14259 29067 14667 29076
rect 575 28632 1189 28633
rect 575 28596 581 28632
rect 633 28596 650 28632
rect 702 28596 719 28632
rect 771 28596 788 28632
rect 575 28540 579 28596
rect 635 28580 650 28596
rect 771 28580 775 28596
rect 840 28580 857 28632
rect 909 28580 926 28632
rect 978 28580 995 28632
rect 1047 28580 1063 28632
rect 1115 28580 1131 28632
rect 1183 28580 1189 28632
rect 635 28558 677 28580
rect 733 28558 775 28580
rect 831 28558 1189 28580
rect 635 28540 650 28558
rect 771 28540 775 28558
rect 575 28515 581 28540
rect 633 28515 650 28540
rect 702 28515 719 28540
rect 771 28515 788 28540
rect 575 28459 579 28515
rect 635 28506 650 28515
rect 771 28506 775 28515
rect 840 28506 857 28558
rect 909 28506 926 28558
rect 978 28506 995 28558
rect 1047 28506 1063 28558
rect 1115 28506 1131 28558
rect 1183 28506 1189 28558
rect 635 28484 677 28506
rect 733 28484 775 28506
rect 831 28484 1189 28506
rect 635 28459 650 28484
rect 771 28459 775 28484
rect 575 28434 581 28459
rect 633 28434 650 28459
rect 702 28434 719 28459
rect 771 28434 788 28459
rect 575 28378 579 28434
rect 635 28432 650 28434
rect 771 28432 775 28434
rect 840 28432 857 28484
rect 909 28432 926 28484
rect 978 28432 995 28484
rect 1047 28432 1063 28484
rect 1115 28432 1131 28484
rect 1183 28432 1189 28484
rect 635 28378 677 28432
rect 733 28378 775 28432
rect 831 28378 1189 28432
rect 575 28353 1189 28378
rect 575 28297 579 28353
rect 635 28297 677 28353
rect 733 28297 775 28353
rect 831 28297 1189 28353
rect 575 28272 1189 28297
rect 575 28216 579 28272
rect 635 28216 677 28272
rect 733 28216 775 28272
rect 831 28216 1189 28272
rect 575 28191 1189 28216
rect 575 28135 579 28191
rect 635 28135 677 28191
rect 733 28135 775 28191
rect 831 28135 1189 28191
rect 575 28110 1189 28135
rect 3472 28581 3478 28633
rect 3530 28620 3546 28633
rect 3598 28581 3614 28633
rect 3666 28581 3682 28633
rect 3734 28581 3750 28633
rect 3802 28581 3818 28633
rect 3870 28581 3886 28633
rect 3938 28581 3954 28633
rect 4006 28581 4021 28633
rect 4073 28581 4088 28633
rect 4140 28581 4155 28633
rect 4207 28581 4222 28633
rect 4274 28581 4289 28633
rect 4341 28581 4356 28633
rect 4408 28581 4423 28633
rect 4475 28620 4490 28633
rect 4475 28581 4485 28620
rect 4542 28581 4557 28633
rect 4609 28581 4615 28633
rect 3472 28564 3494 28581
rect 3550 28564 4485 28581
rect 4541 28564 4615 28581
rect 3472 28559 4615 28564
rect 3472 28507 3478 28559
rect 3530 28507 3546 28559
rect 3598 28507 3614 28559
rect 3666 28507 3682 28559
rect 3734 28507 3750 28559
rect 3802 28507 3818 28559
rect 3870 28507 3886 28559
rect 3938 28507 3954 28559
rect 4006 28507 4021 28559
rect 4073 28507 4088 28559
rect 4140 28507 4155 28559
rect 4207 28507 4222 28559
rect 4274 28507 4289 28559
rect 4341 28507 4356 28559
rect 4408 28507 4423 28559
rect 4475 28507 4490 28559
rect 4542 28507 4557 28559
rect 4609 28507 4615 28559
rect 3472 28485 4615 28507
rect 3472 28433 3478 28485
rect 3530 28451 3546 28485
rect 3598 28433 3614 28485
rect 3666 28433 3682 28485
rect 3734 28433 3750 28485
rect 3802 28433 3818 28485
rect 3870 28433 3886 28485
rect 3938 28433 3954 28485
rect 4006 28433 4021 28485
rect 4073 28433 4088 28485
rect 4140 28433 4155 28485
rect 4207 28433 4222 28485
rect 4274 28433 4289 28485
rect 4341 28433 4356 28485
rect 4408 28433 4423 28485
rect 4475 28451 4490 28485
rect 4475 28433 4485 28451
rect 4542 28433 4557 28485
rect 4609 28433 4615 28485
rect 3472 28395 3494 28433
rect 3550 28395 4485 28433
rect 4541 28395 4615 28433
rect 3472 28282 4615 28395
rect 3472 28226 3494 28282
rect 3550 28226 4485 28282
rect 4541 28226 4615 28282
rect 575 28054 579 28110
rect 635 28054 677 28110
rect 733 28054 775 28110
rect 831 28054 1189 28110
rect 575 28029 1189 28054
rect 575 27973 579 28029
rect 635 27973 677 28029
rect 733 27973 775 28029
rect 831 27973 1189 28029
rect 575 27948 1189 27973
rect 575 27892 579 27948
rect 635 27892 677 27948
rect 733 27892 775 27948
rect 831 27892 1189 27948
rect 575 27867 1189 27892
rect 575 27811 579 27867
rect 635 27811 677 27867
rect 733 27811 775 27867
rect 831 27811 1189 27867
rect 575 27786 1189 27811
rect 575 27730 579 27786
rect 635 27730 677 27786
rect 733 27730 775 27786
rect 831 27730 1189 27786
rect 575 27705 1189 27730
rect 575 27649 579 27705
rect 635 27649 677 27705
rect 733 27649 775 27705
rect 831 27649 1189 27705
rect 575 27624 1189 27649
rect 575 27568 579 27624
rect 635 27568 677 27624
rect 733 27568 775 27624
rect 831 27568 1189 27624
rect 575 27543 1189 27568
rect 575 27487 579 27543
rect 635 27487 677 27543
rect 733 27487 775 27543
rect 831 27487 1189 27543
rect 575 27462 1189 27487
rect 575 27406 579 27462
rect 635 27406 677 27462
rect 733 27406 775 27462
rect 831 27406 1189 27462
rect 575 27381 1189 27406
rect 575 27325 579 27381
rect 635 27325 677 27381
rect 733 27325 775 27381
rect 831 27325 1189 27381
rect 575 27300 1189 27325
rect 575 27244 579 27300
rect 635 27244 677 27300
rect 733 27244 775 27300
rect 831 27244 1189 27300
rect 575 27219 1189 27244
rect 575 27163 579 27219
rect 635 27163 677 27219
rect 733 27163 775 27219
rect 831 27163 1189 27219
rect 575 27138 1189 27163
rect 575 27082 579 27138
rect 635 27082 677 27138
rect 733 27082 775 27138
rect 831 27082 1189 27138
rect 575 27057 1189 27082
rect 575 27001 579 27057
rect 635 27001 677 27057
rect 733 27001 775 27057
rect 831 27001 1189 27057
rect 575 26976 1189 27001
rect 575 26920 579 26976
rect 635 26920 677 26976
rect 733 26920 775 26976
rect 831 26920 1189 26976
rect 575 26894 1189 26920
rect 575 26838 579 26894
rect 635 26838 677 26894
rect 733 26838 775 26894
rect 831 26838 1189 26894
rect 575 26812 1189 26838
rect 575 26756 579 26812
rect 635 26756 677 26812
rect 733 26756 775 26812
rect 831 26756 1189 26812
rect 575 26730 1189 26756
tri 201 26352 575 26726 se
rect 575 26674 579 26730
rect 635 26674 677 26730
rect 733 26674 775 26730
rect 831 26674 1189 26730
rect 575 26648 1189 26674
rect 575 26592 579 26648
rect 635 26592 677 26648
rect 733 26592 775 26648
rect 831 26592 1189 26648
rect 575 26566 1189 26592
rect 575 26510 579 26566
rect 635 26510 677 26566
rect 733 26510 775 26566
rect 831 26510 1189 26566
rect 575 26484 1189 26510
rect 575 26428 579 26484
rect 635 26428 677 26484
rect 733 26428 775 26484
rect 831 26472 1189 26484
rect 831 26428 1069 26472
rect 575 26352 1069 26428
tri 1069 26352 1189 26472 nw
rect 1297 28124 2039 28129
rect 1297 28072 1303 28124
rect 1355 28072 1371 28124
rect 1423 28072 1439 28124
rect 1491 28072 1507 28124
rect 1559 28072 1575 28124
rect 1627 28072 1643 28124
rect 1695 28072 1711 28124
rect 1763 28072 1779 28124
rect 1831 28072 1847 28124
rect 1899 28072 1914 28124
rect 1966 28072 1981 28124
rect 2033 28072 2039 28124
rect 1297 28058 2039 28072
rect 1297 28006 1303 28058
rect 1355 28006 1371 28058
rect 1423 28006 1439 28058
rect 1491 28006 1507 28058
rect 1559 28006 1575 28058
rect 1627 28006 1643 28058
rect 1695 28006 1711 28058
rect 1763 28006 1779 28058
rect 1831 28006 1847 28058
rect 1899 28006 1914 28058
rect 1966 28006 1981 28058
rect 2033 28006 2039 28058
rect 1297 27992 2039 28006
rect 1297 27940 1303 27992
rect 1355 27940 1371 27992
rect 1423 27940 1439 27992
rect 1491 27940 1507 27992
rect 1559 27940 1575 27992
rect 1627 27940 1643 27992
rect 1695 27940 1711 27992
rect 1763 27940 1779 27992
rect 1831 27940 1847 27992
rect 1899 27940 1914 27992
rect 1966 27940 1981 27992
rect 2033 27940 2039 27992
rect 1297 27926 2039 27940
rect 1297 27874 1303 27926
rect 1355 27874 1371 27926
rect 1423 27874 1439 27926
rect 1491 27874 1507 27926
rect 1559 27874 1575 27926
rect 1627 27874 1643 27926
rect 1695 27874 1711 27926
rect 1763 27874 1779 27926
rect 1831 27874 1847 27926
rect 1899 27874 1914 27926
rect 1966 27874 1981 27926
rect 2033 27874 2039 27926
rect 1297 27860 2039 27874
rect 1297 27808 1303 27860
rect 1355 27808 1371 27860
rect 1423 27808 1439 27860
rect 1491 27808 1507 27860
rect 1559 27808 1575 27860
rect 1627 27808 1643 27860
rect 1695 27808 1711 27860
rect 1763 27808 1779 27860
rect 1831 27808 1847 27860
rect 1899 27808 1914 27860
rect 1966 27808 1981 27860
rect 2033 27808 2039 27860
rect 1297 27794 2039 27808
rect 1297 27742 1303 27794
rect 1355 27742 1371 27794
rect 1423 27742 1439 27794
rect 1491 27742 1507 27794
rect 1559 27742 1575 27794
rect 1627 27742 1643 27794
rect 1695 27742 1711 27794
rect 1763 27742 1779 27794
rect 1831 27742 1847 27794
rect 1899 27742 1914 27794
rect 1966 27742 1981 27794
rect 2033 27742 2039 27794
rect 1297 27728 2039 27742
rect 1297 27676 1303 27728
rect 1355 27676 1371 27728
rect 1423 27676 1439 27728
rect 1491 27676 1507 27728
rect 1559 27676 1575 27728
rect 1627 27676 1643 27728
rect 1695 27676 1711 27728
rect 1763 27676 1779 27728
rect 1831 27676 1847 27728
rect 1899 27676 1914 27728
rect 1966 27676 1981 27728
rect 2033 27676 2039 27728
tri 164 26315 201 26352 se
rect 201 26343 904 26352
rect 201 26315 242 26343
rect 164 26287 242 26315
rect 298 26287 334 26343
rect 390 26287 426 26343
rect 482 26287 518 26343
rect 574 26287 610 26343
rect 666 26287 702 26343
rect 758 26287 904 26343
rect 164 26263 904 26287
rect 164 26207 242 26263
rect 298 26207 334 26263
rect 390 26207 426 26263
rect 482 26207 518 26263
rect 574 26207 610 26263
rect 666 26207 702 26263
rect 758 26207 904 26263
rect 164 26187 904 26207
tri 904 26187 1069 26352 nw
rect 164 26183 898 26187
rect 164 26127 242 26183
rect 298 26127 334 26183
rect 390 26127 426 26183
rect 482 26127 518 26183
rect 574 26127 610 26183
rect 666 26127 702 26183
rect 758 26181 898 26183
tri 898 26181 904 26187 nw
rect 758 26129 846 26181
tri 846 26129 898 26181 nw
rect 758 26127 828 26129
rect 164 26111 828 26127
tri 828 26111 846 26129 nw
rect 164 26103 778 26111
rect 164 26047 242 26103
rect 298 26047 334 26103
rect 390 26047 426 26103
rect 482 26047 518 26103
rect 574 26047 610 26103
rect 666 26047 702 26103
rect 758 26047 778 26103
tri 778 26061 828 26111 nw
rect 164 26023 778 26047
rect 164 25967 242 26023
rect 298 25967 334 26023
rect 390 25967 426 26023
rect 482 25967 518 26023
rect 574 25967 610 26023
rect 666 25967 702 26023
rect 758 25967 778 26023
rect 164 25943 778 25967
rect 164 25887 242 25943
rect 298 25887 334 25943
rect 390 25887 426 25943
rect 482 25887 518 25943
rect 574 25887 610 25943
rect 666 25887 702 25943
rect 758 25887 778 25943
rect 164 25863 778 25887
rect 164 25807 242 25863
rect 298 25807 334 25863
rect 390 25807 426 25863
rect 482 25807 518 25863
rect 574 25807 610 25863
rect 666 25807 702 25863
rect 758 25807 778 25863
rect 164 25783 778 25807
rect 164 25727 242 25783
rect 298 25727 334 25783
rect 390 25727 426 25783
rect 482 25727 518 25783
rect 574 25727 610 25783
rect 666 25727 702 25783
rect 758 25727 778 25783
rect 164 25703 778 25727
rect 164 25647 242 25703
rect 298 25647 334 25703
rect 390 25647 426 25703
rect 482 25647 518 25703
rect 574 25647 610 25703
rect 666 25647 702 25703
rect 758 25647 778 25703
rect 164 25623 778 25647
rect 164 25567 242 25623
rect 298 25567 334 25623
rect 390 25567 426 25623
rect 482 25567 518 25623
rect 574 25567 610 25623
rect 666 25567 702 25623
rect 758 25567 778 25623
rect 164 25543 778 25567
rect 164 25487 242 25543
rect 298 25487 334 25543
rect 390 25487 426 25543
rect 482 25487 518 25543
rect 574 25487 610 25543
rect 666 25487 702 25543
rect 758 25487 778 25543
rect 164 25463 778 25487
rect 164 25407 242 25463
rect 298 25407 334 25463
rect 390 25407 426 25463
rect 482 25407 518 25463
rect 574 25407 610 25463
rect 666 25407 702 25463
rect 758 25407 778 25463
rect 164 25383 778 25407
rect 164 25327 242 25383
rect 298 25327 334 25383
rect 390 25327 426 25383
rect 482 25327 518 25383
rect 574 25327 610 25383
rect 666 25327 702 25383
rect 758 25327 778 25383
rect 164 25303 778 25327
rect 164 25247 242 25303
rect 298 25247 334 25303
rect 390 25247 426 25303
rect 482 25247 518 25303
rect 574 25247 610 25303
rect 666 25247 702 25303
rect 758 25247 778 25303
rect 164 25223 778 25247
rect 164 25167 242 25223
rect 298 25167 334 25223
rect 390 25167 426 25223
rect 482 25167 518 25223
rect 574 25167 610 25223
rect 666 25167 702 25223
rect 758 25167 778 25223
rect 164 25143 778 25167
rect 164 25087 242 25143
rect 298 25087 334 25143
rect 390 25087 426 25143
rect 482 25087 518 25143
rect 574 25087 610 25143
rect 666 25087 702 25143
rect 758 25087 778 25143
rect 164 25063 778 25087
rect 164 25007 242 25063
rect 298 25007 334 25063
rect 390 25007 426 25063
rect 482 25007 518 25063
rect 574 25007 610 25063
rect 666 25007 702 25063
rect 758 25007 778 25063
rect 164 24983 778 25007
rect 164 24927 242 24983
rect 298 24927 334 24983
rect 390 24927 426 24983
rect 482 24927 518 24983
rect 574 24927 610 24983
rect 666 24927 702 24983
rect 758 24927 778 24983
rect 164 24903 778 24927
rect 164 24847 242 24903
rect 298 24847 334 24903
rect 390 24847 426 24903
rect 482 24847 518 24903
rect 574 24847 610 24903
rect 666 24847 702 24903
rect 758 24847 778 24903
rect 164 24823 778 24847
rect 164 24767 242 24823
rect 298 24767 334 24823
rect 390 24767 426 24823
rect 482 24767 518 24823
rect 574 24767 610 24823
rect 666 24767 702 24823
rect 758 24767 778 24823
rect 164 24743 778 24767
rect 164 24687 242 24743
rect 298 24687 334 24743
rect 390 24687 426 24743
rect 482 24687 518 24743
rect 574 24687 610 24743
rect 666 24687 702 24743
rect 758 24687 778 24743
rect 164 24663 778 24687
rect 164 24607 242 24663
rect 298 24607 334 24663
rect 390 24607 426 24663
rect 482 24607 518 24663
rect 574 24607 610 24663
rect 666 24607 702 24663
rect 758 24607 778 24663
rect 164 24583 778 24607
rect 164 24527 242 24583
rect 298 24527 334 24583
rect 390 24527 426 24583
rect 482 24527 518 24583
rect 574 24527 610 24583
rect 666 24527 702 24583
rect 758 24527 778 24583
rect 164 24503 778 24527
rect 164 24447 242 24503
rect 298 24447 334 24503
rect 390 24447 426 24503
rect 482 24447 518 24503
rect 574 24447 610 24503
rect 666 24447 702 24503
rect 758 24447 778 24503
rect 1297 25037 2039 27676
rect 3472 28113 4615 28226
rect 3472 28112 4485 28113
rect 3472 28056 3494 28112
rect 3550 28057 4485 28112
rect 4541 28057 4615 28113
rect 3550 28056 4615 28057
rect 3472 27944 4615 28056
rect 3472 27942 4485 27944
rect 3472 27886 3494 27942
rect 3550 27888 4485 27942
rect 4541 27888 4615 27944
rect 3550 27886 4615 27888
rect 3472 27774 4615 27886
rect 3472 27772 4485 27774
rect 3472 27716 3494 27772
rect 3550 27718 4485 27772
rect 4541 27718 4615 27774
rect 3550 27716 4615 27718
rect 3472 27604 4615 27716
rect 3472 27602 4485 27604
rect 3472 27546 3494 27602
rect 3550 27548 4485 27602
rect 4541 27548 4615 27604
rect 3550 27546 4615 27548
rect 3472 27434 4615 27546
rect 3472 27432 4485 27434
rect 3472 27376 3494 27432
rect 3550 27378 4485 27432
rect 4541 27378 4615 27434
rect 3550 27376 4615 27378
rect 3472 27369 4615 27376
rect 3472 27317 3478 27369
rect 3530 27317 3546 27369
rect 3598 27317 3614 27369
rect 3666 27317 3682 27369
rect 3734 27317 3750 27369
rect 3802 27317 3818 27369
rect 3870 27317 3886 27369
rect 3938 27317 3954 27369
rect 4006 27317 4021 27369
rect 4073 27317 4088 27369
rect 4140 27317 4155 27369
rect 4207 27317 4222 27369
rect 4274 27317 4289 27369
rect 4341 27317 4356 27369
rect 4408 27317 4423 27369
rect 4475 27317 4490 27369
rect 4542 27317 4557 27369
rect 4609 27317 4615 27369
rect 3472 27264 4615 27317
rect 3472 27262 4485 27264
rect 3472 27243 3494 27262
rect 3550 27243 4485 27262
rect 4541 27243 4615 27264
rect 3472 27191 3478 27243
rect 3530 27191 3546 27206
rect 3598 27191 3614 27243
rect 3666 27191 3682 27243
rect 3734 27191 3750 27243
rect 3802 27191 3818 27243
rect 3870 27191 3886 27243
rect 3938 27191 3954 27243
rect 4006 27191 4021 27243
rect 4073 27191 4088 27243
rect 4140 27191 4155 27243
rect 4207 27191 4222 27243
rect 4274 27191 4289 27243
rect 4341 27191 4356 27243
rect 4408 27191 4423 27243
rect 4475 27208 4485 27243
rect 4475 27191 4490 27208
rect 4542 27191 4557 27243
rect 4609 27191 4615 27243
rect 5455 28581 5461 28633
rect 5513 28620 5528 28633
rect 5580 28581 5595 28633
rect 5647 28581 5662 28633
rect 5714 28581 5729 28633
rect 5781 28581 5796 28633
rect 5848 28581 5863 28633
rect 5915 28581 5930 28633
rect 5982 28581 5997 28633
rect 6049 28581 6064 28633
rect 6116 28581 6132 28633
rect 6184 28581 6200 28633
rect 6252 28581 6268 28633
rect 6320 28581 6336 28633
rect 6388 28581 6404 28633
rect 6456 28620 6472 28633
rect 6524 28620 6540 28633
rect 6456 28581 6469 28620
rect 6525 28581 6540 28620
rect 6592 28581 6599 28633
rect 5455 28564 5477 28581
rect 5533 28564 6469 28581
rect 6525 28564 6599 28581
rect 5455 28559 6599 28564
rect 5455 28507 5461 28559
rect 5513 28507 5528 28559
rect 5580 28507 5595 28559
rect 5647 28507 5662 28559
rect 5714 28507 5729 28559
rect 5781 28507 5796 28559
rect 5848 28507 5863 28559
rect 5915 28507 5930 28559
rect 5982 28507 5997 28559
rect 6049 28507 6064 28559
rect 6116 28507 6132 28559
rect 6184 28507 6200 28559
rect 6252 28507 6268 28559
rect 6320 28507 6336 28559
rect 6388 28507 6404 28559
rect 6456 28507 6472 28559
rect 6524 28507 6540 28559
rect 6592 28507 6599 28559
rect 5455 28485 6599 28507
rect 5455 28433 5461 28485
rect 5513 28453 5528 28485
rect 5580 28433 5595 28485
rect 5647 28433 5662 28485
rect 5714 28433 5729 28485
rect 5781 28433 5796 28485
rect 5848 28433 5863 28485
rect 5915 28433 5930 28485
rect 5982 28433 5997 28485
rect 6049 28433 6064 28485
rect 6116 28433 6132 28485
rect 6184 28433 6200 28485
rect 6252 28433 6268 28485
rect 6320 28433 6336 28485
rect 6388 28433 6404 28485
rect 6456 28453 6472 28485
rect 6524 28453 6540 28485
rect 6456 28433 6469 28453
rect 6525 28433 6540 28453
rect 6592 28433 6599 28485
rect 5455 28397 5477 28433
rect 5533 28397 6469 28433
rect 6525 28397 6599 28433
rect 5455 28286 6599 28397
rect 5455 28230 5477 28286
rect 5533 28230 6469 28286
rect 6525 28230 6599 28286
rect 5455 28119 6599 28230
rect 5455 28063 5477 28119
rect 5533 28063 6469 28119
rect 6525 28063 6599 28119
rect 5455 27952 6599 28063
rect 5455 27896 5477 27952
rect 5533 27896 6469 27952
rect 6525 27896 6599 27952
rect 5455 27785 6599 27896
rect 5455 27729 5477 27785
rect 5533 27729 6469 27785
rect 6525 27729 6599 27785
rect 5455 27618 6599 27729
rect 5455 27562 5477 27618
rect 5533 27562 6469 27618
rect 6525 27562 6599 27618
rect 5455 27451 6599 27562
rect 5455 27395 5477 27451
rect 5533 27395 6469 27451
rect 6525 27395 6599 27451
rect 5455 27369 6599 27395
rect 5455 27317 5461 27369
rect 5513 27317 5529 27369
rect 5581 27317 5597 27369
rect 5649 27317 5665 27369
rect 5717 27317 5733 27369
rect 5785 27317 5801 27369
rect 5853 27317 5869 27369
rect 5921 27317 5937 27369
rect 5989 27317 6004 27369
rect 6056 27317 6071 27369
rect 6123 27317 6138 27369
rect 6190 27317 6205 27369
rect 6257 27317 6272 27369
rect 6324 27317 6339 27369
rect 6391 27317 6406 27369
rect 6458 27317 6473 27369
rect 6525 27317 6540 27369
rect 6592 27317 6599 27369
rect 5455 27283 6599 27317
rect 5455 27243 5477 27283
rect 5533 27243 6469 27283
rect 6525 27243 6599 27283
rect 5455 27191 5461 27243
rect 5513 27191 5529 27227
rect 5581 27191 5597 27243
rect 5649 27191 5665 27243
rect 5717 27191 5733 27243
rect 5785 27191 5801 27243
rect 5853 27191 5869 27243
rect 5921 27191 5937 27243
rect 5989 27191 6004 27243
rect 6056 27191 6071 27243
rect 6123 27191 6138 27243
rect 6190 27191 6205 27243
rect 6257 27191 6272 27243
rect 6324 27191 6339 27243
rect 6391 27191 6406 27243
rect 6458 27227 6469 27243
rect 6458 27191 6473 27227
rect 6525 27191 6540 27243
rect 6592 27191 6599 27243
rect 7439 28581 7445 28633
rect 7497 28620 7512 28633
rect 7564 28581 7579 28633
rect 7631 28581 7646 28633
rect 7698 28581 7713 28633
rect 7765 28581 7780 28633
rect 7832 28581 7847 28633
rect 7899 28581 7914 28633
rect 7966 28581 7981 28633
rect 8033 28581 8048 28633
rect 8100 28581 8116 28633
rect 8168 28581 8184 28633
rect 8236 28581 8252 28633
rect 8304 28581 8320 28633
rect 8372 28581 8388 28633
rect 8440 28620 8456 28633
rect 8508 28620 8524 28633
rect 8440 28581 8453 28620
rect 8509 28581 8524 28620
rect 8576 28581 8582 28633
rect 7439 28564 7461 28581
rect 7517 28564 8453 28581
rect 8509 28564 8582 28581
rect 7439 28559 8582 28564
rect 7439 28507 7445 28559
rect 7497 28507 7512 28559
rect 7564 28507 7579 28559
rect 7631 28507 7646 28559
rect 7698 28507 7713 28559
rect 7765 28507 7780 28559
rect 7832 28507 7847 28559
rect 7899 28507 7914 28559
rect 7966 28507 7981 28559
rect 8033 28507 8048 28559
rect 8100 28507 8116 28559
rect 8168 28507 8184 28559
rect 8236 28507 8252 28559
rect 8304 28507 8320 28559
rect 8372 28507 8388 28559
rect 8440 28507 8456 28559
rect 8508 28507 8524 28559
rect 8576 28507 8582 28559
rect 7439 28485 8582 28507
rect 7439 28433 7445 28485
rect 7497 28453 7512 28485
rect 7564 28433 7579 28485
rect 7631 28433 7646 28485
rect 7698 28433 7713 28485
rect 7765 28433 7780 28485
rect 7832 28433 7847 28485
rect 7899 28433 7914 28485
rect 7966 28433 7981 28485
rect 8033 28433 8048 28485
rect 8100 28433 8116 28485
rect 8168 28433 8184 28485
rect 8236 28433 8252 28485
rect 8304 28433 8320 28485
rect 8372 28433 8388 28485
rect 8440 28453 8456 28485
rect 8508 28453 8524 28485
rect 8440 28433 8453 28453
rect 8509 28433 8524 28453
rect 8576 28433 8582 28485
rect 7439 28397 7461 28433
rect 7517 28397 8453 28433
rect 8509 28397 8582 28433
rect 7439 28286 8582 28397
rect 7439 28230 7461 28286
rect 7517 28230 8453 28286
rect 8509 28230 8582 28286
rect 7439 28119 8582 28230
rect 7439 28063 7461 28119
rect 7517 28063 8453 28119
rect 8509 28063 8582 28119
rect 7439 27952 8582 28063
rect 7439 27896 7461 27952
rect 7517 27896 8453 27952
rect 8509 27896 8582 27952
rect 7439 27785 8582 27896
rect 7439 27729 7461 27785
rect 7517 27729 8453 27785
rect 8509 27729 8582 27785
rect 7439 27618 8582 27729
rect 7439 27562 7461 27618
rect 7517 27562 8453 27618
rect 8509 27562 8582 27618
rect 7439 27451 8582 27562
rect 7439 27395 7461 27451
rect 7517 27395 8453 27451
rect 8509 27395 8582 27451
rect 7439 27369 8582 27395
rect 7439 27317 7445 27369
rect 7497 27317 7513 27369
rect 7565 27317 7581 27369
rect 7633 27317 7649 27369
rect 7701 27317 7717 27369
rect 7769 27317 7785 27369
rect 7837 27317 7853 27369
rect 7905 27317 7921 27369
rect 7973 27317 7988 27369
rect 8040 27317 8055 27369
rect 8107 27317 8122 27369
rect 8174 27317 8189 27369
rect 8241 27317 8256 27369
rect 8308 27317 8323 27369
rect 8375 27317 8390 27369
rect 8442 27317 8457 27369
rect 8509 27317 8524 27369
rect 8576 27317 8582 27369
rect 7439 27283 8582 27317
rect 7439 27243 7461 27283
rect 7517 27243 8453 27283
rect 8509 27243 8582 27283
rect 7439 27191 7445 27243
rect 7497 27191 7513 27227
rect 7565 27191 7581 27243
rect 7633 27191 7649 27243
rect 7701 27191 7717 27243
rect 7769 27191 7785 27243
rect 7837 27191 7853 27243
rect 7905 27191 7921 27243
rect 7973 27191 7988 27243
rect 8040 27191 8055 27243
rect 8107 27191 8122 27243
rect 8174 27191 8189 27243
rect 8241 27191 8256 27243
rect 8308 27191 8323 27243
rect 8375 27191 8390 27243
rect 8442 27227 8453 27243
rect 8442 27191 8457 27227
rect 8509 27191 8524 27243
rect 8576 27191 8582 27243
rect 9423 28581 9429 28633
rect 9481 28620 9517 28633
rect 9501 28581 9517 28620
rect 9569 28581 9575 28633
rect 9423 28564 9445 28581
rect 9501 28564 9575 28581
rect 9423 28559 9575 28564
rect 9423 28507 9429 28559
rect 9481 28507 9517 28559
rect 9569 28507 9575 28559
rect 9423 28485 9575 28507
rect 9423 28433 9429 28485
rect 9481 28453 9517 28485
rect 9501 28433 9517 28453
rect 9569 28433 9575 28485
rect 9423 28397 9445 28433
rect 9501 28397 9575 28433
rect 9423 28286 9575 28397
rect 9423 28230 9445 28286
rect 9501 28230 9575 28286
rect 9423 28119 9575 28230
rect 14281 28627 14639 28633
rect 14281 28575 14282 28627
rect 14334 28577 14358 28627
rect 14410 28577 14434 28627
rect 14486 28577 14510 28627
rect 14562 28577 14586 28627
rect 14339 28575 14358 28577
rect 14562 28575 14577 28577
rect 14638 28575 14639 28627
rect 14281 28562 14283 28575
rect 14339 28562 14381 28575
rect 14437 28562 14479 28575
rect 14535 28562 14577 28575
rect 14633 28562 14639 28575
rect 14281 28510 14282 28562
rect 14339 28521 14358 28562
rect 14562 28521 14577 28562
rect 14334 28510 14358 28521
rect 14410 28510 14434 28521
rect 14486 28510 14510 28521
rect 14562 28510 14586 28521
rect 14638 28510 14639 28562
rect 14281 28497 14639 28510
rect 14281 28445 14282 28497
rect 14339 28445 14358 28497
rect 14562 28445 14577 28497
rect 14638 28445 14639 28497
rect 14281 28441 14283 28445
rect 14339 28441 14381 28445
rect 14437 28441 14479 28445
rect 14535 28441 14577 28445
rect 14633 28441 14639 28445
rect 14281 28432 14639 28441
rect 14281 28380 14282 28432
rect 14334 28417 14358 28432
rect 14410 28417 14434 28432
rect 14486 28417 14510 28432
rect 14562 28417 14586 28432
rect 14339 28380 14358 28417
rect 14562 28380 14577 28417
rect 14638 28380 14639 28432
rect 14281 28367 14283 28380
rect 14339 28367 14381 28380
rect 14437 28367 14479 28380
rect 14535 28367 14577 28380
rect 14633 28367 14639 28380
rect 14281 28315 14282 28367
rect 14339 28361 14358 28367
rect 14562 28361 14577 28367
rect 14334 28337 14358 28361
rect 14410 28337 14434 28361
rect 14486 28337 14510 28361
rect 14562 28337 14586 28361
rect 14339 28315 14358 28337
rect 14562 28315 14577 28337
rect 14638 28315 14639 28367
rect 14281 28302 14283 28315
rect 14339 28302 14381 28315
rect 14437 28302 14479 28315
rect 14535 28302 14577 28315
rect 14633 28302 14639 28315
rect 14281 28250 14282 28302
rect 14339 28281 14358 28302
rect 14562 28281 14577 28302
rect 14334 28257 14358 28281
rect 14410 28257 14434 28281
rect 14486 28257 14510 28281
rect 14562 28257 14586 28281
rect 14339 28250 14358 28257
rect 14562 28250 14577 28257
rect 14638 28250 14639 28302
rect 14281 28237 14283 28250
rect 14339 28237 14381 28250
rect 14437 28237 14479 28250
rect 14535 28237 14577 28250
rect 14633 28237 14639 28250
rect 14281 28185 14282 28237
rect 14339 28201 14358 28237
rect 14562 28201 14577 28237
rect 14334 28185 14358 28201
rect 14410 28185 14434 28201
rect 14486 28185 14510 28201
rect 14562 28185 14586 28201
rect 14638 28185 14639 28237
rect 14281 28177 14639 28185
rect 14281 28171 14283 28177
rect 14339 28171 14381 28177
rect 14437 28171 14479 28177
rect 14535 28171 14577 28177
rect 14633 28171 14639 28177
rect 9423 28063 9445 28119
rect 9501 28063 9575 28119
rect 9423 27952 9575 28063
rect 9423 27896 9445 27952
rect 9501 27896 9575 27952
rect 9423 27785 9575 27896
rect 9423 27729 9445 27785
rect 9501 27729 9575 27785
rect 9423 27618 9575 27729
rect 9423 27562 9445 27618
rect 9501 27562 9575 27618
rect 9423 27451 9575 27562
rect 9423 27395 9445 27451
rect 9501 27395 9575 27451
rect 9423 27364 9575 27395
rect 9475 27312 9523 27364
rect 9423 27283 9575 27312
rect 9423 27268 9445 27283
rect 9501 27268 9575 27283
rect 9501 27227 9523 27268
rect 9475 27216 9523 27227
rect 9423 27210 9575 27216
rect 12151 28124 12893 28129
rect 12151 28072 12157 28124
rect 12209 28072 12225 28124
rect 12277 28072 12293 28124
rect 12345 28072 12361 28124
rect 12413 28072 12429 28124
rect 12481 28072 12497 28124
rect 12549 28072 12565 28124
rect 12617 28072 12633 28124
rect 12685 28072 12701 28124
rect 12753 28072 12768 28124
rect 12820 28072 12835 28124
rect 12887 28072 12893 28124
rect 12151 28058 12893 28072
rect 12151 28006 12157 28058
rect 12209 28006 12225 28058
rect 12277 28006 12293 28058
rect 12345 28006 12361 28058
rect 12413 28006 12429 28058
rect 12481 28006 12497 28058
rect 12549 28006 12565 28058
rect 12617 28006 12633 28058
rect 12685 28006 12701 28058
rect 12753 28006 12768 28058
rect 12820 28006 12835 28058
rect 12887 28006 12893 28058
rect 12151 27992 12893 28006
rect 12151 27940 12157 27992
rect 12209 27940 12225 27992
rect 12277 27940 12293 27992
rect 12345 27940 12361 27992
rect 12413 27940 12429 27992
rect 12481 27940 12497 27992
rect 12549 27940 12565 27992
rect 12617 27940 12633 27992
rect 12685 27940 12701 27992
rect 12753 27940 12768 27992
rect 12820 27940 12835 27992
rect 12887 27940 12893 27992
rect 12151 27926 12893 27940
rect 12151 27874 12157 27926
rect 12209 27874 12225 27926
rect 12277 27874 12293 27926
rect 12345 27874 12361 27926
rect 12413 27874 12429 27926
rect 12481 27874 12497 27926
rect 12549 27874 12565 27926
rect 12617 27874 12633 27926
rect 12685 27874 12701 27926
rect 12753 27874 12768 27926
rect 12820 27874 12835 27926
rect 12887 27874 12893 27926
rect 12151 27860 12893 27874
rect 12151 27808 12157 27860
rect 12209 27808 12225 27860
rect 12277 27808 12293 27860
rect 12345 27808 12361 27860
rect 12413 27808 12429 27860
rect 12481 27808 12497 27860
rect 12549 27808 12565 27860
rect 12617 27808 12633 27860
rect 12685 27808 12701 27860
rect 12753 27808 12768 27860
rect 12820 27808 12835 27860
rect 12887 27808 12893 27860
rect 12151 27794 12893 27808
rect 12151 27742 12157 27794
rect 12209 27742 12225 27794
rect 12277 27742 12293 27794
rect 12345 27742 12361 27794
rect 12413 27742 12429 27794
rect 12481 27742 12497 27794
rect 12549 27742 12565 27794
rect 12617 27742 12633 27794
rect 12685 27742 12701 27794
rect 12753 27742 12768 27794
rect 12820 27742 12835 27794
rect 12887 27742 12893 27794
rect 12151 27728 12893 27742
rect 12151 27676 12157 27728
rect 12209 27676 12225 27728
rect 12277 27676 12293 27728
rect 12345 27676 12361 27728
rect 12413 27676 12429 27728
rect 12481 27676 12497 27728
rect 12549 27676 12565 27728
rect 12617 27676 12633 27728
rect 12685 27676 12701 27728
rect 12753 27676 12768 27728
rect 12820 27676 12835 27728
rect 12887 27676 12893 27728
rect 2359 27151 2724 27160
rect 2359 27095 2387 27151
rect 2443 27095 2513 27151
rect 2569 27095 2724 27151
rect 2359 27031 2724 27095
rect 2359 27000 2387 27031
rect 2443 27000 2513 27031
rect 2569 27000 2724 27031
rect 2359 26948 2365 27000
rect 2492 26975 2513 27000
rect 2569 26975 2589 27000
rect 2417 26948 2440 26975
rect 2492 26948 2515 26975
rect 2567 26948 2589 26975
rect 2641 26948 2663 27000
rect 2715 26948 2724 27000
rect 2359 26911 2724 26948
rect 2359 26878 2387 26911
rect 2443 26878 2513 26911
rect 2569 26878 2724 26911
rect 2359 26826 2365 26878
rect 2492 26855 2513 26878
rect 2569 26855 2589 26878
rect 2417 26826 2440 26855
rect 2492 26826 2515 26855
rect 2567 26826 2589 26855
rect 2641 26826 2663 26878
rect 2715 26826 2724 26878
rect 2359 26809 2724 26826
rect 2480 26181 2672 26187
rect 2532 26176 2550 26181
rect 2541 26129 2550 26176
rect 2602 26176 2620 26181
rect 2602 26129 2611 26176
rect 2480 26120 2485 26129
rect 2541 26120 2611 26129
rect 2667 26120 2672 26129
rect 2480 26111 2672 26120
rect 2532 26081 2550 26111
rect 2541 26059 2550 26081
rect 2602 26081 2620 26111
rect 2602 26059 2611 26081
rect 2480 26041 2485 26059
rect 2541 26041 2611 26059
rect 2667 26041 2672 26059
rect 2541 26025 2550 26041
rect 2532 25989 2550 26025
rect 2602 26025 2611 26041
rect 2602 25989 2620 26025
rect 2480 25986 2672 25989
rect 2480 25971 2485 25986
rect 2541 25971 2611 25986
rect 2667 25971 2672 25986
rect 2541 25930 2550 25971
rect 2532 25919 2550 25930
rect 2602 25930 2611 25971
rect 2602 25919 2620 25930
rect 2480 25901 2672 25919
rect 2532 25891 2550 25901
rect 2541 25849 2550 25891
rect 2602 25891 2620 25901
rect 2602 25849 2611 25891
rect 2480 25835 2485 25849
rect 2541 25835 2611 25849
rect 2667 25835 2672 25849
rect 2480 25831 2672 25835
rect 2532 25795 2550 25831
rect 2541 25779 2550 25795
rect 2602 25795 2620 25831
rect 2602 25779 2611 25795
rect 2480 25760 2485 25779
rect 2541 25760 2611 25779
rect 2667 25760 2672 25779
rect 2541 25739 2550 25760
rect 2532 25708 2550 25739
rect 2602 25739 2611 25760
rect 2602 25708 2620 25739
rect 2480 25699 2672 25708
rect 2480 25689 2485 25699
rect 2541 25689 2611 25699
rect 2667 25689 2672 25699
rect 2541 25643 2550 25689
rect 2532 25637 2550 25643
rect 2602 25643 2611 25689
rect 2602 25637 2620 25643
rect 2480 25631 2672 25637
rect 3472 26181 3664 26187
rect 3524 26176 3542 26181
rect 3533 26129 3542 26176
rect 3594 26176 3612 26181
rect 3594 26129 3603 26176
rect 3472 26120 3477 26129
rect 3533 26120 3603 26129
rect 3659 26120 3664 26129
rect 3472 26111 3664 26120
rect 3524 26081 3542 26111
rect 3533 26059 3542 26081
rect 3594 26081 3612 26111
rect 3594 26059 3603 26081
rect 3472 26041 3477 26059
rect 3533 26041 3603 26059
rect 3659 26041 3664 26059
rect 3533 26025 3542 26041
rect 3524 25989 3542 26025
rect 3594 26025 3603 26041
rect 3594 25989 3612 26025
rect 3472 25986 3664 25989
rect 3472 25971 3477 25986
rect 3533 25971 3603 25986
rect 3659 25971 3664 25986
rect 3533 25930 3542 25971
rect 3524 25919 3542 25930
rect 3594 25930 3603 25971
rect 3594 25919 3612 25930
rect 3472 25901 3664 25919
rect 3524 25891 3542 25901
rect 3533 25849 3542 25891
rect 3594 25891 3612 25901
rect 3594 25849 3603 25891
rect 3472 25835 3477 25849
rect 3533 25835 3603 25849
rect 3659 25835 3664 25849
rect 3472 25831 3664 25835
rect 3524 25795 3542 25831
rect 3533 25779 3542 25795
rect 3594 25795 3612 25831
rect 3594 25779 3603 25795
rect 3472 25760 3477 25779
rect 3533 25760 3603 25779
rect 3659 25760 3664 25779
rect 3533 25739 3542 25760
rect 3524 25708 3542 25739
rect 3594 25739 3603 25760
rect 3594 25708 3612 25739
rect 3472 25699 3664 25708
rect 3472 25689 3477 25699
rect 3533 25689 3603 25699
rect 3659 25689 3664 25699
rect 3533 25643 3542 25689
rect 3524 25637 3542 25643
rect 3594 25643 3603 25689
rect 3594 25637 3612 25643
rect 3472 25631 3664 25637
rect 4464 26181 4656 26187
rect 4516 26176 4534 26181
rect 4525 26129 4534 26176
rect 4586 26176 4604 26181
rect 4586 26129 4595 26176
rect 4464 26120 4469 26129
rect 4525 26120 4595 26129
rect 4651 26120 4656 26129
rect 4464 26111 4656 26120
rect 4516 26081 4534 26111
rect 4525 26059 4534 26081
rect 4586 26081 4604 26111
rect 4586 26059 4595 26081
rect 4464 26041 4469 26059
rect 4525 26041 4595 26059
rect 4651 26041 4656 26059
rect 4525 26025 4534 26041
rect 4516 25989 4534 26025
rect 4586 26025 4595 26041
rect 4586 25989 4604 26025
rect 4464 25986 4656 25989
rect 4464 25971 4469 25986
rect 4525 25971 4595 25986
rect 4651 25971 4656 25986
rect 4525 25930 4534 25971
rect 4516 25919 4534 25930
rect 4586 25930 4595 25971
rect 4586 25919 4604 25930
rect 4464 25901 4656 25919
rect 4516 25891 4534 25901
rect 4525 25849 4534 25891
rect 4586 25891 4604 25901
rect 4586 25849 4595 25891
rect 4464 25835 4469 25849
rect 4525 25835 4595 25849
rect 4651 25835 4656 25849
rect 4464 25831 4656 25835
rect 4516 25795 4534 25831
rect 4525 25779 4534 25795
rect 4586 25795 4604 25831
rect 4586 25779 4595 25795
rect 4464 25760 4469 25779
rect 4525 25760 4595 25779
rect 4651 25760 4656 25779
rect 4525 25739 4534 25760
rect 4516 25708 4534 25739
rect 4586 25739 4595 25760
rect 4586 25708 4604 25739
rect 4464 25699 4656 25708
rect 4464 25689 4469 25699
rect 4525 25689 4595 25699
rect 4651 25689 4656 25699
rect 4525 25643 4534 25689
rect 4516 25637 4534 25643
rect 4586 25643 4595 25689
rect 4586 25637 4604 25643
rect 4464 25631 4656 25637
rect 5456 26181 5648 26187
rect 5508 26176 5526 26181
rect 5517 26129 5526 26176
rect 5578 26176 5596 26181
rect 5578 26129 5587 26176
rect 5456 26120 5461 26129
rect 5517 26120 5587 26129
rect 5643 26120 5648 26129
rect 5456 26111 5648 26120
rect 5508 26081 5526 26111
rect 5517 26059 5526 26081
rect 5578 26081 5596 26111
rect 5578 26059 5587 26081
rect 5456 26041 5461 26059
rect 5517 26041 5587 26059
rect 5643 26041 5648 26059
rect 5517 26025 5526 26041
rect 5508 25989 5526 26025
rect 5578 26025 5587 26041
rect 5578 25989 5596 26025
rect 5456 25986 5648 25989
rect 5456 25971 5461 25986
rect 5517 25971 5587 25986
rect 5643 25971 5648 25986
rect 5517 25930 5526 25971
rect 5508 25919 5526 25930
rect 5578 25930 5587 25971
rect 5578 25919 5596 25930
rect 5456 25901 5648 25919
rect 5508 25891 5526 25901
rect 5517 25849 5526 25891
rect 5578 25891 5596 25901
rect 5578 25849 5587 25891
rect 5456 25835 5461 25849
rect 5517 25835 5587 25849
rect 5643 25835 5648 25849
rect 5456 25831 5648 25835
rect 5508 25795 5526 25831
rect 5517 25779 5526 25795
rect 5578 25795 5596 25831
rect 5578 25779 5587 25795
rect 5456 25760 5461 25779
rect 5517 25760 5587 25779
rect 5643 25760 5648 25779
rect 5517 25739 5526 25760
rect 5508 25708 5526 25739
rect 5578 25739 5587 25760
rect 5578 25708 5596 25739
rect 5456 25699 5648 25708
rect 5456 25689 5461 25699
rect 5517 25689 5587 25699
rect 5643 25689 5648 25699
rect 5517 25643 5526 25689
rect 5508 25637 5526 25643
rect 5578 25643 5587 25689
rect 5578 25637 5596 25643
rect 5456 25631 5648 25637
rect 6448 26181 6640 26187
rect 6500 26176 6518 26181
rect 6509 26129 6518 26176
rect 6570 26176 6588 26181
rect 6570 26129 6579 26176
rect 6448 26120 6453 26129
rect 6509 26120 6579 26129
rect 6635 26120 6640 26129
rect 6448 26111 6640 26120
rect 6500 26081 6518 26111
rect 6509 26059 6518 26081
rect 6570 26081 6588 26111
rect 6570 26059 6579 26081
rect 6448 26041 6453 26059
rect 6509 26041 6579 26059
rect 6635 26041 6640 26059
rect 6509 26025 6518 26041
rect 6500 25989 6518 26025
rect 6570 26025 6579 26041
rect 6570 25989 6588 26025
rect 6448 25986 6640 25989
rect 6448 25971 6453 25986
rect 6509 25971 6579 25986
rect 6635 25971 6640 25986
rect 6509 25930 6518 25971
rect 6500 25919 6518 25930
rect 6570 25930 6579 25971
rect 6570 25919 6588 25930
rect 6448 25901 6640 25919
rect 6500 25891 6518 25901
rect 6509 25849 6518 25891
rect 6570 25891 6588 25901
rect 6570 25849 6579 25891
rect 6448 25835 6453 25849
rect 6509 25835 6579 25849
rect 6635 25835 6640 25849
rect 6448 25831 6640 25835
rect 6500 25795 6518 25831
rect 6509 25779 6518 25795
rect 6570 25795 6588 25831
rect 6570 25779 6579 25795
rect 6448 25760 6453 25779
rect 6509 25760 6579 25779
rect 6635 25760 6640 25779
rect 6509 25739 6518 25760
rect 6500 25708 6518 25739
rect 6570 25739 6579 25760
rect 6570 25708 6588 25739
rect 6448 25699 6640 25708
rect 6448 25689 6453 25699
rect 6509 25689 6579 25699
rect 6635 25689 6640 25699
rect 6509 25643 6518 25689
rect 6500 25637 6518 25643
rect 6570 25643 6579 25689
rect 6570 25637 6588 25643
rect 6448 25631 6640 25637
rect 7440 26181 7632 26187
rect 7492 26176 7510 26181
rect 7501 26129 7510 26176
rect 7562 26176 7580 26181
rect 7562 26129 7571 26176
rect 7440 26120 7445 26129
rect 7501 26120 7571 26129
rect 7627 26120 7632 26129
rect 7440 26111 7632 26120
rect 7492 26081 7510 26111
rect 7501 26059 7510 26081
rect 7562 26081 7580 26111
rect 7562 26059 7571 26081
rect 7440 26041 7445 26059
rect 7501 26041 7571 26059
rect 7627 26041 7632 26059
rect 7501 26025 7510 26041
rect 7492 25989 7510 26025
rect 7562 26025 7571 26041
rect 7562 25989 7580 26025
rect 7440 25986 7632 25989
rect 7440 25971 7445 25986
rect 7501 25971 7571 25986
rect 7627 25971 7632 25986
rect 7501 25930 7510 25971
rect 7492 25919 7510 25930
rect 7562 25930 7571 25971
rect 7562 25919 7580 25930
rect 7440 25901 7632 25919
rect 7492 25891 7510 25901
rect 7501 25849 7510 25891
rect 7562 25891 7580 25901
rect 7562 25849 7571 25891
rect 7440 25835 7445 25849
rect 7501 25835 7571 25849
rect 7627 25835 7632 25849
rect 7440 25831 7632 25835
rect 7492 25795 7510 25831
rect 7501 25779 7510 25795
rect 7562 25795 7580 25831
rect 7562 25779 7571 25795
rect 7440 25760 7445 25779
rect 7501 25760 7571 25779
rect 7627 25760 7632 25779
rect 7501 25739 7510 25760
rect 7492 25708 7510 25739
rect 7562 25739 7571 25760
rect 7562 25708 7580 25739
rect 7440 25699 7632 25708
rect 7440 25689 7445 25699
rect 7501 25689 7571 25699
rect 7627 25689 7632 25699
rect 7501 25643 7510 25689
rect 7492 25637 7510 25643
rect 7562 25643 7571 25689
rect 7562 25637 7580 25643
rect 7440 25631 7632 25637
rect 8432 26181 8624 26187
rect 8484 26176 8502 26181
rect 8493 26129 8502 26176
rect 8554 26176 8572 26181
rect 8554 26129 8563 26176
rect 8432 26120 8437 26129
rect 8493 26120 8563 26129
rect 8619 26120 8624 26129
rect 8432 26111 8624 26120
rect 8484 26081 8502 26111
rect 8493 26059 8502 26081
rect 8554 26081 8572 26111
rect 8554 26059 8563 26081
rect 8432 26041 8437 26059
rect 8493 26041 8563 26059
rect 8619 26041 8624 26059
rect 8493 26025 8502 26041
rect 8484 25989 8502 26025
rect 8554 26025 8563 26041
rect 8554 25989 8572 26025
rect 8432 25986 8624 25989
rect 8432 25971 8437 25986
rect 8493 25971 8563 25986
rect 8619 25971 8624 25986
rect 8493 25930 8502 25971
rect 8484 25919 8502 25930
rect 8554 25930 8563 25971
rect 8554 25919 8572 25930
rect 8432 25901 8624 25919
rect 8484 25891 8502 25901
rect 8493 25849 8502 25891
rect 8554 25891 8572 25901
rect 8554 25849 8563 25891
rect 8432 25835 8437 25849
rect 8493 25835 8563 25849
rect 8619 25835 8624 25849
rect 8432 25831 8624 25835
rect 8484 25795 8502 25831
rect 8493 25779 8502 25795
rect 8554 25795 8572 25831
rect 8554 25779 8563 25795
rect 8432 25760 8437 25779
rect 8493 25760 8563 25779
rect 8619 25760 8624 25779
rect 8493 25739 8502 25760
rect 8484 25708 8502 25739
rect 8554 25739 8563 25760
rect 8554 25708 8572 25739
rect 8432 25699 8624 25708
rect 8432 25689 8437 25699
rect 8493 25689 8563 25699
rect 8619 25689 8624 25699
rect 8493 25643 8502 25689
rect 8484 25637 8502 25643
rect 8554 25643 8563 25689
rect 8554 25637 8572 25643
rect 8432 25631 8624 25637
rect 9424 26181 9616 26187
rect 9476 26176 9494 26181
rect 9485 26129 9494 26176
rect 9546 26176 9564 26181
rect 9546 26129 9555 26176
rect 9424 26120 9429 26129
rect 9485 26120 9555 26129
rect 9611 26120 9616 26129
rect 9424 26111 9616 26120
rect 9476 26081 9494 26111
rect 9485 26059 9494 26081
rect 9546 26081 9564 26111
rect 9546 26059 9555 26081
rect 9424 26041 9429 26059
rect 9485 26041 9555 26059
rect 9611 26041 9616 26059
rect 9485 26025 9494 26041
rect 9476 25989 9494 26025
rect 9546 26025 9555 26041
rect 9546 25989 9564 26025
rect 9424 25986 9616 25989
rect 9424 25971 9429 25986
rect 9485 25971 9555 25986
rect 9611 25971 9616 25986
rect 9485 25930 9494 25971
rect 9476 25919 9494 25930
rect 9546 25930 9555 25971
rect 9546 25919 9564 25930
rect 9424 25901 9616 25919
rect 9476 25891 9494 25901
rect 9485 25849 9494 25891
rect 9546 25891 9564 25901
rect 9546 25849 9555 25891
rect 9424 25835 9429 25849
rect 9485 25835 9555 25849
rect 9611 25835 9616 25849
rect 9424 25831 9616 25835
rect 9476 25795 9494 25831
rect 9485 25779 9494 25795
rect 9546 25795 9564 25831
rect 9546 25779 9555 25795
rect 9424 25760 9429 25779
rect 9485 25760 9555 25779
rect 9611 25760 9616 25779
rect 9485 25739 9494 25760
rect 9476 25708 9494 25739
rect 9546 25739 9555 25760
rect 9546 25708 9564 25739
rect 9424 25699 9616 25708
rect 9424 25689 9429 25699
rect 9485 25689 9555 25699
rect 9611 25689 9616 25699
rect 9485 25643 9494 25689
rect 9476 25637 9494 25643
rect 9546 25643 9555 25689
rect 9546 25637 9564 25643
rect 9424 25631 9616 25637
rect 1297 24985 1303 25037
rect 1355 24985 1371 25037
rect 1423 24985 1439 25037
rect 1491 24985 1507 25037
rect 1559 24985 1575 25037
rect 1627 24985 1643 25037
rect 1695 24985 1711 25037
rect 1763 24985 1779 25037
rect 1831 24985 1847 25037
rect 1899 24985 1914 25037
rect 1966 24985 1981 25037
rect 2033 24985 2039 25037
rect 1297 24967 2039 24985
rect 1297 24915 1303 24967
rect 1355 24915 1371 24967
rect 1423 24915 1439 24967
rect 1491 24915 1507 24967
rect 1559 24915 1575 24967
rect 1627 24915 1643 24967
rect 1695 24915 1711 24967
rect 1763 24915 1779 24967
rect 1831 24915 1847 24967
rect 1899 24915 1914 24967
rect 1966 24915 1981 24967
rect 2033 24915 2039 24967
rect 1297 24897 2039 24915
rect 1297 24845 1303 24897
rect 1355 24845 1371 24897
rect 1423 24845 1439 24897
rect 1491 24845 1507 24897
rect 1559 24845 1575 24897
rect 1627 24845 1643 24897
rect 1695 24845 1711 24897
rect 1763 24845 1779 24897
rect 1831 24845 1847 24897
rect 1899 24845 1914 24897
rect 1966 24845 1981 24897
rect 2033 24845 2039 24897
rect 1297 24827 2039 24845
rect 1297 24775 1303 24827
rect 1355 24775 1371 24827
rect 1423 24775 1439 24827
rect 1491 24775 1507 24827
rect 1559 24775 1575 24827
rect 1627 24775 1643 24827
rect 1695 24775 1711 24827
rect 1763 24775 1779 24827
rect 1831 24775 1847 24827
rect 1899 24775 1914 24827
rect 1966 24775 1981 24827
rect 2033 24775 2039 24827
rect 1297 24757 2039 24775
rect 1297 24705 1303 24757
rect 1355 24705 1371 24757
rect 1423 24705 1439 24757
rect 1491 24705 1507 24757
rect 1559 24705 1575 24757
rect 1627 24705 1643 24757
rect 1695 24705 1711 24757
rect 1763 24705 1779 24757
rect 1831 24705 1847 24757
rect 1899 24705 1914 24757
rect 1966 24705 1981 24757
rect 2033 24705 2039 24757
rect 1297 24687 2039 24705
rect 1297 24635 1303 24687
rect 1355 24635 1371 24687
rect 1423 24635 1439 24687
rect 1491 24635 1507 24687
rect 1559 24635 1575 24687
rect 1627 24635 1643 24687
rect 1695 24635 1711 24687
rect 1763 24635 1779 24687
rect 1831 24635 1847 24687
rect 1899 24635 1914 24687
rect 1966 24635 1981 24687
rect 2033 24635 2039 24687
rect 1297 24617 2039 24635
rect 1297 24565 1303 24617
rect 1355 24565 1371 24617
rect 1423 24565 1439 24617
rect 1491 24565 1507 24617
rect 1559 24565 1575 24617
rect 1627 24565 1643 24617
rect 1695 24565 1711 24617
rect 1763 24565 1779 24617
rect 1831 24565 1847 24617
rect 1899 24565 1914 24617
rect 1966 24565 1981 24617
rect 2033 24565 2039 24617
rect 1297 24547 2039 24565
rect 1297 24495 1303 24547
rect 1355 24495 1371 24547
rect 1423 24495 1439 24547
rect 1491 24495 1507 24547
rect 1559 24495 1575 24547
rect 1627 24495 1643 24547
rect 1695 24495 1711 24547
rect 1763 24495 1779 24547
rect 1831 24495 1847 24547
rect 1899 24495 1914 24547
rect 1966 24495 1981 24547
rect 2033 24495 2039 24547
rect 1297 24492 2039 24495
rect 12151 25037 12893 27676
rect 14281 28119 14282 28171
rect 14339 28121 14358 28171
rect 14562 28121 14577 28171
rect 14334 28119 14358 28121
rect 14410 28119 14434 28121
rect 14486 28119 14510 28121
rect 14562 28119 14586 28121
rect 14638 28119 14639 28171
rect 14281 28105 14639 28119
rect 14281 28053 14282 28105
rect 14334 28097 14358 28105
rect 14410 28097 14434 28105
rect 14486 28097 14510 28105
rect 14562 28097 14586 28105
rect 14339 28053 14358 28097
rect 14562 28053 14577 28097
rect 14638 28053 14639 28105
rect 14281 28041 14283 28053
rect 14339 28041 14381 28053
rect 14437 28041 14479 28053
rect 14535 28041 14577 28053
rect 14633 28041 14639 28053
rect 14281 28039 14639 28041
rect 14281 27987 14282 28039
rect 14334 28017 14358 28039
rect 14410 28017 14434 28039
rect 14486 28017 14510 28039
rect 14562 28017 14586 28039
rect 14339 27987 14358 28017
rect 14562 27987 14577 28017
rect 14638 27987 14639 28039
rect 14281 27973 14283 27987
rect 14339 27973 14381 27987
rect 14437 27973 14479 27987
rect 14535 27973 14577 27987
rect 14633 27973 14639 27987
rect 14281 27921 14282 27973
rect 14339 27961 14358 27973
rect 14562 27961 14577 27973
rect 14334 27937 14358 27961
rect 14410 27937 14434 27961
rect 14486 27937 14510 27961
rect 14562 27937 14586 27961
rect 14339 27921 14358 27937
rect 14562 27921 14577 27937
rect 14638 27921 14639 27973
rect 14281 27907 14283 27921
rect 14339 27907 14381 27921
rect 14437 27907 14479 27921
rect 14535 27907 14577 27921
rect 14633 27907 14639 27921
rect 14281 27855 14282 27907
rect 14339 27881 14358 27907
rect 14562 27881 14577 27907
rect 14334 27857 14358 27881
rect 14410 27857 14434 27881
rect 14486 27857 14510 27881
rect 14562 27857 14586 27881
rect 14339 27855 14358 27857
rect 14562 27855 14577 27857
rect 14638 27855 14639 27907
rect 14281 27841 14283 27855
rect 14339 27841 14381 27855
rect 14437 27841 14479 27855
rect 14535 27841 14577 27855
rect 14633 27841 14639 27855
rect 14281 27789 14282 27841
rect 14339 27801 14358 27841
rect 14562 27801 14577 27841
rect 14334 27789 14358 27801
rect 14410 27789 14434 27801
rect 14486 27789 14510 27801
rect 14562 27789 14586 27801
rect 14638 27789 14639 27841
rect 14281 27777 14639 27789
rect 14281 27775 14283 27777
rect 14339 27775 14381 27777
rect 14437 27775 14479 27777
rect 14535 27775 14577 27777
rect 14633 27775 14639 27777
rect 14281 27723 14282 27775
rect 14339 27723 14358 27775
rect 14562 27723 14577 27775
rect 14638 27723 14639 27775
rect 14281 27721 14283 27723
rect 14339 27721 14381 27723
rect 14437 27721 14479 27723
rect 14535 27721 14577 27723
rect 14633 27721 14639 27723
rect 14281 27709 14639 27721
rect 14281 27657 14282 27709
rect 14334 27697 14358 27709
rect 14410 27697 14434 27709
rect 14486 27697 14510 27709
rect 14562 27697 14586 27709
rect 14339 27657 14358 27697
rect 14562 27657 14577 27697
rect 14638 27657 14639 27709
rect 14281 27643 14283 27657
rect 14339 27643 14381 27657
rect 14437 27643 14479 27657
rect 14535 27643 14577 27657
rect 14633 27643 14639 27657
rect 14281 27591 14282 27643
rect 14339 27641 14358 27643
rect 14562 27641 14577 27643
rect 14334 27617 14358 27641
rect 14410 27617 14434 27641
rect 14486 27617 14510 27641
rect 14562 27617 14586 27641
rect 14339 27591 14358 27617
rect 14562 27591 14577 27617
rect 14638 27591 14639 27643
rect 14281 27577 14283 27591
rect 14339 27577 14381 27591
rect 14437 27577 14479 27591
rect 14535 27577 14577 27591
rect 14633 27577 14639 27591
rect 14281 27525 14282 27577
rect 14339 27561 14358 27577
rect 14562 27561 14577 27577
rect 14334 27537 14358 27561
rect 14410 27537 14434 27561
rect 14486 27537 14510 27561
rect 14562 27537 14586 27561
rect 14339 27525 14358 27537
rect 14562 27525 14577 27537
rect 14638 27525 14639 27577
rect 14281 27511 14283 27525
rect 14339 27511 14381 27525
rect 14437 27511 14479 27525
rect 14535 27511 14577 27525
rect 14633 27511 14639 27525
rect 14281 27459 14282 27511
rect 14339 27481 14358 27511
rect 14562 27481 14577 27511
rect 14334 27459 14358 27481
rect 14410 27459 14434 27481
rect 14486 27459 14510 27481
rect 14562 27459 14586 27481
rect 14638 27459 14639 27511
rect 14281 27457 14639 27459
rect 14281 27445 14283 27457
rect 14339 27445 14381 27457
rect 14437 27445 14479 27457
rect 14535 27445 14577 27457
rect 14633 27445 14639 27457
rect 14281 27393 14282 27445
rect 14339 27401 14358 27445
rect 14562 27401 14577 27445
rect 14334 27393 14358 27401
rect 14410 27393 14434 27401
rect 14486 27393 14510 27401
rect 14562 27393 14586 27401
rect 14638 27393 14639 27445
rect 14281 27379 14639 27393
rect 14281 27327 14282 27379
rect 14334 27377 14358 27379
rect 14410 27377 14434 27379
rect 14486 27377 14510 27379
rect 14562 27377 14586 27379
rect 14339 27327 14358 27377
rect 14562 27327 14577 27377
rect 14638 27327 14639 27379
rect 14281 27321 14283 27327
rect 14339 27321 14381 27327
rect 14437 27321 14479 27327
rect 14535 27321 14577 27327
rect 14633 27321 14639 27327
rect 14281 27313 14639 27321
rect 14281 27261 14282 27313
rect 14334 27297 14358 27313
rect 14410 27297 14434 27313
rect 14486 27297 14510 27313
rect 14562 27297 14586 27313
rect 14339 27261 14358 27297
rect 14562 27261 14577 27297
rect 14638 27261 14639 27313
rect 14281 27247 14283 27261
rect 14339 27247 14381 27261
rect 14437 27247 14479 27261
rect 14535 27247 14577 27261
rect 14633 27247 14639 27261
rect 14281 27195 14282 27247
rect 14339 27241 14358 27247
rect 14562 27241 14577 27247
rect 14334 27217 14358 27241
rect 14410 27217 14434 27241
rect 14486 27217 14510 27241
rect 14562 27217 14586 27241
rect 14339 27195 14358 27217
rect 14562 27195 14577 27217
rect 14638 27195 14639 27247
rect 14281 27161 14283 27195
rect 14339 27161 14381 27195
rect 14437 27161 14479 27195
rect 14535 27161 14577 27195
rect 14633 27161 14639 27195
rect 14281 27137 14639 27161
rect 14281 27081 14283 27137
rect 14339 27081 14381 27137
rect 14437 27081 14479 27137
rect 14535 27081 14577 27137
rect 14633 27081 14639 27137
rect 14281 27057 14639 27081
rect 14281 27001 14283 27057
rect 14339 27001 14381 27057
rect 14437 27001 14479 27057
rect 14535 27001 14577 27057
rect 14633 27001 14639 27057
rect 14281 26977 14639 27001
rect 14281 26921 14283 26977
rect 14339 26921 14381 26977
rect 14437 26921 14479 26977
rect 14535 26921 14577 26977
rect 14633 26921 14639 26977
rect 14281 26897 14639 26921
rect 13642 26884 14044 26887
rect 13642 26828 13651 26884
rect 13707 26828 13733 26884
rect 13789 26828 13815 26884
rect 13871 26828 13897 26884
rect 13953 26828 13979 26884
rect 14035 26828 14044 26884
rect 13642 26800 14044 26828
rect 13642 26744 13651 26800
rect 13707 26744 13733 26800
rect 13789 26744 13815 26800
rect 13871 26744 13897 26800
rect 13953 26744 13979 26800
rect 14035 26744 14044 26800
rect 13642 26716 14044 26744
rect 13642 26660 13651 26716
rect 13707 26660 13733 26716
rect 13789 26660 13815 26716
rect 13871 26660 13897 26716
rect 13953 26660 13979 26716
rect 14035 26660 14044 26716
rect 13642 26632 14044 26660
rect 13642 26576 13651 26632
rect 13707 26576 13733 26632
rect 13789 26576 13815 26632
rect 13871 26576 13897 26632
rect 13953 26576 13979 26632
rect 14035 26576 14044 26632
rect 13642 26548 14044 26576
rect 13642 26492 13651 26548
rect 13707 26492 13733 26548
rect 13789 26492 13815 26548
rect 13871 26492 13897 26548
rect 13953 26492 13979 26548
rect 14035 26492 14044 26548
rect 13642 26489 14044 26492
rect 14281 26841 14283 26897
rect 14339 26841 14381 26897
rect 14437 26841 14479 26897
rect 14535 26841 14577 26897
rect 14633 26841 14639 26897
rect 14281 26817 14639 26841
rect 14281 26761 14283 26817
rect 14339 26761 14381 26817
rect 14437 26761 14479 26817
rect 14535 26761 14577 26817
rect 14633 26761 14639 26817
rect 14281 26737 14639 26761
rect 14281 26681 14283 26737
rect 14339 26681 14381 26737
rect 14437 26681 14479 26737
rect 14535 26681 14577 26737
rect 14633 26681 14639 26737
rect 14281 26657 14639 26681
rect 14281 26601 14283 26657
rect 14339 26601 14381 26657
rect 14437 26601 14479 26657
rect 14535 26601 14577 26657
rect 14633 26601 14639 26657
rect 14281 26576 14639 26601
rect 14281 26520 14283 26576
rect 14339 26520 14381 26576
rect 14437 26520 14479 26576
rect 14535 26520 14577 26576
rect 14633 26520 14639 26576
rect 14281 26495 14639 26520
rect 12151 24985 12157 25037
rect 12209 24985 12225 25037
rect 12277 24985 12293 25037
rect 12345 24985 12361 25037
rect 12413 24985 12429 25037
rect 12481 24985 12497 25037
rect 12549 24985 12565 25037
rect 12617 24985 12633 25037
rect 12685 24985 12701 25037
rect 12753 24985 12768 25037
rect 12820 24985 12835 25037
rect 12887 24985 12893 25037
rect 12151 24967 12893 24985
rect 12151 24915 12157 24967
rect 12209 24915 12225 24967
rect 12277 24915 12293 24967
rect 12345 24915 12361 24967
rect 12413 24915 12429 24967
rect 12481 24915 12497 24967
rect 12549 24915 12565 24967
rect 12617 24915 12633 24967
rect 12685 24915 12701 24967
rect 12753 24915 12768 24967
rect 12820 24915 12835 24967
rect 12887 24915 12893 24967
rect 12151 24897 12893 24915
rect 12151 24845 12157 24897
rect 12209 24845 12225 24897
rect 12277 24845 12293 24897
rect 12345 24845 12361 24897
rect 12413 24845 12429 24897
rect 12481 24845 12497 24897
rect 12549 24845 12565 24897
rect 12617 24845 12633 24897
rect 12685 24845 12701 24897
rect 12753 24845 12768 24897
rect 12820 24845 12835 24897
rect 12887 24845 12893 24897
rect 12151 24827 12893 24845
rect 12151 24775 12157 24827
rect 12209 24775 12225 24827
rect 12277 24775 12293 24827
rect 12345 24775 12361 24827
rect 12413 24775 12429 24827
rect 12481 24775 12497 24827
rect 12549 24775 12565 24827
rect 12617 24775 12633 24827
rect 12685 24775 12701 24827
rect 12753 24775 12768 24827
rect 12820 24775 12835 24827
rect 12887 24775 12893 24827
rect 12151 24757 12893 24775
rect 12151 24705 12157 24757
rect 12209 24705 12225 24757
rect 12277 24705 12293 24757
rect 12345 24705 12361 24757
rect 12413 24705 12429 24757
rect 12481 24705 12497 24757
rect 12549 24705 12565 24757
rect 12617 24705 12633 24757
rect 12685 24705 12701 24757
rect 12753 24705 12768 24757
rect 12820 24705 12835 24757
rect 12887 24705 12893 24757
rect 12151 24687 12893 24705
rect 12151 24635 12157 24687
rect 12209 24635 12225 24687
rect 12277 24635 12293 24687
rect 12345 24635 12361 24687
rect 12413 24635 12429 24687
rect 12481 24635 12497 24687
rect 12549 24635 12565 24687
rect 12617 24635 12633 24687
rect 12685 24635 12701 24687
rect 12753 24635 12768 24687
rect 12820 24635 12835 24687
rect 12887 24635 12893 24687
rect 12151 24617 12893 24635
rect 12151 24565 12157 24617
rect 12209 24565 12225 24617
rect 12277 24565 12293 24617
rect 12345 24565 12361 24617
rect 12413 24565 12429 24617
rect 12481 24565 12497 24617
rect 12549 24565 12565 24617
rect 12617 24565 12633 24617
rect 12685 24565 12701 24617
rect 12753 24565 12768 24617
rect 12820 24565 12835 24617
rect 12887 24565 12893 24617
rect 12151 24547 12893 24565
rect 12151 24495 12157 24547
rect 12209 24495 12225 24547
rect 12277 24495 12293 24547
rect 12345 24495 12361 24547
rect 12413 24495 12429 24547
rect 12481 24495 12497 24547
rect 12549 24495 12565 24547
rect 12617 24495 12633 24547
rect 12685 24495 12701 24547
rect 12753 24495 12768 24547
rect 12820 24495 12835 24547
rect 12887 24495 12893 24547
rect 12151 24492 12893 24495
rect 14281 26439 14283 26495
rect 14339 26439 14381 26495
rect 14437 26439 14479 26495
rect 14535 26439 14577 26495
rect 14633 26439 14639 26495
rect 14281 26414 14639 26439
rect 14281 26358 14283 26414
rect 14339 26358 14381 26414
rect 14437 26358 14479 26414
rect 14535 26358 14577 26414
rect 14633 26358 14639 26414
rect 14281 26333 14639 26358
rect 14281 26277 14283 26333
rect 14339 26277 14381 26333
rect 14437 26277 14479 26333
rect 14535 26277 14577 26333
rect 14633 26277 14639 26333
rect 14281 26252 14639 26277
rect 14281 26196 14283 26252
rect 14339 26196 14381 26252
rect 14437 26196 14479 26252
rect 14535 26196 14577 26252
rect 14633 26196 14639 26252
rect 14281 26171 14639 26196
rect 14281 26115 14283 26171
rect 14339 26115 14381 26171
rect 14437 26115 14479 26171
rect 14535 26115 14577 26171
rect 14633 26115 14639 26171
rect 14281 26090 14639 26115
rect 14281 26034 14283 26090
rect 14339 26034 14381 26090
rect 14437 26034 14479 26090
rect 14535 26034 14577 26090
rect 14633 26034 14639 26090
rect 14281 26009 14639 26034
rect 14281 25953 14283 26009
rect 14339 25953 14381 26009
rect 14437 25953 14479 26009
rect 14535 25953 14577 26009
rect 14633 25953 14639 26009
rect 14281 25928 14639 25953
rect 14281 25872 14283 25928
rect 14339 25872 14381 25928
rect 14437 25872 14479 25928
rect 14535 25872 14577 25928
rect 14633 25872 14639 25928
rect 14281 25847 14639 25872
rect 14281 25791 14283 25847
rect 14339 25791 14381 25847
rect 14437 25791 14479 25847
rect 14535 25791 14577 25847
rect 14633 25791 14639 25847
rect 14281 25766 14639 25791
rect 14281 25710 14283 25766
rect 14339 25710 14381 25766
rect 14437 25710 14479 25766
rect 14535 25710 14577 25766
rect 14633 25710 14639 25766
rect 14281 25685 14639 25710
rect 14281 25629 14283 25685
rect 14339 25629 14381 25685
rect 14437 25629 14479 25685
rect 14535 25629 14577 25685
rect 14633 25629 14639 25685
rect 14281 25604 14639 25629
rect 14281 25548 14283 25604
rect 14339 25548 14381 25604
rect 14437 25548 14479 25604
rect 14535 25548 14577 25604
rect 14633 25548 14639 25604
rect 14281 25523 14639 25548
rect 14281 25467 14283 25523
rect 14339 25467 14381 25523
rect 14437 25467 14479 25523
rect 14535 25467 14577 25523
rect 14633 25467 14639 25523
rect 14281 25442 14639 25467
rect 14281 25386 14283 25442
rect 14339 25386 14381 25442
rect 14437 25386 14479 25442
rect 14535 25386 14577 25442
rect 14633 25386 14639 25442
rect 14281 25361 14639 25386
rect 14281 25305 14283 25361
rect 14339 25305 14381 25361
rect 14437 25305 14479 25361
rect 14535 25305 14577 25361
rect 14633 25305 14639 25361
rect 14281 25280 14639 25305
rect 14281 25224 14283 25280
rect 14339 25224 14381 25280
rect 14437 25224 14479 25280
rect 14535 25224 14577 25280
rect 14633 25224 14639 25280
rect 14281 25199 14639 25224
rect 14281 25143 14283 25199
rect 14339 25143 14381 25199
rect 14437 25143 14479 25199
rect 14535 25143 14577 25199
rect 14633 25143 14639 25199
rect 14281 25118 14639 25143
rect 14281 25062 14283 25118
rect 14339 25062 14381 25118
rect 14437 25062 14479 25118
rect 14535 25062 14577 25118
rect 14633 25062 14639 25118
rect 14281 25037 14639 25062
rect 14281 24981 14283 25037
rect 14339 24981 14381 25037
rect 14437 24981 14479 25037
rect 14535 24981 14577 25037
rect 14633 24981 14639 25037
rect 14281 24956 14639 24981
rect 14281 24900 14283 24956
rect 14339 24900 14381 24956
rect 14437 24900 14479 24956
rect 14535 24900 14577 24956
rect 14633 24900 14639 24956
rect 14281 24875 14639 24900
rect 14281 24819 14283 24875
rect 14339 24819 14381 24875
rect 14437 24819 14479 24875
rect 14535 24819 14577 24875
rect 14633 24819 14639 24875
rect 14281 24794 14639 24819
rect 14281 24738 14283 24794
rect 14339 24738 14381 24794
rect 14437 24738 14479 24794
rect 14535 24738 14577 24794
rect 14633 24738 14639 24794
rect 14281 24713 14639 24738
rect 14281 24657 14283 24713
rect 14339 24657 14381 24713
rect 14437 24657 14479 24713
rect 14535 24657 14577 24713
rect 14633 24657 14639 24713
rect 14281 24632 14639 24657
rect 14281 24576 14283 24632
rect 14339 24576 14381 24632
rect 14437 24576 14479 24632
rect 14535 24576 14577 24632
rect 14633 24576 14639 24632
rect 14281 24551 14639 24576
rect 14281 24495 14283 24551
rect 14339 24495 14381 24551
rect 14437 24495 14479 24551
rect 14535 24495 14577 24551
rect 14633 24495 14639 24551
rect 164 24423 778 24447
rect 164 24367 242 24423
rect 298 24367 334 24423
rect 390 24367 426 24423
rect 482 24367 518 24423
rect 574 24367 610 24423
rect 666 24367 702 24423
rect 758 24367 778 24423
rect 164 24343 778 24367
rect 164 24287 242 24343
rect 298 24287 334 24343
rect 390 24287 426 24343
rect 482 24287 518 24343
rect 574 24287 610 24343
rect 666 24287 702 24343
rect 758 24287 778 24343
rect 164 24263 778 24287
rect 164 24207 242 24263
rect 298 24207 334 24263
rect 390 24207 426 24263
rect 482 24207 518 24263
rect 574 24207 610 24263
rect 666 24207 702 24263
rect 758 24207 778 24263
rect 164 24183 778 24207
rect 164 24127 242 24183
rect 298 24127 334 24183
rect 390 24127 426 24183
rect 482 24127 518 24183
rect 574 24127 610 24183
rect 666 24127 702 24183
rect 758 24127 778 24183
rect 164 24103 778 24127
rect 164 24047 242 24103
rect 298 24047 334 24103
rect 390 24047 426 24103
rect 482 24047 518 24103
rect 574 24047 610 24103
rect 666 24047 702 24103
rect 758 24047 778 24103
rect 164 24023 778 24047
rect 164 23967 242 24023
rect 298 23967 334 24023
rect 390 23967 426 24023
rect 482 23967 518 24023
rect 574 23967 610 24023
rect 666 23967 702 24023
rect 758 23967 778 24023
rect 164 23943 778 23967
rect 164 23887 242 23943
rect 298 23887 334 23943
rect 390 23887 426 23943
rect 482 23887 518 23943
rect 574 23887 610 23943
rect 666 23887 702 23943
rect 758 23887 778 23943
rect 164 23863 778 23887
rect 164 23807 242 23863
rect 298 23807 334 23863
rect 390 23807 426 23863
rect 482 23807 518 23863
rect 574 23807 610 23863
rect 666 23807 702 23863
rect 758 23807 778 23863
rect 164 23783 778 23807
rect 164 23727 242 23783
rect 298 23727 334 23783
rect 390 23727 426 23783
rect 482 23727 518 23783
rect 574 23727 610 23783
rect 666 23727 702 23783
rect 758 23727 778 23783
rect 164 23703 778 23727
rect 164 23647 242 23703
rect 298 23647 334 23703
rect 390 23647 426 23703
rect 482 23647 518 23703
rect 574 23647 610 23703
rect 666 23647 702 23703
rect 758 23647 778 23703
rect 14281 24470 14639 24495
rect 14281 24414 14283 24470
rect 14339 24414 14381 24470
rect 14437 24414 14479 24470
rect 14535 24414 14577 24470
rect 14633 24414 14639 24470
rect 14281 24389 14639 24414
rect 14281 24333 14283 24389
rect 14339 24333 14381 24389
rect 14437 24333 14479 24389
rect 14535 24333 14577 24389
rect 14633 24333 14639 24389
rect 14281 24308 14639 24333
rect 14281 24252 14283 24308
rect 14339 24252 14381 24308
rect 14437 24252 14479 24308
rect 14535 24252 14577 24308
rect 14633 24252 14639 24308
rect 14281 24227 14639 24252
rect 14281 24171 14283 24227
rect 14339 24171 14381 24227
rect 14437 24171 14479 24227
rect 14535 24171 14577 24227
rect 14633 24171 14639 24227
rect 14281 24146 14639 24171
rect 14281 24090 14283 24146
rect 14339 24090 14381 24146
rect 14437 24090 14479 24146
rect 14535 24090 14577 24146
rect 14633 24090 14639 24146
rect 14281 24065 14639 24090
rect 14281 24009 14283 24065
rect 14339 24009 14381 24065
rect 14437 24009 14479 24065
rect 14535 24009 14577 24065
rect 14633 24009 14639 24065
rect 14281 23984 14639 24009
rect 14281 23928 14283 23984
rect 14339 23928 14381 23984
rect 14437 23928 14479 23984
rect 14535 23928 14577 23984
rect 14633 23928 14639 23984
rect 14281 23903 14639 23928
rect 14281 23847 14283 23903
rect 14339 23847 14381 23903
rect 14437 23847 14479 23903
rect 14535 23847 14577 23903
rect 14633 23847 14639 23903
rect 14281 23822 14639 23847
rect 14281 23766 14283 23822
rect 14339 23766 14381 23822
rect 14437 23766 14479 23822
rect 14535 23766 14577 23822
rect 14633 23766 14639 23822
rect 14281 23741 14639 23766
rect 993 23690 1183 23695
rect 164 23623 778 23647
rect 164 23567 242 23623
rect 298 23567 334 23623
rect 390 23567 426 23623
rect 482 23567 518 23623
rect 574 23567 610 23623
rect 666 23567 702 23623
rect 758 23567 778 23623
rect 164 23543 778 23567
rect 164 23487 242 23543
rect 298 23487 334 23543
rect 390 23487 426 23543
rect 482 23487 518 23543
rect 574 23487 610 23543
rect 666 23487 702 23543
rect 758 23487 778 23543
rect 164 23463 778 23487
rect 164 23407 242 23463
rect 298 23407 334 23463
rect 390 23407 426 23463
rect 482 23407 518 23463
rect 574 23407 610 23463
rect 666 23407 702 23463
rect 758 23407 778 23463
rect 164 23383 778 23407
rect 164 23327 242 23383
rect 298 23327 334 23383
rect 390 23327 426 23383
rect 482 23327 518 23383
rect 574 23327 610 23383
rect 666 23327 702 23383
rect 758 23327 778 23383
rect 164 23303 778 23327
rect 164 23247 242 23303
rect 298 23247 334 23303
rect 390 23247 426 23303
rect 482 23247 518 23303
rect 574 23247 610 23303
rect 666 23247 702 23303
rect 758 23247 778 23303
rect 164 23223 778 23247
rect 164 23167 242 23223
rect 298 23167 334 23223
rect 390 23167 426 23223
rect 482 23167 518 23223
rect 574 23167 610 23223
rect 666 23167 702 23223
rect 758 23167 778 23223
rect 164 23143 778 23167
rect 164 23087 242 23143
rect 298 23087 334 23143
rect 390 23087 426 23143
rect 482 23087 518 23143
rect 574 23087 610 23143
rect 666 23087 702 23143
rect 758 23087 778 23143
rect 164 23063 778 23087
rect 164 23007 242 23063
rect 298 23007 334 23063
rect 390 23007 426 23063
rect 482 23007 518 23063
rect 574 23007 610 23063
rect 666 23007 702 23063
rect 758 23007 778 23063
rect 164 22983 778 23007
rect 164 22927 242 22983
rect 298 22927 334 22983
rect 390 22927 426 22983
rect 482 22927 518 22983
rect 574 22927 610 22983
rect 666 22927 702 22983
rect 758 22927 778 22983
rect 164 22903 778 22927
rect 164 22847 242 22903
rect 298 22847 334 22903
rect 390 22847 426 22903
rect 482 22847 518 22903
rect 574 22847 610 22903
rect 666 22847 702 22903
rect 758 22847 778 22903
rect 164 22822 778 22847
rect 164 22766 242 22822
rect 298 22766 334 22822
rect 390 22766 426 22822
rect 482 22766 518 22822
rect 574 22766 610 22822
rect 666 22766 702 22822
rect 758 22766 778 22822
rect 164 22741 778 22766
rect 164 22685 242 22741
rect 298 22685 334 22741
rect 390 22685 426 22741
rect 482 22685 518 22741
rect 574 22685 610 22741
rect 666 22685 702 22741
rect 758 22685 778 22741
rect 164 22660 778 22685
rect 164 22604 242 22660
rect 298 22604 334 22660
rect 390 22604 426 22660
rect 482 22604 518 22660
rect 574 22604 610 22660
rect 666 22604 702 22660
rect 758 22604 778 22660
rect 164 22579 778 22604
rect 164 22523 242 22579
rect 298 22523 334 22579
rect 390 22523 426 22579
rect 482 22523 518 22579
rect 574 22523 610 22579
rect 666 22523 702 22579
rect 758 22523 778 22579
rect 164 22498 778 22523
rect 164 22442 242 22498
rect 298 22442 334 22498
rect 390 22442 426 22498
rect 482 22442 518 22498
rect 574 22442 610 22498
rect 666 22442 702 22498
rect 758 22442 778 22498
rect 164 22417 778 22442
rect 164 22361 242 22417
rect 298 22361 334 22417
rect 390 22361 426 22417
rect 482 22361 518 22417
rect 574 22361 610 22417
rect 666 22361 702 22417
rect 758 22361 778 22417
rect 164 22336 778 22361
rect 164 22280 242 22336
rect 298 22280 334 22336
rect 390 22280 426 22336
rect 482 22280 518 22336
rect 574 22280 610 22336
rect 666 22280 702 22336
rect 758 22280 778 22336
rect 164 22255 778 22280
rect 164 22199 242 22255
rect 298 22199 334 22255
rect 390 22199 426 22255
rect 482 22199 518 22255
rect 574 22199 610 22255
rect 666 22199 702 22255
rect 758 22199 778 22255
rect 164 22174 778 22199
rect 164 22118 242 22174
rect 298 22118 334 22174
rect 390 22118 426 22174
rect 482 22118 518 22174
rect 574 22118 610 22174
rect 666 22118 702 22174
rect 758 22118 778 22174
rect 164 22093 778 22118
rect 164 22037 242 22093
rect 298 22037 334 22093
rect 390 22037 426 22093
rect 482 22037 518 22093
rect 574 22037 610 22093
rect 666 22037 702 22093
rect 758 22037 778 22093
rect 164 22012 778 22037
rect 164 21956 242 22012
rect 298 21956 334 22012
rect 390 21956 426 22012
rect 482 21956 518 22012
rect 574 21956 610 22012
rect 666 21956 702 22012
rect 758 21956 778 22012
rect 164 21931 778 21956
rect 164 21875 242 21931
rect 298 21875 334 21931
rect 390 21875 426 21931
rect 482 21875 518 21931
rect 574 21875 610 21931
rect 666 21875 702 21931
rect 758 21875 778 21931
rect 164 21850 778 21875
rect 164 21794 242 21850
rect 298 21794 334 21850
rect 390 21794 426 21850
rect 482 21794 518 21850
rect 574 21794 610 21850
rect 666 21794 702 21850
rect 758 21794 778 21850
rect 164 21769 778 21794
rect 164 21713 242 21769
rect 298 21713 334 21769
rect 390 21713 426 21769
rect 482 21713 518 21769
rect 574 21713 610 21769
rect 666 21713 702 21769
rect 758 21713 778 21769
rect 164 21688 778 21713
rect 164 21632 242 21688
rect 298 21632 334 21688
rect 390 21632 426 21688
rect 482 21632 518 21688
rect 574 21632 610 21688
rect 666 21632 702 21688
rect 758 21632 778 21688
rect 164 21607 778 21632
rect 164 21551 242 21607
rect 298 21551 334 21607
rect 390 21551 426 21607
rect 482 21551 518 21607
rect 574 21551 610 21607
rect 666 21551 702 21607
rect 758 21551 778 21607
rect 164 21526 778 21551
rect 164 21470 242 21526
rect 298 21470 334 21526
rect 390 21470 426 21526
rect 482 21470 518 21526
rect 574 21470 610 21526
rect 666 21470 702 21526
rect 758 21470 778 21526
rect 164 21445 778 21470
rect 164 21389 242 21445
rect 298 21389 334 21445
rect 390 21389 426 21445
rect 482 21389 518 21445
rect 574 21389 610 21445
rect 666 21389 702 21445
rect 758 21389 778 21445
rect 164 21364 778 21389
rect 164 21308 242 21364
rect 298 21308 334 21364
rect 390 21308 426 21364
rect 482 21308 518 21364
rect 574 21308 610 21364
rect 666 21308 702 21364
rect 758 21308 778 21364
rect 164 21283 778 21308
rect 164 21227 242 21283
rect 298 21227 334 21283
rect 390 21227 426 21283
rect 482 21227 518 21283
rect 574 21227 610 21283
rect 666 21227 702 21283
rect 758 21227 778 21283
rect 164 21202 778 21227
rect 164 21146 242 21202
rect 298 21146 334 21202
rect 390 21146 426 21202
rect 482 21146 518 21202
rect 574 21146 610 21202
rect 666 21146 702 21202
rect 758 21146 778 21202
rect 164 21121 778 21146
rect 1009 23686 1167 23690
rect 1065 23630 1111 23686
rect 1009 23606 1167 23630
rect 1065 23550 1111 23606
rect 1009 23526 1167 23550
rect 1065 23470 1111 23526
rect 1009 23446 1167 23470
rect 1065 23390 1111 23446
rect 1009 23366 1167 23390
rect 1065 23310 1111 23366
rect 1009 23286 1167 23310
rect 1065 23230 1111 23286
rect 1009 23206 1167 23230
rect 1065 23150 1111 23206
rect 1009 23126 1167 23150
rect 1065 23070 1111 23126
rect 1009 23046 1167 23070
rect 1065 22990 1111 23046
rect 1009 22966 1167 22990
rect 1065 22910 1111 22966
rect 1009 22886 1167 22910
rect 1065 22830 1111 22886
rect 1009 22806 1167 22830
rect 1065 22750 1111 22806
rect 1009 22726 1167 22750
rect 1065 22670 1111 22726
rect 1009 22646 1167 22670
rect 1065 22590 1111 22646
rect 1009 22566 1167 22590
rect 1065 22510 1111 22566
rect 1009 22486 1167 22510
rect 1065 22430 1111 22486
rect 1009 22406 1167 22430
rect 1065 22350 1111 22406
rect 1009 22326 1167 22350
rect 1065 22270 1111 22326
rect 1009 22245 1167 22270
rect 1065 22189 1111 22245
rect 1009 22164 1167 22189
rect 1065 22108 1111 22164
rect 1009 22083 1167 22108
rect 1065 22027 1111 22083
rect 1009 22002 1167 22027
rect 1065 21946 1111 22002
rect 1009 21921 1167 21946
rect 1065 21865 1111 21921
rect 1009 21840 1167 21865
rect 1065 21784 1111 21840
rect 1009 21759 1167 21784
rect 1065 21703 1111 21759
rect 1009 21678 1167 21703
rect 1065 21622 1111 21678
rect 1009 21597 1167 21622
rect 1065 21541 1111 21597
rect 1009 21516 1167 21541
rect 1065 21460 1111 21516
rect 1009 21435 1167 21460
rect 1065 21379 1111 21435
rect 1009 21354 1167 21379
rect 1065 21298 1111 21354
rect 1009 21273 1167 21298
rect 1065 21217 1111 21273
rect 1009 21192 1167 21217
rect 1065 21136 1111 21192
rect 1009 21127 1167 21136
rect 1497 23686 1671 23695
rect 1985 23690 2175 23695
rect 1553 23630 1615 23686
rect 1497 23606 1671 23630
rect 1553 23550 1615 23606
rect 1497 23526 1671 23550
rect 1553 23470 1615 23526
rect 1497 23446 1671 23470
rect 1553 23390 1615 23446
rect 1497 23366 1671 23390
rect 1553 23310 1615 23366
rect 1497 23286 1671 23310
rect 1553 23230 1615 23286
rect 1497 23206 1671 23230
rect 1553 23150 1615 23206
rect 1497 23126 1671 23150
rect 1553 23070 1615 23126
rect 1497 23046 1671 23070
rect 1553 22990 1615 23046
rect 1497 22966 1671 22990
rect 1553 22910 1615 22966
rect 1497 22886 1671 22910
rect 1553 22830 1615 22886
rect 1497 22806 1671 22830
rect 1553 22750 1615 22806
rect 1497 22726 1671 22750
rect 1553 22670 1615 22726
rect 1497 22646 1671 22670
rect 1553 22590 1615 22646
rect 1497 22566 1671 22590
rect 1553 22510 1615 22566
rect 1497 22486 1671 22510
rect 1553 22430 1615 22486
rect 1497 22406 1671 22430
rect 1553 22350 1615 22406
rect 1497 22326 1671 22350
rect 1553 22270 1615 22326
rect 1497 22245 1671 22270
rect 1553 22189 1615 22245
rect 1497 22164 1671 22189
rect 1553 22108 1615 22164
rect 1497 22083 1671 22108
rect 1553 22027 1615 22083
rect 1497 22002 1671 22027
rect 1553 21946 1615 22002
rect 1497 21921 1671 21946
rect 1553 21865 1615 21921
rect 1497 21840 1671 21865
rect 1553 21784 1615 21840
rect 1497 21759 1671 21784
rect 1553 21703 1615 21759
rect 1497 21678 1671 21703
rect 1553 21622 1615 21678
rect 1497 21597 1671 21622
rect 1553 21541 1615 21597
rect 1497 21516 1671 21541
rect 1553 21460 1615 21516
rect 1497 21435 1671 21460
rect 1553 21379 1615 21435
rect 1497 21354 1671 21379
rect 1553 21298 1615 21354
rect 1497 21273 1671 21298
rect 1553 21217 1615 21273
rect 1497 21192 1671 21217
rect 1553 21136 1615 21192
rect 1497 21127 1671 21136
rect 1993 23686 2167 23690
rect 2049 23630 2111 23686
rect 1993 23606 2167 23630
rect 2049 23550 2111 23606
rect 1993 23526 2167 23550
rect 2049 23470 2111 23526
rect 1993 23446 2167 23470
rect 2049 23390 2111 23446
rect 1993 23366 2167 23390
rect 2049 23310 2111 23366
rect 1993 23286 2167 23310
rect 2049 23230 2111 23286
rect 1993 23206 2167 23230
rect 2049 23150 2111 23206
rect 1993 23126 2167 23150
rect 2049 23070 2111 23126
rect 1993 23046 2167 23070
rect 2049 22990 2111 23046
rect 1993 22966 2167 22990
rect 2049 22910 2111 22966
rect 1993 22886 2167 22910
rect 2049 22830 2111 22886
rect 1993 22806 2167 22830
rect 2049 22750 2111 22806
rect 1993 22726 2167 22750
rect 2049 22670 2111 22726
rect 1993 22646 2167 22670
rect 2049 22590 2111 22646
rect 1993 22566 2167 22590
rect 2049 22510 2111 22566
rect 1993 22486 2167 22510
rect 2049 22430 2111 22486
rect 1993 22406 2167 22430
rect 2049 22350 2111 22406
rect 1993 22326 2167 22350
rect 2049 22270 2111 22326
rect 1993 22245 2167 22270
rect 2049 22189 2111 22245
rect 1993 22164 2167 22189
rect 2049 22108 2111 22164
rect 1993 22083 2167 22108
rect 2049 22027 2111 22083
rect 1993 22002 2167 22027
rect 2049 21946 2111 22002
rect 1993 21921 2167 21946
rect 2049 21865 2111 21921
rect 1993 21840 2167 21865
rect 2049 21784 2111 21840
rect 1993 21759 2167 21784
rect 2049 21703 2111 21759
rect 1993 21678 2167 21703
rect 2049 21622 2111 21678
rect 1993 21597 2167 21622
rect 2049 21541 2111 21597
rect 1993 21516 2167 21541
rect 2049 21460 2111 21516
rect 1993 21435 2167 21460
rect 2049 21379 2111 21435
rect 1993 21354 2167 21379
rect 2049 21298 2111 21354
rect 1993 21273 2167 21298
rect 2049 21217 2111 21273
rect 1993 21192 2167 21217
rect 2049 21136 2111 21192
rect 1993 21127 2167 21136
rect 2489 23686 2663 23695
rect 2977 23690 3167 23695
rect 2545 23630 2607 23686
rect 2489 23606 2663 23630
rect 2545 23550 2607 23606
rect 2489 23526 2663 23550
rect 2545 23470 2607 23526
rect 2489 23446 2663 23470
rect 2545 23390 2607 23446
rect 2489 23366 2663 23390
rect 2545 23310 2607 23366
rect 2489 23286 2663 23310
rect 2545 23230 2607 23286
rect 2489 23206 2663 23230
rect 2545 23150 2607 23206
rect 2489 23126 2663 23150
rect 2545 23070 2607 23126
rect 2489 23046 2663 23070
rect 2545 22990 2607 23046
rect 2489 22966 2663 22990
rect 2545 22910 2607 22966
rect 2489 22886 2663 22910
rect 2545 22830 2607 22886
rect 2489 22806 2663 22830
rect 2545 22750 2607 22806
rect 2489 22726 2663 22750
rect 2545 22670 2607 22726
rect 2489 22646 2663 22670
rect 2545 22590 2607 22646
rect 2489 22566 2663 22590
rect 2545 22510 2607 22566
rect 2489 22486 2663 22510
rect 2545 22430 2607 22486
rect 2489 22406 2663 22430
rect 2545 22350 2607 22406
rect 2489 22326 2663 22350
rect 2545 22270 2607 22326
rect 2489 22245 2663 22270
rect 2545 22189 2607 22245
rect 2489 22164 2663 22189
rect 2545 22108 2607 22164
rect 2489 22083 2663 22108
rect 2545 22027 2607 22083
rect 2489 22002 2663 22027
rect 2545 21946 2607 22002
rect 2489 21921 2663 21946
rect 2545 21865 2607 21921
rect 2489 21840 2663 21865
rect 2545 21784 2607 21840
rect 2489 21759 2663 21784
rect 2545 21703 2607 21759
rect 2489 21678 2663 21703
rect 2545 21622 2607 21678
rect 2489 21597 2663 21622
rect 2545 21541 2607 21597
rect 2489 21516 2663 21541
rect 2545 21460 2607 21516
rect 2489 21435 2663 21460
rect 2545 21379 2607 21435
rect 2489 21354 2663 21379
rect 2545 21298 2607 21354
rect 2489 21273 2663 21298
rect 2545 21217 2607 21273
rect 2489 21192 2663 21217
rect 2545 21136 2607 21192
rect 2489 21127 2663 21136
rect 2985 23686 3159 23690
rect 3041 23630 3103 23686
rect 2985 23606 3159 23630
rect 3041 23550 3103 23606
rect 2985 23526 3159 23550
rect 3041 23470 3103 23526
rect 2985 23446 3159 23470
rect 3041 23390 3103 23446
rect 2985 23366 3159 23390
rect 3041 23310 3103 23366
rect 2985 23286 3159 23310
rect 3041 23230 3103 23286
rect 2985 23206 3159 23230
rect 3041 23150 3103 23206
rect 2985 23126 3159 23150
rect 3041 23070 3103 23126
rect 2985 23046 3159 23070
rect 3041 22990 3103 23046
rect 2985 22966 3159 22990
rect 3041 22910 3103 22966
rect 2985 22886 3159 22910
rect 3041 22830 3103 22886
rect 2985 22806 3159 22830
rect 3041 22750 3103 22806
rect 2985 22726 3159 22750
rect 3041 22670 3103 22726
rect 2985 22646 3159 22670
rect 3041 22590 3103 22646
rect 2985 22566 3159 22590
rect 3041 22510 3103 22566
rect 2985 22486 3159 22510
rect 3041 22430 3103 22486
rect 2985 22406 3159 22430
rect 3041 22350 3103 22406
rect 2985 22326 3159 22350
rect 3041 22270 3103 22326
rect 2985 22245 3159 22270
rect 3041 22189 3103 22245
rect 2985 22164 3159 22189
rect 3041 22108 3103 22164
rect 2985 22083 3159 22108
rect 3041 22027 3103 22083
rect 2985 22002 3159 22027
rect 3041 21946 3103 22002
rect 2985 21921 3159 21946
rect 3041 21865 3103 21921
rect 2985 21840 3159 21865
rect 3041 21784 3103 21840
rect 2985 21759 3159 21784
rect 3041 21703 3103 21759
rect 2985 21678 3159 21703
rect 3041 21622 3103 21678
rect 2985 21597 3159 21622
rect 3041 21541 3103 21597
rect 2985 21516 3159 21541
rect 3041 21460 3103 21516
rect 2985 21435 3159 21460
rect 3041 21379 3103 21435
rect 2985 21354 3159 21379
rect 3041 21298 3103 21354
rect 2985 21273 3159 21298
rect 3041 21217 3103 21273
rect 2985 21192 3159 21217
rect 3041 21136 3103 21192
rect 2985 21127 3159 21136
rect 3481 23686 3655 23695
rect 3969 23690 4159 23695
rect 3537 23630 3599 23686
rect 3481 23606 3655 23630
rect 3537 23550 3599 23606
rect 3481 23526 3655 23550
rect 3537 23470 3599 23526
rect 3481 23446 3655 23470
rect 3537 23390 3599 23446
rect 3481 23366 3655 23390
rect 3537 23310 3599 23366
rect 3481 23286 3655 23310
rect 3537 23230 3599 23286
rect 3481 23206 3655 23230
rect 3537 23150 3599 23206
rect 3481 23126 3655 23150
rect 3537 23070 3599 23126
rect 3481 23046 3655 23070
rect 3537 22990 3599 23046
rect 3481 22966 3655 22990
rect 3537 22910 3599 22966
rect 3481 22886 3655 22910
rect 3537 22830 3599 22886
rect 3481 22806 3655 22830
rect 3537 22750 3599 22806
rect 3481 22726 3655 22750
rect 3537 22670 3599 22726
rect 3481 22646 3655 22670
rect 3537 22590 3599 22646
rect 3481 22566 3655 22590
rect 3537 22510 3599 22566
rect 3481 22486 3655 22510
rect 3537 22430 3599 22486
rect 3481 22406 3655 22430
rect 3537 22350 3599 22406
rect 3481 22326 3655 22350
rect 3537 22270 3599 22326
rect 3481 22245 3655 22270
rect 3537 22189 3599 22245
rect 3481 22164 3655 22189
rect 3537 22108 3599 22164
rect 3481 22083 3655 22108
rect 3537 22027 3599 22083
rect 3481 22002 3655 22027
rect 3537 21946 3599 22002
rect 3481 21921 3655 21946
rect 3537 21865 3599 21921
rect 3481 21840 3655 21865
rect 3537 21784 3599 21840
rect 3481 21759 3655 21784
rect 3537 21703 3599 21759
rect 3481 21678 3655 21703
rect 3537 21622 3599 21678
rect 3481 21597 3655 21622
rect 3537 21541 3599 21597
rect 3481 21516 3655 21541
rect 3537 21460 3599 21516
rect 3481 21435 3655 21460
rect 3537 21379 3599 21435
rect 3481 21354 3655 21379
rect 3537 21298 3599 21354
rect 3481 21273 3655 21298
rect 3537 21217 3599 21273
rect 3481 21192 3655 21217
rect 3537 21136 3599 21192
rect 3481 21127 3655 21136
rect 3977 23686 4151 23690
rect 4033 23630 4095 23686
rect 3977 23606 4151 23630
rect 4033 23550 4095 23606
rect 3977 23526 4151 23550
rect 4033 23470 4095 23526
rect 3977 23446 4151 23470
rect 4033 23390 4095 23446
rect 3977 23366 4151 23390
rect 4033 23310 4095 23366
rect 3977 23286 4151 23310
rect 4033 23230 4095 23286
rect 3977 23206 4151 23230
rect 4033 23150 4095 23206
rect 3977 23126 4151 23150
rect 4033 23070 4095 23126
rect 3977 23046 4151 23070
rect 4033 22990 4095 23046
rect 3977 22966 4151 22990
rect 4033 22910 4095 22966
rect 3977 22886 4151 22910
rect 4033 22830 4095 22886
rect 3977 22806 4151 22830
rect 4033 22750 4095 22806
rect 3977 22726 4151 22750
rect 4033 22670 4095 22726
rect 3977 22646 4151 22670
rect 4033 22590 4095 22646
rect 3977 22566 4151 22590
rect 4033 22510 4095 22566
rect 3977 22486 4151 22510
rect 4033 22430 4095 22486
rect 3977 22406 4151 22430
rect 4033 22350 4095 22406
rect 3977 22326 4151 22350
rect 4033 22270 4095 22326
rect 3977 22245 4151 22270
rect 4033 22189 4095 22245
rect 3977 22164 4151 22189
rect 4033 22108 4095 22164
rect 3977 22083 4151 22108
rect 4033 22027 4095 22083
rect 3977 22002 4151 22027
rect 4033 21946 4095 22002
rect 3977 21921 4151 21946
rect 4033 21865 4095 21921
rect 3977 21840 4151 21865
rect 4033 21784 4095 21840
rect 3977 21759 4151 21784
rect 4033 21703 4095 21759
rect 3977 21678 4151 21703
rect 4033 21622 4095 21678
rect 3977 21597 4151 21622
rect 4033 21541 4095 21597
rect 3977 21516 4151 21541
rect 4033 21460 4095 21516
rect 3977 21435 4151 21460
rect 4033 21379 4095 21435
rect 3977 21354 4151 21379
rect 4033 21298 4095 21354
rect 3977 21273 4151 21298
rect 4033 21217 4095 21273
rect 3977 21192 4151 21217
rect 4033 21136 4095 21192
rect 3977 21127 4151 21136
rect 4473 23686 4647 23695
rect 4961 23690 5151 23695
rect 4529 23630 4591 23686
rect 4473 23606 4647 23630
rect 4529 23550 4591 23606
rect 4473 23526 4647 23550
rect 4529 23470 4591 23526
rect 4473 23446 4647 23470
rect 4529 23390 4591 23446
rect 4473 23366 4647 23390
rect 4529 23310 4591 23366
rect 4473 23286 4647 23310
rect 4529 23230 4591 23286
rect 4473 23206 4647 23230
rect 4529 23150 4591 23206
rect 4473 23126 4647 23150
rect 4529 23070 4591 23126
rect 4473 23046 4647 23070
rect 4529 22990 4591 23046
rect 4473 22966 4647 22990
rect 4529 22910 4591 22966
rect 4473 22886 4647 22910
rect 4529 22830 4591 22886
rect 4473 22806 4647 22830
rect 4529 22750 4591 22806
rect 4473 22726 4647 22750
rect 4529 22670 4591 22726
rect 4473 22646 4647 22670
rect 4529 22590 4591 22646
rect 4473 22566 4647 22590
rect 4529 22510 4591 22566
rect 4473 22486 4647 22510
rect 4529 22430 4591 22486
rect 4473 22406 4647 22430
rect 4529 22350 4591 22406
rect 4473 22326 4647 22350
rect 4529 22270 4591 22326
rect 4473 22245 4647 22270
rect 4529 22189 4591 22245
rect 4473 22164 4647 22189
rect 4529 22108 4591 22164
rect 4473 22083 4647 22108
rect 4529 22027 4591 22083
rect 4473 22002 4647 22027
rect 4529 21946 4591 22002
rect 4473 21921 4647 21946
rect 4529 21865 4591 21921
rect 4473 21840 4647 21865
rect 4529 21784 4591 21840
rect 4473 21759 4647 21784
rect 4529 21703 4591 21759
rect 4473 21678 4647 21703
rect 4529 21622 4591 21678
rect 4473 21597 4647 21622
rect 4529 21541 4591 21597
rect 4473 21516 4647 21541
rect 4529 21460 4591 21516
rect 4473 21435 4647 21460
rect 4529 21379 4591 21435
rect 4473 21354 4647 21379
rect 4529 21298 4591 21354
rect 4473 21273 4647 21298
rect 4529 21217 4591 21273
rect 4473 21192 4647 21217
rect 4529 21136 4591 21192
rect 4473 21127 4647 21136
rect 4969 23686 5143 23690
rect 5025 23630 5087 23686
rect 4969 23606 5143 23630
rect 5025 23550 5087 23606
rect 4969 23526 5143 23550
rect 5025 23470 5087 23526
rect 4969 23446 5143 23470
rect 5025 23390 5087 23446
rect 4969 23366 5143 23390
rect 5025 23310 5087 23366
rect 4969 23286 5143 23310
rect 5025 23230 5087 23286
rect 4969 23206 5143 23230
rect 5025 23150 5087 23206
rect 4969 23126 5143 23150
rect 5025 23070 5087 23126
rect 4969 23046 5143 23070
rect 5025 22990 5087 23046
rect 4969 22966 5143 22990
rect 5025 22910 5087 22966
rect 4969 22886 5143 22910
rect 5025 22830 5087 22886
rect 4969 22806 5143 22830
rect 5025 22750 5087 22806
rect 4969 22726 5143 22750
rect 5025 22670 5087 22726
rect 4969 22646 5143 22670
rect 5025 22590 5087 22646
rect 4969 22566 5143 22590
rect 5025 22510 5087 22566
rect 4969 22486 5143 22510
rect 5025 22430 5087 22486
rect 4969 22406 5143 22430
rect 5025 22350 5087 22406
rect 4969 22326 5143 22350
rect 5025 22270 5087 22326
rect 4969 22245 5143 22270
rect 5025 22189 5087 22245
rect 4969 22164 5143 22189
rect 5025 22108 5087 22164
rect 4969 22083 5143 22108
rect 5025 22027 5087 22083
rect 4969 22002 5143 22027
rect 5025 21946 5087 22002
rect 4969 21921 5143 21946
rect 5025 21865 5087 21921
rect 4969 21840 5143 21865
rect 5025 21784 5087 21840
rect 4969 21759 5143 21784
rect 5025 21703 5087 21759
rect 4969 21678 5143 21703
rect 5025 21622 5087 21678
rect 4969 21597 5143 21622
rect 5025 21541 5087 21597
rect 4969 21516 5143 21541
rect 5025 21460 5087 21516
rect 4969 21435 5143 21460
rect 5025 21379 5087 21435
rect 4969 21354 5143 21379
rect 5025 21298 5087 21354
rect 4969 21273 5143 21298
rect 5025 21217 5087 21273
rect 4969 21192 5143 21217
rect 5025 21136 5087 21192
rect 4969 21127 5143 21136
rect 5465 23686 5639 23695
rect 5953 23690 6143 23695
rect 5521 23630 5583 23686
rect 5465 23606 5639 23630
rect 5521 23550 5583 23606
rect 5465 23526 5639 23550
rect 5521 23470 5583 23526
rect 5465 23446 5639 23470
rect 5521 23390 5583 23446
rect 5465 23366 5639 23390
rect 5521 23310 5583 23366
rect 5465 23286 5639 23310
rect 5521 23230 5583 23286
rect 5465 23206 5639 23230
rect 5521 23150 5583 23206
rect 5465 23126 5639 23150
rect 5521 23070 5583 23126
rect 5465 23046 5639 23070
rect 5521 22990 5583 23046
rect 5465 22966 5639 22990
rect 5521 22910 5583 22966
rect 5465 22886 5639 22910
rect 5521 22830 5583 22886
rect 5465 22806 5639 22830
rect 5521 22750 5583 22806
rect 5465 22726 5639 22750
rect 5521 22670 5583 22726
rect 5465 22646 5639 22670
rect 5521 22590 5583 22646
rect 5465 22566 5639 22590
rect 5521 22510 5583 22566
rect 5465 22486 5639 22510
rect 5521 22430 5583 22486
rect 5465 22406 5639 22430
rect 5521 22350 5583 22406
rect 5465 22326 5639 22350
rect 5521 22270 5583 22326
rect 5465 22245 5639 22270
rect 5521 22189 5583 22245
rect 5465 22164 5639 22189
rect 5521 22108 5583 22164
rect 5465 22083 5639 22108
rect 5521 22027 5583 22083
rect 5465 22002 5639 22027
rect 5521 21946 5583 22002
rect 5465 21921 5639 21946
rect 5521 21865 5583 21921
rect 5465 21840 5639 21865
rect 5521 21784 5583 21840
rect 5465 21759 5639 21784
rect 5521 21703 5583 21759
rect 5465 21678 5639 21703
rect 5521 21622 5583 21678
rect 5465 21597 5639 21622
rect 5521 21541 5583 21597
rect 5465 21516 5639 21541
rect 5521 21460 5583 21516
rect 5465 21435 5639 21460
rect 5521 21379 5583 21435
rect 5465 21354 5639 21379
rect 5521 21298 5583 21354
rect 5465 21273 5639 21298
rect 5521 21217 5583 21273
rect 5465 21192 5639 21217
rect 5521 21136 5583 21192
rect 5465 21127 5639 21136
rect 5961 23686 6135 23690
rect 6017 23630 6079 23686
rect 5961 23606 6135 23630
rect 6017 23550 6079 23606
rect 5961 23526 6135 23550
rect 6017 23470 6079 23526
rect 5961 23446 6135 23470
rect 6017 23390 6079 23446
rect 5961 23366 6135 23390
rect 6017 23310 6079 23366
rect 5961 23286 6135 23310
rect 6017 23230 6079 23286
rect 5961 23206 6135 23230
rect 6017 23150 6079 23206
rect 5961 23126 6135 23150
rect 6017 23070 6079 23126
rect 5961 23046 6135 23070
rect 6017 22990 6079 23046
rect 5961 22966 6135 22990
rect 6017 22910 6079 22966
rect 5961 22886 6135 22910
rect 6017 22830 6079 22886
rect 5961 22806 6135 22830
rect 6017 22750 6079 22806
rect 5961 22726 6135 22750
rect 6017 22670 6079 22726
rect 5961 22646 6135 22670
rect 6017 22590 6079 22646
rect 5961 22566 6135 22590
rect 6017 22510 6079 22566
rect 5961 22486 6135 22510
rect 6017 22430 6079 22486
rect 5961 22406 6135 22430
rect 6017 22350 6079 22406
rect 5961 22326 6135 22350
rect 6017 22270 6079 22326
rect 5961 22245 6135 22270
rect 6017 22189 6079 22245
rect 5961 22164 6135 22189
rect 6017 22108 6079 22164
rect 5961 22083 6135 22108
rect 6017 22027 6079 22083
rect 5961 22002 6135 22027
rect 6017 21946 6079 22002
rect 5961 21921 6135 21946
rect 6017 21865 6079 21921
rect 5961 21840 6135 21865
rect 6017 21784 6079 21840
rect 5961 21759 6135 21784
rect 6017 21703 6079 21759
rect 5961 21678 6135 21703
rect 6017 21622 6079 21678
rect 5961 21597 6135 21622
rect 6017 21541 6079 21597
rect 5961 21516 6135 21541
rect 6017 21460 6079 21516
rect 5961 21435 6135 21460
rect 6017 21379 6079 21435
rect 5961 21354 6135 21379
rect 6017 21298 6079 21354
rect 5961 21273 6135 21298
rect 6017 21217 6079 21273
rect 5961 21192 6135 21217
rect 6017 21136 6079 21192
rect 5961 21127 6135 21136
rect 6457 23686 6631 23695
rect 6945 23690 7135 23695
rect 6513 23630 6575 23686
rect 6457 23606 6631 23630
rect 6513 23550 6575 23606
rect 6457 23526 6631 23550
rect 6513 23470 6575 23526
rect 6457 23446 6631 23470
rect 6513 23390 6575 23446
rect 6457 23366 6631 23390
rect 6513 23310 6575 23366
rect 6457 23286 6631 23310
rect 6513 23230 6575 23286
rect 6457 23206 6631 23230
rect 6513 23150 6575 23206
rect 6457 23126 6631 23150
rect 6513 23070 6575 23126
rect 6457 23046 6631 23070
rect 6513 22990 6575 23046
rect 6457 22966 6631 22990
rect 6513 22910 6575 22966
rect 6457 22886 6631 22910
rect 6513 22830 6575 22886
rect 6457 22806 6631 22830
rect 6513 22750 6575 22806
rect 6457 22726 6631 22750
rect 6513 22670 6575 22726
rect 6457 22646 6631 22670
rect 6513 22590 6575 22646
rect 6457 22566 6631 22590
rect 6513 22510 6575 22566
rect 6457 22486 6631 22510
rect 6513 22430 6575 22486
rect 6457 22406 6631 22430
rect 6513 22350 6575 22406
rect 6457 22326 6631 22350
rect 6513 22270 6575 22326
rect 6457 22245 6631 22270
rect 6513 22189 6575 22245
rect 6457 22164 6631 22189
rect 6513 22108 6575 22164
rect 6457 22083 6631 22108
rect 6513 22027 6575 22083
rect 6457 22002 6631 22027
rect 6513 21946 6575 22002
rect 6457 21921 6631 21946
rect 6513 21865 6575 21921
rect 6457 21840 6631 21865
rect 6513 21784 6575 21840
rect 6457 21759 6631 21784
rect 6513 21703 6575 21759
rect 6457 21678 6631 21703
rect 6513 21622 6575 21678
rect 6457 21597 6631 21622
rect 6513 21541 6575 21597
rect 6457 21516 6631 21541
rect 6513 21460 6575 21516
rect 6457 21435 6631 21460
rect 6513 21379 6575 21435
rect 6457 21354 6631 21379
rect 6513 21298 6575 21354
rect 6457 21273 6631 21298
rect 6513 21217 6575 21273
rect 6457 21192 6631 21217
rect 6513 21136 6575 21192
rect 6457 21127 6631 21136
rect 6953 23686 7127 23690
rect 7009 23630 7071 23686
rect 6953 23606 7127 23630
rect 7009 23550 7071 23606
rect 6953 23526 7127 23550
rect 7009 23470 7071 23526
rect 6953 23446 7127 23470
rect 7009 23390 7071 23446
rect 6953 23366 7127 23390
rect 7009 23310 7071 23366
rect 6953 23286 7127 23310
rect 7009 23230 7071 23286
rect 6953 23206 7127 23230
rect 7009 23150 7071 23206
rect 6953 23126 7127 23150
rect 7009 23070 7071 23126
rect 6953 23046 7127 23070
rect 7009 22990 7071 23046
rect 6953 22966 7127 22990
rect 7009 22910 7071 22966
rect 6953 22886 7127 22910
rect 7009 22830 7071 22886
rect 6953 22806 7127 22830
rect 7009 22750 7071 22806
rect 6953 22726 7127 22750
rect 7009 22670 7071 22726
rect 6953 22646 7127 22670
rect 7009 22590 7071 22646
rect 6953 22566 7127 22590
rect 7009 22510 7071 22566
rect 6953 22486 7127 22510
rect 7009 22430 7071 22486
rect 6953 22406 7127 22430
rect 7009 22350 7071 22406
rect 6953 22326 7127 22350
rect 7009 22270 7071 22326
rect 6953 22245 7127 22270
rect 7009 22189 7071 22245
rect 6953 22164 7127 22189
rect 7009 22108 7071 22164
rect 6953 22083 7127 22108
rect 7009 22027 7071 22083
rect 6953 22002 7127 22027
rect 7009 21946 7071 22002
rect 6953 21921 7127 21946
rect 7009 21865 7071 21921
rect 6953 21840 7127 21865
rect 7009 21784 7071 21840
rect 6953 21759 7127 21784
rect 7009 21703 7071 21759
rect 6953 21678 7127 21703
rect 7009 21622 7071 21678
rect 6953 21597 7127 21622
rect 7009 21541 7071 21597
rect 6953 21516 7127 21541
rect 7009 21460 7071 21516
rect 6953 21435 7127 21460
rect 7009 21379 7071 21435
rect 6953 21354 7127 21379
rect 7009 21298 7071 21354
rect 6953 21273 7127 21298
rect 7009 21217 7071 21273
rect 6953 21192 7127 21217
rect 7009 21136 7071 21192
rect 6953 21127 7127 21136
rect 7449 23686 7623 23695
rect 7937 23690 8127 23695
rect 7505 23630 7567 23686
rect 7449 23606 7623 23630
rect 7505 23550 7567 23606
rect 7449 23526 7623 23550
rect 7505 23470 7567 23526
rect 7449 23446 7623 23470
rect 7505 23390 7567 23446
rect 7449 23366 7623 23390
rect 7505 23310 7567 23366
rect 7449 23286 7623 23310
rect 7505 23230 7567 23286
rect 7449 23206 7623 23230
rect 7505 23150 7567 23206
rect 7449 23126 7623 23150
rect 7505 23070 7567 23126
rect 7449 23046 7623 23070
rect 7505 22990 7567 23046
rect 7449 22966 7623 22990
rect 7505 22910 7567 22966
rect 7449 22886 7623 22910
rect 7505 22830 7567 22886
rect 7449 22806 7623 22830
rect 7505 22750 7567 22806
rect 7449 22726 7623 22750
rect 7505 22670 7567 22726
rect 7449 22646 7623 22670
rect 7505 22590 7567 22646
rect 7449 22566 7623 22590
rect 7505 22510 7567 22566
rect 7449 22486 7623 22510
rect 7505 22430 7567 22486
rect 7449 22406 7623 22430
rect 7505 22350 7567 22406
rect 7449 22326 7623 22350
rect 7505 22270 7567 22326
rect 7449 22245 7623 22270
rect 7505 22189 7567 22245
rect 7449 22164 7623 22189
rect 7505 22108 7567 22164
rect 7449 22083 7623 22108
rect 7505 22027 7567 22083
rect 7449 22002 7623 22027
rect 7505 21946 7567 22002
rect 7449 21921 7623 21946
rect 7505 21865 7567 21921
rect 7449 21840 7623 21865
rect 7505 21784 7567 21840
rect 7449 21759 7623 21784
rect 7505 21703 7567 21759
rect 7449 21678 7623 21703
rect 7505 21622 7567 21678
rect 7449 21597 7623 21622
rect 7505 21541 7567 21597
rect 7449 21516 7623 21541
rect 7505 21460 7567 21516
rect 7449 21435 7623 21460
rect 7505 21379 7567 21435
rect 7449 21354 7623 21379
rect 7505 21298 7567 21354
rect 7449 21273 7623 21298
rect 7505 21217 7567 21273
rect 7449 21192 7623 21217
rect 7505 21136 7567 21192
rect 7449 21127 7623 21136
rect 7945 23686 8119 23690
rect 8001 23630 8063 23686
rect 7945 23606 8119 23630
rect 8001 23550 8063 23606
rect 7945 23526 8119 23550
rect 8001 23470 8063 23526
rect 7945 23446 8119 23470
rect 8001 23390 8063 23446
rect 7945 23366 8119 23390
rect 8001 23310 8063 23366
rect 7945 23286 8119 23310
rect 8001 23230 8063 23286
rect 7945 23206 8119 23230
rect 8001 23150 8063 23206
rect 7945 23126 8119 23150
rect 8001 23070 8063 23126
rect 7945 23046 8119 23070
rect 8001 22990 8063 23046
rect 7945 22966 8119 22990
rect 8001 22910 8063 22966
rect 7945 22886 8119 22910
rect 8001 22830 8063 22886
rect 7945 22806 8119 22830
rect 8001 22750 8063 22806
rect 7945 22726 8119 22750
rect 8001 22670 8063 22726
rect 7945 22646 8119 22670
rect 8001 22590 8063 22646
rect 7945 22566 8119 22590
rect 8001 22510 8063 22566
rect 7945 22486 8119 22510
rect 8001 22430 8063 22486
rect 7945 22406 8119 22430
rect 8001 22350 8063 22406
rect 7945 22326 8119 22350
rect 8001 22270 8063 22326
rect 7945 22245 8119 22270
rect 8001 22189 8063 22245
rect 7945 22164 8119 22189
rect 8001 22108 8063 22164
rect 7945 22083 8119 22108
rect 8001 22027 8063 22083
rect 7945 22002 8119 22027
rect 8001 21946 8063 22002
rect 7945 21921 8119 21946
rect 8001 21865 8063 21921
rect 7945 21840 8119 21865
rect 8001 21784 8063 21840
rect 7945 21759 8119 21784
rect 8001 21703 8063 21759
rect 7945 21678 8119 21703
rect 8001 21622 8063 21678
rect 7945 21597 8119 21622
rect 8001 21541 8063 21597
rect 7945 21516 8119 21541
rect 8001 21460 8063 21516
rect 7945 21435 8119 21460
rect 8001 21379 8063 21435
rect 7945 21354 8119 21379
rect 8001 21298 8063 21354
rect 7945 21273 8119 21298
rect 8001 21217 8063 21273
rect 7945 21192 8119 21217
rect 8001 21136 8063 21192
rect 7945 21127 8119 21136
rect 8441 23686 8615 23695
rect 8929 23690 9119 23695
rect 8497 23630 8559 23686
rect 8441 23606 8615 23630
rect 8497 23550 8559 23606
rect 8441 23526 8615 23550
rect 8497 23470 8559 23526
rect 8441 23446 8615 23470
rect 8497 23390 8559 23446
rect 8441 23366 8615 23390
rect 8497 23310 8559 23366
rect 8441 23286 8615 23310
rect 8497 23230 8559 23286
rect 8441 23206 8615 23230
rect 8497 23150 8559 23206
rect 8441 23126 8615 23150
rect 8497 23070 8559 23126
rect 8441 23046 8615 23070
rect 8497 22990 8559 23046
rect 8441 22966 8615 22990
rect 8497 22910 8559 22966
rect 8441 22886 8615 22910
rect 8497 22830 8559 22886
rect 8441 22806 8615 22830
rect 8497 22750 8559 22806
rect 8441 22726 8615 22750
rect 8497 22670 8559 22726
rect 8441 22646 8615 22670
rect 8497 22590 8559 22646
rect 8441 22566 8615 22590
rect 8497 22510 8559 22566
rect 8441 22486 8615 22510
rect 8497 22430 8559 22486
rect 8441 22406 8615 22430
rect 8497 22350 8559 22406
rect 8441 22326 8615 22350
rect 8497 22270 8559 22326
rect 8441 22245 8615 22270
rect 8497 22189 8559 22245
rect 8441 22164 8615 22189
rect 8497 22108 8559 22164
rect 8441 22083 8615 22108
rect 8497 22027 8559 22083
rect 8441 22002 8615 22027
rect 8497 21946 8559 22002
rect 8441 21921 8615 21946
rect 8497 21865 8559 21921
rect 8441 21840 8615 21865
rect 8497 21784 8559 21840
rect 8441 21759 8615 21784
rect 8497 21703 8559 21759
rect 8441 21678 8615 21703
rect 8497 21622 8559 21678
rect 8441 21597 8615 21622
rect 8497 21541 8559 21597
rect 8441 21516 8615 21541
rect 8497 21460 8559 21516
rect 8441 21435 8615 21460
rect 8497 21379 8559 21435
rect 8441 21354 8615 21379
rect 8497 21298 8559 21354
rect 8441 21273 8615 21298
rect 8497 21217 8559 21273
rect 8441 21192 8615 21217
rect 8497 21136 8559 21192
rect 8441 21127 8615 21136
rect 8937 23686 9111 23690
rect 8993 23630 9055 23686
rect 8937 23606 9111 23630
rect 8993 23550 9055 23606
rect 8937 23526 9111 23550
rect 8993 23470 9055 23526
rect 8937 23446 9111 23470
rect 8993 23390 9055 23446
rect 8937 23366 9111 23390
rect 8993 23310 9055 23366
rect 8937 23286 9111 23310
rect 8993 23230 9055 23286
rect 8937 23206 9111 23230
rect 8993 23150 9055 23206
rect 8937 23126 9111 23150
rect 8993 23070 9055 23126
rect 8937 23046 9111 23070
rect 8993 22990 9055 23046
rect 8937 22966 9111 22990
rect 8993 22910 9055 22966
rect 8937 22886 9111 22910
rect 8993 22830 9055 22886
rect 8937 22806 9111 22830
rect 8993 22750 9055 22806
rect 8937 22726 9111 22750
rect 8993 22670 9055 22726
rect 8937 22646 9111 22670
rect 8993 22590 9055 22646
rect 8937 22566 9111 22590
rect 8993 22510 9055 22566
rect 8937 22486 9111 22510
rect 8993 22430 9055 22486
rect 8937 22406 9111 22430
rect 8993 22350 9055 22406
rect 8937 22326 9111 22350
rect 8993 22270 9055 22326
rect 8937 22245 9111 22270
rect 8993 22189 9055 22245
rect 8937 22164 9111 22189
rect 8993 22108 9055 22164
rect 8937 22083 9111 22108
rect 8993 22027 9055 22083
rect 8937 22002 9111 22027
rect 8993 21946 9055 22002
rect 8937 21921 9111 21946
rect 8993 21865 9055 21921
rect 8937 21840 9111 21865
rect 8993 21784 9055 21840
rect 8937 21759 9111 21784
rect 8993 21703 9055 21759
rect 8937 21678 9111 21703
rect 8993 21622 9055 21678
rect 8937 21597 9111 21622
rect 8993 21541 9055 21597
rect 8937 21516 9111 21541
rect 8993 21460 9055 21516
rect 8937 21435 9111 21460
rect 8993 21379 9055 21435
rect 8937 21354 9111 21379
rect 8993 21298 9055 21354
rect 8937 21273 9111 21298
rect 8993 21217 9055 21273
rect 8937 21192 9111 21217
rect 8993 21136 9055 21192
rect 8937 21127 9111 21136
rect 9433 23686 9607 23695
rect 9921 23690 10111 23695
rect 9489 23630 9551 23686
rect 9433 23606 9607 23630
rect 9489 23550 9551 23606
rect 9433 23526 9607 23550
rect 9489 23470 9551 23526
rect 9433 23446 9607 23470
rect 9489 23390 9551 23446
rect 9433 23366 9607 23390
rect 9489 23310 9551 23366
rect 9433 23286 9607 23310
rect 9489 23230 9551 23286
rect 9433 23206 9607 23230
rect 9489 23150 9551 23206
rect 9433 23126 9607 23150
rect 9489 23070 9551 23126
rect 9433 23046 9607 23070
rect 9489 22990 9551 23046
rect 9433 22966 9607 22990
rect 9489 22910 9551 22966
rect 9433 22886 9607 22910
rect 9489 22830 9551 22886
rect 9433 22806 9607 22830
rect 9489 22750 9551 22806
rect 9433 22726 9607 22750
rect 9489 22670 9551 22726
rect 9433 22646 9607 22670
rect 9489 22590 9551 22646
rect 9433 22566 9607 22590
rect 9489 22510 9551 22566
rect 9433 22486 9607 22510
rect 9489 22430 9551 22486
rect 9433 22406 9607 22430
rect 9489 22350 9551 22406
rect 9433 22326 9607 22350
rect 9489 22270 9551 22326
rect 9433 22245 9607 22270
rect 9489 22189 9551 22245
rect 9433 22164 9607 22189
rect 9489 22108 9551 22164
rect 9433 22083 9607 22108
rect 9489 22027 9551 22083
rect 9433 22002 9607 22027
rect 9489 21946 9551 22002
rect 9433 21921 9607 21946
rect 9489 21865 9551 21921
rect 9433 21840 9607 21865
rect 9489 21784 9551 21840
rect 9433 21759 9607 21784
rect 9489 21703 9551 21759
rect 9433 21678 9607 21703
rect 9489 21622 9551 21678
rect 9433 21597 9607 21622
rect 9489 21541 9551 21597
rect 9433 21516 9607 21541
rect 9489 21460 9551 21516
rect 9433 21435 9607 21460
rect 9489 21379 9551 21435
rect 9433 21354 9607 21379
rect 9489 21298 9551 21354
rect 9433 21273 9607 21298
rect 9489 21217 9551 21273
rect 9433 21192 9607 21217
rect 9489 21136 9551 21192
rect 9433 21127 9607 21136
rect 9929 23686 10103 23690
rect 9985 23630 10047 23686
rect 9929 23606 10103 23630
rect 9985 23550 10047 23606
rect 9929 23526 10103 23550
rect 9985 23470 10047 23526
rect 9929 23446 10103 23470
rect 9985 23390 10047 23446
rect 9929 23366 10103 23390
rect 9985 23310 10047 23366
rect 9929 23286 10103 23310
rect 9985 23230 10047 23286
rect 9929 23206 10103 23230
rect 9985 23150 10047 23206
rect 9929 23126 10103 23150
rect 9985 23070 10047 23126
rect 9929 23046 10103 23070
rect 9985 22990 10047 23046
rect 9929 22966 10103 22990
rect 9985 22910 10047 22966
rect 9929 22886 10103 22910
rect 9985 22830 10047 22886
rect 9929 22806 10103 22830
rect 9985 22750 10047 22806
rect 9929 22726 10103 22750
rect 9985 22670 10047 22726
rect 9929 22646 10103 22670
rect 9985 22590 10047 22646
rect 9929 22566 10103 22590
rect 9985 22510 10047 22566
rect 9929 22486 10103 22510
rect 9985 22430 10047 22486
rect 9929 22406 10103 22430
rect 9985 22350 10047 22406
rect 9929 22326 10103 22350
rect 9985 22270 10047 22326
rect 9929 22245 10103 22270
rect 9985 22189 10047 22245
rect 9929 22164 10103 22189
rect 9985 22108 10047 22164
rect 9929 22083 10103 22108
rect 9985 22027 10047 22083
rect 9929 22002 10103 22027
rect 9985 21946 10047 22002
rect 9929 21921 10103 21946
rect 9985 21865 10047 21921
rect 9929 21840 10103 21865
rect 9985 21784 10047 21840
rect 9929 21759 10103 21784
rect 9985 21703 10047 21759
rect 9929 21678 10103 21703
rect 9985 21622 10047 21678
rect 9929 21597 10103 21622
rect 9985 21541 10047 21597
rect 9929 21516 10103 21541
rect 9985 21460 10047 21516
rect 9929 21435 10103 21460
rect 9985 21379 10047 21435
rect 9929 21354 10103 21379
rect 9985 21298 10047 21354
rect 9929 21273 10103 21298
rect 9985 21217 10047 21273
rect 9929 21192 10103 21217
rect 9985 21136 10047 21192
rect 9929 21127 10103 21136
rect 10425 23686 10599 23695
rect 10913 23690 11103 23695
rect 10481 23630 10543 23686
rect 10425 23606 10599 23630
rect 10481 23550 10543 23606
rect 10425 23526 10599 23550
rect 10481 23470 10543 23526
rect 10425 23446 10599 23470
rect 10481 23390 10543 23446
rect 10425 23366 10599 23390
rect 10481 23310 10543 23366
rect 10425 23286 10599 23310
rect 10481 23230 10543 23286
rect 10425 23206 10599 23230
rect 10481 23150 10543 23206
rect 10425 23126 10599 23150
rect 10481 23070 10543 23126
rect 10425 23046 10599 23070
rect 10481 22990 10543 23046
rect 10425 22966 10599 22990
rect 10481 22910 10543 22966
rect 10425 22886 10599 22910
rect 10481 22830 10543 22886
rect 10425 22806 10599 22830
rect 10481 22750 10543 22806
rect 10425 22726 10599 22750
rect 10481 22670 10543 22726
rect 10425 22646 10599 22670
rect 10481 22590 10543 22646
rect 10425 22566 10599 22590
rect 10481 22510 10543 22566
rect 10425 22486 10599 22510
rect 10481 22430 10543 22486
rect 10425 22406 10599 22430
rect 10481 22350 10543 22406
rect 10425 22326 10599 22350
rect 10481 22270 10543 22326
rect 10425 22245 10599 22270
rect 10481 22189 10543 22245
rect 10425 22164 10599 22189
rect 10481 22108 10543 22164
rect 10425 22083 10599 22108
rect 10481 22027 10543 22083
rect 10425 22002 10599 22027
rect 10481 21946 10543 22002
rect 10425 21921 10599 21946
rect 10481 21865 10543 21921
rect 10425 21840 10599 21865
rect 10481 21784 10543 21840
rect 10425 21759 10599 21784
rect 10481 21703 10543 21759
rect 10425 21678 10599 21703
rect 10481 21622 10543 21678
rect 10425 21597 10599 21622
rect 10481 21541 10543 21597
rect 10425 21516 10599 21541
rect 10481 21460 10543 21516
rect 10425 21435 10599 21460
rect 10481 21379 10543 21435
rect 10425 21354 10599 21379
rect 10481 21298 10543 21354
rect 10425 21273 10599 21298
rect 10481 21217 10543 21273
rect 10425 21192 10599 21217
rect 10481 21136 10543 21192
rect 10425 21127 10599 21136
rect 10921 23686 11095 23690
rect 10977 23630 11039 23686
rect 10921 23606 11095 23630
rect 10977 23550 11039 23606
rect 10921 23526 11095 23550
rect 10977 23470 11039 23526
rect 10921 23446 11095 23470
rect 10977 23390 11039 23446
rect 10921 23366 11095 23390
rect 10977 23310 11039 23366
rect 10921 23286 11095 23310
rect 10977 23230 11039 23286
rect 10921 23206 11095 23230
rect 10977 23150 11039 23206
rect 10921 23126 11095 23150
rect 10977 23070 11039 23126
rect 10921 23046 11095 23070
rect 10977 22990 11039 23046
rect 10921 22966 11095 22990
rect 10977 22910 11039 22966
rect 10921 22886 11095 22910
rect 10977 22830 11039 22886
rect 10921 22806 11095 22830
rect 10977 22750 11039 22806
rect 10921 22726 11095 22750
rect 10977 22670 11039 22726
rect 10921 22646 11095 22670
rect 10977 22590 11039 22646
rect 10921 22566 11095 22590
rect 10977 22510 11039 22566
rect 10921 22486 11095 22510
rect 10977 22430 11039 22486
rect 10921 22406 11095 22430
rect 10977 22350 11039 22406
rect 10921 22326 11095 22350
rect 10977 22270 11039 22326
rect 10921 22245 11095 22270
rect 10977 22189 11039 22245
rect 10921 22164 11095 22189
rect 10977 22108 11039 22164
rect 10921 22083 11095 22108
rect 10977 22027 11039 22083
rect 10921 22002 11095 22027
rect 10977 21946 11039 22002
rect 10921 21921 11095 21946
rect 10977 21865 11039 21921
rect 10921 21840 11095 21865
rect 10977 21784 11039 21840
rect 10921 21759 11095 21784
rect 10977 21703 11039 21759
rect 10921 21678 11095 21703
rect 10977 21622 11039 21678
rect 10921 21597 11095 21622
rect 10977 21541 11039 21597
rect 10921 21516 11095 21541
rect 10977 21460 11039 21516
rect 10921 21435 11095 21460
rect 10977 21379 11039 21435
rect 10921 21354 11095 21379
rect 10977 21298 11039 21354
rect 10921 21273 11095 21298
rect 10977 21217 11039 21273
rect 10921 21192 11095 21217
rect 10977 21136 11039 21192
rect 10921 21127 11095 21136
rect 11417 23686 11591 23695
rect 11905 23690 12095 23695
rect 11473 23630 11535 23686
rect 11417 23606 11591 23630
rect 11473 23550 11535 23606
rect 11417 23526 11591 23550
rect 11473 23470 11535 23526
rect 11417 23446 11591 23470
rect 11473 23390 11535 23446
rect 11417 23366 11591 23390
rect 11473 23310 11535 23366
rect 11417 23286 11591 23310
rect 11473 23230 11535 23286
rect 11417 23206 11591 23230
rect 11473 23150 11535 23206
rect 11417 23126 11591 23150
rect 11473 23070 11535 23126
rect 11417 23046 11591 23070
rect 11473 22990 11535 23046
rect 11417 22966 11591 22990
rect 11473 22910 11535 22966
rect 11417 22886 11591 22910
rect 11473 22830 11535 22886
rect 11417 22806 11591 22830
rect 11473 22750 11535 22806
rect 11417 22726 11591 22750
rect 11473 22670 11535 22726
rect 11417 22646 11591 22670
rect 11473 22590 11535 22646
rect 11417 22566 11591 22590
rect 11473 22510 11535 22566
rect 11417 22486 11591 22510
rect 11473 22430 11535 22486
rect 11417 22406 11591 22430
rect 11473 22350 11535 22406
rect 11417 22326 11591 22350
rect 11473 22270 11535 22326
rect 11417 22245 11591 22270
rect 11473 22189 11535 22245
rect 11417 22164 11591 22189
rect 11473 22108 11535 22164
rect 11417 22083 11591 22108
rect 11473 22027 11535 22083
rect 11417 22002 11591 22027
rect 11473 21946 11535 22002
rect 11417 21921 11591 21946
rect 11473 21865 11535 21921
rect 11417 21840 11591 21865
rect 11473 21784 11535 21840
rect 11417 21759 11591 21784
rect 11473 21703 11535 21759
rect 11417 21678 11591 21703
rect 11473 21622 11535 21678
rect 11417 21597 11591 21622
rect 11473 21541 11535 21597
rect 11417 21516 11591 21541
rect 11473 21460 11535 21516
rect 11417 21435 11591 21460
rect 11473 21379 11535 21435
rect 11417 21354 11591 21379
rect 11473 21298 11535 21354
rect 11417 21273 11591 21298
rect 11473 21217 11535 21273
rect 11417 21192 11591 21217
rect 11473 21136 11535 21192
rect 11417 21127 11591 21136
rect 11913 23686 12087 23690
rect 11969 23630 12031 23686
rect 11913 23606 12087 23630
rect 11969 23550 12031 23606
rect 11913 23526 12087 23550
rect 11969 23470 12031 23526
rect 11913 23446 12087 23470
rect 11969 23390 12031 23446
rect 11913 23366 12087 23390
rect 11969 23310 12031 23366
rect 11913 23286 12087 23310
rect 11969 23230 12031 23286
rect 11913 23206 12087 23230
rect 11969 23150 12031 23206
rect 11913 23126 12087 23150
rect 11969 23070 12031 23126
rect 11913 23046 12087 23070
rect 11969 22990 12031 23046
rect 11913 22966 12087 22990
rect 11969 22910 12031 22966
rect 11913 22886 12087 22910
rect 11969 22830 12031 22886
rect 11913 22806 12087 22830
rect 11969 22750 12031 22806
rect 11913 22726 12087 22750
rect 11969 22670 12031 22726
rect 11913 22646 12087 22670
rect 11969 22590 12031 22646
rect 11913 22566 12087 22590
rect 11969 22510 12031 22566
rect 11913 22486 12087 22510
rect 11969 22430 12031 22486
rect 11913 22406 12087 22430
rect 11969 22350 12031 22406
rect 11913 22326 12087 22350
rect 11969 22270 12031 22326
rect 11913 22245 12087 22270
rect 11969 22189 12031 22245
rect 11913 22164 12087 22189
rect 11969 22108 12031 22164
rect 11913 22083 12087 22108
rect 11969 22027 12031 22083
rect 11913 22002 12087 22027
rect 11969 21946 12031 22002
rect 11913 21921 12087 21946
rect 11969 21865 12031 21921
rect 11913 21840 12087 21865
rect 11969 21784 12031 21840
rect 11913 21759 12087 21784
rect 11969 21703 12031 21759
rect 11913 21678 12087 21703
rect 11969 21622 12031 21678
rect 11913 21597 12087 21622
rect 11969 21541 12031 21597
rect 11913 21516 12087 21541
rect 11969 21460 12031 21516
rect 11913 21435 12087 21460
rect 11969 21379 12031 21435
rect 11913 21354 12087 21379
rect 11969 21298 12031 21354
rect 11913 21273 12087 21298
rect 11969 21217 12031 21273
rect 11913 21192 12087 21217
rect 11969 21136 12031 21192
rect 11913 21127 12087 21136
rect 12409 23686 12583 23695
rect 12897 23690 13087 23695
rect 12465 23630 12527 23686
rect 12409 23606 12583 23630
rect 12465 23550 12527 23606
rect 12409 23526 12583 23550
rect 12465 23470 12527 23526
rect 12409 23446 12583 23470
rect 12465 23390 12527 23446
rect 12409 23366 12583 23390
rect 12465 23310 12527 23366
rect 12409 23286 12583 23310
rect 12465 23230 12527 23286
rect 12409 23206 12583 23230
rect 12465 23150 12527 23206
rect 12409 23126 12583 23150
rect 12465 23070 12527 23126
rect 12409 23046 12583 23070
rect 12465 22990 12527 23046
rect 12409 22966 12583 22990
rect 12465 22910 12527 22966
rect 12409 22886 12583 22910
rect 12465 22830 12527 22886
rect 12409 22806 12583 22830
rect 12465 22750 12527 22806
rect 12409 22726 12583 22750
rect 12465 22670 12527 22726
rect 12409 22646 12583 22670
rect 12465 22590 12527 22646
rect 12409 22566 12583 22590
rect 12465 22510 12527 22566
rect 12409 22486 12583 22510
rect 12465 22430 12527 22486
rect 12409 22406 12583 22430
rect 12465 22350 12527 22406
rect 12409 22326 12583 22350
rect 12465 22270 12527 22326
rect 12409 22245 12583 22270
rect 12465 22189 12527 22245
rect 12409 22164 12583 22189
rect 12465 22108 12527 22164
rect 12409 22083 12583 22108
rect 12465 22027 12527 22083
rect 12409 22002 12583 22027
rect 12465 21946 12527 22002
rect 12409 21921 12583 21946
rect 12465 21865 12527 21921
rect 12409 21840 12583 21865
rect 12465 21784 12527 21840
rect 12409 21759 12583 21784
rect 12465 21703 12527 21759
rect 12409 21678 12583 21703
rect 12465 21622 12527 21678
rect 12409 21597 12583 21622
rect 12465 21541 12527 21597
rect 12409 21516 12583 21541
rect 12465 21460 12527 21516
rect 12409 21435 12583 21460
rect 12465 21379 12527 21435
rect 12409 21354 12583 21379
rect 12465 21298 12527 21354
rect 12409 21273 12583 21298
rect 12465 21217 12527 21273
rect 12409 21192 12583 21217
rect 12465 21136 12527 21192
rect 12409 21127 12583 21136
rect 12905 23686 13079 23690
rect 12961 23630 13023 23686
rect 12905 23606 13079 23630
rect 12961 23550 13023 23606
rect 12905 23526 13079 23550
rect 12961 23470 13023 23526
rect 12905 23446 13079 23470
rect 12961 23390 13023 23446
rect 12905 23366 13079 23390
rect 12961 23310 13023 23366
rect 12905 23286 13079 23310
rect 12961 23230 13023 23286
rect 12905 23206 13079 23230
rect 12961 23150 13023 23206
rect 12905 23126 13079 23150
rect 12961 23070 13023 23126
rect 12905 23046 13079 23070
rect 12961 22990 13023 23046
rect 12905 22966 13079 22990
rect 12961 22910 13023 22966
rect 12905 22886 13079 22910
rect 12961 22830 13023 22886
rect 12905 22806 13079 22830
rect 12961 22750 13023 22806
rect 12905 22726 13079 22750
rect 12961 22670 13023 22726
rect 12905 22646 13079 22670
rect 12961 22590 13023 22646
rect 12905 22566 13079 22590
rect 12961 22510 13023 22566
rect 12905 22486 13079 22510
rect 12961 22430 13023 22486
rect 12905 22406 13079 22430
rect 12961 22350 13023 22406
rect 12905 22326 13079 22350
rect 12961 22270 13023 22326
rect 12905 22245 13079 22270
rect 12961 22189 13023 22245
rect 12905 22164 13079 22189
rect 12961 22108 13023 22164
rect 12905 22083 13079 22108
rect 12961 22027 13023 22083
rect 12905 22002 13079 22027
rect 12961 21946 13023 22002
rect 12905 21921 13079 21946
rect 12961 21865 13023 21921
rect 12905 21840 13079 21865
rect 12961 21784 13023 21840
rect 12905 21759 13079 21784
rect 12961 21703 13023 21759
rect 12905 21678 13079 21703
rect 12961 21622 13023 21678
rect 12905 21597 13079 21622
rect 12961 21541 13023 21597
rect 12905 21516 13079 21541
rect 12961 21460 13023 21516
rect 12905 21435 13079 21460
rect 12961 21379 13023 21435
rect 12905 21354 13079 21379
rect 12961 21298 13023 21354
rect 12905 21273 13079 21298
rect 12961 21217 13023 21273
rect 12905 21192 13079 21217
rect 12961 21136 13023 21192
rect 12905 21127 13079 21136
rect 13401 23686 13575 23695
rect 13457 23630 13519 23686
rect 13401 23606 13575 23630
rect 13457 23550 13519 23606
rect 13401 23526 13575 23550
rect 13457 23470 13519 23526
rect 13401 23446 13575 23470
rect 13457 23390 13519 23446
rect 13401 23366 13575 23390
rect 13457 23310 13519 23366
rect 13401 23286 13575 23310
rect 13457 23230 13519 23286
rect 13401 23206 13575 23230
rect 13457 23150 13519 23206
rect 13401 23126 13575 23150
rect 13457 23070 13519 23126
rect 13401 23046 13575 23070
rect 13457 22990 13519 23046
rect 13401 22966 13575 22990
rect 13457 22910 13519 22966
rect 13401 22886 13575 22910
rect 13457 22830 13519 22886
rect 13401 22806 13575 22830
rect 13457 22750 13519 22806
rect 13401 22726 13575 22750
rect 13457 22670 13519 22726
rect 13401 22646 13575 22670
rect 13457 22590 13519 22646
rect 13401 22566 13575 22590
rect 13457 22510 13519 22566
rect 13401 22486 13575 22510
rect 13457 22430 13519 22486
rect 13401 22406 13575 22430
rect 13457 22350 13519 22406
rect 13401 22326 13575 22350
rect 13457 22270 13519 22326
rect 13401 22245 13575 22270
rect 13457 22189 13519 22245
rect 13401 22164 13575 22189
rect 13457 22108 13519 22164
rect 13401 22083 13575 22108
rect 13457 22027 13519 22083
rect 13401 22002 13575 22027
rect 13457 21946 13519 22002
rect 13401 21921 13575 21946
rect 13457 21865 13519 21921
rect 13401 21840 13575 21865
rect 13457 21784 13519 21840
rect 13401 21759 13575 21784
rect 13457 21703 13519 21759
rect 13401 21678 13575 21703
rect 13457 21622 13519 21678
rect 13401 21597 13575 21622
rect 13457 21541 13519 21597
rect 13401 21516 13575 21541
rect 13457 21460 13519 21516
rect 13401 21435 13575 21460
rect 13457 21379 13519 21435
rect 13401 21354 13575 21379
rect 13457 21298 13519 21354
rect 13401 21273 13575 21298
rect 13457 21217 13519 21273
rect 13401 21192 13575 21217
rect 13457 21136 13519 21192
rect 13401 21127 13575 21136
rect 13838 23686 14012 23695
rect 13894 23630 13956 23686
rect 13838 23606 14012 23630
rect 13894 23550 13956 23606
rect 13838 23526 14012 23550
rect 13894 23470 13956 23526
rect 13838 23446 14012 23470
rect 13894 23390 13956 23446
rect 13838 23366 14012 23390
rect 13894 23310 13956 23366
rect 13838 23286 14012 23310
rect 13894 23230 13956 23286
rect 13838 23206 14012 23230
rect 13894 23150 13956 23206
rect 13838 23126 14012 23150
rect 13894 23070 13956 23126
rect 13838 23046 14012 23070
rect 13894 22990 13956 23046
rect 13838 22966 14012 22990
rect 13894 22910 13956 22966
rect 13838 22886 14012 22910
rect 13894 22830 13956 22886
rect 13838 22806 14012 22830
rect 13894 22750 13956 22806
rect 13838 22726 14012 22750
rect 13894 22670 13956 22726
rect 13838 22646 14012 22670
rect 13894 22590 13956 22646
rect 13838 22566 14012 22590
rect 13894 22510 13956 22566
rect 13838 22486 14012 22510
rect 13894 22430 13956 22486
rect 13838 22406 14012 22430
rect 13894 22350 13956 22406
rect 13838 22326 14012 22350
rect 13894 22270 13956 22326
rect 13838 22245 14012 22270
rect 13894 22189 13956 22245
rect 13838 22164 14012 22189
rect 13894 22108 13956 22164
rect 13838 22083 14012 22108
rect 13894 22027 13956 22083
rect 13838 22002 14012 22027
rect 13894 21946 13956 22002
rect 13838 21921 14012 21946
rect 13894 21865 13956 21921
rect 13838 21840 14012 21865
rect 13894 21784 13956 21840
rect 13838 21759 14012 21784
rect 13894 21703 13956 21759
rect 13838 21678 14012 21703
rect 13894 21622 13956 21678
rect 13838 21597 14012 21622
rect 13894 21541 13956 21597
rect 13838 21516 14012 21541
rect 13894 21460 13956 21516
rect 13838 21435 14012 21460
rect 13894 21379 13956 21435
rect 13838 21354 14012 21379
rect 13894 21298 13956 21354
rect 13838 21273 14012 21298
rect 13894 21217 13956 21273
rect 13838 21192 14012 21217
rect 13894 21136 13956 21192
rect 13838 21127 14012 21136
rect 14281 23685 14283 23741
rect 14339 23685 14381 23741
rect 14437 23685 14479 23741
rect 14535 23685 14577 23741
rect 14633 23685 14639 23741
rect 14281 23660 14639 23685
rect 14281 23604 14283 23660
rect 14339 23604 14381 23660
rect 14437 23604 14479 23660
rect 14535 23604 14577 23660
rect 14633 23604 14639 23660
rect 14281 23579 14639 23604
rect 14281 23523 14283 23579
rect 14339 23523 14381 23579
rect 14437 23523 14479 23579
rect 14535 23523 14577 23579
rect 14633 23523 14639 23579
rect 14281 23498 14639 23523
rect 14281 23442 14283 23498
rect 14339 23442 14381 23498
rect 14437 23442 14479 23498
rect 14535 23442 14577 23498
rect 14633 23442 14639 23498
rect 14281 23417 14639 23442
rect 14281 23361 14283 23417
rect 14339 23361 14381 23417
rect 14437 23361 14479 23417
rect 14535 23361 14577 23417
rect 14633 23361 14639 23417
rect 14281 23336 14639 23361
rect 14281 23280 14283 23336
rect 14339 23280 14381 23336
rect 14437 23280 14479 23336
rect 14535 23280 14577 23336
rect 14633 23280 14639 23336
rect 14281 23255 14639 23280
rect 14281 23199 14283 23255
rect 14339 23199 14381 23255
rect 14437 23199 14479 23255
rect 14535 23199 14577 23255
rect 14633 23199 14639 23255
rect 14281 23174 14639 23199
rect 14281 23118 14283 23174
rect 14339 23118 14381 23174
rect 14437 23118 14479 23174
rect 14535 23118 14577 23174
rect 14633 23118 14639 23174
rect 14281 23093 14639 23118
rect 14281 23037 14283 23093
rect 14339 23037 14381 23093
rect 14437 23037 14479 23093
rect 14535 23037 14577 23093
rect 14633 23037 14639 23093
rect 14281 23012 14639 23037
rect 14281 22956 14283 23012
rect 14339 22956 14381 23012
rect 14437 22956 14479 23012
rect 14535 22956 14577 23012
rect 14633 22956 14639 23012
rect 14281 22931 14639 22956
rect 14281 22875 14283 22931
rect 14339 22875 14381 22931
rect 14437 22875 14479 22931
rect 14535 22875 14577 22931
rect 14633 22875 14639 22931
rect 14281 22850 14639 22875
rect 14281 22794 14283 22850
rect 14339 22794 14381 22850
rect 14437 22794 14479 22850
rect 14535 22794 14577 22850
rect 14633 22794 14639 22850
rect 14281 22769 14639 22794
rect 14281 22713 14283 22769
rect 14339 22713 14381 22769
rect 14437 22713 14479 22769
rect 14535 22713 14577 22769
rect 14633 22713 14639 22769
rect 14281 22688 14639 22713
rect 14281 22632 14283 22688
rect 14339 22632 14381 22688
rect 14437 22632 14479 22688
rect 14535 22632 14577 22688
rect 14633 22632 14639 22688
rect 14281 22607 14639 22632
rect 14281 22551 14283 22607
rect 14339 22551 14381 22607
rect 14437 22551 14479 22607
rect 14535 22551 14577 22607
rect 14633 22551 14639 22607
rect 14281 22526 14639 22551
rect 14281 22470 14283 22526
rect 14339 22470 14381 22526
rect 14437 22470 14479 22526
rect 14535 22470 14577 22526
rect 14633 22470 14639 22526
rect 14281 22445 14639 22470
rect 14281 22389 14283 22445
rect 14339 22389 14381 22445
rect 14437 22389 14479 22445
rect 14535 22389 14577 22445
rect 14633 22389 14639 22445
rect 14783 22428 14823 35604
rect 14863 22428 14903 35684
rect 14943 22428 14983 35764
rect 14281 22364 14639 22389
rect 14281 22308 14283 22364
rect 14339 22308 14381 22364
rect 14437 22308 14479 22364
rect 14535 22308 14577 22364
rect 14633 22308 14639 22364
rect 14281 22283 14639 22308
rect 14281 22227 14283 22283
rect 14339 22227 14381 22283
rect 14437 22227 14479 22283
rect 14535 22227 14577 22283
rect 14633 22227 14639 22283
rect 14281 22202 14639 22227
rect 14281 22146 14283 22202
rect 14339 22146 14381 22202
rect 14437 22146 14479 22202
rect 14535 22146 14577 22202
rect 14633 22146 14639 22202
rect 14281 22121 14639 22146
rect 14281 22065 14283 22121
rect 14339 22065 14381 22121
rect 14437 22065 14479 22121
rect 14535 22065 14577 22121
rect 14633 22065 14639 22121
rect 14281 22040 14639 22065
rect 14281 21984 14283 22040
rect 14339 21984 14381 22040
rect 14437 21984 14479 22040
rect 14535 21984 14577 22040
rect 14633 21984 14639 22040
rect 14281 21959 14639 21984
rect 14281 21903 14283 21959
rect 14339 21903 14381 21959
rect 14437 21903 14479 21959
rect 14535 21903 14577 21959
rect 14633 21903 14639 21959
rect 14281 21878 14639 21903
rect 14281 21822 14283 21878
rect 14339 21822 14381 21878
rect 14437 21822 14479 21878
rect 14535 21822 14577 21878
rect 14633 21822 14639 21878
rect 14281 21797 14639 21822
rect 14281 21741 14283 21797
rect 14339 21741 14381 21797
rect 14437 21741 14479 21797
rect 14535 21741 14577 21797
rect 14633 21741 14639 21797
rect 14281 21716 14639 21741
rect 14281 21660 14283 21716
rect 14339 21660 14381 21716
rect 14437 21660 14479 21716
rect 14535 21660 14577 21716
rect 14633 21660 14639 21716
rect 14281 21635 14639 21660
rect 14281 21579 14283 21635
rect 14339 21579 14381 21635
rect 14437 21579 14479 21635
rect 14535 21579 14577 21635
rect 14633 21579 14639 21635
rect 14281 21554 14639 21579
rect 14281 21498 14283 21554
rect 14339 21498 14381 21554
rect 14437 21498 14479 21554
rect 14535 21498 14577 21554
rect 14633 21498 14639 21554
rect 14281 21473 14639 21498
rect 14281 21417 14283 21473
rect 14339 21417 14381 21473
rect 14437 21417 14479 21473
rect 14535 21417 14577 21473
rect 14633 21417 14639 21473
rect 14281 21392 14639 21417
rect 14281 21336 14283 21392
rect 14339 21336 14381 21392
rect 14437 21336 14479 21392
rect 14535 21336 14577 21392
rect 14633 21336 14639 21392
rect 14281 21311 14639 21336
rect 14281 21255 14283 21311
rect 14339 21255 14381 21311
rect 14437 21255 14479 21311
rect 14535 21255 14577 21311
rect 14633 21255 14639 21311
rect 14281 21230 14639 21255
rect 14281 21174 14283 21230
rect 14339 21174 14381 21230
rect 14437 21174 14479 21230
rect 14535 21174 14577 21230
rect 14633 21174 14639 21230
rect 14281 21149 14639 21174
rect 164 21065 242 21121
rect 298 21065 334 21121
rect 390 21065 426 21121
rect 482 21065 518 21121
rect 574 21065 610 21121
rect 666 21065 702 21121
rect 758 21065 778 21121
rect 164 21040 778 21065
rect 164 20984 242 21040
rect 298 20984 334 21040
rect 390 20984 426 21040
rect 482 20984 518 21040
rect 574 20984 610 21040
rect 666 20984 702 21040
rect 758 20984 778 21040
rect 164 20959 778 20984
rect 164 20903 242 20959
rect 298 20903 334 20959
rect 390 20903 426 20959
rect 482 20903 518 20959
rect 574 20903 610 20959
rect 666 20903 702 20959
rect 758 20903 778 20959
rect 164 20878 778 20903
rect 164 20822 242 20878
rect 298 20822 334 20878
rect 390 20822 426 20878
rect 482 20822 518 20878
rect 574 20822 610 20878
rect 666 20822 702 20878
rect 758 20822 778 20878
rect 164 20797 778 20822
rect 164 20741 242 20797
rect 298 20741 334 20797
rect 390 20741 426 20797
rect 482 20741 518 20797
rect 574 20741 610 20797
rect 666 20741 702 20797
rect 758 20741 778 20797
rect 164 20716 778 20741
rect 164 20660 242 20716
rect 298 20660 334 20716
rect 390 20660 426 20716
rect 482 20660 518 20716
rect 574 20660 610 20716
rect 666 20660 702 20716
rect 758 20660 778 20716
rect 164 20635 778 20660
rect 164 20579 242 20635
rect 298 20579 334 20635
rect 390 20579 426 20635
rect 482 20579 518 20635
rect 574 20579 610 20635
rect 666 20579 702 20635
rect 758 20579 778 20635
rect 164 20554 778 20579
rect 164 20498 242 20554
rect 298 20498 334 20554
rect 390 20498 426 20554
rect 482 20498 518 20554
rect 574 20498 610 20554
rect 666 20498 702 20554
rect 758 20498 778 20554
rect 14281 21093 14283 21149
rect 14339 21093 14381 21149
rect 14437 21093 14479 21149
rect 14535 21093 14577 21149
rect 14633 21093 14639 21149
rect 14281 21068 14639 21093
rect 14281 21012 14283 21068
rect 14339 21012 14381 21068
rect 14437 21012 14479 21068
rect 14535 21012 14577 21068
rect 14633 21012 14639 21068
rect 14281 20987 14639 21012
rect 14281 20931 14283 20987
rect 14339 20931 14381 20987
rect 14437 20931 14479 20987
rect 14535 20931 14577 20987
rect 14633 20931 14639 20987
rect 14281 20906 14639 20931
rect 14281 20850 14283 20906
rect 14339 20850 14381 20906
rect 14437 20850 14479 20906
rect 14535 20850 14577 20906
rect 14633 20850 14639 20906
rect 14281 20825 14639 20850
rect 14281 20769 14283 20825
rect 14339 20769 14381 20825
rect 14437 20769 14479 20825
rect 14535 20769 14577 20825
rect 14633 20769 14639 20825
rect 14281 20744 14639 20769
rect 14281 20688 14283 20744
rect 14339 20688 14381 20744
rect 14437 20688 14479 20744
rect 14535 20688 14577 20744
rect 14633 20688 14639 20744
rect 14281 20663 14639 20688
rect 14281 20607 14283 20663
rect 14339 20607 14381 20663
rect 14437 20607 14479 20663
rect 14535 20607 14577 20663
rect 14633 20607 14639 20663
rect 14281 20582 14639 20607
rect 14281 20526 14283 20582
rect 14339 20526 14381 20582
rect 14437 20526 14479 20582
rect 14535 20526 14577 20582
rect 14633 20526 14639 20582
rect 14281 20517 14639 20526
rect 14754 21413 14940 21419
rect 14754 21361 14755 21413
rect 14807 21361 14821 21413
rect 14873 21361 14887 21413
rect 14939 21361 14940 21413
rect 14754 21348 14940 21361
rect 14754 21296 14755 21348
rect 14807 21296 14821 21348
rect 14873 21296 14887 21348
rect 14939 21296 14940 21348
rect 14754 21282 14940 21296
rect 14754 21230 14755 21282
rect 14807 21230 14821 21282
rect 14873 21230 14887 21282
rect 14939 21230 14940 21282
rect 14754 21216 14940 21230
rect 14754 21164 14755 21216
rect 14807 21164 14821 21216
rect 14873 21164 14887 21216
rect 14939 21164 14940 21216
rect 14754 21150 14940 21164
rect 14754 21098 14755 21150
rect 14807 21098 14821 21150
rect 14873 21098 14887 21150
rect 14939 21098 14940 21150
rect 14754 21084 14940 21098
rect 14754 21032 14755 21084
rect 14807 21032 14821 21084
rect 14873 21032 14887 21084
rect 14939 21032 14940 21084
rect 14754 21018 14940 21032
rect 14754 20966 14755 21018
rect 14807 20966 14821 21018
rect 14873 20966 14887 21018
rect 14939 20966 14940 21018
rect 14754 20952 14940 20966
rect 14754 20900 14755 20952
rect 14807 20900 14821 20952
rect 14873 20900 14887 20952
rect 14939 20900 14940 20952
rect 14754 20886 14940 20900
rect 14754 20834 14755 20886
rect 14807 20834 14821 20886
rect 14873 20834 14887 20886
rect 14939 20834 14940 20886
rect 14754 20820 14940 20834
rect 14754 20768 14755 20820
rect 14807 20768 14821 20820
rect 14873 20768 14887 20820
rect 14939 20768 14940 20820
rect 14754 20754 14940 20768
rect 14754 20702 14755 20754
rect 14807 20702 14821 20754
rect 14873 20702 14887 20754
rect 14939 20702 14940 20754
rect 14754 20688 14940 20702
rect 14754 20636 14755 20688
rect 14807 20636 14821 20688
rect 14873 20636 14887 20688
rect 14939 20636 14940 20688
rect 14754 20622 14940 20636
rect 14754 20570 14755 20622
rect 14807 20570 14821 20622
rect 14873 20570 14887 20622
rect 14939 20570 14940 20622
rect 14754 20556 14940 20570
rect 164 20473 778 20498
rect 164 20417 242 20473
rect 298 20417 334 20473
rect 390 20417 426 20473
rect 482 20417 518 20473
rect 574 20417 610 20473
rect 666 20417 702 20473
rect 758 20417 778 20473
rect 164 20387 778 20417
rect 14754 20504 14755 20556
rect 14807 20504 14821 20556
rect 14873 20504 14887 20556
rect 14939 20504 14940 20556
rect 14754 20490 14940 20504
rect 14754 20438 14755 20490
rect 14807 20438 14821 20490
rect 14873 20438 14887 20490
rect 14939 20438 14940 20490
rect 14754 20424 14940 20438
rect 14754 20372 14755 20424
rect 14807 20372 14821 20424
rect 14873 20372 14887 20424
rect 14939 20372 14940 20424
rect 14754 20358 14940 20372
rect 14754 20306 14755 20358
rect 14807 20306 14821 20358
rect 14873 20306 14887 20358
rect 14939 20306 14940 20358
rect 14754 20292 14940 20306
rect 14754 20240 14755 20292
rect 14807 20240 14821 20292
rect 14873 20240 14887 20292
rect 14939 20240 14940 20292
rect 14754 20226 14940 20240
rect 14754 20174 14755 20226
rect 14807 20174 14821 20226
rect 14873 20174 14887 20226
rect 14939 20174 14940 20226
rect 14754 20160 14940 20174
rect 14754 20108 14755 20160
rect 14807 20108 14821 20160
rect 14873 20108 14887 20160
rect 14939 20108 14940 20160
rect 14754 20094 14940 20108
rect 14754 20042 14755 20094
rect 14807 20042 14821 20094
rect 14873 20042 14887 20094
rect 14939 20042 14940 20094
rect 14754 20028 14940 20042
rect 14754 19976 14755 20028
rect 14807 19976 14821 20028
rect 14873 19976 14887 20028
rect 14939 19976 14940 20028
rect 194 19964 1266 19967
rect 194 19912 201 19964
rect 253 19912 269 19964
rect 321 19912 337 19964
rect 389 19912 404 19964
rect 456 19912 471 19964
rect 523 19912 538 19964
rect 590 19912 605 19964
rect 657 19912 672 19964
rect 724 19912 739 19964
rect 791 19912 806 19964
rect 858 19912 873 19964
rect 925 19912 940 19964
rect 992 19912 1007 19964
rect 1059 19912 1074 19964
rect 1126 19912 1141 19964
rect 1193 19912 1208 19964
rect 1260 19912 1266 19964
rect 194 19896 1266 19912
rect 194 19844 201 19896
rect 253 19844 269 19896
rect 321 19844 337 19896
rect 389 19844 404 19896
rect 456 19844 471 19896
rect 523 19844 538 19896
rect 590 19844 605 19896
rect 657 19844 672 19896
rect 724 19844 739 19896
rect 791 19844 806 19896
rect 858 19844 873 19896
rect 925 19844 940 19896
rect 992 19844 1007 19896
rect 1059 19844 1074 19896
rect 1126 19844 1141 19896
rect 1193 19844 1208 19896
rect 1260 19844 1266 19896
rect 194 19828 1266 19844
rect 194 19776 201 19828
rect 253 19776 269 19828
rect 321 19776 337 19828
rect 389 19776 404 19828
rect 456 19776 471 19828
rect 523 19776 538 19828
rect 590 19776 605 19828
rect 657 19776 672 19828
rect 724 19776 739 19828
rect 791 19776 806 19828
rect 858 19776 873 19828
rect 925 19776 940 19828
rect 992 19776 1007 19828
rect 1059 19776 1074 19828
rect 1126 19776 1141 19828
rect 1193 19776 1208 19828
rect 1260 19776 1266 19828
rect 194 19760 1266 19776
rect 194 19708 201 19760
rect 253 19708 269 19760
rect 321 19708 337 19760
rect 389 19708 404 19760
rect 456 19708 471 19760
rect 523 19708 538 19760
rect 590 19708 605 19760
rect 657 19708 672 19760
rect 724 19708 739 19760
rect 791 19708 806 19760
rect 858 19708 873 19760
rect 925 19708 940 19760
rect 992 19708 1007 19760
rect 1059 19708 1074 19760
rect 1126 19708 1141 19760
rect 1193 19708 1208 19760
rect 1260 19708 1266 19760
rect 194 19692 1266 19708
rect 194 19640 201 19692
rect 253 19640 269 19692
rect 321 19640 337 19692
rect 389 19640 404 19692
rect 456 19640 471 19692
rect 523 19640 538 19692
rect 590 19640 605 19692
rect 657 19640 672 19692
rect 724 19640 739 19692
rect 791 19640 806 19692
rect 858 19640 873 19692
rect 925 19640 940 19692
rect 992 19640 1007 19692
rect 1059 19640 1074 19692
rect 1126 19640 1141 19692
rect 1193 19640 1208 19692
rect 1260 19640 1266 19692
rect 194 19624 1266 19640
rect 194 19572 201 19624
rect 253 19572 269 19624
rect 321 19572 337 19624
rect 389 19572 404 19624
rect 456 19572 471 19624
rect 523 19572 538 19624
rect 590 19572 605 19624
rect 657 19572 672 19624
rect 724 19572 739 19624
rect 791 19572 806 19624
rect 858 19572 873 19624
rect 925 19572 940 19624
rect 992 19572 1007 19624
rect 1059 19572 1074 19624
rect 1126 19572 1141 19624
rect 1193 19572 1208 19624
rect 1260 19572 1266 19624
rect 194 18387 1266 19572
rect 194 18335 201 18387
rect 253 18335 269 18387
rect 321 18335 337 18387
rect 389 18335 404 18387
rect 456 18335 471 18387
rect 523 18335 538 18387
rect 590 18335 605 18387
rect 657 18335 672 18387
rect 724 18335 739 18387
rect 791 18335 806 18387
rect 858 18335 873 18387
rect 925 18335 940 18387
rect 992 18335 1007 18387
rect 1059 18335 1074 18387
rect 1126 18335 1141 18387
rect 1193 18335 1208 18387
rect 1260 18335 1266 18387
rect 194 18323 1266 18335
rect 194 18271 201 18323
rect 253 18271 269 18323
rect 321 18271 337 18323
rect 389 18271 404 18323
rect 456 18271 471 18323
rect 523 18271 538 18323
rect 590 18271 605 18323
rect 657 18271 672 18323
rect 724 18271 739 18323
rect 791 18271 806 18323
rect 858 18271 873 18323
rect 925 18271 940 18323
rect 992 18271 1007 18323
rect 1059 18271 1074 18323
rect 1126 18271 1141 18323
rect 1193 18271 1208 18323
rect 1260 18271 1266 18323
rect 194 18259 1266 18271
rect 194 18207 201 18259
rect 253 18207 269 18259
rect 321 18207 337 18259
rect 389 18207 404 18259
rect 456 18207 471 18259
rect 523 18207 538 18259
rect 590 18207 605 18259
rect 657 18207 672 18259
rect 724 18207 739 18259
rect 791 18207 806 18259
rect 858 18207 873 18259
rect 925 18207 940 18259
rect 992 18207 1007 18259
rect 1059 18207 1074 18259
rect 1126 18207 1141 18259
rect 1193 18207 1208 18259
rect 1260 18207 1266 18259
rect 194 18195 1266 18207
rect 194 18143 201 18195
rect 253 18143 269 18195
rect 321 18143 337 18195
rect 389 18143 404 18195
rect 456 18143 471 18195
rect 523 18143 538 18195
rect 590 18143 605 18195
rect 657 18143 672 18195
rect 724 18143 739 18195
rect 791 18143 806 18195
rect 858 18143 873 18195
rect 925 18143 940 18195
rect 992 18143 1007 18195
rect 1059 18143 1074 18195
rect 1126 18143 1141 18195
rect 1193 18143 1208 18195
rect 1260 18143 1266 18195
rect 194 18131 1266 18143
rect 194 18079 201 18131
rect 253 18079 269 18131
rect 321 18079 337 18131
rect 389 18079 404 18131
rect 456 18079 471 18131
rect 523 18079 538 18131
rect 590 18079 605 18131
rect 657 18079 672 18131
rect 724 18079 739 18131
rect 791 18079 806 18131
rect 858 18079 873 18131
rect 925 18079 940 18131
rect 992 18079 1007 18131
rect 1059 18079 1074 18131
rect 1126 18079 1141 18131
rect 1193 18079 1208 18131
rect 1260 18079 1266 18131
rect 194 18067 1266 18079
rect 194 18015 201 18067
rect 253 18015 269 18067
rect 321 18015 337 18067
rect 389 18015 404 18067
rect 456 18015 471 18067
rect 523 18015 538 18067
rect 590 18015 605 18067
rect 657 18015 672 18067
rect 724 18015 739 18067
rect 791 18015 806 18067
rect 858 18015 873 18067
rect 925 18015 940 18067
rect 992 18015 1007 18067
rect 1059 18015 1074 18067
rect 1126 18015 1141 18067
rect 1193 18015 1208 18067
rect 1260 18015 1266 18067
rect 194 18003 1266 18015
rect 194 17951 201 18003
rect 253 17951 269 18003
rect 321 17951 337 18003
rect 389 17951 404 18003
rect 456 17951 471 18003
rect 523 17951 538 18003
rect 590 17951 605 18003
rect 657 17951 672 18003
rect 724 17951 739 18003
rect 791 17951 806 18003
rect 858 17951 873 18003
rect 925 17951 940 18003
rect 992 17951 1007 18003
rect 1059 17951 1074 18003
rect 1126 17951 1141 18003
rect 1193 17951 1208 18003
rect 1260 17951 1266 18003
rect 194 17939 1266 17951
rect 194 17887 201 17939
rect 253 17887 269 17939
rect 321 17887 337 17939
rect 389 17887 404 17939
rect 456 17887 471 17939
rect 523 17887 538 17939
rect 590 17887 605 17939
rect 657 17887 672 17939
rect 724 17887 739 17939
rect 791 17887 806 17939
rect 858 17887 873 17939
rect 925 17887 940 17939
rect 992 17887 1007 17939
rect 1059 17887 1074 17939
rect 1126 17887 1141 17939
rect 1193 17887 1208 17939
rect 1260 17887 1266 17939
rect 194 8841 1266 17887
rect 194 8785 203 8841
rect 259 8785 287 8841
rect 343 8785 371 8841
rect 427 8785 454 8841
rect 510 8785 537 8841
rect 593 8785 620 8841
rect 676 8785 703 8841
rect 759 8785 786 8841
rect 842 8785 869 8841
rect 925 8785 952 8841
rect 1008 8785 1035 8841
rect 1091 8785 1118 8841
rect 1174 8785 1201 8841
rect 1257 8785 1266 8841
rect 194 8755 1266 8785
rect 194 8699 203 8755
rect 259 8699 287 8755
rect 343 8699 371 8755
rect 427 8699 454 8755
rect 510 8699 537 8755
rect 593 8699 620 8755
rect 676 8699 703 8755
rect 759 8699 786 8755
rect 842 8699 869 8755
rect 925 8699 952 8755
rect 1008 8699 1035 8755
rect 1091 8699 1118 8755
rect 1174 8699 1201 8755
rect 1257 8699 1266 8755
rect 194 8669 1266 8699
rect 194 8613 203 8669
rect 259 8613 287 8669
rect 343 8613 371 8669
rect 427 8613 454 8669
rect 510 8613 537 8669
rect 593 8613 620 8669
rect 676 8613 703 8669
rect 759 8613 786 8669
rect 842 8613 869 8669
rect 925 8613 952 8669
rect 1008 8613 1035 8669
rect 1091 8613 1118 8669
rect 1174 8613 1201 8669
rect 1257 8613 1266 8669
rect 194 8583 1266 8613
rect 194 8527 203 8583
rect 259 8527 287 8583
rect 343 8527 371 8583
rect 427 8527 454 8583
rect 510 8527 537 8583
rect 593 8527 620 8583
rect 676 8527 703 8583
rect 759 8527 786 8583
rect 842 8527 869 8583
rect 925 8527 952 8583
rect 1008 8527 1035 8583
rect 1091 8527 1118 8583
rect 1174 8527 1201 8583
rect 1257 8527 1266 8583
rect 194 8497 1266 8527
rect 194 8441 203 8497
rect 259 8441 287 8497
rect 343 8441 371 8497
rect 427 8441 454 8497
rect 510 8441 537 8497
rect 593 8441 620 8497
rect 676 8441 703 8497
rect 759 8441 786 8497
rect 842 8441 869 8497
rect 925 8441 952 8497
rect 1008 8441 1035 8497
rect 1091 8441 1118 8497
rect 1174 8441 1201 8497
rect 1257 8441 1266 8497
rect 194 8411 1266 8441
rect 194 8355 203 8411
rect 259 8355 287 8411
rect 343 8355 371 8411
rect 427 8355 454 8411
rect 510 8355 537 8411
rect 593 8355 620 8411
rect 676 8355 703 8411
rect 759 8355 786 8411
rect 842 8355 869 8411
rect 925 8355 952 8411
rect 1008 8355 1035 8411
rect 1091 8355 1118 8411
rect 1174 8355 1201 8411
rect 1257 8355 1266 8411
rect 194 8325 1266 8355
rect 194 8269 203 8325
rect 259 8269 287 8325
rect 343 8269 371 8325
rect 427 8269 454 8325
rect 510 8269 537 8325
rect 593 8269 620 8325
rect 676 8269 703 8325
rect 759 8269 786 8325
rect 842 8269 869 8325
rect 925 8269 952 8325
rect 1008 8269 1035 8325
rect 1091 8269 1118 8325
rect 1174 8269 1201 8325
rect 1257 8269 1266 8325
rect 194 8239 1266 8269
rect 194 8183 203 8239
rect 259 8183 287 8239
rect 343 8183 371 8239
rect 427 8183 454 8239
rect 510 8183 537 8239
rect 593 8183 620 8239
rect 676 8183 703 8239
rect 759 8183 786 8239
rect 842 8183 869 8239
rect 925 8183 952 8239
rect 1008 8183 1035 8239
rect 1091 8183 1118 8239
rect 1174 8183 1201 8239
rect 1257 8183 1266 8239
rect 194 8153 1266 8183
rect 194 8097 203 8153
rect 259 8097 287 8153
rect 343 8097 371 8153
rect 427 8097 454 8153
rect 510 8097 537 8153
rect 593 8097 620 8153
rect 676 8097 703 8153
rect 759 8097 786 8153
rect 842 8097 869 8153
rect 925 8097 952 8153
rect 1008 8097 1035 8153
rect 1091 8097 1118 8153
rect 1174 8097 1201 8153
rect 1257 8097 1266 8153
rect 194 8067 1266 8097
rect 194 8011 203 8067
rect 259 8011 287 8067
rect 343 8011 371 8067
rect 427 8011 454 8067
rect 510 8011 537 8067
rect 593 8011 620 8067
rect 676 8011 703 8067
rect 759 8011 786 8067
rect 842 8011 869 8067
rect 925 8011 952 8067
rect 1008 8011 1035 8067
rect 1091 8011 1118 8067
rect 1174 8011 1201 8067
rect 1257 8011 1266 8067
rect 194 7981 1266 8011
rect 194 7925 203 7981
rect 259 7925 287 7981
rect 343 7925 371 7981
rect 427 7925 454 7981
rect 510 7925 537 7981
rect 593 7925 620 7981
rect 676 7925 703 7981
rect 759 7925 786 7981
rect 842 7925 869 7981
rect 925 7925 952 7981
rect 1008 7925 1035 7981
rect 1091 7925 1118 7981
rect 1174 7925 1201 7981
rect 1257 7925 1266 7981
rect 194 7916 1266 7925
rect 8194 19964 9265 19967
rect 8194 19912 8200 19964
rect 8252 19912 8268 19964
rect 8320 19912 8336 19964
rect 8388 19912 8403 19964
rect 8455 19912 8470 19964
rect 8522 19912 8537 19964
rect 8589 19912 8604 19964
rect 8656 19912 8671 19964
rect 8723 19912 8738 19964
rect 8790 19912 8805 19964
rect 8857 19912 8872 19964
rect 8924 19912 8939 19964
rect 8991 19912 9006 19964
rect 9058 19912 9073 19964
rect 9125 19912 9140 19964
rect 9192 19912 9207 19964
rect 9259 19912 9265 19964
rect 8194 19896 9265 19912
rect 8194 19844 8200 19896
rect 8252 19844 8268 19896
rect 8320 19844 8336 19896
rect 8388 19844 8403 19896
rect 8455 19844 8470 19896
rect 8522 19844 8537 19896
rect 8589 19844 8604 19896
rect 8656 19844 8671 19896
rect 8723 19844 8738 19896
rect 8790 19844 8805 19896
rect 8857 19844 8872 19896
rect 8924 19844 8939 19896
rect 8991 19844 9006 19896
rect 9058 19844 9073 19896
rect 9125 19844 9140 19896
rect 9192 19844 9207 19896
rect 9259 19844 9265 19896
rect 8194 19828 9265 19844
rect 8194 19776 8200 19828
rect 8252 19776 8268 19828
rect 8320 19776 8336 19828
rect 8388 19776 8403 19828
rect 8455 19776 8470 19828
rect 8522 19776 8537 19828
rect 8589 19776 8604 19828
rect 8656 19776 8671 19828
rect 8723 19776 8738 19828
rect 8790 19776 8805 19828
rect 8857 19776 8872 19828
rect 8924 19776 8939 19828
rect 8991 19776 9006 19828
rect 9058 19776 9073 19828
rect 9125 19776 9140 19828
rect 9192 19776 9207 19828
rect 9259 19776 9265 19828
rect 8194 19760 9265 19776
rect 8194 19708 8200 19760
rect 8252 19708 8268 19760
rect 8320 19708 8336 19760
rect 8388 19708 8403 19760
rect 8455 19708 8470 19760
rect 8522 19708 8537 19760
rect 8589 19708 8604 19760
rect 8656 19708 8671 19760
rect 8723 19708 8738 19760
rect 8790 19708 8805 19760
rect 8857 19708 8872 19760
rect 8924 19708 8939 19760
rect 8991 19708 9006 19760
rect 9058 19708 9073 19760
rect 9125 19708 9140 19760
rect 9192 19708 9207 19760
rect 9259 19708 9265 19760
rect 8194 19692 9265 19708
rect 8194 19640 8200 19692
rect 8252 19640 8268 19692
rect 8320 19640 8336 19692
rect 8388 19640 8403 19692
rect 8455 19640 8470 19692
rect 8522 19640 8537 19692
rect 8589 19640 8604 19692
rect 8656 19640 8671 19692
rect 8723 19640 8738 19692
rect 8790 19640 8805 19692
rect 8857 19640 8872 19692
rect 8924 19640 8939 19692
rect 8991 19640 9006 19692
rect 9058 19640 9073 19692
rect 9125 19640 9140 19692
rect 9192 19640 9207 19692
rect 9259 19640 9265 19692
rect 8194 19624 9265 19640
rect 8194 19572 8200 19624
rect 8252 19572 8268 19624
rect 8320 19572 8336 19624
rect 8388 19572 8403 19624
rect 8455 19572 8470 19624
rect 8522 19572 8537 19624
rect 8589 19572 8604 19624
rect 8656 19572 8671 19624
rect 8723 19572 8738 19624
rect 8790 19572 8805 19624
rect 8857 19572 8872 19624
rect 8924 19572 8939 19624
rect 8991 19572 9006 19624
rect 9058 19572 9073 19624
rect 9125 19572 9140 19624
rect 9192 19572 9207 19624
rect 9259 19572 9265 19624
rect 14754 19962 14940 19976
rect 14754 19910 14755 19962
rect 14807 19910 14821 19962
rect 14873 19910 14887 19962
rect 14939 19910 14940 19962
rect 14754 19896 14940 19910
rect 14754 19844 14755 19896
rect 14807 19844 14821 19896
rect 14873 19844 14887 19896
rect 14939 19844 14940 19896
rect 14754 19830 14940 19844
rect 14754 19778 14755 19830
rect 14807 19778 14821 19830
rect 14873 19778 14887 19830
rect 14939 19778 14940 19830
rect 14754 19764 14940 19778
rect 14754 19712 14755 19764
rect 14807 19712 14821 19764
rect 14873 19712 14887 19764
rect 14939 19712 14940 19764
rect 14754 19698 14940 19712
rect 14754 19646 14755 19698
rect 14807 19646 14821 19698
rect 14873 19646 14887 19698
rect 14939 19646 14940 19698
rect 14754 19632 14940 19646
rect 14754 19580 14755 19632
rect 14807 19580 14821 19632
rect 14873 19580 14887 19632
rect 14939 19580 14940 19632
rect 14754 19574 14940 19580
rect 8194 8841 9265 19572
rect 12610 18817 12740 18850
rect 12610 18765 12616 18817
rect 12668 18765 12682 18817
rect 12734 18765 12740 18817
rect 12610 18737 12740 18765
rect 12610 18685 12616 18737
rect 12668 18685 12682 18737
rect 12734 18685 12740 18737
rect 8194 8785 8203 8841
rect 8259 8785 8287 8841
rect 8343 8785 8370 8841
rect 8426 8785 8453 8841
rect 8509 8785 8536 8841
rect 8592 8785 8619 8841
rect 8675 8785 8702 8841
rect 8758 8785 8785 8841
rect 8841 8785 8868 8841
rect 8924 8785 8951 8841
rect 9007 8785 9034 8841
rect 9090 8785 9117 8841
rect 9173 8785 9200 8841
rect 9256 8785 9265 8841
rect 8194 8755 9265 8785
rect 8194 8699 8203 8755
rect 8259 8699 8287 8755
rect 8343 8699 8370 8755
rect 8426 8699 8453 8755
rect 8509 8699 8536 8755
rect 8592 8699 8619 8755
rect 8675 8699 8702 8755
rect 8758 8699 8785 8755
rect 8841 8699 8868 8755
rect 8924 8699 8951 8755
rect 9007 8699 9034 8755
rect 9090 8699 9117 8755
rect 9173 8699 9200 8755
rect 9256 8699 9265 8755
rect 8194 8669 9265 8699
rect 8194 8613 8203 8669
rect 8259 8613 8287 8669
rect 8343 8613 8370 8669
rect 8426 8613 8453 8669
rect 8509 8613 8536 8669
rect 8592 8613 8619 8669
rect 8675 8613 8702 8669
rect 8758 8613 8785 8669
rect 8841 8613 8868 8669
rect 8924 8613 8951 8669
rect 9007 8613 9034 8669
rect 9090 8613 9117 8669
rect 9173 8613 9200 8669
rect 9256 8613 9265 8669
rect 8194 8583 9265 8613
rect 8194 8527 8203 8583
rect 8259 8527 8287 8583
rect 8343 8527 8370 8583
rect 8426 8527 8453 8583
rect 8509 8527 8536 8583
rect 8592 8527 8619 8583
rect 8675 8527 8702 8583
rect 8758 8527 8785 8583
rect 8841 8527 8868 8583
rect 8924 8527 8951 8583
rect 9007 8527 9034 8583
rect 9090 8527 9117 8583
rect 9173 8527 9200 8583
rect 9256 8527 9265 8583
rect 8194 8497 9265 8527
rect 8194 8441 8203 8497
rect 8259 8441 8287 8497
rect 8343 8441 8370 8497
rect 8426 8441 8453 8497
rect 8509 8441 8536 8497
rect 8592 8441 8619 8497
rect 8675 8441 8702 8497
rect 8758 8441 8785 8497
rect 8841 8441 8868 8497
rect 8924 8441 8951 8497
rect 9007 8441 9034 8497
rect 9090 8441 9117 8497
rect 9173 8441 9200 8497
rect 9256 8441 9265 8497
rect 8194 8411 9265 8441
rect 8194 8355 8203 8411
rect 8259 8355 8287 8411
rect 8343 8355 8370 8411
rect 8426 8355 8453 8411
rect 8509 8355 8536 8411
rect 8592 8355 8619 8411
rect 8675 8355 8702 8411
rect 8758 8355 8785 8411
rect 8841 8355 8868 8411
rect 8924 8355 8951 8411
rect 9007 8355 9034 8411
rect 9090 8355 9117 8411
rect 9173 8355 9200 8411
rect 9256 8355 9265 8411
rect 8194 8325 9265 8355
rect 8194 8269 8203 8325
rect 8259 8269 8287 8325
rect 8343 8269 8370 8325
rect 8426 8269 8453 8325
rect 8509 8269 8536 8325
rect 8592 8269 8619 8325
rect 8675 8269 8702 8325
rect 8758 8269 8785 8325
rect 8841 8269 8868 8325
rect 8924 8269 8951 8325
rect 9007 8269 9034 8325
rect 9090 8269 9117 8325
rect 9173 8269 9200 8325
rect 9256 8269 9265 8325
rect 8194 8239 9265 8269
rect 8194 8183 8203 8239
rect 8259 8183 8287 8239
rect 8343 8183 8370 8239
rect 8426 8183 8453 8239
rect 8509 8183 8536 8239
rect 8592 8183 8619 8239
rect 8675 8183 8702 8239
rect 8758 8183 8785 8239
rect 8841 8183 8868 8239
rect 8924 8183 8951 8239
rect 9007 8183 9034 8239
rect 9090 8183 9117 8239
rect 9173 8183 9200 8239
rect 9256 8183 9265 8239
rect 8194 8153 9265 8183
rect 8194 8097 8203 8153
rect 8259 8097 8287 8153
rect 8343 8097 8370 8153
rect 8426 8097 8453 8153
rect 8509 8097 8536 8153
rect 8592 8097 8619 8153
rect 8675 8097 8702 8153
rect 8758 8097 8785 8153
rect 8841 8097 8868 8153
rect 8924 8097 8951 8153
rect 9007 8097 9034 8153
rect 9090 8097 9117 8153
rect 9173 8097 9200 8153
rect 9256 8097 9265 8153
rect 8194 8067 9265 8097
rect 8194 8011 8203 8067
rect 8259 8011 8287 8067
rect 8343 8011 8370 8067
rect 8426 8011 8453 8067
rect 8509 8011 8536 8067
rect 8592 8011 8619 8067
rect 8675 8011 8702 8067
rect 8758 8011 8785 8067
rect 8841 8011 8868 8067
rect 8924 8011 8951 8067
rect 9007 8011 9034 8067
rect 9090 8011 9117 8067
rect 9173 8011 9200 8067
rect 9256 8011 9265 8067
rect 8194 7981 9265 8011
rect 8194 7925 8203 7981
rect 8259 7925 8287 7981
rect 8343 7925 8370 7981
rect 8426 7925 8453 7981
rect 8509 7925 8536 7981
rect 8592 7925 8619 7981
rect 8675 7925 8702 7981
rect 8758 7925 8785 7981
rect 8841 7925 8868 7981
rect 8924 7925 8951 7981
rect 9007 7925 9034 7981
rect 9090 7925 9117 7981
rect 9173 7925 9200 7981
rect 9256 7925 9265 7981
rect 8194 7916 9265 7925
<< via2 >>
rect 465 32708 521 32764
rect 623 32708 679 32764
rect 465 32627 521 32683
rect 623 32627 679 32683
rect 465 32545 521 32601
rect 623 32545 679 32601
rect 465 32463 521 32519
rect 623 32463 679 32519
rect 465 32381 521 32437
rect 623 32381 679 32437
rect 465 32299 521 32355
rect 623 32299 679 32355
rect 465 32217 521 32273
rect 623 32217 679 32273
rect 465 32135 521 32191
rect 623 32135 679 32191
rect 465 32053 521 32109
rect 623 32053 679 32109
rect 14259 32705 14315 32761
rect 14347 32705 14403 32761
rect 14435 32705 14491 32761
rect 14523 32705 14579 32761
rect 14611 32705 14667 32761
rect 14259 32625 14315 32681
rect 14347 32625 14403 32681
rect 14435 32625 14491 32681
rect 14523 32625 14579 32681
rect 14611 32625 14667 32681
rect 14259 32545 14315 32601
rect 14347 32545 14403 32601
rect 14435 32545 14491 32601
rect 14523 32545 14579 32601
rect 14611 32545 14667 32601
rect 14259 32465 14315 32521
rect 14347 32465 14403 32521
rect 14435 32465 14491 32521
rect 14523 32465 14579 32521
rect 14611 32465 14667 32521
rect 14259 32385 14315 32441
rect 14347 32385 14403 32441
rect 14435 32385 14491 32441
rect 14523 32385 14579 32441
rect 14611 32385 14667 32441
rect 14259 32305 14315 32361
rect 14347 32305 14403 32361
rect 14435 32305 14491 32361
rect 14523 32305 14579 32361
rect 14611 32305 14667 32361
rect 14259 32225 14315 32281
rect 14347 32225 14403 32281
rect 14435 32225 14491 32281
rect 14523 32225 14579 32281
rect 14611 32225 14667 32281
rect 14259 32145 14315 32201
rect 14347 32145 14403 32201
rect 14435 32145 14491 32201
rect 14523 32145 14579 32201
rect 14611 32145 14667 32201
rect 14259 32065 14315 32121
rect 14347 32065 14403 32121
rect 14435 32065 14491 32121
rect 14523 32065 14579 32121
rect 14611 32065 14667 32121
rect 465 31971 521 32027
rect 623 31971 679 32027
rect 465 31889 521 31945
rect 623 31889 679 31945
rect 465 31807 521 31863
rect 623 31807 679 31863
rect 465 31725 521 31781
rect 623 31725 679 31781
rect 465 31643 521 31699
rect 623 31643 679 31699
rect 465 31561 521 31617
rect 623 31561 679 31617
rect 465 31479 521 31535
rect 623 31479 679 31535
rect 465 31397 521 31453
rect 623 31397 679 31453
rect 465 31315 521 31371
rect 623 31315 679 31371
rect 465 31233 521 31289
rect 623 31233 679 31289
rect 465 31151 521 31207
rect 623 31151 679 31207
rect 465 31069 521 31125
rect 623 31069 679 31125
rect 465 30987 521 31043
rect 623 30987 679 31043
rect 465 30905 521 30961
rect 623 30905 679 30961
rect 465 30823 521 30879
rect 623 30823 679 30879
rect 465 30741 521 30797
rect 623 30741 679 30797
rect 465 30659 521 30715
rect 623 30659 679 30715
rect 465 30577 521 30633
rect 623 30577 679 30633
rect 465 30495 521 30551
rect 623 30495 679 30551
rect 465 30413 521 30469
rect 623 30413 679 30469
rect 465 30331 521 30387
rect 623 30331 679 30387
rect 465 30249 521 30305
rect 623 30249 679 30305
rect 465 30167 521 30223
rect 623 30167 679 30223
rect 465 30085 521 30141
rect 623 30085 679 30141
rect 465 30003 521 30059
rect 623 30003 679 30059
rect 465 29921 521 29977
rect 623 29921 679 29977
rect 465 29839 521 29895
rect 623 29839 679 29895
rect 465 29757 521 29813
rect 623 29757 679 29813
rect 465 29675 521 29731
rect 623 29675 679 29731
rect 465 29593 521 29649
rect 623 29593 679 29649
rect 465 29511 521 29567
rect 623 29511 679 29567
rect 465 29429 521 29485
rect 623 29429 679 29485
rect 862 31962 918 32018
rect 996 31962 1052 32018
rect 862 31880 918 31936
rect 996 31880 1052 31936
rect 862 31798 918 31854
rect 996 31798 1052 31854
rect 862 31716 918 31772
rect 996 31716 1052 31772
rect 862 31634 918 31690
rect 996 31634 1052 31690
rect 862 31552 918 31608
rect 996 31552 1052 31608
rect 862 31470 918 31526
rect 996 31470 1052 31526
rect 862 31388 918 31444
rect 996 31388 1052 31444
rect 862 31306 918 31362
rect 996 31306 1052 31362
rect 862 31224 918 31280
rect 996 31224 1052 31280
rect 862 31142 918 31198
rect 996 31142 1052 31198
rect 862 31060 918 31116
rect 996 31060 1052 31116
rect 862 30978 918 31034
rect 996 30978 1052 31034
rect 862 30896 918 30952
rect 996 30896 1052 30952
rect 862 30814 918 30870
rect 996 30814 1052 30870
rect 862 30732 918 30788
rect 996 30732 1052 30788
rect 862 30650 918 30706
rect 996 30650 1052 30706
rect 862 30568 918 30624
rect 996 30568 1052 30624
rect 862 30486 918 30542
rect 996 30486 1052 30542
rect 862 30404 918 30460
rect 996 30404 1052 30460
rect 862 30322 918 30378
rect 996 30322 1052 30378
rect 862 30240 918 30296
rect 996 30240 1052 30296
rect 862 30158 918 30214
rect 996 30158 1052 30214
rect 862 30076 918 30132
rect 996 30076 1052 30132
rect 862 29994 918 30050
rect 996 29994 1052 30050
rect 862 29912 918 29968
rect 996 29912 1052 29968
rect 862 29830 918 29886
rect 996 29830 1052 29886
rect 862 29748 918 29804
rect 996 29748 1052 29804
rect 862 29666 918 29722
rect 996 29666 1052 29722
rect 862 29584 918 29640
rect 996 29584 1052 29640
rect 862 29502 918 29558
rect 996 29502 1052 29558
rect 862 29420 918 29476
rect 996 29420 1052 29476
rect 1395 31962 1451 32018
rect 1521 31962 1577 32018
rect 1395 31881 1451 31937
rect 1521 31881 1577 31937
rect 1395 31800 1451 31856
rect 1521 31800 1577 31856
rect 1395 31719 1451 31775
rect 1521 31719 1577 31775
rect 1395 31638 1451 31694
rect 1521 31638 1577 31694
rect 1395 31557 1451 31613
rect 1521 31557 1577 31613
rect 1395 31476 1451 31532
rect 1521 31476 1577 31532
rect 1395 31395 1451 31451
rect 1521 31395 1577 31451
rect 1395 31314 1451 31370
rect 1521 31314 1577 31370
rect 1395 31233 1451 31289
rect 1521 31233 1577 31289
rect 1395 31151 1451 31207
rect 1521 31151 1577 31207
rect 1395 31069 1451 31125
rect 1521 31069 1577 31125
rect 1395 30987 1451 31043
rect 1521 30987 1577 31043
rect 1395 30905 1451 30961
rect 1521 30905 1577 30961
rect 1395 30823 1451 30879
rect 1521 30823 1577 30879
rect 1395 30741 1451 30797
rect 1521 30741 1577 30797
rect 1395 30659 1451 30715
rect 1521 30659 1577 30715
rect 1395 30577 1451 30633
rect 1521 30577 1577 30633
rect 1395 30495 1451 30551
rect 1521 30495 1577 30551
rect 1395 30413 1451 30469
rect 1521 30413 1577 30469
rect 1395 30331 1451 30387
rect 1521 30331 1577 30387
rect 1395 30249 1451 30305
rect 1521 30249 1577 30305
rect 1395 30167 1451 30223
rect 1521 30167 1577 30223
rect 1395 30085 1451 30141
rect 1521 30085 1577 30141
rect 1395 30003 1451 30059
rect 1521 30003 1577 30059
rect 1395 29921 1451 29977
rect 1521 29921 1577 29977
rect 1395 29839 1451 29895
rect 1521 29839 1577 29895
rect 1395 29757 1451 29813
rect 1521 29757 1577 29813
rect 1395 29675 1451 29731
rect 1521 29675 1577 29731
rect 1395 29593 1451 29649
rect 1521 29593 1577 29649
rect 1395 29511 1451 29567
rect 1521 29511 1577 29567
rect 1395 29429 1451 29485
rect 1521 29429 1577 29485
rect 1891 31962 1947 32018
rect 2017 31962 2073 32018
rect 1891 31880 1947 31936
rect 2017 31880 2073 31936
rect 1891 31798 1947 31854
rect 2017 31798 2073 31854
rect 1891 31716 1947 31772
rect 2017 31716 2073 31772
rect 1891 31634 1947 31690
rect 2017 31634 2073 31690
rect 1891 31552 1947 31608
rect 2017 31552 2073 31608
rect 1891 31470 1947 31526
rect 2017 31470 2073 31526
rect 1891 31388 1947 31444
rect 2017 31388 2073 31444
rect 1891 31306 1947 31362
rect 2017 31306 2073 31362
rect 1891 31224 1947 31280
rect 2017 31224 2073 31280
rect 1891 31142 1947 31198
rect 2017 31142 2073 31198
rect 1891 31060 1947 31116
rect 2017 31060 2073 31116
rect 1891 30978 1947 31034
rect 2017 30978 2073 31034
rect 1891 30896 1947 30952
rect 2017 30896 2073 30952
rect 1891 30814 1947 30870
rect 2017 30814 2073 30870
rect 1891 30732 1947 30788
rect 2017 30732 2073 30788
rect 1891 30650 1947 30706
rect 2017 30650 2073 30706
rect 1891 30568 1947 30624
rect 2017 30568 2073 30624
rect 1891 30486 1947 30542
rect 2017 30486 2073 30542
rect 1891 30404 1947 30460
rect 2017 30404 2073 30460
rect 1891 30322 1947 30378
rect 2017 30322 2073 30378
rect 1891 30240 1947 30296
rect 2017 30240 2073 30296
rect 1891 30158 1947 30214
rect 2017 30158 2073 30214
rect 1891 30076 1947 30132
rect 2017 30076 2073 30132
rect 1891 29994 1947 30050
rect 2017 29994 2073 30050
rect 1891 29912 1947 29968
rect 2017 29912 2073 29968
rect 1891 29830 1947 29886
rect 2017 29830 2073 29886
rect 1891 29748 1947 29804
rect 2017 29748 2073 29804
rect 1891 29666 1947 29722
rect 2017 29666 2073 29722
rect 1891 29584 1947 29640
rect 2017 29584 2073 29640
rect 1891 29502 1947 29558
rect 2017 29502 2073 29558
rect 1891 29420 1947 29476
rect 2017 29420 2073 29476
rect 2387 31962 2443 32018
rect 2513 31962 2569 32018
rect 2387 31880 2443 31936
rect 2513 31880 2569 31936
rect 2387 31798 2443 31854
rect 2513 31798 2569 31854
rect 2387 31716 2443 31772
rect 2513 31716 2569 31772
rect 2387 31634 2443 31690
rect 2513 31634 2569 31690
rect 2387 31552 2443 31608
rect 2513 31552 2569 31608
rect 2387 31470 2443 31526
rect 2513 31470 2569 31526
rect 2387 31388 2443 31444
rect 2513 31388 2569 31444
rect 2387 31306 2443 31362
rect 2513 31306 2569 31362
rect 2387 31224 2443 31280
rect 2513 31224 2569 31280
rect 2387 31142 2443 31198
rect 2513 31142 2569 31198
rect 2387 31060 2443 31116
rect 2513 31060 2569 31116
rect 2387 30978 2443 31034
rect 2513 30978 2569 31034
rect 2387 30896 2443 30952
rect 2513 30896 2569 30952
rect 2387 30814 2443 30870
rect 2513 30814 2569 30870
rect 2387 30732 2443 30788
rect 2513 30732 2569 30788
rect 2387 30650 2443 30706
rect 2513 30650 2569 30706
rect 2387 30568 2443 30624
rect 2513 30568 2569 30624
rect 2387 30486 2443 30542
rect 2513 30486 2569 30542
rect 2387 30404 2443 30460
rect 2513 30404 2569 30460
rect 2387 30322 2443 30378
rect 2513 30322 2569 30378
rect 2387 30240 2443 30296
rect 2513 30240 2569 30296
rect 2387 30158 2443 30214
rect 2513 30158 2569 30214
rect 2387 30076 2443 30132
rect 2513 30076 2569 30132
rect 2387 29994 2443 30050
rect 2513 29994 2569 30050
rect 2387 29912 2443 29968
rect 2513 29912 2569 29968
rect 2387 29830 2443 29886
rect 2513 29830 2569 29886
rect 2387 29748 2443 29804
rect 2513 29748 2569 29804
rect 2387 29666 2443 29722
rect 2513 29666 2569 29722
rect 2387 29584 2443 29640
rect 2513 29584 2569 29640
rect 2387 29502 2443 29558
rect 2513 29502 2569 29558
rect 2387 29420 2443 29476
rect 2513 29420 2569 29476
rect 2883 31962 2939 32018
rect 3009 31962 3065 32018
rect 2883 31880 2939 31936
rect 3009 31880 3065 31936
rect 2883 31798 2939 31854
rect 3009 31798 3065 31854
rect 2883 31716 2939 31772
rect 3009 31716 3065 31772
rect 2883 31634 2939 31690
rect 3009 31634 3065 31690
rect 2883 31552 2939 31608
rect 3009 31552 3065 31608
rect 2883 31470 2939 31526
rect 3009 31470 3065 31526
rect 2883 31388 2939 31444
rect 3009 31388 3065 31444
rect 2883 31306 2939 31362
rect 3009 31306 3065 31362
rect 2883 31224 2939 31280
rect 3009 31224 3065 31280
rect 2883 31142 2939 31198
rect 3009 31142 3065 31198
rect 2883 31060 2939 31116
rect 3009 31060 3065 31116
rect 2883 30978 2939 31034
rect 3009 30978 3065 31034
rect 2883 30896 2939 30952
rect 3009 30896 3065 30952
rect 2883 30814 2939 30870
rect 3009 30814 3065 30870
rect 2883 30732 2939 30788
rect 3009 30732 3065 30788
rect 2883 30650 2939 30706
rect 3009 30650 3065 30706
rect 2883 30568 2939 30624
rect 3009 30568 3065 30624
rect 2883 30486 2939 30542
rect 3009 30486 3065 30542
rect 2883 30404 2939 30460
rect 3009 30404 3065 30460
rect 2883 30322 2939 30378
rect 3009 30322 3065 30378
rect 2883 30240 2939 30296
rect 3009 30240 3065 30296
rect 2883 30158 2939 30214
rect 3009 30158 3065 30214
rect 2883 30076 2939 30132
rect 3009 30076 3065 30132
rect 2883 29994 2939 30050
rect 3009 29994 3065 30050
rect 2883 29912 2939 29968
rect 3009 29912 3065 29968
rect 2883 29830 2939 29886
rect 3009 29830 3065 29886
rect 2883 29748 2939 29804
rect 3009 29748 3065 29804
rect 2883 29666 2939 29722
rect 3009 29666 3065 29722
rect 2883 29584 2939 29640
rect 3009 29584 3065 29640
rect 2883 29502 2939 29558
rect 3009 29502 3065 29558
rect 2883 29420 2939 29476
rect 3009 29420 3065 29476
rect 3379 31962 3435 32018
rect 3505 31962 3561 32018
rect 3379 31880 3435 31936
rect 3505 31880 3561 31936
rect 3379 31798 3435 31854
rect 3505 31798 3561 31854
rect 3379 31716 3435 31772
rect 3505 31716 3561 31772
rect 3379 31634 3435 31690
rect 3505 31634 3561 31690
rect 3379 31552 3435 31608
rect 3505 31552 3561 31608
rect 3379 31470 3435 31526
rect 3505 31470 3561 31526
rect 3379 31388 3435 31444
rect 3505 31388 3561 31444
rect 3379 31306 3435 31362
rect 3505 31306 3561 31362
rect 3379 31224 3435 31280
rect 3505 31224 3561 31280
rect 3379 31142 3435 31198
rect 3505 31142 3561 31198
rect 3379 31060 3435 31116
rect 3505 31060 3561 31116
rect 3379 30978 3435 31034
rect 3505 30978 3561 31034
rect 3379 30896 3435 30952
rect 3505 30896 3561 30952
rect 3379 30814 3435 30870
rect 3505 30814 3561 30870
rect 3379 30732 3435 30788
rect 3505 30732 3561 30788
rect 3379 30650 3435 30706
rect 3505 30650 3561 30706
rect 3379 30568 3435 30624
rect 3505 30568 3561 30624
rect 3379 30486 3435 30542
rect 3505 30486 3561 30542
rect 3379 30404 3435 30460
rect 3505 30404 3561 30460
rect 3379 30322 3435 30378
rect 3505 30322 3561 30378
rect 3379 30240 3435 30296
rect 3505 30240 3561 30296
rect 3379 30158 3435 30214
rect 3505 30158 3561 30214
rect 3379 30076 3435 30132
rect 3505 30076 3561 30132
rect 3379 29994 3435 30050
rect 3505 29994 3561 30050
rect 3379 29912 3435 29968
rect 3505 29912 3561 29968
rect 3379 29830 3435 29886
rect 3505 29830 3561 29886
rect 3379 29748 3435 29804
rect 3505 29748 3561 29804
rect 3379 29666 3435 29722
rect 3505 29666 3561 29722
rect 3379 29584 3435 29640
rect 3505 29584 3561 29640
rect 3379 29502 3435 29558
rect 3505 29502 3561 29558
rect 3379 29420 3435 29476
rect 3505 29420 3561 29476
rect 3875 31962 3931 32018
rect 4001 31962 4057 32018
rect 3875 31880 3931 31936
rect 4001 31880 4057 31936
rect 3875 31798 3931 31854
rect 4001 31798 4057 31854
rect 3875 31716 3931 31772
rect 4001 31716 4057 31772
rect 3875 31634 3931 31690
rect 4001 31634 4057 31690
rect 3875 31552 3931 31608
rect 4001 31552 4057 31608
rect 3875 31470 3931 31526
rect 4001 31470 4057 31526
rect 3875 31388 3931 31444
rect 4001 31388 4057 31444
rect 3875 31306 3931 31362
rect 4001 31306 4057 31362
rect 3875 31224 3931 31280
rect 4001 31224 4057 31280
rect 3875 31142 3931 31198
rect 4001 31142 4057 31198
rect 3875 31060 3931 31116
rect 4001 31060 4057 31116
rect 3875 30978 3931 31034
rect 4001 30978 4057 31034
rect 3875 30896 3931 30952
rect 4001 30896 4057 30952
rect 3875 30814 3931 30870
rect 4001 30814 4057 30870
rect 3875 30732 3931 30788
rect 4001 30732 4057 30788
rect 3875 30650 3931 30706
rect 4001 30650 4057 30706
rect 3875 30568 3931 30624
rect 4001 30568 4057 30624
rect 3875 30486 3931 30542
rect 4001 30486 4057 30542
rect 3875 30404 3931 30460
rect 4001 30404 4057 30460
rect 3875 30322 3931 30378
rect 4001 30322 4057 30378
rect 3875 30240 3931 30296
rect 4001 30240 4057 30296
rect 3875 30158 3931 30214
rect 4001 30158 4057 30214
rect 3875 30076 3931 30132
rect 4001 30076 4057 30132
rect 3875 29994 3931 30050
rect 4001 29994 4057 30050
rect 3875 29912 3931 29968
rect 4001 29912 4057 29968
rect 3875 29830 3931 29886
rect 4001 29830 4057 29886
rect 3875 29748 3931 29804
rect 4001 29748 4057 29804
rect 3875 29666 3931 29722
rect 4001 29666 4057 29722
rect 3875 29584 3931 29640
rect 4001 29584 4057 29640
rect 3875 29502 3931 29558
rect 4001 29502 4057 29558
rect 3875 29420 3931 29476
rect 4001 29420 4057 29476
rect 4371 31962 4427 32018
rect 4497 31962 4553 32018
rect 4371 31880 4427 31936
rect 4497 31880 4553 31936
rect 4371 31798 4427 31854
rect 4497 31798 4553 31854
rect 4371 31716 4427 31772
rect 4497 31716 4553 31772
rect 4371 31634 4427 31690
rect 4497 31634 4553 31690
rect 4371 31552 4427 31608
rect 4497 31552 4553 31608
rect 4371 31470 4427 31526
rect 4497 31470 4553 31526
rect 4371 31388 4427 31444
rect 4497 31388 4553 31444
rect 4371 31306 4427 31362
rect 4497 31306 4553 31362
rect 4371 31224 4427 31280
rect 4497 31224 4553 31280
rect 4371 31142 4427 31198
rect 4497 31142 4553 31198
rect 4371 31060 4427 31116
rect 4497 31060 4553 31116
rect 4371 30978 4427 31034
rect 4497 30978 4553 31034
rect 4371 30896 4427 30952
rect 4497 30896 4553 30952
rect 4371 30814 4427 30870
rect 4497 30814 4553 30870
rect 4371 30732 4427 30788
rect 4497 30732 4553 30788
rect 4371 30650 4427 30706
rect 4497 30650 4553 30706
rect 4371 30568 4427 30624
rect 4497 30568 4553 30624
rect 4371 30486 4427 30542
rect 4497 30486 4553 30542
rect 4371 30404 4427 30460
rect 4497 30404 4553 30460
rect 4371 30322 4427 30378
rect 4497 30322 4553 30378
rect 4371 30240 4427 30296
rect 4497 30240 4553 30296
rect 4371 30158 4427 30214
rect 4497 30158 4553 30214
rect 4371 30076 4427 30132
rect 4497 30076 4553 30132
rect 4371 29994 4427 30050
rect 4497 29994 4553 30050
rect 4371 29912 4427 29968
rect 4497 29912 4553 29968
rect 4371 29830 4427 29886
rect 4497 29830 4553 29886
rect 4371 29748 4427 29804
rect 4497 29748 4553 29804
rect 4371 29666 4427 29722
rect 4497 29666 4553 29722
rect 4371 29584 4427 29640
rect 4497 29584 4553 29640
rect 4371 29502 4427 29558
rect 4497 29502 4553 29558
rect 4371 29420 4427 29476
rect 4497 29420 4553 29476
rect 4867 31962 4923 32018
rect 4993 31962 5049 32018
rect 4867 31880 4923 31936
rect 4993 31880 5049 31936
rect 4867 31798 4923 31854
rect 4993 31798 5049 31854
rect 4867 31716 4923 31772
rect 4993 31716 5049 31772
rect 4867 31634 4923 31690
rect 4993 31634 5049 31690
rect 4867 31552 4923 31608
rect 4993 31552 5049 31608
rect 4867 31470 4923 31526
rect 4993 31470 5049 31526
rect 4867 31388 4923 31444
rect 4993 31388 5049 31444
rect 4867 31306 4923 31362
rect 4993 31306 5049 31362
rect 4867 31224 4923 31280
rect 4993 31224 5049 31280
rect 4867 31142 4923 31198
rect 4993 31142 5049 31198
rect 4867 31060 4923 31116
rect 4993 31060 5049 31116
rect 4867 30978 4923 31034
rect 4993 30978 5049 31034
rect 4867 30896 4923 30952
rect 4993 30896 5049 30952
rect 4867 30814 4923 30870
rect 4993 30814 5049 30870
rect 4867 30732 4923 30788
rect 4993 30732 5049 30788
rect 4867 30650 4923 30706
rect 4993 30650 5049 30706
rect 4867 30568 4923 30624
rect 4993 30568 5049 30624
rect 4867 30486 4923 30542
rect 4993 30486 5049 30542
rect 4867 30404 4923 30460
rect 4993 30404 5049 30460
rect 4867 30322 4923 30378
rect 4993 30322 5049 30378
rect 4867 30240 4923 30296
rect 4993 30240 5049 30296
rect 4867 30158 4923 30214
rect 4993 30158 5049 30214
rect 4867 30076 4923 30132
rect 4993 30076 5049 30132
rect 4867 29994 4923 30050
rect 4993 29994 5049 30050
rect 4867 29912 4923 29968
rect 4993 29912 5049 29968
rect 4867 29830 4923 29886
rect 4993 29830 5049 29886
rect 4867 29748 4923 29804
rect 4993 29748 5049 29804
rect 4867 29666 4923 29722
rect 4993 29666 5049 29722
rect 4867 29584 4923 29640
rect 4993 29584 5049 29640
rect 4867 29502 4923 29558
rect 4993 29502 5049 29558
rect 4867 29420 4923 29476
rect 4993 29420 5049 29476
rect 5363 31962 5419 32018
rect 5489 31962 5545 32018
rect 5363 31880 5419 31936
rect 5489 31880 5545 31936
rect 5363 31798 5419 31854
rect 5489 31798 5545 31854
rect 5363 31716 5419 31772
rect 5489 31716 5545 31772
rect 5363 31634 5419 31690
rect 5489 31634 5545 31690
rect 5363 31552 5419 31608
rect 5489 31552 5545 31608
rect 5363 31470 5419 31526
rect 5489 31470 5545 31526
rect 5363 31388 5419 31444
rect 5489 31388 5545 31444
rect 5363 31306 5419 31362
rect 5489 31306 5545 31362
rect 5363 31224 5419 31280
rect 5489 31224 5545 31280
rect 5363 31142 5419 31198
rect 5489 31142 5545 31198
rect 5363 31060 5419 31116
rect 5489 31060 5545 31116
rect 5363 30978 5419 31034
rect 5489 30978 5545 31034
rect 5363 30896 5419 30952
rect 5489 30896 5545 30952
rect 5363 30814 5419 30870
rect 5489 30814 5545 30870
rect 5363 30732 5419 30788
rect 5489 30732 5545 30788
rect 5363 30650 5419 30706
rect 5489 30650 5545 30706
rect 5363 30568 5419 30624
rect 5489 30568 5545 30624
rect 5363 30486 5419 30542
rect 5489 30486 5545 30542
rect 5363 30404 5419 30460
rect 5489 30404 5545 30460
rect 5363 30322 5419 30378
rect 5489 30322 5545 30378
rect 5363 30240 5419 30296
rect 5489 30240 5545 30296
rect 5363 30158 5419 30214
rect 5489 30158 5545 30214
rect 5363 30076 5419 30132
rect 5489 30076 5545 30132
rect 5363 29994 5419 30050
rect 5489 29994 5545 30050
rect 5363 29912 5419 29968
rect 5489 29912 5545 29968
rect 5363 29830 5419 29886
rect 5489 29830 5545 29886
rect 5363 29748 5419 29804
rect 5489 29748 5545 29804
rect 5363 29666 5419 29722
rect 5489 29666 5545 29722
rect 5363 29584 5419 29640
rect 5489 29584 5545 29640
rect 5363 29502 5419 29558
rect 5489 29502 5545 29558
rect 5363 29420 5419 29476
rect 5489 29420 5545 29476
rect 5859 31962 5915 32018
rect 5985 31962 6041 32018
rect 5859 31880 5915 31936
rect 5985 31880 6041 31936
rect 5859 31798 5915 31854
rect 5985 31798 6041 31854
rect 5859 31716 5915 31772
rect 5985 31716 6041 31772
rect 5859 31634 5915 31690
rect 5985 31634 6041 31690
rect 5859 31552 5915 31608
rect 5985 31552 6041 31608
rect 5859 31470 5915 31526
rect 5985 31470 6041 31526
rect 5859 31388 5915 31444
rect 5985 31388 6041 31444
rect 5859 31306 5915 31362
rect 5985 31306 6041 31362
rect 5859 31224 5915 31280
rect 5985 31224 6041 31280
rect 5859 31142 5915 31198
rect 5985 31142 6041 31198
rect 5859 31060 5915 31116
rect 5985 31060 6041 31116
rect 5859 30978 5915 31034
rect 5985 30978 6041 31034
rect 5859 30896 5915 30952
rect 5985 30896 6041 30952
rect 5859 30814 5915 30870
rect 5985 30814 6041 30870
rect 5859 30732 5915 30788
rect 5985 30732 6041 30788
rect 5859 30650 5915 30706
rect 5985 30650 6041 30706
rect 5859 30568 5915 30624
rect 5985 30568 6041 30624
rect 5859 30486 5915 30542
rect 5985 30486 6041 30542
rect 5859 30404 5915 30460
rect 5985 30404 6041 30460
rect 5859 30322 5915 30378
rect 5985 30322 6041 30378
rect 5859 30240 5915 30296
rect 5985 30240 6041 30296
rect 5859 30158 5915 30214
rect 5985 30158 6041 30214
rect 5859 30076 5915 30132
rect 5985 30076 6041 30132
rect 5859 29994 5915 30050
rect 5985 29994 6041 30050
rect 5859 29912 5915 29968
rect 5985 29912 6041 29968
rect 5859 29830 5915 29886
rect 5985 29830 6041 29886
rect 5859 29748 5915 29804
rect 5985 29748 6041 29804
rect 5859 29666 5915 29722
rect 5985 29666 6041 29722
rect 5859 29584 5915 29640
rect 5985 29584 6041 29640
rect 5859 29502 5915 29558
rect 5985 29502 6041 29558
rect 5859 29420 5915 29476
rect 5985 29420 6041 29476
rect 6355 31962 6411 32018
rect 6481 31962 6537 32018
rect 6355 31880 6411 31936
rect 6481 31880 6537 31936
rect 6355 31798 6411 31854
rect 6481 31798 6537 31854
rect 6355 31716 6411 31772
rect 6481 31716 6537 31772
rect 6355 31634 6411 31690
rect 6481 31634 6537 31690
rect 6355 31552 6411 31608
rect 6481 31552 6537 31608
rect 6355 31470 6411 31526
rect 6481 31470 6537 31526
rect 6355 31388 6411 31444
rect 6481 31388 6537 31444
rect 6355 31306 6411 31362
rect 6481 31306 6537 31362
rect 6355 31224 6411 31280
rect 6481 31224 6537 31280
rect 6355 31142 6411 31198
rect 6481 31142 6537 31198
rect 6355 31060 6411 31116
rect 6481 31060 6537 31116
rect 6355 30978 6411 31034
rect 6481 30978 6537 31034
rect 6355 30896 6411 30952
rect 6481 30896 6537 30952
rect 6355 30814 6411 30870
rect 6481 30814 6537 30870
rect 6355 30732 6411 30788
rect 6481 30732 6537 30788
rect 6355 30650 6411 30706
rect 6481 30650 6537 30706
rect 6355 30568 6411 30624
rect 6481 30568 6537 30624
rect 6355 30486 6411 30542
rect 6481 30486 6537 30542
rect 6355 30404 6411 30460
rect 6481 30404 6537 30460
rect 6355 30322 6411 30378
rect 6481 30322 6537 30378
rect 6355 30240 6411 30296
rect 6481 30240 6537 30296
rect 6355 30158 6411 30214
rect 6481 30158 6537 30214
rect 6355 30076 6411 30132
rect 6481 30076 6537 30132
rect 6355 29994 6411 30050
rect 6481 29994 6537 30050
rect 6355 29912 6411 29968
rect 6481 29912 6537 29968
rect 6355 29830 6411 29886
rect 6481 29830 6537 29886
rect 6355 29748 6411 29804
rect 6481 29748 6537 29804
rect 6355 29666 6411 29722
rect 6481 29666 6537 29722
rect 6355 29584 6411 29640
rect 6481 29584 6537 29640
rect 6355 29502 6411 29558
rect 6481 29502 6537 29558
rect 6355 29420 6411 29476
rect 6481 29420 6537 29476
rect 6851 31962 6907 32018
rect 6977 31962 7033 32018
rect 6851 31880 6907 31936
rect 6977 31880 7033 31936
rect 6851 31798 6907 31854
rect 6977 31798 7033 31854
rect 6851 31716 6907 31772
rect 6977 31716 7033 31772
rect 6851 31634 6907 31690
rect 6977 31634 7033 31690
rect 6851 31552 6907 31608
rect 6977 31552 7033 31608
rect 6851 31470 6907 31526
rect 6977 31470 7033 31526
rect 6851 31388 6907 31444
rect 6977 31388 7033 31444
rect 6851 31306 6907 31362
rect 6977 31306 7033 31362
rect 6851 31224 6907 31280
rect 6977 31224 7033 31280
rect 6851 31142 6907 31198
rect 6977 31142 7033 31198
rect 6851 31060 6907 31116
rect 6977 31060 7033 31116
rect 6851 30978 6907 31034
rect 6977 30978 7033 31034
rect 6851 30896 6907 30952
rect 6977 30896 7033 30952
rect 6851 30814 6907 30870
rect 6977 30814 7033 30870
rect 6851 30732 6907 30788
rect 6977 30732 7033 30788
rect 6851 30650 6907 30706
rect 6977 30650 7033 30706
rect 6851 30568 6907 30624
rect 6977 30568 7033 30624
rect 6851 30486 6907 30542
rect 6977 30486 7033 30542
rect 6851 30404 6907 30460
rect 6977 30404 7033 30460
rect 6851 30322 6907 30378
rect 6977 30322 7033 30378
rect 6851 30240 6907 30296
rect 6977 30240 7033 30296
rect 6851 30158 6907 30214
rect 6977 30158 7033 30214
rect 6851 30076 6907 30132
rect 6977 30076 7033 30132
rect 6851 29994 6907 30050
rect 6977 29994 7033 30050
rect 6851 29912 6907 29968
rect 6977 29912 7033 29968
rect 6851 29830 6907 29886
rect 6977 29830 7033 29886
rect 6851 29748 6907 29804
rect 6977 29748 7033 29804
rect 6851 29666 6907 29722
rect 6977 29666 7033 29722
rect 6851 29584 6907 29640
rect 6977 29584 7033 29640
rect 6851 29502 6907 29558
rect 6977 29502 7033 29558
rect 6851 29420 6907 29476
rect 6977 29420 7033 29476
rect 7347 31962 7403 32018
rect 7473 31962 7529 32018
rect 7347 31880 7403 31936
rect 7473 31880 7529 31936
rect 7347 31798 7403 31854
rect 7473 31798 7529 31854
rect 7347 31716 7403 31772
rect 7473 31716 7529 31772
rect 7347 31634 7403 31690
rect 7473 31634 7529 31690
rect 7347 31552 7403 31608
rect 7473 31552 7529 31608
rect 7347 31470 7403 31526
rect 7473 31470 7529 31526
rect 7347 31388 7403 31444
rect 7473 31388 7529 31444
rect 7347 31306 7403 31362
rect 7473 31306 7529 31362
rect 7347 31224 7403 31280
rect 7473 31224 7529 31280
rect 7347 31142 7403 31198
rect 7473 31142 7529 31198
rect 7347 31060 7403 31116
rect 7473 31060 7529 31116
rect 7347 30978 7403 31034
rect 7473 30978 7529 31034
rect 7347 30896 7403 30952
rect 7473 30896 7529 30952
rect 7347 30814 7403 30870
rect 7473 30814 7529 30870
rect 7347 30732 7403 30788
rect 7473 30732 7529 30788
rect 7347 30650 7403 30706
rect 7473 30650 7529 30706
rect 7347 30568 7403 30624
rect 7473 30568 7529 30624
rect 7347 30486 7403 30542
rect 7473 30486 7529 30542
rect 7347 30404 7403 30460
rect 7473 30404 7529 30460
rect 7347 30322 7403 30378
rect 7473 30322 7529 30378
rect 7347 30240 7403 30296
rect 7473 30240 7529 30296
rect 7347 30158 7403 30214
rect 7473 30158 7529 30214
rect 7347 30076 7403 30132
rect 7473 30076 7529 30132
rect 7347 29994 7403 30050
rect 7473 29994 7529 30050
rect 7347 29912 7403 29968
rect 7473 29912 7529 29968
rect 7347 29830 7403 29886
rect 7473 29830 7529 29886
rect 7347 29748 7403 29804
rect 7473 29748 7529 29804
rect 7347 29666 7403 29722
rect 7473 29666 7529 29722
rect 7347 29584 7403 29640
rect 7473 29584 7529 29640
rect 7347 29502 7403 29558
rect 7473 29502 7529 29558
rect 7347 29420 7403 29476
rect 7473 29420 7529 29476
rect 7843 31962 7899 32018
rect 7969 31962 8025 32018
rect 7843 31880 7899 31936
rect 7969 31880 8025 31936
rect 7843 31798 7899 31854
rect 7969 31798 8025 31854
rect 7843 31716 7899 31772
rect 7969 31716 8025 31772
rect 7843 31634 7899 31690
rect 7969 31634 8025 31690
rect 7843 31552 7899 31608
rect 7969 31552 8025 31608
rect 7843 31470 7899 31526
rect 7969 31470 8025 31526
rect 7843 31388 7899 31444
rect 7969 31388 8025 31444
rect 7843 31306 7899 31362
rect 7969 31306 8025 31362
rect 7843 31224 7899 31280
rect 7969 31224 8025 31280
rect 7843 31142 7899 31198
rect 7969 31142 8025 31198
rect 7843 31060 7899 31116
rect 7969 31060 8025 31116
rect 7843 30978 7899 31034
rect 7969 30978 8025 31034
rect 7843 30896 7899 30952
rect 7969 30896 8025 30952
rect 7843 30814 7899 30870
rect 7969 30814 8025 30870
rect 7843 30732 7899 30788
rect 7969 30732 8025 30788
rect 7843 30650 7899 30706
rect 7969 30650 8025 30706
rect 7843 30568 7899 30624
rect 7969 30568 8025 30624
rect 7843 30486 7899 30542
rect 7969 30486 8025 30542
rect 7843 30404 7899 30460
rect 7969 30404 8025 30460
rect 7843 30322 7899 30378
rect 7969 30322 8025 30378
rect 7843 30240 7899 30296
rect 7969 30240 8025 30296
rect 7843 30158 7899 30214
rect 7969 30158 8025 30214
rect 7843 30076 7899 30132
rect 7969 30076 8025 30132
rect 7843 29994 7899 30050
rect 7969 29994 8025 30050
rect 7843 29912 7899 29968
rect 7969 29912 8025 29968
rect 7843 29830 7899 29886
rect 7969 29830 8025 29886
rect 7843 29748 7899 29804
rect 7969 29748 8025 29804
rect 7843 29666 7899 29722
rect 7969 29666 8025 29722
rect 7843 29584 7899 29640
rect 7969 29584 8025 29640
rect 7843 29502 7899 29558
rect 7969 29502 8025 29558
rect 7843 29420 7899 29476
rect 7969 29420 8025 29476
rect 8339 31962 8395 32018
rect 8465 31962 8521 32018
rect 8339 31880 8395 31936
rect 8465 31880 8521 31936
rect 8339 31798 8395 31854
rect 8465 31798 8521 31854
rect 8339 31716 8395 31772
rect 8465 31716 8521 31772
rect 8339 31634 8395 31690
rect 8465 31634 8521 31690
rect 8339 31552 8395 31608
rect 8465 31552 8521 31608
rect 8339 31470 8395 31526
rect 8465 31470 8521 31526
rect 8339 31388 8395 31444
rect 8465 31388 8521 31444
rect 8339 31306 8395 31362
rect 8465 31306 8521 31362
rect 8339 31224 8395 31280
rect 8465 31224 8521 31280
rect 8339 31142 8395 31198
rect 8465 31142 8521 31198
rect 8339 31060 8395 31116
rect 8465 31060 8521 31116
rect 8339 30978 8395 31034
rect 8465 30978 8521 31034
rect 8339 30896 8395 30952
rect 8465 30896 8521 30952
rect 8339 30814 8395 30870
rect 8465 30814 8521 30870
rect 8339 30732 8395 30788
rect 8465 30732 8521 30788
rect 8339 30650 8395 30706
rect 8465 30650 8521 30706
rect 8339 30568 8395 30624
rect 8465 30568 8521 30624
rect 8339 30486 8395 30542
rect 8465 30486 8521 30542
rect 8339 30404 8395 30460
rect 8465 30404 8521 30460
rect 8339 30322 8395 30378
rect 8465 30322 8521 30378
rect 8339 30240 8395 30296
rect 8465 30240 8521 30296
rect 8339 30158 8395 30214
rect 8465 30158 8521 30214
rect 8339 30076 8395 30132
rect 8465 30076 8521 30132
rect 8339 29994 8395 30050
rect 8465 29994 8521 30050
rect 8339 29912 8395 29968
rect 8465 29912 8521 29968
rect 8339 29830 8395 29886
rect 8465 29830 8521 29886
rect 8339 29748 8395 29804
rect 8465 29748 8521 29804
rect 8339 29666 8395 29722
rect 8465 29666 8521 29722
rect 8339 29584 8395 29640
rect 8465 29584 8521 29640
rect 8339 29502 8395 29558
rect 8465 29502 8521 29558
rect 8339 29420 8395 29476
rect 8465 29420 8521 29476
rect 8835 31962 8891 32018
rect 8961 31962 9017 32018
rect 8835 31880 8891 31936
rect 8961 31880 9017 31936
rect 8835 31798 8891 31854
rect 8961 31798 9017 31854
rect 8835 31716 8891 31772
rect 8961 31716 9017 31772
rect 8835 31634 8891 31690
rect 8961 31634 9017 31690
rect 8835 31552 8891 31608
rect 8961 31552 9017 31608
rect 8835 31470 8891 31526
rect 8961 31470 9017 31526
rect 8835 31388 8891 31444
rect 8961 31388 9017 31444
rect 8835 31306 8891 31362
rect 8961 31306 9017 31362
rect 8835 31224 8891 31280
rect 8961 31224 9017 31280
rect 8835 31142 8891 31198
rect 8961 31142 9017 31198
rect 8835 31060 8891 31116
rect 8961 31060 9017 31116
rect 8835 30978 8891 31034
rect 8961 30978 9017 31034
rect 8835 30896 8891 30952
rect 8961 30896 9017 30952
rect 8835 30814 8891 30870
rect 8961 30814 9017 30870
rect 8835 30732 8891 30788
rect 8961 30732 9017 30788
rect 8835 30650 8891 30706
rect 8961 30650 9017 30706
rect 8835 30568 8891 30624
rect 8961 30568 9017 30624
rect 8835 30486 8891 30542
rect 8961 30486 9017 30542
rect 8835 30404 8891 30460
rect 8961 30404 9017 30460
rect 8835 30322 8891 30378
rect 8961 30322 9017 30378
rect 8835 30240 8891 30296
rect 8961 30240 9017 30296
rect 8835 30158 8891 30214
rect 8961 30158 9017 30214
rect 8835 30076 8891 30132
rect 8961 30076 9017 30132
rect 8835 29994 8891 30050
rect 8961 29994 9017 30050
rect 8835 29912 8891 29968
rect 8961 29912 9017 29968
rect 8835 29830 8891 29886
rect 8961 29830 9017 29886
rect 8835 29748 8891 29804
rect 8961 29748 9017 29804
rect 8835 29666 8891 29722
rect 8961 29666 9017 29722
rect 8835 29584 8891 29640
rect 8961 29584 9017 29640
rect 8835 29502 8891 29558
rect 8961 29502 9017 29558
rect 8835 29420 8891 29476
rect 8961 29420 9017 29476
rect 9331 31962 9387 32018
rect 9457 31962 9513 32018
rect 9331 31880 9387 31936
rect 9457 31880 9513 31936
rect 9331 31798 9387 31854
rect 9457 31798 9513 31854
rect 9331 31716 9387 31772
rect 9457 31716 9513 31772
rect 9331 31634 9387 31690
rect 9457 31634 9513 31690
rect 9331 31552 9387 31608
rect 9457 31552 9513 31608
rect 9331 31470 9387 31526
rect 9457 31470 9513 31526
rect 9331 31388 9387 31444
rect 9457 31388 9513 31444
rect 9331 31306 9387 31362
rect 9457 31306 9513 31362
rect 9331 31224 9387 31280
rect 9457 31224 9513 31280
rect 9331 31142 9387 31198
rect 9457 31142 9513 31198
rect 9331 31060 9387 31116
rect 9457 31060 9513 31116
rect 9331 30978 9387 31034
rect 9457 30978 9513 31034
rect 9331 30896 9387 30952
rect 9457 30896 9513 30952
rect 9331 30814 9387 30870
rect 9457 30814 9513 30870
rect 9331 30732 9387 30788
rect 9457 30732 9513 30788
rect 9331 30650 9387 30706
rect 9457 30650 9513 30706
rect 9331 30568 9387 30624
rect 9457 30568 9513 30624
rect 9331 30486 9387 30542
rect 9457 30486 9513 30542
rect 9331 30404 9387 30460
rect 9457 30404 9513 30460
rect 9331 30322 9387 30378
rect 9457 30322 9513 30378
rect 9331 30240 9387 30296
rect 9457 30240 9513 30296
rect 9331 30158 9387 30214
rect 9457 30158 9513 30214
rect 9331 30076 9387 30132
rect 9457 30076 9513 30132
rect 9331 29994 9387 30050
rect 9457 29994 9513 30050
rect 9331 29912 9387 29968
rect 9457 29912 9513 29968
rect 9331 29830 9387 29886
rect 9457 29830 9513 29886
rect 9331 29748 9387 29804
rect 9457 29748 9513 29804
rect 9331 29666 9387 29722
rect 9457 29666 9513 29722
rect 9331 29584 9387 29640
rect 9457 29584 9513 29640
rect 9331 29502 9387 29558
rect 9457 29502 9513 29558
rect 9331 29420 9387 29476
rect 9457 29420 9513 29476
rect 9827 31962 9883 32018
rect 9953 31962 10009 32018
rect 9827 31880 9883 31936
rect 9953 31880 10009 31936
rect 9827 31798 9883 31854
rect 9953 31798 10009 31854
rect 9827 31716 9883 31772
rect 9953 31716 10009 31772
rect 9827 31634 9883 31690
rect 9953 31634 10009 31690
rect 9827 31552 9883 31608
rect 9953 31552 10009 31608
rect 9827 31470 9883 31526
rect 9953 31470 10009 31526
rect 9827 31388 9883 31444
rect 9953 31388 10009 31444
rect 9827 31306 9883 31362
rect 9953 31306 10009 31362
rect 9827 31224 9883 31280
rect 9953 31224 10009 31280
rect 9827 31142 9883 31198
rect 9953 31142 10009 31198
rect 9827 31060 9883 31116
rect 9953 31060 10009 31116
rect 9827 30978 9883 31034
rect 9953 30978 10009 31034
rect 9827 30896 9883 30952
rect 9953 30896 10009 30952
rect 9827 30814 9883 30870
rect 9953 30814 10009 30870
rect 9827 30732 9883 30788
rect 9953 30732 10009 30788
rect 9827 30650 9883 30706
rect 9953 30650 10009 30706
rect 9827 30568 9883 30624
rect 9953 30568 10009 30624
rect 9827 30486 9883 30542
rect 9953 30486 10009 30542
rect 9827 30404 9883 30460
rect 9953 30404 10009 30460
rect 9827 30322 9883 30378
rect 9953 30322 10009 30378
rect 9827 30240 9883 30296
rect 9953 30240 10009 30296
rect 9827 30158 9883 30214
rect 9953 30158 10009 30214
rect 9827 30076 9883 30132
rect 9953 30076 10009 30132
rect 9827 29994 9883 30050
rect 9953 29994 10009 30050
rect 9827 29912 9883 29968
rect 9953 29912 10009 29968
rect 9827 29830 9883 29886
rect 9953 29830 10009 29886
rect 9827 29748 9883 29804
rect 9953 29748 10009 29804
rect 9827 29666 9883 29722
rect 9953 29666 10009 29722
rect 9827 29584 9883 29640
rect 9953 29584 10009 29640
rect 9827 29502 9883 29558
rect 9953 29502 10009 29558
rect 9827 29420 9883 29476
rect 9953 29420 10009 29476
rect 10323 31962 10379 32018
rect 10449 31962 10505 32018
rect 10323 31880 10379 31936
rect 10449 31880 10505 31936
rect 10323 31798 10379 31854
rect 10449 31798 10505 31854
rect 10323 31716 10379 31772
rect 10449 31716 10505 31772
rect 10323 31634 10379 31690
rect 10449 31634 10505 31690
rect 10323 31552 10379 31608
rect 10449 31552 10505 31608
rect 10323 31470 10379 31526
rect 10449 31470 10505 31526
rect 10323 31388 10379 31444
rect 10449 31388 10505 31444
rect 10323 31306 10379 31362
rect 10449 31306 10505 31362
rect 10323 31224 10379 31280
rect 10449 31224 10505 31280
rect 10323 31142 10379 31198
rect 10449 31142 10505 31198
rect 10323 31060 10379 31116
rect 10449 31060 10505 31116
rect 10323 30978 10379 31034
rect 10449 30978 10505 31034
rect 10323 30896 10379 30952
rect 10449 30896 10505 30952
rect 10323 30814 10379 30870
rect 10449 30814 10505 30870
rect 10323 30732 10379 30788
rect 10449 30732 10505 30788
rect 10323 30650 10379 30706
rect 10449 30650 10505 30706
rect 10323 30568 10379 30624
rect 10449 30568 10505 30624
rect 10323 30486 10379 30542
rect 10449 30486 10505 30542
rect 10323 30404 10379 30460
rect 10449 30404 10505 30460
rect 10323 30322 10379 30378
rect 10449 30322 10505 30378
rect 10323 30240 10379 30296
rect 10449 30240 10505 30296
rect 10323 30158 10379 30214
rect 10449 30158 10505 30214
rect 10323 30076 10379 30132
rect 10449 30076 10505 30132
rect 10323 29994 10379 30050
rect 10449 29994 10505 30050
rect 10323 29912 10379 29968
rect 10449 29912 10505 29968
rect 10323 29830 10379 29886
rect 10449 29830 10505 29886
rect 10323 29748 10379 29804
rect 10449 29748 10505 29804
rect 10323 29666 10379 29722
rect 10449 29666 10505 29722
rect 10323 29584 10379 29640
rect 10449 29584 10505 29640
rect 10323 29502 10379 29558
rect 10449 29502 10505 29558
rect 10323 29420 10379 29476
rect 10449 29420 10505 29476
rect 10819 31962 10875 32018
rect 10945 31962 11001 32018
rect 10819 31880 10875 31936
rect 10945 31880 11001 31936
rect 10819 31798 10875 31854
rect 10945 31798 11001 31854
rect 10819 31716 10875 31772
rect 10945 31716 11001 31772
rect 10819 31634 10875 31690
rect 10945 31634 11001 31690
rect 10819 31552 10875 31608
rect 10945 31552 11001 31608
rect 10819 31470 10875 31526
rect 10945 31470 11001 31526
rect 10819 31388 10875 31444
rect 10945 31388 11001 31444
rect 10819 31306 10875 31362
rect 10945 31306 11001 31362
rect 10819 31224 10875 31280
rect 10945 31224 11001 31280
rect 10819 31142 10875 31198
rect 10945 31142 11001 31198
rect 10819 31060 10875 31116
rect 10945 31060 11001 31116
rect 10819 30978 10875 31034
rect 10945 30978 11001 31034
rect 10819 30896 10875 30952
rect 10945 30896 11001 30952
rect 10819 30814 10875 30870
rect 10945 30814 11001 30870
rect 10819 30732 10875 30788
rect 10945 30732 11001 30788
rect 10819 30650 10875 30706
rect 10945 30650 11001 30706
rect 10819 30568 10875 30624
rect 10945 30568 11001 30624
rect 10819 30486 10875 30542
rect 10945 30486 11001 30542
rect 10819 30404 10875 30460
rect 10945 30404 11001 30460
rect 10819 30322 10875 30378
rect 10945 30322 11001 30378
rect 10819 30240 10875 30296
rect 10945 30240 11001 30296
rect 10819 30158 10875 30214
rect 10945 30158 11001 30214
rect 10819 30076 10875 30132
rect 10945 30076 11001 30132
rect 10819 29994 10875 30050
rect 10945 29994 11001 30050
rect 10819 29912 10875 29968
rect 10945 29912 11001 29968
rect 10819 29830 10875 29886
rect 10945 29830 11001 29886
rect 10819 29748 10875 29804
rect 10945 29748 11001 29804
rect 10819 29666 10875 29722
rect 10945 29666 11001 29722
rect 10819 29584 10875 29640
rect 10945 29584 11001 29640
rect 10819 29502 10875 29558
rect 10945 29502 11001 29558
rect 10819 29420 10875 29476
rect 10945 29420 11001 29476
rect 11315 31962 11371 32018
rect 11441 31962 11497 32018
rect 11315 31880 11371 31936
rect 11441 31880 11497 31936
rect 11315 31798 11371 31854
rect 11441 31798 11497 31854
rect 11315 31716 11371 31772
rect 11441 31716 11497 31772
rect 11315 31634 11371 31690
rect 11441 31634 11497 31690
rect 11315 31552 11371 31608
rect 11441 31552 11497 31608
rect 11315 31470 11371 31526
rect 11441 31470 11497 31526
rect 11315 31388 11371 31444
rect 11441 31388 11497 31444
rect 11315 31306 11371 31362
rect 11441 31306 11497 31362
rect 11315 31224 11371 31280
rect 11441 31224 11497 31280
rect 11315 31142 11371 31198
rect 11441 31142 11497 31198
rect 11315 31060 11371 31116
rect 11441 31060 11497 31116
rect 11315 30978 11371 31034
rect 11441 30978 11497 31034
rect 11315 30896 11371 30952
rect 11441 30896 11497 30952
rect 11315 30814 11371 30870
rect 11441 30814 11497 30870
rect 11315 30732 11371 30788
rect 11441 30732 11497 30788
rect 11315 30650 11371 30706
rect 11441 30650 11497 30706
rect 11315 30568 11371 30624
rect 11441 30568 11497 30624
rect 11315 30486 11371 30542
rect 11441 30486 11497 30542
rect 11315 30404 11371 30460
rect 11441 30404 11497 30460
rect 11315 30322 11371 30378
rect 11441 30322 11497 30378
rect 11315 30240 11371 30296
rect 11441 30240 11497 30296
rect 11315 30158 11371 30214
rect 11441 30158 11497 30214
rect 11315 30076 11371 30132
rect 11441 30076 11497 30132
rect 11315 29994 11371 30050
rect 11441 29994 11497 30050
rect 11315 29912 11371 29968
rect 11441 29912 11497 29968
rect 11315 29830 11371 29886
rect 11441 29830 11497 29886
rect 11315 29748 11371 29804
rect 11441 29748 11497 29804
rect 11315 29666 11371 29722
rect 11441 29666 11497 29722
rect 11315 29584 11371 29640
rect 11441 29584 11497 29640
rect 11315 29502 11371 29558
rect 11441 29502 11497 29558
rect 11315 29420 11371 29476
rect 11441 29420 11497 29476
rect 11811 31962 11867 32018
rect 11937 31962 11993 32018
rect 11811 31880 11867 31936
rect 11937 31880 11993 31936
rect 11811 31798 11867 31854
rect 11937 31798 11993 31854
rect 11811 31716 11867 31772
rect 11937 31716 11993 31772
rect 11811 31634 11867 31690
rect 11937 31634 11993 31690
rect 11811 31552 11867 31608
rect 11937 31552 11993 31608
rect 11811 31470 11867 31526
rect 11937 31470 11993 31526
rect 11811 31388 11867 31444
rect 11937 31388 11993 31444
rect 11811 31306 11867 31362
rect 11937 31306 11993 31362
rect 11811 31224 11867 31280
rect 11937 31224 11993 31280
rect 11811 31142 11867 31198
rect 11937 31142 11993 31198
rect 11811 31060 11867 31116
rect 11937 31060 11993 31116
rect 11811 30978 11867 31034
rect 11937 30978 11993 31034
rect 11811 30896 11867 30952
rect 11937 30896 11993 30952
rect 11811 30814 11867 30870
rect 11937 30814 11993 30870
rect 11811 30732 11867 30788
rect 11937 30732 11993 30788
rect 11811 30650 11867 30706
rect 11937 30650 11993 30706
rect 11811 30568 11867 30624
rect 11937 30568 11993 30624
rect 11811 30486 11867 30542
rect 11937 30486 11993 30542
rect 11811 30404 11867 30460
rect 11937 30404 11993 30460
rect 11811 30322 11867 30378
rect 11937 30322 11993 30378
rect 11811 30240 11867 30296
rect 11937 30240 11993 30296
rect 11811 30158 11867 30214
rect 11937 30158 11993 30214
rect 11811 30076 11867 30132
rect 11937 30076 11993 30132
rect 11811 29994 11867 30050
rect 11937 29994 11993 30050
rect 11811 29912 11867 29968
rect 11937 29912 11993 29968
rect 11811 29830 11867 29886
rect 11937 29830 11993 29886
rect 11811 29748 11867 29804
rect 11937 29748 11993 29804
rect 11811 29666 11867 29722
rect 11937 29666 11993 29722
rect 11811 29584 11867 29640
rect 11937 29584 11993 29640
rect 11811 29502 11867 29558
rect 11937 29502 11993 29558
rect 11811 29420 11867 29476
rect 11937 29420 11993 29476
rect 12307 31962 12363 32018
rect 12433 31962 12489 32018
rect 12307 31880 12363 31936
rect 12433 31880 12489 31936
rect 12307 31798 12363 31854
rect 12433 31798 12489 31854
rect 12307 31716 12363 31772
rect 12433 31716 12489 31772
rect 12307 31634 12363 31690
rect 12433 31634 12489 31690
rect 12307 31552 12363 31608
rect 12433 31552 12489 31608
rect 12307 31470 12363 31526
rect 12433 31470 12489 31526
rect 12307 31388 12363 31444
rect 12433 31388 12489 31444
rect 12307 31306 12363 31362
rect 12433 31306 12489 31362
rect 12307 31224 12363 31280
rect 12433 31224 12489 31280
rect 12307 31142 12363 31198
rect 12433 31142 12489 31198
rect 12307 31060 12363 31116
rect 12433 31060 12489 31116
rect 12307 30978 12363 31034
rect 12433 30978 12489 31034
rect 12307 30896 12363 30952
rect 12433 30896 12489 30952
rect 12307 30814 12363 30870
rect 12433 30814 12489 30870
rect 12307 30732 12363 30788
rect 12433 30732 12489 30788
rect 12307 30650 12363 30706
rect 12433 30650 12489 30706
rect 12307 30568 12363 30624
rect 12433 30568 12489 30624
rect 12307 30486 12363 30542
rect 12433 30486 12489 30542
rect 12307 30404 12363 30460
rect 12433 30404 12489 30460
rect 12307 30322 12363 30378
rect 12433 30322 12489 30378
rect 12307 30240 12363 30296
rect 12433 30240 12489 30296
rect 12307 30158 12363 30214
rect 12433 30158 12489 30214
rect 12307 30076 12363 30132
rect 12433 30076 12489 30132
rect 12307 29994 12363 30050
rect 12433 29994 12489 30050
rect 12307 29912 12363 29968
rect 12433 29912 12489 29968
rect 12307 29830 12363 29886
rect 12433 29830 12489 29886
rect 12307 29748 12363 29804
rect 12433 29748 12489 29804
rect 12307 29666 12363 29722
rect 12433 29666 12489 29722
rect 12307 29584 12363 29640
rect 12433 29584 12489 29640
rect 12307 29502 12363 29558
rect 12433 29502 12489 29558
rect 12307 29420 12363 29476
rect 12433 29420 12489 29476
rect 12803 31962 12859 32018
rect 12929 31962 12985 32018
rect 12803 31880 12859 31936
rect 12929 31880 12985 31936
rect 12803 31798 12859 31854
rect 12929 31798 12985 31854
rect 12803 31716 12859 31772
rect 12929 31716 12985 31772
rect 12803 31634 12859 31690
rect 12929 31634 12985 31690
rect 12803 31552 12859 31608
rect 12929 31552 12985 31608
rect 12803 31470 12859 31526
rect 12929 31470 12985 31526
rect 12803 31388 12859 31444
rect 12929 31388 12985 31444
rect 12803 31306 12859 31362
rect 12929 31306 12985 31362
rect 12803 31224 12859 31280
rect 12929 31224 12985 31280
rect 12803 31142 12859 31198
rect 12929 31142 12985 31198
rect 12803 31060 12859 31116
rect 12929 31060 12985 31116
rect 12803 30978 12859 31034
rect 12929 30978 12985 31034
rect 12803 30896 12859 30952
rect 12929 30896 12985 30952
rect 12803 30814 12859 30870
rect 12929 30814 12985 30870
rect 12803 30732 12859 30788
rect 12929 30732 12985 30788
rect 12803 30650 12859 30706
rect 12929 30650 12985 30706
rect 12803 30568 12859 30624
rect 12929 30568 12985 30624
rect 12803 30486 12859 30542
rect 12929 30486 12985 30542
rect 12803 30404 12859 30460
rect 12929 30404 12985 30460
rect 12803 30322 12859 30378
rect 12929 30322 12985 30378
rect 12803 30240 12859 30296
rect 12929 30240 12985 30296
rect 12803 30158 12859 30214
rect 12929 30158 12985 30214
rect 12803 30076 12859 30132
rect 12929 30076 12985 30132
rect 12803 29994 12859 30050
rect 12929 29994 12985 30050
rect 12803 29912 12859 29968
rect 12929 29912 12985 29968
rect 12803 29830 12859 29886
rect 12929 29830 12985 29886
rect 12803 29748 12859 29804
rect 12929 29748 12985 29804
rect 12803 29666 12859 29722
rect 12929 29666 12985 29722
rect 12803 29584 12859 29640
rect 12929 29584 12985 29640
rect 12803 29502 12859 29558
rect 12929 29502 12985 29558
rect 12803 29420 12859 29476
rect 12929 29420 12985 29476
rect 13299 31962 13355 32018
rect 13425 31962 13481 32018
rect 13299 31880 13355 31936
rect 13425 31880 13481 31936
rect 13299 31798 13355 31854
rect 13425 31798 13481 31854
rect 13299 31716 13355 31772
rect 13425 31716 13481 31772
rect 13299 31634 13355 31690
rect 13425 31634 13481 31690
rect 13299 31552 13355 31608
rect 13425 31552 13481 31608
rect 13299 31470 13355 31526
rect 13425 31470 13481 31526
rect 13299 31388 13355 31444
rect 13425 31388 13481 31444
rect 13299 31306 13355 31362
rect 13425 31306 13481 31362
rect 13299 31224 13355 31280
rect 13425 31224 13481 31280
rect 13299 31142 13355 31198
rect 13425 31142 13481 31198
rect 13299 31060 13355 31116
rect 13425 31060 13481 31116
rect 13299 30978 13355 31034
rect 13425 30978 13481 31034
rect 13299 30896 13355 30952
rect 13425 30896 13481 30952
rect 13299 30814 13355 30870
rect 13425 30814 13481 30870
rect 13299 30732 13355 30788
rect 13425 30732 13481 30788
rect 13299 30650 13355 30706
rect 13425 30650 13481 30706
rect 13299 30568 13355 30624
rect 13425 30568 13481 30624
rect 13299 30486 13355 30542
rect 13425 30486 13481 30542
rect 13299 30404 13355 30460
rect 13425 30404 13481 30460
rect 13299 30322 13355 30378
rect 13425 30322 13481 30378
rect 13299 30240 13355 30296
rect 13425 30240 13481 30296
rect 13299 30158 13355 30214
rect 13425 30158 13481 30214
rect 13299 30076 13355 30132
rect 13425 30076 13481 30132
rect 13299 29994 13355 30050
rect 13425 29994 13481 30050
rect 13299 29912 13355 29968
rect 13425 29912 13481 29968
rect 13299 29830 13355 29886
rect 13425 29830 13481 29886
rect 13299 29748 13355 29804
rect 13425 29748 13481 29804
rect 13299 29666 13355 29722
rect 13425 29666 13481 29722
rect 13299 29584 13355 29640
rect 13425 29584 13481 29640
rect 13299 29502 13355 29558
rect 13425 29502 13481 29558
rect 13299 29420 13355 29476
rect 13425 29420 13481 29476
rect 13795 31962 13851 32018
rect 13921 31962 13977 32018
rect 13795 31880 13851 31936
rect 13921 31880 13977 31936
rect 13795 31798 13851 31854
rect 13921 31798 13977 31854
rect 13795 31716 13851 31772
rect 13921 31716 13977 31772
rect 13795 31634 13851 31690
rect 13921 31634 13977 31690
rect 13795 31552 13851 31608
rect 13921 31552 13977 31608
rect 13795 31470 13851 31526
rect 13921 31470 13977 31526
rect 13795 31388 13851 31444
rect 13921 31388 13977 31444
rect 13795 31306 13851 31362
rect 13921 31306 13977 31362
rect 13795 31224 13851 31280
rect 13921 31224 13977 31280
rect 13795 31142 13851 31198
rect 13921 31142 13977 31198
rect 13795 31060 13851 31116
rect 13921 31060 13977 31116
rect 13795 30978 13851 31034
rect 13921 30978 13977 31034
rect 13795 30896 13851 30952
rect 13921 30896 13977 30952
rect 13795 30814 13851 30870
rect 13921 30814 13977 30870
rect 13795 30732 13851 30788
rect 13921 30732 13977 30788
rect 13795 30650 13851 30706
rect 13921 30650 13977 30706
rect 13795 30568 13851 30624
rect 13921 30568 13977 30624
rect 13795 30486 13851 30542
rect 13921 30486 13977 30542
rect 13795 30404 13851 30460
rect 13921 30404 13977 30460
rect 13795 30322 13851 30378
rect 13921 30322 13977 30378
rect 13795 30240 13851 30296
rect 13921 30240 13977 30296
rect 13795 30158 13851 30214
rect 13921 30158 13977 30214
rect 13795 30076 13851 30132
rect 13921 30076 13977 30132
rect 13795 29994 13851 30050
rect 13921 29994 13977 30050
rect 13795 29912 13851 29968
rect 13921 29912 13977 29968
rect 13795 29830 13851 29886
rect 13921 29830 13977 29886
rect 13795 29748 13851 29804
rect 13921 29748 13977 29804
rect 13795 29666 13851 29722
rect 13921 29666 13977 29722
rect 13795 29584 13851 29640
rect 13921 29584 13977 29640
rect 13795 29502 13851 29558
rect 13921 29502 13977 29558
rect 13795 29420 13851 29476
rect 13921 29420 13977 29476
rect 14259 31985 14315 32041
rect 14347 31985 14403 32041
rect 14435 31985 14491 32041
rect 14523 31985 14579 32041
rect 14611 31985 14667 32041
rect 14259 31905 14315 31961
rect 14347 31905 14403 31961
rect 14435 31905 14491 31961
rect 14523 31905 14579 31961
rect 14611 31905 14667 31961
rect 14259 31825 14315 31881
rect 14347 31825 14403 31881
rect 14435 31825 14491 31881
rect 14523 31825 14579 31881
rect 14611 31825 14667 31881
rect 14259 31745 14315 31801
rect 14347 31745 14403 31801
rect 14435 31745 14491 31801
rect 14523 31745 14579 31801
rect 14611 31745 14667 31801
rect 14259 31665 14315 31721
rect 14347 31665 14403 31721
rect 14435 31665 14491 31721
rect 14523 31665 14579 31721
rect 14611 31665 14667 31721
rect 14259 31585 14315 31641
rect 14347 31585 14403 31641
rect 14435 31585 14491 31641
rect 14523 31585 14579 31641
rect 14611 31585 14667 31641
rect 14259 31505 14315 31561
rect 14347 31505 14403 31561
rect 14435 31505 14491 31561
rect 14523 31505 14579 31561
rect 14611 31505 14667 31561
rect 14259 31425 14315 31481
rect 14347 31425 14403 31481
rect 14435 31425 14491 31481
rect 14523 31425 14579 31481
rect 14611 31425 14667 31481
rect 14259 31344 14315 31400
rect 14347 31344 14403 31400
rect 14435 31344 14491 31400
rect 14523 31344 14579 31400
rect 14611 31344 14667 31400
rect 14259 31263 14315 31319
rect 14347 31263 14403 31319
rect 14435 31263 14491 31319
rect 14523 31263 14579 31319
rect 14611 31263 14667 31319
rect 14259 31182 14315 31238
rect 14347 31182 14403 31238
rect 14435 31182 14491 31238
rect 14523 31182 14579 31238
rect 14611 31182 14667 31238
rect 14259 31101 14315 31157
rect 14347 31101 14403 31157
rect 14435 31101 14491 31157
rect 14523 31101 14579 31157
rect 14611 31101 14667 31157
rect 14259 31020 14315 31076
rect 14347 31020 14403 31076
rect 14435 31020 14491 31076
rect 14523 31020 14579 31076
rect 14611 31020 14667 31076
rect 14259 30939 14315 30995
rect 14347 30939 14403 30995
rect 14435 30939 14491 30995
rect 14523 30939 14579 30995
rect 14611 30939 14667 30995
rect 14259 30858 14315 30914
rect 14347 30858 14403 30914
rect 14435 30858 14491 30914
rect 14523 30858 14579 30914
rect 14611 30858 14667 30914
rect 14259 30777 14315 30833
rect 14347 30777 14403 30833
rect 14435 30777 14491 30833
rect 14523 30777 14579 30833
rect 14611 30777 14667 30833
rect 14259 30696 14315 30752
rect 14347 30696 14403 30752
rect 14435 30696 14491 30752
rect 14523 30696 14579 30752
rect 14611 30696 14667 30752
rect 14259 30615 14315 30671
rect 14347 30615 14403 30671
rect 14435 30615 14491 30671
rect 14523 30615 14579 30671
rect 14611 30615 14667 30671
rect 14259 30534 14315 30590
rect 14347 30534 14403 30590
rect 14435 30534 14491 30590
rect 14523 30534 14579 30590
rect 14611 30534 14667 30590
rect 14259 30453 14315 30509
rect 14347 30453 14403 30509
rect 14435 30453 14491 30509
rect 14523 30453 14579 30509
rect 14611 30453 14667 30509
rect 14259 30372 14315 30428
rect 14347 30372 14403 30428
rect 14435 30372 14491 30428
rect 14523 30372 14579 30428
rect 14611 30372 14667 30428
rect 14259 30291 14315 30347
rect 14347 30291 14403 30347
rect 14435 30291 14491 30347
rect 14523 30291 14579 30347
rect 14611 30291 14667 30347
rect 14259 30210 14315 30266
rect 14347 30210 14403 30266
rect 14435 30210 14491 30266
rect 14523 30210 14579 30266
rect 14611 30210 14667 30266
rect 14259 30129 14315 30185
rect 14347 30129 14403 30185
rect 14435 30129 14491 30185
rect 14523 30129 14579 30185
rect 14611 30129 14667 30185
rect 14259 30048 14315 30104
rect 14347 30048 14403 30104
rect 14435 30048 14491 30104
rect 14523 30048 14579 30104
rect 14611 30048 14667 30104
rect 14259 29967 14315 30023
rect 14347 29967 14403 30023
rect 14435 29967 14491 30023
rect 14523 29967 14579 30023
rect 14611 29967 14667 30023
rect 14259 29886 14315 29942
rect 14347 29886 14403 29942
rect 14435 29886 14491 29942
rect 14523 29886 14579 29942
rect 14611 29886 14667 29942
rect 14259 29805 14315 29861
rect 14347 29805 14403 29861
rect 14435 29805 14491 29861
rect 14523 29805 14579 29861
rect 14611 29805 14667 29861
rect 14259 29724 14315 29780
rect 14347 29724 14403 29780
rect 14435 29724 14491 29780
rect 14523 29724 14579 29780
rect 14611 29724 14667 29780
rect 14259 29643 14315 29699
rect 14347 29643 14403 29699
rect 14435 29643 14491 29699
rect 14523 29643 14579 29699
rect 14611 29643 14667 29699
rect 14259 29562 14315 29618
rect 14347 29562 14403 29618
rect 14435 29562 14491 29618
rect 14523 29562 14579 29618
rect 14611 29562 14667 29618
rect 14259 29481 14315 29537
rect 14347 29481 14403 29537
rect 14435 29481 14491 29537
rect 14523 29481 14579 29537
rect 14611 29481 14667 29537
rect 14259 29400 14315 29456
rect 14347 29400 14403 29456
rect 14435 29400 14491 29456
rect 14523 29400 14579 29456
rect 14611 29400 14667 29456
rect 14259 29319 14315 29375
rect 14347 29319 14403 29375
rect 14435 29319 14491 29375
rect 14523 29319 14579 29375
rect 14611 29319 14667 29375
rect 14259 29238 14315 29294
rect 14347 29238 14403 29294
rect 14435 29238 14491 29294
rect 14523 29238 14579 29294
rect 14611 29238 14667 29294
rect 14259 29157 14315 29213
rect 14347 29157 14403 29213
rect 14435 29157 14491 29213
rect 14523 29157 14579 29213
rect 14611 29157 14667 29213
rect 14259 29076 14315 29132
rect 14347 29076 14403 29132
rect 14435 29076 14491 29132
rect 14523 29076 14579 29132
rect 14611 29076 14667 29132
rect 579 28580 581 28596
rect 581 28580 633 28596
rect 633 28580 635 28596
rect 677 28580 702 28596
rect 702 28580 719 28596
rect 719 28580 733 28596
rect 775 28580 788 28596
rect 788 28580 831 28596
rect 579 28558 635 28580
rect 677 28558 733 28580
rect 775 28558 831 28580
rect 579 28540 581 28558
rect 581 28540 633 28558
rect 633 28540 635 28558
rect 677 28540 702 28558
rect 702 28540 719 28558
rect 719 28540 733 28558
rect 775 28540 788 28558
rect 788 28540 831 28558
rect 579 28506 581 28515
rect 581 28506 633 28515
rect 633 28506 635 28515
rect 677 28506 702 28515
rect 702 28506 719 28515
rect 719 28506 733 28515
rect 775 28506 788 28515
rect 788 28506 831 28515
rect 579 28484 635 28506
rect 677 28484 733 28506
rect 775 28484 831 28506
rect 579 28459 581 28484
rect 581 28459 633 28484
rect 633 28459 635 28484
rect 677 28459 702 28484
rect 702 28459 719 28484
rect 719 28459 733 28484
rect 775 28459 788 28484
rect 788 28459 831 28484
rect 579 28432 581 28434
rect 581 28432 633 28434
rect 633 28432 635 28434
rect 677 28432 702 28434
rect 702 28432 719 28434
rect 719 28432 733 28434
rect 775 28432 788 28434
rect 788 28432 831 28434
rect 579 28378 635 28432
rect 677 28378 733 28432
rect 775 28378 831 28432
rect 579 28297 635 28353
rect 677 28297 733 28353
rect 775 28297 831 28353
rect 579 28216 635 28272
rect 677 28216 733 28272
rect 775 28216 831 28272
rect 579 28135 635 28191
rect 677 28135 733 28191
rect 775 28135 831 28191
rect 3494 28581 3530 28620
rect 3530 28581 3546 28620
rect 3546 28581 3550 28620
rect 4485 28581 4490 28620
rect 4490 28581 4541 28620
rect 3494 28564 3550 28581
rect 4485 28564 4541 28581
rect 3494 28433 3530 28451
rect 3530 28433 3546 28451
rect 3546 28433 3550 28451
rect 4485 28433 4490 28451
rect 4490 28433 4541 28451
rect 3494 28395 3550 28433
rect 4485 28395 4541 28433
rect 3494 28226 3550 28282
rect 4485 28226 4541 28282
rect 579 28054 635 28110
rect 677 28054 733 28110
rect 775 28054 831 28110
rect 579 27973 635 28029
rect 677 27973 733 28029
rect 775 27973 831 28029
rect 579 27892 635 27948
rect 677 27892 733 27948
rect 775 27892 831 27948
rect 579 27811 635 27867
rect 677 27811 733 27867
rect 775 27811 831 27867
rect 579 27730 635 27786
rect 677 27730 733 27786
rect 775 27730 831 27786
rect 579 27649 635 27705
rect 677 27649 733 27705
rect 775 27649 831 27705
rect 579 27568 635 27624
rect 677 27568 733 27624
rect 775 27568 831 27624
rect 579 27487 635 27543
rect 677 27487 733 27543
rect 775 27487 831 27543
rect 579 27406 635 27462
rect 677 27406 733 27462
rect 775 27406 831 27462
rect 579 27325 635 27381
rect 677 27325 733 27381
rect 775 27325 831 27381
rect 579 27244 635 27300
rect 677 27244 733 27300
rect 775 27244 831 27300
rect 579 27163 635 27219
rect 677 27163 733 27219
rect 775 27163 831 27219
rect 579 27082 635 27138
rect 677 27082 733 27138
rect 775 27082 831 27138
rect 579 27001 635 27057
rect 677 27001 733 27057
rect 775 27001 831 27057
rect 579 26920 635 26976
rect 677 26920 733 26976
rect 775 26920 831 26976
rect 579 26838 635 26894
rect 677 26838 733 26894
rect 775 26838 831 26894
rect 579 26756 635 26812
rect 677 26756 733 26812
rect 775 26756 831 26812
rect 579 26674 635 26730
rect 677 26674 733 26730
rect 775 26674 831 26730
rect 579 26592 635 26648
rect 677 26592 733 26648
rect 775 26592 831 26648
rect 579 26510 635 26566
rect 677 26510 733 26566
rect 775 26510 831 26566
rect 579 26428 635 26484
rect 677 26428 733 26484
rect 775 26428 831 26484
rect 242 26287 298 26343
rect 334 26287 390 26343
rect 426 26287 482 26343
rect 518 26287 574 26343
rect 610 26287 666 26343
rect 702 26287 758 26343
rect 242 26207 298 26263
rect 334 26207 390 26263
rect 426 26207 482 26263
rect 518 26207 574 26263
rect 610 26207 666 26263
rect 702 26207 758 26263
rect 242 26127 298 26183
rect 334 26127 390 26183
rect 426 26127 482 26183
rect 518 26127 574 26183
rect 610 26127 666 26183
rect 702 26127 758 26183
rect 242 26047 298 26103
rect 334 26047 390 26103
rect 426 26047 482 26103
rect 518 26047 574 26103
rect 610 26047 666 26103
rect 702 26047 758 26103
rect 242 25967 298 26023
rect 334 25967 390 26023
rect 426 25967 482 26023
rect 518 25967 574 26023
rect 610 25967 666 26023
rect 702 25967 758 26023
rect 242 25887 298 25943
rect 334 25887 390 25943
rect 426 25887 482 25943
rect 518 25887 574 25943
rect 610 25887 666 25943
rect 702 25887 758 25943
rect 242 25807 298 25863
rect 334 25807 390 25863
rect 426 25807 482 25863
rect 518 25807 574 25863
rect 610 25807 666 25863
rect 702 25807 758 25863
rect 242 25727 298 25783
rect 334 25727 390 25783
rect 426 25727 482 25783
rect 518 25727 574 25783
rect 610 25727 666 25783
rect 702 25727 758 25783
rect 242 25647 298 25703
rect 334 25647 390 25703
rect 426 25647 482 25703
rect 518 25647 574 25703
rect 610 25647 666 25703
rect 702 25647 758 25703
rect 242 25567 298 25623
rect 334 25567 390 25623
rect 426 25567 482 25623
rect 518 25567 574 25623
rect 610 25567 666 25623
rect 702 25567 758 25623
rect 242 25487 298 25543
rect 334 25487 390 25543
rect 426 25487 482 25543
rect 518 25487 574 25543
rect 610 25487 666 25543
rect 702 25487 758 25543
rect 242 25407 298 25463
rect 334 25407 390 25463
rect 426 25407 482 25463
rect 518 25407 574 25463
rect 610 25407 666 25463
rect 702 25407 758 25463
rect 242 25327 298 25383
rect 334 25327 390 25383
rect 426 25327 482 25383
rect 518 25327 574 25383
rect 610 25327 666 25383
rect 702 25327 758 25383
rect 242 25247 298 25303
rect 334 25247 390 25303
rect 426 25247 482 25303
rect 518 25247 574 25303
rect 610 25247 666 25303
rect 702 25247 758 25303
rect 242 25167 298 25223
rect 334 25167 390 25223
rect 426 25167 482 25223
rect 518 25167 574 25223
rect 610 25167 666 25223
rect 702 25167 758 25223
rect 242 25087 298 25143
rect 334 25087 390 25143
rect 426 25087 482 25143
rect 518 25087 574 25143
rect 610 25087 666 25143
rect 702 25087 758 25143
rect 242 25007 298 25063
rect 334 25007 390 25063
rect 426 25007 482 25063
rect 518 25007 574 25063
rect 610 25007 666 25063
rect 702 25007 758 25063
rect 242 24927 298 24983
rect 334 24927 390 24983
rect 426 24927 482 24983
rect 518 24927 574 24983
rect 610 24927 666 24983
rect 702 24927 758 24983
rect 242 24847 298 24903
rect 334 24847 390 24903
rect 426 24847 482 24903
rect 518 24847 574 24903
rect 610 24847 666 24903
rect 702 24847 758 24903
rect 242 24767 298 24823
rect 334 24767 390 24823
rect 426 24767 482 24823
rect 518 24767 574 24823
rect 610 24767 666 24823
rect 702 24767 758 24823
rect 242 24687 298 24743
rect 334 24687 390 24743
rect 426 24687 482 24743
rect 518 24687 574 24743
rect 610 24687 666 24743
rect 702 24687 758 24743
rect 242 24607 298 24663
rect 334 24607 390 24663
rect 426 24607 482 24663
rect 518 24607 574 24663
rect 610 24607 666 24663
rect 702 24607 758 24663
rect 242 24527 298 24583
rect 334 24527 390 24583
rect 426 24527 482 24583
rect 518 24527 574 24583
rect 610 24527 666 24583
rect 702 24527 758 24583
rect 242 24447 298 24503
rect 334 24447 390 24503
rect 426 24447 482 24503
rect 518 24447 574 24503
rect 610 24447 666 24503
rect 702 24447 758 24503
rect 3494 28056 3550 28112
rect 4485 28057 4541 28113
rect 3494 27886 3550 27942
rect 4485 27888 4541 27944
rect 3494 27716 3550 27772
rect 4485 27718 4541 27774
rect 3494 27546 3550 27602
rect 4485 27548 4541 27604
rect 3494 27376 3550 27432
rect 4485 27378 4541 27434
rect 3494 27243 3550 27262
rect 4485 27243 4541 27264
rect 3494 27206 3530 27243
rect 3530 27206 3546 27243
rect 3546 27206 3550 27243
rect 4485 27208 4490 27243
rect 4490 27208 4541 27243
rect 5477 28581 5513 28620
rect 5513 28581 5528 28620
rect 5528 28581 5533 28620
rect 6469 28581 6472 28620
rect 6472 28581 6524 28620
rect 6524 28581 6525 28620
rect 5477 28564 5533 28581
rect 6469 28564 6525 28581
rect 5477 28433 5513 28453
rect 5513 28433 5528 28453
rect 5528 28433 5533 28453
rect 6469 28433 6472 28453
rect 6472 28433 6524 28453
rect 6524 28433 6525 28453
rect 5477 28397 5533 28433
rect 6469 28397 6525 28433
rect 5477 28230 5533 28286
rect 6469 28230 6525 28286
rect 5477 28063 5533 28119
rect 6469 28063 6525 28119
rect 5477 27896 5533 27952
rect 6469 27896 6525 27952
rect 5477 27729 5533 27785
rect 6469 27729 6525 27785
rect 5477 27562 5533 27618
rect 6469 27562 6525 27618
rect 5477 27395 5533 27451
rect 6469 27395 6525 27451
rect 5477 27243 5533 27283
rect 6469 27243 6525 27283
rect 5477 27227 5513 27243
rect 5513 27227 5529 27243
rect 5529 27227 5533 27243
rect 6469 27227 6473 27243
rect 6473 27227 6525 27243
rect 7461 28581 7497 28620
rect 7497 28581 7512 28620
rect 7512 28581 7517 28620
rect 8453 28581 8456 28620
rect 8456 28581 8508 28620
rect 8508 28581 8509 28620
rect 7461 28564 7517 28581
rect 8453 28564 8509 28581
rect 7461 28433 7497 28453
rect 7497 28433 7512 28453
rect 7512 28433 7517 28453
rect 8453 28433 8456 28453
rect 8456 28433 8508 28453
rect 8508 28433 8509 28453
rect 7461 28397 7517 28433
rect 8453 28397 8509 28433
rect 7461 28230 7517 28286
rect 8453 28230 8509 28286
rect 7461 28063 7517 28119
rect 8453 28063 8509 28119
rect 7461 27896 7517 27952
rect 8453 27896 8509 27952
rect 7461 27729 7517 27785
rect 8453 27729 8509 27785
rect 7461 27562 7517 27618
rect 8453 27562 8509 27618
rect 7461 27395 7517 27451
rect 8453 27395 8509 27451
rect 7461 27243 7517 27283
rect 8453 27243 8509 27283
rect 7461 27227 7497 27243
rect 7497 27227 7513 27243
rect 7513 27227 7517 27243
rect 8453 27227 8457 27243
rect 8457 27227 8509 27243
rect 9445 28581 9481 28620
rect 9481 28581 9501 28620
rect 9445 28564 9501 28581
rect 9445 28433 9481 28453
rect 9481 28433 9501 28453
rect 9445 28397 9501 28433
rect 9445 28230 9501 28286
rect 14283 28575 14334 28577
rect 14334 28575 14339 28577
rect 14381 28575 14410 28577
rect 14410 28575 14434 28577
rect 14434 28575 14437 28577
rect 14479 28575 14486 28577
rect 14486 28575 14510 28577
rect 14510 28575 14535 28577
rect 14577 28575 14586 28577
rect 14586 28575 14633 28577
rect 14283 28562 14339 28575
rect 14381 28562 14437 28575
rect 14479 28562 14535 28575
rect 14577 28562 14633 28575
rect 14283 28521 14334 28562
rect 14334 28521 14339 28562
rect 14381 28521 14410 28562
rect 14410 28521 14434 28562
rect 14434 28521 14437 28562
rect 14479 28521 14486 28562
rect 14486 28521 14510 28562
rect 14510 28521 14535 28562
rect 14577 28521 14586 28562
rect 14586 28521 14633 28562
rect 14283 28445 14334 28497
rect 14334 28445 14339 28497
rect 14381 28445 14410 28497
rect 14410 28445 14434 28497
rect 14434 28445 14437 28497
rect 14479 28445 14486 28497
rect 14486 28445 14510 28497
rect 14510 28445 14535 28497
rect 14577 28445 14586 28497
rect 14586 28445 14633 28497
rect 14283 28441 14339 28445
rect 14381 28441 14437 28445
rect 14479 28441 14535 28445
rect 14577 28441 14633 28445
rect 14283 28380 14334 28417
rect 14334 28380 14339 28417
rect 14381 28380 14410 28417
rect 14410 28380 14434 28417
rect 14434 28380 14437 28417
rect 14479 28380 14486 28417
rect 14486 28380 14510 28417
rect 14510 28380 14535 28417
rect 14577 28380 14586 28417
rect 14586 28380 14633 28417
rect 14283 28367 14339 28380
rect 14381 28367 14437 28380
rect 14479 28367 14535 28380
rect 14577 28367 14633 28380
rect 14283 28361 14334 28367
rect 14334 28361 14339 28367
rect 14381 28361 14410 28367
rect 14410 28361 14434 28367
rect 14434 28361 14437 28367
rect 14479 28361 14486 28367
rect 14486 28361 14510 28367
rect 14510 28361 14535 28367
rect 14577 28361 14586 28367
rect 14586 28361 14633 28367
rect 14283 28315 14334 28337
rect 14334 28315 14339 28337
rect 14381 28315 14410 28337
rect 14410 28315 14434 28337
rect 14434 28315 14437 28337
rect 14479 28315 14486 28337
rect 14486 28315 14510 28337
rect 14510 28315 14535 28337
rect 14577 28315 14586 28337
rect 14586 28315 14633 28337
rect 14283 28302 14339 28315
rect 14381 28302 14437 28315
rect 14479 28302 14535 28315
rect 14577 28302 14633 28315
rect 14283 28281 14334 28302
rect 14334 28281 14339 28302
rect 14381 28281 14410 28302
rect 14410 28281 14434 28302
rect 14434 28281 14437 28302
rect 14479 28281 14486 28302
rect 14486 28281 14510 28302
rect 14510 28281 14535 28302
rect 14577 28281 14586 28302
rect 14586 28281 14633 28302
rect 14283 28250 14334 28257
rect 14334 28250 14339 28257
rect 14381 28250 14410 28257
rect 14410 28250 14434 28257
rect 14434 28250 14437 28257
rect 14479 28250 14486 28257
rect 14486 28250 14510 28257
rect 14510 28250 14535 28257
rect 14577 28250 14586 28257
rect 14586 28250 14633 28257
rect 14283 28237 14339 28250
rect 14381 28237 14437 28250
rect 14479 28237 14535 28250
rect 14577 28237 14633 28250
rect 14283 28201 14334 28237
rect 14334 28201 14339 28237
rect 14381 28201 14410 28237
rect 14410 28201 14434 28237
rect 14434 28201 14437 28237
rect 14479 28201 14486 28237
rect 14486 28201 14510 28237
rect 14510 28201 14535 28237
rect 14577 28201 14586 28237
rect 14586 28201 14633 28237
rect 14283 28171 14339 28177
rect 14381 28171 14437 28177
rect 14479 28171 14535 28177
rect 14577 28171 14633 28177
rect 9445 28063 9501 28119
rect 9445 27896 9501 27952
rect 9445 27729 9501 27785
rect 9445 27562 9501 27618
rect 9445 27395 9501 27451
rect 9445 27268 9501 27283
rect 9445 27227 9475 27268
rect 9475 27227 9501 27268
rect 2387 27095 2443 27151
rect 2513 27095 2569 27151
rect 2387 27000 2443 27031
rect 2513 27000 2569 27031
rect 2387 26975 2417 27000
rect 2417 26975 2440 27000
rect 2440 26975 2443 27000
rect 2513 26975 2515 27000
rect 2515 26975 2567 27000
rect 2567 26975 2569 27000
rect 2387 26878 2443 26911
rect 2513 26878 2569 26911
rect 2387 26855 2417 26878
rect 2417 26855 2440 26878
rect 2440 26855 2443 26878
rect 2513 26855 2515 26878
rect 2515 26855 2567 26878
rect 2567 26855 2569 26878
rect 2485 26129 2532 26176
rect 2532 26129 2541 26176
rect 2611 26129 2620 26176
rect 2620 26129 2667 26176
rect 2485 26120 2541 26129
rect 2611 26120 2667 26129
rect 2485 26059 2532 26081
rect 2532 26059 2541 26081
rect 2611 26059 2620 26081
rect 2620 26059 2667 26081
rect 2485 26041 2541 26059
rect 2611 26041 2667 26059
rect 2485 26025 2532 26041
rect 2532 26025 2541 26041
rect 2611 26025 2620 26041
rect 2620 26025 2667 26041
rect 2485 25971 2541 25986
rect 2611 25971 2667 25986
rect 2485 25930 2532 25971
rect 2532 25930 2541 25971
rect 2611 25930 2620 25971
rect 2620 25930 2667 25971
rect 2485 25849 2532 25891
rect 2532 25849 2541 25891
rect 2611 25849 2620 25891
rect 2620 25849 2667 25891
rect 2485 25835 2541 25849
rect 2611 25835 2667 25849
rect 2485 25779 2532 25795
rect 2532 25779 2541 25795
rect 2611 25779 2620 25795
rect 2620 25779 2667 25795
rect 2485 25760 2541 25779
rect 2611 25760 2667 25779
rect 2485 25739 2532 25760
rect 2532 25739 2541 25760
rect 2611 25739 2620 25760
rect 2620 25739 2667 25760
rect 2485 25689 2541 25699
rect 2611 25689 2667 25699
rect 2485 25643 2532 25689
rect 2532 25643 2541 25689
rect 2611 25643 2620 25689
rect 2620 25643 2667 25689
rect 3477 26129 3524 26176
rect 3524 26129 3533 26176
rect 3603 26129 3612 26176
rect 3612 26129 3659 26176
rect 3477 26120 3533 26129
rect 3603 26120 3659 26129
rect 3477 26059 3524 26081
rect 3524 26059 3533 26081
rect 3603 26059 3612 26081
rect 3612 26059 3659 26081
rect 3477 26041 3533 26059
rect 3603 26041 3659 26059
rect 3477 26025 3524 26041
rect 3524 26025 3533 26041
rect 3603 26025 3612 26041
rect 3612 26025 3659 26041
rect 3477 25971 3533 25986
rect 3603 25971 3659 25986
rect 3477 25930 3524 25971
rect 3524 25930 3533 25971
rect 3603 25930 3612 25971
rect 3612 25930 3659 25971
rect 3477 25849 3524 25891
rect 3524 25849 3533 25891
rect 3603 25849 3612 25891
rect 3612 25849 3659 25891
rect 3477 25835 3533 25849
rect 3603 25835 3659 25849
rect 3477 25779 3524 25795
rect 3524 25779 3533 25795
rect 3603 25779 3612 25795
rect 3612 25779 3659 25795
rect 3477 25760 3533 25779
rect 3603 25760 3659 25779
rect 3477 25739 3524 25760
rect 3524 25739 3533 25760
rect 3603 25739 3612 25760
rect 3612 25739 3659 25760
rect 3477 25689 3533 25699
rect 3603 25689 3659 25699
rect 3477 25643 3524 25689
rect 3524 25643 3533 25689
rect 3603 25643 3612 25689
rect 3612 25643 3659 25689
rect 4469 26129 4516 26176
rect 4516 26129 4525 26176
rect 4595 26129 4604 26176
rect 4604 26129 4651 26176
rect 4469 26120 4525 26129
rect 4595 26120 4651 26129
rect 4469 26059 4516 26081
rect 4516 26059 4525 26081
rect 4595 26059 4604 26081
rect 4604 26059 4651 26081
rect 4469 26041 4525 26059
rect 4595 26041 4651 26059
rect 4469 26025 4516 26041
rect 4516 26025 4525 26041
rect 4595 26025 4604 26041
rect 4604 26025 4651 26041
rect 4469 25971 4525 25986
rect 4595 25971 4651 25986
rect 4469 25930 4516 25971
rect 4516 25930 4525 25971
rect 4595 25930 4604 25971
rect 4604 25930 4651 25971
rect 4469 25849 4516 25891
rect 4516 25849 4525 25891
rect 4595 25849 4604 25891
rect 4604 25849 4651 25891
rect 4469 25835 4525 25849
rect 4595 25835 4651 25849
rect 4469 25779 4516 25795
rect 4516 25779 4525 25795
rect 4595 25779 4604 25795
rect 4604 25779 4651 25795
rect 4469 25760 4525 25779
rect 4595 25760 4651 25779
rect 4469 25739 4516 25760
rect 4516 25739 4525 25760
rect 4595 25739 4604 25760
rect 4604 25739 4651 25760
rect 4469 25689 4525 25699
rect 4595 25689 4651 25699
rect 4469 25643 4516 25689
rect 4516 25643 4525 25689
rect 4595 25643 4604 25689
rect 4604 25643 4651 25689
rect 5461 26129 5508 26176
rect 5508 26129 5517 26176
rect 5587 26129 5596 26176
rect 5596 26129 5643 26176
rect 5461 26120 5517 26129
rect 5587 26120 5643 26129
rect 5461 26059 5508 26081
rect 5508 26059 5517 26081
rect 5587 26059 5596 26081
rect 5596 26059 5643 26081
rect 5461 26041 5517 26059
rect 5587 26041 5643 26059
rect 5461 26025 5508 26041
rect 5508 26025 5517 26041
rect 5587 26025 5596 26041
rect 5596 26025 5643 26041
rect 5461 25971 5517 25986
rect 5587 25971 5643 25986
rect 5461 25930 5508 25971
rect 5508 25930 5517 25971
rect 5587 25930 5596 25971
rect 5596 25930 5643 25971
rect 5461 25849 5508 25891
rect 5508 25849 5517 25891
rect 5587 25849 5596 25891
rect 5596 25849 5643 25891
rect 5461 25835 5517 25849
rect 5587 25835 5643 25849
rect 5461 25779 5508 25795
rect 5508 25779 5517 25795
rect 5587 25779 5596 25795
rect 5596 25779 5643 25795
rect 5461 25760 5517 25779
rect 5587 25760 5643 25779
rect 5461 25739 5508 25760
rect 5508 25739 5517 25760
rect 5587 25739 5596 25760
rect 5596 25739 5643 25760
rect 5461 25689 5517 25699
rect 5587 25689 5643 25699
rect 5461 25643 5508 25689
rect 5508 25643 5517 25689
rect 5587 25643 5596 25689
rect 5596 25643 5643 25689
rect 6453 26129 6500 26176
rect 6500 26129 6509 26176
rect 6579 26129 6588 26176
rect 6588 26129 6635 26176
rect 6453 26120 6509 26129
rect 6579 26120 6635 26129
rect 6453 26059 6500 26081
rect 6500 26059 6509 26081
rect 6579 26059 6588 26081
rect 6588 26059 6635 26081
rect 6453 26041 6509 26059
rect 6579 26041 6635 26059
rect 6453 26025 6500 26041
rect 6500 26025 6509 26041
rect 6579 26025 6588 26041
rect 6588 26025 6635 26041
rect 6453 25971 6509 25986
rect 6579 25971 6635 25986
rect 6453 25930 6500 25971
rect 6500 25930 6509 25971
rect 6579 25930 6588 25971
rect 6588 25930 6635 25971
rect 6453 25849 6500 25891
rect 6500 25849 6509 25891
rect 6579 25849 6588 25891
rect 6588 25849 6635 25891
rect 6453 25835 6509 25849
rect 6579 25835 6635 25849
rect 6453 25779 6500 25795
rect 6500 25779 6509 25795
rect 6579 25779 6588 25795
rect 6588 25779 6635 25795
rect 6453 25760 6509 25779
rect 6579 25760 6635 25779
rect 6453 25739 6500 25760
rect 6500 25739 6509 25760
rect 6579 25739 6588 25760
rect 6588 25739 6635 25760
rect 6453 25689 6509 25699
rect 6579 25689 6635 25699
rect 6453 25643 6500 25689
rect 6500 25643 6509 25689
rect 6579 25643 6588 25689
rect 6588 25643 6635 25689
rect 7445 26129 7492 26176
rect 7492 26129 7501 26176
rect 7571 26129 7580 26176
rect 7580 26129 7627 26176
rect 7445 26120 7501 26129
rect 7571 26120 7627 26129
rect 7445 26059 7492 26081
rect 7492 26059 7501 26081
rect 7571 26059 7580 26081
rect 7580 26059 7627 26081
rect 7445 26041 7501 26059
rect 7571 26041 7627 26059
rect 7445 26025 7492 26041
rect 7492 26025 7501 26041
rect 7571 26025 7580 26041
rect 7580 26025 7627 26041
rect 7445 25971 7501 25986
rect 7571 25971 7627 25986
rect 7445 25930 7492 25971
rect 7492 25930 7501 25971
rect 7571 25930 7580 25971
rect 7580 25930 7627 25971
rect 7445 25849 7492 25891
rect 7492 25849 7501 25891
rect 7571 25849 7580 25891
rect 7580 25849 7627 25891
rect 7445 25835 7501 25849
rect 7571 25835 7627 25849
rect 7445 25779 7492 25795
rect 7492 25779 7501 25795
rect 7571 25779 7580 25795
rect 7580 25779 7627 25795
rect 7445 25760 7501 25779
rect 7571 25760 7627 25779
rect 7445 25739 7492 25760
rect 7492 25739 7501 25760
rect 7571 25739 7580 25760
rect 7580 25739 7627 25760
rect 7445 25689 7501 25699
rect 7571 25689 7627 25699
rect 7445 25643 7492 25689
rect 7492 25643 7501 25689
rect 7571 25643 7580 25689
rect 7580 25643 7627 25689
rect 8437 26129 8484 26176
rect 8484 26129 8493 26176
rect 8563 26129 8572 26176
rect 8572 26129 8619 26176
rect 8437 26120 8493 26129
rect 8563 26120 8619 26129
rect 8437 26059 8484 26081
rect 8484 26059 8493 26081
rect 8563 26059 8572 26081
rect 8572 26059 8619 26081
rect 8437 26041 8493 26059
rect 8563 26041 8619 26059
rect 8437 26025 8484 26041
rect 8484 26025 8493 26041
rect 8563 26025 8572 26041
rect 8572 26025 8619 26041
rect 8437 25971 8493 25986
rect 8563 25971 8619 25986
rect 8437 25930 8484 25971
rect 8484 25930 8493 25971
rect 8563 25930 8572 25971
rect 8572 25930 8619 25971
rect 8437 25849 8484 25891
rect 8484 25849 8493 25891
rect 8563 25849 8572 25891
rect 8572 25849 8619 25891
rect 8437 25835 8493 25849
rect 8563 25835 8619 25849
rect 8437 25779 8484 25795
rect 8484 25779 8493 25795
rect 8563 25779 8572 25795
rect 8572 25779 8619 25795
rect 8437 25760 8493 25779
rect 8563 25760 8619 25779
rect 8437 25739 8484 25760
rect 8484 25739 8493 25760
rect 8563 25739 8572 25760
rect 8572 25739 8619 25760
rect 8437 25689 8493 25699
rect 8563 25689 8619 25699
rect 8437 25643 8484 25689
rect 8484 25643 8493 25689
rect 8563 25643 8572 25689
rect 8572 25643 8619 25689
rect 9429 26129 9476 26176
rect 9476 26129 9485 26176
rect 9555 26129 9564 26176
rect 9564 26129 9611 26176
rect 9429 26120 9485 26129
rect 9555 26120 9611 26129
rect 9429 26059 9476 26081
rect 9476 26059 9485 26081
rect 9555 26059 9564 26081
rect 9564 26059 9611 26081
rect 9429 26041 9485 26059
rect 9555 26041 9611 26059
rect 9429 26025 9476 26041
rect 9476 26025 9485 26041
rect 9555 26025 9564 26041
rect 9564 26025 9611 26041
rect 9429 25971 9485 25986
rect 9555 25971 9611 25986
rect 9429 25930 9476 25971
rect 9476 25930 9485 25971
rect 9555 25930 9564 25971
rect 9564 25930 9611 25971
rect 9429 25849 9476 25891
rect 9476 25849 9485 25891
rect 9555 25849 9564 25891
rect 9564 25849 9611 25891
rect 9429 25835 9485 25849
rect 9555 25835 9611 25849
rect 9429 25779 9476 25795
rect 9476 25779 9485 25795
rect 9555 25779 9564 25795
rect 9564 25779 9611 25795
rect 9429 25760 9485 25779
rect 9555 25760 9611 25779
rect 9429 25739 9476 25760
rect 9476 25739 9485 25760
rect 9555 25739 9564 25760
rect 9564 25739 9611 25760
rect 9429 25689 9485 25699
rect 9555 25689 9611 25699
rect 9429 25643 9476 25689
rect 9476 25643 9485 25689
rect 9555 25643 9564 25689
rect 9564 25643 9611 25689
rect 14283 28121 14334 28171
rect 14334 28121 14339 28171
rect 14381 28121 14410 28171
rect 14410 28121 14434 28171
rect 14434 28121 14437 28171
rect 14479 28121 14486 28171
rect 14486 28121 14510 28171
rect 14510 28121 14535 28171
rect 14577 28121 14586 28171
rect 14586 28121 14633 28171
rect 14283 28053 14334 28097
rect 14334 28053 14339 28097
rect 14381 28053 14410 28097
rect 14410 28053 14434 28097
rect 14434 28053 14437 28097
rect 14479 28053 14486 28097
rect 14486 28053 14510 28097
rect 14510 28053 14535 28097
rect 14577 28053 14586 28097
rect 14586 28053 14633 28097
rect 14283 28041 14339 28053
rect 14381 28041 14437 28053
rect 14479 28041 14535 28053
rect 14577 28041 14633 28053
rect 14283 27987 14334 28017
rect 14334 27987 14339 28017
rect 14381 27987 14410 28017
rect 14410 27987 14434 28017
rect 14434 27987 14437 28017
rect 14479 27987 14486 28017
rect 14486 27987 14510 28017
rect 14510 27987 14535 28017
rect 14577 27987 14586 28017
rect 14586 27987 14633 28017
rect 14283 27973 14339 27987
rect 14381 27973 14437 27987
rect 14479 27973 14535 27987
rect 14577 27973 14633 27987
rect 14283 27961 14334 27973
rect 14334 27961 14339 27973
rect 14381 27961 14410 27973
rect 14410 27961 14434 27973
rect 14434 27961 14437 27973
rect 14479 27961 14486 27973
rect 14486 27961 14510 27973
rect 14510 27961 14535 27973
rect 14577 27961 14586 27973
rect 14586 27961 14633 27973
rect 14283 27921 14334 27937
rect 14334 27921 14339 27937
rect 14381 27921 14410 27937
rect 14410 27921 14434 27937
rect 14434 27921 14437 27937
rect 14479 27921 14486 27937
rect 14486 27921 14510 27937
rect 14510 27921 14535 27937
rect 14577 27921 14586 27937
rect 14586 27921 14633 27937
rect 14283 27907 14339 27921
rect 14381 27907 14437 27921
rect 14479 27907 14535 27921
rect 14577 27907 14633 27921
rect 14283 27881 14334 27907
rect 14334 27881 14339 27907
rect 14381 27881 14410 27907
rect 14410 27881 14434 27907
rect 14434 27881 14437 27907
rect 14479 27881 14486 27907
rect 14486 27881 14510 27907
rect 14510 27881 14535 27907
rect 14577 27881 14586 27907
rect 14586 27881 14633 27907
rect 14283 27855 14334 27857
rect 14334 27855 14339 27857
rect 14381 27855 14410 27857
rect 14410 27855 14434 27857
rect 14434 27855 14437 27857
rect 14479 27855 14486 27857
rect 14486 27855 14510 27857
rect 14510 27855 14535 27857
rect 14577 27855 14586 27857
rect 14586 27855 14633 27857
rect 14283 27841 14339 27855
rect 14381 27841 14437 27855
rect 14479 27841 14535 27855
rect 14577 27841 14633 27855
rect 14283 27801 14334 27841
rect 14334 27801 14339 27841
rect 14381 27801 14410 27841
rect 14410 27801 14434 27841
rect 14434 27801 14437 27841
rect 14479 27801 14486 27841
rect 14486 27801 14510 27841
rect 14510 27801 14535 27841
rect 14577 27801 14586 27841
rect 14586 27801 14633 27841
rect 14283 27775 14339 27777
rect 14381 27775 14437 27777
rect 14479 27775 14535 27777
rect 14577 27775 14633 27777
rect 14283 27723 14334 27775
rect 14334 27723 14339 27775
rect 14381 27723 14410 27775
rect 14410 27723 14434 27775
rect 14434 27723 14437 27775
rect 14479 27723 14486 27775
rect 14486 27723 14510 27775
rect 14510 27723 14535 27775
rect 14577 27723 14586 27775
rect 14586 27723 14633 27775
rect 14283 27721 14339 27723
rect 14381 27721 14437 27723
rect 14479 27721 14535 27723
rect 14577 27721 14633 27723
rect 14283 27657 14334 27697
rect 14334 27657 14339 27697
rect 14381 27657 14410 27697
rect 14410 27657 14434 27697
rect 14434 27657 14437 27697
rect 14479 27657 14486 27697
rect 14486 27657 14510 27697
rect 14510 27657 14535 27697
rect 14577 27657 14586 27697
rect 14586 27657 14633 27697
rect 14283 27643 14339 27657
rect 14381 27643 14437 27657
rect 14479 27643 14535 27657
rect 14577 27643 14633 27657
rect 14283 27641 14334 27643
rect 14334 27641 14339 27643
rect 14381 27641 14410 27643
rect 14410 27641 14434 27643
rect 14434 27641 14437 27643
rect 14479 27641 14486 27643
rect 14486 27641 14510 27643
rect 14510 27641 14535 27643
rect 14577 27641 14586 27643
rect 14586 27641 14633 27643
rect 14283 27591 14334 27617
rect 14334 27591 14339 27617
rect 14381 27591 14410 27617
rect 14410 27591 14434 27617
rect 14434 27591 14437 27617
rect 14479 27591 14486 27617
rect 14486 27591 14510 27617
rect 14510 27591 14535 27617
rect 14577 27591 14586 27617
rect 14586 27591 14633 27617
rect 14283 27577 14339 27591
rect 14381 27577 14437 27591
rect 14479 27577 14535 27591
rect 14577 27577 14633 27591
rect 14283 27561 14334 27577
rect 14334 27561 14339 27577
rect 14381 27561 14410 27577
rect 14410 27561 14434 27577
rect 14434 27561 14437 27577
rect 14479 27561 14486 27577
rect 14486 27561 14510 27577
rect 14510 27561 14535 27577
rect 14577 27561 14586 27577
rect 14586 27561 14633 27577
rect 14283 27525 14334 27537
rect 14334 27525 14339 27537
rect 14381 27525 14410 27537
rect 14410 27525 14434 27537
rect 14434 27525 14437 27537
rect 14479 27525 14486 27537
rect 14486 27525 14510 27537
rect 14510 27525 14535 27537
rect 14577 27525 14586 27537
rect 14586 27525 14633 27537
rect 14283 27511 14339 27525
rect 14381 27511 14437 27525
rect 14479 27511 14535 27525
rect 14577 27511 14633 27525
rect 14283 27481 14334 27511
rect 14334 27481 14339 27511
rect 14381 27481 14410 27511
rect 14410 27481 14434 27511
rect 14434 27481 14437 27511
rect 14479 27481 14486 27511
rect 14486 27481 14510 27511
rect 14510 27481 14535 27511
rect 14577 27481 14586 27511
rect 14586 27481 14633 27511
rect 14283 27445 14339 27457
rect 14381 27445 14437 27457
rect 14479 27445 14535 27457
rect 14577 27445 14633 27457
rect 14283 27401 14334 27445
rect 14334 27401 14339 27445
rect 14381 27401 14410 27445
rect 14410 27401 14434 27445
rect 14434 27401 14437 27445
rect 14479 27401 14486 27445
rect 14486 27401 14510 27445
rect 14510 27401 14535 27445
rect 14577 27401 14586 27445
rect 14586 27401 14633 27445
rect 14283 27327 14334 27377
rect 14334 27327 14339 27377
rect 14381 27327 14410 27377
rect 14410 27327 14434 27377
rect 14434 27327 14437 27377
rect 14479 27327 14486 27377
rect 14486 27327 14510 27377
rect 14510 27327 14535 27377
rect 14577 27327 14586 27377
rect 14586 27327 14633 27377
rect 14283 27321 14339 27327
rect 14381 27321 14437 27327
rect 14479 27321 14535 27327
rect 14577 27321 14633 27327
rect 14283 27261 14334 27297
rect 14334 27261 14339 27297
rect 14381 27261 14410 27297
rect 14410 27261 14434 27297
rect 14434 27261 14437 27297
rect 14479 27261 14486 27297
rect 14486 27261 14510 27297
rect 14510 27261 14535 27297
rect 14577 27261 14586 27297
rect 14586 27261 14633 27297
rect 14283 27247 14339 27261
rect 14381 27247 14437 27261
rect 14479 27247 14535 27261
rect 14577 27247 14633 27261
rect 14283 27241 14334 27247
rect 14334 27241 14339 27247
rect 14381 27241 14410 27247
rect 14410 27241 14434 27247
rect 14434 27241 14437 27247
rect 14479 27241 14486 27247
rect 14486 27241 14510 27247
rect 14510 27241 14535 27247
rect 14577 27241 14586 27247
rect 14586 27241 14633 27247
rect 14283 27195 14334 27217
rect 14334 27195 14339 27217
rect 14381 27195 14410 27217
rect 14410 27195 14434 27217
rect 14434 27195 14437 27217
rect 14479 27195 14486 27217
rect 14486 27195 14510 27217
rect 14510 27195 14535 27217
rect 14577 27195 14586 27217
rect 14586 27195 14633 27217
rect 14283 27161 14339 27195
rect 14381 27161 14437 27195
rect 14479 27161 14535 27195
rect 14577 27161 14633 27195
rect 14283 27081 14339 27137
rect 14381 27081 14437 27137
rect 14479 27081 14535 27137
rect 14577 27081 14633 27137
rect 14283 27001 14339 27057
rect 14381 27001 14437 27057
rect 14479 27001 14535 27057
rect 14577 27001 14633 27057
rect 14283 26921 14339 26977
rect 14381 26921 14437 26977
rect 14479 26921 14535 26977
rect 14577 26921 14633 26977
rect 13651 26828 13707 26884
rect 13733 26828 13789 26884
rect 13815 26828 13871 26884
rect 13897 26828 13953 26884
rect 13979 26828 14035 26884
rect 13651 26744 13707 26800
rect 13733 26744 13789 26800
rect 13815 26744 13871 26800
rect 13897 26744 13953 26800
rect 13979 26744 14035 26800
rect 13651 26660 13707 26716
rect 13733 26660 13789 26716
rect 13815 26660 13871 26716
rect 13897 26660 13953 26716
rect 13979 26660 14035 26716
rect 13651 26576 13707 26632
rect 13733 26576 13789 26632
rect 13815 26576 13871 26632
rect 13897 26576 13953 26632
rect 13979 26576 14035 26632
rect 13651 26492 13707 26548
rect 13733 26492 13789 26548
rect 13815 26492 13871 26548
rect 13897 26492 13953 26548
rect 13979 26492 14035 26548
rect 14283 26841 14339 26897
rect 14381 26841 14437 26897
rect 14479 26841 14535 26897
rect 14577 26841 14633 26897
rect 14283 26761 14339 26817
rect 14381 26761 14437 26817
rect 14479 26761 14535 26817
rect 14577 26761 14633 26817
rect 14283 26681 14339 26737
rect 14381 26681 14437 26737
rect 14479 26681 14535 26737
rect 14577 26681 14633 26737
rect 14283 26601 14339 26657
rect 14381 26601 14437 26657
rect 14479 26601 14535 26657
rect 14577 26601 14633 26657
rect 14283 26520 14339 26576
rect 14381 26520 14437 26576
rect 14479 26520 14535 26576
rect 14577 26520 14633 26576
rect 14283 26439 14339 26495
rect 14381 26439 14437 26495
rect 14479 26439 14535 26495
rect 14577 26439 14633 26495
rect 14283 26358 14339 26414
rect 14381 26358 14437 26414
rect 14479 26358 14535 26414
rect 14577 26358 14633 26414
rect 14283 26277 14339 26333
rect 14381 26277 14437 26333
rect 14479 26277 14535 26333
rect 14577 26277 14633 26333
rect 14283 26196 14339 26252
rect 14381 26196 14437 26252
rect 14479 26196 14535 26252
rect 14577 26196 14633 26252
rect 14283 26115 14339 26171
rect 14381 26115 14437 26171
rect 14479 26115 14535 26171
rect 14577 26115 14633 26171
rect 14283 26034 14339 26090
rect 14381 26034 14437 26090
rect 14479 26034 14535 26090
rect 14577 26034 14633 26090
rect 14283 25953 14339 26009
rect 14381 25953 14437 26009
rect 14479 25953 14535 26009
rect 14577 25953 14633 26009
rect 14283 25872 14339 25928
rect 14381 25872 14437 25928
rect 14479 25872 14535 25928
rect 14577 25872 14633 25928
rect 14283 25791 14339 25847
rect 14381 25791 14437 25847
rect 14479 25791 14535 25847
rect 14577 25791 14633 25847
rect 14283 25710 14339 25766
rect 14381 25710 14437 25766
rect 14479 25710 14535 25766
rect 14577 25710 14633 25766
rect 14283 25629 14339 25685
rect 14381 25629 14437 25685
rect 14479 25629 14535 25685
rect 14577 25629 14633 25685
rect 14283 25548 14339 25604
rect 14381 25548 14437 25604
rect 14479 25548 14535 25604
rect 14577 25548 14633 25604
rect 14283 25467 14339 25523
rect 14381 25467 14437 25523
rect 14479 25467 14535 25523
rect 14577 25467 14633 25523
rect 14283 25386 14339 25442
rect 14381 25386 14437 25442
rect 14479 25386 14535 25442
rect 14577 25386 14633 25442
rect 14283 25305 14339 25361
rect 14381 25305 14437 25361
rect 14479 25305 14535 25361
rect 14577 25305 14633 25361
rect 14283 25224 14339 25280
rect 14381 25224 14437 25280
rect 14479 25224 14535 25280
rect 14577 25224 14633 25280
rect 14283 25143 14339 25199
rect 14381 25143 14437 25199
rect 14479 25143 14535 25199
rect 14577 25143 14633 25199
rect 14283 25062 14339 25118
rect 14381 25062 14437 25118
rect 14479 25062 14535 25118
rect 14577 25062 14633 25118
rect 14283 24981 14339 25037
rect 14381 24981 14437 25037
rect 14479 24981 14535 25037
rect 14577 24981 14633 25037
rect 14283 24900 14339 24956
rect 14381 24900 14437 24956
rect 14479 24900 14535 24956
rect 14577 24900 14633 24956
rect 14283 24819 14339 24875
rect 14381 24819 14437 24875
rect 14479 24819 14535 24875
rect 14577 24819 14633 24875
rect 14283 24738 14339 24794
rect 14381 24738 14437 24794
rect 14479 24738 14535 24794
rect 14577 24738 14633 24794
rect 14283 24657 14339 24713
rect 14381 24657 14437 24713
rect 14479 24657 14535 24713
rect 14577 24657 14633 24713
rect 14283 24576 14339 24632
rect 14381 24576 14437 24632
rect 14479 24576 14535 24632
rect 14577 24576 14633 24632
rect 14283 24495 14339 24551
rect 14381 24495 14437 24551
rect 14479 24495 14535 24551
rect 14577 24495 14633 24551
rect 242 24367 298 24423
rect 334 24367 390 24423
rect 426 24367 482 24423
rect 518 24367 574 24423
rect 610 24367 666 24423
rect 702 24367 758 24423
rect 242 24287 298 24343
rect 334 24287 390 24343
rect 426 24287 482 24343
rect 518 24287 574 24343
rect 610 24287 666 24343
rect 702 24287 758 24343
rect 242 24207 298 24263
rect 334 24207 390 24263
rect 426 24207 482 24263
rect 518 24207 574 24263
rect 610 24207 666 24263
rect 702 24207 758 24263
rect 242 24127 298 24183
rect 334 24127 390 24183
rect 426 24127 482 24183
rect 518 24127 574 24183
rect 610 24127 666 24183
rect 702 24127 758 24183
rect 242 24047 298 24103
rect 334 24047 390 24103
rect 426 24047 482 24103
rect 518 24047 574 24103
rect 610 24047 666 24103
rect 702 24047 758 24103
rect 242 23967 298 24023
rect 334 23967 390 24023
rect 426 23967 482 24023
rect 518 23967 574 24023
rect 610 23967 666 24023
rect 702 23967 758 24023
rect 242 23887 298 23943
rect 334 23887 390 23943
rect 426 23887 482 23943
rect 518 23887 574 23943
rect 610 23887 666 23943
rect 702 23887 758 23943
rect 242 23807 298 23863
rect 334 23807 390 23863
rect 426 23807 482 23863
rect 518 23807 574 23863
rect 610 23807 666 23863
rect 702 23807 758 23863
rect 242 23727 298 23783
rect 334 23727 390 23783
rect 426 23727 482 23783
rect 518 23727 574 23783
rect 610 23727 666 23783
rect 702 23727 758 23783
rect 242 23647 298 23703
rect 334 23647 390 23703
rect 426 23647 482 23703
rect 518 23647 574 23703
rect 610 23647 666 23703
rect 702 23647 758 23703
rect 14283 24414 14339 24470
rect 14381 24414 14437 24470
rect 14479 24414 14535 24470
rect 14577 24414 14633 24470
rect 14283 24333 14339 24389
rect 14381 24333 14437 24389
rect 14479 24333 14535 24389
rect 14577 24333 14633 24389
rect 14283 24252 14339 24308
rect 14381 24252 14437 24308
rect 14479 24252 14535 24308
rect 14577 24252 14633 24308
rect 14283 24171 14339 24227
rect 14381 24171 14437 24227
rect 14479 24171 14535 24227
rect 14577 24171 14633 24227
rect 14283 24090 14339 24146
rect 14381 24090 14437 24146
rect 14479 24090 14535 24146
rect 14577 24090 14633 24146
rect 14283 24009 14339 24065
rect 14381 24009 14437 24065
rect 14479 24009 14535 24065
rect 14577 24009 14633 24065
rect 14283 23928 14339 23984
rect 14381 23928 14437 23984
rect 14479 23928 14535 23984
rect 14577 23928 14633 23984
rect 14283 23847 14339 23903
rect 14381 23847 14437 23903
rect 14479 23847 14535 23903
rect 14577 23847 14633 23903
rect 14283 23766 14339 23822
rect 14381 23766 14437 23822
rect 14479 23766 14535 23822
rect 14577 23766 14633 23822
rect 242 23567 298 23623
rect 334 23567 390 23623
rect 426 23567 482 23623
rect 518 23567 574 23623
rect 610 23567 666 23623
rect 702 23567 758 23623
rect 242 23487 298 23543
rect 334 23487 390 23543
rect 426 23487 482 23543
rect 518 23487 574 23543
rect 610 23487 666 23543
rect 702 23487 758 23543
rect 242 23407 298 23463
rect 334 23407 390 23463
rect 426 23407 482 23463
rect 518 23407 574 23463
rect 610 23407 666 23463
rect 702 23407 758 23463
rect 242 23327 298 23383
rect 334 23327 390 23383
rect 426 23327 482 23383
rect 518 23327 574 23383
rect 610 23327 666 23383
rect 702 23327 758 23383
rect 242 23247 298 23303
rect 334 23247 390 23303
rect 426 23247 482 23303
rect 518 23247 574 23303
rect 610 23247 666 23303
rect 702 23247 758 23303
rect 242 23167 298 23223
rect 334 23167 390 23223
rect 426 23167 482 23223
rect 518 23167 574 23223
rect 610 23167 666 23223
rect 702 23167 758 23223
rect 242 23087 298 23143
rect 334 23087 390 23143
rect 426 23087 482 23143
rect 518 23087 574 23143
rect 610 23087 666 23143
rect 702 23087 758 23143
rect 242 23007 298 23063
rect 334 23007 390 23063
rect 426 23007 482 23063
rect 518 23007 574 23063
rect 610 23007 666 23063
rect 702 23007 758 23063
rect 242 22927 298 22983
rect 334 22927 390 22983
rect 426 22927 482 22983
rect 518 22927 574 22983
rect 610 22927 666 22983
rect 702 22927 758 22983
rect 242 22847 298 22903
rect 334 22847 390 22903
rect 426 22847 482 22903
rect 518 22847 574 22903
rect 610 22847 666 22903
rect 702 22847 758 22903
rect 242 22766 298 22822
rect 334 22766 390 22822
rect 426 22766 482 22822
rect 518 22766 574 22822
rect 610 22766 666 22822
rect 702 22766 758 22822
rect 242 22685 298 22741
rect 334 22685 390 22741
rect 426 22685 482 22741
rect 518 22685 574 22741
rect 610 22685 666 22741
rect 702 22685 758 22741
rect 242 22604 298 22660
rect 334 22604 390 22660
rect 426 22604 482 22660
rect 518 22604 574 22660
rect 610 22604 666 22660
rect 702 22604 758 22660
rect 242 22523 298 22579
rect 334 22523 390 22579
rect 426 22523 482 22579
rect 518 22523 574 22579
rect 610 22523 666 22579
rect 702 22523 758 22579
rect 242 22442 298 22498
rect 334 22442 390 22498
rect 426 22442 482 22498
rect 518 22442 574 22498
rect 610 22442 666 22498
rect 702 22442 758 22498
rect 242 22361 298 22417
rect 334 22361 390 22417
rect 426 22361 482 22417
rect 518 22361 574 22417
rect 610 22361 666 22417
rect 702 22361 758 22417
rect 242 22280 298 22336
rect 334 22280 390 22336
rect 426 22280 482 22336
rect 518 22280 574 22336
rect 610 22280 666 22336
rect 702 22280 758 22336
rect 242 22199 298 22255
rect 334 22199 390 22255
rect 426 22199 482 22255
rect 518 22199 574 22255
rect 610 22199 666 22255
rect 702 22199 758 22255
rect 242 22118 298 22174
rect 334 22118 390 22174
rect 426 22118 482 22174
rect 518 22118 574 22174
rect 610 22118 666 22174
rect 702 22118 758 22174
rect 242 22037 298 22093
rect 334 22037 390 22093
rect 426 22037 482 22093
rect 518 22037 574 22093
rect 610 22037 666 22093
rect 702 22037 758 22093
rect 242 21956 298 22012
rect 334 21956 390 22012
rect 426 21956 482 22012
rect 518 21956 574 22012
rect 610 21956 666 22012
rect 702 21956 758 22012
rect 242 21875 298 21931
rect 334 21875 390 21931
rect 426 21875 482 21931
rect 518 21875 574 21931
rect 610 21875 666 21931
rect 702 21875 758 21931
rect 242 21794 298 21850
rect 334 21794 390 21850
rect 426 21794 482 21850
rect 518 21794 574 21850
rect 610 21794 666 21850
rect 702 21794 758 21850
rect 242 21713 298 21769
rect 334 21713 390 21769
rect 426 21713 482 21769
rect 518 21713 574 21769
rect 610 21713 666 21769
rect 702 21713 758 21769
rect 242 21632 298 21688
rect 334 21632 390 21688
rect 426 21632 482 21688
rect 518 21632 574 21688
rect 610 21632 666 21688
rect 702 21632 758 21688
rect 242 21551 298 21607
rect 334 21551 390 21607
rect 426 21551 482 21607
rect 518 21551 574 21607
rect 610 21551 666 21607
rect 702 21551 758 21607
rect 242 21470 298 21526
rect 334 21470 390 21526
rect 426 21470 482 21526
rect 518 21470 574 21526
rect 610 21470 666 21526
rect 702 21470 758 21526
rect 242 21389 298 21445
rect 334 21389 390 21445
rect 426 21389 482 21445
rect 518 21389 574 21445
rect 610 21389 666 21445
rect 702 21389 758 21445
rect 242 21308 298 21364
rect 334 21308 390 21364
rect 426 21308 482 21364
rect 518 21308 574 21364
rect 610 21308 666 21364
rect 702 21308 758 21364
rect 242 21227 298 21283
rect 334 21227 390 21283
rect 426 21227 482 21283
rect 518 21227 574 21283
rect 610 21227 666 21283
rect 702 21227 758 21283
rect 242 21146 298 21202
rect 334 21146 390 21202
rect 426 21146 482 21202
rect 518 21146 574 21202
rect 610 21146 666 21202
rect 702 21146 758 21202
rect 1009 23630 1065 23686
rect 1111 23630 1167 23686
rect 1009 23550 1065 23606
rect 1111 23550 1167 23606
rect 1009 23470 1065 23526
rect 1111 23470 1167 23526
rect 1009 23390 1065 23446
rect 1111 23390 1167 23446
rect 1009 23310 1065 23366
rect 1111 23310 1167 23366
rect 1009 23230 1065 23286
rect 1111 23230 1167 23286
rect 1009 23150 1065 23206
rect 1111 23150 1167 23206
rect 1009 23070 1065 23126
rect 1111 23070 1167 23126
rect 1009 22990 1065 23046
rect 1111 22990 1167 23046
rect 1009 22910 1065 22966
rect 1111 22910 1167 22966
rect 1009 22830 1065 22886
rect 1111 22830 1167 22886
rect 1009 22750 1065 22806
rect 1111 22750 1167 22806
rect 1009 22670 1065 22726
rect 1111 22670 1167 22726
rect 1009 22590 1065 22646
rect 1111 22590 1167 22646
rect 1009 22510 1065 22566
rect 1111 22510 1167 22566
rect 1009 22430 1065 22486
rect 1111 22430 1167 22486
rect 1009 22350 1065 22406
rect 1111 22350 1167 22406
rect 1009 22270 1065 22326
rect 1111 22270 1167 22326
rect 1009 22189 1065 22245
rect 1111 22189 1167 22245
rect 1009 22108 1065 22164
rect 1111 22108 1167 22164
rect 1009 22027 1065 22083
rect 1111 22027 1167 22083
rect 1009 21946 1065 22002
rect 1111 21946 1167 22002
rect 1009 21865 1065 21921
rect 1111 21865 1167 21921
rect 1009 21784 1065 21840
rect 1111 21784 1167 21840
rect 1009 21703 1065 21759
rect 1111 21703 1167 21759
rect 1009 21622 1065 21678
rect 1111 21622 1167 21678
rect 1009 21541 1065 21597
rect 1111 21541 1167 21597
rect 1009 21460 1065 21516
rect 1111 21460 1167 21516
rect 1009 21379 1065 21435
rect 1111 21379 1167 21435
rect 1009 21298 1065 21354
rect 1111 21298 1167 21354
rect 1009 21217 1065 21273
rect 1111 21217 1167 21273
rect 1009 21136 1065 21192
rect 1111 21136 1167 21192
rect 1497 23630 1553 23686
rect 1615 23630 1671 23686
rect 1497 23550 1553 23606
rect 1615 23550 1671 23606
rect 1497 23470 1553 23526
rect 1615 23470 1671 23526
rect 1497 23390 1553 23446
rect 1615 23390 1671 23446
rect 1497 23310 1553 23366
rect 1615 23310 1671 23366
rect 1497 23230 1553 23286
rect 1615 23230 1671 23286
rect 1497 23150 1553 23206
rect 1615 23150 1671 23206
rect 1497 23070 1553 23126
rect 1615 23070 1671 23126
rect 1497 22990 1553 23046
rect 1615 22990 1671 23046
rect 1497 22910 1553 22966
rect 1615 22910 1671 22966
rect 1497 22830 1553 22886
rect 1615 22830 1671 22886
rect 1497 22750 1553 22806
rect 1615 22750 1671 22806
rect 1497 22670 1553 22726
rect 1615 22670 1671 22726
rect 1497 22590 1553 22646
rect 1615 22590 1671 22646
rect 1497 22510 1553 22566
rect 1615 22510 1671 22566
rect 1497 22430 1553 22486
rect 1615 22430 1671 22486
rect 1497 22350 1553 22406
rect 1615 22350 1671 22406
rect 1497 22270 1553 22326
rect 1615 22270 1671 22326
rect 1497 22189 1553 22245
rect 1615 22189 1671 22245
rect 1497 22108 1553 22164
rect 1615 22108 1671 22164
rect 1497 22027 1553 22083
rect 1615 22027 1671 22083
rect 1497 21946 1553 22002
rect 1615 21946 1671 22002
rect 1497 21865 1553 21921
rect 1615 21865 1671 21921
rect 1497 21784 1553 21840
rect 1615 21784 1671 21840
rect 1497 21703 1553 21759
rect 1615 21703 1671 21759
rect 1497 21622 1553 21678
rect 1615 21622 1671 21678
rect 1497 21541 1553 21597
rect 1615 21541 1671 21597
rect 1497 21460 1553 21516
rect 1615 21460 1671 21516
rect 1497 21379 1553 21435
rect 1615 21379 1671 21435
rect 1497 21298 1553 21354
rect 1615 21298 1671 21354
rect 1497 21217 1553 21273
rect 1615 21217 1671 21273
rect 1497 21136 1553 21192
rect 1615 21136 1671 21192
rect 1993 23630 2049 23686
rect 2111 23630 2167 23686
rect 1993 23550 2049 23606
rect 2111 23550 2167 23606
rect 1993 23470 2049 23526
rect 2111 23470 2167 23526
rect 1993 23390 2049 23446
rect 2111 23390 2167 23446
rect 1993 23310 2049 23366
rect 2111 23310 2167 23366
rect 1993 23230 2049 23286
rect 2111 23230 2167 23286
rect 1993 23150 2049 23206
rect 2111 23150 2167 23206
rect 1993 23070 2049 23126
rect 2111 23070 2167 23126
rect 1993 22990 2049 23046
rect 2111 22990 2167 23046
rect 1993 22910 2049 22966
rect 2111 22910 2167 22966
rect 1993 22830 2049 22886
rect 2111 22830 2167 22886
rect 1993 22750 2049 22806
rect 2111 22750 2167 22806
rect 1993 22670 2049 22726
rect 2111 22670 2167 22726
rect 1993 22590 2049 22646
rect 2111 22590 2167 22646
rect 1993 22510 2049 22566
rect 2111 22510 2167 22566
rect 1993 22430 2049 22486
rect 2111 22430 2167 22486
rect 1993 22350 2049 22406
rect 2111 22350 2167 22406
rect 1993 22270 2049 22326
rect 2111 22270 2167 22326
rect 1993 22189 2049 22245
rect 2111 22189 2167 22245
rect 1993 22108 2049 22164
rect 2111 22108 2167 22164
rect 1993 22027 2049 22083
rect 2111 22027 2167 22083
rect 1993 21946 2049 22002
rect 2111 21946 2167 22002
rect 1993 21865 2049 21921
rect 2111 21865 2167 21921
rect 1993 21784 2049 21840
rect 2111 21784 2167 21840
rect 1993 21703 2049 21759
rect 2111 21703 2167 21759
rect 1993 21622 2049 21678
rect 2111 21622 2167 21678
rect 1993 21541 2049 21597
rect 2111 21541 2167 21597
rect 1993 21460 2049 21516
rect 2111 21460 2167 21516
rect 1993 21379 2049 21435
rect 2111 21379 2167 21435
rect 1993 21298 2049 21354
rect 2111 21298 2167 21354
rect 1993 21217 2049 21273
rect 2111 21217 2167 21273
rect 1993 21136 2049 21192
rect 2111 21136 2167 21192
rect 2489 23630 2545 23686
rect 2607 23630 2663 23686
rect 2489 23550 2545 23606
rect 2607 23550 2663 23606
rect 2489 23470 2545 23526
rect 2607 23470 2663 23526
rect 2489 23390 2545 23446
rect 2607 23390 2663 23446
rect 2489 23310 2545 23366
rect 2607 23310 2663 23366
rect 2489 23230 2545 23286
rect 2607 23230 2663 23286
rect 2489 23150 2545 23206
rect 2607 23150 2663 23206
rect 2489 23070 2545 23126
rect 2607 23070 2663 23126
rect 2489 22990 2545 23046
rect 2607 22990 2663 23046
rect 2489 22910 2545 22966
rect 2607 22910 2663 22966
rect 2489 22830 2545 22886
rect 2607 22830 2663 22886
rect 2489 22750 2545 22806
rect 2607 22750 2663 22806
rect 2489 22670 2545 22726
rect 2607 22670 2663 22726
rect 2489 22590 2545 22646
rect 2607 22590 2663 22646
rect 2489 22510 2545 22566
rect 2607 22510 2663 22566
rect 2489 22430 2545 22486
rect 2607 22430 2663 22486
rect 2489 22350 2545 22406
rect 2607 22350 2663 22406
rect 2489 22270 2545 22326
rect 2607 22270 2663 22326
rect 2489 22189 2545 22245
rect 2607 22189 2663 22245
rect 2489 22108 2545 22164
rect 2607 22108 2663 22164
rect 2489 22027 2545 22083
rect 2607 22027 2663 22083
rect 2489 21946 2545 22002
rect 2607 21946 2663 22002
rect 2489 21865 2545 21921
rect 2607 21865 2663 21921
rect 2489 21784 2545 21840
rect 2607 21784 2663 21840
rect 2489 21703 2545 21759
rect 2607 21703 2663 21759
rect 2489 21622 2545 21678
rect 2607 21622 2663 21678
rect 2489 21541 2545 21597
rect 2607 21541 2663 21597
rect 2489 21460 2545 21516
rect 2607 21460 2663 21516
rect 2489 21379 2545 21435
rect 2607 21379 2663 21435
rect 2489 21298 2545 21354
rect 2607 21298 2663 21354
rect 2489 21217 2545 21273
rect 2607 21217 2663 21273
rect 2489 21136 2545 21192
rect 2607 21136 2663 21192
rect 2985 23630 3041 23686
rect 3103 23630 3159 23686
rect 2985 23550 3041 23606
rect 3103 23550 3159 23606
rect 2985 23470 3041 23526
rect 3103 23470 3159 23526
rect 2985 23390 3041 23446
rect 3103 23390 3159 23446
rect 2985 23310 3041 23366
rect 3103 23310 3159 23366
rect 2985 23230 3041 23286
rect 3103 23230 3159 23286
rect 2985 23150 3041 23206
rect 3103 23150 3159 23206
rect 2985 23070 3041 23126
rect 3103 23070 3159 23126
rect 2985 22990 3041 23046
rect 3103 22990 3159 23046
rect 2985 22910 3041 22966
rect 3103 22910 3159 22966
rect 2985 22830 3041 22886
rect 3103 22830 3159 22886
rect 2985 22750 3041 22806
rect 3103 22750 3159 22806
rect 2985 22670 3041 22726
rect 3103 22670 3159 22726
rect 2985 22590 3041 22646
rect 3103 22590 3159 22646
rect 2985 22510 3041 22566
rect 3103 22510 3159 22566
rect 2985 22430 3041 22486
rect 3103 22430 3159 22486
rect 2985 22350 3041 22406
rect 3103 22350 3159 22406
rect 2985 22270 3041 22326
rect 3103 22270 3159 22326
rect 2985 22189 3041 22245
rect 3103 22189 3159 22245
rect 2985 22108 3041 22164
rect 3103 22108 3159 22164
rect 2985 22027 3041 22083
rect 3103 22027 3159 22083
rect 2985 21946 3041 22002
rect 3103 21946 3159 22002
rect 2985 21865 3041 21921
rect 3103 21865 3159 21921
rect 2985 21784 3041 21840
rect 3103 21784 3159 21840
rect 2985 21703 3041 21759
rect 3103 21703 3159 21759
rect 2985 21622 3041 21678
rect 3103 21622 3159 21678
rect 2985 21541 3041 21597
rect 3103 21541 3159 21597
rect 2985 21460 3041 21516
rect 3103 21460 3159 21516
rect 2985 21379 3041 21435
rect 3103 21379 3159 21435
rect 2985 21298 3041 21354
rect 3103 21298 3159 21354
rect 2985 21217 3041 21273
rect 3103 21217 3159 21273
rect 2985 21136 3041 21192
rect 3103 21136 3159 21192
rect 3481 23630 3537 23686
rect 3599 23630 3655 23686
rect 3481 23550 3537 23606
rect 3599 23550 3655 23606
rect 3481 23470 3537 23526
rect 3599 23470 3655 23526
rect 3481 23390 3537 23446
rect 3599 23390 3655 23446
rect 3481 23310 3537 23366
rect 3599 23310 3655 23366
rect 3481 23230 3537 23286
rect 3599 23230 3655 23286
rect 3481 23150 3537 23206
rect 3599 23150 3655 23206
rect 3481 23070 3537 23126
rect 3599 23070 3655 23126
rect 3481 22990 3537 23046
rect 3599 22990 3655 23046
rect 3481 22910 3537 22966
rect 3599 22910 3655 22966
rect 3481 22830 3537 22886
rect 3599 22830 3655 22886
rect 3481 22750 3537 22806
rect 3599 22750 3655 22806
rect 3481 22670 3537 22726
rect 3599 22670 3655 22726
rect 3481 22590 3537 22646
rect 3599 22590 3655 22646
rect 3481 22510 3537 22566
rect 3599 22510 3655 22566
rect 3481 22430 3537 22486
rect 3599 22430 3655 22486
rect 3481 22350 3537 22406
rect 3599 22350 3655 22406
rect 3481 22270 3537 22326
rect 3599 22270 3655 22326
rect 3481 22189 3537 22245
rect 3599 22189 3655 22245
rect 3481 22108 3537 22164
rect 3599 22108 3655 22164
rect 3481 22027 3537 22083
rect 3599 22027 3655 22083
rect 3481 21946 3537 22002
rect 3599 21946 3655 22002
rect 3481 21865 3537 21921
rect 3599 21865 3655 21921
rect 3481 21784 3537 21840
rect 3599 21784 3655 21840
rect 3481 21703 3537 21759
rect 3599 21703 3655 21759
rect 3481 21622 3537 21678
rect 3599 21622 3655 21678
rect 3481 21541 3537 21597
rect 3599 21541 3655 21597
rect 3481 21460 3537 21516
rect 3599 21460 3655 21516
rect 3481 21379 3537 21435
rect 3599 21379 3655 21435
rect 3481 21298 3537 21354
rect 3599 21298 3655 21354
rect 3481 21217 3537 21273
rect 3599 21217 3655 21273
rect 3481 21136 3537 21192
rect 3599 21136 3655 21192
rect 3977 23630 4033 23686
rect 4095 23630 4151 23686
rect 3977 23550 4033 23606
rect 4095 23550 4151 23606
rect 3977 23470 4033 23526
rect 4095 23470 4151 23526
rect 3977 23390 4033 23446
rect 4095 23390 4151 23446
rect 3977 23310 4033 23366
rect 4095 23310 4151 23366
rect 3977 23230 4033 23286
rect 4095 23230 4151 23286
rect 3977 23150 4033 23206
rect 4095 23150 4151 23206
rect 3977 23070 4033 23126
rect 4095 23070 4151 23126
rect 3977 22990 4033 23046
rect 4095 22990 4151 23046
rect 3977 22910 4033 22966
rect 4095 22910 4151 22966
rect 3977 22830 4033 22886
rect 4095 22830 4151 22886
rect 3977 22750 4033 22806
rect 4095 22750 4151 22806
rect 3977 22670 4033 22726
rect 4095 22670 4151 22726
rect 3977 22590 4033 22646
rect 4095 22590 4151 22646
rect 3977 22510 4033 22566
rect 4095 22510 4151 22566
rect 3977 22430 4033 22486
rect 4095 22430 4151 22486
rect 3977 22350 4033 22406
rect 4095 22350 4151 22406
rect 3977 22270 4033 22326
rect 4095 22270 4151 22326
rect 3977 22189 4033 22245
rect 4095 22189 4151 22245
rect 3977 22108 4033 22164
rect 4095 22108 4151 22164
rect 3977 22027 4033 22083
rect 4095 22027 4151 22083
rect 3977 21946 4033 22002
rect 4095 21946 4151 22002
rect 3977 21865 4033 21921
rect 4095 21865 4151 21921
rect 3977 21784 4033 21840
rect 4095 21784 4151 21840
rect 3977 21703 4033 21759
rect 4095 21703 4151 21759
rect 3977 21622 4033 21678
rect 4095 21622 4151 21678
rect 3977 21541 4033 21597
rect 4095 21541 4151 21597
rect 3977 21460 4033 21516
rect 4095 21460 4151 21516
rect 3977 21379 4033 21435
rect 4095 21379 4151 21435
rect 3977 21298 4033 21354
rect 4095 21298 4151 21354
rect 3977 21217 4033 21273
rect 4095 21217 4151 21273
rect 3977 21136 4033 21192
rect 4095 21136 4151 21192
rect 4473 23630 4529 23686
rect 4591 23630 4647 23686
rect 4473 23550 4529 23606
rect 4591 23550 4647 23606
rect 4473 23470 4529 23526
rect 4591 23470 4647 23526
rect 4473 23390 4529 23446
rect 4591 23390 4647 23446
rect 4473 23310 4529 23366
rect 4591 23310 4647 23366
rect 4473 23230 4529 23286
rect 4591 23230 4647 23286
rect 4473 23150 4529 23206
rect 4591 23150 4647 23206
rect 4473 23070 4529 23126
rect 4591 23070 4647 23126
rect 4473 22990 4529 23046
rect 4591 22990 4647 23046
rect 4473 22910 4529 22966
rect 4591 22910 4647 22966
rect 4473 22830 4529 22886
rect 4591 22830 4647 22886
rect 4473 22750 4529 22806
rect 4591 22750 4647 22806
rect 4473 22670 4529 22726
rect 4591 22670 4647 22726
rect 4473 22590 4529 22646
rect 4591 22590 4647 22646
rect 4473 22510 4529 22566
rect 4591 22510 4647 22566
rect 4473 22430 4529 22486
rect 4591 22430 4647 22486
rect 4473 22350 4529 22406
rect 4591 22350 4647 22406
rect 4473 22270 4529 22326
rect 4591 22270 4647 22326
rect 4473 22189 4529 22245
rect 4591 22189 4647 22245
rect 4473 22108 4529 22164
rect 4591 22108 4647 22164
rect 4473 22027 4529 22083
rect 4591 22027 4647 22083
rect 4473 21946 4529 22002
rect 4591 21946 4647 22002
rect 4473 21865 4529 21921
rect 4591 21865 4647 21921
rect 4473 21784 4529 21840
rect 4591 21784 4647 21840
rect 4473 21703 4529 21759
rect 4591 21703 4647 21759
rect 4473 21622 4529 21678
rect 4591 21622 4647 21678
rect 4473 21541 4529 21597
rect 4591 21541 4647 21597
rect 4473 21460 4529 21516
rect 4591 21460 4647 21516
rect 4473 21379 4529 21435
rect 4591 21379 4647 21435
rect 4473 21298 4529 21354
rect 4591 21298 4647 21354
rect 4473 21217 4529 21273
rect 4591 21217 4647 21273
rect 4473 21136 4529 21192
rect 4591 21136 4647 21192
rect 4969 23630 5025 23686
rect 5087 23630 5143 23686
rect 4969 23550 5025 23606
rect 5087 23550 5143 23606
rect 4969 23470 5025 23526
rect 5087 23470 5143 23526
rect 4969 23390 5025 23446
rect 5087 23390 5143 23446
rect 4969 23310 5025 23366
rect 5087 23310 5143 23366
rect 4969 23230 5025 23286
rect 5087 23230 5143 23286
rect 4969 23150 5025 23206
rect 5087 23150 5143 23206
rect 4969 23070 5025 23126
rect 5087 23070 5143 23126
rect 4969 22990 5025 23046
rect 5087 22990 5143 23046
rect 4969 22910 5025 22966
rect 5087 22910 5143 22966
rect 4969 22830 5025 22886
rect 5087 22830 5143 22886
rect 4969 22750 5025 22806
rect 5087 22750 5143 22806
rect 4969 22670 5025 22726
rect 5087 22670 5143 22726
rect 4969 22590 5025 22646
rect 5087 22590 5143 22646
rect 4969 22510 5025 22566
rect 5087 22510 5143 22566
rect 4969 22430 5025 22486
rect 5087 22430 5143 22486
rect 4969 22350 5025 22406
rect 5087 22350 5143 22406
rect 4969 22270 5025 22326
rect 5087 22270 5143 22326
rect 4969 22189 5025 22245
rect 5087 22189 5143 22245
rect 4969 22108 5025 22164
rect 5087 22108 5143 22164
rect 4969 22027 5025 22083
rect 5087 22027 5143 22083
rect 4969 21946 5025 22002
rect 5087 21946 5143 22002
rect 4969 21865 5025 21921
rect 5087 21865 5143 21921
rect 4969 21784 5025 21840
rect 5087 21784 5143 21840
rect 4969 21703 5025 21759
rect 5087 21703 5143 21759
rect 4969 21622 5025 21678
rect 5087 21622 5143 21678
rect 4969 21541 5025 21597
rect 5087 21541 5143 21597
rect 4969 21460 5025 21516
rect 5087 21460 5143 21516
rect 4969 21379 5025 21435
rect 5087 21379 5143 21435
rect 4969 21298 5025 21354
rect 5087 21298 5143 21354
rect 4969 21217 5025 21273
rect 5087 21217 5143 21273
rect 4969 21136 5025 21192
rect 5087 21136 5143 21192
rect 5465 23630 5521 23686
rect 5583 23630 5639 23686
rect 5465 23550 5521 23606
rect 5583 23550 5639 23606
rect 5465 23470 5521 23526
rect 5583 23470 5639 23526
rect 5465 23390 5521 23446
rect 5583 23390 5639 23446
rect 5465 23310 5521 23366
rect 5583 23310 5639 23366
rect 5465 23230 5521 23286
rect 5583 23230 5639 23286
rect 5465 23150 5521 23206
rect 5583 23150 5639 23206
rect 5465 23070 5521 23126
rect 5583 23070 5639 23126
rect 5465 22990 5521 23046
rect 5583 22990 5639 23046
rect 5465 22910 5521 22966
rect 5583 22910 5639 22966
rect 5465 22830 5521 22886
rect 5583 22830 5639 22886
rect 5465 22750 5521 22806
rect 5583 22750 5639 22806
rect 5465 22670 5521 22726
rect 5583 22670 5639 22726
rect 5465 22590 5521 22646
rect 5583 22590 5639 22646
rect 5465 22510 5521 22566
rect 5583 22510 5639 22566
rect 5465 22430 5521 22486
rect 5583 22430 5639 22486
rect 5465 22350 5521 22406
rect 5583 22350 5639 22406
rect 5465 22270 5521 22326
rect 5583 22270 5639 22326
rect 5465 22189 5521 22245
rect 5583 22189 5639 22245
rect 5465 22108 5521 22164
rect 5583 22108 5639 22164
rect 5465 22027 5521 22083
rect 5583 22027 5639 22083
rect 5465 21946 5521 22002
rect 5583 21946 5639 22002
rect 5465 21865 5521 21921
rect 5583 21865 5639 21921
rect 5465 21784 5521 21840
rect 5583 21784 5639 21840
rect 5465 21703 5521 21759
rect 5583 21703 5639 21759
rect 5465 21622 5521 21678
rect 5583 21622 5639 21678
rect 5465 21541 5521 21597
rect 5583 21541 5639 21597
rect 5465 21460 5521 21516
rect 5583 21460 5639 21516
rect 5465 21379 5521 21435
rect 5583 21379 5639 21435
rect 5465 21298 5521 21354
rect 5583 21298 5639 21354
rect 5465 21217 5521 21273
rect 5583 21217 5639 21273
rect 5465 21136 5521 21192
rect 5583 21136 5639 21192
rect 5961 23630 6017 23686
rect 6079 23630 6135 23686
rect 5961 23550 6017 23606
rect 6079 23550 6135 23606
rect 5961 23470 6017 23526
rect 6079 23470 6135 23526
rect 5961 23390 6017 23446
rect 6079 23390 6135 23446
rect 5961 23310 6017 23366
rect 6079 23310 6135 23366
rect 5961 23230 6017 23286
rect 6079 23230 6135 23286
rect 5961 23150 6017 23206
rect 6079 23150 6135 23206
rect 5961 23070 6017 23126
rect 6079 23070 6135 23126
rect 5961 22990 6017 23046
rect 6079 22990 6135 23046
rect 5961 22910 6017 22966
rect 6079 22910 6135 22966
rect 5961 22830 6017 22886
rect 6079 22830 6135 22886
rect 5961 22750 6017 22806
rect 6079 22750 6135 22806
rect 5961 22670 6017 22726
rect 6079 22670 6135 22726
rect 5961 22590 6017 22646
rect 6079 22590 6135 22646
rect 5961 22510 6017 22566
rect 6079 22510 6135 22566
rect 5961 22430 6017 22486
rect 6079 22430 6135 22486
rect 5961 22350 6017 22406
rect 6079 22350 6135 22406
rect 5961 22270 6017 22326
rect 6079 22270 6135 22326
rect 5961 22189 6017 22245
rect 6079 22189 6135 22245
rect 5961 22108 6017 22164
rect 6079 22108 6135 22164
rect 5961 22027 6017 22083
rect 6079 22027 6135 22083
rect 5961 21946 6017 22002
rect 6079 21946 6135 22002
rect 5961 21865 6017 21921
rect 6079 21865 6135 21921
rect 5961 21784 6017 21840
rect 6079 21784 6135 21840
rect 5961 21703 6017 21759
rect 6079 21703 6135 21759
rect 5961 21622 6017 21678
rect 6079 21622 6135 21678
rect 5961 21541 6017 21597
rect 6079 21541 6135 21597
rect 5961 21460 6017 21516
rect 6079 21460 6135 21516
rect 5961 21379 6017 21435
rect 6079 21379 6135 21435
rect 5961 21298 6017 21354
rect 6079 21298 6135 21354
rect 5961 21217 6017 21273
rect 6079 21217 6135 21273
rect 5961 21136 6017 21192
rect 6079 21136 6135 21192
rect 6457 23630 6513 23686
rect 6575 23630 6631 23686
rect 6457 23550 6513 23606
rect 6575 23550 6631 23606
rect 6457 23470 6513 23526
rect 6575 23470 6631 23526
rect 6457 23390 6513 23446
rect 6575 23390 6631 23446
rect 6457 23310 6513 23366
rect 6575 23310 6631 23366
rect 6457 23230 6513 23286
rect 6575 23230 6631 23286
rect 6457 23150 6513 23206
rect 6575 23150 6631 23206
rect 6457 23070 6513 23126
rect 6575 23070 6631 23126
rect 6457 22990 6513 23046
rect 6575 22990 6631 23046
rect 6457 22910 6513 22966
rect 6575 22910 6631 22966
rect 6457 22830 6513 22886
rect 6575 22830 6631 22886
rect 6457 22750 6513 22806
rect 6575 22750 6631 22806
rect 6457 22670 6513 22726
rect 6575 22670 6631 22726
rect 6457 22590 6513 22646
rect 6575 22590 6631 22646
rect 6457 22510 6513 22566
rect 6575 22510 6631 22566
rect 6457 22430 6513 22486
rect 6575 22430 6631 22486
rect 6457 22350 6513 22406
rect 6575 22350 6631 22406
rect 6457 22270 6513 22326
rect 6575 22270 6631 22326
rect 6457 22189 6513 22245
rect 6575 22189 6631 22245
rect 6457 22108 6513 22164
rect 6575 22108 6631 22164
rect 6457 22027 6513 22083
rect 6575 22027 6631 22083
rect 6457 21946 6513 22002
rect 6575 21946 6631 22002
rect 6457 21865 6513 21921
rect 6575 21865 6631 21921
rect 6457 21784 6513 21840
rect 6575 21784 6631 21840
rect 6457 21703 6513 21759
rect 6575 21703 6631 21759
rect 6457 21622 6513 21678
rect 6575 21622 6631 21678
rect 6457 21541 6513 21597
rect 6575 21541 6631 21597
rect 6457 21460 6513 21516
rect 6575 21460 6631 21516
rect 6457 21379 6513 21435
rect 6575 21379 6631 21435
rect 6457 21298 6513 21354
rect 6575 21298 6631 21354
rect 6457 21217 6513 21273
rect 6575 21217 6631 21273
rect 6457 21136 6513 21192
rect 6575 21136 6631 21192
rect 6953 23630 7009 23686
rect 7071 23630 7127 23686
rect 6953 23550 7009 23606
rect 7071 23550 7127 23606
rect 6953 23470 7009 23526
rect 7071 23470 7127 23526
rect 6953 23390 7009 23446
rect 7071 23390 7127 23446
rect 6953 23310 7009 23366
rect 7071 23310 7127 23366
rect 6953 23230 7009 23286
rect 7071 23230 7127 23286
rect 6953 23150 7009 23206
rect 7071 23150 7127 23206
rect 6953 23070 7009 23126
rect 7071 23070 7127 23126
rect 6953 22990 7009 23046
rect 7071 22990 7127 23046
rect 6953 22910 7009 22966
rect 7071 22910 7127 22966
rect 6953 22830 7009 22886
rect 7071 22830 7127 22886
rect 6953 22750 7009 22806
rect 7071 22750 7127 22806
rect 6953 22670 7009 22726
rect 7071 22670 7127 22726
rect 6953 22590 7009 22646
rect 7071 22590 7127 22646
rect 6953 22510 7009 22566
rect 7071 22510 7127 22566
rect 6953 22430 7009 22486
rect 7071 22430 7127 22486
rect 6953 22350 7009 22406
rect 7071 22350 7127 22406
rect 6953 22270 7009 22326
rect 7071 22270 7127 22326
rect 6953 22189 7009 22245
rect 7071 22189 7127 22245
rect 6953 22108 7009 22164
rect 7071 22108 7127 22164
rect 6953 22027 7009 22083
rect 7071 22027 7127 22083
rect 6953 21946 7009 22002
rect 7071 21946 7127 22002
rect 6953 21865 7009 21921
rect 7071 21865 7127 21921
rect 6953 21784 7009 21840
rect 7071 21784 7127 21840
rect 6953 21703 7009 21759
rect 7071 21703 7127 21759
rect 6953 21622 7009 21678
rect 7071 21622 7127 21678
rect 6953 21541 7009 21597
rect 7071 21541 7127 21597
rect 6953 21460 7009 21516
rect 7071 21460 7127 21516
rect 6953 21379 7009 21435
rect 7071 21379 7127 21435
rect 6953 21298 7009 21354
rect 7071 21298 7127 21354
rect 6953 21217 7009 21273
rect 7071 21217 7127 21273
rect 6953 21136 7009 21192
rect 7071 21136 7127 21192
rect 7449 23630 7505 23686
rect 7567 23630 7623 23686
rect 7449 23550 7505 23606
rect 7567 23550 7623 23606
rect 7449 23470 7505 23526
rect 7567 23470 7623 23526
rect 7449 23390 7505 23446
rect 7567 23390 7623 23446
rect 7449 23310 7505 23366
rect 7567 23310 7623 23366
rect 7449 23230 7505 23286
rect 7567 23230 7623 23286
rect 7449 23150 7505 23206
rect 7567 23150 7623 23206
rect 7449 23070 7505 23126
rect 7567 23070 7623 23126
rect 7449 22990 7505 23046
rect 7567 22990 7623 23046
rect 7449 22910 7505 22966
rect 7567 22910 7623 22966
rect 7449 22830 7505 22886
rect 7567 22830 7623 22886
rect 7449 22750 7505 22806
rect 7567 22750 7623 22806
rect 7449 22670 7505 22726
rect 7567 22670 7623 22726
rect 7449 22590 7505 22646
rect 7567 22590 7623 22646
rect 7449 22510 7505 22566
rect 7567 22510 7623 22566
rect 7449 22430 7505 22486
rect 7567 22430 7623 22486
rect 7449 22350 7505 22406
rect 7567 22350 7623 22406
rect 7449 22270 7505 22326
rect 7567 22270 7623 22326
rect 7449 22189 7505 22245
rect 7567 22189 7623 22245
rect 7449 22108 7505 22164
rect 7567 22108 7623 22164
rect 7449 22027 7505 22083
rect 7567 22027 7623 22083
rect 7449 21946 7505 22002
rect 7567 21946 7623 22002
rect 7449 21865 7505 21921
rect 7567 21865 7623 21921
rect 7449 21784 7505 21840
rect 7567 21784 7623 21840
rect 7449 21703 7505 21759
rect 7567 21703 7623 21759
rect 7449 21622 7505 21678
rect 7567 21622 7623 21678
rect 7449 21541 7505 21597
rect 7567 21541 7623 21597
rect 7449 21460 7505 21516
rect 7567 21460 7623 21516
rect 7449 21379 7505 21435
rect 7567 21379 7623 21435
rect 7449 21298 7505 21354
rect 7567 21298 7623 21354
rect 7449 21217 7505 21273
rect 7567 21217 7623 21273
rect 7449 21136 7505 21192
rect 7567 21136 7623 21192
rect 7945 23630 8001 23686
rect 8063 23630 8119 23686
rect 7945 23550 8001 23606
rect 8063 23550 8119 23606
rect 7945 23470 8001 23526
rect 8063 23470 8119 23526
rect 7945 23390 8001 23446
rect 8063 23390 8119 23446
rect 7945 23310 8001 23366
rect 8063 23310 8119 23366
rect 7945 23230 8001 23286
rect 8063 23230 8119 23286
rect 7945 23150 8001 23206
rect 8063 23150 8119 23206
rect 7945 23070 8001 23126
rect 8063 23070 8119 23126
rect 7945 22990 8001 23046
rect 8063 22990 8119 23046
rect 7945 22910 8001 22966
rect 8063 22910 8119 22966
rect 7945 22830 8001 22886
rect 8063 22830 8119 22886
rect 7945 22750 8001 22806
rect 8063 22750 8119 22806
rect 7945 22670 8001 22726
rect 8063 22670 8119 22726
rect 7945 22590 8001 22646
rect 8063 22590 8119 22646
rect 7945 22510 8001 22566
rect 8063 22510 8119 22566
rect 7945 22430 8001 22486
rect 8063 22430 8119 22486
rect 7945 22350 8001 22406
rect 8063 22350 8119 22406
rect 7945 22270 8001 22326
rect 8063 22270 8119 22326
rect 7945 22189 8001 22245
rect 8063 22189 8119 22245
rect 7945 22108 8001 22164
rect 8063 22108 8119 22164
rect 7945 22027 8001 22083
rect 8063 22027 8119 22083
rect 7945 21946 8001 22002
rect 8063 21946 8119 22002
rect 7945 21865 8001 21921
rect 8063 21865 8119 21921
rect 7945 21784 8001 21840
rect 8063 21784 8119 21840
rect 7945 21703 8001 21759
rect 8063 21703 8119 21759
rect 7945 21622 8001 21678
rect 8063 21622 8119 21678
rect 7945 21541 8001 21597
rect 8063 21541 8119 21597
rect 7945 21460 8001 21516
rect 8063 21460 8119 21516
rect 7945 21379 8001 21435
rect 8063 21379 8119 21435
rect 7945 21298 8001 21354
rect 8063 21298 8119 21354
rect 7945 21217 8001 21273
rect 8063 21217 8119 21273
rect 7945 21136 8001 21192
rect 8063 21136 8119 21192
rect 8441 23630 8497 23686
rect 8559 23630 8615 23686
rect 8441 23550 8497 23606
rect 8559 23550 8615 23606
rect 8441 23470 8497 23526
rect 8559 23470 8615 23526
rect 8441 23390 8497 23446
rect 8559 23390 8615 23446
rect 8441 23310 8497 23366
rect 8559 23310 8615 23366
rect 8441 23230 8497 23286
rect 8559 23230 8615 23286
rect 8441 23150 8497 23206
rect 8559 23150 8615 23206
rect 8441 23070 8497 23126
rect 8559 23070 8615 23126
rect 8441 22990 8497 23046
rect 8559 22990 8615 23046
rect 8441 22910 8497 22966
rect 8559 22910 8615 22966
rect 8441 22830 8497 22886
rect 8559 22830 8615 22886
rect 8441 22750 8497 22806
rect 8559 22750 8615 22806
rect 8441 22670 8497 22726
rect 8559 22670 8615 22726
rect 8441 22590 8497 22646
rect 8559 22590 8615 22646
rect 8441 22510 8497 22566
rect 8559 22510 8615 22566
rect 8441 22430 8497 22486
rect 8559 22430 8615 22486
rect 8441 22350 8497 22406
rect 8559 22350 8615 22406
rect 8441 22270 8497 22326
rect 8559 22270 8615 22326
rect 8441 22189 8497 22245
rect 8559 22189 8615 22245
rect 8441 22108 8497 22164
rect 8559 22108 8615 22164
rect 8441 22027 8497 22083
rect 8559 22027 8615 22083
rect 8441 21946 8497 22002
rect 8559 21946 8615 22002
rect 8441 21865 8497 21921
rect 8559 21865 8615 21921
rect 8441 21784 8497 21840
rect 8559 21784 8615 21840
rect 8441 21703 8497 21759
rect 8559 21703 8615 21759
rect 8441 21622 8497 21678
rect 8559 21622 8615 21678
rect 8441 21541 8497 21597
rect 8559 21541 8615 21597
rect 8441 21460 8497 21516
rect 8559 21460 8615 21516
rect 8441 21379 8497 21435
rect 8559 21379 8615 21435
rect 8441 21298 8497 21354
rect 8559 21298 8615 21354
rect 8441 21217 8497 21273
rect 8559 21217 8615 21273
rect 8441 21136 8497 21192
rect 8559 21136 8615 21192
rect 8937 23630 8993 23686
rect 9055 23630 9111 23686
rect 8937 23550 8993 23606
rect 9055 23550 9111 23606
rect 8937 23470 8993 23526
rect 9055 23470 9111 23526
rect 8937 23390 8993 23446
rect 9055 23390 9111 23446
rect 8937 23310 8993 23366
rect 9055 23310 9111 23366
rect 8937 23230 8993 23286
rect 9055 23230 9111 23286
rect 8937 23150 8993 23206
rect 9055 23150 9111 23206
rect 8937 23070 8993 23126
rect 9055 23070 9111 23126
rect 8937 22990 8993 23046
rect 9055 22990 9111 23046
rect 8937 22910 8993 22966
rect 9055 22910 9111 22966
rect 8937 22830 8993 22886
rect 9055 22830 9111 22886
rect 8937 22750 8993 22806
rect 9055 22750 9111 22806
rect 8937 22670 8993 22726
rect 9055 22670 9111 22726
rect 8937 22590 8993 22646
rect 9055 22590 9111 22646
rect 8937 22510 8993 22566
rect 9055 22510 9111 22566
rect 8937 22430 8993 22486
rect 9055 22430 9111 22486
rect 8937 22350 8993 22406
rect 9055 22350 9111 22406
rect 8937 22270 8993 22326
rect 9055 22270 9111 22326
rect 8937 22189 8993 22245
rect 9055 22189 9111 22245
rect 8937 22108 8993 22164
rect 9055 22108 9111 22164
rect 8937 22027 8993 22083
rect 9055 22027 9111 22083
rect 8937 21946 8993 22002
rect 9055 21946 9111 22002
rect 8937 21865 8993 21921
rect 9055 21865 9111 21921
rect 8937 21784 8993 21840
rect 9055 21784 9111 21840
rect 8937 21703 8993 21759
rect 9055 21703 9111 21759
rect 8937 21622 8993 21678
rect 9055 21622 9111 21678
rect 8937 21541 8993 21597
rect 9055 21541 9111 21597
rect 8937 21460 8993 21516
rect 9055 21460 9111 21516
rect 8937 21379 8993 21435
rect 9055 21379 9111 21435
rect 8937 21298 8993 21354
rect 9055 21298 9111 21354
rect 8937 21217 8993 21273
rect 9055 21217 9111 21273
rect 8937 21136 8993 21192
rect 9055 21136 9111 21192
rect 9433 23630 9489 23686
rect 9551 23630 9607 23686
rect 9433 23550 9489 23606
rect 9551 23550 9607 23606
rect 9433 23470 9489 23526
rect 9551 23470 9607 23526
rect 9433 23390 9489 23446
rect 9551 23390 9607 23446
rect 9433 23310 9489 23366
rect 9551 23310 9607 23366
rect 9433 23230 9489 23286
rect 9551 23230 9607 23286
rect 9433 23150 9489 23206
rect 9551 23150 9607 23206
rect 9433 23070 9489 23126
rect 9551 23070 9607 23126
rect 9433 22990 9489 23046
rect 9551 22990 9607 23046
rect 9433 22910 9489 22966
rect 9551 22910 9607 22966
rect 9433 22830 9489 22886
rect 9551 22830 9607 22886
rect 9433 22750 9489 22806
rect 9551 22750 9607 22806
rect 9433 22670 9489 22726
rect 9551 22670 9607 22726
rect 9433 22590 9489 22646
rect 9551 22590 9607 22646
rect 9433 22510 9489 22566
rect 9551 22510 9607 22566
rect 9433 22430 9489 22486
rect 9551 22430 9607 22486
rect 9433 22350 9489 22406
rect 9551 22350 9607 22406
rect 9433 22270 9489 22326
rect 9551 22270 9607 22326
rect 9433 22189 9489 22245
rect 9551 22189 9607 22245
rect 9433 22108 9489 22164
rect 9551 22108 9607 22164
rect 9433 22027 9489 22083
rect 9551 22027 9607 22083
rect 9433 21946 9489 22002
rect 9551 21946 9607 22002
rect 9433 21865 9489 21921
rect 9551 21865 9607 21921
rect 9433 21784 9489 21840
rect 9551 21784 9607 21840
rect 9433 21703 9489 21759
rect 9551 21703 9607 21759
rect 9433 21622 9489 21678
rect 9551 21622 9607 21678
rect 9433 21541 9489 21597
rect 9551 21541 9607 21597
rect 9433 21460 9489 21516
rect 9551 21460 9607 21516
rect 9433 21379 9489 21435
rect 9551 21379 9607 21435
rect 9433 21298 9489 21354
rect 9551 21298 9607 21354
rect 9433 21217 9489 21273
rect 9551 21217 9607 21273
rect 9433 21136 9489 21192
rect 9551 21136 9607 21192
rect 9929 23630 9985 23686
rect 10047 23630 10103 23686
rect 9929 23550 9985 23606
rect 10047 23550 10103 23606
rect 9929 23470 9985 23526
rect 10047 23470 10103 23526
rect 9929 23390 9985 23446
rect 10047 23390 10103 23446
rect 9929 23310 9985 23366
rect 10047 23310 10103 23366
rect 9929 23230 9985 23286
rect 10047 23230 10103 23286
rect 9929 23150 9985 23206
rect 10047 23150 10103 23206
rect 9929 23070 9985 23126
rect 10047 23070 10103 23126
rect 9929 22990 9985 23046
rect 10047 22990 10103 23046
rect 9929 22910 9985 22966
rect 10047 22910 10103 22966
rect 9929 22830 9985 22886
rect 10047 22830 10103 22886
rect 9929 22750 9985 22806
rect 10047 22750 10103 22806
rect 9929 22670 9985 22726
rect 10047 22670 10103 22726
rect 9929 22590 9985 22646
rect 10047 22590 10103 22646
rect 9929 22510 9985 22566
rect 10047 22510 10103 22566
rect 9929 22430 9985 22486
rect 10047 22430 10103 22486
rect 9929 22350 9985 22406
rect 10047 22350 10103 22406
rect 9929 22270 9985 22326
rect 10047 22270 10103 22326
rect 9929 22189 9985 22245
rect 10047 22189 10103 22245
rect 9929 22108 9985 22164
rect 10047 22108 10103 22164
rect 9929 22027 9985 22083
rect 10047 22027 10103 22083
rect 9929 21946 9985 22002
rect 10047 21946 10103 22002
rect 9929 21865 9985 21921
rect 10047 21865 10103 21921
rect 9929 21784 9985 21840
rect 10047 21784 10103 21840
rect 9929 21703 9985 21759
rect 10047 21703 10103 21759
rect 9929 21622 9985 21678
rect 10047 21622 10103 21678
rect 9929 21541 9985 21597
rect 10047 21541 10103 21597
rect 9929 21460 9985 21516
rect 10047 21460 10103 21516
rect 9929 21379 9985 21435
rect 10047 21379 10103 21435
rect 9929 21298 9985 21354
rect 10047 21298 10103 21354
rect 9929 21217 9985 21273
rect 10047 21217 10103 21273
rect 9929 21136 9985 21192
rect 10047 21136 10103 21192
rect 10425 23630 10481 23686
rect 10543 23630 10599 23686
rect 10425 23550 10481 23606
rect 10543 23550 10599 23606
rect 10425 23470 10481 23526
rect 10543 23470 10599 23526
rect 10425 23390 10481 23446
rect 10543 23390 10599 23446
rect 10425 23310 10481 23366
rect 10543 23310 10599 23366
rect 10425 23230 10481 23286
rect 10543 23230 10599 23286
rect 10425 23150 10481 23206
rect 10543 23150 10599 23206
rect 10425 23070 10481 23126
rect 10543 23070 10599 23126
rect 10425 22990 10481 23046
rect 10543 22990 10599 23046
rect 10425 22910 10481 22966
rect 10543 22910 10599 22966
rect 10425 22830 10481 22886
rect 10543 22830 10599 22886
rect 10425 22750 10481 22806
rect 10543 22750 10599 22806
rect 10425 22670 10481 22726
rect 10543 22670 10599 22726
rect 10425 22590 10481 22646
rect 10543 22590 10599 22646
rect 10425 22510 10481 22566
rect 10543 22510 10599 22566
rect 10425 22430 10481 22486
rect 10543 22430 10599 22486
rect 10425 22350 10481 22406
rect 10543 22350 10599 22406
rect 10425 22270 10481 22326
rect 10543 22270 10599 22326
rect 10425 22189 10481 22245
rect 10543 22189 10599 22245
rect 10425 22108 10481 22164
rect 10543 22108 10599 22164
rect 10425 22027 10481 22083
rect 10543 22027 10599 22083
rect 10425 21946 10481 22002
rect 10543 21946 10599 22002
rect 10425 21865 10481 21921
rect 10543 21865 10599 21921
rect 10425 21784 10481 21840
rect 10543 21784 10599 21840
rect 10425 21703 10481 21759
rect 10543 21703 10599 21759
rect 10425 21622 10481 21678
rect 10543 21622 10599 21678
rect 10425 21541 10481 21597
rect 10543 21541 10599 21597
rect 10425 21460 10481 21516
rect 10543 21460 10599 21516
rect 10425 21379 10481 21435
rect 10543 21379 10599 21435
rect 10425 21298 10481 21354
rect 10543 21298 10599 21354
rect 10425 21217 10481 21273
rect 10543 21217 10599 21273
rect 10425 21136 10481 21192
rect 10543 21136 10599 21192
rect 10921 23630 10977 23686
rect 11039 23630 11095 23686
rect 10921 23550 10977 23606
rect 11039 23550 11095 23606
rect 10921 23470 10977 23526
rect 11039 23470 11095 23526
rect 10921 23390 10977 23446
rect 11039 23390 11095 23446
rect 10921 23310 10977 23366
rect 11039 23310 11095 23366
rect 10921 23230 10977 23286
rect 11039 23230 11095 23286
rect 10921 23150 10977 23206
rect 11039 23150 11095 23206
rect 10921 23070 10977 23126
rect 11039 23070 11095 23126
rect 10921 22990 10977 23046
rect 11039 22990 11095 23046
rect 10921 22910 10977 22966
rect 11039 22910 11095 22966
rect 10921 22830 10977 22886
rect 11039 22830 11095 22886
rect 10921 22750 10977 22806
rect 11039 22750 11095 22806
rect 10921 22670 10977 22726
rect 11039 22670 11095 22726
rect 10921 22590 10977 22646
rect 11039 22590 11095 22646
rect 10921 22510 10977 22566
rect 11039 22510 11095 22566
rect 10921 22430 10977 22486
rect 11039 22430 11095 22486
rect 10921 22350 10977 22406
rect 11039 22350 11095 22406
rect 10921 22270 10977 22326
rect 11039 22270 11095 22326
rect 10921 22189 10977 22245
rect 11039 22189 11095 22245
rect 10921 22108 10977 22164
rect 11039 22108 11095 22164
rect 10921 22027 10977 22083
rect 11039 22027 11095 22083
rect 10921 21946 10977 22002
rect 11039 21946 11095 22002
rect 10921 21865 10977 21921
rect 11039 21865 11095 21921
rect 10921 21784 10977 21840
rect 11039 21784 11095 21840
rect 10921 21703 10977 21759
rect 11039 21703 11095 21759
rect 10921 21622 10977 21678
rect 11039 21622 11095 21678
rect 10921 21541 10977 21597
rect 11039 21541 11095 21597
rect 10921 21460 10977 21516
rect 11039 21460 11095 21516
rect 10921 21379 10977 21435
rect 11039 21379 11095 21435
rect 10921 21298 10977 21354
rect 11039 21298 11095 21354
rect 10921 21217 10977 21273
rect 11039 21217 11095 21273
rect 10921 21136 10977 21192
rect 11039 21136 11095 21192
rect 11417 23630 11473 23686
rect 11535 23630 11591 23686
rect 11417 23550 11473 23606
rect 11535 23550 11591 23606
rect 11417 23470 11473 23526
rect 11535 23470 11591 23526
rect 11417 23390 11473 23446
rect 11535 23390 11591 23446
rect 11417 23310 11473 23366
rect 11535 23310 11591 23366
rect 11417 23230 11473 23286
rect 11535 23230 11591 23286
rect 11417 23150 11473 23206
rect 11535 23150 11591 23206
rect 11417 23070 11473 23126
rect 11535 23070 11591 23126
rect 11417 22990 11473 23046
rect 11535 22990 11591 23046
rect 11417 22910 11473 22966
rect 11535 22910 11591 22966
rect 11417 22830 11473 22886
rect 11535 22830 11591 22886
rect 11417 22750 11473 22806
rect 11535 22750 11591 22806
rect 11417 22670 11473 22726
rect 11535 22670 11591 22726
rect 11417 22590 11473 22646
rect 11535 22590 11591 22646
rect 11417 22510 11473 22566
rect 11535 22510 11591 22566
rect 11417 22430 11473 22486
rect 11535 22430 11591 22486
rect 11417 22350 11473 22406
rect 11535 22350 11591 22406
rect 11417 22270 11473 22326
rect 11535 22270 11591 22326
rect 11417 22189 11473 22245
rect 11535 22189 11591 22245
rect 11417 22108 11473 22164
rect 11535 22108 11591 22164
rect 11417 22027 11473 22083
rect 11535 22027 11591 22083
rect 11417 21946 11473 22002
rect 11535 21946 11591 22002
rect 11417 21865 11473 21921
rect 11535 21865 11591 21921
rect 11417 21784 11473 21840
rect 11535 21784 11591 21840
rect 11417 21703 11473 21759
rect 11535 21703 11591 21759
rect 11417 21622 11473 21678
rect 11535 21622 11591 21678
rect 11417 21541 11473 21597
rect 11535 21541 11591 21597
rect 11417 21460 11473 21516
rect 11535 21460 11591 21516
rect 11417 21379 11473 21435
rect 11535 21379 11591 21435
rect 11417 21298 11473 21354
rect 11535 21298 11591 21354
rect 11417 21217 11473 21273
rect 11535 21217 11591 21273
rect 11417 21136 11473 21192
rect 11535 21136 11591 21192
rect 11913 23630 11969 23686
rect 12031 23630 12087 23686
rect 11913 23550 11969 23606
rect 12031 23550 12087 23606
rect 11913 23470 11969 23526
rect 12031 23470 12087 23526
rect 11913 23390 11969 23446
rect 12031 23390 12087 23446
rect 11913 23310 11969 23366
rect 12031 23310 12087 23366
rect 11913 23230 11969 23286
rect 12031 23230 12087 23286
rect 11913 23150 11969 23206
rect 12031 23150 12087 23206
rect 11913 23070 11969 23126
rect 12031 23070 12087 23126
rect 11913 22990 11969 23046
rect 12031 22990 12087 23046
rect 11913 22910 11969 22966
rect 12031 22910 12087 22966
rect 11913 22830 11969 22886
rect 12031 22830 12087 22886
rect 11913 22750 11969 22806
rect 12031 22750 12087 22806
rect 11913 22670 11969 22726
rect 12031 22670 12087 22726
rect 11913 22590 11969 22646
rect 12031 22590 12087 22646
rect 11913 22510 11969 22566
rect 12031 22510 12087 22566
rect 11913 22430 11969 22486
rect 12031 22430 12087 22486
rect 11913 22350 11969 22406
rect 12031 22350 12087 22406
rect 11913 22270 11969 22326
rect 12031 22270 12087 22326
rect 11913 22189 11969 22245
rect 12031 22189 12087 22245
rect 11913 22108 11969 22164
rect 12031 22108 12087 22164
rect 11913 22027 11969 22083
rect 12031 22027 12087 22083
rect 11913 21946 11969 22002
rect 12031 21946 12087 22002
rect 11913 21865 11969 21921
rect 12031 21865 12087 21921
rect 11913 21784 11969 21840
rect 12031 21784 12087 21840
rect 11913 21703 11969 21759
rect 12031 21703 12087 21759
rect 11913 21622 11969 21678
rect 12031 21622 12087 21678
rect 11913 21541 11969 21597
rect 12031 21541 12087 21597
rect 11913 21460 11969 21516
rect 12031 21460 12087 21516
rect 11913 21379 11969 21435
rect 12031 21379 12087 21435
rect 11913 21298 11969 21354
rect 12031 21298 12087 21354
rect 11913 21217 11969 21273
rect 12031 21217 12087 21273
rect 11913 21136 11969 21192
rect 12031 21136 12087 21192
rect 12409 23630 12465 23686
rect 12527 23630 12583 23686
rect 12409 23550 12465 23606
rect 12527 23550 12583 23606
rect 12409 23470 12465 23526
rect 12527 23470 12583 23526
rect 12409 23390 12465 23446
rect 12527 23390 12583 23446
rect 12409 23310 12465 23366
rect 12527 23310 12583 23366
rect 12409 23230 12465 23286
rect 12527 23230 12583 23286
rect 12409 23150 12465 23206
rect 12527 23150 12583 23206
rect 12409 23070 12465 23126
rect 12527 23070 12583 23126
rect 12409 22990 12465 23046
rect 12527 22990 12583 23046
rect 12409 22910 12465 22966
rect 12527 22910 12583 22966
rect 12409 22830 12465 22886
rect 12527 22830 12583 22886
rect 12409 22750 12465 22806
rect 12527 22750 12583 22806
rect 12409 22670 12465 22726
rect 12527 22670 12583 22726
rect 12409 22590 12465 22646
rect 12527 22590 12583 22646
rect 12409 22510 12465 22566
rect 12527 22510 12583 22566
rect 12409 22430 12465 22486
rect 12527 22430 12583 22486
rect 12409 22350 12465 22406
rect 12527 22350 12583 22406
rect 12409 22270 12465 22326
rect 12527 22270 12583 22326
rect 12409 22189 12465 22245
rect 12527 22189 12583 22245
rect 12409 22108 12465 22164
rect 12527 22108 12583 22164
rect 12409 22027 12465 22083
rect 12527 22027 12583 22083
rect 12409 21946 12465 22002
rect 12527 21946 12583 22002
rect 12409 21865 12465 21921
rect 12527 21865 12583 21921
rect 12409 21784 12465 21840
rect 12527 21784 12583 21840
rect 12409 21703 12465 21759
rect 12527 21703 12583 21759
rect 12409 21622 12465 21678
rect 12527 21622 12583 21678
rect 12409 21541 12465 21597
rect 12527 21541 12583 21597
rect 12409 21460 12465 21516
rect 12527 21460 12583 21516
rect 12409 21379 12465 21435
rect 12527 21379 12583 21435
rect 12409 21298 12465 21354
rect 12527 21298 12583 21354
rect 12409 21217 12465 21273
rect 12527 21217 12583 21273
rect 12409 21136 12465 21192
rect 12527 21136 12583 21192
rect 12905 23630 12961 23686
rect 13023 23630 13079 23686
rect 12905 23550 12961 23606
rect 13023 23550 13079 23606
rect 12905 23470 12961 23526
rect 13023 23470 13079 23526
rect 12905 23390 12961 23446
rect 13023 23390 13079 23446
rect 12905 23310 12961 23366
rect 13023 23310 13079 23366
rect 12905 23230 12961 23286
rect 13023 23230 13079 23286
rect 12905 23150 12961 23206
rect 13023 23150 13079 23206
rect 12905 23070 12961 23126
rect 13023 23070 13079 23126
rect 12905 22990 12961 23046
rect 13023 22990 13079 23046
rect 12905 22910 12961 22966
rect 13023 22910 13079 22966
rect 12905 22830 12961 22886
rect 13023 22830 13079 22886
rect 12905 22750 12961 22806
rect 13023 22750 13079 22806
rect 12905 22670 12961 22726
rect 13023 22670 13079 22726
rect 12905 22590 12961 22646
rect 13023 22590 13079 22646
rect 12905 22510 12961 22566
rect 13023 22510 13079 22566
rect 12905 22430 12961 22486
rect 13023 22430 13079 22486
rect 12905 22350 12961 22406
rect 13023 22350 13079 22406
rect 12905 22270 12961 22326
rect 13023 22270 13079 22326
rect 12905 22189 12961 22245
rect 13023 22189 13079 22245
rect 12905 22108 12961 22164
rect 13023 22108 13079 22164
rect 12905 22027 12961 22083
rect 13023 22027 13079 22083
rect 12905 21946 12961 22002
rect 13023 21946 13079 22002
rect 12905 21865 12961 21921
rect 13023 21865 13079 21921
rect 12905 21784 12961 21840
rect 13023 21784 13079 21840
rect 12905 21703 12961 21759
rect 13023 21703 13079 21759
rect 12905 21622 12961 21678
rect 13023 21622 13079 21678
rect 12905 21541 12961 21597
rect 13023 21541 13079 21597
rect 12905 21460 12961 21516
rect 13023 21460 13079 21516
rect 12905 21379 12961 21435
rect 13023 21379 13079 21435
rect 12905 21298 12961 21354
rect 13023 21298 13079 21354
rect 12905 21217 12961 21273
rect 13023 21217 13079 21273
rect 12905 21136 12961 21192
rect 13023 21136 13079 21192
rect 13401 23630 13457 23686
rect 13519 23630 13575 23686
rect 13401 23550 13457 23606
rect 13519 23550 13575 23606
rect 13401 23470 13457 23526
rect 13519 23470 13575 23526
rect 13401 23390 13457 23446
rect 13519 23390 13575 23446
rect 13401 23310 13457 23366
rect 13519 23310 13575 23366
rect 13401 23230 13457 23286
rect 13519 23230 13575 23286
rect 13401 23150 13457 23206
rect 13519 23150 13575 23206
rect 13401 23070 13457 23126
rect 13519 23070 13575 23126
rect 13401 22990 13457 23046
rect 13519 22990 13575 23046
rect 13401 22910 13457 22966
rect 13519 22910 13575 22966
rect 13401 22830 13457 22886
rect 13519 22830 13575 22886
rect 13401 22750 13457 22806
rect 13519 22750 13575 22806
rect 13401 22670 13457 22726
rect 13519 22670 13575 22726
rect 13401 22590 13457 22646
rect 13519 22590 13575 22646
rect 13401 22510 13457 22566
rect 13519 22510 13575 22566
rect 13401 22430 13457 22486
rect 13519 22430 13575 22486
rect 13401 22350 13457 22406
rect 13519 22350 13575 22406
rect 13401 22270 13457 22326
rect 13519 22270 13575 22326
rect 13401 22189 13457 22245
rect 13519 22189 13575 22245
rect 13401 22108 13457 22164
rect 13519 22108 13575 22164
rect 13401 22027 13457 22083
rect 13519 22027 13575 22083
rect 13401 21946 13457 22002
rect 13519 21946 13575 22002
rect 13401 21865 13457 21921
rect 13519 21865 13575 21921
rect 13401 21784 13457 21840
rect 13519 21784 13575 21840
rect 13401 21703 13457 21759
rect 13519 21703 13575 21759
rect 13401 21622 13457 21678
rect 13519 21622 13575 21678
rect 13401 21541 13457 21597
rect 13519 21541 13575 21597
rect 13401 21460 13457 21516
rect 13519 21460 13575 21516
rect 13401 21379 13457 21435
rect 13519 21379 13575 21435
rect 13401 21298 13457 21354
rect 13519 21298 13575 21354
rect 13401 21217 13457 21273
rect 13519 21217 13575 21273
rect 13401 21136 13457 21192
rect 13519 21136 13575 21192
rect 13838 23630 13894 23686
rect 13956 23630 14012 23686
rect 13838 23550 13894 23606
rect 13956 23550 14012 23606
rect 13838 23470 13894 23526
rect 13956 23470 14012 23526
rect 13838 23390 13894 23446
rect 13956 23390 14012 23446
rect 13838 23310 13894 23366
rect 13956 23310 14012 23366
rect 13838 23230 13894 23286
rect 13956 23230 14012 23286
rect 13838 23150 13894 23206
rect 13956 23150 14012 23206
rect 13838 23070 13894 23126
rect 13956 23070 14012 23126
rect 13838 22990 13894 23046
rect 13956 22990 14012 23046
rect 13838 22910 13894 22966
rect 13956 22910 14012 22966
rect 13838 22830 13894 22886
rect 13956 22830 14012 22886
rect 13838 22750 13894 22806
rect 13956 22750 14012 22806
rect 13838 22670 13894 22726
rect 13956 22670 14012 22726
rect 13838 22590 13894 22646
rect 13956 22590 14012 22646
rect 13838 22510 13894 22566
rect 13956 22510 14012 22566
rect 13838 22430 13894 22486
rect 13956 22430 14012 22486
rect 13838 22350 13894 22406
rect 13956 22350 14012 22406
rect 13838 22270 13894 22326
rect 13956 22270 14012 22326
rect 13838 22189 13894 22245
rect 13956 22189 14012 22245
rect 13838 22108 13894 22164
rect 13956 22108 14012 22164
rect 13838 22027 13894 22083
rect 13956 22027 14012 22083
rect 13838 21946 13894 22002
rect 13956 21946 14012 22002
rect 13838 21865 13894 21921
rect 13956 21865 14012 21921
rect 13838 21784 13894 21840
rect 13956 21784 14012 21840
rect 13838 21703 13894 21759
rect 13956 21703 14012 21759
rect 13838 21622 13894 21678
rect 13956 21622 14012 21678
rect 13838 21541 13894 21597
rect 13956 21541 14012 21597
rect 13838 21460 13894 21516
rect 13956 21460 14012 21516
rect 13838 21379 13894 21435
rect 13956 21379 14012 21435
rect 13838 21298 13894 21354
rect 13956 21298 14012 21354
rect 13838 21217 13894 21273
rect 13956 21217 14012 21273
rect 13838 21136 13894 21192
rect 13956 21136 14012 21192
rect 14283 23685 14339 23741
rect 14381 23685 14437 23741
rect 14479 23685 14535 23741
rect 14577 23685 14633 23741
rect 14283 23604 14339 23660
rect 14381 23604 14437 23660
rect 14479 23604 14535 23660
rect 14577 23604 14633 23660
rect 14283 23523 14339 23579
rect 14381 23523 14437 23579
rect 14479 23523 14535 23579
rect 14577 23523 14633 23579
rect 14283 23442 14339 23498
rect 14381 23442 14437 23498
rect 14479 23442 14535 23498
rect 14577 23442 14633 23498
rect 14283 23361 14339 23417
rect 14381 23361 14437 23417
rect 14479 23361 14535 23417
rect 14577 23361 14633 23417
rect 14283 23280 14339 23336
rect 14381 23280 14437 23336
rect 14479 23280 14535 23336
rect 14577 23280 14633 23336
rect 14283 23199 14339 23255
rect 14381 23199 14437 23255
rect 14479 23199 14535 23255
rect 14577 23199 14633 23255
rect 14283 23118 14339 23174
rect 14381 23118 14437 23174
rect 14479 23118 14535 23174
rect 14577 23118 14633 23174
rect 14283 23037 14339 23093
rect 14381 23037 14437 23093
rect 14479 23037 14535 23093
rect 14577 23037 14633 23093
rect 14283 22956 14339 23012
rect 14381 22956 14437 23012
rect 14479 22956 14535 23012
rect 14577 22956 14633 23012
rect 14283 22875 14339 22931
rect 14381 22875 14437 22931
rect 14479 22875 14535 22931
rect 14577 22875 14633 22931
rect 14283 22794 14339 22850
rect 14381 22794 14437 22850
rect 14479 22794 14535 22850
rect 14577 22794 14633 22850
rect 14283 22713 14339 22769
rect 14381 22713 14437 22769
rect 14479 22713 14535 22769
rect 14577 22713 14633 22769
rect 14283 22632 14339 22688
rect 14381 22632 14437 22688
rect 14479 22632 14535 22688
rect 14577 22632 14633 22688
rect 14283 22551 14339 22607
rect 14381 22551 14437 22607
rect 14479 22551 14535 22607
rect 14577 22551 14633 22607
rect 14283 22470 14339 22526
rect 14381 22470 14437 22526
rect 14479 22470 14535 22526
rect 14577 22470 14633 22526
rect 14283 22389 14339 22445
rect 14381 22389 14437 22445
rect 14479 22389 14535 22445
rect 14577 22389 14633 22445
rect 14283 22308 14339 22364
rect 14381 22308 14437 22364
rect 14479 22308 14535 22364
rect 14577 22308 14633 22364
rect 14283 22227 14339 22283
rect 14381 22227 14437 22283
rect 14479 22227 14535 22283
rect 14577 22227 14633 22283
rect 14283 22146 14339 22202
rect 14381 22146 14437 22202
rect 14479 22146 14535 22202
rect 14577 22146 14633 22202
rect 14283 22065 14339 22121
rect 14381 22065 14437 22121
rect 14479 22065 14535 22121
rect 14577 22065 14633 22121
rect 14283 21984 14339 22040
rect 14381 21984 14437 22040
rect 14479 21984 14535 22040
rect 14577 21984 14633 22040
rect 14283 21903 14339 21959
rect 14381 21903 14437 21959
rect 14479 21903 14535 21959
rect 14577 21903 14633 21959
rect 14283 21822 14339 21878
rect 14381 21822 14437 21878
rect 14479 21822 14535 21878
rect 14577 21822 14633 21878
rect 14283 21741 14339 21797
rect 14381 21741 14437 21797
rect 14479 21741 14535 21797
rect 14577 21741 14633 21797
rect 14283 21660 14339 21716
rect 14381 21660 14437 21716
rect 14479 21660 14535 21716
rect 14577 21660 14633 21716
rect 14283 21579 14339 21635
rect 14381 21579 14437 21635
rect 14479 21579 14535 21635
rect 14577 21579 14633 21635
rect 14283 21498 14339 21554
rect 14381 21498 14437 21554
rect 14479 21498 14535 21554
rect 14577 21498 14633 21554
rect 14283 21417 14339 21473
rect 14381 21417 14437 21473
rect 14479 21417 14535 21473
rect 14577 21417 14633 21473
rect 14283 21336 14339 21392
rect 14381 21336 14437 21392
rect 14479 21336 14535 21392
rect 14577 21336 14633 21392
rect 14283 21255 14339 21311
rect 14381 21255 14437 21311
rect 14479 21255 14535 21311
rect 14577 21255 14633 21311
rect 14283 21174 14339 21230
rect 14381 21174 14437 21230
rect 14479 21174 14535 21230
rect 14577 21174 14633 21230
rect 242 21065 298 21121
rect 334 21065 390 21121
rect 426 21065 482 21121
rect 518 21065 574 21121
rect 610 21065 666 21121
rect 702 21065 758 21121
rect 242 20984 298 21040
rect 334 20984 390 21040
rect 426 20984 482 21040
rect 518 20984 574 21040
rect 610 20984 666 21040
rect 702 20984 758 21040
rect 242 20903 298 20959
rect 334 20903 390 20959
rect 426 20903 482 20959
rect 518 20903 574 20959
rect 610 20903 666 20959
rect 702 20903 758 20959
rect 242 20822 298 20878
rect 334 20822 390 20878
rect 426 20822 482 20878
rect 518 20822 574 20878
rect 610 20822 666 20878
rect 702 20822 758 20878
rect 242 20741 298 20797
rect 334 20741 390 20797
rect 426 20741 482 20797
rect 518 20741 574 20797
rect 610 20741 666 20797
rect 702 20741 758 20797
rect 242 20660 298 20716
rect 334 20660 390 20716
rect 426 20660 482 20716
rect 518 20660 574 20716
rect 610 20660 666 20716
rect 702 20660 758 20716
rect 242 20579 298 20635
rect 334 20579 390 20635
rect 426 20579 482 20635
rect 518 20579 574 20635
rect 610 20579 666 20635
rect 702 20579 758 20635
rect 242 20498 298 20554
rect 334 20498 390 20554
rect 426 20498 482 20554
rect 518 20498 574 20554
rect 610 20498 666 20554
rect 702 20498 758 20554
rect 14283 21093 14339 21149
rect 14381 21093 14437 21149
rect 14479 21093 14535 21149
rect 14577 21093 14633 21149
rect 14283 21012 14339 21068
rect 14381 21012 14437 21068
rect 14479 21012 14535 21068
rect 14577 21012 14633 21068
rect 14283 20931 14339 20987
rect 14381 20931 14437 20987
rect 14479 20931 14535 20987
rect 14577 20931 14633 20987
rect 14283 20850 14339 20906
rect 14381 20850 14437 20906
rect 14479 20850 14535 20906
rect 14577 20850 14633 20906
rect 14283 20769 14339 20825
rect 14381 20769 14437 20825
rect 14479 20769 14535 20825
rect 14577 20769 14633 20825
rect 14283 20688 14339 20744
rect 14381 20688 14437 20744
rect 14479 20688 14535 20744
rect 14577 20688 14633 20744
rect 14283 20607 14339 20663
rect 14381 20607 14437 20663
rect 14479 20607 14535 20663
rect 14577 20607 14633 20663
rect 14283 20526 14339 20582
rect 14381 20526 14437 20582
rect 14479 20526 14535 20582
rect 14577 20526 14633 20582
rect 242 20417 298 20473
rect 334 20417 390 20473
rect 426 20417 482 20473
rect 518 20417 574 20473
rect 610 20417 666 20473
rect 702 20417 758 20473
rect 203 8785 259 8841
rect 287 8785 343 8841
rect 371 8785 427 8841
rect 454 8785 510 8841
rect 537 8785 593 8841
rect 620 8785 676 8841
rect 703 8785 759 8841
rect 786 8785 842 8841
rect 869 8785 925 8841
rect 952 8785 1008 8841
rect 1035 8785 1091 8841
rect 1118 8785 1174 8841
rect 1201 8785 1257 8841
rect 203 8699 259 8755
rect 287 8699 343 8755
rect 371 8699 427 8755
rect 454 8699 510 8755
rect 537 8699 593 8755
rect 620 8699 676 8755
rect 703 8699 759 8755
rect 786 8699 842 8755
rect 869 8699 925 8755
rect 952 8699 1008 8755
rect 1035 8699 1091 8755
rect 1118 8699 1174 8755
rect 1201 8699 1257 8755
rect 203 8613 259 8669
rect 287 8613 343 8669
rect 371 8613 427 8669
rect 454 8613 510 8669
rect 537 8613 593 8669
rect 620 8613 676 8669
rect 703 8613 759 8669
rect 786 8613 842 8669
rect 869 8613 925 8669
rect 952 8613 1008 8669
rect 1035 8613 1091 8669
rect 1118 8613 1174 8669
rect 1201 8613 1257 8669
rect 203 8527 259 8583
rect 287 8527 343 8583
rect 371 8527 427 8583
rect 454 8527 510 8583
rect 537 8527 593 8583
rect 620 8527 676 8583
rect 703 8527 759 8583
rect 786 8527 842 8583
rect 869 8527 925 8583
rect 952 8527 1008 8583
rect 1035 8527 1091 8583
rect 1118 8527 1174 8583
rect 1201 8527 1257 8583
rect 203 8441 259 8497
rect 287 8441 343 8497
rect 371 8441 427 8497
rect 454 8441 510 8497
rect 537 8441 593 8497
rect 620 8441 676 8497
rect 703 8441 759 8497
rect 786 8441 842 8497
rect 869 8441 925 8497
rect 952 8441 1008 8497
rect 1035 8441 1091 8497
rect 1118 8441 1174 8497
rect 1201 8441 1257 8497
rect 203 8355 259 8411
rect 287 8355 343 8411
rect 371 8355 427 8411
rect 454 8355 510 8411
rect 537 8355 593 8411
rect 620 8355 676 8411
rect 703 8355 759 8411
rect 786 8355 842 8411
rect 869 8355 925 8411
rect 952 8355 1008 8411
rect 1035 8355 1091 8411
rect 1118 8355 1174 8411
rect 1201 8355 1257 8411
rect 203 8269 259 8325
rect 287 8269 343 8325
rect 371 8269 427 8325
rect 454 8269 510 8325
rect 537 8269 593 8325
rect 620 8269 676 8325
rect 703 8269 759 8325
rect 786 8269 842 8325
rect 869 8269 925 8325
rect 952 8269 1008 8325
rect 1035 8269 1091 8325
rect 1118 8269 1174 8325
rect 1201 8269 1257 8325
rect 203 8183 259 8239
rect 287 8183 343 8239
rect 371 8183 427 8239
rect 454 8183 510 8239
rect 537 8183 593 8239
rect 620 8183 676 8239
rect 703 8183 759 8239
rect 786 8183 842 8239
rect 869 8183 925 8239
rect 952 8183 1008 8239
rect 1035 8183 1091 8239
rect 1118 8183 1174 8239
rect 1201 8183 1257 8239
rect 203 8097 259 8153
rect 287 8097 343 8153
rect 371 8097 427 8153
rect 454 8097 510 8153
rect 537 8097 593 8153
rect 620 8097 676 8153
rect 703 8097 759 8153
rect 786 8097 842 8153
rect 869 8097 925 8153
rect 952 8097 1008 8153
rect 1035 8097 1091 8153
rect 1118 8097 1174 8153
rect 1201 8097 1257 8153
rect 203 8011 259 8067
rect 287 8011 343 8067
rect 371 8011 427 8067
rect 454 8011 510 8067
rect 537 8011 593 8067
rect 620 8011 676 8067
rect 703 8011 759 8067
rect 786 8011 842 8067
rect 869 8011 925 8067
rect 952 8011 1008 8067
rect 1035 8011 1091 8067
rect 1118 8011 1174 8067
rect 1201 8011 1257 8067
rect 203 7925 259 7981
rect 287 7925 343 7981
rect 371 7925 427 7981
rect 454 7925 510 7981
rect 537 7925 593 7981
rect 620 7925 676 7981
rect 703 7925 759 7981
rect 786 7925 842 7981
rect 869 7925 925 7981
rect 952 7925 1008 7981
rect 1035 7925 1091 7981
rect 1118 7925 1174 7981
rect 1201 7925 1257 7981
rect 8203 8785 8259 8841
rect 8287 8785 8343 8841
rect 8370 8785 8426 8841
rect 8453 8785 8509 8841
rect 8536 8785 8592 8841
rect 8619 8785 8675 8841
rect 8702 8785 8758 8841
rect 8785 8785 8841 8841
rect 8868 8785 8924 8841
rect 8951 8785 9007 8841
rect 9034 8785 9090 8841
rect 9117 8785 9173 8841
rect 9200 8785 9256 8841
rect 8203 8699 8259 8755
rect 8287 8699 8343 8755
rect 8370 8699 8426 8755
rect 8453 8699 8509 8755
rect 8536 8699 8592 8755
rect 8619 8699 8675 8755
rect 8702 8699 8758 8755
rect 8785 8699 8841 8755
rect 8868 8699 8924 8755
rect 8951 8699 9007 8755
rect 9034 8699 9090 8755
rect 9117 8699 9173 8755
rect 9200 8699 9256 8755
rect 8203 8613 8259 8669
rect 8287 8613 8343 8669
rect 8370 8613 8426 8669
rect 8453 8613 8509 8669
rect 8536 8613 8592 8669
rect 8619 8613 8675 8669
rect 8702 8613 8758 8669
rect 8785 8613 8841 8669
rect 8868 8613 8924 8669
rect 8951 8613 9007 8669
rect 9034 8613 9090 8669
rect 9117 8613 9173 8669
rect 9200 8613 9256 8669
rect 8203 8527 8259 8583
rect 8287 8527 8343 8583
rect 8370 8527 8426 8583
rect 8453 8527 8509 8583
rect 8536 8527 8592 8583
rect 8619 8527 8675 8583
rect 8702 8527 8758 8583
rect 8785 8527 8841 8583
rect 8868 8527 8924 8583
rect 8951 8527 9007 8583
rect 9034 8527 9090 8583
rect 9117 8527 9173 8583
rect 9200 8527 9256 8583
rect 8203 8441 8259 8497
rect 8287 8441 8343 8497
rect 8370 8441 8426 8497
rect 8453 8441 8509 8497
rect 8536 8441 8592 8497
rect 8619 8441 8675 8497
rect 8702 8441 8758 8497
rect 8785 8441 8841 8497
rect 8868 8441 8924 8497
rect 8951 8441 9007 8497
rect 9034 8441 9090 8497
rect 9117 8441 9173 8497
rect 9200 8441 9256 8497
rect 8203 8355 8259 8411
rect 8287 8355 8343 8411
rect 8370 8355 8426 8411
rect 8453 8355 8509 8411
rect 8536 8355 8592 8411
rect 8619 8355 8675 8411
rect 8702 8355 8758 8411
rect 8785 8355 8841 8411
rect 8868 8355 8924 8411
rect 8951 8355 9007 8411
rect 9034 8355 9090 8411
rect 9117 8355 9173 8411
rect 9200 8355 9256 8411
rect 8203 8269 8259 8325
rect 8287 8269 8343 8325
rect 8370 8269 8426 8325
rect 8453 8269 8509 8325
rect 8536 8269 8592 8325
rect 8619 8269 8675 8325
rect 8702 8269 8758 8325
rect 8785 8269 8841 8325
rect 8868 8269 8924 8325
rect 8951 8269 9007 8325
rect 9034 8269 9090 8325
rect 9117 8269 9173 8325
rect 9200 8269 9256 8325
rect 8203 8183 8259 8239
rect 8287 8183 8343 8239
rect 8370 8183 8426 8239
rect 8453 8183 8509 8239
rect 8536 8183 8592 8239
rect 8619 8183 8675 8239
rect 8702 8183 8758 8239
rect 8785 8183 8841 8239
rect 8868 8183 8924 8239
rect 8951 8183 9007 8239
rect 9034 8183 9090 8239
rect 9117 8183 9173 8239
rect 9200 8183 9256 8239
rect 8203 8097 8259 8153
rect 8287 8097 8343 8153
rect 8370 8097 8426 8153
rect 8453 8097 8509 8153
rect 8536 8097 8592 8153
rect 8619 8097 8675 8153
rect 8702 8097 8758 8153
rect 8785 8097 8841 8153
rect 8868 8097 8924 8153
rect 8951 8097 9007 8153
rect 9034 8097 9090 8153
rect 9117 8097 9173 8153
rect 9200 8097 9256 8153
rect 8203 8011 8259 8067
rect 8287 8011 8343 8067
rect 8370 8011 8426 8067
rect 8453 8011 8509 8067
rect 8536 8011 8592 8067
rect 8619 8011 8675 8067
rect 8702 8011 8758 8067
rect 8785 8011 8841 8067
rect 8868 8011 8924 8067
rect 8951 8011 9007 8067
rect 9034 8011 9090 8067
rect 9117 8011 9173 8067
rect 9200 8011 9256 8067
rect 8203 7925 8259 7981
rect 8287 7925 8343 7981
rect 8370 7925 8426 7981
rect 8453 7925 8509 7981
rect 8536 7925 8592 7981
rect 8619 7925 8675 7981
rect 8702 7925 8758 7981
rect 8785 7925 8841 7981
rect 8868 7925 8924 7981
rect 8951 7925 9007 7981
rect 9034 7925 9090 7981
rect 9117 7925 9173 7981
rect 9200 7925 9256 7981
<< metal3 >>
rect 460 39592 684 39600
rect 460 39528 462 39592
rect 526 39528 620 39592
rect 460 39512 684 39528
rect 460 39448 462 39512
rect 526 39448 620 39512
rect 460 39432 684 39448
rect 460 39368 462 39432
rect 526 39368 620 39432
rect 460 39352 684 39368
rect 460 39288 462 39352
rect 526 39288 620 39352
rect 460 39272 684 39288
rect 460 39208 462 39272
rect 526 39208 620 39272
rect 460 39192 684 39208
rect 460 39128 462 39192
rect 526 39128 620 39192
rect 460 39112 684 39128
rect 460 39048 462 39112
rect 526 39048 620 39112
rect 460 39032 684 39048
rect 460 38968 462 39032
rect 526 38968 620 39032
rect 460 38952 684 38968
rect 460 38888 462 38952
rect 526 38888 620 38952
rect 460 38872 684 38888
rect 460 38808 462 38872
rect 526 38808 620 38872
rect 460 38792 684 38808
rect 460 38728 462 38792
rect 526 38728 620 38792
rect 460 38712 684 38728
rect 460 38648 462 38712
rect 526 38648 620 38712
rect 460 38632 684 38648
rect 460 38568 462 38632
rect 526 38568 620 38632
rect 460 38552 684 38568
rect 460 38488 462 38552
rect 526 38488 620 38552
rect 460 38472 684 38488
rect 460 38408 462 38472
rect 526 38408 620 38472
rect 460 38392 684 38408
rect 460 38328 462 38392
rect 526 38328 620 38392
rect 460 38311 684 38328
rect 460 38247 462 38311
rect 526 38247 620 38311
rect 460 38230 684 38247
rect 460 38166 462 38230
rect 526 38166 620 38230
rect 460 38149 684 38166
rect 460 38085 462 38149
rect 526 38085 620 38149
rect 460 38068 684 38085
rect 460 38004 462 38068
rect 526 38004 620 38068
rect 460 37987 684 38004
rect 460 37923 462 37987
rect 526 37923 620 37987
rect 460 37906 684 37923
rect 460 37842 462 37906
rect 526 37842 620 37906
rect 460 37825 684 37842
rect 460 37761 462 37825
rect 526 37761 620 37825
rect 460 37744 684 37761
rect 460 37680 462 37744
rect 526 37680 620 37744
rect 460 37663 684 37680
rect 460 37599 462 37663
rect 526 37599 620 37663
rect 460 37582 684 37599
rect 460 37518 462 37582
rect 526 37518 620 37582
rect 460 37501 684 37518
rect 460 37437 462 37501
rect 526 37437 620 37501
rect 460 37420 684 37437
rect 460 37356 462 37420
rect 526 37356 620 37420
rect 460 37339 684 37356
rect 460 37275 462 37339
rect 526 37275 620 37339
rect 460 37258 684 37275
rect 460 37194 462 37258
rect 526 37194 620 37258
rect 460 37177 684 37194
rect 460 37113 462 37177
rect 526 37113 620 37177
rect 460 37096 684 37113
rect 460 37032 462 37096
rect 526 37032 620 37096
rect 460 37015 684 37032
rect 460 36951 462 37015
rect 526 36951 620 37015
rect 460 36934 684 36951
rect 460 36870 462 36934
rect 526 36870 620 36934
rect 460 36853 684 36870
rect 460 36789 462 36853
rect 526 36789 620 36853
rect 460 36772 684 36789
rect 460 36708 462 36772
rect 526 36708 620 36772
rect 460 36691 684 36708
rect 460 36627 462 36691
rect 526 36627 620 36691
rect 460 36610 684 36627
rect 460 36546 462 36610
rect 526 36546 620 36610
rect 460 36529 684 36546
rect 460 36465 462 36529
rect 526 36465 620 36529
rect 460 36448 684 36465
rect 460 36384 462 36448
rect 526 36384 620 36448
rect 460 36367 684 36384
rect 460 36303 462 36367
rect 526 36303 620 36367
rect 460 36286 684 36303
rect 460 36222 462 36286
rect 526 36222 620 36286
rect 460 36205 684 36222
rect 460 36141 462 36205
rect 526 36141 620 36205
rect 460 36124 684 36141
rect 460 36060 462 36124
rect 526 36060 620 36124
rect 460 36043 684 36060
rect 460 35979 462 36043
rect 526 35979 620 36043
rect 460 35962 684 35979
rect 460 35898 462 35962
rect 526 35898 620 35962
rect 460 35881 684 35898
rect 460 35817 462 35881
rect 526 35817 620 35881
rect 460 35800 684 35817
rect 460 35736 462 35800
rect 526 35736 620 35800
rect 460 35719 684 35736
rect 460 35655 462 35719
rect 526 35655 620 35719
rect 460 35638 684 35655
rect 460 35574 462 35638
rect 526 35574 620 35638
rect 460 35557 684 35574
rect 460 35493 462 35557
rect 526 35493 620 35557
rect 460 35476 684 35493
rect 460 35412 462 35476
rect 526 35412 620 35476
rect 460 35395 684 35412
rect 460 35331 462 35395
rect 526 35331 620 35395
rect 460 35314 684 35331
rect 460 35250 462 35314
rect 526 35250 620 35314
rect 460 35233 684 35250
rect 460 35169 462 35233
rect 526 35169 620 35233
rect 460 35152 684 35169
rect 460 35088 462 35152
rect 526 35088 620 35152
rect 460 35071 684 35088
rect 460 35007 462 35071
rect 526 35007 620 35071
rect 460 34990 684 35007
rect 460 34926 462 34990
rect 526 34926 620 34990
rect 460 34909 684 34926
rect 460 34845 462 34909
rect 526 34845 620 34909
rect 460 34828 684 34845
rect 460 34764 462 34828
rect 526 34764 620 34828
rect 460 32764 684 34764
rect 460 32708 465 32764
rect 521 32708 623 32764
rect 679 32708 684 32764
rect 460 32683 684 32708
rect 460 32627 465 32683
rect 521 32627 623 32683
rect 679 32627 684 32683
rect 460 32601 684 32627
rect 460 32545 465 32601
rect 521 32545 623 32601
rect 679 32545 684 32601
rect 460 32519 684 32545
rect 460 32463 465 32519
rect 521 32463 623 32519
rect 679 32463 684 32519
rect 460 32437 684 32463
rect 460 32381 465 32437
rect 521 32381 623 32437
rect 679 32381 684 32437
rect 460 32355 684 32381
rect 460 32299 465 32355
rect 521 32299 623 32355
rect 679 32299 684 32355
rect 460 32273 684 32299
rect 460 32217 465 32273
rect 521 32217 623 32273
rect 679 32217 684 32273
rect 460 32191 684 32217
rect 460 32135 465 32191
rect 521 32135 623 32191
rect 679 32135 684 32191
rect 460 32109 684 32135
rect 460 32053 465 32109
rect 521 32053 623 32109
rect 679 32053 684 32109
rect 460 32027 684 32053
rect 460 31971 465 32027
rect 521 31971 623 32027
rect 679 31971 684 32027
rect 1390 39592 1582 39600
rect 1454 39528 1518 39592
rect 1390 39512 1582 39528
rect 1454 39448 1518 39512
rect 1390 39432 1582 39448
rect 1454 39368 1518 39432
rect 1390 39352 1582 39368
rect 1454 39288 1518 39352
rect 1390 39272 1582 39288
rect 1454 39208 1518 39272
rect 1390 39192 1582 39208
rect 1454 39128 1518 39192
rect 1390 39112 1582 39128
rect 1454 39048 1518 39112
rect 1390 39032 1582 39048
rect 1454 38968 1518 39032
rect 1390 38952 1582 38968
rect 1454 38888 1518 38952
rect 1390 38872 1582 38888
rect 1454 38808 1518 38872
rect 1390 38792 1582 38808
rect 1454 38728 1518 38792
rect 1390 38712 1582 38728
rect 1454 38648 1518 38712
rect 1390 38632 1582 38648
rect 1454 38568 1518 38632
rect 1390 38552 1582 38568
rect 1454 38488 1518 38552
rect 1390 38472 1582 38488
rect 1454 38408 1518 38472
rect 1390 38392 1582 38408
rect 1454 38328 1518 38392
rect 1390 38311 1582 38328
rect 1454 38247 1518 38311
rect 1390 38230 1582 38247
rect 1454 38166 1518 38230
rect 1390 38149 1582 38166
rect 1454 38085 1518 38149
rect 1390 38068 1582 38085
rect 1454 38004 1518 38068
rect 1390 37987 1582 38004
rect 1454 37923 1518 37987
rect 1390 37906 1582 37923
rect 1454 37842 1518 37906
rect 1390 37825 1582 37842
rect 1454 37761 1518 37825
rect 1390 37744 1582 37761
rect 1454 37680 1518 37744
rect 1390 37663 1582 37680
rect 1454 37599 1518 37663
rect 1390 37582 1582 37599
rect 1454 37518 1518 37582
rect 1390 37501 1582 37518
rect 1454 37437 1518 37501
rect 1390 37420 1582 37437
rect 1454 37356 1518 37420
rect 1390 37339 1582 37356
rect 1454 37275 1518 37339
rect 1390 37258 1582 37275
rect 1454 37194 1518 37258
rect 1390 37177 1582 37194
rect 1454 37113 1518 37177
rect 1390 37096 1582 37113
rect 1454 37032 1518 37096
rect 1390 37015 1582 37032
rect 1454 36951 1518 37015
rect 1390 36934 1582 36951
rect 1454 36870 1518 36934
rect 1390 36853 1582 36870
rect 1454 36789 1518 36853
rect 1390 36772 1582 36789
rect 1454 36708 1518 36772
rect 1390 36691 1582 36708
rect 1454 36627 1518 36691
rect 1390 36610 1582 36627
rect 1454 36546 1518 36610
rect 1390 36529 1582 36546
rect 1454 36465 1518 36529
rect 1390 36448 1582 36465
rect 1454 36384 1518 36448
rect 1390 36367 1582 36384
rect 1454 36303 1518 36367
rect 1390 36286 1582 36303
rect 1454 36222 1518 36286
rect 1390 36205 1582 36222
rect 1454 36141 1518 36205
rect 1390 36124 1582 36141
rect 1454 36060 1518 36124
rect 1390 36043 1582 36060
rect 1454 35979 1518 36043
rect 1390 35962 1582 35979
rect 1454 35898 1518 35962
rect 1390 35881 1582 35898
rect 1454 35817 1518 35881
rect 1390 35800 1582 35817
rect 1454 35736 1518 35800
rect 1390 35719 1582 35736
rect 1454 35655 1518 35719
rect 1390 35638 1582 35655
rect 1454 35574 1518 35638
rect 1390 35557 1582 35574
rect 1454 35493 1518 35557
rect 1390 35476 1582 35493
rect 1454 35412 1518 35476
rect 1390 35395 1582 35412
rect 1454 35331 1518 35395
rect 1390 35314 1582 35331
rect 1454 35250 1518 35314
rect 1390 35233 1582 35250
rect 1454 35169 1518 35233
rect 1390 35152 1582 35169
rect 1454 35088 1518 35152
rect 1390 35071 1582 35088
rect 1454 35007 1518 35071
rect 1390 34990 1582 35007
rect 1454 34926 1518 34990
rect 1390 34909 1582 34926
rect 1454 34845 1518 34909
rect 1390 34828 1582 34845
rect 1454 34764 1518 34828
rect 460 31945 684 31971
rect 460 31889 465 31945
rect 521 31889 623 31945
rect 679 31889 684 31945
rect 460 31863 684 31889
rect 460 31807 465 31863
rect 521 31807 623 31863
rect 679 31807 684 31863
rect 460 31781 684 31807
rect 460 31725 465 31781
rect 521 31725 623 31781
rect 679 31725 684 31781
rect 460 31699 684 31725
rect 460 31643 465 31699
rect 521 31643 623 31699
rect 679 31643 684 31699
rect 460 31617 684 31643
rect 460 31561 465 31617
rect 521 31561 623 31617
rect 679 31561 684 31617
rect 460 31535 684 31561
rect 460 31479 465 31535
rect 521 31479 623 31535
rect 679 31479 684 31535
rect 460 31453 684 31479
rect 460 31397 465 31453
rect 521 31397 623 31453
rect 679 31397 684 31453
rect 460 31371 684 31397
rect 460 31315 465 31371
rect 521 31315 623 31371
rect 679 31315 684 31371
rect 460 31289 684 31315
rect 460 31233 465 31289
rect 521 31233 623 31289
rect 679 31233 684 31289
rect 460 31207 684 31233
rect 460 31151 465 31207
rect 521 31151 623 31207
rect 679 31151 684 31207
rect 460 31125 684 31151
rect 460 31069 465 31125
rect 521 31069 623 31125
rect 679 31069 684 31125
rect 460 31043 684 31069
rect 460 30987 465 31043
rect 521 30987 623 31043
rect 679 30987 684 31043
rect 460 30961 684 30987
rect 460 30905 465 30961
rect 521 30905 623 30961
rect 679 30905 684 30961
rect 460 30879 684 30905
rect 460 30823 465 30879
rect 521 30823 623 30879
rect 679 30823 684 30879
rect 460 30797 684 30823
rect 460 30741 465 30797
rect 521 30741 623 30797
rect 679 30741 684 30797
rect 460 30715 684 30741
rect 460 30659 465 30715
rect 521 30659 623 30715
rect 679 30659 684 30715
rect 460 30633 684 30659
rect 460 30577 465 30633
rect 521 30577 623 30633
rect 679 30577 684 30633
rect 460 30551 684 30577
rect 460 30495 465 30551
rect 521 30495 623 30551
rect 679 30495 684 30551
rect 460 30469 684 30495
rect 460 30413 465 30469
rect 521 30413 623 30469
rect 679 30413 684 30469
rect 460 30387 684 30413
rect 460 30331 465 30387
rect 521 30331 623 30387
rect 679 30331 684 30387
rect 460 30305 684 30331
rect 460 30249 465 30305
rect 521 30249 623 30305
rect 679 30249 684 30305
rect 460 30223 684 30249
rect 460 30167 465 30223
rect 521 30167 623 30223
rect 679 30167 684 30223
rect 460 30141 684 30167
rect 460 30085 465 30141
rect 521 30085 623 30141
rect 679 30085 684 30141
rect 460 30059 684 30085
rect 460 30003 465 30059
rect 521 30003 623 30059
rect 679 30003 684 30059
rect 460 29977 684 30003
rect 460 29921 465 29977
rect 521 29921 623 29977
rect 679 29921 684 29977
rect 460 29895 684 29921
rect 460 29839 465 29895
rect 521 29839 623 29895
rect 679 29839 684 29895
rect 460 29813 684 29839
rect 460 29757 465 29813
rect 521 29757 623 29813
rect 679 29757 684 29813
rect 460 29731 684 29757
rect 460 29675 465 29731
rect 521 29675 623 29731
rect 679 29675 684 29731
rect 460 29649 684 29675
rect 460 29593 465 29649
rect 521 29593 623 29649
rect 679 29593 684 29649
rect 460 29567 684 29593
rect 460 29511 465 29567
rect 521 29511 623 29567
rect 679 29511 684 29567
rect 460 29485 684 29511
rect 460 29429 465 29485
rect 521 29429 623 29485
rect 679 29429 684 29485
rect 460 29424 684 29429
rect 857 32018 1057 32023
rect 857 31953 862 32018
rect 918 32017 996 32018
rect 1052 32017 1057 32018
rect 926 31953 990 32017
rect 1054 31953 1057 32017
rect 857 31936 1057 31953
rect 857 31872 862 31936
rect 926 31872 990 31936
rect 1054 31872 1057 31936
rect 857 31855 1057 31872
rect 857 31791 862 31855
rect 926 31791 990 31855
rect 1054 31791 1057 31855
rect 857 31774 1057 31791
rect 857 31710 862 31774
rect 926 31710 990 31774
rect 1054 31710 1057 31774
rect 857 31693 1057 31710
rect 857 31629 862 31693
rect 926 31629 990 31693
rect 1054 31629 1057 31693
rect 857 31612 1057 31629
rect 857 31548 862 31612
rect 926 31548 990 31612
rect 1054 31548 1057 31612
rect 857 31531 1057 31548
rect 857 31467 862 31531
rect 926 31467 990 31531
rect 1054 31467 1057 31531
rect 857 31450 1057 31467
rect 857 31386 862 31450
rect 926 31386 990 31450
rect 1054 31386 1057 31450
rect 857 31369 1057 31386
rect 857 31305 862 31369
rect 926 31305 990 31369
rect 1054 31305 1057 31369
rect 857 31288 1057 31305
rect 857 31224 862 31288
rect 926 31224 990 31288
rect 1054 31224 1057 31288
rect 857 31207 1057 31224
rect 857 31142 862 31207
rect 926 31143 990 31207
rect 1054 31143 1057 31207
rect 918 31142 996 31143
rect 1052 31142 1057 31143
rect 857 31125 1057 31142
rect 857 31060 862 31125
rect 926 31061 990 31125
rect 1054 31061 1057 31125
rect 918 31060 996 31061
rect 1052 31060 1057 31061
rect 857 31043 1057 31060
rect 857 30978 862 31043
rect 926 30979 990 31043
rect 1054 30979 1057 31043
rect 918 30978 996 30979
rect 1052 30978 1057 30979
rect 857 30961 1057 30978
rect 857 30896 862 30961
rect 926 30897 990 30961
rect 1054 30897 1057 30961
rect 918 30896 996 30897
rect 1052 30896 1057 30897
rect 857 30879 1057 30896
rect 857 30814 862 30879
rect 926 30815 990 30879
rect 1054 30815 1057 30879
rect 918 30814 996 30815
rect 1052 30814 1057 30815
rect 857 30797 1057 30814
rect 857 30732 862 30797
rect 926 30733 990 30797
rect 1054 30733 1057 30797
rect 918 30732 996 30733
rect 1052 30732 1057 30733
rect 857 30715 1057 30732
rect 857 30650 862 30715
rect 926 30651 990 30715
rect 1054 30651 1057 30715
rect 918 30650 996 30651
rect 1052 30650 1057 30651
rect 857 30633 1057 30650
rect 857 30568 862 30633
rect 926 30569 990 30633
rect 1054 30569 1057 30633
rect 918 30568 996 30569
rect 1052 30568 1057 30569
rect 857 30551 1057 30568
rect 857 30486 862 30551
rect 926 30487 990 30551
rect 1054 30487 1057 30551
rect 918 30486 996 30487
rect 1052 30486 1057 30487
rect 857 30469 1057 30486
rect 857 30404 862 30469
rect 926 30405 990 30469
rect 1054 30405 1057 30469
rect 918 30404 996 30405
rect 1052 30404 1057 30405
rect 857 30387 1057 30404
rect 857 30322 862 30387
rect 926 30323 990 30387
rect 1054 30323 1057 30387
rect 918 30322 996 30323
rect 1052 30322 1057 30323
rect 857 30305 1057 30322
rect 857 30240 862 30305
rect 926 30241 990 30305
rect 1054 30241 1057 30305
rect 918 30240 996 30241
rect 1052 30240 1057 30241
rect 857 30223 1057 30240
rect 857 30158 862 30223
rect 926 30159 990 30223
rect 1054 30159 1057 30223
rect 918 30158 996 30159
rect 1052 30158 1057 30159
rect 857 30141 1057 30158
rect 857 30076 862 30141
rect 926 30077 990 30141
rect 1054 30077 1057 30141
rect 918 30076 996 30077
rect 1052 30076 1057 30077
rect 857 30059 1057 30076
rect 857 29994 862 30059
rect 926 29995 990 30059
rect 1054 29995 1057 30059
rect 918 29994 996 29995
rect 1052 29994 1057 29995
rect 857 29977 1057 29994
rect 857 29912 862 29977
rect 926 29913 990 29977
rect 1054 29913 1057 29977
rect 918 29912 996 29913
rect 1052 29912 1057 29913
rect 857 29895 1057 29912
rect 857 29830 862 29895
rect 926 29831 990 29895
rect 1054 29831 1057 29895
rect 918 29830 996 29831
rect 1052 29830 1057 29831
rect 857 29813 1057 29830
rect 857 29748 862 29813
rect 926 29749 990 29813
rect 1054 29749 1057 29813
rect 918 29748 996 29749
rect 1052 29748 1057 29749
rect 857 29731 1057 29748
rect 857 29666 862 29731
rect 926 29667 990 29731
rect 1054 29667 1057 29731
rect 918 29666 996 29667
rect 1052 29666 1057 29667
rect 857 29649 1057 29666
rect 857 29584 862 29649
rect 926 29585 990 29649
rect 1054 29585 1057 29649
rect 918 29584 996 29585
rect 1052 29584 1057 29585
rect 857 29567 1057 29584
rect 857 29502 862 29567
rect 926 29503 990 29567
rect 1054 29503 1057 29567
rect 918 29502 996 29503
rect 1052 29502 1057 29503
rect 857 29485 1057 29502
rect 857 29420 862 29485
rect 926 29421 990 29485
rect 1054 29421 1057 29485
rect 1390 32018 1582 34764
rect 2382 39592 2574 39600
rect 2446 39528 2510 39592
rect 2382 39512 2574 39528
rect 2446 39448 2510 39512
rect 2382 39432 2574 39448
rect 2446 39368 2510 39432
rect 2382 39352 2574 39368
rect 2446 39288 2510 39352
rect 2382 39272 2574 39288
rect 2446 39208 2510 39272
rect 2382 39192 2574 39208
rect 2446 39128 2510 39192
rect 2382 39112 2574 39128
rect 2446 39048 2510 39112
rect 2382 39032 2574 39048
rect 2446 38968 2510 39032
rect 2382 38952 2574 38968
rect 2446 38888 2510 38952
rect 2382 38872 2574 38888
rect 2446 38808 2510 38872
rect 2382 38792 2574 38808
rect 2446 38728 2510 38792
rect 2382 38712 2574 38728
rect 2446 38648 2510 38712
rect 2382 38632 2574 38648
rect 2446 38568 2510 38632
rect 2382 38552 2574 38568
rect 2446 38488 2510 38552
rect 2382 38472 2574 38488
rect 2446 38408 2510 38472
rect 2382 38392 2574 38408
rect 2446 38328 2510 38392
rect 2382 38311 2574 38328
rect 2446 38247 2510 38311
rect 2382 38230 2574 38247
rect 2446 38166 2510 38230
rect 2382 38149 2574 38166
rect 2446 38085 2510 38149
rect 2382 38068 2574 38085
rect 2446 38004 2510 38068
rect 2382 37987 2574 38004
rect 2446 37923 2510 37987
rect 2382 37906 2574 37923
rect 2446 37842 2510 37906
rect 2382 37825 2574 37842
rect 2446 37761 2510 37825
rect 2382 37744 2574 37761
rect 2446 37680 2510 37744
rect 2382 37663 2574 37680
rect 2446 37599 2510 37663
rect 2382 37582 2574 37599
rect 2446 37518 2510 37582
rect 2382 37501 2574 37518
rect 2446 37437 2510 37501
rect 2382 37420 2574 37437
rect 2446 37356 2510 37420
rect 2382 37339 2574 37356
rect 2446 37275 2510 37339
rect 2382 37258 2574 37275
rect 2446 37194 2510 37258
rect 2382 37177 2574 37194
rect 2446 37113 2510 37177
rect 2382 37096 2574 37113
rect 2446 37032 2510 37096
rect 2382 37015 2574 37032
rect 2446 36951 2510 37015
rect 2382 36934 2574 36951
rect 2446 36870 2510 36934
rect 2382 36853 2574 36870
rect 2446 36789 2510 36853
rect 2382 36772 2574 36789
rect 2446 36708 2510 36772
rect 2382 36691 2574 36708
rect 2446 36627 2510 36691
rect 2382 36610 2574 36627
rect 2446 36546 2510 36610
rect 2382 36529 2574 36546
rect 2446 36465 2510 36529
rect 2382 36448 2574 36465
rect 2446 36384 2510 36448
rect 2382 36367 2574 36384
rect 2446 36303 2510 36367
rect 2382 36286 2574 36303
rect 2446 36222 2510 36286
rect 2382 36205 2574 36222
rect 2446 36141 2510 36205
rect 2382 36124 2574 36141
rect 2446 36060 2510 36124
rect 2382 36043 2574 36060
rect 2446 35979 2510 36043
rect 2382 35962 2574 35979
rect 2446 35898 2510 35962
rect 2382 35881 2574 35898
rect 2446 35817 2510 35881
rect 2382 35800 2574 35817
rect 2446 35736 2510 35800
rect 2382 35719 2574 35736
rect 2446 35655 2510 35719
rect 2382 35638 2574 35655
rect 2446 35574 2510 35638
rect 2382 35557 2574 35574
rect 2446 35493 2510 35557
rect 2382 35476 2574 35493
rect 2446 35412 2510 35476
rect 2382 35395 2574 35412
rect 2446 35331 2510 35395
rect 2382 35314 2574 35331
rect 2446 35250 2510 35314
rect 2382 35233 2574 35250
rect 2446 35169 2510 35233
rect 2382 35152 2574 35169
rect 2446 35088 2510 35152
rect 2382 35071 2574 35088
rect 2446 35007 2510 35071
rect 2382 34990 2574 35007
rect 2446 34926 2510 34990
rect 2382 34909 2574 34926
rect 2446 34845 2510 34909
rect 2382 34828 2574 34845
rect 2446 34764 2510 34828
rect 1390 31962 1395 32018
rect 1451 31962 1521 32018
rect 1577 31962 1582 32018
rect 1390 31937 1582 31962
rect 1390 31881 1395 31937
rect 1451 31881 1521 31937
rect 1577 31881 1582 31937
rect 1390 31856 1582 31881
rect 1390 31800 1395 31856
rect 1451 31800 1521 31856
rect 1577 31800 1582 31856
rect 1390 31775 1582 31800
rect 1390 31719 1395 31775
rect 1451 31719 1521 31775
rect 1577 31719 1582 31775
rect 1390 31694 1582 31719
rect 1390 31638 1395 31694
rect 1451 31638 1521 31694
rect 1577 31638 1582 31694
rect 1390 31613 1582 31638
rect 1390 31557 1395 31613
rect 1451 31557 1521 31613
rect 1577 31557 1582 31613
rect 1390 31532 1582 31557
rect 1390 31476 1395 31532
rect 1451 31476 1521 31532
rect 1577 31476 1582 31532
rect 1390 31451 1582 31476
rect 1390 31395 1395 31451
rect 1451 31395 1521 31451
rect 1577 31395 1582 31451
rect 1390 31370 1582 31395
rect 1390 31314 1395 31370
rect 1451 31314 1521 31370
rect 1577 31314 1582 31370
rect 1390 31289 1582 31314
rect 1390 31233 1395 31289
rect 1451 31233 1521 31289
rect 1577 31233 1582 31289
rect 1390 31207 1582 31233
rect 1390 31151 1395 31207
rect 1451 31151 1521 31207
rect 1577 31151 1582 31207
rect 1390 31125 1582 31151
rect 1390 31069 1395 31125
rect 1451 31069 1521 31125
rect 1577 31069 1582 31125
rect 1390 31043 1582 31069
rect 1390 30987 1395 31043
rect 1451 30987 1521 31043
rect 1577 30987 1582 31043
rect 1390 30961 1582 30987
rect 1390 30905 1395 30961
rect 1451 30905 1521 30961
rect 1577 30905 1582 30961
rect 1390 30879 1582 30905
rect 1390 30823 1395 30879
rect 1451 30823 1521 30879
rect 1577 30823 1582 30879
rect 1390 30797 1582 30823
rect 1390 30741 1395 30797
rect 1451 30741 1521 30797
rect 1577 30741 1582 30797
rect 1390 30715 1582 30741
rect 1390 30659 1395 30715
rect 1451 30659 1521 30715
rect 1577 30659 1582 30715
rect 1390 30633 1582 30659
rect 1390 30577 1395 30633
rect 1451 30577 1521 30633
rect 1577 30577 1582 30633
rect 1390 30551 1582 30577
rect 1390 30495 1395 30551
rect 1451 30495 1521 30551
rect 1577 30495 1582 30551
rect 1390 30469 1582 30495
rect 1390 30413 1395 30469
rect 1451 30413 1521 30469
rect 1577 30413 1582 30469
rect 1390 30387 1582 30413
rect 1390 30331 1395 30387
rect 1451 30331 1521 30387
rect 1577 30331 1582 30387
rect 1390 30305 1582 30331
rect 1390 30249 1395 30305
rect 1451 30249 1521 30305
rect 1577 30249 1582 30305
rect 1390 30223 1582 30249
rect 1390 30167 1395 30223
rect 1451 30167 1521 30223
rect 1577 30167 1582 30223
rect 1390 30141 1582 30167
rect 1390 30085 1395 30141
rect 1451 30085 1521 30141
rect 1577 30085 1582 30141
rect 1390 30059 1582 30085
rect 1390 30003 1395 30059
rect 1451 30003 1521 30059
rect 1577 30003 1582 30059
rect 1390 29977 1582 30003
rect 1390 29921 1395 29977
rect 1451 29921 1521 29977
rect 1577 29921 1582 29977
rect 1390 29895 1582 29921
rect 1390 29839 1395 29895
rect 1451 29839 1521 29895
rect 1577 29839 1582 29895
rect 1390 29813 1582 29839
rect 1390 29757 1395 29813
rect 1451 29757 1521 29813
rect 1577 29757 1582 29813
rect 1390 29731 1582 29757
rect 1390 29675 1395 29731
rect 1451 29675 1521 29731
rect 1577 29675 1582 29731
rect 1390 29649 1582 29675
rect 1390 29593 1395 29649
rect 1451 29593 1521 29649
rect 1577 29593 1582 29649
rect 1390 29567 1582 29593
rect 1390 29511 1395 29567
rect 1451 29511 1521 29567
rect 1577 29511 1582 29567
rect 1390 29485 1582 29511
rect 1390 29429 1395 29485
rect 1451 29429 1521 29485
rect 1577 29429 1582 29485
rect 1390 29424 1582 29429
rect 1886 33831 2078 33844
rect 1950 33767 2014 33831
rect 1886 33749 2078 33767
rect 1950 33685 2014 33749
rect 1886 33666 2078 33685
rect 1950 33602 2014 33666
rect 1886 33583 2078 33602
rect 1950 33519 2014 33583
rect 1886 33500 2078 33519
rect 1950 33436 2014 33500
rect 1886 33417 2078 33436
rect 1950 33353 2014 33417
rect 1886 33334 2078 33353
rect 1950 33270 2014 33334
rect 1886 32018 2078 33270
rect 1886 31962 1891 32018
rect 1947 31962 2017 32018
rect 2073 31962 2078 32018
rect 1886 31936 2078 31962
rect 1886 31880 1891 31936
rect 1947 31880 2017 31936
rect 2073 31880 2078 31936
rect 1886 31854 2078 31880
rect 1886 31798 1891 31854
rect 1947 31798 2017 31854
rect 2073 31798 2078 31854
rect 1886 31772 2078 31798
rect 1886 31716 1891 31772
rect 1947 31716 2017 31772
rect 2073 31716 2078 31772
rect 1886 31690 2078 31716
rect 1886 31634 1891 31690
rect 1947 31634 2017 31690
rect 2073 31634 2078 31690
rect 1886 31608 2078 31634
rect 1886 31552 1891 31608
rect 1947 31552 2017 31608
rect 2073 31552 2078 31608
rect 1886 31526 2078 31552
rect 1886 31470 1891 31526
rect 1947 31470 2017 31526
rect 2073 31470 2078 31526
rect 1886 31444 2078 31470
rect 1886 31388 1891 31444
rect 1947 31388 2017 31444
rect 2073 31388 2078 31444
rect 1886 31362 2078 31388
rect 1886 31306 1891 31362
rect 1947 31306 2017 31362
rect 2073 31306 2078 31362
rect 1886 31280 2078 31306
rect 1886 31224 1891 31280
rect 1947 31224 2017 31280
rect 2073 31224 2078 31280
rect 1886 31198 2078 31224
rect 1886 31142 1891 31198
rect 1947 31142 2017 31198
rect 2073 31142 2078 31198
rect 1886 31116 2078 31142
rect 1886 31060 1891 31116
rect 1947 31060 2017 31116
rect 2073 31060 2078 31116
rect 1886 31034 2078 31060
rect 1886 30978 1891 31034
rect 1947 30978 2017 31034
rect 2073 30978 2078 31034
rect 1886 30952 2078 30978
rect 1886 30896 1891 30952
rect 1947 30896 2017 30952
rect 2073 30896 2078 30952
rect 1886 30870 2078 30896
rect 1886 30814 1891 30870
rect 1947 30814 2017 30870
rect 2073 30814 2078 30870
rect 1886 30788 2078 30814
rect 1886 30732 1891 30788
rect 1947 30732 2017 30788
rect 2073 30732 2078 30788
rect 1886 30706 2078 30732
rect 1886 30650 1891 30706
rect 1947 30650 2017 30706
rect 2073 30650 2078 30706
rect 1886 30624 2078 30650
rect 1886 30568 1891 30624
rect 1947 30568 2017 30624
rect 2073 30568 2078 30624
rect 1886 30542 2078 30568
rect 1886 30486 1891 30542
rect 1947 30486 2017 30542
rect 2073 30486 2078 30542
rect 1886 30460 2078 30486
rect 1886 30404 1891 30460
rect 1947 30404 2017 30460
rect 2073 30404 2078 30460
rect 1886 30378 2078 30404
rect 1886 30322 1891 30378
rect 1947 30322 2017 30378
rect 2073 30322 2078 30378
rect 1886 30296 2078 30322
rect 1886 30240 1891 30296
rect 1947 30240 2017 30296
rect 2073 30240 2078 30296
rect 1886 30214 2078 30240
rect 1886 30158 1891 30214
rect 1947 30158 2017 30214
rect 2073 30158 2078 30214
rect 1886 30132 2078 30158
rect 1886 30076 1891 30132
rect 1947 30076 2017 30132
rect 2073 30076 2078 30132
rect 1886 30050 2078 30076
rect 1886 29994 1891 30050
rect 1947 29994 2017 30050
rect 2073 29994 2078 30050
rect 1886 29968 2078 29994
rect 1886 29912 1891 29968
rect 1947 29912 2017 29968
rect 2073 29912 2078 29968
rect 1886 29886 2078 29912
rect 1886 29830 1891 29886
rect 1947 29830 2017 29886
rect 2073 29830 2078 29886
rect 1886 29804 2078 29830
rect 1886 29748 1891 29804
rect 1947 29748 2017 29804
rect 2073 29748 2078 29804
rect 1886 29722 2078 29748
rect 1886 29666 1891 29722
rect 1947 29666 2017 29722
rect 2073 29666 2078 29722
rect 1886 29640 2078 29666
rect 1886 29584 1891 29640
rect 1947 29584 2017 29640
rect 2073 29584 2078 29640
rect 1886 29558 2078 29584
rect 1886 29502 1891 29558
rect 1947 29502 2017 29558
rect 2073 29502 2078 29558
rect 1886 29476 2078 29502
rect 918 29420 996 29421
rect 1052 29420 1057 29421
rect 857 29415 1057 29420
rect 1886 29420 1891 29476
rect 1947 29420 2017 29476
rect 2073 29420 2078 29476
tri 1834 29238 1886 29290 se
rect 1886 29238 2078 29420
tri 1809 29213 1834 29238 se
rect 1834 29213 2078 29238
tri 1753 29157 1809 29213 se
rect 1809 29157 2078 29213
tri 1728 29132 1753 29157 se
rect 1753 29132 2078 29157
tri 1672 29076 1728 29132 se
rect 1728 29076 2078 29132
tri 1229 28633 1672 29076 se
rect 1672 28633 2078 29076
rect 219 28596 836 28633
tri 1216 28620 1229 28633 se
rect 1229 28620 2078 28633
rect 219 28540 579 28596
rect 635 28540 677 28596
rect 733 28540 775 28596
rect 831 28540 836 28596
tri 1160 28564 1216 28620 se
rect 1216 28564 2078 28620
rect 219 28515 836 28540
tri 1117 28521 1160 28564 se
rect 1160 28521 2078 28564
rect 219 28459 579 28515
rect 635 28459 677 28515
rect 733 28459 775 28515
rect 831 28459 836 28515
tri 1093 28497 1117 28521 se
rect 1117 28497 2078 28521
rect 219 28434 836 28459
tri 1049 28453 1093 28497 se
rect 1093 28453 2078 28497
tri 1047 28451 1049 28453 se
rect 1049 28451 2078 28453
rect 219 28378 579 28434
rect 635 28378 677 28434
rect 733 28378 775 28434
rect 831 28378 836 28434
tri 991 28395 1047 28451 se
rect 1047 28395 2078 28451
rect 219 28353 836 28378
rect 219 28297 579 28353
rect 635 28297 677 28353
rect 733 28297 775 28353
rect 831 28297 836 28353
rect 219 28272 836 28297
rect 219 28216 579 28272
rect 635 28216 677 28272
rect 733 28216 775 28272
rect 831 28216 836 28272
rect 219 28191 836 28216
rect 219 28135 579 28191
rect 635 28135 677 28191
rect 733 28135 775 28191
rect 831 28135 836 28191
rect 219 28110 836 28135
rect 219 28054 579 28110
rect 635 28054 677 28110
rect 733 28054 775 28110
rect 831 28054 836 28110
rect 219 28029 836 28054
rect 219 27973 579 28029
rect 635 27973 677 28029
rect 733 27973 775 28029
rect 831 27973 836 28029
rect 219 27948 836 27973
rect 219 27892 579 27948
rect 635 27892 677 27948
rect 733 27892 775 27948
rect 831 27892 836 27948
rect 219 27867 836 27892
rect 219 27811 579 27867
rect 635 27811 677 27867
rect 733 27811 775 27867
rect 831 27811 836 27867
rect 219 27786 836 27811
rect 219 27730 579 27786
rect 635 27730 677 27786
rect 733 27730 775 27786
rect 831 27730 836 27786
rect 219 27705 836 27730
rect 219 27649 579 27705
rect 635 27649 677 27705
rect 733 27649 775 27705
rect 831 27649 836 27705
rect 219 27624 836 27649
rect 219 27568 579 27624
rect 635 27568 677 27624
rect 733 27568 775 27624
rect 831 27568 836 27624
rect 219 27543 836 27568
rect 219 27487 579 27543
rect 635 27487 677 27543
rect 733 27487 775 27543
rect 831 27487 836 27543
rect 219 27462 836 27487
rect 219 27406 579 27462
rect 635 27406 677 27462
rect 733 27406 775 27462
rect 831 27406 836 27462
rect 219 27381 836 27406
rect 219 27325 579 27381
rect 635 27325 677 27381
rect 733 27325 775 27381
rect 831 27325 836 27381
rect 219 27300 836 27325
rect 219 27244 579 27300
rect 635 27244 677 27300
rect 733 27244 775 27300
rect 831 27244 836 27300
rect 219 27219 836 27244
rect 219 27163 579 27219
rect 635 27163 677 27219
rect 733 27163 775 27219
rect 831 27163 836 27219
rect 219 27138 836 27163
rect 219 27082 579 27138
rect 635 27082 677 27138
rect 733 27082 775 27138
rect 831 27082 836 27138
rect 219 27057 836 27082
rect 219 27001 579 27057
rect 635 27001 677 27057
rect 733 27001 775 27057
rect 831 27001 836 27057
rect 219 26976 836 27001
rect 219 26920 579 26976
rect 635 26920 677 26976
rect 733 26920 775 26976
rect 831 26920 836 26976
rect 219 26894 836 26920
rect 219 26838 579 26894
rect 635 26838 677 26894
rect 733 26838 775 26894
rect 831 26838 836 26894
rect 219 26812 836 26838
rect 219 26756 579 26812
rect 635 26756 677 26812
rect 733 26756 775 26812
rect 831 26756 836 26812
rect 219 26730 836 26756
rect 219 26674 579 26730
rect 635 26674 677 26730
rect 733 26674 775 26730
rect 831 26674 836 26730
rect 219 26648 836 26674
rect 219 26592 579 26648
rect 635 26592 677 26648
rect 733 26592 775 26648
rect 831 26592 836 26648
rect 219 26566 836 26592
rect 219 26510 579 26566
rect 635 26510 677 26566
rect 733 26510 775 26566
rect 831 26510 836 26566
rect 219 26484 836 26510
rect 219 26428 579 26484
rect 635 26428 677 26484
rect 733 26428 775 26484
rect 831 26428 836 26484
rect 219 26343 836 26428
rect 219 26287 242 26343
rect 298 26287 334 26343
rect 390 26287 426 26343
rect 482 26287 518 26343
rect 574 26287 610 26343
rect 666 26287 702 26343
rect 758 26287 836 26343
rect 219 26263 836 26287
rect 219 26207 242 26263
rect 298 26207 334 26263
rect 390 26207 426 26263
rect 482 26207 518 26263
rect 574 26207 610 26263
rect 666 26207 702 26263
rect 758 26207 836 26263
rect 219 26183 836 26207
rect 219 26127 242 26183
rect 298 26127 334 26183
rect 390 26127 426 26183
rect 482 26127 518 26183
rect 574 26127 610 26183
rect 666 26127 702 26183
rect 758 26127 836 26183
rect 219 26103 836 26127
rect 219 26047 242 26103
rect 298 26047 334 26103
rect 390 26047 426 26103
rect 482 26047 518 26103
rect 574 26047 610 26103
rect 666 26047 702 26103
rect 758 26047 836 26103
rect 219 26023 836 26047
rect 219 25967 242 26023
rect 298 25967 334 26023
rect 390 25967 426 26023
rect 482 25967 518 26023
rect 574 25967 610 26023
rect 666 25967 702 26023
rect 758 25967 836 26023
rect 219 25943 836 25967
rect 219 25887 242 25943
rect 298 25887 334 25943
rect 390 25887 426 25943
rect 482 25887 518 25943
rect 574 25887 610 25943
rect 666 25887 702 25943
rect 758 25887 836 25943
rect 219 25863 836 25887
rect 219 25807 242 25863
rect 298 25807 334 25863
rect 390 25807 426 25863
rect 482 25807 518 25863
rect 574 25807 610 25863
rect 666 25807 702 25863
rect 758 25807 836 25863
rect 219 25783 836 25807
rect 219 25727 242 25783
rect 298 25727 334 25783
rect 390 25727 426 25783
rect 482 25727 518 25783
rect 574 25727 610 25783
rect 666 25727 702 25783
rect 758 25727 836 25783
rect 219 25703 836 25727
rect 219 25647 242 25703
rect 298 25647 334 25703
rect 390 25647 426 25703
rect 482 25647 518 25703
rect 574 25647 610 25703
rect 666 25647 702 25703
rect 758 25647 836 25703
rect 219 25623 836 25647
rect 219 25567 242 25623
rect 298 25567 334 25623
rect 390 25567 426 25623
rect 482 25567 518 25623
rect 574 25567 610 25623
rect 666 25567 702 25623
rect 758 25567 836 25623
rect 219 25543 836 25567
rect 219 25487 242 25543
rect 298 25487 334 25543
rect 390 25487 426 25543
rect 482 25487 518 25543
rect 574 25487 610 25543
rect 666 25487 702 25543
rect 758 25487 836 25543
rect 219 25463 836 25487
rect 219 25407 242 25463
rect 298 25407 334 25463
rect 390 25407 426 25463
rect 482 25407 518 25463
rect 574 25407 610 25463
rect 666 25407 702 25463
rect 758 25407 836 25463
rect 219 25383 836 25407
rect 219 25327 242 25383
rect 298 25327 334 25383
rect 390 25327 426 25383
rect 482 25327 518 25383
rect 574 25327 610 25383
rect 666 25327 702 25383
rect 758 25327 836 25383
rect 219 25303 836 25327
rect 219 25247 242 25303
rect 298 25247 334 25303
rect 390 25247 426 25303
rect 482 25247 518 25303
rect 574 25247 610 25303
rect 666 25247 702 25303
rect 758 25247 836 25303
rect 219 25223 836 25247
rect 219 25167 242 25223
rect 298 25167 334 25223
rect 390 25167 426 25223
rect 482 25167 518 25223
rect 574 25167 610 25223
rect 666 25167 702 25223
rect 758 25167 836 25223
rect 219 25143 836 25167
rect 219 25087 242 25143
rect 298 25087 334 25143
rect 390 25087 426 25143
rect 482 25087 518 25143
rect 574 25087 610 25143
rect 666 25087 702 25143
rect 758 25087 836 25143
rect 219 25063 836 25087
rect 219 25007 242 25063
rect 298 25007 334 25063
rect 390 25007 426 25063
rect 482 25007 518 25063
rect 574 25007 610 25063
rect 666 25007 702 25063
rect 758 25007 836 25063
rect 219 24983 836 25007
rect 219 24927 242 24983
rect 298 24927 334 24983
rect 390 24927 426 24983
rect 482 24927 518 24983
rect 574 24927 610 24983
rect 666 24927 702 24983
rect 758 24927 836 24983
rect 219 24903 836 24927
rect 219 24847 242 24903
rect 298 24847 334 24903
rect 390 24847 426 24903
rect 482 24847 518 24903
rect 574 24847 610 24903
rect 666 24847 702 24903
rect 758 24847 836 24903
tri 961 28365 991 28395 se
rect 991 28365 2078 28395
rect 961 28348 2078 28365
rect 961 28284 963 28348
rect 1027 28284 1057 28348
rect 1121 28284 1151 28348
rect 1215 28284 1245 28348
rect 1309 28284 1339 28348
rect 1403 28284 1433 28348
rect 1497 28284 2078 28348
rect 961 28268 2078 28284
rect 961 28204 963 28268
rect 1027 28204 1057 28268
rect 1121 28204 1151 28268
rect 1215 28204 1245 28268
rect 1309 28204 1339 28268
rect 1403 28204 1433 28268
rect 1497 28204 2078 28268
rect 961 28188 2078 28204
rect 961 28124 963 28188
rect 1027 28124 1057 28188
rect 1121 28124 1151 28188
rect 1215 28124 1245 28188
rect 1309 28124 1339 28188
rect 1403 28124 1433 28188
rect 1497 28124 2078 28188
rect 961 28108 2078 28124
rect 961 28044 963 28108
rect 1027 28044 1057 28108
rect 1121 28044 1151 28108
rect 1215 28044 1245 28108
rect 1309 28044 1339 28108
rect 1403 28044 1433 28108
rect 1497 28044 2078 28108
rect 961 28028 2078 28044
rect 961 27964 963 28028
rect 1027 27964 1057 28028
rect 1121 27964 1151 28028
rect 1215 27964 1245 28028
rect 1309 27964 1339 28028
rect 1403 27964 1433 28028
rect 1497 27964 2078 28028
rect 961 27948 2078 27964
rect 961 27884 963 27948
rect 1027 27884 1057 27948
rect 1121 27884 1151 27948
rect 1215 27884 1245 27948
rect 1309 27884 1339 27948
rect 1403 27884 1433 27948
rect 1497 27884 2078 27948
rect 961 27867 2078 27884
rect 961 27803 963 27867
rect 1027 27803 1057 27867
rect 1121 27803 1151 27867
rect 1215 27803 1245 27867
rect 1309 27803 1339 27867
rect 1403 27803 1433 27867
rect 1497 27803 2078 27867
rect 961 27786 2078 27803
rect 961 27722 963 27786
rect 1027 27722 1057 27786
rect 1121 27722 1151 27786
rect 1215 27722 1245 27786
rect 1309 27722 1339 27786
rect 1403 27722 1433 27786
rect 1497 27722 2078 27786
rect 961 27705 2078 27722
rect 961 27641 963 27705
rect 1027 27641 1057 27705
rect 1121 27641 1151 27705
rect 1215 27641 1245 27705
rect 1309 27641 1339 27705
rect 1403 27641 1433 27705
rect 1497 27641 2078 27705
rect 961 27624 2078 27641
rect 961 27560 963 27624
rect 1027 27560 1057 27624
rect 1121 27560 1151 27624
rect 1215 27560 1245 27624
rect 1309 27560 1339 27624
rect 1403 27560 1433 27624
rect 1497 27560 2078 27624
rect 961 27543 2078 27560
rect 961 27479 963 27543
rect 1027 27479 1057 27543
rect 1121 27479 1151 27543
rect 1215 27479 1245 27543
rect 1309 27479 1339 27543
rect 1403 27479 1433 27543
rect 1497 27479 2078 27543
rect 961 27462 2078 27479
rect 961 27398 963 27462
rect 1027 27398 1057 27462
rect 1121 27398 1151 27462
rect 1215 27398 1245 27462
rect 1309 27398 1339 27462
rect 1403 27398 1433 27462
rect 1497 27398 2078 27462
rect 961 27381 2078 27398
rect 961 27317 963 27381
rect 1027 27317 1057 27381
rect 1121 27317 1151 27381
rect 1215 27317 1245 27381
rect 1309 27317 1339 27381
rect 1403 27317 1433 27381
rect 1497 27317 2078 27381
rect 961 27300 2078 27317
rect 961 27236 963 27300
rect 1027 27236 1057 27300
rect 1121 27236 1151 27300
rect 1215 27236 1245 27300
rect 1309 27236 1339 27300
rect 1403 27236 1433 27300
rect 1497 27236 2078 27300
rect 961 27219 2078 27236
rect 961 27155 963 27219
rect 1027 27155 1057 27219
rect 1121 27155 1151 27219
rect 1215 27155 1245 27219
rect 1309 27155 1339 27219
rect 1403 27155 1433 27219
rect 1497 27155 2078 27219
rect 961 27138 2078 27155
rect 961 27074 963 27138
rect 1027 27074 1057 27138
rect 1121 27074 1151 27138
rect 1215 27074 1245 27138
rect 1309 27074 1339 27138
rect 1403 27074 1433 27138
rect 1497 27074 2078 27138
rect 961 27057 2078 27074
rect 961 26993 963 27057
rect 1027 26993 1057 27057
rect 1121 26993 1151 27057
rect 1215 26993 1245 27057
rect 1309 26993 1339 27057
rect 1403 26993 1433 27057
rect 1497 26993 2078 27057
rect 961 26976 2078 26993
rect 961 26912 963 26976
rect 1027 26912 1057 26976
rect 1121 26912 1151 26976
rect 1215 26912 1245 26976
rect 1309 26912 1339 26976
rect 1403 26912 1433 26976
rect 1497 26912 2078 26976
rect 961 26895 2078 26912
rect 961 26831 963 26895
rect 1027 26831 1057 26895
rect 1121 26831 1151 26895
rect 1215 26831 1245 26895
rect 1309 26831 1339 26895
rect 1403 26831 1433 26895
rect 1497 26831 2078 26895
rect 2382 32018 2574 34764
rect 3374 39592 3566 39600
rect 3438 39528 3502 39592
rect 3374 39512 3566 39528
rect 3438 39448 3502 39512
rect 3374 39432 3566 39448
rect 3438 39368 3502 39432
rect 3374 39352 3566 39368
rect 3438 39288 3502 39352
rect 3374 39272 3566 39288
rect 3438 39208 3502 39272
rect 3374 39192 3566 39208
rect 3438 39128 3502 39192
rect 3374 39112 3566 39128
rect 3438 39048 3502 39112
rect 3374 39032 3566 39048
rect 3438 38968 3502 39032
rect 3374 38952 3566 38968
rect 3438 38888 3502 38952
rect 3374 38872 3566 38888
rect 3438 38808 3502 38872
rect 3374 38792 3566 38808
rect 3438 38728 3502 38792
rect 3374 38712 3566 38728
rect 3438 38648 3502 38712
rect 3374 38632 3566 38648
rect 3438 38568 3502 38632
rect 3374 38552 3566 38568
rect 3438 38488 3502 38552
rect 3374 38472 3566 38488
rect 3438 38408 3502 38472
rect 3374 38392 3566 38408
rect 3438 38328 3502 38392
rect 3374 38311 3566 38328
rect 3438 38247 3502 38311
rect 3374 38230 3566 38247
rect 3438 38166 3502 38230
rect 3374 38149 3566 38166
rect 3438 38085 3502 38149
rect 3374 38068 3566 38085
rect 3438 38004 3502 38068
rect 3374 37987 3566 38004
rect 3438 37923 3502 37987
rect 3374 37906 3566 37923
rect 3438 37842 3502 37906
rect 3374 37825 3566 37842
rect 3438 37761 3502 37825
rect 3374 37744 3566 37761
rect 3438 37680 3502 37744
rect 3374 37663 3566 37680
rect 3438 37599 3502 37663
rect 3374 37582 3566 37599
rect 3438 37518 3502 37582
rect 3374 37501 3566 37518
rect 3438 37437 3502 37501
rect 3374 37420 3566 37437
rect 3438 37356 3502 37420
rect 3374 37339 3566 37356
rect 3438 37275 3502 37339
rect 3374 37258 3566 37275
rect 3438 37194 3502 37258
rect 3374 37177 3566 37194
rect 3438 37113 3502 37177
rect 3374 37096 3566 37113
rect 3438 37032 3502 37096
rect 3374 37015 3566 37032
rect 3438 36951 3502 37015
rect 3374 36934 3566 36951
rect 3438 36870 3502 36934
rect 3374 36853 3566 36870
rect 3438 36789 3502 36853
rect 3374 36772 3566 36789
rect 3438 36708 3502 36772
rect 3374 36691 3566 36708
rect 3438 36627 3502 36691
rect 3374 36610 3566 36627
rect 3438 36546 3502 36610
rect 3374 36529 3566 36546
rect 3438 36465 3502 36529
rect 3374 36448 3566 36465
rect 3438 36384 3502 36448
rect 3374 36367 3566 36384
rect 3438 36303 3502 36367
rect 3374 36286 3566 36303
rect 3438 36222 3502 36286
rect 3374 36205 3566 36222
rect 3438 36141 3502 36205
rect 3374 36124 3566 36141
rect 3438 36060 3502 36124
rect 3374 36043 3566 36060
rect 3438 35979 3502 36043
rect 3374 35962 3566 35979
rect 3438 35898 3502 35962
rect 3374 35881 3566 35898
rect 3438 35817 3502 35881
rect 3374 35800 3566 35817
rect 3438 35736 3502 35800
rect 3374 35719 3566 35736
rect 3438 35655 3502 35719
rect 3374 35638 3566 35655
rect 3438 35574 3502 35638
rect 3374 35557 3566 35574
rect 3438 35493 3502 35557
rect 3374 35476 3566 35493
rect 3438 35412 3502 35476
rect 3374 35395 3566 35412
rect 3438 35331 3502 35395
rect 3374 35314 3566 35331
rect 3438 35250 3502 35314
rect 3374 35233 3566 35250
rect 3438 35169 3502 35233
rect 3374 35152 3566 35169
rect 3438 35088 3502 35152
rect 3374 35071 3566 35088
rect 3438 35007 3502 35071
rect 3374 34990 3566 35007
rect 3438 34926 3502 34990
rect 3374 34909 3566 34926
rect 3438 34845 3502 34909
rect 3374 34828 3566 34845
rect 3438 34764 3502 34828
rect 2382 31962 2387 32018
rect 2443 31962 2513 32018
rect 2569 31962 2574 32018
rect 2382 31936 2574 31962
rect 2382 31880 2387 31936
rect 2443 31880 2513 31936
rect 2569 31880 2574 31936
rect 2382 31854 2574 31880
rect 2382 31798 2387 31854
rect 2443 31798 2513 31854
rect 2569 31798 2574 31854
rect 2382 31772 2574 31798
rect 2382 31716 2387 31772
rect 2443 31716 2513 31772
rect 2569 31716 2574 31772
rect 2382 31690 2574 31716
rect 2382 31634 2387 31690
rect 2443 31634 2513 31690
rect 2569 31634 2574 31690
rect 2382 31608 2574 31634
rect 2382 31552 2387 31608
rect 2443 31552 2513 31608
rect 2569 31552 2574 31608
rect 2382 31526 2574 31552
rect 2382 31470 2387 31526
rect 2443 31470 2513 31526
rect 2569 31470 2574 31526
rect 2382 31444 2574 31470
rect 2382 31388 2387 31444
rect 2443 31388 2513 31444
rect 2569 31388 2574 31444
rect 2382 31362 2574 31388
rect 2382 31306 2387 31362
rect 2443 31306 2513 31362
rect 2569 31306 2574 31362
rect 2382 31280 2574 31306
rect 2382 31224 2387 31280
rect 2443 31224 2513 31280
rect 2569 31224 2574 31280
rect 2382 31198 2574 31224
rect 2382 31142 2387 31198
rect 2443 31142 2513 31198
rect 2569 31142 2574 31198
rect 2382 31116 2574 31142
rect 2382 31060 2387 31116
rect 2443 31060 2513 31116
rect 2569 31060 2574 31116
rect 2382 31034 2574 31060
rect 2382 30978 2387 31034
rect 2443 30978 2513 31034
rect 2569 30978 2574 31034
rect 2382 30952 2574 30978
rect 2382 30896 2387 30952
rect 2443 30896 2513 30952
rect 2569 30896 2574 30952
rect 2382 30870 2574 30896
rect 2382 30814 2387 30870
rect 2443 30814 2513 30870
rect 2569 30814 2574 30870
rect 2382 30788 2574 30814
rect 2382 30732 2387 30788
rect 2443 30732 2513 30788
rect 2569 30732 2574 30788
rect 2382 30706 2574 30732
rect 2382 30650 2387 30706
rect 2443 30650 2513 30706
rect 2569 30650 2574 30706
rect 2382 30624 2574 30650
rect 2382 30568 2387 30624
rect 2443 30568 2513 30624
rect 2569 30568 2574 30624
rect 2382 30542 2574 30568
rect 2382 30486 2387 30542
rect 2443 30486 2513 30542
rect 2569 30486 2574 30542
rect 2382 30460 2574 30486
rect 2382 30404 2387 30460
rect 2443 30404 2513 30460
rect 2569 30404 2574 30460
rect 2382 30378 2574 30404
rect 2382 30322 2387 30378
rect 2443 30322 2513 30378
rect 2569 30322 2574 30378
rect 2382 30296 2574 30322
rect 2382 30240 2387 30296
rect 2443 30240 2513 30296
rect 2569 30240 2574 30296
rect 2382 30214 2574 30240
rect 2382 30158 2387 30214
rect 2443 30158 2513 30214
rect 2569 30158 2574 30214
rect 2382 30132 2574 30158
rect 2382 30076 2387 30132
rect 2443 30076 2513 30132
rect 2569 30076 2574 30132
rect 2382 30050 2574 30076
rect 2382 29994 2387 30050
rect 2443 29994 2513 30050
rect 2569 29994 2574 30050
rect 2382 29968 2574 29994
rect 2382 29912 2387 29968
rect 2443 29912 2513 29968
rect 2569 29912 2574 29968
rect 2382 29886 2574 29912
rect 2382 29830 2387 29886
rect 2443 29830 2513 29886
rect 2569 29830 2574 29886
rect 2382 29804 2574 29830
rect 2382 29748 2387 29804
rect 2443 29748 2513 29804
rect 2569 29748 2574 29804
rect 2382 29722 2574 29748
rect 2382 29666 2387 29722
rect 2443 29666 2513 29722
rect 2569 29666 2574 29722
rect 2382 29640 2574 29666
rect 2382 29584 2387 29640
rect 2443 29584 2513 29640
rect 2569 29584 2574 29640
rect 2382 29558 2574 29584
rect 2382 29502 2387 29558
rect 2443 29502 2513 29558
rect 2569 29502 2574 29558
rect 2382 29476 2574 29502
rect 2382 29420 2387 29476
rect 2443 29420 2513 29476
rect 2569 29420 2574 29476
rect 2382 27151 2574 29420
rect 2382 27095 2387 27151
rect 2443 27095 2513 27151
rect 2569 27095 2574 27151
rect 2382 27031 2574 27095
rect 2382 26975 2387 27031
rect 2443 26975 2513 27031
rect 2569 26975 2574 27031
rect 2382 26911 2574 26975
rect 2382 26855 2387 26911
rect 2443 26855 2513 26911
rect 2569 26855 2574 26911
rect 2382 26845 2574 26855
rect 2878 34219 3070 34225
rect 2942 34155 3006 34219
rect 2878 34125 3070 34155
rect 2942 34061 3006 34125
rect 2878 34030 3070 34061
rect 2942 33966 3006 34030
rect 2878 33935 3070 33966
rect 2942 33871 3006 33935
rect 2878 33840 3070 33871
rect 2942 33776 3006 33840
rect 2878 33745 3070 33776
rect 2942 33681 3006 33745
rect 2878 32018 3070 33681
rect 2878 31962 2883 32018
rect 2939 31962 3009 32018
rect 3065 31962 3070 32018
rect 2878 31936 3070 31962
rect 2878 31880 2883 31936
rect 2939 31880 3009 31936
rect 3065 31880 3070 31936
rect 2878 31854 3070 31880
rect 2878 31798 2883 31854
rect 2939 31798 3009 31854
rect 3065 31798 3070 31854
rect 2878 31772 3070 31798
rect 2878 31716 2883 31772
rect 2939 31716 3009 31772
rect 3065 31716 3070 31772
rect 2878 31690 3070 31716
rect 2878 31634 2883 31690
rect 2939 31634 3009 31690
rect 3065 31634 3070 31690
rect 2878 31608 3070 31634
rect 2878 31552 2883 31608
rect 2939 31552 3009 31608
rect 3065 31552 3070 31608
rect 2878 31526 3070 31552
rect 2878 31470 2883 31526
rect 2939 31470 3009 31526
rect 3065 31470 3070 31526
rect 2878 31444 3070 31470
rect 2878 31388 2883 31444
rect 2939 31388 3009 31444
rect 3065 31388 3070 31444
rect 2878 31362 3070 31388
rect 2878 31306 2883 31362
rect 2939 31306 3009 31362
rect 3065 31306 3070 31362
rect 2878 31280 3070 31306
rect 2878 31224 2883 31280
rect 2939 31224 3009 31280
rect 3065 31224 3070 31280
rect 2878 31198 3070 31224
rect 2878 31142 2883 31198
rect 2939 31142 3009 31198
rect 3065 31142 3070 31198
rect 2878 31116 3070 31142
rect 2878 31060 2883 31116
rect 2939 31060 3009 31116
rect 3065 31060 3070 31116
rect 2878 31034 3070 31060
rect 2878 30978 2883 31034
rect 2939 30978 3009 31034
rect 3065 30978 3070 31034
rect 2878 30952 3070 30978
rect 2878 30896 2883 30952
rect 2939 30896 3009 30952
rect 3065 30896 3070 30952
rect 2878 30870 3070 30896
rect 2878 30814 2883 30870
rect 2939 30814 3009 30870
rect 3065 30814 3070 30870
rect 2878 30788 3070 30814
rect 2878 30732 2883 30788
rect 2939 30732 3009 30788
rect 3065 30732 3070 30788
rect 2878 30706 3070 30732
rect 2878 30650 2883 30706
rect 2939 30650 3009 30706
rect 3065 30650 3070 30706
rect 2878 30624 3070 30650
rect 2878 30568 2883 30624
rect 2939 30568 3009 30624
rect 3065 30568 3070 30624
rect 2878 30542 3070 30568
rect 2878 30486 2883 30542
rect 2939 30486 3009 30542
rect 3065 30486 3070 30542
rect 2878 30460 3070 30486
rect 2878 30404 2883 30460
rect 2939 30404 3009 30460
rect 3065 30404 3070 30460
rect 2878 30378 3070 30404
rect 2878 30322 2883 30378
rect 2939 30322 3009 30378
rect 3065 30322 3070 30378
rect 2878 30296 3070 30322
rect 2878 30240 2883 30296
rect 2939 30240 3009 30296
rect 3065 30240 3070 30296
rect 2878 30214 3070 30240
rect 2878 30158 2883 30214
rect 2939 30158 3009 30214
rect 3065 30158 3070 30214
rect 2878 30132 3070 30158
rect 2878 30076 2883 30132
rect 2939 30076 3009 30132
rect 3065 30076 3070 30132
rect 2878 30050 3070 30076
rect 2878 29994 2883 30050
rect 2939 29994 3009 30050
rect 3065 29994 3070 30050
rect 2878 29968 3070 29994
rect 2878 29912 2883 29968
rect 2939 29912 3009 29968
rect 3065 29912 3070 29968
rect 2878 29886 3070 29912
rect 2878 29830 2883 29886
rect 2939 29830 3009 29886
rect 3065 29830 3070 29886
rect 2878 29804 3070 29830
rect 2878 29748 2883 29804
rect 2939 29748 3009 29804
rect 3065 29748 3070 29804
rect 2878 29722 3070 29748
rect 2878 29666 2883 29722
rect 2939 29666 3009 29722
rect 3065 29666 3070 29722
rect 2878 29640 3070 29666
rect 2878 29584 2883 29640
rect 2939 29584 3009 29640
rect 3065 29584 3070 29640
rect 2878 29558 3070 29584
rect 2878 29502 2883 29558
rect 2939 29502 3009 29558
rect 3065 29502 3070 29558
rect 2878 29476 3070 29502
rect 2878 29420 2883 29476
rect 2939 29420 3009 29476
rect 3065 29420 3070 29476
rect 2878 26921 3070 29420
rect 3374 32018 3566 34764
rect 4366 39592 4558 39600
rect 4430 39528 4494 39592
rect 4366 39512 4558 39528
rect 4430 39448 4494 39512
rect 4366 39432 4558 39448
rect 4430 39368 4494 39432
rect 4366 39352 4558 39368
rect 4430 39288 4494 39352
rect 4366 39272 4558 39288
rect 4430 39208 4494 39272
rect 4366 39192 4558 39208
rect 4430 39128 4494 39192
rect 4366 39112 4558 39128
rect 4430 39048 4494 39112
rect 4366 39032 4558 39048
rect 4430 38968 4494 39032
rect 4366 38952 4558 38968
rect 4430 38888 4494 38952
rect 4366 38872 4558 38888
rect 4430 38808 4494 38872
rect 4366 38792 4558 38808
rect 4430 38728 4494 38792
rect 4366 38712 4558 38728
rect 4430 38648 4494 38712
rect 4366 38632 4558 38648
rect 4430 38568 4494 38632
rect 4366 38552 4558 38568
rect 4430 38488 4494 38552
rect 4366 38472 4558 38488
rect 4430 38408 4494 38472
rect 4366 38392 4558 38408
rect 4430 38328 4494 38392
rect 4366 38311 4558 38328
rect 4430 38247 4494 38311
rect 4366 38230 4558 38247
rect 4430 38166 4494 38230
rect 4366 38149 4558 38166
rect 4430 38085 4494 38149
rect 4366 38068 4558 38085
rect 4430 38004 4494 38068
rect 4366 37987 4558 38004
rect 4430 37923 4494 37987
rect 4366 37906 4558 37923
rect 4430 37842 4494 37906
rect 4366 37825 4558 37842
rect 4430 37761 4494 37825
rect 4366 37744 4558 37761
rect 4430 37680 4494 37744
rect 4366 37663 4558 37680
rect 4430 37599 4494 37663
rect 4366 37582 4558 37599
rect 4430 37518 4494 37582
rect 4366 37501 4558 37518
rect 4430 37437 4494 37501
rect 4366 37420 4558 37437
rect 4430 37356 4494 37420
rect 4366 37339 4558 37356
rect 4430 37275 4494 37339
rect 4366 37258 4558 37275
rect 4430 37194 4494 37258
rect 4366 37177 4558 37194
rect 4430 37113 4494 37177
rect 4366 37096 4558 37113
rect 4430 37032 4494 37096
rect 4366 37015 4558 37032
rect 4430 36951 4494 37015
rect 4366 36934 4558 36951
rect 4430 36870 4494 36934
rect 4366 36853 4558 36870
rect 4430 36789 4494 36853
rect 4366 36772 4558 36789
rect 4430 36708 4494 36772
rect 4366 36691 4558 36708
rect 4430 36627 4494 36691
rect 4366 36610 4558 36627
rect 4430 36546 4494 36610
rect 4366 36529 4558 36546
rect 4430 36465 4494 36529
rect 4366 36448 4558 36465
rect 4430 36384 4494 36448
rect 4366 36367 4558 36384
rect 4430 36303 4494 36367
rect 4366 36286 4558 36303
rect 4430 36222 4494 36286
rect 4366 36205 4558 36222
rect 4430 36141 4494 36205
rect 4366 36124 4558 36141
rect 4430 36060 4494 36124
rect 4366 36043 4558 36060
rect 4430 35979 4494 36043
rect 4366 35962 4558 35979
rect 4430 35898 4494 35962
rect 4366 35881 4558 35898
rect 4430 35817 4494 35881
rect 4366 35800 4558 35817
rect 4430 35736 4494 35800
rect 4366 35719 4558 35736
rect 4430 35655 4494 35719
rect 4366 35638 4558 35655
rect 4430 35574 4494 35638
rect 4366 35557 4558 35574
rect 4430 35493 4494 35557
rect 4366 35476 4558 35493
rect 4430 35412 4494 35476
rect 4366 35395 4558 35412
rect 4430 35331 4494 35395
rect 4366 35314 4558 35331
rect 4430 35250 4494 35314
rect 4366 35233 4558 35250
rect 4430 35169 4494 35233
rect 4366 35152 4558 35169
rect 4430 35088 4494 35152
rect 4366 35071 4558 35088
rect 4430 35007 4494 35071
rect 4366 34990 4558 35007
rect 4430 34926 4494 34990
rect 4366 34909 4558 34926
rect 4430 34845 4494 34909
rect 4366 34828 4558 34845
rect 4430 34764 4494 34828
rect 3374 31962 3379 32018
rect 3435 31962 3505 32018
rect 3561 31962 3566 32018
rect 3374 31936 3566 31962
rect 3374 31880 3379 31936
rect 3435 31880 3505 31936
rect 3561 31880 3566 31936
rect 3374 31854 3566 31880
rect 3374 31798 3379 31854
rect 3435 31798 3505 31854
rect 3561 31798 3566 31854
rect 3374 31772 3566 31798
rect 3374 31716 3379 31772
rect 3435 31716 3505 31772
rect 3561 31716 3566 31772
rect 3374 31690 3566 31716
rect 3374 31634 3379 31690
rect 3435 31634 3505 31690
rect 3561 31634 3566 31690
rect 3374 31608 3566 31634
rect 3374 31552 3379 31608
rect 3435 31552 3505 31608
rect 3561 31552 3566 31608
rect 3374 31526 3566 31552
rect 3374 31470 3379 31526
rect 3435 31470 3505 31526
rect 3561 31470 3566 31526
rect 3374 31444 3566 31470
rect 3374 31388 3379 31444
rect 3435 31388 3505 31444
rect 3561 31388 3566 31444
rect 3374 31362 3566 31388
rect 3374 31306 3379 31362
rect 3435 31306 3505 31362
rect 3561 31306 3566 31362
rect 3374 31280 3566 31306
rect 3374 31224 3379 31280
rect 3435 31224 3505 31280
rect 3561 31224 3566 31280
rect 3374 31198 3566 31224
rect 3374 31142 3379 31198
rect 3435 31142 3505 31198
rect 3561 31142 3566 31198
rect 3374 31116 3566 31142
rect 3374 31060 3379 31116
rect 3435 31060 3505 31116
rect 3561 31060 3566 31116
rect 3374 31034 3566 31060
rect 3374 30978 3379 31034
rect 3435 30978 3505 31034
rect 3561 30978 3566 31034
rect 3374 30952 3566 30978
rect 3374 30896 3379 30952
rect 3435 30896 3505 30952
rect 3561 30896 3566 30952
rect 3374 30870 3566 30896
rect 3374 30814 3379 30870
rect 3435 30814 3505 30870
rect 3561 30814 3566 30870
rect 3374 30788 3566 30814
rect 3374 30732 3379 30788
rect 3435 30732 3505 30788
rect 3561 30732 3566 30788
rect 3374 30706 3566 30732
rect 3374 30650 3379 30706
rect 3435 30650 3505 30706
rect 3561 30650 3566 30706
rect 3374 30624 3566 30650
rect 3374 30568 3379 30624
rect 3435 30568 3505 30624
rect 3561 30568 3566 30624
rect 3374 30542 3566 30568
rect 3374 30486 3379 30542
rect 3435 30486 3505 30542
rect 3561 30486 3566 30542
rect 3374 30460 3566 30486
rect 3374 30404 3379 30460
rect 3435 30404 3505 30460
rect 3561 30404 3566 30460
rect 3374 30378 3566 30404
rect 3374 30322 3379 30378
rect 3435 30322 3505 30378
rect 3561 30322 3566 30378
rect 3374 30296 3566 30322
rect 3374 30240 3379 30296
rect 3435 30240 3505 30296
rect 3561 30240 3566 30296
rect 3374 30214 3566 30240
rect 3374 30158 3379 30214
rect 3435 30158 3505 30214
rect 3561 30158 3566 30214
rect 3374 30132 3566 30158
rect 3374 30076 3379 30132
rect 3435 30076 3505 30132
rect 3561 30076 3566 30132
rect 3374 30050 3566 30076
rect 3374 29994 3379 30050
rect 3435 29994 3505 30050
rect 3561 29994 3566 30050
rect 3374 29968 3566 29994
rect 3374 29912 3379 29968
rect 3435 29912 3505 29968
rect 3561 29912 3566 29968
rect 3374 29886 3566 29912
rect 3374 29830 3379 29886
rect 3435 29830 3505 29886
rect 3561 29830 3566 29886
rect 3374 29804 3566 29830
rect 3374 29748 3379 29804
rect 3435 29748 3505 29804
rect 3561 29748 3566 29804
rect 3374 29722 3566 29748
rect 3374 29666 3379 29722
rect 3435 29666 3505 29722
rect 3561 29666 3566 29722
rect 3374 29640 3566 29666
rect 3374 29584 3379 29640
rect 3435 29584 3505 29640
rect 3561 29584 3566 29640
rect 3374 29558 3566 29584
rect 3374 29502 3379 29558
rect 3435 29502 3505 29558
rect 3561 29502 3566 29558
rect 3374 29476 3566 29502
rect 3374 29420 3379 29476
rect 3435 29420 3505 29476
rect 3561 29420 3566 29476
rect 3374 29415 3566 29420
rect 3870 34219 4062 34225
rect 3934 34155 3998 34219
rect 3870 34125 4062 34155
rect 3934 34061 3998 34125
rect 3870 34030 4062 34061
rect 3934 33966 3998 34030
rect 3870 33935 4062 33966
rect 3934 33871 3998 33935
rect 3870 33840 4062 33871
rect 3934 33776 3998 33840
rect 3870 33745 4062 33776
rect 3934 33681 3998 33745
rect 3870 32018 4062 33681
rect 3870 31962 3875 32018
rect 3931 31962 4001 32018
rect 4057 31962 4062 32018
rect 3870 31936 4062 31962
rect 3870 31880 3875 31936
rect 3931 31880 4001 31936
rect 4057 31880 4062 31936
rect 3870 31854 4062 31880
rect 3870 31798 3875 31854
rect 3931 31798 4001 31854
rect 4057 31798 4062 31854
rect 3870 31772 4062 31798
rect 3870 31716 3875 31772
rect 3931 31716 4001 31772
rect 4057 31716 4062 31772
rect 3870 31690 4062 31716
rect 3870 31634 3875 31690
rect 3931 31634 4001 31690
rect 4057 31634 4062 31690
rect 3870 31608 4062 31634
rect 3870 31552 3875 31608
rect 3931 31552 4001 31608
rect 4057 31552 4062 31608
rect 3870 31526 4062 31552
rect 3870 31470 3875 31526
rect 3931 31470 4001 31526
rect 4057 31470 4062 31526
rect 3870 31444 4062 31470
rect 3870 31388 3875 31444
rect 3931 31388 4001 31444
rect 4057 31388 4062 31444
rect 3870 31362 4062 31388
rect 3870 31306 3875 31362
rect 3931 31306 4001 31362
rect 4057 31306 4062 31362
rect 3870 31280 4062 31306
rect 3870 31224 3875 31280
rect 3931 31224 4001 31280
rect 4057 31224 4062 31280
rect 3870 31198 4062 31224
rect 3870 31142 3875 31198
rect 3931 31142 4001 31198
rect 4057 31142 4062 31198
rect 3870 31116 4062 31142
rect 3870 31060 3875 31116
rect 3931 31060 4001 31116
rect 4057 31060 4062 31116
rect 3870 31034 4062 31060
rect 3870 30978 3875 31034
rect 3931 30978 4001 31034
rect 4057 30978 4062 31034
rect 3870 30952 4062 30978
rect 3870 30896 3875 30952
rect 3931 30896 4001 30952
rect 4057 30896 4062 30952
rect 3870 30870 4062 30896
rect 3870 30814 3875 30870
rect 3931 30814 4001 30870
rect 4057 30814 4062 30870
rect 3870 30788 4062 30814
rect 3870 30732 3875 30788
rect 3931 30732 4001 30788
rect 4057 30732 4062 30788
rect 3870 30706 4062 30732
rect 3870 30650 3875 30706
rect 3931 30650 4001 30706
rect 4057 30650 4062 30706
rect 3870 30624 4062 30650
rect 3870 30568 3875 30624
rect 3931 30568 4001 30624
rect 4057 30568 4062 30624
rect 3870 30542 4062 30568
rect 3870 30486 3875 30542
rect 3931 30486 4001 30542
rect 4057 30486 4062 30542
rect 3870 30460 4062 30486
rect 3870 30404 3875 30460
rect 3931 30404 4001 30460
rect 4057 30404 4062 30460
rect 3870 30378 4062 30404
rect 3870 30322 3875 30378
rect 3931 30322 4001 30378
rect 4057 30322 4062 30378
rect 3870 30296 4062 30322
rect 3870 30240 3875 30296
rect 3931 30240 4001 30296
rect 4057 30240 4062 30296
rect 3870 30214 4062 30240
rect 3870 30158 3875 30214
rect 3931 30158 4001 30214
rect 4057 30158 4062 30214
rect 3870 30132 4062 30158
rect 3870 30076 3875 30132
rect 3931 30076 4001 30132
rect 4057 30076 4062 30132
rect 3870 30050 4062 30076
rect 3870 29994 3875 30050
rect 3931 29994 4001 30050
rect 4057 29994 4062 30050
rect 3870 29968 4062 29994
rect 3870 29912 3875 29968
rect 3931 29912 4001 29968
rect 4057 29912 4062 29968
rect 3870 29886 4062 29912
rect 3870 29830 3875 29886
rect 3931 29830 4001 29886
rect 4057 29830 4062 29886
rect 3870 29804 4062 29830
rect 3870 29748 3875 29804
rect 3931 29748 4001 29804
rect 4057 29748 4062 29804
rect 3870 29722 4062 29748
rect 3870 29666 3875 29722
rect 3931 29666 4001 29722
rect 4057 29666 4062 29722
rect 3870 29640 4062 29666
rect 3870 29584 3875 29640
rect 3931 29584 4001 29640
rect 4057 29584 4062 29640
rect 3870 29558 4062 29584
rect 3870 29502 3875 29558
rect 3931 29502 4001 29558
rect 4057 29502 4062 29558
rect 3870 29476 4062 29502
rect 3870 29420 3875 29476
rect 3931 29420 4001 29476
rect 4057 29420 4062 29476
rect 3472 28620 3570 28633
rect 3472 28564 3494 28620
rect 3550 28564 3570 28620
rect 3472 28451 3570 28564
rect 3472 28395 3494 28451
rect 3550 28395 3570 28451
rect 3472 28282 3570 28395
rect 3472 28226 3494 28282
rect 3550 28226 3570 28282
rect 3472 28112 3570 28226
rect 3472 28056 3494 28112
rect 3550 28056 3570 28112
rect 3472 27942 3570 28056
rect 3472 27886 3494 27942
rect 3550 27886 3570 27942
rect 3472 27772 3570 27886
rect 3472 27716 3494 27772
rect 3550 27716 3570 27772
rect 3472 27602 3570 27716
rect 3472 27546 3494 27602
rect 3550 27546 3570 27602
rect 3472 27432 3570 27546
rect 3472 27376 3494 27432
rect 3550 27376 3570 27432
rect 3472 27262 3570 27376
rect 3472 27206 3494 27262
rect 3550 27206 3570 27262
tri 3070 26921 3101 26952 sw
rect 2878 26897 3101 26921
tri 3101 26897 3125 26921 sw
rect 2878 26884 3125 26897
tri 3125 26884 3138 26897 sw
rect 2878 26858 3138 26884
tri 3138 26858 3164 26884 sw
rect 961 26814 2078 26831
rect 961 26750 963 26814
rect 1027 26750 1057 26814
rect 1121 26750 1151 26814
rect 1215 26750 1245 26814
rect 1309 26750 1339 26814
rect 1403 26750 1433 26814
rect 1497 26750 2078 26814
rect 961 26733 2078 26750
rect 961 26669 963 26733
rect 1027 26669 1057 26733
rect 1121 26669 1151 26733
rect 1215 26669 1245 26733
rect 1309 26669 1339 26733
rect 1403 26669 1433 26733
rect 1497 26669 2078 26733
rect 961 26652 2078 26669
rect 961 26588 963 26652
rect 1027 26588 1057 26652
rect 1121 26588 1151 26652
rect 1215 26588 1245 26652
rect 1309 26588 1339 26652
rect 1403 26588 1433 26652
rect 1497 26588 2078 26652
rect 961 26571 2078 26588
rect 961 26507 963 26571
rect 1027 26507 1057 26571
rect 1121 26507 1151 26571
rect 1215 26507 1245 26571
rect 1309 26507 1339 26571
rect 1403 26507 1433 26571
rect 1497 26507 2078 26571
rect 2878 26566 3164 26858
tri 2878 26548 2896 26566 ne
rect 2896 26548 3164 26566
rect 961 26490 2078 26507
tri 2896 26492 2952 26548 ne
rect 2952 26492 3164 26548
rect 961 26426 963 26490
rect 1027 26426 1057 26490
rect 1121 26426 1151 26490
rect 1215 26426 1245 26490
rect 1309 26426 1339 26490
rect 1403 26426 1433 26490
rect 1497 26426 2078 26490
tri 2952 26464 2980 26492 ne
rect 961 26409 2078 26426
rect 961 26345 963 26409
rect 1027 26345 1057 26409
rect 1121 26345 1151 26409
rect 1215 26345 1245 26409
rect 1309 26345 1339 26409
rect 1403 26345 1433 26409
rect 1497 26345 2078 26409
rect 961 26328 2078 26345
rect 961 26264 963 26328
rect 1027 26264 1057 26328
rect 1121 26264 1151 26328
rect 1215 26264 1245 26328
rect 1309 26264 1339 26328
rect 1403 26264 1433 26328
rect 1497 26264 2078 26328
rect 961 26247 2078 26264
rect 961 26183 963 26247
rect 1027 26183 1057 26247
rect 1121 26183 1151 26247
rect 1215 26183 1245 26247
rect 1309 26183 1339 26247
rect 1403 26183 1433 26247
rect 1497 26183 2078 26247
rect 961 26166 2078 26183
rect 961 26102 963 26166
rect 1027 26102 1057 26166
rect 1121 26102 1151 26166
rect 1215 26102 1245 26166
rect 1309 26102 1339 26166
rect 1403 26102 1433 26166
rect 1497 26102 2078 26166
rect 961 26085 2078 26102
rect 961 26021 963 26085
rect 1027 26021 1057 26085
rect 1121 26021 1151 26085
rect 1215 26021 1245 26085
rect 1309 26021 1339 26085
rect 1403 26021 1433 26085
rect 1497 26021 2078 26085
rect 961 26004 2078 26021
rect 961 25940 963 26004
rect 1027 25940 1057 26004
rect 1121 25940 1151 26004
rect 1215 25940 1245 26004
rect 1309 25940 1339 26004
rect 1403 25940 1433 26004
rect 1497 25940 2078 26004
rect 961 25923 2078 25940
rect 961 25859 963 25923
rect 1027 25859 1057 25923
rect 1121 25859 1151 25923
rect 1215 25859 1245 25923
rect 1309 25859 1339 25923
rect 1403 25859 1433 25923
rect 1497 25859 2078 25923
rect 961 25842 2078 25859
rect 961 25778 963 25842
rect 1027 25778 1057 25842
rect 1121 25778 1151 25842
rect 1215 25778 1245 25842
rect 1309 25778 1339 25842
rect 1403 25778 1433 25842
rect 1497 25778 2078 25842
rect 961 25761 2078 25778
rect 961 25697 963 25761
rect 1027 25697 1057 25761
rect 1121 25697 1151 25761
rect 1215 25697 1245 25761
rect 1309 25697 1339 25761
rect 1403 25697 1433 25761
rect 1497 25697 2078 25761
rect 961 25680 2078 25697
rect 961 25616 963 25680
rect 1027 25616 1057 25680
rect 1121 25616 1151 25680
rect 1215 25616 1245 25680
rect 1309 25616 1339 25680
rect 1403 25616 1433 25680
rect 1497 25616 2078 25680
rect 961 25599 2078 25616
rect 961 25535 963 25599
rect 1027 25535 1057 25599
rect 1121 25535 1151 25599
rect 1215 25535 1245 25599
rect 1309 25535 1339 25599
rect 1403 25535 1433 25599
rect 1497 25535 2078 25599
rect 961 25518 2078 25535
rect 961 25454 963 25518
rect 1027 25454 1057 25518
rect 1121 25454 1151 25518
rect 1215 25454 1245 25518
rect 1309 25454 1339 25518
rect 1403 25454 1433 25518
rect 1497 25454 2078 25518
rect 961 25437 2078 25454
rect 961 25373 963 25437
rect 1027 25373 1057 25437
rect 1121 25373 1151 25437
rect 1215 25373 1245 25437
rect 1309 25373 1339 25437
rect 1403 25373 1433 25437
rect 1497 25373 2078 25437
rect 961 25356 2078 25373
rect 961 25292 963 25356
rect 1027 25292 1057 25356
rect 1121 25292 1151 25356
rect 1215 25292 1245 25356
rect 1309 25292 1339 25356
rect 1403 25292 1433 25356
rect 1497 25292 2078 25356
rect 961 25275 2078 25292
rect 961 25211 963 25275
rect 1027 25211 1057 25275
rect 1121 25211 1151 25275
rect 1215 25211 1245 25275
rect 1309 25211 1339 25275
rect 1403 25211 1433 25275
rect 1497 25211 2078 25275
rect 961 25194 2078 25211
rect 961 25130 963 25194
rect 1027 25130 1057 25194
rect 1121 25130 1151 25194
rect 1215 25130 1245 25194
rect 1309 25130 1339 25194
rect 1403 25130 1433 25194
rect 1497 25130 2078 25194
rect 961 25113 2078 25130
rect 961 25049 963 25113
rect 1027 25049 1057 25113
rect 1121 25049 1151 25113
rect 1215 25049 1245 25113
rect 1309 25049 1339 25113
rect 1403 25049 1433 25113
rect 1497 25049 2078 25113
rect 961 25032 2078 25049
rect 961 24968 963 25032
rect 1027 24968 1057 25032
rect 1121 24968 1151 25032
rect 1215 24968 1245 25032
rect 1309 24968 1339 25032
rect 1403 24968 1433 25032
rect 1497 24968 2078 25032
rect 961 24951 2078 24968
rect 961 24887 963 24951
rect 1027 24887 1057 24951
rect 1121 24887 1151 24951
rect 1215 24887 1245 24951
rect 1309 24887 1339 24951
rect 1403 24887 1433 24951
rect 1497 24887 2078 24951
rect 961 24881 2078 24887
tri 962 24875 968 24881 ne
rect 968 24875 2078 24881
rect 219 24823 836 24847
rect 219 24767 242 24823
rect 298 24767 334 24823
rect 390 24767 426 24823
rect 482 24767 518 24823
rect 574 24767 610 24823
rect 666 24767 702 24823
rect 758 24767 836 24823
tri 968 24819 1024 24875 ne
rect 1024 24819 2078 24875
tri 1024 24794 1049 24819 ne
rect 1049 24794 2078 24819
rect 219 24743 836 24767
rect 219 24687 242 24743
rect 298 24687 334 24743
rect 390 24687 426 24743
rect 482 24687 518 24743
rect 574 24687 610 24743
rect 666 24687 702 24743
rect 758 24687 836 24743
tri 1049 24738 1105 24794 ne
rect 1105 24738 2078 24794
tri 1105 24713 1130 24738 ne
rect 1130 24713 2078 24738
rect 219 24663 836 24687
rect 219 24607 242 24663
rect 298 24607 334 24663
rect 390 24607 426 24663
rect 482 24607 518 24663
rect 574 24607 610 24663
rect 666 24607 702 24663
rect 758 24607 836 24663
tri 1130 24657 1186 24713 ne
rect 1186 24657 2078 24713
tri 1186 24632 1211 24657 ne
rect 1211 24632 2078 24657
tri 1211 24618 1225 24632 ne
rect 1225 24618 2078 24632
rect 2480 26176 2672 26187
rect 2480 26120 2485 26176
rect 2541 26120 2611 26176
rect 2667 26120 2672 26176
rect 2480 26081 2672 26120
rect 2480 26025 2485 26081
rect 2541 26025 2611 26081
rect 2667 26025 2672 26081
rect 2480 25986 2672 26025
rect 2480 25930 2485 25986
rect 2541 25930 2611 25986
rect 2667 25930 2672 25986
rect 2480 25891 2672 25930
rect 2480 25835 2485 25891
rect 2541 25835 2611 25891
rect 2667 25835 2672 25891
rect 2480 25795 2672 25835
rect 2480 25739 2485 25795
rect 2541 25739 2611 25795
rect 2667 25739 2672 25795
rect 2480 25699 2672 25739
rect 2480 25643 2485 25699
rect 2541 25643 2611 25699
rect 2667 25643 2672 25699
rect 219 24583 836 24607
rect 219 24527 242 24583
rect 298 24527 334 24583
rect 390 24527 426 24583
rect 482 24527 518 24583
rect 574 24527 610 24583
rect 666 24527 702 24583
rect 758 24527 836 24583
tri 1225 24576 1267 24618 ne
rect 1267 24576 2078 24618
tri 2078 24576 2120 24618 sw
tri 1267 24551 1292 24576 ne
rect 1292 24551 2120 24576
tri 2120 24551 2145 24576 sw
rect 219 24503 836 24527
tri 1292 24524 1319 24551 ne
rect 1319 24524 2145 24551
tri 2145 24524 2172 24551 sw
rect 219 24447 242 24503
rect 298 24447 334 24503
rect 390 24447 426 24503
rect 482 24447 518 24503
rect 574 24447 610 24503
rect 666 24447 702 24503
rect 758 24447 836 24503
tri 1319 24495 1348 24524 ne
rect 1348 24495 2172 24524
tri 1348 24470 1373 24495 ne
rect 1373 24470 2172 24495
rect 219 24423 836 24447
rect 219 24367 242 24423
rect 298 24367 334 24423
rect 390 24367 426 24423
rect 482 24367 518 24423
rect 574 24367 610 24423
rect 666 24367 702 24423
rect 758 24367 836 24423
tri 1373 24414 1429 24470 ne
rect 1429 24414 2172 24470
tri 1429 24389 1454 24414 ne
rect 1454 24389 2172 24414
rect 219 24343 836 24367
rect 219 24287 242 24343
rect 298 24287 334 24343
rect 390 24287 426 24343
rect 482 24287 518 24343
rect 574 24287 610 24343
rect 666 24287 702 24343
rect 758 24287 836 24343
tri 1454 24333 1510 24389 ne
rect 1510 24333 2172 24389
tri 1510 24308 1535 24333 ne
rect 1535 24308 2172 24333
rect 219 24263 836 24287
rect 219 24207 242 24263
rect 298 24207 334 24263
rect 390 24207 426 24263
rect 482 24207 518 24263
rect 574 24207 610 24263
rect 666 24207 702 24263
rect 758 24207 836 24263
tri 1535 24252 1591 24308 ne
rect 1591 24252 2172 24308
tri 1591 24227 1616 24252 ne
rect 1616 24227 2172 24252
rect 219 24183 836 24207
rect 219 24127 242 24183
rect 298 24127 334 24183
rect 390 24127 426 24183
rect 482 24127 518 24183
rect 574 24127 610 24183
rect 666 24127 702 24183
rect 758 24127 836 24183
tri 1616 24171 1672 24227 ne
rect 1672 24171 2172 24227
tri 1672 24146 1697 24171 ne
rect 1697 24146 2172 24171
rect 219 24103 836 24127
rect 219 24047 242 24103
rect 298 24047 334 24103
rect 390 24047 426 24103
rect 482 24047 518 24103
rect 574 24047 610 24103
rect 666 24047 702 24103
rect 758 24047 836 24103
tri 1697 24090 1753 24146 ne
rect 1753 24090 2172 24146
tri 1753 24065 1778 24090 ne
rect 1778 24065 2172 24090
rect 219 24023 836 24047
rect 219 23967 242 24023
rect 298 23967 334 24023
rect 390 23967 426 24023
rect 482 23967 518 24023
rect 574 23967 610 24023
rect 666 23967 702 24023
rect 758 23967 836 24023
tri 1778 24009 1834 24065 ne
rect 1834 24009 2172 24065
tri 1834 23984 1859 24009 ne
rect 1859 23984 2172 24009
rect 219 23943 836 23967
rect 219 23887 242 23943
rect 298 23887 334 23943
rect 390 23887 426 23943
rect 482 23887 518 23943
rect 574 23887 610 23943
rect 666 23887 702 23943
rect 758 23887 836 23943
tri 1859 23928 1915 23984 ne
rect 1915 23928 2172 23984
tri 1915 23903 1940 23928 ne
rect 1940 23903 2172 23928
rect 219 23863 836 23887
rect 219 23807 242 23863
rect 298 23807 334 23863
rect 390 23807 426 23863
rect 482 23807 518 23863
rect 574 23807 610 23863
rect 666 23807 702 23863
rect 758 23807 836 23863
tri 1940 23861 1982 23903 ne
rect 219 23783 836 23807
rect 219 23727 242 23783
rect 298 23727 334 23783
rect 390 23727 426 23783
rect 482 23727 518 23783
rect 574 23727 610 23783
rect 666 23727 702 23783
rect 758 23727 836 23783
rect 219 23703 836 23727
rect 219 23647 242 23703
rect 298 23647 334 23703
rect 390 23647 426 23703
rect 482 23647 518 23703
rect 574 23647 610 23703
rect 666 23647 702 23703
rect 758 23647 836 23703
rect 219 23623 836 23647
rect 219 23567 242 23623
rect 298 23567 334 23623
rect 390 23567 426 23623
rect 482 23567 518 23623
rect 574 23567 610 23623
rect 666 23567 702 23623
rect 758 23567 836 23623
rect 219 23543 836 23567
rect 219 23487 242 23543
rect 298 23487 334 23543
rect 390 23487 426 23543
rect 482 23487 518 23543
rect 574 23487 610 23543
rect 666 23487 702 23543
rect 758 23487 836 23543
rect 219 23463 836 23487
rect 219 23407 242 23463
rect 298 23407 334 23463
rect 390 23407 426 23463
rect 482 23407 518 23463
rect 574 23407 610 23463
rect 666 23407 702 23463
rect 758 23407 836 23463
rect 219 23383 836 23407
rect 219 23327 242 23383
rect 298 23327 334 23383
rect 390 23327 426 23383
rect 482 23327 518 23383
rect 574 23327 610 23383
rect 666 23327 702 23383
rect 758 23327 836 23383
rect 219 23303 836 23327
rect 219 23247 242 23303
rect 298 23247 334 23303
rect 390 23247 426 23303
rect 482 23247 518 23303
rect 574 23247 610 23303
rect 666 23247 702 23303
rect 758 23247 836 23303
rect 219 23223 836 23247
rect 219 23167 242 23223
rect 298 23167 334 23223
rect 390 23167 426 23223
rect 482 23167 518 23223
rect 574 23167 610 23223
rect 666 23167 702 23223
rect 758 23167 836 23223
rect 219 23143 836 23167
rect 219 23087 242 23143
rect 298 23087 334 23143
rect 390 23087 426 23143
rect 482 23087 518 23143
rect 574 23087 610 23143
rect 666 23087 702 23143
rect 758 23087 836 23143
rect 219 23063 836 23087
rect 219 23007 242 23063
rect 298 23007 334 23063
rect 390 23007 426 23063
rect 482 23007 518 23063
rect 574 23007 610 23063
rect 666 23007 702 23063
rect 758 23007 836 23063
rect 219 22983 836 23007
rect 219 22927 242 22983
rect 298 22927 334 22983
rect 390 22927 426 22983
rect 482 22927 518 22983
rect 574 22927 610 22983
rect 666 22927 702 22983
rect 758 22927 836 22983
rect 219 22903 836 22927
rect 219 22847 242 22903
rect 298 22847 334 22903
rect 390 22847 426 22903
rect 482 22847 518 22903
rect 574 22847 610 22903
rect 666 22847 702 22903
rect 758 22847 836 22903
rect 219 22822 836 22847
rect 219 22766 242 22822
rect 298 22766 334 22822
rect 390 22766 426 22822
rect 482 22766 518 22822
rect 574 22766 610 22822
rect 666 22766 702 22822
rect 758 22766 836 22822
rect 219 22741 836 22766
rect 219 22685 242 22741
rect 298 22685 334 22741
rect 390 22685 426 22741
rect 482 22685 518 22741
rect 574 22685 610 22741
rect 666 22685 702 22741
rect 758 22685 836 22741
rect 219 22660 836 22685
rect 219 22604 242 22660
rect 298 22604 334 22660
rect 390 22604 426 22660
rect 482 22604 518 22660
rect 574 22604 610 22660
rect 666 22604 702 22660
rect 758 22604 836 22660
rect 219 22579 836 22604
rect 219 22523 242 22579
rect 298 22523 334 22579
rect 390 22523 426 22579
rect 482 22523 518 22579
rect 574 22523 610 22579
rect 666 22523 702 22579
rect 758 22523 836 22579
rect 219 22498 836 22523
rect 219 22442 242 22498
rect 298 22442 334 22498
rect 390 22442 426 22498
rect 482 22442 518 22498
rect 574 22442 610 22498
rect 666 22442 702 22498
rect 758 22442 836 22498
rect 219 22417 836 22442
rect 219 22361 242 22417
rect 298 22361 334 22417
rect 390 22361 426 22417
rect 482 22361 518 22417
rect 574 22361 610 22417
rect 666 22361 702 22417
rect 758 22361 836 22417
rect 219 22336 836 22361
rect 219 22280 242 22336
rect 298 22280 334 22336
rect 390 22280 426 22336
rect 482 22280 518 22336
rect 574 22280 610 22336
rect 666 22280 702 22336
rect 758 22280 836 22336
rect 219 22255 836 22280
rect 219 22199 242 22255
rect 298 22199 334 22255
rect 390 22199 426 22255
rect 482 22199 518 22255
rect 574 22199 610 22255
rect 666 22199 702 22255
rect 758 22199 836 22255
rect 219 22174 836 22199
rect 219 22118 242 22174
rect 298 22118 334 22174
rect 390 22118 426 22174
rect 482 22118 518 22174
rect 574 22118 610 22174
rect 666 22118 702 22174
rect 758 22118 836 22174
rect 219 22093 836 22118
rect 219 22037 242 22093
rect 298 22037 334 22093
rect 390 22037 426 22093
rect 482 22037 518 22093
rect 574 22037 610 22093
rect 666 22037 702 22093
rect 758 22037 836 22093
rect 219 22012 836 22037
rect 219 21956 242 22012
rect 298 21956 334 22012
rect 390 21956 426 22012
rect 482 21956 518 22012
rect 574 21956 610 22012
rect 666 21956 702 22012
rect 758 21956 836 22012
rect 219 21931 836 21956
rect 219 21875 242 21931
rect 298 21875 334 21931
rect 390 21875 426 21931
rect 482 21875 518 21931
rect 574 21875 610 21931
rect 666 21875 702 21931
rect 758 21875 836 21931
rect 219 21850 836 21875
rect 219 21794 242 21850
rect 298 21794 334 21850
rect 390 21794 426 21850
rect 482 21794 518 21850
rect 574 21794 610 21850
rect 666 21794 702 21850
rect 758 21794 836 21850
rect 219 21769 836 21794
rect 219 21713 242 21769
rect 298 21713 334 21769
rect 390 21713 426 21769
rect 482 21713 518 21769
rect 574 21713 610 21769
rect 666 21713 702 21769
rect 758 21713 836 21769
rect 219 21688 836 21713
rect 219 21632 242 21688
rect 298 21632 334 21688
rect 390 21632 426 21688
rect 482 21632 518 21688
rect 574 21632 610 21688
rect 666 21632 702 21688
rect 758 21632 836 21688
rect 219 21607 836 21632
rect 219 21551 242 21607
rect 298 21551 334 21607
rect 390 21551 426 21607
rect 482 21551 518 21607
rect 574 21551 610 21607
rect 666 21551 702 21607
rect 758 21551 836 21607
rect 219 21526 836 21551
rect 219 21470 242 21526
rect 298 21470 334 21526
rect 390 21470 426 21526
rect 482 21470 518 21526
rect 574 21470 610 21526
rect 666 21470 702 21526
rect 758 21470 836 21526
rect 219 21445 836 21470
rect 219 21389 242 21445
rect 298 21389 334 21445
rect 390 21389 426 21445
rect 482 21389 518 21445
rect 574 21389 610 21445
rect 666 21389 702 21445
rect 758 21389 836 21445
rect 219 21364 836 21389
rect 219 21308 242 21364
rect 298 21308 334 21364
rect 390 21308 426 21364
rect 482 21308 518 21364
rect 574 21308 610 21364
rect 666 21308 702 21364
rect 758 21308 836 21364
rect 219 21283 836 21308
rect 219 21227 242 21283
rect 298 21227 334 21283
rect 390 21227 426 21283
rect 482 21227 518 21283
rect 574 21227 610 21283
rect 666 21227 702 21283
rect 758 21227 836 21283
rect 219 21202 836 21227
rect 219 21146 242 21202
rect 298 21146 334 21202
rect 390 21146 426 21202
rect 482 21146 518 21202
rect 574 21146 610 21202
rect 666 21146 702 21202
rect 758 21146 836 21202
rect 219 21121 836 21146
rect 1004 23686 1172 23691
rect 1004 23621 1009 23686
rect 1065 23685 1111 23686
rect 1073 23621 1103 23685
rect 1167 23621 1172 23686
rect 1004 23606 1172 23621
rect 1004 23540 1009 23606
rect 1065 23604 1111 23606
rect 1073 23540 1103 23604
rect 1167 23540 1172 23606
rect 1004 23526 1172 23540
rect 1004 23458 1009 23526
rect 1065 23522 1111 23526
rect 1073 23458 1103 23522
rect 1167 23458 1172 23526
rect 1004 23446 1172 23458
rect 1004 23376 1009 23446
rect 1065 23440 1111 23446
rect 1073 23376 1103 23440
rect 1167 23376 1172 23446
rect 1004 23366 1172 23376
rect 1004 23294 1009 23366
rect 1065 23358 1111 23366
rect 1073 23294 1103 23358
rect 1167 23294 1172 23366
rect 1004 23286 1172 23294
rect 1004 23212 1009 23286
rect 1065 23276 1111 23286
rect 1073 23212 1103 23276
rect 1167 23212 1172 23286
rect 1004 23206 1172 23212
rect 1004 23130 1009 23206
rect 1065 23194 1111 23206
rect 1073 23130 1103 23194
rect 1167 23130 1172 23206
rect 1004 23126 1172 23130
rect 1004 23048 1009 23126
rect 1065 23112 1111 23126
rect 1073 23048 1103 23112
rect 1167 23048 1172 23126
rect 1004 23046 1172 23048
rect 1004 21784 1009 23046
rect 1065 23030 1111 23046
rect 1073 22966 1103 23030
rect 1065 22948 1111 22966
rect 1073 22884 1103 22948
rect 1065 22866 1111 22884
rect 1073 22802 1103 22866
rect 1065 22784 1111 22802
rect 1073 22720 1103 22784
rect 1065 22702 1111 22720
rect 1073 22638 1103 22702
rect 1065 22620 1111 22638
rect 1073 22556 1103 22620
rect 1065 22538 1111 22556
rect 1073 22474 1103 22538
rect 1065 22456 1111 22474
rect 1073 22392 1103 22456
rect 1065 22374 1111 22392
rect 1073 22310 1103 22374
rect 1065 22292 1111 22310
rect 1073 22228 1103 22292
rect 1065 22210 1111 22228
rect 1073 22146 1103 22210
rect 1065 22128 1111 22146
rect 1073 22064 1103 22128
rect 1065 22046 1111 22064
rect 1073 21982 1103 22046
rect 1065 21964 1111 21982
rect 1073 21900 1103 21964
rect 1065 21882 1111 21900
rect 1073 21818 1103 21882
rect 1065 21784 1111 21818
rect 1167 21784 1172 23046
rect 1004 21759 1172 21784
rect 1004 21703 1009 21759
rect 1065 21703 1111 21759
rect 1167 21703 1172 21759
rect 1004 21678 1172 21703
rect 1004 21622 1009 21678
rect 1065 21622 1111 21678
rect 1167 21622 1172 21678
rect 1004 21597 1172 21622
rect 1004 21541 1009 21597
rect 1065 21541 1111 21597
rect 1167 21541 1172 21597
rect 1004 21516 1172 21541
rect 1004 21460 1009 21516
rect 1065 21460 1111 21516
rect 1167 21460 1172 21516
rect 1004 21435 1172 21460
rect 1004 21379 1009 21435
rect 1065 21379 1111 21435
rect 1167 21379 1172 21435
rect 1004 21354 1172 21379
rect 1004 21298 1009 21354
rect 1065 21298 1111 21354
rect 1167 21298 1172 21354
rect 1004 21273 1172 21298
rect 1004 21217 1009 21273
rect 1065 21217 1111 21273
rect 1167 21217 1172 21273
rect 1004 21192 1172 21217
rect 1004 21136 1009 21192
rect 1065 21136 1111 21192
rect 1167 21136 1172 21192
rect 1004 21131 1172 21136
rect 1488 23686 1680 23721
rect 1488 23630 1497 23686
rect 1553 23630 1615 23686
rect 1671 23630 1680 23686
rect 1488 23606 1680 23630
rect 1488 23550 1497 23606
rect 1553 23550 1615 23606
rect 1671 23550 1680 23606
rect 1488 23526 1680 23550
rect 1488 23470 1497 23526
rect 1553 23470 1615 23526
rect 1671 23470 1680 23526
rect 1488 23446 1680 23470
rect 1488 23390 1497 23446
rect 1553 23390 1615 23446
rect 1671 23390 1680 23446
rect 1488 23366 1680 23390
rect 1488 23310 1497 23366
rect 1553 23310 1615 23366
rect 1671 23310 1680 23366
rect 1488 23286 1680 23310
rect 1488 23230 1497 23286
rect 1553 23230 1615 23286
rect 1671 23230 1680 23286
rect 1488 23206 1680 23230
rect 1488 23150 1497 23206
rect 1553 23150 1615 23206
rect 1671 23150 1680 23206
rect 1488 23126 1680 23150
rect 1488 23070 1497 23126
rect 1553 23070 1615 23126
rect 1671 23070 1680 23126
rect 1488 23046 1680 23070
rect 1488 22990 1497 23046
rect 1553 22990 1615 23046
rect 1671 22990 1680 23046
rect 1488 22966 1680 22990
rect 1488 22910 1497 22966
rect 1553 22910 1615 22966
rect 1671 22910 1680 22966
rect 1488 22886 1680 22910
rect 1488 22830 1497 22886
rect 1553 22830 1615 22886
rect 1671 22830 1680 22886
rect 1488 22806 1680 22830
rect 1488 22750 1497 22806
rect 1553 22750 1615 22806
rect 1671 22750 1680 22806
rect 1488 22726 1680 22750
rect 1488 22670 1497 22726
rect 1553 22670 1615 22726
rect 1671 22670 1680 22726
rect 1488 22646 1680 22670
rect 1488 22590 1497 22646
rect 1553 22590 1615 22646
rect 1671 22590 1680 22646
rect 1488 22566 1680 22590
rect 1488 22510 1497 22566
rect 1553 22510 1615 22566
rect 1671 22510 1680 22566
rect 1488 22486 1680 22510
rect 1488 22430 1497 22486
rect 1553 22430 1615 22486
rect 1671 22430 1680 22486
rect 1488 22406 1680 22430
rect 1488 22350 1497 22406
rect 1553 22350 1615 22406
rect 1671 22350 1680 22406
rect 1488 22326 1680 22350
rect 1488 22270 1497 22326
rect 1553 22270 1615 22326
rect 1671 22270 1680 22326
rect 1488 22245 1680 22270
rect 1488 22189 1497 22245
rect 1553 22189 1615 22245
rect 1671 22189 1680 22245
rect 1488 22164 1680 22189
rect 1488 22108 1497 22164
rect 1553 22108 1615 22164
rect 1671 22108 1680 22164
rect 1488 22083 1680 22108
rect 1488 22027 1497 22083
rect 1553 22027 1615 22083
rect 1671 22027 1680 22083
rect 1488 22002 1680 22027
rect 1488 21946 1497 22002
rect 1553 21946 1615 22002
rect 1671 21946 1680 22002
rect 1488 21921 1680 21946
rect 1488 21865 1497 21921
rect 1553 21865 1615 21921
rect 1671 21865 1680 21921
rect 1488 21840 1680 21865
rect 1488 21784 1497 21840
rect 1553 21784 1615 21840
rect 1671 21784 1680 21840
rect 1488 21759 1680 21784
rect 1488 21703 1497 21759
rect 1553 21703 1615 21759
rect 1671 21703 1680 21759
rect 1488 21678 1680 21703
rect 1488 21622 1497 21678
rect 1553 21622 1615 21678
rect 1671 21622 1680 21678
rect 1488 21597 1680 21622
rect 1488 21541 1497 21597
rect 1553 21541 1615 21597
rect 1671 21541 1680 21597
rect 1488 21516 1680 21541
rect 1488 21460 1497 21516
rect 1553 21460 1615 21516
rect 1671 21460 1680 21516
rect 1488 21435 1680 21460
rect 1488 21379 1497 21435
rect 1553 21379 1615 21435
rect 1671 21379 1680 21435
rect 1488 21354 1680 21379
rect 1488 21298 1497 21354
rect 1553 21298 1615 21354
rect 1671 21298 1680 21354
rect 1488 21273 1680 21298
rect 1488 21217 1497 21273
rect 1553 21217 1615 21273
rect 1671 21217 1680 21273
rect 1488 21192 1680 21217
rect 1488 21136 1497 21192
rect 1553 21136 1615 21192
rect 1671 21136 1680 21192
rect 219 21065 242 21121
rect 298 21065 334 21121
rect 390 21065 426 21121
rect 482 21065 518 21121
rect 574 21065 610 21121
rect 666 21065 702 21121
rect 758 21065 836 21121
rect 219 21040 836 21065
rect 219 20984 242 21040
rect 298 20984 334 21040
rect 390 20984 426 21040
rect 482 20984 518 21040
rect 574 20984 610 21040
rect 666 20984 702 21040
rect 758 20984 836 21040
rect 219 20959 836 20984
rect 219 20903 242 20959
rect 298 20903 334 20959
rect 390 20903 426 20959
rect 482 20903 518 20959
rect 574 20903 610 20959
rect 666 20903 702 20959
rect 758 20903 836 20959
rect 219 20878 836 20903
rect 219 20822 242 20878
rect 298 20822 334 20878
rect 390 20822 426 20878
rect 482 20822 518 20878
rect 574 20822 610 20878
rect 666 20822 702 20878
rect 758 20822 836 20878
rect 219 20797 836 20822
rect 219 20741 242 20797
rect 298 20741 334 20797
rect 390 20741 426 20797
rect 482 20741 518 20797
rect 574 20741 610 20797
rect 666 20741 702 20797
rect 758 20741 836 20797
rect 219 20716 836 20741
rect 219 20660 242 20716
rect 298 20660 334 20716
rect 390 20660 426 20716
rect 482 20660 518 20716
rect 574 20660 610 20716
rect 666 20660 702 20716
rect 758 20660 836 20716
rect 219 20635 836 20660
rect 219 20579 242 20635
rect 298 20579 334 20635
rect 390 20579 426 20635
rect 482 20579 518 20635
rect 574 20579 610 20635
rect 666 20579 702 20635
rect 758 20607 836 20635
tri 836 20607 853 20624 sw
rect 758 20582 853 20607
tri 853 20582 878 20607 sw
rect 758 20579 878 20582
rect 219 20554 878 20579
rect 219 20498 242 20554
rect 298 20498 334 20554
rect 390 20498 426 20554
rect 482 20498 518 20554
rect 574 20498 610 20554
rect 666 20498 702 20554
rect 758 20531 878 20554
tri 878 20531 929 20582 sw
rect 758 20526 929 20531
tri 929 20526 934 20531 sw
rect 758 20498 934 20526
rect 219 20473 934 20498
rect 219 20417 242 20473
rect 298 20417 334 20473
rect 390 20417 426 20473
rect 482 20417 518 20473
rect 574 20417 610 20473
rect 666 20417 702 20473
rect 758 20417 934 20473
rect 219 20412 934 20417
tri 934 20412 1048 20526 sw
rect 219 20293 1048 20412
tri 1048 20293 1167 20412 sw
rect 219 20131 1167 20293
tri 219 19902 448 20131 ne
rect 448 18588 1167 20131
tri 1484 19923 1488 19927 se
rect 1488 19923 1680 21136
rect 1982 23686 2172 23903
rect 1982 23630 1993 23686
rect 2049 23630 2111 23686
rect 2167 23630 2172 23686
rect 1982 23606 2172 23630
rect 1982 23550 1993 23606
rect 2049 23550 2111 23606
rect 2167 23550 2172 23606
rect 1982 23526 2172 23550
rect 1982 23470 1993 23526
rect 2049 23470 2111 23526
rect 2167 23470 2172 23526
rect 1982 23446 2172 23470
rect 1982 23390 1993 23446
rect 2049 23390 2111 23446
rect 2167 23390 2172 23446
rect 1982 23366 2172 23390
rect 1982 23310 1993 23366
rect 2049 23310 2111 23366
rect 2167 23310 2172 23366
rect 1982 23286 2172 23310
rect 1982 23230 1993 23286
rect 2049 23230 2111 23286
rect 2167 23230 2172 23286
rect 1982 23206 2172 23230
rect 1982 23150 1993 23206
rect 2049 23150 2111 23206
rect 2167 23150 2172 23206
rect 1982 23126 2172 23150
rect 1982 23070 1993 23126
rect 2049 23070 2111 23126
rect 2167 23070 2172 23126
rect 1982 23046 2172 23070
rect 1982 22990 1993 23046
rect 2049 22990 2111 23046
rect 2167 22990 2172 23046
rect 1982 22966 2172 22990
rect 1982 22910 1993 22966
rect 2049 22910 2111 22966
rect 2167 22910 2172 22966
rect 1982 22886 2172 22910
rect 1982 22830 1993 22886
rect 2049 22830 2111 22886
rect 2167 22830 2172 22886
rect 1982 22806 2172 22830
rect 1982 22750 1993 22806
rect 2049 22750 2111 22806
rect 2167 22750 2172 22806
rect 1982 22726 2172 22750
rect 1982 22670 1993 22726
rect 2049 22670 2111 22726
rect 2167 22670 2172 22726
rect 1982 22646 2172 22670
rect 1982 22590 1993 22646
rect 2049 22590 2111 22646
rect 2167 22590 2172 22646
rect 1982 22566 2172 22590
rect 1982 22510 1993 22566
rect 2049 22510 2111 22566
rect 2167 22510 2172 22566
rect 1982 22486 2172 22510
rect 1982 22430 1993 22486
rect 2049 22430 2111 22486
rect 2167 22430 2172 22486
rect 1982 22406 2172 22430
rect 1982 22350 1993 22406
rect 2049 22350 2111 22406
rect 2167 22350 2172 22406
rect 1982 22326 2172 22350
rect 1982 22270 1993 22326
rect 2049 22270 2111 22326
rect 2167 22270 2172 22326
rect 1982 22245 2172 22270
rect 1982 22189 1993 22245
rect 2049 22189 2111 22245
rect 2167 22189 2172 22245
rect 1982 22164 2172 22189
rect 1982 22108 1993 22164
rect 2049 22108 2111 22164
rect 2167 22108 2172 22164
rect 1982 22083 2172 22108
rect 1982 22027 1993 22083
rect 2049 22027 2111 22083
rect 2167 22027 2172 22083
rect 1982 22002 2172 22027
rect 1982 21946 1993 22002
rect 2049 21946 2111 22002
rect 2167 21946 2172 22002
rect 1982 21921 2172 21946
rect 1982 21865 1993 21921
rect 2049 21865 2111 21921
rect 2167 21865 2172 21921
rect 1982 21840 2172 21865
rect 1982 21784 1993 21840
rect 2049 21784 2111 21840
rect 2167 21784 2172 21840
rect 1982 21759 2172 21784
rect 1982 21703 1993 21759
rect 2049 21703 2111 21759
rect 2167 21703 2172 21759
rect 1982 21678 2172 21703
rect 1982 21622 1993 21678
rect 2049 21622 2111 21678
rect 2167 21622 2172 21678
rect 1982 21597 2172 21622
rect 1982 21541 1993 21597
rect 2049 21541 2111 21597
rect 2167 21541 2172 21597
rect 1982 21516 2172 21541
rect 1982 21460 1993 21516
rect 2049 21460 2111 21516
rect 2167 21460 2172 21516
rect 1982 21435 2172 21460
rect 1982 21379 1993 21435
rect 2049 21379 2111 21435
rect 2167 21379 2172 21435
rect 1982 21354 2172 21379
rect 1982 21298 1993 21354
rect 2049 21298 2111 21354
rect 2167 21298 2172 21354
rect 1982 21273 2172 21298
rect 1982 21217 1993 21273
rect 2049 21217 2111 21273
rect 2167 21217 2172 21273
rect 1982 21192 2172 21217
rect 1982 21136 1993 21192
rect 2049 21136 2111 21192
rect 2167 21136 2172 21192
rect 1982 19990 2172 21136
rect 1982 19926 1986 19990
rect 2050 19926 2102 19990
rect 2166 19926 2172 19990
rect 448 15484 456 18588
rect 1160 15484 1167 18588
rect 448 15467 1167 15484
rect 448 15403 456 15467
rect 520 15403 536 15467
rect 600 15403 616 15467
rect 680 15403 696 15467
rect 760 15403 776 15467
rect 840 15403 856 15467
rect 920 15403 936 15467
rect 1000 15403 1016 15467
rect 1080 15403 1096 15467
rect 1160 15403 1167 15467
rect 448 15386 1167 15403
rect 448 15322 456 15386
rect 520 15322 536 15386
rect 600 15322 616 15386
rect 680 15322 696 15386
rect 760 15322 776 15386
rect 840 15322 856 15386
rect 920 15322 936 15386
rect 1000 15322 1016 15386
rect 1080 15322 1096 15386
rect 1160 15322 1167 15386
rect 448 15305 1167 15322
rect 448 15241 456 15305
rect 520 15241 536 15305
rect 600 15241 616 15305
rect 680 15241 696 15305
rect 760 15241 776 15305
rect 840 15241 856 15305
rect 920 15241 936 15305
rect 1000 15241 1016 15305
rect 1080 15241 1096 15305
rect 1160 15241 1167 15305
rect 448 15224 1167 15241
rect 448 15160 456 15224
rect 520 15160 536 15224
rect 600 15160 616 15224
rect 680 15160 696 15224
rect 760 15160 776 15224
rect 840 15160 856 15224
rect 920 15160 936 15224
rect 1000 15160 1016 15224
rect 1080 15160 1096 15224
rect 1160 15160 1167 15224
rect 448 15143 1167 15160
rect 448 15079 456 15143
rect 520 15079 536 15143
rect 600 15079 616 15143
rect 680 15079 696 15143
rect 760 15079 776 15143
rect 840 15079 856 15143
rect 920 15079 936 15143
rect 1000 15079 1016 15143
rect 1080 15079 1096 15143
rect 1160 15079 1167 15143
rect 448 15062 1167 15079
rect 448 14998 456 15062
rect 520 14998 536 15062
rect 600 14998 616 15062
rect 680 14998 696 15062
rect 760 14998 776 15062
rect 840 14998 856 15062
rect 920 14998 936 15062
rect 1000 14998 1016 15062
rect 1080 14998 1096 15062
rect 1160 14998 1167 15062
rect 448 14981 1167 14998
rect 448 14917 456 14981
rect 520 14917 536 14981
rect 600 14917 616 14981
rect 680 14917 696 14981
rect 760 14917 776 14981
rect 840 14917 856 14981
rect 920 14917 936 14981
rect 1000 14917 1016 14981
rect 1080 14917 1096 14981
rect 1160 14917 1167 14981
rect 448 14900 1167 14917
rect 448 14836 456 14900
rect 520 14836 536 14900
rect 600 14836 616 14900
rect 680 14836 696 14900
rect 760 14836 776 14900
rect 840 14836 856 14900
rect 920 14836 936 14900
rect 1000 14836 1016 14900
rect 1080 14836 1096 14900
rect 1160 14836 1167 14900
rect 448 14819 1167 14836
rect 448 14755 456 14819
rect 520 14755 536 14819
rect 600 14755 616 14819
rect 680 14755 696 14819
rect 760 14755 776 14819
rect 840 14755 856 14819
rect 920 14755 936 14819
rect 1000 14755 1016 14819
rect 1080 14755 1096 14819
rect 1160 14755 1167 14819
rect 448 14738 1167 14755
rect 448 14674 456 14738
rect 520 14674 536 14738
rect 600 14674 616 14738
rect 680 14674 696 14738
rect 760 14674 776 14738
rect 840 14674 856 14738
rect 920 14674 936 14738
rect 1000 14674 1016 14738
rect 1080 14674 1096 14738
rect 1160 14674 1167 14738
rect 448 14657 1167 14674
rect 448 14593 456 14657
rect 520 14593 536 14657
rect 600 14593 616 14657
rect 680 14593 696 14657
rect 760 14593 776 14657
rect 840 14593 856 14657
rect 920 14593 936 14657
rect 1000 14593 1016 14657
rect 1080 14593 1096 14657
rect 1160 14593 1167 14657
rect 448 14576 1167 14593
rect 448 14512 456 14576
rect 520 14512 536 14576
rect 600 14512 616 14576
rect 680 14512 696 14576
rect 760 14512 776 14576
rect 840 14512 856 14576
rect 920 14512 936 14576
rect 1000 14512 1016 14576
rect 1080 14512 1096 14576
rect 1160 14512 1167 14576
rect 448 14495 1167 14512
rect 448 14431 456 14495
rect 520 14431 536 14495
rect 600 14431 616 14495
rect 680 14431 696 14495
rect 760 14431 776 14495
rect 840 14431 856 14495
rect 920 14431 936 14495
rect 1000 14431 1016 14495
rect 1080 14431 1096 14495
rect 1160 14431 1167 14495
rect 448 14414 1167 14431
rect 448 14350 456 14414
rect 520 14350 536 14414
rect 600 14350 616 14414
rect 680 14350 696 14414
rect 760 14350 776 14414
rect 840 14350 856 14414
rect 920 14350 936 14414
rect 1000 14350 1016 14414
rect 1080 14350 1096 14414
rect 1160 14350 1167 14414
rect 448 14333 1167 14350
rect 448 14269 456 14333
rect 520 14269 536 14333
rect 600 14269 616 14333
rect 680 14269 696 14333
rect 760 14269 776 14333
rect 840 14269 856 14333
rect 920 14269 936 14333
rect 1000 14269 1016 14333
rect 1080 14269 1096 14333
rect 1160 14269 1167 14333
rect 448 14252 1167 14269
rect 448 14188 456 14252
rect 520 14188 536 14252
rect 600 14188 616 14252
rect 680 14188 696 14252
rect 760 14188 776 14252
rect 840 14188 856 14252
rect 920 14188 936 14252
rect 1000 14188 1016 14252
rect 1080 14188 1096 14252
rect 1160 14188 1167 14252
rect 448 14171 1167 14188
rect 448 14107 456 14171
rect 520 14107 536 14171
rect 600 14107 616 14171
rect 680 14107 696 14171
rect 760 14107 776 14171
rect 840 14107 856 14171
rect 920 14107 936 14171
rect 1000 14107 1016 14171
rect 1080 14107 1096 14171
rect 1160 14107 1167 14171
rect 448 14090 1167 14107
rect 448 14026 456 14090
rect 520 14026 536 14090
rect 600 14026 616 14090
rect 680 14026 696 14090
rect 760 14026 776 14090
rect 840 14026 856 14090
rect 920 14026 936 14090
rect 1000 14026 1016 14090
rect 1080 14026 1096 14090
rect 1160 14026 1167 14090
rect 448 14009 1167 14026
rect 448 13945 456 14009
rect 520 13945 536 14009
rect 600 13945 616 14009
rect 680 13945 696 14009
rect 760 13945 776 14009
rect 840 13945 856 14009
rect 920 13945 936 14009
rect 1000 13945 1016 14009
rect 1080 13945 1096 14009
rect 1160 13945 1167 14009
rect 448 13928 1167 13945
rect 448 13864 456 13928
rect 520 13864 536 13928
rect 600 13864 616 13928
rect 680 13864 696 13928
rect 760 13864 776 13928
rect 840 13864 856 13928
rect 920 13864 936 13928
rect 1000 13864 1016 13928
rect 1080 13864 1096 13928
rect 1160 13864 1167 13928
rect 448 13847 1167 13864
rect 448 13783 456 13847
rect 520 13783 536 13847
rect 600 13783 616 13847
rect 680 13783 696 13847
rect 760 13783 776 13847
rect 840 13783 856 13847
rect 920 13783 936 13847
rect 1000 13783 1016 13847
rect 1080 13783 1096 13847
rect 1160 13783 1167 13847
rect 448 13766 1167 13783
rect 448 13702 456 13766
rect 520 13702 536 13766
rect 600 13702 616 13766
rect 680 13702 696 13766
rect 760 13702 776 13766
rect 840 13702 856 13766
rect 920 13702 936 13766
rect 1000 13702 1016 13766
rect 1080 13702 1096 13766
rect 1160 13702 1167 13766
rect 448 13685 1167 13702
rect 448 13621 456 13685
rect 520 13621 536 13685
rect 600 13621 616 13685
rect 680 13621 696 13685
rect 760 13621 776 13685
rect 840 13621 856 13685
rect 920 13621 936 13685
rect 1000 13621 1016 13685
rect 1080 13621 1096 13685
rect 1160 13621 1167 13685
rect 448 13607 1167 13621
tri 1275 19714 1484 19923 se
rect 1484 19714 1680 19923
tri 1680 19714 1889 19923 sw
rect 1275 18586 1889 19714
rect 1275 18522 1287 18586
rect 1351 18522 1375 18586
rect 1439 18522 1463 18586
rect 1527 18522 1551 18586
rect 1615 18522 1639 18586
rect 1703 18522 1727 18586
rect 1791 18522 1815 18586
rect 1879 18522 1889 18586
rect 1275 18506 1889 18522
rect 1275 18442 1287 18506
rect 1351 18442 1375 18506
rect 1439 18442 1463 18506
rect 1527 18442 1551 18506
rect 1615 18442 1639 18506
rect 1703 18442 1727 18506
rect 1791 18442 1815 18506
rect 1879 18442 1889 18506
rect 1275 18426 1889 18442
rect 1275 18362 1287 18426
rect 1351 18362 1375 18426
rect 1439 18362 1463 18426
rect 1527 18362 1551 18426
rect 1615 18362 1639 18426
rect 1703 18362 1727 18426
rect 1791 18362 1815 18426
rect 1879 18362 1889 18426
rect 1275 18346 1889 18362
rect 1275 18282 1287 18346
rect 1351 18282 1375 18346
rect 1439 18282 1463 18346
rect 1527 18282 1551 18346
rect 1615 18282 1639 18346
rect 1703 18282 1727 18346
rect 1791 18282 1815 18346
rect 1879 18282 1889 18346
rect 1275 18266 1889 18282
rect 1275 18202 1287 18266
rect 1351 18202 1375 18266
rect 1439 18202 1463 18266
rect 1527 18202 1551 18266
rect 1615 18202 1639 18266
rect 1703 18202 1727 18266
rect 1791 18202 1815 18266
rect 1879 18202 1889 18266
rect 1275 18186 1889 18202
rect 1275 18122 1287 18186
rect 1351 18122 1375 18186
rect 1439 18122 1463 18186
rect 1527 18122 1551 18186
rect 1615 18122 1639 18186
rect 1703 18122 1727 18186
rect 1791 18122 1815 18186
rect 1879 18122 1889 18186
rect 1275 18106 1889 18122
rect 1275 18042 1287 18106
rect 1351 18042 1375 18106
rect 1439 18042 1463 18106
rect 1527 18042 1551 18106
rect 1615 18042 1639 18106
rect 1703 18042 1727 18106
rect 1791 18042 1815 18106
rect 1879 18042 1889 18106
rect 1275 18026 1889 18042
rect 1275 17962 1287 18026
rect 1351 17962 1375 18026
rect 1439 17962 1463 18026
rect 1527 17962 1551 18026
rect 1615 17962 1639 18026
rect 1703 17962 1727 18026
rect 1791 17962 1815 18026
rect 1879 17962 1889 18026
rect 1275 17946 1889 17962
rect 1275 17882 1287 17946
rect 1351 17882 1375 17946
rect 1439 17882 1463 17946
rect 1527 17882 1551 17946
rect 1615 17882 1639 17946
rect 1703 17882 1727 17946
rect 1791 17882 1815 17946
rect 1879 17882 1889 17946
rect 1275 17866 1889 17882
rect 1275 17802 1287 17866
rect 1351 17802 1375 17866
rect 1439 17802 1463 17866
rect 1527 17802 1551 17866
rect 1615 17802 1639 17866
rect 1703 17802 1727 17866
rect 1791 17802 1815 17866
rect 1879 17802 1889 17866
rect 1275 17786 1889 17802
rect 1275 17722 1287 17786
rect 1351 17722 1375 17786
rect 1439 17722 1463 17786
rect 1527 17722 1551 17786
rect 1615 17722 1639 17786
rect 1703 17722 1727 17786
rect 1791 17722 1815 17786
rect 1879 17722 1889 17786
rect 1275 17706 1889 17722
rect 1275 17642 1287 17706
rect 1351 17642 1375 17706
rect 1439 17642 1463 17706
rect 1527 17642 1551 17706
rect 1615 17642 1639 17706
rect 1703 17642 1727 17706
rect 1791 17642 1815 17706
rect 1879 17642 1889 17706
rect 1275 17626 1889 17642
rect 1275 17562 1287 17626
rect 1351 17562 1375 17626
rect 1439 17562 1463 17626
rect 1527 17562 1551 17626
rect 1615 17562 1639 17626
rect 1703 17562 1727 17626
rect 1791 17562 1815 17626
rect 1879 17562 1889 17626
rect 1275 17546 1889 17562
rect 1275 17482 1287 17546
rect 1351 17482 1375 17546
rect 1439 17482 1463 17546
rect 1527 17482 1551 17546
rect 1615 17482 1639 17546
rect 1703 17482 1727 17546
rect 1791 17482 1815 17546
rect 1879 17482 1889 17546
rect 1275 17466 1889 17482
rect 1275 17402 1287 17466
rect 1351 17402 1375 17466
rect 1439 17402 1463 17466
rect 1527 17402 1551 17466
rect 1615 17402 1639 17466
rect 1703 17402 1727 17466
rect 1791 17402 1815 17466
rect 1879 17402 1889 17466
rect 1275 17386 1889 17402
rect 1275 17322 1287 17386
rect 1351 17322 1375 17386
rect 1439 17322 1463 17386
rect 1527 17322 1551 17386
rect 1615 17322 1639 17386
rect 1703 17322 1727 17386
rect 1791 17322 1815 17386
rect 1879 17322 1889 17386
rect 1275 17306 1889 17322
rect 1275 17242 1287 17306
rect 1351 17242 1375 17306
rect 1439 17242 1463 17306
rect 1527 17242 1551 17306
rect 1615 17242 1639 17306
rect 1703 17242 1727 17306
rect 1791 17242 1815 17306
rect 1879 17242 1889 17306
rect 1275 17226 1889 17242
rect 1275 17162 1287 17226
rect 1351 17162 1375 17226
rect 1439 17162 1463 17226
rect 1527 17162 1551 17226
rect 1615 17162 1639 17226
rect 1703 17162 1727 17226
rect 1791 17162 1815 17226
rect 1879 17162 1889 17226
rect 1275 17146 1889 17162
rect 1275 17082 1287 17146
rect 1351 17082 1375 17146
rect 1439 17082 1463 17146
rect 1527 17082 1551 17146
rect 1615 17082 1639 17146
rect 1703 17082 1727 17146
rect 1791 17082 1815 17146
rect 1879 17082 1889 17146
rect 1275 17066 1889 17082
rect 1275 17002 1287 17066
rect 1351 17002 1375 17066
rect 1439 17002 1463 17066
rect 1527 17002 1551 17066
rect 1615 17002 1639 17066
rect 1703 17002 1727 17066
rect 1791 17002 1815 17066
rect 1879 17002 1889 17066
rect 1275 16986 1889 17002
rect 1275 16922 1287 16986
rect 1351 16922 1375 16986
rect 1439 16922 1463 16986
rect 1527 16922 1551 16986
rect 1615 16922 1639 16986
rect 1703 16922 1727 16986
rect 1791 16922 1815 16986
rect 1879 16922 1889 16986
rect 1275 16906 1889 16922
rect 1275 16842 1287 16906
rect 1351 16842 1375 16906
rect 1439 16842 1463 16906
rect 1527 16842 1551 16906
rect 1615 16842 1639 16906
rect 1703 16842 1727 16906
rect 1791 16842 1815 16906
rect 1879 16842 1889 16906
rect 1275 16826 1889 16842
rect 1275 16762 1287 16826
rect 1351 16762 1375 16826
rect 1439 16762 1463 16826
rect 1527 16762 1551 16826
rect 1615 16762 1639 16826
rect 1703 16762 1727 16826
rect 1791 16762 1815 16826
rect 1879 16762 1889 16826
rect 1275 16746 1889 16762
rect 1275 16682 1287 16746
rect 1351 16682 1375 16746
rect 1439 16682 1463 16746
rect 1527 16682 1551 16746
rect 1615 16682 1639 16746
rect 1703 16682 1727 16746
rect 1791 16682 1815 16746
rect 1879 16682 1889 16746
rect 1275 16666 1889 16682
rect 1275 16602 1287 16666
rect 1351 16602 1375 16666
rect 1439 16602 1463 16666
rect 1527 16602 1551 16666
rect 1615 16602 1639 16666
rect 1703 16602 1727 16666
rect 1791 16602 1815 16666
rect 1879 16602 1889 16666
rect 1275 16586 1889 16602
rect 1275 16522 1287 16586
rect 1351 16522 1375 16586
rect 1439 16522 1463 16586
rect 1527 16522 1551 16586
rect 1615 16522 1639 16586
rect 1703 16522 1727 16586
rect 1791 16522 1815 16586
rect 1879 16522 1889 16586
rect 1275 16506 1889 16522
rect 1275 16442 1287 16506
rect 1351 16442 1375 16506
rect 1439 16442 1463 16506
rect 1527 16442 1551 16506
rect 1615 16442 1639 16506
rect 1703 16442 1727 16506
rect 1791 16442 1815 16506
rect 1879 16442 1889 16506
rect 1275 16426 1889 16442
rect 1275 16362 1287 16426
rect 1351 16362 1375 16426
rect 1439 16362 1463 16426
rect 1527 16362 1551 16426
rect 1615 16362 1639 16426
rect 1703 16362 1727 16426
rect 1791 16362 1815 16426
rect 1879 16362 1889 16426
rect 1275 16346 1889 16362
rect 1275 16282 1287 16346
rect 1351 16282 1375 16346
rect 1439 16282 1463 16346
rect 1527 16282 1551 16346
rect 1615 16282 1639 16346
rect 1703 16282 1727 16346
rect 1791 16282 1815 16346
rect 1879 16282 1889 16346
rect 1275 16266 1889 16282
rect 1275 16202 1287 16266
rect 1351 16202 1375 16266
rect 1439 16202 1463 16266
rect 1527 16202 1551 16266
rect 1615 16202 1639 16266
rect 1703 16202 1727 16266
rect 1791 16202 1815 16266
rect 1879 16202 1889 16266
rect 1275 16186 1889 16202
rect 1275 16122 1287 16186
rect 1351 16122 1375 16186
rect 1439 16122 1463 16186
rect 1527 16122 1551 16186
rect 1615 16122 1639 16186
rect 1703 16122 1727 16186
rect 1791 16122 1815 16186
rect 1879 16122 1889 16186
rect 1275 16106 1889 16122
rect 1275 16042 1287 16106
rect 1351 16042 1375 16106
rect 1439 16042 1463 16106
rect 1527 16042 1551 16106
rect 1615 16042 1639 16106
rect 1703 16042 1727 16106
rect 1791 16042 1815 16106
rect 1879 16042 1889 16106
rect 1275 16026 1889 16042
rect 1275 15962 1287 16026
rect 1351 15962 1375 16026
rect 1439 15962 1463 16026
rect 1527 15962 1551 16026
rect 1615 15962 1639 16026
rect 1703 15962 1727 16026
rect 1791 15962 1815 16026
rect 1879 15962 1889 16026
rect 1275 15946 1889 15962
rect 1275 15882 1287 15946
rect 1351 15882 1375 15946
rect 1439 15882 1463 15946
rect 1527 15882 1551 15946
rect 1615 15882 1639 15946
rect 1703 15882 1727 15946
rect 1791 15882 1815 15946
rect 1879 15882 1889 15946
rect 1275 15866 1889 15882
rect 1275 15802 1287 15866
rect 1351 15802 1375 15866
rect 1439 15802 1463 15866
rect 1527 15802 1551 15866
rect 1615 15802 1639 15866
rect 1703 15802 1727 15866
rect 1791 15802 1815 15866
rect 1879 15802 1889 15866
rect 1275 15786 1889 15802
rect 1275 15722 1287 15786
rect 1351 15722 1375 15786
rect 1439 15722 1463 15786
rect 1527 15722 1551 15786
rect 1615 15722 1639 15786
rect 1703 15722 1727 15786
rect 1791 15722 1815 15786
rect 1879 15722 1889 15786
rect 1275 15706 1889 15722
rect 1275 15642 1287 15706
rect 1351 15642 1375 15706
rect 1439 15642 1463 15706
rect 1527 15642 1551 15706
rect 1615 15642 1639 15706
rect 1703 15642 1727 15706
rect 1791 15642 1815 15706
rect 1879 15642 1889 15706
rect 1275 15626 1889 15642
rect 1275 15562 1287 15626
rect 1351 15562 1375 15626
rect 1439 15562 1463 15626
rect 1527 15562 1551 15626
rect 1615 15562 1639 15626
rect 1703 15562 1727 15626
rect 1791 15562 1815 15626
rect 1879 15562 1889 15626
rect 1275 15546 1889 15562
rect 1275 15482 1287 15546
rect 1351 15482 1375 15546
rect 1439 15482 1463 15546
rect 1527 15482 1551 15546
rect 1615 15482 1639 15546
rect 1703 15482 1727 15546
rect 1791 15482 1815 15546
rect 1879 15482 1889 15546
rect 1275 15466 1889 15482
rect 1275 15402 1287 15466
rect 1351 15402 1375 15466
rect 1439 15402 1463 15466
rect 1527 15402 1551 15466
rect 1615 15402 1639 15466
rect 1703 15402 1727 15466
rect 1791 15402 1815 15466
rect 1879 15402 1889 15466
rect 1275 15386 1889 15402
rect 1275 15322 1287 15386
rect 1351 15322 1375 15386
rect 1439 15322 1463 15386
rect 1527 15322 1551 15386
rect 1615 15322 1639 15386
rect 1703 15322 1727 15386
rect 1791 15322 1815 15386
rect 1879 15322 1889 15386
rect 1275 15306 1889 15322
rect 1275 15242 1287 15306
rect 1351 15242 1375 15306
rect 1439 15242 1463 15306
rect 1527 15242 1551 15306
rect 1615 15242 1639 15306
rect 1703 15242 1727 15306
rect 1791 15242 1815 15306
rect 1879 15242 1889 15306
rect 1275 15226 1889 15242
rect 1275 15162 1287 15226
rect 1351 15162 1375 15226
rect 1439 15162 1463 15226
rect 1527 15162 1551 15226
rect 1615 15162 1639 15226
rect 1703 15162 1727 15226
rect 1791 15162 1815 15226
rect 1879 15162 1889 15226
rect 1275 15146 1889 15162
rect 1275 15082 1287 15146
rect 1351 15082 1375 15146
rect 1439 15082 1463 15146
rect 1527 15082 1551 15146
rect 1615 15082 1639 15146
rect 1703 15082 1727 15146
rect 1791 15082 1815 15146
rect 1879 15082 1889 15146
rect 1275 15066 1889 15082
rect 1275 15002 1287 15066
rect 1351 15002 1375 15066
rect 1439 15002 1463 15066
rect 1527 15002 1551 15066
rect 1615 15002 1639 15066
rect 1703 15002 1727 15066
rect 1791 15002 1815 15066
rect 1879 15002 1889 15066
rect 1275 14986 1889 15002
rect 1275 14922 1287 14986
rect 1351 14922 1375 14986
rect 1439 14922 1463 14986
rect 1527 14922 1551 14986
rect 1615 14922 1639 14986
rect 1703 14922 1727 14986
rect 1791 14922 1815 14986
rect 1879 14922 1889 14986
rect 1275 14906 1889 14922
rect 1275 14842 1287 14906
rect 1351 14842 1375 14906
rect 1439 14842 1463 14906
rect 1527 14842 1551 14906
rect 1615 14842 1639 14906
rect 1703 14842 1727 14906
rect 1791 14842 1815 14906
rect 1879 14842 1889 14906
rect 1275 14826 1889 14842
rect 1275 14762 1287 14826
rect 1351 14762 1375 14826
rect 1439 14762 1463 14826
rect 1527 14762 1551 14826
rect 1615 14762 1639 14826
rect 1703 14762 1727 14826
rect 1791 14762 1815 14826
rect 1879 14762 1889 14826
rect 1275 14746 1889 14762
rect 1275 14682 1287 14746
rect 1351 14682 1375 14746
rect 1439 14682 1463 14746
rect 1527 14682 1551 14746
rect 1615 14682 1639 14746
rect 1703 14682 1727 14746
rect 1791 14682 1815 14746
rect 1879 14682 1889 14746
rect 1275 14666 1889 14682
rect 1275 14602 1287 14666
rect 1351 14602 1375 14666
rect 1439 14602 1463 14666
rect 1527 14602 1551 14666
rect 1615 14602 1639 14666
rect 1703 14602 1727 14666
rect 1791 14602 1815 14666
rect 1879 14602 1889 14666
rect 1275 14586 1889 14602
rect 1275 14522 1287 14586
rect 1351 14522 1375 14586
rect 1439 14522 1463 14586
rect 1527 14522 1551 14586
rect 1615 14522 1639 14586
rect 1703 14522 1727 14586
rect 1791 14522 1815 14586
rect 1879 14522 1889 14586
rect 1275 14505 1889 14522
rect 1275 14441 1287 14505
rect 1351 14441 1375 14505
rect 1439 14441 1463 14505
rect 1527 14441 1551 14505
rect 1615 14441 1639 14505
rect 1703 14441 1727 14505
rect 1791 14441 1815 14505
rect 1879 14441 1889 14505
rect 1275 14424 1889 14441
rect 1275 14360 1287 14424
rect 1351 14360 1375 14424
rect 1439 14360 1463 14424
rect 1527 14360 1551 14424
rect 1615 14360 1639 14424
rect 1703 14360 1727 14424
rect 1791 14360 1815 14424
rect 1879 14360 1889 14424
rect 1275 14343 1889 14360
rect 1275 14279 1287 14343
rect 1351 14279 1375 14343
rect 1439 14279 1463 14343
rect 1527 14279 1551 14343
rect 1615 14279 1639 14343
rect 1703 14279 1727 14343
rect 1791 14279 1815 14343
rect 1879 14279 1889 14343
rect 1275 14262 1889 14279
rect 1275 14198 1287 14262
rect 1351 14198 1375 14262
rect 1439 14198 1463 14262
rect 1527 14198 1551 14262
rect 1615 14198 1639 14262
rect 1703 14198 1727 14262
rect 1791 14198 1815 14262
rect 1879 14198 1889 14262
rect 1275 14181 1889 14198
rect 1275 14117 1287 14181
rect 1351 14117 1375 14181
rect 1439 14117 1463 14181
rect 1527 14117 1551 14181
rect 1615 14117 1639 14181
rect 1703 14117 1727 14181
rect 1791 14117 1815 14181
rect 1879 14117 1889 14181
rect 1275 14100 1889 14117
rect 1275 14036 1287 14100
rect 1351 14036 1375 14100
rect 1439 14036 1463 14100
rect 1527 14036 1551 14100
rect 1615 14036 1639 14100
rect 1703 14036 1727 14100
rect 1791 14036 1815 14100
rect 1879 14036 1889 14100
rect 1275 14019 1889 14036
rect 1275 13955 1287 14019
rect 1351 13955 1375 14019
rect 1439 13955 1463 14019
rect 1527 13955 1551 14019
rect 1615 13955 1639 14019
rect 1703 13955 1727 14019
rect 1791 13955 1815 14019
rect 1879 13955 1889 14019
rect 1275 13938 1889 13955
rect 1275 13874 1287 13938
rect 1351 13874 1375 13938
rect 1439 13874 1463 13938
rect 1527 13874 1551 13938
rect 1615 13874 1639 13938
rect 1703 13874 1727 13938
rect 1791 13874 1815 13938
rect 1879 13874 1889 13938
rect 1275 13857 1889 13874
rect 1275 13793 1287 13857
rect 1351 13793 1375 13857
rect 1439 13793 1463 13857
rect 1527 13793 1551 13857
rect 1615 13793 1639 13857
rect 1703 13793 1727 13857
rect 1791 13793 1815 13857
rect 1879 13793 1889 13857
rect 1275 13776 1889 13793
rect 1275 13712 1287 13776
rect 1351 13712 1375 13776
rect 1439 13712 1463 13776
rect 1527 13712 1551 13776
rect 1615 13712 1639 13776
rect 1703 13712 1727 13776
rect 1791 13712 1815 13776
rect 1879 13712 1889 13776
rect 1275 13695 1889 13712
rect 1275 13631 1287 13695
rect 1351 13631 1375 13695
rect 1439 13631 1463 13695
rect 1527 13631 1551 13695
rect 1615 13631 1639 13695
rect 1703 13631 1727 13695
rect 1791 13631 1815 13695
rect 1879 13631 1889 13695
rect 1275 13607 1889 13631
rect 1982 19907 2172 19926
rect 1982 19843 1986 19907
rect 2050 19843 2102 19907
rect 2166 19843 2172 19907
rect 1982 19823 2172 19843
rect 1982 19759 1986 19823
rect 2050 19759 2102 19823
rect 2166 19759 2172 19823
rect 1982 19739 2172 19759
rect 1982 19675 1986 19739
rect 2050 19675 2102 19739
rect 2166 19675 2172 19739
rect 1982 19655 2172 19675
rect 1982 19591 1986 19655
rect 2050 19591 2102 19655
rect 2166 19591 2172 19655
rect 1982 19571 2172 19591
rect 1982 19507 1986 19571
rect 2050 19507 2102 19571
rect 2166 19507 2172 19571
rect 1982 19487 2172 19507
rect 1982 19423 1986 19487
rect 2050 19423 2102 19487
rect 2166 19423 2172 19487
rect 1982 12887 2172 19423
rect 2480 23686 2672 25643
rect 2480 23630 2489 23686
rect 2545 23630 2607 23686
rect 2663 23630 2672 23686
rect 2480 23606 2672 23630
rect 2480 23550 2489 23606
rect 2545 23550 2607 23606
rect 2663 23550 2672 23606
rect 2480 23526 2672 23550
rect 2480 23470 2489 23526
rect 2545 23470 2607 23526
rect 2663 23470 2672 23526
rect 2480 23446 2672 23470
rect 2480 23390 2489 23446
rect 2545 23390 2607 23446
rect 2663 23390 2672 23446
rect 2480 23366 2672 23390
rect 2480 23310 2489 23366
rect 2545 23310 2607 23366
rect 2663 23310 2672 23366
rect 2480 23286 2672 23310
rect 2480 23230 2489 23286
rect 2545 23230 2607 23286
rect 2663 23230 2672 23286
rect 2480 23206 2672 23230
rect 2480 23150 2489 23206
rect 2545 23150 2607 23206
rect 2663 23150 2672 23206
rect 2480 23126 2672 23150
rect 2480 23070 2489 23126
rect 2545 23070 2607 23126
rect 2663 23070 2672 23126
rect 2480 23046 2672 23070
rect 2480 22990 2489 23046
rect 2545 22990 2607 23046
rect 2663 22990 2672 23046
rect 2480 22966 2672 22990
rect 2480 22910 2489 22966
rect 2545 22910 2607 22966
rect 2663 22910 2672 22966
rect 2480 22886 2672 22910
rect 2480 22830 2489 22886
rect 2545 22830 2607 22886
rect 2663 22830 2672 22886
rect 2480 22806 2672 22830
rect 2480 22750 2489 22806
rect 2545 22750 2607 22806
rect 2663 22750 2672 22806
rect 2480 22726 2672 22750
rect 2480 22670 2489 22726
rect 2545 22670 2607 22726
rect 2663 22670 2672 22726
rect 2480 22646 2672 22670
rect 2480 22590 2489 22646
rect 2545 22590 2607 22646
rect 2663 22590 2672 22646
rect 2480 22566 2672 22590
rect 2480 22510 2489 22566
rect 2545 22510 2607 22566
rect 2663 22510 2672 22566
rect 2480 22486 2672 22510
rect 2480 22430 2489 22486
rect 2545 22430 2607 22486
rect 2663 22430 2672 22486
rect 2480 22406 2672 22430
rect 2480 22350 2489 22406
rect 2545 22350 2607 22406
rect 2663 22350 2672 22406
rect 2480 22326 2672 22350
rect 2480 22270 2489 22326
rect 2545 22270 2607 22326
rect 2663 22270 2672 22326
rect 2480 22245 2672 22270
rect 2480 22189 2489 22245
rect 2545 22189 2607 22245
rect 2663 22189 2672 22245
rect 2480 22164 2672 22189
rect 2480 22108 2489 22164
rect 2545 22108 2607 22164
rect 2663 22108 2672 22164
rect 2480 22083 2672 22108
rect 2480 22027 2489 22083
rect 2545 22027 2607 22083
rect 2663 22027 2672 22083
rect 2480 22002 2672 22027
rect 2480 21946 2489 22002
rect 2545 21946 2607 22002
rect 2663 21946 2672 22002
rect 2480 21921 2672 21946
rect 2480 21865 2489 21921
rect 2545 21865 2607 21921
rect 2663 21865 2672 21921
rect 2480 21840 2672 21865
rect 2480 21784 2489 21840
rect 2545 21784 2607 21840
rect 2663 21784 2672 21840
rect 2480 21759 2672 21784
rect 2480 21703 2489 21759
rect 2545 21703 2607 21759
rect 2663 21703 2672 21759
rect 2480 21678 2672 21703
rect 2480 21622 2489 21678
rect 2545 21622 2607 21678
rect 2663 21622 2672 21678
rect 2480 21597 2672 21622
rect 2480 21541 2489 21597
rect 2545 21541 2607 21597
rect 2663 21541 2672 21597
rect 2480 21516 2672 21541
rect 2480 21460 2489 21516
rect 2545 21460 2607 21516
rect 2663 21460 2672 21516
rect 2480 21435 2672 21460
rect 2480 21379 2489 21435
rect 2545 21379 2607 21435
rect 2663 21379 2672 21435
rect 2480 21354 2672 21379
rect 2480 21298 2489 21354
rect 2545 21298 2607 21354
rect 2663 21298 2672 21354
rect 2480 21273 2672 21298
rect 2480 21217 2489 21273
rect 2545 21217 2607 21273
rect 2663 21217 2672 21273
rect 2480 21192 2672 21217
rect 2480 21136 2489 21192
rect 2545 21136 2607 21192
rect 2663 21136 2672 21192
rect 2480 18592 2672 21136
rect 2544 18528 2608 18592
rect 2480 18512 2672 18528
rect 2544 18448 2608 18512
rect 2480 18432 2672 18448
rect 2544 18368 2608 18432
rect 2480 18352 2672 18368
rect 2544 18288 2608 18352
rect 2480 18272 2672 18288
rect 2544 18208 2608 18272
rect 2480 18192 2672 18208
rect 2544 18128 2608 18192
rect 2480 18112 2672 18128
rect 2544 18048 2608 18112
rect 2480 18032 2672 18048
rect 2544 17968 2608 18032
rect 2480 17952 2672 17968
rect 2544 17888 2608 17952
rect 2480 17872 2672 17888
rect 2544 17808 2608 17872
rect 2480 17792 2672 17808
rect 2544 17728 2608 17792
rect 2480 17712 2672 17728
rect 2544 17648 2608 17712
rect 2480 17632 2672 17648
rect 2544 17568 2608 17632
rect 2480 17552 2672 17568
rect 2544 17488 2608 17552
rect 2480 17472 2672 17488
rect 2544 17408 2608 17472
rect 2480 17392 2672 17408
rect 2544 17328 2608 17392
rect 2480 17312 2672 17328
rect 2544 17248 2608 17312
rect 2480 17232 2672 17248
rect 2544 17168 2608 17232
rect 2480 17152 2672 17168
rect 2544 17088 2608 17152
rect 2480 17072 2672 17088
rect 2544 17008 2608 17072
rect 2480 16992 2672 17008
rect 2544 16928 2608 16992
rect 2480 16912 2672 16928
rect 2544 16848 2608 16912
rect 2480 16832 2672 16848
rect 2544 16768 2608 16832
rect 2480 16752 2672 16768
rect 2544 16688 2608 16752
rect 2480 16672 2672 16688
rect 2544 16608 2608 16672
rect 2480 16592 2672 16608
rect 2544 16528 2608 16592
rect 2480 16512 2672 16528
rect 2544 16448 2608 16512
rect 2480 16432 2672 16448
rect 2544 16368 2608 16432
rect 2480 16351 2672 16368
rect 2544 16287 2608 16351
rect 2480 16270 2672 16287
rect 2544 16206 2608 16270
rect 2480 16189 2672 16206
rect 2544 16125 2608 16189
rect 2480 16108 2672 16125
rect 2544 16044 2608 16108
rect 2480 16027 2672 16044
rect 2544 15963 2608 16027
rect 2480 15946 2672 15963
rect 2544 15882 2608 15946
rect 2480 15865 2672 15882
rect 2544 15801 2608 15865
rect 2480 15784 2672 15801
rect 2544 15720 2608 15784
rect 2480 15703 2672 15720
rect 2544 15639 2608 15703
rect 2480 15622 2672 15639
rect 2544 15558 2608 15622
rect 2480 15541 2672 15558
rect 2544 15477 2608 15541
rect 2480 15460 2672 15477
rect 2544 15396 2608 15460
rect 2480 15379 2672 15396
rect 2544 15315 2608 15379
rect 2480 15298 2672 15315
rect 2544 15234 2608 15298
rect 2480 15217 2672 15234
rect 2544 15153 2608 15217
rect 2480 15136 2672 15153
rect 2544 15072 2608 15136
rect 2480 15055 2672 15072
rect 2544 14991 2608 15055
rect 2480 14974 2672 14991
rect 2544 14910 2608 14974
rect 2480 14893 2672 14910
rect 2544 14829 2608 14893
rect 2480 14812 2672 14829
rect 2544 14748 2608 14812
rect 2480 14731 2672 14748
rect 2544 14667 2608 14731
rect 2480 14650 2672 14667
rect 2544 14586 2608 14650
rect 2480 14569 2672 14586
rect 2544 14505 2608 14569
rect 2480 14488 2672 14505
rect 2544 14424 2608 14488
rect 2480 14407 2672 14424
rect 2544 14343 2608 14407
rect 2480 14326 2672 14343
rect 2544 14262 2608 14326
rect 2480 14245 2672 14262
rect 2544 14181 2608 14245
rect 2480 14164 2672 14181
rect 2544 14100 2608 14164
rect 2480 14083 2672 14100
rect 2544 14019 2608 14083
rect 2480 14002 2672 14019
rect 2544 13938 2608 14002
rect 2480 13921 2672 13938
rect 2544 13857 2608 13921
rect 2480 13840 2672 13857
rect 2544 13776 2608 13840
rect 2480 13759 2672 13776
rect 2544 13695 2608 13759
rect 2480 13678 2672 13695
rect 2544 13614 2608 13678
rect 2480 13607 2672 13614
rect 2980 23686 3164 26492
rect 2980 23630 2985 23686
rect 3041 23630 3103 23686
rect 3159 23630 3164 23686
rect 2980 23606 3164 23630
rect 2980 23550 2985 23606
rect 3041 23550 3103 23606
rect 3159 23550 3164 23606
rect 2980 23526 3164 23550
rect 2980 23470 2985 23526
rect 3041 23470 3103 23526
rect 3159 23470 3164 23526
rect 2980 23446 3164 23470
rect 2980 23390 2985 23446
rect 3041 23390 3103 23446
rect 3159 23390 3164 23446
rect 2980 23366 3164 23390
rect 2980 23310 2985 23366
rect 3041 23310 3103 23366
rect 3159 23310 3164 23366
rect 2980 23286 3164 23310
rect 2980 23230 2985 23286
rect 3041 23230 3103 23286
rect 3159 23230 3164 23286
rect 2980 23206 3164 23230
rect 2980 23150 2985 23206
rect 3041 23150 3103 23206
rect 3159 23150 3164 23206
rect 2980 23126 3164 23150
rect 2980 23070 2985 23126
rect 3041 23070 3103 23126
rect 3159 23070 3164 23126
rect 2980 23046 3164 23070
rect 2980 22990 2985 23046
rect 3041 22990 3103 23046
rect 3159 22990 3164 23046
rect 2980 22966 3164 22990
rect 2980 22910 2985 22966
rect 3041 22910 3103 22966
rect 3159 22910 3164 22966
rect 2980 22886 3164 22910
rect 2980 22830 2985 22886
rect 3041 22830 3103 22886
rect 3159 22830 3164 22886
rect 2980 22806 3164 22830
rect 2980 22750 2985 22806
rect 3041 22750 3103 22806
rect 3159 22750 3164 22806
rect 2980 22726 3164 22750
rect 2980 22670 2985 22726
rect 3041 22670 3103 22726
rect 3159 22670 3164 22726
rect 2980 22646 3164 22670
rect 2980 22590 2985 22646
rect 3041 22590 3103 22646
rect 3159 22590 3164 22646
rect 2980 22566 3164 22590
rect 2980 22510 2985 22566
rect 3041 22510 3103 22566
rect 3159 22510 3164 22566
rect 2980 22486 3164 22510
rect 2980 22430 2985 22486
rect 3041 22430 3103 22486
rect 3159 22430 3164 22486
rect 2980 22406 3164 22430
rect 2980 22350 2985 22406
rect 3041 22350 3103 22406
rect 3159 22350 3164 22406
rect 2980 22326 3164 22350
rect 2980 22270 2985 22326
rect 3041 22270 3103 22326
rect 3159 22270 3164 22326
rect 2980 22245 3164 22270
rect 2980 22189 2985 22245
rect 3041 22189 3103 22245
rect 3159 22189 3164 22245
rect 2980 22164 3164 22189
rect 2980 22108 2985 22164
rect 3041 22108 3103 22164
rect 3159 22108 3164 22164
rect 2980 22083 3164 22108
rect 2980 22027 2985 22083
rect 3041 22027 3103 22083
rect 3159 22027 3164 22083
rect 2980 22002 3164 22027
rect 2980 21946 2985 22002
rect 3041 21946 3103 22002
rect 3159 21946 3164 22002
rect 2980 21921 3164 21946
rect 2980 21865 2985 21921
rect 3041 21865 3103 21921
rect 3159 21865 3164 21921
rect 2980 21840 3164 21865
rect 2980 21784 2985 21840
rect 3041 21784 3103 21840
rect 3159 21784 3164 21840
rect 2980 21759 3164 21784
rect 2980 21703 2985 21759
rect 3041 21703 3103 21759
rect 3159 21703 3164 21759
rect 2980 21678 3164 21703
rect 2980 21622 2985 21678
rect 3041 21622 3103 21678
rect 3159 21622 3164 21678
rect 2980 21597 3164 21622
rect 2980 21541 2985 21597
rect 3041 21541 3103 21597
rect 3159 21541 3164 21597
rect 2980 21516 3164 21541
rect 2980 21460 2985 21516
rect 3041 21460 3103 21516
rect 3159 21460 3164 21516
rect 2980 21435 3164 21460
rect 2980 21379 2985 21435
rect 3041 21379 3103 21435
rect 3159 21379 3164 21435
rect 2980 21354 3164 21379
rect 2980 21298 2985 21354
rect 3041 21298 3103 21354
rect 3159 21298 3164 21354
rect 2980 21273 3164 21298
rect 2980 21217 2985 21273
rect 3041 21217 3103 21273
rect 3159 21217 3164 21273
rect 2980 21192 3164 21217
rect 2980 21136 2985 21192
rect 3041 21136 3103 21192
rect 3159 21136 3164 21192
rect 2980 19673 3164 21136
rect 3044 19609 3100 19673
rect 2980 19581 3164 19609
rect 3044 19517 3100 19581
rect 2980 19489 3164 19517
rect 3044 19425 3100 19489
rect 2980 19397 3164 19425
rect 3044 19333 3100 19397
rect 2980 19305 3164 19333
rect 3044 19241 3100 19305
rect 2980 19212 3164 19241
rect 3044 19148 3100 19212
tri 2974 13058 2980 13064 se
rect 2980 13058 3164 19148
rect 3472 26492 3570 27206
rect 3870 27161 4062 29420
rect 4366 32018 4558 34764
rect 5358 39592 5550 39600
rect 5422 39528 5486 39592
rect 5358 39512 5550 39528
rect 5422 39448 5486 39512
rect 5358 39432 5550 39448
rect 5422 39368 5486 39432
rect 5358 39352 5550 39368
rect 5422 39288 5486 39352
rect 5358 39272 5550 39288
rect 5422 39208 5486 39272
rect 5358 39192 5550 39208
rect 5422 39128 5486 39192
rect 5358 39112 5550 39128
rect 5422 39048 5486 39112
rect 5358 39032 5550 39048
rect 5422 38968 5486 39032
rect 5358 38952 5550 38968
rect 5422 38888 5486 38952
rect 5358 38872 5550 38888
rect 5422 38808 5486 38872
rect 5358 38792 5550 38808
rect 5422 38728 5486 38792
rect 5358 38712 5550 38728
rect 5422 38648 5486 38712
rect 5358 38632 5550 38648
rect 5422 38568 5486 38632
rect 5358 38552 5550 38568
rect 5422 38488 5486 38552
rect 5358 38472 5550 38488
rect 5422 38408 5486 38472
rect 5358 38392 5550 38408
rect 5422 38328 5486 38392
rect 5358 38311 5550 38328
rect 5422 38247 5486 38311
rect 5358 38230 5550 38247
rect 5422 38166 5486 38230
rect 5358 38149 5550 38166
rect 5422 38085 5486 38149
rect 5358 38068 5550 38085
rect 5422 38004 5486 38068
rect 5358 37987 5550 38004
rect 5422 37923 5486 37987
rect 5358 37906 5550 37923
rect 5422 37842 5486 37906
rect 5358 37825 5550 37842
rect 5422 37761 5486 37825
rect 5358 37744 5550 37761
rect 5422 37680 5486 37744
rect 5358 37663 5550 37680
rect 5422 37599 5486 37663
rect 5358 37582 5550 37599
rect 5422 37518 5486 37582
rect 5358 37501 5550 37518
rect 5422 37437 5486 37501
rect 5358 37420 5550 37437
rect 5422 37356 5486 37420
rect 5358 37339 5550 37356
rect 5422 37275 5486 37339
rect 5358 37258 5550 37275
rect 5422 37194 5486 37258
rect 5358 37177 5550 37194
rect 5422 37113 5486 37177
rect 5358 37096 5550 37113
rect 5422 37032 5486 37096
rect 5358 37015 5550 37032
rect 5422 36951 5486 37015
rect 5358 36934 5550 36951
rect 5422 36870 5486 36934
rect 5358 36853 5550 36870
rect 5422 36789 5486 36853
rect 5358 36772 5550 36789
rect 5422 36708 5486 36772
rect 5358 36691 5550 36708
rect 5422 36627 5486 36691
rect 5358 36610 5550 36627
rect 5422 36546 5486 36610
rect 5358 36529 5550 36546
rect 5422 36465 5486 36529
rect 5358 36448 5550 36465
rect 5422 36384 5486 36448
rect 5358 36367 5550 36384
rect 5422 36303 5486 36367
rect 5358 36286 5550 36303
rect 5422 36222 5486 36286
rect 5358 36205 5550 36222
rect 5422 36141 5486 36205
rect 5358 36124 5550 36141
rect 5422 36060 5486 36124
rect 5358 36043 5550 36060
rect 5422 35979 5486 36043
rect 5358 35962 5550 35979
rect 5422 35898 5486 35962
rect 5358 35881 5550 35898
rect 5422 35817 5486 35881
rect 5358 35800 5550 35817
rect 5422 35736 5486 35800
rect 5358 35719 5550 35736
rect 5422 35655 5486 35719
rect 5358 35638 5550 35655
rect 5422 35574 5486 35638
rect 5358 35557 5550 35574
rect 5422 35493 5486 35557
rect 5358 35476 5550 35493
rect 5422 35412 5486 35476
rect 5358 35395 5550 35412
rect 5422 35331 5486 35395
rect 5358 35314 5550 35331
rect 5422 35250 5486 35314
rect 5358 35233 5550 35250
rect 5422 35169 5486 35233
rect 5358 35152 5550 35169
rect 5422 35088 5486 35152
rect 5358 35071 5550 35088
rect 5422 35007 5486 35071
rect 5358 34990 5550 35007
rect 5422 34926 5486 34990
rect 5358 34909 5550 34926
rect 5422 34845 5486 34909
rect 5358 34828 5550 34845
rect 5422 34764 5486 34828
rect 4366 31962 4371 32018
rect 4427 31962 4497 32018
rect 4553 31962 4558 32018
rect 4366 31936 4558 31962
rect 4366 31880 4371 31936
rect 4427 31880 4497 31936
rect 4553 31880 4558 31936
rect 4366 31854 4558 31880
rect 4366 31798 4371 31854
rect 4427 31798 4497 31854
rect 4553 31798 4558 31854
rect 4366 31772 4558 31798
rect 4366 31716 4371 31772
rect 4427 31716 4497 31772
rect 4553 31716 4558 31772
rect 4366 31690 4558 31716
rect 4366 31634 4371 31690
rect 4427 31634 4497 31690
rect 4553 31634 4558 31690
rect 4366 31608 4558 31634
rect 4366 31552 4371 31608
rect 4427 31552 4497 31608
rect 4553 31552 4558 31608
rect 4366 31526 4558 31552
rect 4366 31470 4371 31526
rect 4427 31470 4497 31526
rect 4553 31470 4558 31526
rect 4366 31444 4558 31470
rect 4366 31388 4371 31444
rect 4427 31388 4497 31444
rect 4553 31388 4558 31444
rect 4366 31362 4558 31388
rect 4366 31306 4371 31362
rect 4427 31306 4497 31362
rect 4553 31306 4558 31362
rect 4366 31280 4558 31306
rect 4366 31224 4371 31280
rect 4427 31224 4497 31280
rect 4553 31224 4558 31280
rect 4366 31198 4558 31224
rect 4366 31142 4371 31198
rect 4427 31142 4497 31198
rect 4553 31142 4558 31198
rect 4366 31116 4558 31142
rect 4366 31060 4371 31116
rect 4427 31060 4497 31116
rect 4553 31060 4558 31116
rect 4366 31034 4558 31060
rect 4366 30978 4371 31034
rect 4427 30978 4497 31034
rect 4553 30978 4558 31034
rect 4366 30952 4558 30978
rect 4366 30896 4371 30952
rect 4427 30896 4497 30952
rect 4553 30896 4558 30952
rect 4366 30870 4558 30896
rect 4366 30814 4371 30870
rect 4427 30814 4497 30870
rect 4553 30814 4558 30870
rect 4366 30788 4558 30814
rect 4366 30732 4371 30788
rect 4427 30732 4497 30788
rect 4553 30732 4558 30788
rect 4366 30706 4558 30732
rect 4366 30650 4371 30706
rect 4427 30650 4497 30706
rect 4553 30650 4558 30706
rect 4366 30624 4558 30650
rect 4366 30568 4371 30624
rect 4427 30568 4497 30624
rect 4553 30568 4558 30624
rect 4366 30542 4558 30568
rect 4366 30486 4371 30542
rect 4427 30486 4497 30542
rect 4553 30486 4558 30542
rect 4366 30460 4558 30486
rect 4366 30404 4371 30460
rect 4427 30404 4497 30460
rect 4553 30404 4558 30460
rect 4366 30378 4558 30404
rect 4366 30322 4371 30378
rect 4427 30322 4497 30378
rect 4553 30322 4558 30378
rect 4366 30296 4558 30322
rect 4366 30240 4371 30296
rect 4427 30240 4497 30296
rect 4553 30240 4558 30296
rect 4366 30214 4558 30240
rect 4366 30158 4371 30214
rect 4427 30158 4497 30214
rect 4553 30158 4558 30214
rect 4366 30132 4558 30158
rect 4366 30076 4371 30132
rect 4427 30076 4497 30132
rect 4553 30076 4558 30132
rect 4366 30050 4558 30076
rect 4366 29994 4371 30050
rect 4427 29994 4497 30050
rect 4553 29994 4558 30050
rect 4366 29968 4558 29994
rect 4366 29912 4371 29968
rect 4427 29912 4497 29968
rect 4553 29912 4558 29968
rect 4366 29886 4558 29912
rect 4366 29830 4371 29886
rect 4427 29830 4497 29886
rect 4553 29830 4558 29886
rect 4366 29804 4558 29830
rect 4366 29748 4371 29804
rect 4427 29748 4497 29804
rect 4553 29748 4558 29804
rect 4366 29722 4558 29748
rect 4366 29666 4371 29722
rect 4427 29666 4497 29722
rect 4553 29666 4558 29722
rect 4366 29640 4558 29666
rect 4366 29584 4371 29640
rect 4427 29584 4497 29640
rect 4553 29584 4558 29640
rect 4366 29558 4558 29584
rect 4366 29502 4371 29558
rect 4427 29502 4497 29558
rect 4553 29502 4558 29558
rect 4366 29476 4558 29502
rect 4366 29420 4371 29476
rect 4427 29420 4497 29476
rect 4553 29420 4558 29476
rect 4366 29415 4558 29420
rect 4862 34219 5054 34225
rect 4926 34155 4990 34219
rect 4862 34125 5054 34155
rect 4926 34061 4990 34125
rect 4862 34030 5054 34061
rect 4926 33966 4990 34030
rect 4862 33935 5054 33966
rect 4926 33871 4990 33935
rect 4862 33840 5054 33871
rect 4926 33776 4990 33840
rect 4862 33745 5054 33776
rect 4926 33681 4990 33745
rect 4862 32018 5054 33681
rect 4862 31962 4867 32018
rect 4923 31962 4993 32018
rect 5049 31962 5054 32018
rect 4862 31936 5054 31962
rect 4862 31880 4867 31936
rect 4923 31880 4993 31936
rect 5049 31880 5054 31936
rect 4862 31854 5054 31880
rect 4862 31798 4867 31854
rect 4923 31798 4993 31854
rect 5049 31798 5054 31854
rect 4862 31772 5054 31798
rect 4862 31716 4867 31772
rect 4923 31716 4993 31772
rect 5049 31716 5054 31772
rect 4862 31690 5054 31716
rect 4862 31634 4867 31690
rect 4923 31634 4993 31690
rect 5049 31634 5054 31690
rect 4862 31608 5054 31634
rect 4862 31552 4867 31608
rect 4923 31552 4993 31608
rect 5049 31552 5054 31608
rect 4862 31526 5054 31552
rect 4862 31470 4867 31526
rect 4923 31470 4993 31526
rect 5049 31470 5054 31526
rect 4862 31444 5054 31470
rect 4862 31388 4867 31444
rect 4923 31388 4993 31444
rect 5049 31388 5054 31444
rect 4862 31362 5054 31388
rect 4862 31306 4867 31362
rect 4923 31306 4993 31362
rect 5049 31306 5054 31362
rect 4862 31280 5054 31306
rect 4862 31224 4867 31280
rect 4923 31224 4993 31280
rect 5049 31224 5054 31280
rect 4862 31198 5054 31224
rect 4862 31142 4867 31198
rect 4923 31142 4993 31198
rect 5049 31142 5054 31198
rect 4862 31116 5054 31142
rect 4862 31060 4867 31116
rect 4923 31060 4993 31116
rect 5049 31060 5054 31116
rect 4862 31034 5054 31060
rect 4862 30978 4867 31034
rect 4923 30978 4993 31034
rect 5049 30978 5054 31034
rect 4862 30952 5054 30978
rect 4862 30896 4867 30952
rect 4923 30896 4993 30952
rect 5049 30896 5054 30952
rect 4862 30870 5054 30896
rect 4862 30814 4867 30870
rect 4923 30814 4993 30870
rect 5049 30814 5054 30870
rect 4862 30788 5054 30814
rect 4862 30732 4867 30788
rect 4923 30732 4993 30788
rect 5049 30732 5054 30788
rect 4862 30706 5054 30732
rect 4862 30650 4867 30706
rect 4923 30650 4993 30706
rect 5049 30650 5054 30706
rect 4862 30624 5054 30650
rect 4862 30568 4867 30624
rect 4923 30568 4993 30624
rect 5049 30568 5054 30624
rect 4862 30542 5054 30568
rect 4862 30486 4867 30542
rect 4923 30486 4993 30542
rect 5049 30486 5054 30542
rect 4862 30460 5054 30486
rect 4862 30404 4867 30460
rect 4923 30404 4993 30460
rect 5049 30404 5054 30460
rect 4862 30378 5054 30404
rect 4862 30322 4867 30378
rect 4923 30322 4993 30378
rect 5049 30322 5054 30378
rect 4862 30296 5054 30322
rect 4862 30240 4867 30296
rect 4923 30240 4993 30296
rect 5049 30240 5054 30296
rect 4862 30214 5054 30240
rect 4862 30158 4867 30214
rect 4923 30158 4993 30214
rect 5049 30158 5054 30214
rect 4862 30132 5054 30158
rect 4862 30076 4867 30132
rect 4923 30076 4993 30132
rect 5049 30076 5054 30132
rect 4862 30050 5054 30076
rect 4862 29994 4867 30050
rect 4923 29994 4993 30050
rect 5049 29994 5054 30050
rect 4862 29968 5054 29994
rect 4862 29912 4867 29968
rect 4923 29912 4993 29968
rect 5049 29912 5054 29968
rect 4862 29886 5054 29912
rect 4862 29830 4867 29886
rect 4923 29830 4993 29886
rect 5049 29830 5054 29886
rect 4862 29804 5054 29830
rect 4862 29748 4867 29804
rect 4923 29748 4993 29804
rect 5049 29748 5054 29804
rect 4862 29722 5054 29748
rect 4862 29666 4867 29722
rect 4923 29666 4993 29722
rect 5049 29666 5054 29722
rect 4862 29640 5054 29666
rect 4862 29584 4867 29640
rect 4923 29584 4993 29640
rect 5049 29584 5054 29640
rect 4862 29558 5054 29584
rect 4862 29502 4867 29558
rect 4923 29502 4993 29558
rect 5049 29502 5054 29558
rect 4862 29476 5054 29502
rect 4862 29420 4867 29476
rect 4923 29420 4993 29476
rect 5049 29420 5054 29476
rect 4464 28620 4562 28633
rect 4464 28564 4485 28620
rect 4541 28564 4562 28620
rect 4464 28451 4562 28564
rect 4464 28395 4485 28451
rect 4541 28395 4562 28451
rect 4464 28282 4562 28395
rect 4464 28226 4485 28282
rect 4541 28226 4562 28282
rect 4464 28113 4562 28226
rect 4464 28057 4485 28113
rect 4541 28057 4562 28113
rect 4464 27944 4562 28057
rect 4464 27888 4485 27944
rect 4541 27888 4562 27944
rect 4464 27774 4562 27888
rect 4464 27718 4485 27774
rect 4541 27718 4562 27774
rect 4464 27604 4562 27718
rect 4464 27548 4485 27604
rect 4541 27548 4562 27604
rect 4464 27434 4562 27548
rect 4464 27378 4485 27434
rect 4541 27378 4562 27434
rect 4464 27264 4562 27378
rect 4464 27208 4485 27264
rect 4541 27208 4562 27264
tri 4062 27161 4096 27195 sw
rect 3870 27137 4096 27161
tri 4096 27137 4120 27161 sw
rect 3870 27101 4120 27137
tri 4120 27101 4156 27137 sw
rect 3870 26726 4156 27101
tri 3870 26716 3880 26726 ne
rect 3880 26716 4156 26726
tri 3880 26660 3936 26716 ne
rect 3936 26660 4156 26716
tri 3936 26657 3939 26660 ne
rect 3939 26657 4156 26660
tri 3939 26632 3964 26657 ne
rect 3964 26632 4156 26657
tri 3964 26624 3972 26632 ne
tri 3570 26492 3626 26548 sw
rect 3472 26454 3626 26492
tri 3626 26454 3664 26492 sw
rect 3472 26176 3664 26454
rect 3472 26120 3477 26176
rect 3533 26120 3603 26176
rect 3659 26120 3664 26176
rect 3472 26081 3664 26120
rect 3472 26025 3477 26081
rect 3533 26025 3603 26081
rect 3659 26025 3664 26081
rect 3472 25986 3664 26025
rect 3472 25930 3477 25986
rect 3533 25930 3603 25986
rect 3659 25930 3664 25986
rect 3472 25891 3664 25930
rect 3472 25835 3477 25891
rect 3533 25835 3603 25891
rect 3659 25835 3664 25891
rect 3472 25795 3664 25835
rect 3472 25739 3477 25795
rect 3533 25739 3603 25795
rect 3659 25739 3664 25795
rect 3472 25699 3664 25739
rect 3472 25643 3477 25699
rect 3533 25643 3603 25699
rect 3659 25643 3664 25699
rect 3472 23686 3664 25643
rect 3472 23630 3481 23686
rect 3537 23630 3599 23686
rect 3655 23630 3664 23686
rect 3472 23606 3664 23630
rect 3472 23550 3481 23606
rect 3537 23550 3599 23606
rect 3655 23550 3664 23606
rect 3472 23526 3664 23550
rect 3472 23470 3481 23526
rect 3537 23470 3599 23526
rect 3655 23470 3664 23526
rect 3472 23446 3664 23470
rect 3472 23390 3481 23446
rect 3537 23390 3599 23446
rect 3655 23390 3664 23446
rect 3472 23366 3664 23390
rect 3472 23310 3481 23366
rect 3537 23310 3599 23366
rect 3655 23310 3664 23366
rect 3472 23286 3664 23310
rect 3472 23230 3481 23286
rect 3537 23230 3599 23286
rect 3655 23230 3664 23286
rect 3472 23206 3664 23230
rect 3472 23150 3481 23206
rect 3537 23150 3599 23206
rect 3655 23150 3664 23206
rect 3472 23126 3664 23150
rect 3472 23070 3481 23126
rect 3537 23070 3599 23126
rect 3655 23070 3664 23126
rect 3472 23046 3664 23070
rect 3472 22990 3481 23046
rect 3537 22990 3599 23046
rect 3655 22990 3664 23046
rect 3472 22966 3664 22990
rect 3472 22910 3481 22966
rect 3537 22910 3599 22966
rect 3655 22910 3664 22966
rect 3472 22886 3664 22910
rect 3472 22830 3481 22886
rect 3537 22830 3599 22886
rect 3655 22830 3664 22886
rect 3472 22806 3664 22830
rect 3472 22750 3481 22806
rect 3537 22750 3599 22806
rect 3655 22750 3664 22806
rect 3472 22726 3664 22750
rect 3472 22670 3481 22726
rect 3537 22670 3599 22726
rect 3655 22670 3664 22726
rect 3472 22646 3664 22670
rect 3472 22590 3481 22646
rect 3537 22590 3599 22646
rect 3655 22590 3664 22646
rect 3472 22566 3664 22590
rect 3472 22510 3481 22566
rect 3537 22510 3599 22566
rect 3655 22510 3664 22566
rect 3472 22486 3664 22510
rect 3472 22430 3481 22486
rect 3537 22430 3599 22486
rect 3655 22430 3664 22486
rect 3472 22406 3664 22430
rect 3472 22350 3481 22406
rect 3537 22350 3599 22406
rect 3655 22350 3664 22406
rect 3472 22326 3664 22350
rect 3472 22270 3481 22326
rect 3537 22270 3599 22326
rect 3655 22270 3664 22326
rect 3472 22245 3664 22270
rect 3472 22189 3481 22245
rect 3537 22189 3599 22245
rect 3655 22189 3664 22245
rect 3472 22164 3664 22189
rect 3472 22108 3481 22164
rect 3537 22108 3599 22164
rect 3655 22108 3664 22164
rect 3472 22083 3664 22108
rect 3472 22027 3481 22083
rect 3537 22027 3599 22083
rect 3655 22027 3664 22083
rect 3472 22002 3664 22027
rect 3472 21946 3481 22002
rect 3537 21946 3599 22002
rect 3655 21946 3664 22002
rect 3472 21921 3664 21946
rect 3472 21865 3481 21921
rect 3537 21865 3599 21921
rect 3655 21865 3664 21921
rect 3472 21840 3664 21865
rect 3472 21784 3481 21840
rect 3537 21784 3599 21840
rect 3655 21784 3664 21840
rect 3472 21759 3664 21784
rect 3472 21703 3481 21759
rect 3537 21703 3599 21759
rect 3655 21703 3664 21759
rect 3472 21678 3664 21703
rect 3472 21622 3481 21678
rect 3537 21622 3599 21678
rect 3655 21622 3664 21678
rect 3472 21597 3664 21622
rect 3472 21541 3481 21597
rect 3537 21541 3599 21597
rect 3655 21541 3664 21597
rect 3472 21516 3664 21541
rect 3472 21460 3481 21516
rect 3537 21460 3599 21516
rect 3655 21460 3664 21516
rect 3472 21435 3664 21460
rect 3472 21379 3481 21435
rect 3537 21379 3599 21435
rect 3655 21379 3664 21435
rect 3472 21354 3664 21379
rect 3472 21298 3481 21354
rect 3537 21298 3599 21354
rect 3655 21298 3664 21354
rect 3472 21273 3664 21298
rect 3472 21217 3481 21273
rect 3537 21217 3599 21273
rect 3655 21217 3664 21273
rect 3472 21192 3664 21217
rect 3472 21136 3481 21192
rect 3537 21136 3599 21192
rect 3655 21136 3664 21192
rect 3472 18592 3664 21136
rect 3536 18528 3600 18592
rect 3472 18512 3664 18528
rect 3536 18448 3600 18512
rect 3472 18432 3664 18448
rect 3536 18368 3600 18432
rect 3472 18352 3664 18368
rect 3536 18288 3600 18352
rect 3472 18272 3664 18288
rect 3536 18208 3600 18272
rect 3472 18192 3664 18208
rect 3536 18128 3600 18192
rect 3472 18112 3664 18128
rect 3536 18048 3600 18112
rect 3472 18032 3664 18048
rect 3536 17968 3600 18032
rect 3472 17952 3664 17968
rect 3536 17888 3600 17952
rect 3472 17872 3664 17888
rect 3536 17808 3600 17872
rect 3472 17792 3664 17808
rect 3536 17728 3600 17792
rect 3472 17712 3664 17728
rect 3536 17648 3600 17712
rect 3472 17632 3664 17648
rect 3536 17568 3600 17632
rect 3472 17552 3664 17568
rect 3536 17488 3600 17552
rect 3472 17472 3664 17488
rect 3536 17408 3600 17472
rect 3472 17392 3664 17408
rect 3536 17328 3600 17392
rect 3472 17312 3664 17328
rect 3536 17248 3600 17312
rect 3472 17232 3664 17248
rect 3536 17168 3600 17232
rect 3472 17152 3664 17168
rect 3536 17088 3600 17152
rect 3472 17072 3664 17088
rect 3536 17008 3600 17072
rect 3472 16992 3664 17008
rect 3536 16928 3600 16992
rect 3472 16912 3664 16928
rect 3536 16848 3600 16912
rect 3472 16832 3664 16848
rect 3536 16768 3600 16832
rect 3472 16752 3664 16768
rect 3536 16688 3600 16752
rect 3472 16672 3664 16688
rect 3536 16608 3600 16672
rect 3472 16592 3664 16608
rect 3536 16528 3600 16592
rect 3472 16512 3664 16528
rect 3536 16448 3600 16512
rect 3472 16432 3664 16448
rect 3536 16368 3600 16432
rect 3472 16351 3664 16368
rect 3536 16287 3600 16351
rect 3472 16270 3664 16287
rect 3536 16206 3600 16270
rect 3472 16189 3664 16206
rect 3536 16125 3600 16189
rect 3472 16108 3664 16125
rect 3536 16044 3600 16108
rect 3472 16027 3664 16044
rect 3536 15963 3600 16027
rect 3472 15946 3664 15963
rect 3536 15882 3600 15946
rect 3472 15865 3664 15882
rect 3536 15801 3600 15865
rect 3472 15784 3664 15801
rect 3536 15720 3600 15784
rect 3472 15703 3664 15720
rect 3536 15639 3600 15703
rect 3472 15622 3664 15639
rect 3536 15558 3600 15622
rect 3472 15541 3664 15558
rect 3536 15477 3600 15541
rect 3472 15460 3664 15477
rect 3536 15396 3600 15460
rect 3472 15379 3664 15396
rect 3536 15315 3600 15379
rect 3472 15298 3664 15315
rect 3536 15234 3600 15298
rect 3472 15217 3664 15234
rect 3536 15153 3600 15217
rect 3472 15136 3664 15153
rect 3536 15072 3600 15136
rect 3472 15055 3664 15072
rect 3536 14991 3600 15055
rect 3472 14974 3664 14991
rect 3536 14910 3600 14974
rect 3472 14893 3664 14910
rect 3536 14829 3600 14893
rect 3472 14812 3664 14829
rect 3536 14748 3600 14812
rect 3472 14731 3664 14748
rect 3536 14667 3600 14731
rect 3472 14650 3664 14667
rect 3536 14586 3600 14650
rect 3472 14569 3664 14586
rect 3536 14505 3600 14569
rect 3472 14488 3664 14505
rect 3536 14424 3600 14488
rect 3472 14407 3664 14424
rect 3536 14343 3600 14407
rect 3472 14326 3664 14343
rect 3536 14262 3600 14326
rect 3472 14245 3664 14262
rect 3536 14181 3600 14245
rect 3472 14164 3664 14181
rect 3536 14100 3600 14164
rect 3472 14083 3664 14100
rect 3536 14019 3600 14083
rect 3472 14002 3664 14019
rect 3536 13938 3600 14002
rect 3472 13921 3664 13938
rect 3536 13857 3600 13921
rect 3472 13840 3664 13857
rect 3536 13776 3600 13840
rect 3472 13759 3664 13776
rect 3536 13695 3600 13759
rect 3472 13678 3664 13695
rect 3536 13614 3600 13678
rect 3472 13607 3664 13614
rect 3972 23686 4156 26632
rect 3972 23630 3977 23686
rect 4033 23630 4095 23686
rect 4151 23630 4156 23686
rect 3972 23606 4156 23630
rect 3972 23550 3977 23606
rect 4033 23550 4095 23606
rect 4151 23550 4156 23606
rect 3972 23526 4156 23550
rect 3972 23470 3977 23526
rect 4033 23470 4095 23526
rect 4151 23470 4156 23526
rect 3972 23446 4156 23470
rect 3972 23390 3977 23446
rect 4033 23390 4095 23446
rect 4151 23390 4156 23446
rect 3972 23366 4156 23390
rect 3972 23310 3977 23366
rect 4033 23310 4095 23366
rect 4151 23310 4156 23366
rect 3972 23286 4156 23310
rect 3972 23230 3977 23286
rect 4033 23230 4095 23286
rect 4151 23230 4156 23286
rect 3972 23206 4156 23230
rect 3972 23150 3977 23206
rect 4033 23150 4095 23206
rect 4151 23150 4156 23206
rect 3972 23126 4156 23150
rect 3972 23070 3977 23126
rect 4033 23070 4095 23126
rect 4151 23070 4156 23126
rect 3972 23046 4156 23070
rect 3972 22990 3977 23046
rect 4033 22990 4095 23046
rect 4151 22990 4156 23046
rect 3972 22966 4156 22990
rect 3972 22910 3977 22966
rect 4033 22910 4095 22966
rect 4151 22910 4156 22966
rect 3972 22886 4156 22910
rect 3972 22830 3977 22886
rect 4033 22830 4095 22886
rect 4151 22830 4156 22886
rect 3972 22806 4156 22830
rect 3972 22750 3977 22806
rect 4033 22750 4095 22806
rect 4151 22750 4156 22806
rect 3972 22726 4156 22750
rect 3972 22670 3977 22726
rect 4033 22670 4095 22726
rect 4151 22670 4156 22726
rect 3972 22646 4156 22670
rect 3972 22590 3977 22646
rect 4033 22590 4095 22646
rect 4151 22590 4156 22646
rect 3972 22566 4156 22590
rect 3972 22510 3977 22566
rect 4033 22510 4095 22566
rect 4151 22510 4156 22566
rect 3972 22486 4156 22510
rect 3972 22430 3977 22486
rect 4033 22430 4095 22486
rect 4151 22430 4156 22486
rect 3972 22406 4156 22430
rect 3972 22350 3977 22406
rect 4033 22350 4095 22406
rect 4151 22350 4156 22406
rect 3972 22326 4156 22350
rect 3972 22270 3977 22326
rect 4033 22270 4095 22326
rect 4151 22270 4156 22326
rect 3972 22245 4156 22270
rect 3972 22189 3977 22245
rect 4033 22189 4095 22245
rect 4151 22189 4156 22245
rect 3972 22164 4156 22189
rect 3972 22108 3977 22164
rect 4033 22108 4095 22164
rect 4151 22108 4156 22164
rect 3972 22083 4156 22108
rect 3972 22027 3977 22083
rect 4033 22027 4095 22083
rect 4151 22027 4156 22083
rect 3972 22002 4156 22027
rect 3972 21946 3977 22002
rect 4033 21946 4095 22002
rect 4151 21946 4156 22002
rect 3972 21921 4156 21946
rect 3972 21865 3977 21921
rect 4033 21865 4095 21921
rect 4151 21865 4156 21921
rect 3972 21840 4156 21865
rect 3972 21784 3977 21840
rect 4033 21784 4095 21840
rect 4151 21784 4156 21840
rect 3972 21759 4156 21784
rect 3972 21703 3977 21759
rect 4033 21703 4095 21759
rect 4151 21703 4156 21759
rect 3972 21678 4156 21703
rect 3972 21622 3977 21678
rect 4033 21622 4095 21678
rect 4151 21622 4156 21678
rect 3972 21597 4156 21622
rect 3972 21541 3977 21597
rect 4033 21541 4095 21597
rect 4151 21541 4156 21597
rect 3972 21516 4156 21541
rect 3972 21460 3977 21516
rect 4033 21460 4095 21516
rect 4151 21460 4156 21516
rect 3972 21435 4156 21460
rect 3972 21379 3977 21435
rect 4033 21379 4095 21435
rect 4151 21379 4156 21435
rect 3972 21354 4156 21379
rect 3972 21298 3977 21354
rect 4033 21298 4095 21354
rect 4151 21298 4156 21354
rect 3972 21273 4156 21298
rect 3972 21217 3977 21273
rect 4033 21217 4095 21273
rect 4151 21217 4156 21273
rect 3972 21192 4156 21217
rect 3972 21136 3977 21192
rect 4033 21136 4095 21192
rect 4151 21136 4156 21192
rect 3972 19673 4156 21136
rect 4036 19609 4092 19673
rect 3972 19581 4156 19609
rect 4036 19517 4092 19581
rect 3972 19488 4156 19517
rect 4036 19424 4092 19488
rect 3972 19395 4156 19424
rect 4036 19331 4092 19395
rect 3972 19302 4156 19331
rect 4036 19238 4092 19302
rect 3972 19209 4156 19238
rect 4036 19145 4092 19209
tri 3966 13058 3972 13064 se
rect 3972 13060 4156 19145
rect 4464 26548 4562 27208
rect 4862 27161 5054 29420
rect 5358 32018 5550 34764
rect 6350 39592 6542 39600
rect 6414 39528 6478 39592
rect 6350 39512 6542 39528
rect 6414 39448 6478 39512
rect 6350 39432 6542 39448
rect 6414 39368 6478 39432
rect 6350 39352 6542 39368
rect 6414 39288 6478 39352
rect 6350 39272 6542 39288
rect 6414 39208 6478 39272
rect 6350 39192 6542 39208
rect 6414 39128 6478 39192
rect 6350 39112 6542 39128
rect 6414 39048 6478 39112
rect 6350 39032 6542 39048
rect 6414 38968 6478 39032
rect 6350 38952 6542 38968
rect 6414 38888 6478 38952
rect 6350 38872 6542 38888
rect 6414 38808 6478 38872
rect 6350 38792 6542 38808
rect 6414 38728 6478 38792
rect 6350 38712 6542 38728
rect 6414 38648 6478 38712
rect 6350 38632 6542 38648
rect 6414 38568 6478 38632
rect 6350 38552 6542 38568
rect 6414 38488 6478 38552
rect 6350 38472 6542 38488
rect 6414 38408 6478 38472
rect 6350 38392 6542 38408
rect 6414 38328 6478 38392
rect 6350 38311 6542 38328
rect 6414 38247 6478 38311
rect 6350 38230 6542 38247
rect 6414 38166 6478 38230
rect 6350 38149 6542 38166
rect 6414 38085 6478 38149
rect 6350 38068 6542 38085
rect 6414 38004 6478 38068
rect 6350 37987 6542 38004
rect 6414 37923 6478 37987
rect 6350 37906 6542 37923
rect 6414 37842 6478 37906
rect 6350 37825 6542 37842
rect 6414 37761 6478 37825
rect 6350 37744 6542 37761
rect 6414 37680 6478 37744
rect 6350 37663 6542 37680
rect 6414 37599 6478 37663
rect 6350 37582 6542 37599
rect 6414 37518 6478 37582
rect 6350 37501 6542 37518
rect 6414 37437 6478 37501
rect 6350 37420 6542 37437
rect 6414 37356 6478 37420
rect 6350 37339 6542 37356
rect 6414 37275 6478 37339
rect 6350 37258 6542 37275
rect 6414 37194 6478 37258
rect 6350 37177 6542 37194
rect 6414 37113 6478 37177
rect 6350 37096 6542 37113
rect 6414 37032 6478 37096
rect 6350 37015 6542 37032
rect 6414 36951 6478 37015
rect 6350 36934 6542 36951
rect 6414 36870 6478 36934
rect 6350 36853 6542 36870
rect 6414 36789 6478 36853
rect 6350 36772 6542 36789
rect 6414 36708 6478 36772
rect 6350 36691 6542 36708
rect 6414 36627 6478 36691
rect 6350 36610 6542 36627
rect 6414 36546 6478 36610
rect 6350 36529 6542 36546
rect 6414 36465 6478 36529
rect 6350 36448 6542 36465
rect 6414 36384 6478 36448
rect 6350 36367 6542 36384
rect 6414 36303 6478 36367
rect 6350 36286 6542 36303
rect 6414 36222 6478 36286
rect 6350 36205 6542 36222
rect 6414 36141 6478 36205
rect 6350 36124 6542 36141
rect 6414 36060 6478 36124
rect 6350 36043 6542 36060
rect 6414 35979 6478 36043
rect 6350 35962 6542 35979
rect 6414 35898 6478 35962
rect 6350 35881 6542 35898
rect 6414 35817 6478 35881
rect 6350 35800 6542 35817
rect 6414 35736 6478 35800
rect 6350 35719 6542 35736
rect 6414 35655 6478 35719
rect 6350 35638 6542 35655
rect 6414 35574 6478 35638
rect 6350 35557 6542 35574
rect 6414 35493 6478 35557
rect 6350 35476 6542 35493
rect 6414 35412 6478 35476
rect 6350 35395 6542 35412
rect 6414 35331 6478 35395
rect 6350 35314 6542 35331
rect 6414 35250 6478 35314
rect 6350 35233 6542 35250
rect 6414 35169 6478 35233
rect 6350 35152 6542 35169
rect 6414 35088 6478 35152
rect 6350 35071 6542 35088
rect 6414 35007 6478 35071
rect 6350 34990 6542 35007
rect 6414 34926 6478 34990
rect 6350 34909 6542 34926
rect 6414 34845 6478 34909
rect 6350 34828 6542 34845
rect 6414 34764 6478 34828
rect 5358 31962 5363 32018
rect 5419 31962 5489 32018
rect 5545 31962 5550 32018
rect 5358 31936 5550 31962
rect 5358 31880 5363 31936
rect 5419 31880 5489 31936
rect 5545 31880 5550 31936
rect 5358 31854 5550 31880
rect 5358 31798 5363 31854
rect 5419 31798 5489 31854
rect 5545 31798 5550 31854
rect 5358 31772 5550 31798
rect 5358 31716 5363 31772
rect 5419 31716 5489 31772
rect 5545 31716 5550 31772
rect 5358 31690 5550 31716
rect 5358 31634 5363 31690
rect 5419 31634 5489 31690
rect 5545 31634 5550 31690
rect 5358 31608 5550 31634
rect 5358 31552 5363 31608
rect 5419 31552 5489 31608
rect 5545 31552 5550 31608
rect 5358 31526 5550 31552
rect 5358 31470 5363 31526
rect 5419 31470 5489 31526
rect 5545 31470 5550 31526
rect 5358 31444 5550 31470
rect 5358 31388 5363 31444
rect 5419 31388 5489 31444
rect 5545 31388 5550 31444
rect 5358 31362 5550 31388
rect 5358 31306 5363 31362
rect 5419 31306 5489 31362
rect 5545 31306 5550 31362
rect 5358 31280 5550 31306
rect 5358 31224 5363 31280
rect 5419 31224 5489 31280
rect 5545 31224 5550 31280
rect 5358 31198 5550 31224
rect 5358 31142 5363 31198
rect 5419 31142 5489 31198
rect 5545 31142 5550 31198
rect 5358 31116 5550 31142
rect 5358 31060 5363 31116
rect 5419 31060 5489 31116
rect 5545 31060 5550 31116
rect 5358 31034 5550 31060
rect 5358 30978 5363 31034
rect 5419 30978 5489 31034
rect 5545 30978 5550 31034
rect 5358 30952 5550 30978
rect 5358 30896 5363 30952
rect 5419 30896 5489 30952
rect 5545 30896 5550 30952
rect 5358 30870 5550 30896
rect 5358 30814 5363 30870
rect 5419 30814 5489 30870
rect 5545 30814 5550 30870
rect 5358 30788 5550 30814
rect 5358 30732 5363 30788
rect 5419 30732 5489 30788
rect 5545 30732 5550 30788
rect 5358 30706 5550 30732
rect 5358 30650 5363 30706
rect 5419 30650 5489 30706
rect 5545 30650 5550 30706
rect 5358 30624 5550 30650
rect 5358 30568 5363 30624
rect 5419 30568 5489 30624
rect 5545 30568 5550 30624
rect 5358 30542 5550 30568
rect 5358 30486 5363 30542
rect 5419 30486 5489 30542
rect 5545 30486 5550 30542
rect 5358 30460 5550 30486
rect 5358 30404 5363 30460
rect 5419 30404 5489 30460
rect 5545 30404 5550 30460
rect 5358 30378 5550 30404
rect 5358 30322 5363 30378
rect 5419 30322 5489 30378
rect 5545 30322 5550 30378
rect 5358 30296 5550 30322
rect 5358 30240 5363 30296
rect 5419 30240 5489 30296
rect 5545 30240 5550 30296
rect 5358 30214 5550 30240
rect 5358 30158 5363 30214
rect 5419 30158 5489 30214
rect 5545 30158 5550 30214
rect 5358 30132 5550 30158
rect 5358 30076 5363 30132
rect 5419 30076 5489 30132
rect 5545 30076 5550 30132
rect 5358 30050 5550 30076
rect 5358 29994 5363 30050
rect 5419 29994 5489 30050
rect 5545 29994 5550 30050
rect 5358 29968 5550 29994
rect 5358 29912 5363 29968
rect 5419 29912 5489 29968
rect 5545 29912 5550 29968
rect 5358 29886 5550 29912
rect 5358 29830 5363 29886
rect 5419 29830 5489 29886
rect 5545 29830 5550 29886
rect 5358 29804 5550 29830
rect 5358 29748 5363 29804
rect 5419 29748 5489 29804
rect 5545 29748 5550 29804
rect 5358 29722 5550 29748
rect 5358 29666 5363 29722
rect 5419 29666 5489 29722
rect 5545 29666 5550 29722
rect 5358 29640 5550 29666
rect 5358 29584 5363 29640
rect 5419 29584 5489 29640
rect 5545 29584 5550 29640
rect 5358 29558 5550 29584
rect 5358 29502 5363 29558
rect 5419 29502 5489 29558
rect 5545 29502 5550 29558
rect 5358 29476 5550 29502
rect 5358 29420 5363 29476
rect 5419 29420 5489 29476
rect 5545 29420 5550 29476
rect 5358 29415 5550 29420
rect 5854 34219 6046 34225
rect 5918 34155 5982 34219
rect 5854 34125 6046 34155
rect 5918 34061 5982 34125
rect 5854 34030 6046 34061
rect 5918 33966 5982 34030
rect 5854 33935 6046 33966
rect 5918 33871 5982 33935
rect 5854 33840 6046 33871
rect 5918 33776 5982 33840
rect 5854 33745 6046 33776
rect 5918 33681 5982 33745
rect 5854 32018 6046 33681
rect 5854 31962 5859 32018
rect 5915 31962 5985 32018
rect 6041 31962 6046 32018
rect 5854 31936 6046 31962
rect 5854 31880 5859 31936
rect 5915 31880 5985 31936
rect 6041 31880 6046 31936
rect 5854 31854 6046 31880
rect 5854 31798 5859 31854
rect 5915 31798 5985 31854
rect 6041 31798 6046 31854
rect 5854 31772 6046 31798
rect 5854 31716 5859 31772
rect 5915 31716 5985 31772
rect 6041 31716 6046 31772
rect 5854 31690 6046 31716
rect 5854 31634 5859 31690
rect 5915 31634 5985 31690
rect 6041 31634 6046 31690
rect 5854 31608 6046 31634
rect 5854 31552 5859 31608
rect 5915 31552 5985 31608
rect 6041 31552 6046 31608
rect 5854 31526 6046 31552
rect 5854 31470 5859 31526
rect 5915 31470 5985 31526
rect 6041 31470 6046 31526
rect 5854 31444 6046 31470
rect 5854 31388 5859 31444
rect 5915 31388 5985 31444
rect 6041 31388 6046 31444
rect 5854 31362 6046 31388
rect 5854 31306 5859 31362
rect 5915 31306 5985 31362
rect 6041 31306 6046 31362
rect 5854 31280 6046 31306
rect 5854 31224 5859 31280
rect 5915 31224 5985 31280
rect 6041 31224 6046 31280
rect 5854 31198 6046 31224
rect 5854 31142 5859 31198
rect 5915 31142 5985 31198
rect 6041 31142 6046 31198
rect 5854 31116 6046 31142
rect 5854 31060 5859 31116
rect 5915 31060 5985 31116
rect 6041 31060 6046 31116
rect 5854 31034 6046 31060
rect 5854 30978 5859 31034
rect 5915 30978 5985 31034
rect 6041 30978 6046 31034
rect 5854 30952 6046 30978
rect 5854 30896 5859 30952
rect 5915 30896 5985 30952
rect 6041 30896 6046 30952
rect 5854 30870 6046 30896
rect 5854 30814 5859 30870
rect 5915 30814 5985 30870
rect 6041 30814 6046 30870
rect 5854 30788 6046 30814
rect 5854 30732 5859 30788
rect 5915 30732 5985 30788
rect 6041 30732 6046 30788
rect 5854 30706 6046 30732
rect 5854 30650 5859 30706
rect 5915 30650 5985 30706
rect 6041 30650 6046 30706
rect 5854 30624 6046 30650
rect 5854 30568 5859 30624
rect 5915 30568 5985 30624
rect 6041 30568 6046 30624
rect 5854 30542 6046 30568
rect 5854 30486 5859 30542
rect 5915 30486 5985 30542
rect 6041 30486 6046 30542
rect 5854 30460 6046 30486
rect 5854 30404 5859 30460
rect 5915 30404 5985 30460
rect 6041 30404 6046 30460
rect 5854 30378 6046 30404
rect 5854 30322 5859 30378
rect 5915 30322 5985 30378
rect 6041 30322 6046 30378
rect 5854 30296 6046 30322
rect 5854 30240 5859 30296
rect 5915 30240 5985 30296
rect 6041 30240 6046 30296
rect 5854 30214 6046 30240
rect 5854 30158 5859 30214
rect 5915 30158 5985 30214
rect 6041 30158 6046 30214
rect 5854 30132 6046 30158
rect 5854 30076 5859 30132
rect 5915 30076 5985 30132
rect 6041 30076 6046 30132
rect 5854 30050 6046 30076
rect 5854 29994 5859 30050
rect 5915 29994 5985 30050
rect 6041 29994 6046 30050
rect 5854 29968 6046 29994
rect 5854 29912 5859 29968
rect 5915 29912 5985 29968
rect 6041 29912 6046 29968
rect 5854 29886 6046 29912
rect 5854 29830 5859 29886
rect 5915 29830 5985 29886
rect 6041 29830 6046 29886
rect 5854 29804 6046 29830
rect 5854 29748 5859 29804
rect 5915 29748 5985 29804
rect 6041 29748 6046 29804
rect 5854 29722 6046 29748
rect 5854 29666 5859 29722
rect 5915 29666 5985 29722
rect 6041 29666 6046 29722
rect 5854 29640 6046 29666
rect 5854 29584 5859 29640
rect 5915 29584 5985 29640
rect 6041 29584 6046 29640
rect 5854 29558 6046 29584
rect 5854 29502 5859 29558
rect 5915 29502 5985 29558
rect 6041 29502 6046 29558
rect 5854 29476 6046 29502
rect 5854 29420 5859 29476
rect 5915 29420 5985 29476
rect 6041 29420 6046 29476
rect 5456 28620 5554 28633
rect 5456 28564 5477 28620
rect 5533 28564 5554 28620
rect 5456 28453 5554 28564
rect 5456 28397 5477 28453
rect 5533 28397 5554 28453
rect 5456 28286 5554 28397
rect 5456 28230 5477 28286
rect 5533 28230 5554 28286
rect 5456 28119 5554 28230
rect 5456 28063 5477 28119
rect 5533 28063 5554 28119
rect 5456 27952 5554 28063
rect 5456 27896 5477 27952
rect 5533 27896 5554 27952
rect 5456 27785 5554 27896
rect 5456 27729 5477 27785
rect 5533 27729 5554 27785
rect 5456 27618 5554 27729
rect 5456 27562 5477 27618
rect 5533 27562 5554 27618
rect 5456 27451 5554 27562
rect 5456 27395 5477 27451
rect 5533 27395 5554 27451
rect 5456 27283 5554 27395
rect 5456 27227 5477 27283
rect 5533 27227 5554 27283
tri 5054 27161 5092 27199 sw
rect 4862 27137 5092 27161
tri 5092 27137 5116 27161 sw
rect 4862 27101 5116 27137
tri 5116 27101 5152 27137 sw
rect 4862 26730 5152 27101
tri 4862 26716 4876 26730 ne
rect 4876 26716 5152 26730
tri 4876 26660 4932 26716 ne
rect 4932 26660 5152 26716
tri 4932 26657 4935 26660 ne
rect 4935 26657 5152 26660
tri 4935 26632 4960 26657 ne
tri 4562 26548 4566 26552 sw
rect 4464 26492 4566 26548
tri 4566 26492 4622 26548 sw
rect 4464 26458 4622 26492
tri 4622 26458 4656 26492 sw
rect 4464 26176 4656 26458
rect 4464 26120 4469 26176
rect 4525 26120 4595 26176
rect 4651 26120 4656 26176
rect 4464 26081 4656 26120
rect 4464 26025 4469 26081
rect 4525 26025 4595 26081
rect 4651 26025 4656 26081
rect 4464 25986 4656 26025
rect 4464 25930 4469 25986
rect 4525 25930 4595 25986
rect 4651 25930 4656 25986
rect 4464 25891 4656 25930
rect 4464 25835 4469 25891
rect 4525 25835 4595 25891
rect 4651 25835 4656 25891
rect 4464 25795 4656 25835
rect 4464 25739 4469 25795
rect 4525 25739 4595 25795
rect 4651 25739 4656 25795
rect 4464 25699 4656 25739
rect 4464 25643 4469 25699
rect 4525 25643 4595 25699
rect 4651 25643 4656 25699
rect 4464 23686 4656 25643
rect 4464 23630 4473 23686
rect 4529 23630 4591 23686
rect 4647 23630 4656 23686
rect 4464 23606 4656 23630
rect 4464 23550 4473 23606
rect 4529 23550 4591 23606
rect 4647 23550 4656 23606
rect 4464 23526 4656 23550
rect 4464 23470 4473 23526
rect 4529 23470 4591 23526
rect 4647 23470 4656 23526
rect 4464 23446 4656 23470
rect 4464 23390 4473 23446
rect 4529 23390 4591 23446
rect 4647 23390 4656 23446
rect 4464 23366 4656 23390
rect 4464 23310 4473 23366
rect 4529 23310 4591 23366
rect 4647 23310 4656 23366
rect 4464 23286 4656 23310
rect 4464 23230 4473 23286
rect 4529 23230 4591 23286
rect 4647 23230 4656 23286
rect 4464 23206 4656 23230
rect 4464 23150 4473 23206
rect 4529 23150 4591 23206
rect 4647 23150 4656 23206
rect 4464 23126 4656 23150
rect 4464 23070 4473 23126
rect 4529 23070 4591 23126
rect 4647 23070 4656 23126
rect 4464 23046 4656 23070
rect 4464 22990 4473 23046
rect 4529 22990 4591 23046
rect 4647 22990 4656 23046
rect 4464 22966 4656 22990
rect 4464 22910 4473 22966
rect 4529 22910 4591 22966
rect 4647 22910 4656 22966
rect 4464 22886 4656 22910
rect 4464 22830 4473 22886
rect 4529 22830 4591 22886
rect 4647 22830 4656 22886
rect 4464 22806 4656 22830
rect 4464 22750 4473 22806
rect 4529 22750 4591 22806
rect 4647 22750 4656 22806
rect 4464 22726 4656 22750
rect 4464 22670 4473 22726
rect 4529 22670 4591 22726
rect 4647 22670 4656 22726
rect 4464 22646 4656 22670
rect 4464 22590 4473 22646
rect 4529 22590 4591 22646
rect 4647 22590 4656 22646
rect 4464 22566 4656 22590
rect 4464 22510 4473 22566
rect 4529 22510 4591 22566
rect 4647 22510 4656 22566
rect 4464 22486 4656 22510
rect 4464 22430 4473 22486
rect 4529 22430 4591 22486
rect 4647 22430 4656 22486
rect 4464 22406 4656 22430
rect 4464 22350 4473 22406
rect 4529 22350 4591 22406
rect 4647 22350 4656 22406
rect 4464 22326 4656 22350
rect 4464 22270 4473 22326
rect 4529 22270 4591 22326
rect 4647 22270 4656 22326
rect 4464 22245 4656 22270
rect 4464 22189 4473 22245
rect 4529 22189 4591 22245
rect 4647 22189 4656 22245
rect 4464 22164 4656 22189
rect 4464 22108 4473 22164
rect 4529 22108 4591 22164
rect 4647 22108 4656 22164
rect 4464 22083 4656 22108
rect 4464 22027 4473 22083
rect 4529 22027 4591 22083
rect 4647 22027 4656 22083
rect 4464 22002 4656 22027
rect 4464 21946 4473 22002
rect 4529 21946 4591 22002
rect 4647 21946 4656 22002
rect 4464 21921 4656 21946
rect 4464 21865 4473 21921
rect 4529 21865 4591 21921
rect 4647 21865 4656 21921
rect 4464 21840 4656 21865
rect 4464 21784 4473 21840
rect 4529 21784 4591 21840
rect 4647 21784 4656 21840
rect 4464 21759 4656 21784
rect 4464 21703 4473 21759
rect 4529 21703 4591 21759
rect 4647 21703 4656 21759
rect 4464 21678 4656 21703
rect 4464 21622 4473 21678
rect 4529 21622 4591 21678
rect 4647 21622 4656 21678
rect 4464 21597 4656 21622
rect 4464 21541 4473 21597
rect 4529 21541 4591 21597
rect 4647 21541 4656 21597
rect 4464 21516 4656 21541
rect 4464 21460 4473 21516
rect 4529 21460 4591 21516
rect 4647 21460 4656 21516
rect 4464 21435 4656 21460
rect 4464 21379 4473 21435
rect 4529 21379 4591 21435
rect 4647 21379 4656 21435
rect 4464 21354 4656 21379
rect 4464 21298 4473 21354
rect 4529 21298 4591 21354
rect 4647 21298 4656 21354
rect 4464 21273 4656 21298
rect 4464 21217 4473 21273
rect 4529 21217 4591 21273
rect 4647 21217 4656 21273
rect 4464 21192 4656 21217
rect 4464 21136 4473 21192
rect 4529 21136 4591 21192
rect 4647 21136 4656 21192
rect 4464 18592 4656 21136
rect 4528 18528 4592 18592
rect 4464 18512 4656 18528
rect 4528 18448 4592 18512
rect 4464 18432 4656 18448
rect 4528 18368 4592 18432
rect 4464 18352 4656 18368
rect 4528 18288 4592 18352
rect 4464 18272 4656 18288
rect 4528 18208 4592 18272
rect 4464 18192 4656 18208
rect 4528 18128 4592 18192
rect 4464 18112 4656 18128
rect 4528 18048 4592 18112
rect 4464 18032 4656 18048
rect 4528 17968 4592 18032
rect 4464 17952 4656 17968
rect 4528 17888 4592 17952
rect 4464 17872 4656 17888
rect 4528 17808 4592 17872
rect 4464 17792 4656 17808
rect 4528 17728 4592 17792
rect 4464 17712 4656 17728
rect 4528 17648 4592 17712
rect 4464 17632 4656 17648
rect 4528 17568 4592 17632
rect 4464 17552 4656 17568
rect 4528 17488 4592 17552
rect 4464 17472 4656 17488
rect 4528 17408 4592 17472
rect 4464 17392 4656 17408
rect 4528 17328 4592 17392
rect 4464 17312 4656 17328
rect 4528 17248 4592 17312
rect 4464 17232 4656 17248
rect 4528 17168 4592 17232
rect 4464 17152 4656 17168
rect 4528 17088 4592 17152
rect 4464 17072 4656 17088
rect 4528 17008 4592 17072
rect 4464 16992 4656 17008
rect 4528 16928 4592 16992
rect 4464 16912 4656 16928
rect 4528 16848 4592 16912
rect 4464 16832 4656 16848
rect 4528 16768 4592 16832
rect 4464 16752 4656 16768
rect 4528 16688 4592 16752
rect 4464 16672 4656 16688
rect 4528 16608 4592 16672
rect 4464 16592 4656 16608
rect 4528 16528 4592 16592
rect 4464 16512 4656 16528
rect 4528 16448 4592 16512
rect 4464 16432 4656 16448
rect 4528 16368 4592 16432
rect 4464 16351 4656 16368
rect 4528 16287 4592 16351
rect 4464 16270 4656 16287
rect 4528 16206 4592 16270
rect 4464 16189 4656 16206
rect 4528 16125 4592 16189
rect 4464 16108 4656 16125
rect 4528 16044 4592 16108
rect 4464 16027 4656 16044
rect 4528 15963 4592 16027
rect 4464 15946 4656 15963
rect 4528 15882 4592 15946
rect 4464 15865 4656 15882
rect 4528 15801 4592 15865
rect 4464 15784 4656 15801
rect 4528 15720 4592 15784
rect 4464 15703 4656 15720
rect 4528 15639 4592 15703
rect 4464 15622 4656 15639
rect 4528 15558 4592 15622
rect 4464 15541 4656 15558
rect 4528 15477 4592 15541
rect 4464 15460 4656 15477
rect 4528 15396 4592 15460
rect 4464 15379 4656 15396
rect 4528 15315 4592 15379
rect 4464 15298 4656 15315
rect 4528 15234 4592 15298
rect 4464 15217 4656 15234
rect 4528 15153 4592 15217
rect 4464 15136 4656 15153
rect 4528 15072 4592 15136
rect 4464 15055 4656 15072
rect 4528 14991 4592 15055
rect 4464 14974 4656 14991
rect 4528 14910 4592 14974
rect 4464 14893 4656 14910
rect 4528 14829 4592 14893
rect 4464 14812 4656 14829
rect 4528 14748 4592 14812
rect 4464 14731 4656 14748
rect 4528 14667 4592 14731
rect 4464 14650 4656 14667
rect 4528 14586 4592 14650
rect 4464 14569 4656 14586
rect 4528 14505 4592 14569
rect 4464 14488 4656 14505
rect 4528 14424 4592 14488
rect 4464 14407 4656 14424
rect 4528 14343 4592 14407
rect 4464 14326 4656 14343
rect 4528 14262 4592 14326
rect 4464 14245 4656 14262
rect 4528 14181 4592 14245
rect 4464 14164 4656 14181
rect 4528 14100 4592 14164
rect 4464 14083 4656 14100
rect 4528 14019 4592 14083
rect 4464 14002 4656 14019
rect 4528 13938 4592 14002
rect 4464 13921 4656 13938
rect 4528 13857 4592 13921
rect 4464 13840 4656 13857
rect 4528 13776 4592 13840
rect 4464 13759 4656 13776
rect 4528 13695 4592 13759
rect 4464 13678 4656 13695
rect 4528 13614 4592 13678
rect 4464 13607 4656 13614
rect 4960 23686 5152 26657
rect 4960 23630 4969 23686
rect 5025 23630 5087 23686
rect 5143 23630 5152 23686
rect 4960 23606 5152 23630
rect 4960 23550 4969 23606
rect 5025 23550 5087 23606
rect 5143 23550 5152 23606
rect 4960 23526 5152 23550
rect 4960 23470 4969 23526
rect 5025 23470 5087 23526
rect 5143 23470 5152 23526
rect 4960 23446 5152 23470
rect 4960 23390 4969 23446
rect 5025 23390 5087 23446
rect 5143 23390 5152 23446
rect 4960 23366 5152 23390
rect 4960 23310 4969 23366
rect 5025 23310 5087 23366
rect 5143 23310 5152 23366
rect 4960 23286 5152 23310
rect 4960 23230 4969 23286
rect 5025 23230 5087 23286
rect 5143 23230 5152 23286
rect 4960 23206 5152 23230
rect 4960 23150 4969 23206
rect 5025 23150 5087 23206
rect 5143 23150 5152 23206
rect 4960 23126 5152 23150
rect 4960 23070 4969 23126
rect 5025 23070 5087 23126
rect 5143 23070 5152 23126
rect 4960 23046 5152 23070
rect 4960 22990 4969 23046
rect 5025 22990 5087 23046
rect 5143 22990 5152 23046
rect 4960 22966 5152 22990
rect 4960 22910 4969 22966
rect 5025 22910 5087 22966
rect 5143 22910 5152 22966
rect 4960 22886 5152 22910
rect 4960 22830 4969 22886
rect 5025 22830 5087 22886
rect 5143 22830 5152 22886
rect 4960 22806 5152 22830
rect 4960 22750 4969 22806
rect 5025 22750 5087 22806
rect 5143 22750 5152 22806
rect 4960 22726 5152 22750
rect 4960 22670 4969 22726
rect 5025 22670 5087 22726
rect 5143 22670 5152 22726
rect 4960 22646 5152 22670
rect 4960 22590 4969 22646
rect 5025 22590 5087 22646
rect 5143 22590 5152 22646
rect 4960 22566 5152 22590
rect 4960 22510 4969 22566
rect 5025 22510 5087 22566
rect 5143 22510 5152 22566
rect 4960 22486 5152 22510
rect 4960 22430 4969 22486
rect 5025 22430 5087 22486
rect 5143 22430 5152 22486
rect 4960 22406 5152 22430
rect 4960 22350 4969 22406
rect 5025 22350 5087 22406
rect 5143 22350 5152 22406
rect 4960 22326 5152 22350
rect 4960 22270 4969 22326
rect 5025 22270 5087 22326
rect 5143 22270 5152 22326
rect 4960 22245 5152 22270
rect 4960 22189 4969 22245
rect 5025 22189 5087 22245
rect 5143 22189 5152 22245
rect 4960 22164 5152 22189
rect 4960 22108 4969 22164
rect 5025 22108 5087 22164
rect 5143 22108 5152 22164
rect 4960 22083 5152 22108
rect 4960 22027 4969 22083
rect 5025 22027 5087 22083
rect 5143 22027 5152 22083
rect 4960 22002 5152 22027
rect 4960 21946 4969 22002
rect 5025 21946 5087 22002
rect 5143 21946 5152 22002
rect 4960 21921 5152 21946
rect 4960 21865 4969 21921
rect 5025 21865 5087 21921
rect 5143 21865 5152 21921
rect 4960 21840 5152 21865
rect 4960 21784 4969 21840
rect 5025 21784 5087 21840
rect 5143 21784 5152 21840
rect 4960 21759 5152 21784
rect 4960 21703 4969 21759
rect 5025 21703 5087 21759
rect 5143 21703 5152 21759
rect 4960 21678 5152 21703
rect 4960 21622 4969 21678
rect 5025 21622 5087 21678
rect 5143 21622 5152 21678
rect 4960 21597 5152 21622
rect 4960 21541 4969 21597
rect 5025 21541 5087 21597
rect 5143 21541 5152 21597
rect 4960 21516 5152 21541
rect 4960 21460 4969 21516
rect 5025 21460 5087 21516
rect 5143 21460 5152 21516
rect 4960 21435 5152 21460
rect 4960 21379 4969 21435
rect 5025 21379 5087 21435
rect 5143 21379 5152 21435
rect 4960 21354 5152 21379
rect 4960 21298 4969 21354
rect 5025 21298 5087 21354
rect 5143 21298 5152 21354
rect 4960 21273 5152 21298
rect 4960 21217 4969 21273
rect 5025 21217 5087 21273
rect 5143 21217 5152 21273
rect 4960 21192 5152 21217
rect 4960 21136 4969 21192
rect 5025 21136 5087 21192
rect 5143 21136 5152 21192
rect 4960 19673 5152 21136
rect 4960 19609 4964 19673
rect 5028 19609 5084 19673
rect 5148 19609 5152 19673
rect 4960 19581 5152 19609
rect 4960 19517 4964 19581
rect 5028 19517 5084 19581
rect 5148 19517 5152 19581
rect 4960 19489 5152 19517
rect 4960 19425 4964 19489
rect 5028 19425 5084 19489
rect 5148 19425 5152 19489
rect 4960 19397 5152 19425
rect 4960 19333 4964 19397
rect 5028 19333 5084 19397
rect 5148 19333 5152 19397
rect 4960 19305 5152 19333
rect 4960 19241 4964 19305
rect 5028 19241 5084 19305
rect 5148 19241 5152 19305
rect 4960 19212 5152 19241
rect 4960 19148 4964 19212
rect 5028 19148 5084 19212
rect 5148 19148 5152 19212
tri 4156 13060 4160 13064 sw
tri 4956 13060 4960 13064 se
rect 4960 13060 5152 19148
rect 5456 26548 5554 27227
rect 5854 27161 6046 29420
rect 6350 32018 6542 34764
rect 7342 39592 7534 39600
rect 7406 39528 7470 39592
rect 7342 39512 7534 39528
rect 7406 39448 7470 39512
rect 7342 39432 7534 39448
rect 7406 39368 7470 39432
rect 7342 39352 7534 39368
rect 7406 39288 7470 39352
rect 7342 39272 7534 39288
rect 7406 39208 7470 39272
rect 7342 39192 7534 39208
rect 7406 39128 7470 39192
rect 7342 39112 7534 39128
rect 7406 39048 7470 39112
rect 7342 39032 7534 39048
rect 7406 38968 7470 39032
rect 7342 38952 7534 38968
rect 7406 38888 7470 38952
rect 7342 38872 7534 38888
rect 7406 38808 7470 38872
rect 7342 38792 7534 38808
rect 7406 38728 7470 38792
rect 7342 38712 7534 38728
rect 7406 38648 7470 38712
rect 7342 38632 7534 38648
rect 7406 38568 7470 38632
rect 7342 38552 7534 38568
rect 7406 38488 7470 38552
rect 7342 38472 7534 38488
rect 7406 38408 7470 38472
rect 7342 38392 7534 38408
rect 7406 38328 7470 38392
rect 7342 38311 7534 38328
rect 7406 38247 7470 38311
rect 7342 38230 7534 38247
rect 7406 38166 7470 38230
rect 7342 38149 7534 38166
rect 7406 38085 7470 38149
rect 7342 38068 7534 38085
rect 7406 38004 7470 38068
rect 7342 37987 7534 38004
rect 7406 37923 7470 37987
rect 7342 37906 7534 37923
rect 7406 37842 7470 37906
rect 7342 37825 7534 37842
rect 7406 37761 7470 37825
rect 7342 37744 7534 37761
rect 7406 37680 7470 37744
rect 7342 37663 7534 37680
rect 7406 37599 7470 37663
rect 7342 37582 7534 37599
rect 7406 37518 7470 37582
rect 7342 37501 7534 37518
rect 7406 37437 7470 37501
rect 7342 37420 7534 37437
rect 7406 37356 7470 37420
rect 7342 37339 7534 37356
rect 7406 37275 7470 37339
rect 7342 37258 7534 37275
rect 7406 37194 7470 37258
rect 7342 37177 7534 37194
rect 7406 37113 7470 37177
rect 7342 37096 7534 37113
rect 7406 37032 7470 37096
rect 7342 37015 7534 37032
rect 7406 36951 7470 37015
rect 7342 36934 7534 36951
rect 7406 36870 7470 36934
rect 7342 36853 7534 36870
rect 7406 36789 7470 36853
rect 7342 36772 7534 36789
rect 7406 36708 7470 36772
rect 7342 36691 7534 36708
rect 7406 36627 7470 36691
rect 7342 36610 7534 36627
rect 7406 36546 7470 36610
rect 7342 36529 7534 36546
rect 7406 36465 7470 36529
rect 7342 36448 7534 36465
rect 7406 36384 7470 36448
rect 7342 36367 7534 36384
rect 7406 36303 7470 36367
rect 7342 36286 7534 36303
rect 7406 36222 7470 36286
rect 7342 36205 7534 36222
rect 7406 36141 7470 36205
rect 7342 36124 7534 36141
rect 7406 36060 7470 36124
rect 7342 36043 7534 36060
rect 7406 35979 7470 36043
rect 7342 35962 7534 35979
rect 7406 35898 7470 35962
rect 7342 35881 7534 35898
rect 7406 35817 7470 35881
rect 7342 35800 7534 35817
rect 7406 35736 7470 35800
rect 7342 35719 7534 35736
rect 7406 35655 7470 35719
rect 7342 35638 7534 35655
rect 7406 35574 7470 35638
rect 7342 35557 7534 35574
rect 7406 35493 7470 35557
rect 7342 35476 7534 35493
rect 7406 35412 7470 35476
rect 7342 35395 7534 35412
rect 7406 35331 7470 35395
rect 7342 35314 7534 35331
rect 7406 35250 7470 35314
rect 7342 35233 7534 35250
rect 7406 35169 7470 35233
rect 7342 35152 7534 35169
rect 7406 35088 7470 35152
rect 7342 35071 7534 35088
rect 7406 35007 7470 35071
rect 7342 34990 7534 35007
rect 7406 34926 7470 34990
rect 7342 34909 7534 34926
rect 7406 34845 7470 34909
rect 7342 34828 7534 34845
rect 7406 34764 7470 34828
rect 6350 31962 6355 32018
rect 6411 31962 6481 32018
rect 6537 31962 6542 32018
rect 6350 31936 6542 31962
rect 6350 31880 6355 31936
rect 6411 31880 6481 31936
rect 6537 31880 6542 31936
rect 6350 31854 6542 31880
rect 6350 31798 6355 31854
rect 6411 31798 6481 31854
rect 6537 31798 6542 31854
rect 6350 31772 6542 31798
rect 6350 31716 6355 31772
rect 6411 31716 6481 31772
rect 6537 31716 6542 31772
rect 6350 31690 6542 31716
rect 6350 31634 6355 31690
rect 6411 31634 6481 31690
rect 6537 31634 6542 31690
rect 6350 31608 6542 31634
rect 6350 31552 6355 31608
rect 6411 31552 6481 31608
rect 6537 31552 6542 31608
rect 6350 31526 6542 31552
rect 6350 31470 6355 31526
rect 6411 31470 6481 31526
rect 6537 31470 6542 31526
rect 6350 31444 6542 31470
rect 6350 31388 6355 31444
rect 6411 31388 6481 31444
rect 6537 31388 6542 31444
rect 6350 31362 6542 31388
rect 6350 31306 6355 31362
rect 6411 31306 6481 31362
rect 6537 31306 6542 31362
rect 6350 31280 6542 31306
rect 6350 31224 6355 31280
rect 6411 31224 6481 31280
rect 6537 31224 6542 31280
rect 6350 31198 6542 31224
rect 6350 31142 6355 31198
rect 6411 31142 6481 31198
rect 6537 31142 6542 31198
rect 6350 31116 6542 31142
rect 6350 31060 6355 31116
rect 6411 31060 6481 31116
rect 6537 31060 6542 31116
rect 6350 31034 6542 31060
rect 6350 30978 6355 31034
rect 6411 30978 6481 31034
rect 6537 30978 6542 31034
rect 6350 30952 6542 30978
rect 6350 30896 6355 30952
rect 6411 30896 6481 30952
rect 6537 30896 6542 30952
rect 6350 30870 6542 30896
rect 6350 30814 6355 30870
rect 6411 30814 6481 30870
rect 6537 30814 6542 30870
rect 6350 30788 6542 30814
rect 6350 30732 6355 30788
rect 6411 30732 6481 30788
rect 6537 30732 6542 30788
rect 6350 30706 6542 30732
rect 6350 30650 6355 30706
rect 6411 30650 6481 30706
rect 6537 30650 6542 30706
rect 6350 30624 6542 30650
rect 6350 30568 6355 30624
rect 6411 30568 6481 30624
rect 6537 30568 6542 30624
rect 6350 30542 6542 30568
rect 6350 30486 6355 30542
rect 6411 30486 6481 30542
rect 6537 30486 6542 30542
rect 6350 30460 6542 30486
rect 6350 30404 6355 30460
rect 6411 30404 6481 30460
rect 6537 30404 6542 30460
rect 6350 30378 6542 30404
rect 6350 30322 6355 30378
rect 6411 30322 6481 30378
rect 6537 30322 6542 30378
rect 6350 30296 6542 30322
rect 6350 30240 6355 30296
rect 6411 30240 6481 30296
rect 6537 30240 6542 30296
rect 6350 30214 6542 30240
rect 6350 30158 6355 30214
rect 6411 30158 6481 30214
rect 6537 30158 6542 30214
rect 6350 30132 6542 30158
rect 6350 30076 6355 30132
rect 6411 30076 6481 30132
rect 6537 30076 6542 30132
rect 6350 30050 6542 30076
rect 6350 29994 6355 30050
rect 6411 29994 6481 30050
rect 6537 29994 6542 30050
rect 6350 29968 6542 29994
rect 6350 29912 6355 29968
rect 6411 29912 6481 29968
rect 6537 29912 6542 29968
rect 6350 29886 6542 29912
rect 6350 29830 6355 29886
rect 6411 29830 6481 29886
rect 6537 29830 6542 29886
rect 6350 29804 6542 29830
rect 6350 29748 6355 29804
rect 6411 29748 6481 29804
rect 6537 29748 6542 29804
rect 6350 29722 6542 29748
rect 6350 29666 6355 29722
rect 6411 29666 6481 29722
rect 6537 29666 6542 29722
rect 6350 29640 6542 29666
rect 6350 29584 6355 29640
rect 6411 29584 6481 29640
rect 6537 29584 6542 29640
rect 6350 29558 6542 29584
rect 6350 29502 6355 29558
rect 6411 29502 6481 29558
rect 6537 29502 6542 29558
rect 6350 29476 6542 29502
rect 6350 29420 6355 29476
rect 6411 29420 6481 29476
rect 6537 29420 6542 29476
rect 6350 29415 6542 29420
rect 6846 34219 7042 34225
rect 6910 34155 6974 34219
rect 7038 34155 7042 34219
rect 6846 34125 7042 34155
rect 6910 34061 6974 34125
rect 7038 34061 7042 34125
rect 6846 34030 7042 34061
rect 6910 33966 6974 34030
rect 7038 33966 7042 34030
rect 6846 33935 7042 33966
rect 6910 33871 6974 33935
rect 7038 33871 7042 33935
rect 6846 33840 7042 33871
rect 6910 33776 6974 33840
rect 7038 33776 7042 33840
rect 6846 33745 7042 33776
rect 6910 33681 6974 33745
rect 7038 33681 7042 33745
rect 6846 32018 7042 33681
rect 6846 31962 6851 32018
rect 6907 31962 6977 32018
rect 7033 31962 7042 32018
rect 6846 31936 7042 31962
rect 6846 31880 6851 31936
rect 6907 31880 6977 31936
rect 7033 31880 7042 31936
rect 6846 31854 7042 31880
rect 6846 31798 6851 31854
rect 6907 31798 6977 31854
rect 7033 31798 7042 31854
rect 6846 31772 7042 31798
rect 6846 31716 6851 31772
rect 6907 31716 6977 31772
rect 7033 31716 7042 31772
rect 6846 31690 7042 31716
rect 6846 31634 6851 31690
rect 6907 31634 6977 31690
rect 7033 31634 7042 31690
rect 6846 31608 7042 31634
rect 6846 31552 6851 31608
rect 6907 31552 6977 31608
rect 7033 31552 7042 31608
rect 6846 31526 7042 31552
rect 6846 31470 6851 31526
rect 6907 31470 6977 31526
rect 7033 31470 7042 31526
rect 6846 31444 7042 31470
rect 6846 31388 6851 31444
rect 6907 31388 6977 31444
rect 7033 31388 7042 31444
rect 6846 31362 7042 31388
rect 6846 31306 6851 31362
rect 6907 31306 6977 31362
rect 7033 31306 7042 31362
rect 6846 31280 7042 31306
rect 6846 31224 6851 31280
rect 6907 31224 6977 31280
rect 7033 31224 7042 31280
rect 6846 31198 7042 31224
rect 6846 31142 6851 31198
rect 6907 31142 6977 31198
rect 7033 31142 7042 31198
rect 6846 31116 7042 31142
rect 6846 31060 6851 31116
rect 6907 31060 6977 31116
rect 7033 31060 7042 31116
rect 6846 31034 7042 31060
rect 6846 30978 6851 31034
rect 6907 30978 6977 31034
rect 7033 30978 7042 31034
rect 6846 30952 7042 30978
rect 6846 30896 6851 30952
rect 6907 30896 6977 30952
rect 7033 30896 7042 30952
rect 6846 30870 7042 30896
rect 6846 30814 6851 30870
rect 6907 30814 6977 30870
rect 7033 30814 7042 30870
rect 6846 30788 7042 30814
rect 6846 30732 6851 30788
rect 6907 30732 6977 30788
rect 7033 30732 7042 30788
rect 6846 30706 7042 30732
rect 6846 30650 6851 30706
rect 6907 30650 6977 30706
rect 7033 30650 7042 30706
rect 6846 30624 7042 30650
rect 6846 30568 6851 30624
rect 6907 30568 6977 30624
rect 7033 30568 7042 30624
rect 6846 30542 7042 30568
rect 6846 30486 6851 30542
rect 6907 30486 6977 30542
rect 7033 30486 7042 30542
rect 6846 30460 7042 30486
rect 6846 30404 6851 30460
rect 6907 30404 6977 30460
rect 7033 30404 7042 30460
rect 6846 30378 7042 30404
rect 6846 30322 6851 30378
rect 6907 30322 6977 30378
rect 7033 30322 7042 30378
rect 6846 30296 7042 30322
rect 6846 30240 6851 30296
rect 6907 30240 6977 30296
rect 7033 30240 7042 30296
rect 6846 30214 7042 30240
rect 6846 30158 6851 30214
rect 6907 30158 6977 30214
rect 7033 30158 7042 30214
rect 6846 30132 7042 30158
rect 6846 30076 6851 30132
rect 6907 30076 6977 30132
rect 7033 30076 7042 30132
rect 6846 30050 7042 30076
rect 6846 29994 6851 30050
rect 6907 29994 6977 30050
rect 7033 29994 7042 30050
rect 6846 29968 7042 29994
rect 6846 29912 6851 29968
rect 6907 29912 6977 29968
rect 7033 29912 7042 29968
rect 6846 29886 7042 29912
rect 6846 29830 6851 29886
rect 6907 29830 6977 29886
rect 7033 29830 7042 29886
rect 6846 29804 7042 29830
rect 6846 29748 6851 29804
rect 6907 29748 6977 29804
rect 7033 29748 7042 29804
rect 6846 29722 7042 29748
rect 6846 29666 6851 29722
rect 6907 29666 6977 29722
rect 7033 29666 7042 29722
rect 6846 29640 7042 29666
rect 6846 29584 6851 29640
rect 6907 29584 6977 29640
rect 7033 29584 7042 29640
rect 6846 29558 7042 29584
rect 6846 29502 6851 29558
rect 6907 29502 6977 29558
rect 7033 29502 7042 29558
rect 6846 29476 7042 29502
rect 6846 29420 6851 29476
rect 6907 29420 6977 29476
rect 7033 29420 7042 29476
rect 6448 28620 6546 28633
rect 6448 28564 6469 28620
rect 6525 28564 6546 28620
rect 6448 28453 6546 28564
rect 6448 28397 6469 28453
rect 6525 28397 6546 28453
rect 6448 28286 6546 28397
rect 6448 28230 6469 28286
rect 6525 28230 6546 28286
rect 6448 28119 6546 28230
rect 6448 28063 6469 28119
rect 6525 28063 6546 28119
rect 6448 27952 6546 28063
rect 6448 27896 6469 27952
rect 6525 27896 6546 27952
rect 6448 27785 6546 27896
rect 6448 27729 6469 27785
rect 6525 27729 6546 27785
rect 6448 27618 6546 27729
rect 6448 27562 6469 27618
rect 6525 27562 6546 27618
rect 6448 27451 6546 27562
rect 6448 27395 6469 27451
rect 6525 27395 6546 27451
rect 6448 27283 6546 27395
rect 6448 27227 6469 27283
rect 6525 27227 6546 27283
tri 6046 27161 6080 27195 sw
rect 5854 27137 6080 27161
tri 6080 27137 6104 27161 sw
rect 5854 27097 6104 27137
tri 6104 27097 6144 27137 sw
rect 5854 26726 6144 27097
tri 5854 26716 5864 26726 ne
rect 5864 26716 6144 26726
tri 5864 26660 5920 26716 ne
rect 5920 26660 6144 26716
tri 5920 26657 5923 26660 ne
rect 5923 26657 6144 26660
tri 5923 26632 5948 26657 ne
rect 5948 26632 6144 26657
tri 5948 26628 5952 26632 ne
tri 5554 26548 5558 26552 sw
rect 5456 26492 5558 26548
tri 5558 26492 5614 26548 sw
rect 5456 26458 5614 26492
tri 5614 26458 5648 26492 sw
rect 5456 26176 5648 26458
rect 5456 26120 5461 26176
rect 5517 26120 5587 26176
rect 5643 26120 5648 26176
rect 5456 26081 5648 26120
rect 5456 26025 5461 26081
rect 5517 26025 5587 26081
rect 5643 26025 5648 26081
rect 5456 25986 5648 26025
rect 5456 25930 5461 25986
rect 5517 25930 5587 25986
rect 5643 25930 5648 25986
rect 5456 25891 5648 25930
rect 5456 25835 5461 25891
rect 5517 25835 5587 25891
rect 5643 25835 5648 25891
rect 5456 25795 5648 25835
rect 5456 25739 5461 25795
rect 5517 25739 5587 25795
rect 5643 25739 5648 25795
rect 5456 25699 5648 25739
rect 5456 25643 5461 25699
rect 5517 25643 5587 25699
rect 5643 25643 5648 25699
rect 5456 23686 5648 25643
rect 5456 23630 5465 23686
rect 5521 23630 5583 23686
rect 5639 23630 5648 23686
rect 5456 23606 5648 23630
rect 5456 23550 5465 23606
rect 5521 23550 5583 23606
rect 5639 23550 5648 23606
rect 5456 23526 5648 23550
rect 5456 23470 5465 23526
rect 5521 23470 5583 23526
rect 5639 23470 5648 23526
rect 5456 23446 5648 23470
rect 5456 23390 5465 23446
rect 5521 23390 5583 23446
rect 5639 23390 5648 23446
rect 5456 23366 5648 23390
rect 5456 23310 5465 23366
rect 5521 23310 5583 23366
rect 5639 23310 5648 23366
rect 5456 23286 5648 23310
rect 5456 23230 5465 23286
rect 5521 23230 5583 23286
rect 5639 23230 5648 23286
rect 5456 23206 5648 23230
rect 5456 23150 5465 23206
rect 5521 23150 5583 23206
rect 5639 23150 5648 23206
rect 5456 23126 5648 23150
rect 5456 23070 5465 23126
rect 5521 23070 5583 23126
rect 5639 23070 5648 23126
rect 5456 23046 5648 23070
rect 5456 22990 5465 23046
rect 5521 22990 5583 23046
rect 5639 22990 5648 23046
rect 5456 22966 5648 22990
rect 5456 22910 5465 22966
rect 5521 22910 5583 22966
rect 5639 22910 5648 22966
rect 5456 22886 5648 22910
rect 5456 22830 5465 22886
rect 5521 22830 5583 22886
rect 5639 22830 5648 22886
rect 5456 22806 5648 22830
rect 5456 22750 5465 22806
rect 5521 22750 5583 22806
rect 5639 22750 5648 22806
rect 5456 22726 5648 22750
rect 5456 22670 5465 22726
rect 5521 22670 5583 22726
rect 5639 22670 5648 22726
rect 5456 22646 5648 22670
rect 5456 22590 5465 22646
rect 5521 22590 5583 22646
rect 5639 22590 5648 22646
rect 5456 22566 5648 22590
rect 5456 22510 5465 22566
rect 5521 22510 5583 22566
rect 5639 22510 5648 22566
rect 5456 22486 5648 22510
rect 5456 22430 5465 22486
rect 5521 22430 5583 22486
rect 5639 22430 5648 22486
rect 5456 22406 5648 22430
rect 5456 22350 5465 22406
rect 5521 22350 5583 22406
rect 5639 22350 5648 22406
rect 5456 22326 5648 22350
rect 5456 22270 5465 22326
rect 5521 22270 5583 22326
rect 5639 22270 5648 22326
rect 5456 22245 5648 22270
rect 5456 22189 5465 22245
rect 5521 22189 5583 22245
rect 5639 22189 5648 22245
rect 5456 22164 5648 22189
rect 5456 22108 5465 22164
rect 5521 22108 5583 22164
rect 5639 22108 5648 22164
rect 5456 22083 5648 22108
rect 5456 22027 5465 22083
rect 5521 22027 5583 22083
rect 5639 22027 5648 22083
rect 5456 22002 5648 22027
rect 5456 21946 5465 22002
rect 5521 21946 5583 22002
rect 5639 21946 5648 22002
rect 5456 21921 5648 21946
rect 5456 21865 5465 21921
rect 5521 21865 5583 21921
rect 5639 21865 5648 21921
rect 5456 21840 5648 21865
rect 5456 21784 5465 21840
rect 5521 21784 5583 21840
rect 5639 21784 5648 21840
rect 5456 21759 5648 21784
rect 5456 21703 5465 21759
rect 5521 21703 5583 21759
rect 5639 21703 5648 21759
rect 5456 21678 5648 21703
rect 5456 21622 5465 21678
rect 5521 21622 5583 21678
rect 5639 21622 5648 21678
rect 5456 21597 5648 21622
rect 5456 21541 5465 21597
rect 5521 21541 5583 21597
rect 5639 21541 5648 21597
rect 5456 21516 5648 21541
rect 5456 21460 5465 21516
rect 5521 21460 5583 21516
rect 5639 21460 5648 21516
rect 5456 21435 5648 21460
rect 5456 21379 5465 21435
rect 5521 21379 5583 21435
rect 5639 21379 5648 21435
rect 5456 21354 5648 21379
rect 5456 21298 5465 21354
rect 5521 21298 5583 21354
rect 5639 21298 5648 21354
rect 5456 21273 5648 21298
rect 5456 21217 5465 21273
rect 5521 21217 5583 21273
rect 5639 21217 5648 21273
rect 5456 21192 5648 21217
rect 5456 21136 5465 21192
rect 5521 21136 5583 21192
rect 5639 21136 5648 21192
rect 5456 18592 5648 21136
rect 5520 18528 5584 18592
rect 5456 18512 5648 18528
rect 5520 18448 5584 18512
rect 5456 18432 5648 18448
rect 5520 18368 5584 18432
rect 5456 18352 5648 18368
rect 5520 18288 5584 18352
rect 5456 18272 5648 18288
rect 5520 18208 5584 18272
rect 5456 18192 5648 18208
rect 5520 18128 5584 18192
rect 5456 18112 5648 18128
rect 5520 18048 5584 18112
rect 5456 18032 5648 18048
rect 5520 17968 5584 18032
rect 5456 17952 5648 17968
rect 5520 17888 5584 17952
rect 5456 17872 5648 17888
rect 5520 17808 5584 17872
rect 5456 17792 5648 17808
rect 5520 17728 5584 17792
rect 5456 17712 5648 17728
rect 5520 17648 5584 17712
rect 5456 17632 5648 17648
rect 5520 17568 5584 17632
rect 5456 17552 5648 17568
rect 5520 17488 5584 17552
rect 5456 17472 5648 17488
rect 5520 17408 5584 17472
rect 5456 17392 5648 17408
rect 5520 17328 5584 17392
rect 5456 17312 5648 17328
rect 5520 17248 5584 17312
rect 5456 17232 5648 17248
rect 5520 17168 5584 17232
rect 5456 17152 5648 17168
rect 5520 17088 5584 17152
rect 5456 17072 5648 17088
rect 5520 17008 5584 17072
rect 5456 16992 5648 17008
rect 5520 16928 5584 16992
rect 5456 16912 5648 16928
rect 5520 16848 5584 16912
rect 5456 16832 5648 16848
rect 5520 16768 5584 16832
rect 5456 16752 5648 16768
rect 5520 16688 5584 16752
rect 5456 16672 5648 16688
rect 5520 16608 5584 16672
rect 5456 16592 5648 16608
rect 5520 16528 5584 16592
rect 5456 16512 5648 16528
rect 5520 16448 5584 16512
rect 5456 16431 5648 16448
rect 5520 16367 5584 16431
rect 5456 16350 5648 16367
rect 5520 16286 5584 16350
rect 5456 16269 5648 16286
rect 5520 16205 5584 16269
rect 5456 16188 5648 16205
rect 5520 16124 5584 16188
rect 5456 16107 5648 16124
rect 5520 16043 5584 16107
rect 5456 16026 5648 16043
rect 5520 15962 5584 16026
rect 5456 15945 5648 15962
rect 5520 15881 5584 15945
rect 5456 15864 5648 15881
rect 5520 15800 5584 15864
rect 5456 15783 5648 15800
rect 5520 15719 5584 15783
rect 5456 15702 5648 15719
rect 5520 15638 5584 15702
rect 5456 15621 5648 15638
rect 5520 15557 5584 15621
rect 5456 15540 5648 15557
rect 5520 15476 5584 15540
rect 5456 15459 5648 15476
rect 5520 15395 5584 15459
rect 5456 15378 5648 15395
rect 5520 15314 5584 15378
rect 5456 15297 5648 15314
rect 5520 15233 5584 15297
rect 5456 15216 5648 15233
rect 5520 15152 5584 15216
rect 5456 15135 5648 15152
rect 5520 15071 5584 15135
rect 5456 15054 5648 15071
rect 5520 14990 5584 15054
rect 5456 14973 5648 14990
rect 5520 14909 5584 14973
rect 5456 14892 5648 14909
rect 5520 14828 5584 14892
rect 5456 14811 5648 14828
rect 5520 14747 5584 14811
rect 5456 14730 5648 14747
rect 5520 14666 5584 14730
rect 5456 14649 5648 14666
rect 5520 14585 5584 14649
rect 5456 14568 5648 14585
rect 5520 14504 5584 14568
rect 5456 14487 5648 14504
rect 5520 14423 5584 14487
rect 5456 14406 5648 14423
rect 5520 14342 5584 14406
rect 5456 14325 5648 14342
rect 5520 14261 5584 14325
rect 5456 14244 5648 14261
rect 5520 14180 5584 14244
rect 5456 14163 5648 14180
rect 5520 14099 5584 14163
rect 5456 14082 5648 14099
rect 5520 14018 5584 14082
rect 5456 14001 5648 14018
rect 5520 13937 5584 14001
rect 5456 13920 5648 13937
rect 5520 13856 5584 13920
rect 5456 13839 5648 13856
rect 5520 13775 5584 13839
rect 5456 13758 5648 13775
rect 5520 13694 5584 13758
rect 5456 13677 5648 13694
rect 5520 13613 5584 13677
rect 5456 13607 5648 13613
rect 5952 23686 6144 26632
rect 5952 23630 5961 23686
rect 6017 23630 6079 23686
rect 6135 23630 6144 23686
rect 5952 23606 6144 23630
rect 5952 23550 5961 23606
rect 6017 23550 6079 23606
rect 6135 23550 6144 23606
rect 5952 23526 6144 23550
rect 5952 23470 5961 23526
rect 6017 23470 6079 23526
rect 6135 23470 6144 23526
rect 5952 23446 6144 23470
rect 5952 23390 5961 23446
rect 6017 23390 6079 23446
rect 6135 23390 6144 23446
rect 5952 23366 6144 23390
rect 5952 23310 5961 23366
rect 6017 23310 6079 23366
rect 6135 23310 6144 23366
rect 5952 23286 6144 23310
rect 5952 23230 5961 23286
rect 6017 23230 6079 23286
rect 6135 23230 6144 23286
rect 5952 23206 6144 23230
rect 5952 23150 5961 23206
rect 6017 23150 6079 23206
rect 6135 23150 6144 23206
rect 5952 23126 6144 23150
rect 5952 23070 5961 23126
rect 6017 23070 6079 23126
rect 6135 23070 6144 23126
rect 5952 23046 6144 23070
rect 5952 22990 5961 23046
rect 6017 22990 6079 23046
rect 6135 22990 6144 23046
rect 5952 22966 6144 22990
rect 5952 22910 5961 22966
rect 6017 22910 6079 22966
rect 6135 22910 6144 22966
rect 5952 22886 6144 22910
rect 5952 22830 5961 22886
rect 6017 22830 6079 22886
rect 6135 22830 6144 22886
rect 5952 22806 6144 22830
rect 5952 22750 5961 22806
rect 6017 22750 6079 22806
rect 6135 22750 6144 22806
rect 5952 22726 6144 22750
rect 5952 22670 5961 22726
rect 6017 22670 6079 22726
rect 6135 22670 6144 22726
rect 5952 22646 6144 22670
rect 5952 22590 5961 22646
rect 6017 22590 6079 22646
rect 6135 22590 6144 22646
rect 5952 22566 6144 22590
rect 5952 22510 5961 22566
rect 6017 22510 6079 22566
rect 6135 22510 6144 22566
rect 5952 22486 6144 22510
rect 5952 22430 5961 22486
rect 6017 22430 6079 22486
rect 6135 22430 6144 22486
rect 5952 22406 6144 22430
rect 5952 22350 5961 22406
rect 6017 22350 6079 22406
rect 6135 22350 6144 22406
rect 5952 22326 6144 22350
rect 5952 22270 5961 22326
rect 6017 22270 6079 22326
rect 6135 22270 6144 22326
rect 5952 22245 6144 22270
rect 5952 22189 5961 22245
rect 6017 22189 6079 22245
rect 6135 22189 6144 22245
rect 5952 22164 6144 22189
rect 5952 22108 5961 22164
rect 6017 22108 6079 22164
rect 6135 22108 6144 22164
rect 5952 22083 6144 22108
rect 5952 22027 5961 22083
rect 6017 22027 6079 22083
rect 6135 22027 6144 22083
rect 5952 22002 6144 22027
rect 5952 21946 5961 22002
rect 6017 21946 6079 22002
rect 6135 21946 6144 22002
rect 5952 21921 6144 21946
rect 5952 21865 5961 21921
rect 6017 21865 6079 21921
rect 6135 21865 6144 21921
rect 5952 21840 6144 21865
rect 5952 21784 5961 21840
rect 6017 21784 6079 21840
rect 6135 21784 6144 21840
rect 5952 21759 6144 21784
rect 5952 21703 5961 21759
rect 6017 21703 6079 21759
rect 6135 21703 6144 21759
rect 5952 21678 6144 21703
rect 5952 21622 5961 21678
rect 6017 21622 6079 21678
rect 6135 21622 6144 21678
rect 5952 21597 6144 21622
rect 5952 21541 5961 21597
rect 6017 21541 6079 21597
rect 6135 21541 6144 21597
rect 5952 21516 6144 21541
rect 5952 21460 5961 21516
rect 6017 21460 6079 21516
rect 6135 21460 6144 21516
rect 5952 21435 6144 21460
rect 5952 21379 5961 21435
rect 6017 21379 6079 21435
rect 6135 21379 6144 21435
rect 5952 21354 6144 21379
rect 5952 21298 5961 21354
rect 6017 21298 6079 21354
rect 6135 21298 6144 21354
rect 5952 21273 6144 21298
rect 5952 21217 5961 21273
rect 6017 21217 6079 21273
rect 6135 21217 6144 21273
rect 5952 21192 6144 21217
rect 5952 21136 5961 21192
rect 6017 21136 6079 21192
rect 6135 21136 6144 21192
rect 5952 19673 6144 21136
rect 5952 19609 5953 19673
rect 6017 19609 6073 19673
rect 6137 19609 6144 19673
rect 5952 19581 6144 19609
rect 5952 19517 5953 19581
rect 6017 19517 6073 19581
rect 6137 19517 6144 19581
rect 5952 19489 6144 19517
rect 5952 19425 5953 19489
rect 6017 19425 6073 19489
rect 6137 19425 6144 19489
rect 5952 19397 6144 19425
rect 5952 19333 5953 19397
rect 6017 19333 6073 19397
rect 6137 19333 6144 19397
rect 5952 19305 6144 19333
rect 5952 19241 5953 19305
rect 6017 19241 6073 19305
rect 6137 19241 6144 19305
rect 5952 19212 6144 19241
rect 5952 19148 5953 19212
rect 6017 19148 6073 19212
rect 6137 19148 6144 19212
tri 5948 13060 5952 13064 se
rect 5952 13060 6144 19148
rect 6448 26548 6546 27227
rect 6846 27161 7042 29420
rect 7342 32018 7534 34764
rect 8334 39592 8526 39600
rect 8398 39528 8462 39592
rect 8334 39512 8526 39528
rect 8398 39448 8462 39512
rect 8334 39432 8526 39448
rect 8398 39368 8462 39432
rect 8334 39352 8526 39368
rect 8398 39288 8462 39352
rect 8334 39272 8526 39288
rect 8398 39208 8462 39272
rect 8334 39192 8526 39208
rect 8398 39128 8462 39192
rect 8334 39112 8526 39128
rect 8398 39048 8462 39112
rect 8334 39032 8526 39048
rect 8398 38968 8462 39032
rect 8334 38952 8526 38968
rect 8398 38888 8462 38952
rect 8334 38872 8526 38888
rect 8398 38808 8462 38872
rect 8334 38792 8526 38808
rect 8398 38728 8462 38792
rect 8334 38712 8526 38728
rect 8398 38648 8462 38712
rect 8334 38632 8526 38648
rect 8398 38568 8462 38632
rect 8334 38552 8526 38568
rect 8398 38488 8462 38552
rect 8334 38472 8526 38488
rect 8398 38408 8462 38472
rect 8334 38392 8526 38408
rect 8398 38328 8462 38392
rect 8334 38311 8526 38328
rect 8398 38247 8462 38311
rect 8334 38230 8526 38247
rect 8398 38166 8462 38230
rect 8334 38149 8526 38166
rect 8398 38085 8462 38149
rect 8334 38068 8526 38085
rect 8398 38004 8462 38068
rect 8334 37987 8526 38004
rect 8398 37923 8462 37987
rect 8334 37906 8526 37923
rect 8398 37842 8462 37906
rect 8334 37825 8526 37842
rect 8398 37761 8462 37825
rect 8334 37744 8526 37761
rect 8398 37680 8462 37744
rect 8334 37663 8526 37680
rect 8398 37599 8462 37663
rect 8334 37582 8526 37599
rect 8398 37518 8462 37582
rect 8334 37501 8526 37518
rect 8398 37437 8462 37501
rect 8334 37420 8526 37437
rect 8398 37356 8462 37420
rect 8334 37339 8526 37356
rect 8398 37275 8462 37339
rect 8334 37258 8526 37275
rect 8398 37194 8462 37258
rect 8334 37177 8526 37194
rect 8398 37113 8462 37177
rect 8334 37096 8526 37113
rect 8398 37032 8462 37096
rect 8334 37015 8526 37032
rect 8398 36951 8462 37015
rect 8334 36934 8526 36951
rect 8398 36870 8462 36934
rect 8334 36853 8526 36870
rect 8398 36789 8462 36853
rect 8334 36772 8526 36789
rect 8398 36708 8462 36772
rect 8334 36691 8526 36708
rect 8398 36627 8462 36691
rect 8334 36610 8526 36627
rect 8398 36546 8462 36610
rect 8334 36529 8526 36546
rect 8398 36465 8462 36529
rect 8334 36448 8526 36465
rect 8398 36384 8462 36448
rect 8334 36367 8526 36384
rect 8398 36303 8462 36367
rect 8334 36286 8526 36303
rect 8398 36222 8462 36286
rect 8334 36205 8526 36222
rect 8398 36141 8462 36205
rect 8334 36124 8526 36141
rect 8398 36060 8462 36124
rect 8334 36043 8526 36060
rect 8398 35979 8462 36043
rect 8334 35962 8526 35979
rect 8398 35898 8462 35962
rect 8334 35881 8526 35898
rect 8398 35817 8462 35881
rect 8334 35800 8526 35817
rect 8398 35736 8462 35800
rect 8334 35719 8526 35736
rect 8398 35655 8462 35719
rect 8334 35638 8526 35655
rect 8398 35574 8462 35638
rect 8334 35557 8526 35574
rect 8398 35493 8462 35557
rect 8334 35476 8526 35493
rect 8398 35412 8462 35476
rect 8334 35395 8526 35412
rect 8398 35331 8462 35395
rect 8334 35314 8526 35331
rect 8398 35250 8462 35314
rect 8334 35233 8526 35250
rect 8398 35169 8462 35233
rect 8334 35152 8526 35169
rect 8398 35088 8462 35152
rect 8334 35071 8526 35088
rect 8398 35007 8462 35071
rect 8334 34990 8526 35007
rect 8398 34926 8462 34990
rect 8334 34909 8526 34926
rect 8398 34845 8462 34909
rect 8334 34828 8526 34845
rect 8398 34764 8462 34828
rect 7342 31962 7347 32018
rect 7403 31962 7473 32018
rect 7529 31962 7534 32018
rect 7342 31936 7534 31962
rect 7342 31880 7347 31936
rect 7403 31880 7473 31936
rect 7529 31880 7534 31936
rect 7342 31854 7534 31880
rect 7342 31798 7347 31854
rect 7403 31798 7473 31854
rect 7529 31798 7534 31854
rect 7342 31772 7534 31798
rect 7342 31716 7347 31772
rect 7403 31716 7473 31772
rect 7529 31716 7534 31772
rect 7342 31690 7534 31716
rect 7342 31634 7347 31690
rect 7403 31634 7473 31690
rect 7529 31634 7534 31690
rect 7342 31608 7534 31634
rect 7342 31552 7347 31608
rect 7403 31552 7473 31608
rect 7529 31552 7534 31608
rect 7342 31526 7534 31552
rect 7342 31470 7347 31526
rect 7403 31470 7473 31526
rect 7529 31470 7534 31526
rect 7342 31444 7534 31470
rect 7342 31388 7347 31444
rect 7403 31388 7473 31444
rect 7529 31388 7534 31444
rect 7342 31362 7534 31388
rect 7342 31306 7347 31362
rect 7403 31306 7473 31362
rect 7529 31306 7534 31362
rect 7342 31280 7534 31306
rect 7342 31224 7347 31280
rect 7403 31224 7473 31280
rect 7529 31224 7534 31280
rect 7342 31198 7534 31224
rect 7342 31142 7347 31198
rect 7403 31142 7473 31198
rect 7529 31142 7534 31198
rect 7342 31116 7534 31142
rect 7342 31060 7347 31116
rect 7403 31060 7473 31116
rect 7529 31060 7534 31116
rect 7342 31034 7534 31060
rect 7342 30978 7347 31034
rect 7403 30978 7473 31034
rect 7529 30978 7534 31034
rect 7342 30952 7534 30978
rect 7342 30896 7347 30952
rect 7403 30896 7473 30952
rect 7529 30896 7534 30952
rect 7342 30870 7534 30896
rect 7342 30814 7347 30870
rect 7403 30814 7473 30870
rect 7529 30814 7534 30870
rect 7342 30788 7534 30814
rect 7342 30732 7347 30788
rect 7403 30732 7473 30788
rect 7529 30732 7534 30788
rect 7342 30706 7534 30732
rect 7342 30650 7347 30706
rect 7403 30650 7473 30706
rect 7529 30650 7534 30706
rect 7342 30624 7534 30650
rect 7342 30568 7347 30624
rect 7403 30568 7473 30624
rect 7529 30568 7534 30624
rect 7342 30542 7534 30568
rect 7342 30486 7347 30542
rect 7403 30486 7473 30542
rect 7529 30486 7534 30542
rect 7342 30460 7534 30486
rect 7342 30404 7347 30460
rect 7403 30404 7473 30460
rect 7529 30404 7534 30460
rect 7342 30378 7534 30404
rect 7342 30322 7347 30378
rect 7403 30322 7473 30378
rect 7529 30322 7534 30378
rect 7342 30296 7534 30322
rect 7342 30240 7347 30296
rect 7403 30240 7473 30296
rect 7529 30240 7534 30296
rect 7342 30214 7534 30240
rect 7342 30158 7347 30214
rect 7403 30158 7473 30214
rect 7529 30158 7534 30214
rect 7342 30132 7534 30158
rect 7342 30076 7347 30132
rect 7403 30076 7473 30132
rect 7529 30076 7534 30132
rect 7342 30050 7534 30076
rect 7342 29994 7347 30050
rect 7403 29994 7473 30050
rect 7529 29994 7534 30050
rect 7342 29968 7534 29994
rect 7342 29912 7347 29968
rect 7403 29912 7473 29968
rect 7529 29912 7534 29968
rect 7342 29886 7534 29912
rect 7342 29830 7347 29886
rect 7403 29830 7473 29886
rect 7529 29830 7534 29886
rect 7342 29804 7534 29830
rect 7342 29748 7347 29804
rect 7403 29748 7473 29804
rect 7529 29748 7534 29804
rect 7342 29722 7534 29748
rect 7342 29666 7347 29722
rect 7403 29666 7473 29722
rect 7529 29666 7534 29722
rect 7342 29640 7534 29666
rect 7342 29584 7347 29640
rect 7403 29584 7473 29640
rect 7529 29584 7534 29640
rect 7342 29558 7534 29584
rect 7342 29502 7347 29558
rect 7403 29502 7473 29558
rect 7529 29502 7534 29558
rect 7342 29476 7534 29502
rect 7342 29420 7347 29476
rect 7403 29420 7473 29476
rect 7529 29420 7534 29476
rect 7342 29415 7534 29420
rect 7838 34219 8030 34225
rect 7902 34155 7966 34219
rect 7838 34125 8030 34155
rect 7902 34061 7966 34125
rect 7838 34030 8030 34061
rect 7902 33966 7966 34030
rect 7838 33935 8030 33966
rect 7902 33871 7966 33935
rect 7838 33840 8030 33871
rect 7902 33776 7966 33840
rect 7838 33745 8030 33776
rect 7902 33681 7966 33745
rect 7838 32018 8030 33681
rect 7838 31962 7843 32018
rect 7899 31962 7969 32018
rect 8025 31962 8030 32018
rect 7838 31936 8030 31962
rect 7838 31880 7843 31936
rect 7899 31880 7969 31936
rect 8025 31880 8030 31936
rect 7838 31854 8030 31880
rect 7838 31798 7843 31854
rect 7899 31798 7969 31854
rect 8025 31798 8030 31854
rect 7838 31772 8030 31798
rect 7838 31716 7843 31772
rect 7899 31716 7969 31772
rect 8025 31716 8030 31772
rect 7838 31690 8030 31716
rect 7838 31634 7843 31690
rect 7899 31634 7969 31690
rect 8025 31634 8030 31690
rect 7838 31608 8030 31634
rect 7838 31552 7843 31608
rect 7899 31552 7969 31608
rect 8025 31552 8030 31608
rect 7838 31526 8030 31552
rect 7838 31470 7843 31526
rect 7899 31470 7969 31526
rect 8025 31470 8030 31526
rect 7838 31444 8030 31470
rect 7838 31388 7843 31444
rect 7899 31388 7969 31444
rect 8025 31388 8030 31444
rect 7838 31362 8030 31388
rect 7838 31306 7843 31362
rect 7899 31306 7969 31362
rect 8025 31306 8030 31362
rect 7838 31280 8030 31306
rect 7838 31224 7843 31280
rect 7899 31224 7969 31280
rect 8025 31224 8030 31280
rect 7838 31198 8030 31224
rect 7838 31142 7843 31198
rect 7899 31142 7969 31198
rect 8025 31142 8030 31198
rect 7838 31116 8030 31142
rect 7838 31060 7843 31116
rect 7899 31060 7969 31116
rect 8025 31060 8030 31116
rect 7838 31034 8030 31060
rect 7838 30978 7843 31034
rect 7899 30978 7969 31034
rect 8025 30978 8030 31034
rect 7838 30952 8030 30978
rect 7838 30896 7843 30952
rect 7899 30896 7969 30952
rect 8025 30896 8030 30952
rect 7838 30870 8030 30896
rect 7838 30814 7843 30870
rect 7899 30814 7969 30870
rect 8025 30814 8030 30870
rect 7838 30788 8030 30814
rect 7838 30732 7843 30788
rect 7899 30732 7969 30788
rect 8025 30732 8030 30788
rect 7838 30706 8030 30732
rect 7838 30650 7843 30706
rect 7899 30650 7969 30706
rect 8025 30650 8030 30706
rect 7838 30624 8030 30650
rect 7838 30568 7843 30624
rect 7899 30568 7969 30624
rect 8025 30568 8030 30624
rect 7838 30542 8030 30568
rect 7838 30486 7843 30542
rect 7899 30486 7969 30542
rect 8025 30486 8030 30542
rect 7838 30460 8030 30486
rect 7838 30404 7843 30460
rect 7899 30404 7969 30460
rect 8025 30404 8030 30460
rect 7838 30378 8030 30404
rect 7838 30322 7843 30378
rect 7899 30322 7969 30378
rect 8025 30322 8030 30378
rect 7838 30296 8030 30322
rect 7838 30240 7843 30296
rect 7899 30240 7969 30296
rect 8025 30240 8030 30296
rect 7838 30214 8030 30240
rect 7838 30158 7843 30214
rect 7899 30158 7969 30214
rect 8025 30158 8030 30214
rect 7838 30132 8030 30158
rect 7838 30076 7843 30132
rect 7899 30076 7969 30132
rect 8025 30076 8030 30132
rect 7838 30050 8030 30076
rect 7838 29994 7843 30050
rect 7899 29994 7969 30050
rect 8025 29994 8030 30050
rect 7838 29968 8030 29994
rect 7838 29912 7843 29968
rect 7899 29912 7969 29968
rect 8025 29912 8030 29968
rect 7838 29886 8030 29912
rect 7838 29830 7843 29886
rect 7899 29830 7969 29886
rect 8025 29830 8030 29886
rect 7838 29804 8030 29830
rect 7838 29748 7843 29804
rect 7899 29748 7969 29804
rect 8025 29748 8030 29804
rect 7838 29722 8030 29748
rect 7838 29666 7843 29722
rect 7899 29666 7969 29722
rect 8025 29666 8030 29722
rect 7838 29640 8030 29666
rect 7838 29584 7843 29640
rect 7899 29584 7969 29640
rect 8025 29584 8030 29640
rect 7838 29558 8030 29584
rect 7838 29502 7843 29558
rect 7899 29502 7969 29558
rect 8025 29502 8030 29558
rect 7838 29476 8030 29502
rect 7838 29420 7843 29476
rect 7899 29420 7969 29476
rect 8025 29420 8030 29476
rect 7440 28620 7538 28633
rect 7440 28564 7461 28620
rect 7517 28564 7538 28620
rect 7440 28453 7538 28564
rect 7440 28397 7461 28453
rect 7517 28397 7538 28453
rect 7440 28286 7538 28397
rect 7440 28230 7461 28286
rect 7517 28230 7538 28286
rect 7440 28119 7538 28230
rect 7440 28063 7461 28119
rect 7517 28063 7538 28119
rect 7440 27952 7538 28063
rect 7440 27896 7461 27952
rect 7517 27896 7538 27952
rect 7440 27785 7538 27896
rect 7440 27729 7461 27785
rect 7517 27729 7538 27785
rect 7440 27618 7538 27729
rect 7440 27562 7461 27618
rect 7517 27562 7538 27618
rect 7440 27451 7538 27562
rect 7440 27395 7461 27451
rect 7517 27395 7538 27451
rect 7440 27283 7538 27395
rect 7440 27227 7461 27283
rect 7517 27227 7538 27283
tri 7042 27161 7076 27195 sw
rect 6846 27137 7076 27161
tri 7076 27137 7100 27161 sw
rect 6846 27101 7100 27137
tri 7100 27101 7136 27137 sw
rect 6846 26730 7136 27101
tri 6846 26716 6860 26730 ne
rect 6860 26716 7136 26730
tri 6860 26660 6916 26716 ne
rect 6916 26660 7136 26716
tri 6916 26657 6919 26660 ne
rect 6919 26657 7136 26660
tri 6919 26632 6944 26657 ne
tri 6546 26548 6550 26552 sw
rect 6448 26492 6550 26548
tri 6550 26492 6606 26548 sw
rect 6448 26458 6606 26492
tri 6606 26458 6640 26492 sw
rect 6448 26176 6640 26458
rect 6448 26120 6453 26176
rect 6509 26120 6579 26176
rect 6635 26120 6640 26176
rect 6448 26081 6640 26120
rect 6448 26025 6453 26081
rect 6509 26025 6579 26081
rect 6635 26025 6640 26081
rect 6448 25986 6640 26025
rect 6448 25930 6453 25986
rect 6509 25930 6579 25986
rect 6635 25930 6640 25986
rect 6448 25891 6640 25930
rect 6448 25835 6453 25891
rect 6509 25835 6579 25891
rect 6635 25835 6640 25891
rect 6448 25795 6640 25835
rect 6448 25739 6453 25795
rect 6509 25739 6579 25795
rect 6635 25739 6640 25795
rect 6448 25699 6640 25739
rect 6448 25643 6453 25699
rect 6509 25643 6579 25699
rect 6635 25643 6640 25699
rect 6448 23686 6640 25643
rect 6448 23630 6457 23686
rect 6513 23630 6575 23686
rect 6631 23630 6640 23686
rect 6448 23606 6640 23630
rect 6448 23550 6457 23606
rect 6513 23550 6575 23606
rect 6631 23550 6640 23606
rect 6448 23526 6640 23550
rect 6448 23470 6457 23526
rect 6513 23470 6575 23526
rect 6631 23470 6640 23526
rect 6448 23446 6640 23470
rect 6448 23390 6457 23446
rect 6513 23390 6575 23446
rect 6631 23390 6640 23446
rect 6448 23366 6640 23390
rect 6448 23310 6457 23366
rect 6513 23310 6575 23366
rect 6631 23310 6640 23366
rect 6448 23286 6640 23310
rect 6448 23230 6457 23286
rect 6513 23230 6575 23286
rect 6631 23230 6640 23286
rect 6448 23206 6640 23230
rect 6448 23150 6457 23206
rect 6513 23150 6575 23206
rect 6631 23150 6640 23206
rect 6448 23126 6640 23150
rect 6448 23070 6457 23126
rect 6513 23070 6575 23126
rect 6631 23070 6640 23126
rect 6448 23046 6640 23070
rect 6448 22990 6457 23046
rect 6513 22990 6575 23046
rect 6631 22990 6640 23046
rect 6448 22966 6640 22990
rect 6448 22910 6457 22966
rect 6513 22910 6575 22966
rect 6631 22910 6640 22966
rect 6448 22886 6640 22910
rect 6448 22830 6457 22886
rect 6513 22830 6575 22886
rect 6631 22830 6640 22886
rect 6448 22806 6640 22830
rect 6448 22750 6457 22806
rect 6513 22750 6575 22806
rect 6631 22750 6640 22806
rect 6448 22726 6640 22750
rect 6448 22670 6457 22726
rect 6513 22670 6575 22726
rect 6631 22670 6640 22726
rect 6448 22646 6640 22670
rect 6448 22590 6457 22646
rect 6513 22590 6575 22646
rect 6631 22590 6640 22646
rect 6448 22566 6640 22590
rect 6448 22510 6457 22566
rect 6513 22510 6575 22566
rect 6631 22510 6640 22566
rect 6448 22486 6640 22510
rect 6448 22430 6457 22486
rect 6513 22430 6575 22486
rect 6631 22430 6640 22486
rect 6448 22406 6640 22430
rect 6448 22350 6457 22406
rect 6513 22350 6575 22406
rect 6631 22350 6640 22406
rect 6448 22326 6640 22350
rect 6448 22270 6457 22326
rect 6513 22270 6575 22326
rect 6631 22270 6640 22326
rect 6448 22245 6640 22270
rect 6448 22189 6457 22245
rect 6513 22189 6575 22245
rect 6631 22189 6640 22245
rect 6448 22164 6640 22189
rect 6448 22108 6457 22164
rect 6513 22108 6575 22164
rect 6631 22108 6640 22164
rect 6448 22083 6640 22108
rect 6448 22027 6457 22083
rect 6513 22027 6575 22083
rect 6631 22027 6640 22083
rect 6448 22002 6640 22027
rect 6448 21946 6457 22002
rect 6513 21946 6575 22002
rect 6631 21946 6640 22002
rect 6448 21921 6640 21946
rect 6448 21865 6457 21921
rect 6513 21865 6575 21921
rect 6631 21865 6640 21921
rect 6448 21840 6640 21865
rect 6448 21784 6457 21840
rect 6513 21784 6575 21840
rect 6631 21784 6640 21840
rect 6448 21759 6640 21784
rect 6448 21703 6457 21759
rect 6513 21703 6575 21759
rect 6631 21703 6640 21759
rect 6448 21678 6640 21703
rect 6448 21622 6457 21678
rect 6513 21622 6575 21678
rect 6631 21622 6640 21678
rect 6448 21597 6640 21622
rect 6448 21541 6457 21597
rect 6513 21541 6575 21597
rect 6631 21541 6640 21597
rect 6448 21516 6640 21541
rect 6448 21460 6457 21516
rect 6513 21460 6575 21516
rect 6631 21460 6640 21516
rect 6448 21435 6640 21460
rect 6448 21379 6457 21435
rect 6513 21379 6575 21435
rect 6631 21379 6640 21435
rect 6448 21354 6640 21379
rect 6448 21298 6457 21354
rect 6513 21298 6575 21354
rect 6631 21298 6640 21354
rect 6448 21273 6640 21298
rect 6448 21217 6457 21273
rect 6513 21217 6575 21273
rect 6631 21217 6640 21273
rect 6448 21192 6640 21217
rect 6448 21136 6457 21192
rect 6513 21136 6575 21192
rect 6631 21136 6640 21192
rect 6448 18592 6640 21136
rect 6512 18528 6576 18592
rect 6448 18512 6640 18528
rect 6512 18448 6576 18512
rect 6448 18432 6640 18448
rect 6512 18368 6576 18432
rect 6448 18352 6640 18368
rect 6512 18288 6576 18352
rect 6448 18272 6640 18288
rect 6512 18208 6576 18272
rect 6448 18192 6640 18208
rect 6512 18128 6576 18192
rect 6448 18112 6640 18128
rect 6512 18048 6576 18112
rect 6448 18032 6640 18048
rect 6512 17968 6576 18032
rect 6448 17952 6640 17968
rect 6512 17888 6576 17952
rect 6448 17872 6640 17888
rect 6512 17808 6576 17872
rect 6448 17792 6640 17808
rect 6512 17728 6576 17792
rect 6448 17712 6640 17728
rect 6512 17648 6576 17712
rect 6448 17632 6640 17648
rect 6512 17568 6576 17632
rect 6448 17552 6640 17568
rect 6512 17488 6576 17552
rect 6448 17472 6640 17488
rect 6512 17408 6576 17472
rect 6448 17392 6640 17408
rect 6512 17328 6576 17392
rect 6448 17312 6640 17328
rect 6512 17248 6576 17312
rect 6448 17232 6640 17248
rect 6512 17168 6576 17232
rect 6448 17152 6640 17168
rect 6512 17088 6576 17152
rect 6448 17072 6640 17088
rect 6512 17008 6576 17072
rect 6448 16992 6640 17008
rect 6512 16928 6576 16992
rect 6448 16912 6640 16928
rect 6512 16848 6576 16912
rect 6448 16832 6640 16848
rect 6512 16768 6576 16832
rect 6448 16752 6640 16768
rect 6512 16688 6576 16752
rect 6448 16672 6640 16688
rect 6512 16608 6576 16672
rect 6448 16592 6640 16608
rect 6512 16528 6576 16592
rect 6448 16512 6640 16528
rect 6512 16448 6576 16512
rect 6448 16432 6640 16448
rect 6512 16368 6576 16432
rect 6448 16351 6640 16368
rect 6512 16287 6576 16351
rect 6448 16270 6640 16287
rect 6512 16206 6576 16270
rect 6448 16189 6640 16206
rect 6512 16125 6576 16189
rect 6448 16108 6640 16125
rect 6512 16044 6576 16108
rect 6448 16027 6640 16044
rect 6512 15963 6576 16027
rect 6448 15946 6640 15963
rect 6512 15882 6576 15946
rect 6448 15865 6640 15882
rect 6512 15801 6576 15865
rect 6448 15784 6640 15801
rect 6512 15720 6576 15784
rect 6448 15703 6640 15720
rect 6512 15639 6576 15703
rect 6448 15622 6640 15639
rect 6512 15558 6576 15622
rect 6448 15541 6640 15558
rect 6512 15477 6576 15541
rect 6448 15460 6640 15477
rect 6512 15396 6576 15460
rect 6448 15379 6640 15396
rect 6512 15315 6576 15379
rect 6448 15298 6640 15315
rect 6512 15234 6576 15298
rect 6448 15217 6640 15234
rect 6512 15153 6576 15217
rect 6448 15136 6640 15153
rect 6512 15072 6576 15136
rect 6448 15055 6640 15072
rect 6512 14991 6576 15055
rect 6448 14974 6640 14991
rect 6512 14910 6576 14974
rect 6448 14893 6640 14910
rect 6512 14829 6576 14893
rect 6448 14812 6640 14829
rect 6512 14748 6576 14812
rect 6448 14731 6640 14748
rect 6512 14667 6576 14731
rect 6448 14650 6640 14667
rect 6512 14586 6576 14650
rect 6448 14569 6640 14586
rect 6512 14505 6576 14569
rect 6448 14488 6640 14505
rect 6512 14424 6576 14488
rect 6448 14407 6640 14424
rect 6512 14343 6576 14407
rect 6448 14326 6640 14343
rect 6512 14262 6576 14326
rect 6448 14245 6640 14262
rect 6512 14181 6576 14245
rect 6448 14164 6640 14181
rect 6512 14100 6576 14164
rect 6448 14083 6640 14100
rect 6512 14019 6576 14083
rect 6448 14002 6640 14019
rect 6512 13938 6576 14002
rect 6448 13921 6640 13938
rect 6512 13857 6576 13921
rect 6448 13840 6640 13857
rect 6512 13776 6576 13840
rect 6448 13759 6640 13776
rect 6512 13695 6576 13759
rect 6448 13678 6640 13695
rect 6512 13614 6576 13678
rect 6448 13607 6640 13614
rect 6944 23686 7136 26657
rect 6944 23630 6953 23686
rect 7009 23630 7071 23686
rect 7127 23630 7136 23686
rect 6944 23606 7136 23630
rect 6944 23550 6953 23606
rect 7009 23550 7071 23606
rect 7127 23550 7136 23606
rect 6944 23526 7136 23550
rect 6944 23470 6953 23526
rect 7009 23470 7071 23526
rect 7127 23470 7136 23526
rect 6944 23446 7136 23470
rect 6944 23390 6953 23446
rect 7009 23390 7071 23446
rect 7127 23390 7136 23446
rect 6944 23366 7136 23390
rect 6944 23310 6953 23366
rect 7009 23310 7071 23366
rect 7127 23310 7136 23366
rect 6944 23286 7136 23310
rect 6944 23230 6953 23286
rect 7009 23230 7071 23286
rect 7127 23230 7136 23286
rect 6944 23206 7136 23230
rect 6944 23150 6953 23206
rect 7009 23150 7071 23206
rect 7127 23150 7136 23206
rect 6944 23126 7136 23150
rect 6944 23070 6953 23126
rect 7009 23070 7071 23126
rect 7127 23070 7136 23126
rect 6944 23046 7136 23070
rect 6944 22990 6953 23046
rect 7009 22990 7071 23046
rect 7127 22990 7136 23046
rect 6944 22966 7136 22990
rect 6944 22910 6953 22966
rect 7009 22910 7071 22966
rect 7127 22910 7136 22966
rect 6944 22886 7136 22910
rect 6944 22830 6953 22886
rect 7009 22830 7071 22886
rect 7127 22830 7136 22886
rect 6944 22806 7136 22830
rect 6944 22750 6953 22806
rect 7009 22750 7071 22806
rect 7127 22750 7136 22806
rect 6944 22726 7136 22750
rect 6944 22670 6953 22726
rect 7009 22670 7071 22726
rect 7127 22670 7136 22726
rect 6944 22646 7136 22670
rect 6944 22590 6953 22646
rect 7009 22590 7071 22646
rect 7127 22590 7136 22646
rect 6944 22566 7136 22590
rect 6944 22510 6953 22566
rect 7009 22510 7071 22566
rect 7127 22510 7136 22566
rect 6944 22486 7136 22510
rect 6944 22430 6953 22486
rect 7009 22430 7071 22486
rect 7127 22430 7136 22486
rect 6944 22406 7136 22430
rect 6944 22350 6953 22406
rect 7009 22350 7071 22406
rect 7127 22350 7136 22406
rect 6944 22326 7136 22350
rect 6944 22270 6953 22326
rect 7009 22270 7071 22326
rect 7127 22270 7136 22326
rect 6944 22245 7136 22270
rect 6944 22189 6953 22245
rect 7009 22189 7071 22245
rect 7127 22189 7136 22245
rect 6944 22164 7136 22189
rect 6944 22108 6953 22164
rect 7009 22108 7071 22164
rect 7127 22108 7136 22164
rect 6944 22083 7136 22108
rect 6944 22027 6953 22083
rect 7009 22027 7071 22083
rect 7127 22027 7136 22083
rect 6944 22002 7136 22027
rect 6944 21946 6953 22002
rect 7009 21946 7071 22002
rect 7127 21946 7136 22002
rect 6944 21921 7136 21946
rect 6944 21865 6953 21921
rect 7009 21865 7071 21921
rect 7127 21865 7136 21921
rect 6944 21840 7136 21865
rect 6944 21784 6953 21840
rect 7009 21784 7071 21840
rect 7127 21784 7136 21840
rect 6944 21759 7136 21784
rect 6944 21703 6953 21759
rect 7009 21703 7071 21759
rect 7127 21703 7136 21759
rect 6944 21678 7136 21703
rect 6944 21622 6953 21678
rect 7009 21622 7071 21678
rect 7127 21622 7136 21678
rect 6944 21597 7136 21622
rect 6944 21541 6953 21597
rect 7009 21541 7071 21597
rect 7127 21541 7136 21597
rect 6944 21516 7136 21541
rect 6944 21460 6953 21516
rect 7009 21460 7071 21516
rect 7127 21460 7136 21516
rect 6944 21435 7136 21460
rect 6944 21379 6953 21435
rect 7009 21379 7071 21435
rect 7127 21379 7136 21435
rect 6944 21354 7136 21379
rect 6944 21298 6953 21354
rect 7009 21298 7071 21354
rect 7127 21298 7136 21354
rect 6944 21273 7136 21298
rect 6944 21217 6953 21273
rect 7009 21217 7071 21273
rect 7127 21217 7136 21273
rect 6944 21192 7136 21217
rect 6944 21136 6953 21192
rect 7009 21136 7071 21192
rect 7127 21136 7136 21192
rect 6944 19673 7136 21136
rect 6944 19609 6945 19673
rect 7009 19609 7065 19673
rect 7129 19609 7136 19673
rect 6944 19581 7136 19609
rect 6944 19517 6945 19581
rect 7009 19517 7065 19581
rect 7129 19517 7136 19581
rect 6944 19489 7136 19517
rect 6944 19425 6945 19489
rect 7009 19425 7065 19489
rect 7129 19425 7136 19489
rect 6944 19397 7136 19425
rect 6944 19333 6945 19397
rect 7009 19333 7065 19397
rect 7129 19333 7136 19397
rect 6944 19305 7136 19333
rect 6944 19241 6945 19305
rect 7009 19241 7065 19305
rect 7129 19241 7136 19305
rect 6944 19212 7136 19241
rect 6944 19148 6945 19212
rect 7009 19148 7065 19212
rect 7129 19148 7136 19212
rect 3972 13058 4160 13060
tri 2172 12887 2343 13058 sw
tri 2803 12887 2974 13058 se
rect 2974 12887 3164 13058
tri 3164 12887 3335 13058 sw
tri 3795 12887 3966 13058 se
rect 3966 12887 4160 13058
tri 4160 12887 4333 13060 sw
tri 4783 12887 4956 13060 se
rect 4956 12887 5152 13060
tri 5152 12887 5325 13060 sw
tri 5775 12887 5948 13060 se
rect 5948 12887 6144 13060
tri 6144 12887 6321 13064 sw
tri 6767 12887 6944 13064 se
rect 6944 12887 7136 19148
rect 7440 26548 7538 27227
rect 7838 27161 8030 29420
rect 8334 32018 8526 34764
rect 9326 39592 9518 39600
rect 9390 39528 9454 39592
rect 9326 39512 9518 39528
rect 9390 39448 9454 39512
rect 9326 39432 9518 39448
rect 9390 39368 9454 39432
rect 9326 39352 9518 39368
rect 9390 39288 9454 39352
rect 9326 39272 9518 39288
rect 9390 39208 9454 39272
rect 9326 39192 9518 39208
rect 9390 39128 9454 39192
rect 9326 39112 9518 39128
rect 9390 39048 9454 39112
rect 9326 39032 9518 39048
rect 9390 38968 9454 39032
rect 9326 38952 9518 38968
rect 9390 38888 9454 38952
rect 9326 38872 9518 38888
rect 9390 38808 9454 38872
rect 9326 38792 9518 38808
rect 9390 38728 9454 38792
rect 9326 38712 9518 38728
rect 9390 38648 9454 38712
rect 9326 38632 9518 38648
rect 9390 38568 9454 38632
rect 9326 38552 9518 38568
rect 9390 38488 9454 38552
rect 9326 38472 9518 38488
rect 9390 38408 9454 38472
rect 9326 38392 9518 38408
rect 9390 38328 9454 38392
rect 9326 38311 9518 38328
rect 9390 38247 9454 38311
rect 9326 38230 9518 38247
rect 9390 38166 9454 38230
rect 9326 38149 9518 38166
rect 9390 38085 9454 38149
rect 9326 38068 9518 38085
rect 9390 38004 9454 38068
rect 9326 37987 9518 38004
rect 9390 37923 9454 37987
rect 9326 37906 9518 37923
rect 9390 37842 9454 37906
rect 9326 37825 9518 37842
rect 9390 37761 9454 37825
rect 9326 37744 9518 37761
rect 9390 37680 9454 37744
rect 9326 37663 9518 37680
rect 9390 37599 9454 37663
rect 9326 37582 9518 37599
rect 9390 37518 9454 37582
rect 9326 37501 9518 37518
rect 9390 37437 9454 37501
rect 9326 37420 9518 37437
rect 9390 37356 9454 37420
rect 9326 37339 9518 37356
rect 9390 37275 9454 37339
rect 9326 37258 9518 37275
rect 9390 37194 9454 37258
rect 9326 37177 9518 37194
rect 9390 37113 9454 37177
rect 9326 37096 9518 37113
rect 9390 37032 9454 37096
rect 9326 37015 9518 37032
rect 9390 36951 9454 37015
rect 9326 36934 9518 36951
rect 9390 36870 9454 36934
rect 9326 36853 9518 36870
rect 9390 36789 9454 36853
rect 9326 36772 9518 36789
rect 9390 36708 9454 36772
rect 9326 36691 9518 36708
rect 9390 36627 9454 36691
rect 9326 36610 9518 36627
rect 9390 36546 9454 36610
rect 9326 36529 9518 36546
rect 9390 36465 9454 36529
rect 9326 36448 9518 36465
rect 9390 36384 9454 36448
rect 9326 36367 9518 36384
rect 9390 36303 9454 36367
rect 9326 36286 9518 36303
rect 9390 36222 9454 36286
rect 9326 36205 9518 36222
rect 9390 36141 9454 36205
rect 9326 36124 9518 36141
rect 9390 36060 9454 36124
rect 9326 36043 9518 36060
rect 9390 35979 9454 36043
rect 9326 35962 9518 35979
rect 9390 35898 9454 35962
rect 9326 35881 9518 35898
rect 9390 35817 9454 35881
rect 9326 35800 9518 35817
rect 9390 35736 9454 35800
rect 9326 35719 9518 35736
rect 9390 35655 9454 35719
rect 9326 35638 9518 35655
rect 9390 35574 9454 35638
rect 9326 35557 9518 35574
rect 9390 35493 9454 35557
rect 9326 35476 9518 35493
rect 9390 35412 9454 35476
rect 9326 35395 9518 35412
rect 9390 35331 9454 35395
rect 9326 35314 9518 35331
rect 9390 35250 9454 35314
rect 9326 35233 9518 35250
rect 9390 35169 9454 35233
rect 9326 35152 9518 35169
rect 9390 35088 9454 35152
rect 9326 35071 9518 35088
rect 9390 35007 9454 35071
rect 9326 34990 9518 35007
rect 9390 34926 9454 34990
rect 9326 34909 9518 34926
rect 9390 34845 9454 34909
rect 9326 34828 9518 34845
rect 9390 34764 9454 34828
rect 8334 31962 8339 32018
rect 8395 31962 8465 32018
rect 8521 31962 8526 32018
rect 8334 31936 8526 31962
rect 8334 31880 8339 31936
rect 8395 31880 8465 31936
rect 8521 31880 8526 31936
rect 8334 31854 8526 31880
rect 8334 31798 8339 31854
rect 8395 31798 8465 31854
rect 8521 31798 8526 31854
rect 8334 31772 8526 31798
rect 8334 31716 8339 31772
rect 8395 31716 8465 31772
rect 8521 31716 8526 31772
rect 8334 31690 8526 31716
rect 8334 31634 8339 31690
rect 8395 31634 8465 31690
rect 8521 31634 8526 31690
rect 8334 31608 8526 31634
rect 8334 31552 8339 31608
rect 8395 31552 8465 31608
rect 8521 31552 8526 31608
rect 8334 31526 8526 31552
rect 8334 31470 8339 31526
rect 8395 31470 8465 31526
rect 8521 31470 8526 31526
rect 8334 31444 8526 31470
rect 8334 31388 8339 31444
rect 8395 31388 8465 31444
rect 8521 31388 8526 31444
rect 8334 31362 8526 31388
rect 8334 31306 8339 31362
rect 8395 31306 8465 31362
rect 8521 31306 8526 31362
rect 8334 31280 8526 31306
rect 8334 31224 8339 31280
rect 8395 31224 8465 31280
rect 8521 31224 8526 31280
rect 8334 31198 8526 31224
rect 8334 31142 8339 31198
rect 8395 31142 8465 31198
rect 8521 31142 8526 31198
rect 8334 31116 8526 31142
rect 8334 31060 8339 31116
rect 8395 31060 8465 31116
rect 8521 31060 8526 31116
rect 8334 31034 8526 31060
rect 8334 30978 8339 31034
rect 8395 30978 8465 31034
rect 8521 30978 8526 31034
rect 8334 30952 8526 30978
rect 8334 30896 8339 30952
rect 8395 30896 8465 30952
rect 8521 30896 8526 30952
rect 8334 30870 8526 30896
rect 8334 30814 8339 30870
rect 8395 30814 8465 30870
rect 8521 30814 8526 30870
rect 8334 30788 8526 30814
rect 8334 30732 8339 30788
rect 8395 30732 8465 30788
rect 8521 30732 8526 30788
rect 8334 30706 8526 30732
rect 8334 30650 8339 30706
rect 8395 30650 8465 30706
rect 8521 30650 8526 30706
rect 8334 30624 8526 30650
rect 8334 30568 8339 30624
rect 8395 30568 8465 30624
rect 8521 30568 8526 30624
rect 8334 30542 8526 30568
rect 8334 30486 8339 30542
rect 8395 30486 8465 30542
rect 8521 30486 8526 30542
rect 8334 30460 8526 30486
rect 8334 30404 8339 30460
rect 8395 30404 8465 30460
rect 8521 30404 8526 30460
rect 8334 30378 8526 30404
rect 8334 30322 8339 30378
rect 8395 30322 8465 30378
rect 8521 30322 8526 30378
rect 8334 30296 8526 30322
rect 8334 30240 8339 30296
rect 8395 30240 8465 30296
rect 8521 30240 8526 30296
rect 8334 30214 8526 30240
rect 8334 30158 8339 30214
rect 8395 30158 8465 30214
rect 8521 30158 8526 30214
rect 8334 30132 8526 30158
rect 8334 30076 8339 30132
rect 8395 30076 8465 30132
rect 8521 30076 8526 30132
rect 8334 30050 8526 30076
rect 8334 29994 8339 30050
rect 8395 29994 8465 30050
rect 8521 29994 8526 30050
rect 8334 29968 8526 29994
rect 8334 29912 8339 29968
rect 8395 29912 8465 29968
rect 8521 29912 8526 29968
rect 8334 29886 8526 29912
rect 8334 29830 8339 29886
rect 8395 29830 8465 29886
rect 8521 29830 8526 29886
rect 8334 29804 8526 29830
rect 8334 29748 8339 29804
rect 8395 29748 8465 29804
rect 8521 29748 8526 29804
rect 8334 29722 8526 29748
rect 8334 29666 8339 29722
rect 8395 29666 8465 29722
rect 8521 29666 8526 29722
rect 8334 29640 8526 29666
rect 8334 29584 8339 29640
rect 8395 29584 8465 29640
rect 8521 29584 8526 29640
rect 8334 29558 8526 29584
rect 8334 29502 8339 29558
rect 8395 29502 8465 29558
rect 8521 29502 8526 29558
rect 8334 29476 8526 29502
rect 8334 29420 8339 29476
rect 8395 29420 8465 29476
rect 8521 29420 8526 29476
rect 8334 29415 8526 29420
rect 8830 34219 9022 34225
rect 8894 34155 8958 34219
rect 8830 34125 9022 34155
rect 8894 34061 8958 34125
rect 8830 34030 9022 34061
rect 8894 33966 8958 34030
rect 8830 33935 9022 33966
rect 8894 33871 8958 33935
rect 8830 33840 9022 33871
rect 8894 33776 8958 33840
rect 8830 33745 9022 33776
rect 8894 33681 8958 33745
rect 8830 32018 9022 33681
rect 8830 31962 8835 32018
rect 8891 31962 8961 32018
rect 9017 31962 9022 32018
rect 8830 31936 9022 31962
rect 8830 31880 8835 31936
rect 8891 31880 8961 31936
rect 9017 31880 9022 31936
rect 8830 31854 9022 31880
rect 8830 31798 8835 31854
rect 8891 31798 8961 31854
rect 9017 31798 9022 31854
rect 8830 31772 9022 31798
rect 8830 31716 8835 31772
rect 8891 31716 8961 31772
rect 9017 31716 9022 31772
rect 8830 31690 9022 31716
rect 8830 31634 8835 31690
rect 8891 31634 8961 31690
rect 9017 31634 9022 31690
rect 8830 31608 9022 31634
rect 8830 31552 8835 31608
rect 8891 31552 8961 31608
rect 9017 31552 9022 31608
rect 8830 31526 9022 31552
rect 8830 31470 8835 31526
rect 8891 31470 8961 31526
rect 9017 31470 9022 31526
rect 8830 31444 9022 31470
rect 8830 31388 8835 31444
rect 8891 31388 8961 31444
rect 9017 31388 9022 31444
rect 8830 31362 9022 31388
rect 8830 31306 8835 31362
rect 8891 31306 8961 31362
rect 9017 31306 9022 31362
rect 8830 31280 9022 31306
rect 8830 31224 8835 31280
rect 8891 31224 8961 31280
rect 9017 31224 9022 31280
rect 8830 31198 9022 31224
rect 8830 31142 8835 31198
rect 8891 31142 8961 31198
rect 9017 31142 9022 31198
rect 8830 31116 9022 31142
rect 8830 31060 8835 31116
rect 8891 31060 8961 31116
rect 9017 31060 9022 31116
rect 8830 31034 9022 31060
rect 8830 30978 8835 31034
rect 8891 30978 8961 31034
rect 9017 30978 9022 31034
rect 8830 30952 9022 30978
rect 8830 30896 8835 30952
rect 8891 30896 8961 30952
rect 9017 30896 9022 30952
rect 8830 30870 9022 30896
rect 8830 30814 8835 30870
rect 8891 30814 8961 30870
rect 9017 30814 9022 30870
rect 8830 30788 9022 30814
rect 8830 30732 8835 30788
rect 8891 30732 8961 30788
rect 9017 30732 9022 30788
rect 8830 30706 9022 30732
rect 8830 30650 8835 30706
rect 8891 30650 8961 30706
rect 9017 30650 9022 30706
rect 8830 30624 9022 30650
rect 8830 30568 8835 30624
rect 8891 30568 8961 30624
rect 9017 30568 9022 30624
rect 8830 30542 9022 30568
rect 8830 30486 8835 30542
rect 8891 30486 8961 30542
rect 9017 30486 9022 30542
rect 8830 30460 9022 30486
rect 8830 30404 8835 30460
rect 8891 30404 8961 30460
rect 9017 30404 9022 30460
rect 8830 30378 9022 30404
rect 8830 30322 8835 30378
rect 8891 30322 8961 30378
rect 9017 30322 9022 30378
rect 8830 30296 9022 30322
rect 8830 30240 8835 30296
rect 8891 30240 8961 30296
rect 9017 30240 9022 30296
rect 8830 30214 9022 30240
rect 8830 30158 8835 30214
rect 8891 30158 8961 30214
rect 9017 30158 9022 30214
rect 8830 30132 9022 30158
rect 8830 30076 8835 30132
rect 8891 30076 8961 30132
rect 9017 30076 9022 30132
rect 8830 30050 9022 30076
rect 8830 29994 8835 30050
rect 8891 29994 8961 30050
rect 9017 29994 9022 30050
rect 8830 29968 9022 29994
rect 8830 29912 8835 29968
rect 8891 29912 8961 29968
rect 9017 29912 9022 29968
rect 8830 29886 9022 29912
rect 8830 29830 8835 29886
rect 8891 29830 8961 29886
rect 9017 29830 9022 29886
rect 8830 29804 9022 29830
rect 8830 29748 8835 29804
rect 8891 29748 8961 29804
rect 9017 29748 9022 29804
rect 8830 29722 9022 29748
rect 8830 29666 8835 29722
rect 8891 29666 8961 29722
rect 9017 29666 9022 29722
rect 8830 29640 9022 29666
rect 8830 29584 8835 29640
rect 8891 29584 8961 29640
rect 9017 29584 9022 29640
rect 8830 29558 9022 29584
rect 8830 29502 8835 29558
rect 8891 29502 8961 29558
rect 9017 29502 9022 29558
rect 8830 29476 9022 29502
rect 8830 29420 8835 29476
rect 8891 29420 8961 29476
rect 9017 29420 9022 29476
rect 8432 28620 8530 28633
rect 8432 28564 8453 28620
rect 8509 28564 8530 28620
rect 8432 28453 8530 28564
rect 8432 28397 8453 28453
rect 8509 28397 8530 28453
rect 8432 28286 8530 28397
rect 8432 28230 8453 28286
rect 8509 28230 8530 28286
rect 8432 28119 8530 28230
rect 8432 28063 8453 28119
rect 8509 28063 8530 28119
rect 8432 27952 8530 28063
rect 8432 27896 8453 27952
rect 8509 27896 8530 27952
rect 8432 27785 8530 27896
rect 8432 27729 8453 27785
rect 8509 27729 8530 27785
rect 8432 27618 8530 27729
rect 8432 27562 8453 27618
rect 8509 27562 8530 27618
rect 8432 27451 8530 27562
rect 8432 27395 8453 27451
rect 8509 27395 8530 27451
rect 8432 27283 8530 27395
rect 8432 27227 8453 27283
rect 8509 27227 8530 27283
tri 8030 27161 8064 27195 sw
rect 7838 27137 8064 27161
tri 8064 27137 8088 27161 sw
rect 7838 27101 8088 27137
tri 8088 27101 8124 27137 sw
rect 7838 26726 8124 27101
tri 7838 26716 7848 26726 ne
rect 7848 26716 8124 26726
tri 7848 26660 7904 26716 ne
rect 7904 26660 8124 26716
tri 7904 26657 7907 26660 ne
rect 7907 26657 8124 26660
tri 7907 26632 7932 26657 ne
rect 7932 26632 8124 26657
tri 7932 26624 7940 26632 ne
tri 7538 26548 7542 26552 sw
rect 7440 26492 7542 26548
tri 7542 26492 7598 26548 sw
rect 7440 26458 7598 26492
tri 7598 26458 7632 26492 sw
rect 7440 26176 7632 26458
rect 7440 26120 7445 26176
rect 7501 26120 7571 26176
rect 7627 26120 7632 26176
rect 7440 26081 7632 26120
rect 7440 26025 7445 26081
rect 7501 26025 7571 26081
rect 7627 26025 7632 26081
rect 7440 25986 7632 26025
rect 7440 25930 7445 25986
rect 7501 25930 7571 25986
rect 7627 25930 7632 25986
rect 7440 25891 7632 25930
rect 7440 25835 7445 25891
rect 7501 25835 7571 25891
rect 7627 25835 7632 25891
rect 7440 25795 7632 25835
rect 7440 25739 7445 25795
rect 7501 25739 7571 25795
rect 7627 25739 7632 25795
rect 7440 25699 7632 25739
rect 7440 25643 7445 25699
rect 7501 25643 7571 25699
rect 7627 25643 7632 25699
rect 7440 23686 7632 25643
rect 7440 23630 7449 23686
rect 7505 23630 7567 23686
rect 7623 23630 7632 23686
rect 7440 23606 7632 23630
rect 7440 23550 7449 23606
rect 7505 23550 7567 23606
rect 7623 23550 7632 23606
rect 7440 23526 7632 23550
rect 7440 23470 7449 23526
rect 7505 23470 7567 23526
rect 7623 23470 7632 23526
rect 7440 23446 7632 23470
rect 7440 23390 7449 23446
rect 7505 23390 7567 23446
rect 7623 23390 7632 23446
rect 7440 23366 7632 23390
rect 7440 23310 7449 23366
rect 7505 23310 7567 23366
rect 7623 23310 7632 23366
rect 7440 23286 7632 23310
rect 7440 23230 7449 23286
rect 7505 23230 7567 23286
rect 7623 23230 7632 23286
rect 7440 23206 7632 23230
rect 7440 23150 7449 23206
rect 7505 23150 7567 23206
rect 7623 23150 7632 23206
rect 7440 23126 7632 23150
rect 7440 23070 7449 23126
rect 7505 23070 7567 23126
rect 7623 23070 7632 23126
rect 7440 23046 7632 23070
rect 7440 22990 7449 23046
rect 7505 22990 7567 23046
rect 7623 22990 7632 23046
rect 7440 22966 7632 22990
rect 7440 22910 7449 22966
rect 7505 22910 7567 22966
rect 7623 22910 7632 22966
rect 7440 22886 7632 22910
rect 7440 22830 7449 22886
rect 7505 22830 7567 22886
rect 7623 22830 7632 22886
rect 7440 22806 7632 22830
rect 7440 22750 7449 22806
rect 7505 22750 7567 22806
rect 7623 22750 7632 22806
rect 7440 22726 7632 22750
rect 7440 22670 7449 22726
rect 7505 22670 7567 22726
rect 7623 22670 7632 22726
rect 7440 22646 7632 22670
rect 7440 22590 7449 22646
rect 7505 22590 7567 22646
rect 7623 22590 7632 22646
rect 7440 22566 7632 22590
rect 7440 22510 7449 22566
rect 7505 22510 7567 22566
rect 7623 22510 7632 22566
rect 7440 22486 7632 22510
rect 7440 22430 7449 22486
rect 7505 22430 7567 22486
rect 7623 22430 7632 22486
rect 7440 22406 7632 22430
rect 7440 22350 7449 22406
rect 7505 22350 7567 22406
rect 7623 22350 7632 22406
rect 7440 22326 7632 22350
rect 7440 22270 7449 22326
rect 7505 22270 7567 22326
rect 7623 22270 7632 22326
rect 7440 22245 7632 22270
rect 7440 22189 7449 22245
rect 7505 22189 7567 22245
rect 7623 22189 7632 22245
rect 7440 22164 7632 22189
rect 7440 22108 7449 22164
rect 7505 22108 7567 22164
rect 7623 22108 7632 22164
rect 7440 22083 7632 22108
rect 7440 22027 7449 22083
rect 7505 22027 7567 22083
rect 7623 22027 7632 22083
rect 7440 22002 7632 22027
rect 7440 21946 7449 22002
rect 7505 21946 7567 22002
rect 7623 21946 7632 22002
rect 7440 21921 7632 21946
rect 7440 21865 7449 21921
rect 7505 21865 7567 21921
rect 7623 21865 7632 21921
rect 7440 21840 7632 21865
rect 7440 21784 7449 21840
rect 7505 21784 7567 21840
rect 7623 21784 7632 21840
rect 7440 21759 7632 21784
rect 7440 21703 7449 21759
rect 7505 21703 7567 21759
rect 7623 21703 7632 21759
rect 7440 21678 7632 21703
rect 7440 21622 7449 21678
rect 7505 21622 7567 21678
rect 7623 21622 7632 21678
rect 7440 21597 7632 21622
rect 7440 21541 7449 21597
rect 7505 21541 7567 21597
rect 7623 21541 7632 21597
rect 7440 21516 7632 21541
rect 7440 21460 7449 21516
rect 7505 21460 7567 21516
rect 7623 21460 7632 21516
rect 7440 21435 7632 21460
rect 7440 21379 7449 21435
rect 7505 21379 7567 21435
rect 7623 21379 7632 21435
rect 7440 21354 7632 21379
rect 7440 21298 7449 21354
rect 7505 21298 7567 21354
rect 7623 21298 7632 21354
rect 7440 21273 7632 21298
rect 7440 21217 7449 21273
rect 7505 21217 7567 21273
rect 7623 21217 7632 21273
rect 7440 21192 7632 21217
rect 7440 21136 7449 21192
rect 7505 21136 7567 21192
rect 7623 21136 7632 21192
rect 7440 18592 7632 21136
rect 7504 18528 7568 18592
rect 7440 18512 7632 18528
rect 7504 18448 7568 18512
rect 7440 18432 7632 18448
rect 7504 18368 7568 18432
rect 7440 18352 7632 18368
rect 7504 18288 7568 18352
rect 7440 18272 7632 18288
rect 7504 18208 7568 18272
rect 7440 18192 7632 18208
rect 7504 18128 7568 18192
rect 7440 18112 7632 18128
rect 7504 18048 7568 18112
rect 7440 18032 7632 18048
rect 7504 17968 7568 18032
rect 7440 17952 7632 17968
rect 7504 17888 7568 17952
rect 7440 17872 7632 17888
rect 7504 17808 7568 17872
rect 7440 17792 7632 17808
rect 7504 17728 7568 17792
rect 7440 17712 7632 17728
rect 7504 17648 7568 17712
rect 7440 17632 7632 17648
rect 7504 17568 7568 17632
rect 7440 17552 7632 17568
rect 7504 17488 7568 17552
rect 7440 17472 7632 17488
rect 7504 17408 7568 17472
rect 7440 17392 7632 17408
rect 7504 17328 7568 17392
rect 7440 17312 7632 17328
rect 7504 17248 7568 17312
rect 7440 17232 7632 17248
rect 7504 17168 7568 17232
rect 7440 17152 7632 17168
rect 7504 17088 7568 17152
rect 7440 17072 7632 17088
rect 7504 17008 7568 17072
rect 7440 16992 7632 17008
rect 7504 16928 7568 16992
rect 7440 16912 7632 16928
rect 7504 16848 7568 16912
rect 7440 16832 7632 16848
rect 7504 16768 7568 16832
rect 7440 16752 7632 16768
rect 7504 16688 7568 16752
rect 7440 16672 7632 16688
rect 7504 16608 7568 16672
rect 7440 16592 7632 16608
rect 7504 16528 7568 16592
rect 7440 16512 7632 16528
rect 7504 16448 7568 16512
rect 7440 16432 7632 16448
rect 7504 16368 7568 16432
rect 7440 16351 7632 16368
rect 7504 16287 7568 16351
rect 7440 16270 7632 16287
rect 7504 16206 7568 16270
rect 7440 16189 7632 16206
rect 7504 16125 7568 16189
rect 7440 16108 7632 16125
rect 7504 16044 7568 16108
rect 7440 16027 7632 16044
rect 7504 15963 7568 16027
rect 7440 15946 7632 15963
rect 7504 15882 7568 15946
rect 7440 15865 7632 15882
rect 7504 15801 7568 15865
rect 7440 15784 7632 15801
rect 7504 15720 7568 15784
rect 7440 15703 7632 15720
rect 7504 15639 7568 15703
rect 7440 15622 7632 15639
rect 7504 15558 7568 15622
rect 7440 15541 7632 15558
rect 7504 15477 7568 15541
rect 7440 15460 7632 15477
rect 7504 15396 7568 15460
rect 7440 15379 7632 15396
rect 7504 15315 7568 15379
rect 7440 15298 7632 15315
rect 7504 15234 7568 15298
rect 7440 15217 7632 15234
rect 7504 15153 7568 15217
rect 7440 15136 7632 15153
rect 7504 15072 7568 15136
rect 7440 15055 7632 15072
rect 7504 14991 7568 15055
rect 7440 14974 7632 14991
rect 7504 14910 7568 14974
rect 7440 14893 7632 14910
rect 7504 14829 7568 14893
rect 7440 14812 7632 14829
rect 7504 14748 7568 14812
rect 7440 14731 7632 14748
rect 7504 14667 7568 14731
rect 7440 14650 7632 14667
rect 7504 14586 7568 14650
rect 7440 14569 7632 14586
rect 7504 14505 7568 14569
rect 7440 14488 7632 14505
rect 7504 14424 7568 14488
rect 7440 14407 7632 14424
rect 7504 14343 7568 14407
rect 7440 14326 7632 14343
rect 7504 14262 7568 14326
rect 7440 14245 7632 14262
rect 7504 14181 7568 14245
rect 7440 14164 7632 14181
rect 7504 14100 7568 14164
rect 7440 14083 7632 14100
rect 7504 14019 7568 14083
rect 7440 14002 7632 14019
rect 7504 13938 7568 14002
rect 7440 13921 7632 13938
rect 7504 13857 7568 13921
rect 7440 13840 7632 13857
rect 7504 13776 7568 13840
rect 7440 13759 7632 13776
rect 7504 13695 7568 13759
rect 7440 13678 7632 13695
rect 7504 13614 7568 13678
rect 7440 13607 7632 13614
rect 7940 23686 8124 26632
rect 7940 23630 7945 23686
rect 8001 23630 8063 23686
rect 8119 23630 8124 23686
rect 7940 23606 8124 23630
rect 7940 23550 7945 23606
rect 8001 23550 8063 23606
rect 8119 23550 8124 23606
rect 7940 23526 8124 23550
rect 7940 23470 7945 23526
rect 8001 23470 8063 23526
rect 8119 23470 8124 23526
rect 7940 23446 8124 23470
rect 7940 23390 7945 23446
rect 8001 23390 8063 23446
rect 8119 23390 8124 23446
rect 7940 23366 8124 23390
rect 7940 23310 7945 23366
rect 8001 23310 8063 23366
rect 8119 23310 8124 23366
rect 7940 23286 8124 23310
rect 7940 23230 7945 23286
rect 8001 23230 8063 23286
rect 8119 23230 8124 23286
rect 7940 23206 8124 23230
rect 7940 23150 7945 23206
rect 8001 23150 8063 23206
rect 8119 23150 8124 23206
rect 7940 23126 8124 23150
rect 7940 23070 7945 23126
rect 8001 23070 8063 23126
rect 8119 23070 8124 23126
rect 7940 23046 8124 23070
rect 7940 22990 7945 23046
rect 8001 22990 8063 23046
rect 8119 22990 8124 23046
rect 7940 22966 8124 22990
rect 7940 22910 7945 22966
rect 8001 22910 8063 22966
rect 8119 22910 8124 22966
rect 7940 22886 8124 22910
rect 7940 22830 7945 22886
rect 8001 22830 8063 22886
rect 8119 22830 8124 22886
rect 7940 22806 8124 22830
rect 7940 22750 7945 22806
rect 8001 22750 8063 22806
rect 8119 22750 8124 22806
rect 7940 22726 8124 22750
rect 7940 22670 7945 22726
rect 8001 22670 8063 22726
rect 8119 22670 8124 22726
rect 7940 22646 8124 22670
rect 7940 22590 7945 22646
rect 8001 22590 8063 22646
rect 8119 22590 8124 22646
rect 7940 22566 8124 22590
rect 7940 22510 7945 22566
rect 8001 22510 8063 22566
rect 8119 22510 8124 22566
rect 7940 22486 8124 22510
rect 7940 22430 7945 22486
rect 8001 22430 8063 22486
rect 8119 22430 8124 22486
rect 7940 22406 8124 22430
rect 7940 22350 7945 22406
rect 8001 22350 8063 22406
rect 8119 22350 8124 22406
rect 7940 22326 8124 22350
rect 7940 22270 7945 22326
rect 8001 22270 8063 22326
rect 8119 22270 8124 22326
rect 7940 22245 8124 22270
rect 7940 22189 7945 22245
rect 8001 22189 8063 22245
rect 8119 22189 8124 22245
rect 7940 22164 8124 22189
rect 7940 22108 7945 22164
rect 8001 22108 8063 22164
rect 8119 22108 8124 22164
rect 7940 22083 8124 22108
rect 7940 22027 7945 22083
rect 8001 22027 8063 22083
rect 8119 22027 8124 22083
rect 7940 22002 8124 22027
rect 7940 21946 7945 22002
rect 8001 21946 8063 22002
rect 8119 21946 8124 22002
rect 7940 21921 8124 21946
rect 7940 21865 7945 21921
rect 8001 21865 8063 21921
rect 8119 21865 8124 21921
rect 7940 21840 8124 21865
rect 7940 21784 7945 21840
rect 8001 21784 8063 21840
rect 8119 21784 8124 21840
rect 7940 21759 8124 21784
rect 7940 21703 7945 21759
rect 8001 21703 8063 21759
rect 8119 21703 8124 21759
rect 7940 21678 8124 21703
rect 7940 21622 7945 21678
rect 8001 21622 8063 21678
rect 8119 21622 8124 21678
rect 7940 21597 8124 21622
rect 7940 21541 7945 21597
rect 8001 21541 8063 21597
rect 8119 21541 8124 21597
rect 7940 21516 8124 21541
rect 7940 21460 7945 21516
rect 8001 21460 8063 21516
rect 8119 21460 8124 21516
rect 7940 21435 8124 21460
rect 7940 21379 7945 21435
rect 8001 21379 8063 21435
rect 8119 21379 8124 21435
rect 7940 21354 8124 21379
rect 7940 21298 7945 21354
rect 8001 21298 8063 21354
rect 8119 21298 8124 21354
rect 7940 21273 8124 21298
rect 7940 21217 7945 21273
rect 8001 21217 8063 21273
rect 8119 21217 8124 21273
rect 7940 21192 8124 21217
rect 7940 21136 7945 21192
rect 8001 21136 8063 21192
rect 8119 21136 8124 21192
rect 7940 19673 8124 21136
rect 8004 19609 8060 19673
rect 7940 19581 8124 19609
rect 8004 19517 8060 19581
rect 7940 19489 8124 19517
rect 8004 19425 8060 19489
rect 7940 19397 8124 19425
rect 8004 19333 8060 19397
rect 7940 19305 8124 19333
rect 8004 19241 8060 19305
rect 7940 19212 8124 19241
rect 8004 19148 8060 19212
tri 7136 12887 7313 13064 sw
tri 7763 12887 7940 13064 se
rect 7940 12887 8124 19148
rect 8432 26548 8530 27227
rect 8830 27161 9022 29420
rect 9326 32018 9518 34764
rect 10318 39592 10510 39600
rect 10382 39528 10446 39592
rect 10318 39512 10510 39528
rect 10382 39448 10446 39512
rect 10318 39432 10510 39448
rect 10382 39368 10446 39432
rect 10318 39352 10510 39368
rect 10382 39288 10446 39352
rect 10318 39272 10510 39288
rect 10382 39208 10446 39272
rect 10318 39192 10510 39208
rect 10382 39128 10446 39192
rect 10318 39112 10510 39128
rect 10382 39048 10446 39112
rect 10318 39032 10510 39048
rect 10382 38968 10446 39032
rect 10318 38952 10510 38968
rect 10382 38888 10446 38952
rect 10318 38872 10510 38888
rect 10382 38808 10446 38872
rect 10318 38792 10510 38808
rect 10382 38728 10446 38792
rect 10318 38712 10510 38728
rect 10382 38648 10446 38712
rect 10318 38632 10510 38648
rect 10382 38568 10446 38632
rect 10318 38552 10510 38568
rect 10382 38488 10446 38552
rect 10318 38472 10510 38488
rect 10382 38408 10446 38472
rect 10318 38392 10510 38408
rect 10382 38328 10446 38392
rect 10318 38311 10510 38328
rect 10382 38247 10446 38311
rect 10318 38230 10510 38247
rect 10382 38166 10446 38230
rect 10318 38149 10510 38166
rect 10382 38085 10446 38149
rect 10318 38068 10510 38085
rect 10382 38004 10446 38068
rect 10318 37987 10510 38004
rect 10382 37923 10446 37987
rect 10318 37906 10510 37923
rect 10382 37842 10446 37906
rect 10318 37825 10510 37842
rect 10382 37761 10446 37825
rect 10318 37744 10510 37761
rect 10382 37680 10446 37744
rect 10318 37663 10510 37680
rect 10382 37599 10446 37663
rect 10318 37582 10510 37599
rect 10382 37518 10446 37582
rect 10318 37501 10510 37518
rect 10382 37437 10446 37501
rect 10318 37420 10510 37437
rect 10382 37356 10446 37420
rect 10318 37339 10510 37356
rect 10382 37275 10446 37339
rect 10318 37258 10510 37275
rect 10382 37194 10446 37258
rect 10318 37177 10510 37194
rect 10382 37113 10446 37177
rect 10318 37096 10510 37113
rect 10382 37032 10446 37096
rect 10318 37015 10510 37032
rect 10382 36951 10446 37015
rect 10318 36934 10510 36951
rect 10382 36870 10446 36934
rect 10318 36853 10510 36870
rect 10382 36789 10446 36853
rect 10318 36772 10510 36789
rect 10382 36708 10446 36772
rect 10318 36691 10510 36708
rect 10382 36627 10446 36691
rect 10318 36610 10510 36627
rect 10382 36546 10446 36610
rect 10318 36529 10510 36546
rect 10382 36465 10446 36529
rect 10318 36448 10510 36465
rect 10382 36384 10446 36448
rect 10318 36367 10510 36384
rect 10382 36303 10446 36367
rect 10318 36286 10510 36303
rect 10382 36222 10446 36286
rect 10318 36205 10510 36222
rect 10382 36141 10446 36205
rect 10318 36124 10510 36141
rect 10382 36060 10446 36124
rect 10318 36043 10510 36060
rect 10382 35979 10446 36043
rect 10318 35962 10510 35979
rect 10382 35898 10446 35962
rect 10318 35881 10510 35898
rect 10382 35817 10446 35881
rect 10318 35800 10510 35817
rect 10382 35736 10446 35800
rect 10318 35719 10510 35736
rect 10382 35655 10446 35719
rect 10318 35638 10510 35655
rect 10382 35574 10446 35638
rect 10318 35557 10510 35574
rect 10382 35493 10446 35557
rect 10318 35476 10510 35493
rect 10382 35412 10446 35476
rect 10318 35395 10510 35412
rect 10382 35331 10446 35395
rect 10318 35314 10510 35331
rect 10382 35250 10446 35314
rect 10318 35233 10510 35250
rect 10382 35169 10446 35233
rect 10318 35152 10510 35169
rect 10382 35088 10446 35152
rect 10318 35071 10510 35088
rect 10382 35007 10446 35071
rect 10318 34990 10510 35007
rect 10382 34926 10446 34990
rect 10318 34909 10510 34926
rect 10382 34845 10446 34909
rect 10318 34828 10510 34845
rect 10382 34764 10446 34828
rect 9326 31962 9331 32018
rect 9387 31962 9457 32018
rect 9513 31962 9518 32018
rect 9326 31936 9518 31962
rect 9326 31880 9331 31936
rect 9387 31880 9457 31936
rect 9513 31880 9518 31936
rect 9326 31854 9518 31880
rect 9326 31798 9331 31854
rect 9387 31798 9457 31854
rect 9513 31798 9518 31854
rect 9326 31772 9518 31798
rect 9326 31716 9331 31772
rect 9387 31716 9457 31772
rect 9513 31716 9518 31772
rect 9326 31690 9518 31716
rect 9326 31634 9331 31690
rect 9387 31634 9457 31690
rect 9513 31634 9518 31690
rect 9326 31608 9518 31634
rect 9326 31552 9331 31608
rect 9387 31552 9457 31608
rect 9513 31552 9518 31608
rect 9326 31526 9518 31552
rect 9326 31470 9331 31526
rect 9387 31470 9457 31526
rect 9513 31470 9518 31526
rect 9326 31444 9518 31470
rect 9326 31388 9331 31444
rect 9387 31388 9457 31444
rect 9513 31388 9518 31444
rect 9326 31362 9518 31388
rect 9326 31306 9331 31362
rect 9387 31306 9457 31362
rect 9513 31306 9518 31362
rect 9326 31280 9518 31306
rect 9326 31224 9331 31280
rect 9387 31224 9457 31280
rect 9513 31224 9518 31280
rect 9326 31198 9518 31224
rect 9326 31142 9331 31198
rect 9387 31142 9457 31198
rect 9513 31142 9518 31198
rect 9326 31116 9518 31142
rect 9326 31060 9331 31116
rect 9387 31060 9457 31116
rect 9513 31060 9518 31116
rect 9326 31034 9518 31060
rect 9326 30978 9331 31034
rect 9387 30978 9457 31034
rect 9513 30978 9518 31034
rect 9326 30952 9518 30978
rect 9326 30896 9331 30952
rect 9387 30896 9457 30952
rect 9513 30896 9518 30952
rect 9326 30870 9518 30896
rect 9326 30814 9331 30870
rect 9387 30814 9457 30870
rect 9513 30814 9518 30870
rect 9326 30788 9518 30814
rect 9326 30732 9331 30788
rect 9387 30732 9457 30788
rect 9513 30732 9518 30788
rect 9326 30706 9518 30732
rect 9326 30650 9331 30706
rect 9387 30650 9457 30706
rect 9513 30650 9518 30706
rect 9326 30624 9518 30650
rect 9326 30568 9331 30624
rect 9387 30568 9457 30624
rect 9513 30568 9518 30624
rect 9326 30542 9518 30568
rect 9326 30486 9331 30542
rect 9387 30486 9457 30542
rect 9513 30486 9518 30542
rect 9326 30460 9518 30486
rect 9326 30404 9331 30460
rect 9387 30404 9457 30460
rect 9513 30404 9518 30460
rect 9326 30378 9518 30404
rect 9326 30322 9331 30378
rect 9387 30322 9457 30378
rect 9513 30322 9518 30378
rect 9326 30296 9518 30322
rect 9326 30240 9331 30296
rect 9387 30240 9457 30296
rect 9513 30240 9518 30296
rect 9326 30214 9518 30240
rect 9326 30158 9331 30214
rect 9387 30158 9457 30214
rect 9513 30158 9518 30214
rect 9326 30132 9518 30158
rect 9326 30076 9331 30132
rect 9387 30076 9457 30132
rect 9513 30076 9518 30132
rect 9326 30050 9518 30076
rect 9326 29994 9331 30050
rect 9387 29994 9457 30050
rect 9513 29994 9518 30050
rect 9326 29968 9518 29994
rect 9326 29912 9331 29968
rect 9387 29912 9457 29968
rect 9513 29912 9518 29968
rect 9326 29886 9518 29912
rect 9326 29830 9331 29886
rect 9387 29830 9457 29886
rect 9513 29830 9518 29886
rect 9326 29804 9518 29830
rect 9326 29748 9331 29804
rect 9387 29748 9457 29804
rect 9513 29748 9518 29804
rect 9326 29722 9518 29748
rect 9326 29666 9331 29722
rect 9387 29666 9457 29722
rect 9513 29666 9518 29722
rect 9326 29640 9518 29666
rect 9326 29584 9331 29640
rect 9387 29584 9457 29640
rect 9513 29584 9518 29640
rect 9326 29558 9518 29584
rect 9326 29502 9331 29558
rect 9387 29502 9457 29558
rect 9513 29502 9518 29558
rect 9326 29476 9518 29502
rect 9326 29420 9331 29476
rect 9387 29420 9457 29476
rect 9513 29420 9518 29476
rect 9326 29415 9518 29420
rect 9822 34219 10014 34225
rect 9886 34155 9950 34219
rect 9822 34125 10014 34155
rect 9886 34061 9950 34125
rect 9822 34030 10014 34061
rect 9886 33966 9950 34030
rect 9822 33935 10014 33966
rect 9886 33871 9950 33935
rect 9822 33840 10014 33871
rect 9886 33776 9950 33840
rect 9822 33745 10014 33776
rect 9886 33681 9950 33745
rect 9822 32018 10014 33681
rect 9822 31962 9827 32018
rect 9883 31962 9953 32018
rect 10009 31962 10014 32018
rect 9822 31936 10014 31962
rect 9822 31880 9827 31936
rect 9883 31880 9953 31936
rect 10009 31880 10014 31936
rect 9822 31854 10014 31880
rect 9822 31798 9827 31854
rect 9883 31798 9953 31854
rect 10009 31798 10014 31854
rect 9822 31772 10014 31798
rect 9822 31716 9827 31772
rect 9883 31716 9953 31772
rect 10009 31716 10014 31772
rect 9822 31690 10014 31716
rect 9822 31634 9827 31690
rect 9883 31634 9953 31690
rect 10009 31634 10014 31690
rect 9822 31608 10014 31634
rect 9822 31552 9827 31608
rect 9883 31552 9953 31608
rect 10009 31552 10014 31608
rect 9822 31526 10014 31552
rect 9822 31470 9827 31526
rect 9883 31470 9953 31526
rect 10009 31470 10014 31526
rect 9822 31444 10014 31470
rect 9822 31388 9827 31444
rect 9883 31388 9953 31444
rect 10009 31388 10014 31444
rect 9822 31362 10014 31388
rect 9822 31306 9827 31362
rect 9883 31306 9953 31362
rect 10009 31306 10014 31362
rect 9822 31280 10014 31306
rect 9822 31224 9827 31280
rect 9883 31224 9953 31280
rect 10009 31224 10014 31280
rect 9822 31198 10014 31224
rect 9822 31142 9827 31198
rect 9883 31142 9953 31198
rect 10009 31142 10014 31198
rect 9822 31116 10014 31142
rect 9822 31060 9827 31116
rect 9883 31060 9953 31116
rect 10009 31060 10014 31116
rect 9822 31034 10014 31060
rect 9822 30978 9827 31034
rect 9883 30978 9953 31034
rect 10009 30978 10014 31034
rect 9822 30952 10014 30978
rect 9822 30896 9827 30952
rect 9883 30896 9953 30952
rect 10009 30896 10014 30952
rect 9822 30870 10014 30896
rect 9822 30814 9827 30870
rect 9883 30814 9953 30870
rect 10009 30814 10014 30870
rect 9822 30788 10014 30814
rect 9822 30732 9827 30788
rect 9883 30732 9953 30788
rect 10009 30732 10014 30788
rect 9822 30706 10014 30732
rect 9822 30650 9827 30706
rect 9883 30650 9953 30706
rect 10009 30650 10014 30706
rect 9822 30624 10014 30650
rect 9822 30568 9827 30624
rect 9883 30568 9953 30624
rect 10009 30568 10014 30624
rect 9822 30542 10014 30568
rect 9822 30486 9827 30542
rect 9883 30486 9953 30542
rect 10009 30486 10014 30542
rect 9822 30460 10014 30486
rect 9822 30404 9827 30460
rect 9883 30404 9953 30460
rect 10009 30404 10014 30460
rect 9822 30378 10014 30404
rect 9822 30322 9827 30378
rect 9883 30322 9953 30378
rect 10009 30322 10014 30378
rect 9822 30296 10014 30322
rect 9822 30240 9827 30296
rect 9883 30240 9953 30296
rect 10009 30240 10014 30296
rect 9822 30214 10014 30240
rect 9822 30158 9827 30214
rect 9883 30158 9953 30214
rect 10009 30158 10014 30214
rect 9822 30132 10014 30158
rect 9822 30076 9827 30132
rect 9883 30076 9953 30132
rect 10009 30076 10014 30132
rect 9822 30050 10014 30076
rect 9822 29994 9827 30050
rect 9883 29994 9953 30050
rect 10009 29994 10014 30050
rect 9822 29968 10014 29994
rect 9822 29912 9827 29968
rect 9883 29912 9953 29968
rect 10009 29912 10014 29968
rect 9822 29886 10014 29912
rect 9822 29830 9827 29886
rect 9883 29830 9953 29886
rect 10009 29830 10014 29886
rect 9822 29804 10014 29830
rect 9822 29748 9827 29804
rect 9883 29748 9953 29804
rect 10009 29748 10014 29804
rect 9822 29722 10014 29748
rect 9822 29666 9827 29722
rect 9883 29666 9953 29722
rect 10009 29666 10014 29722
rect 9822 29640 10014 29666
rect 9822 29584 9827 29640
rect 9883 29584 9953 29640
rect 10009 29584 10014 29640
rect 9822 29558 10014 29584
rect 9822 29502 9827 29558
rect 9883 29502 9953 29558
rect 10009 29502 10014 29558
rect 9822 29476 10014 29502
rect 9822 29420 9827 29476
rect 9883 29420 9953 29476
rect 10009 29420 10014 29476
rect 9424 28620 9522 28633
rect 9424 28564 9445 28620
rect 9501 28564 9522 28620
rect 9424 28453 9522 28564
rect 9424 28397 9445 28453
rect 9501 28397 9522 28453
rect 9424 28286 9522 28397
rect 9424 28230 9445 28286
rect 9501 28230 9522 28286
rect 9424 28119 9522 28230
rect 9424 28063 9445 28119
rect 9501 28063 9522 28119
rect 9424 27952 9522 28063
rect 9424 27896 9445 27952
rect 9501 27896 9522 27952
rect 9424 27785 9522 27896
rect 9424 27729 9445 27785
rect 9501 27729 9522 27785
rect 9424 27618 9522 27729
rect 9424 27562 9445 27618
rect 9501 27562 9522 27618
rect 9424 27451 9522 27562
rect 9424 27395 9445 27451
rect 9501 27395 9522 27451
rect 9424 27283 9522 27395
rect 9424 27227 9445 27283
rect 9501 27227 9522 27283
tri 9022 27161 9056 27195 sw
rect 8830 27137 9056 27161
tri 9056 27137 9080 27161 sw
rect 8830 27101 9080 27137
tri 9080 27101 9116 27137 sw
rect 8830 26726 9116 27101
tri 8830 26716 8840 26726 ne
rect 8840 26716 9116 26726
tri 8840 26660 8896 26716 ne
rect 8896 26660 9116 26716
tri 8896 26657 8899 26660 ne
rect 8899 26657 9116 26660
tri 8899 26632 8924 26657 ne
rect 8924 26632 9116 26657
tri 8924 26624 8932 26632 ne
tri 8530 26548 8534 26552 sw
rect 8432 26492 8534 26548
tri 8534 26492 8590 26548 sw
rect 8432 26458 8590 26492
tri 8590 26458 8624 26492 sw
rect 8432 26176 8624 26458
rect 8432 26120 8437 26176
rect 8493 26120 8563 26176
rect 8619 26120 8624 26176
rect 8432 26081 8624 26120
rect 8432 26025 8437 26081
rect 8493 26025 8563 26081
rect 8619 26025 8624 26081
rect 8432 25986 8624 26025
rect 8432 25930 8437 25986
rect 8493 25930 8563 25986
rect 8619 25930 8624 25986
rect 8432 25891 8624 25930
rect 8432 25835 8437 25891
rect 8493 25835 8563 25891
rect 8619 25835 8624 25891
rect 8432 25795 8624 25835
rect 8432 25739 8437 25795
rect 8493 25739 8563 25795
rect 8619 25739 8624 25795
rect 8432 25699 8624 25739
rect 8432 25643 8437 25699
rect 8493 25643 8563 25699
rect 8619 25643 8624 25699
rect 8432 23686 8624 25643
rect 8432 23630 8441 23686
rect 8497 23630 8559 23686
rect 8615 23630 8624 23686
rect 8432 23606 8624 23630
rect 8432 23550 8441 23606
rect 8497 23550 8559 23606
rect 8615 23550 8624 23606
rect 8432 23526 8624 23550
rect 8432 23470 8441 23526
rect 8497 23470 8559 23526
rect 8615 23470 8624 23526
rect 8432 23446 8624 23470
rect 8432 23390 8441 23446
rect 8497 23390 8559 23446
rect 8615 23390 8624 23446
rect 8432 23366 8624 23390
rect 8432 23310 8441 23366
rect 8497 23310 8559 23366
rect 8615 23310 8624 23366
rect 8432 23286 8624 23310
rect 8432 23230 8441 23286
rect 8497 23230 8559 23286
rect 8615 23230 8624 23286
rect 8432 23206 8624 23230
rect 8432 23150 8441 23206
rect 8497 23150 8559 23206
rect 8615 23150 8624 23206
rect 8432 23126 8624 23150
rect 8432 23070 8441 23126
rect 8497 23070 8559 23126
rect 8615 23070 8624 23126
rect 8432 23046 8624 23070
rect 8432 22990 8441 23046
rect 8497 22990 8559 23046
rect 8615 22990 8624 23046
rect 8432 22966 8624 22990
rect 8432 22910 8441 22966
rect 8497 22910 8559 22966
rect 8615 22910 8624 22966
rect 8432 22886 8624 22910
rect 8432 22830 8441 22886
rect 8497 22830 8559 22886
rect 8615 22830 8624 22886
rect 8432 22806 8624 22830
rect 8432 22750 8441 22806
rect 8497 22750 8559 22806
rect 8615 22750 8624 22806
rect 8432 22726 8624 22750
rect 8432 22670 8441 22726
rect 8497 22670 8559 22726
rect 8615 22670 8624 22726
rect 8432 22646 8624 22670
rect 8432 22590 8441 22646
rect 8497 22590 8559 22646
rect 8615 22590 8624 22646
rect 8432 22566 8624 22590
rect 8432 22510 8441 22566
rect 8497 22510 8559 22566
rect 8615 22510 8624 22566
rect 8432 22486 8624 22510
rect 8432 22430 8441 22486
rect 8497 22430 8559 22486
rect 8615 22430 8624 22486
rect 8432 22406 8624 22430
rect 8432 22350 8441 22406
rect 8497 22350 8559 22406
rect 8615 22350 8624 22406
rect 8432 22326 8624 22350
rect 8432 22270 8441 22326
rect 8497 22270 8559 22326
rect 8615 22270 8624 22326
rect 8432 22245 8624 22270
rect 8432 22189 8441 22245
rect 8497 22189 8559 22245
rect 8615 22189 8624 22245
rect 8432 22164 8624 22189
rect 8432 22108 8441 22164
rect 8497 22108 8559 22164
rect 8615 22108 8624 22164
rect 8432 22083 8624 22108
rect 8432 22027 8441 22083
rect 8497 22027 8559 22083
rect 8615 22027 8624 22083
rect 8432 22002 8624 22027
rect 8432 21946 8441 22002
rect 8497 21946 8559 22002
rect 8615 21946 8624 22002
rect 8432 21921 8624 21946
rect 8432 21865 8441 21921
rect 8497 21865 8559 21921
rect 8615 21865 8624 21921
rect 8432 21840 8624 21865
rect 8432 21784 8441 21840
rect 8497 21784 8559 21840
rect 8615 21784 8624 21840
rect 8432 21759 8624 21784
rect 8432 21703 8441 21759
rect 8497 21703 8559 21759
rect 8615 21703 8624 21759
rect 8432 21678 8624 21703
rect 8432 21622 8441 21678
rect 8497 21622 8559 21678
rect 8615 21622 8624 21678
rect 8432 21597 8624 21622
rect 8432 21541 8441 21597
rect 8497 21541 8559 21597
rect 8615 21541 8624 21597
rect 8432 21516 8624 21541
rect 8432 21460 8441 21516
rect 8497 21460 8559 21516
rect 8615 21460 8624 21516
rect 8432 21435 8624 21460
rect 8432 21379 8441 21435
rect 8497 21379 8559 21435
rect 8615 21379 8624 21435
rect 8432 21354 8624 21379
rect 8432 21298 8441 21354
rect 8497 21298 8559 21354
rect 8615 21298 8624 21354
rect 8432 21273 8624 21298
rect 8432 21217 8441 21273
rect 8497 21217 8559 21273
rect 8615 21217 8624 21273
rect 8432 21192 8624 21217
rect 8432 21136 8441 21192
rect 8497 21136 8559 21192
rect 8615 21136 8624 21192
rect 8432 18592 8624 21136
rect 8932 23686 9116 26632
rect 8932 23630 8937 23686
rect 8993 23630 9055 23686
rect 9111 23630 9116 23686
rect 8932 23606 9116 23630
rect 8932 23550 8937 23606
rect 8993 23550 9055 23606
rect 9111 23550 9116 23606
rect 8932 23526 9116 23550
rect 8932 23470 8937 23526
rect 8993 23470 9055 23526
rect 9111 23470 9116 23526
rect 8932 23446 9116 23470
rect 8932 23390 8937 23446
rect 8993 23390 9055 23446
rect 9111 23390 9116 23446
rect 8932 23366 9116 23390
rect 8932 23310 8937 23366
rect 8993 23310 9055 23366
rect 9111 23310 9116 23366
rect 8932 23286 9116 23310
rect 8932 23230 8937 23286
rect 8993 23230 9055 23286
rect 9111 23230 9116 23286
rect 8932 23206 9116 23230
rect 8932 23150 8937 23206
rect 8993 23150 9055 23206
rect 9111 23150 9116 23206
rect 8932 23126 9116 23150
rect 8932 23070 8937 23126
rect 8993 23070 9055 23126
rect 9111 23070 9116 23126
rect 8932 23046 9116 23070
rect 8932 22990 8937 23046
rect 8993 22990 9055 23046
rect 9111 22990 9116 23046
rect 8932 22966 9116 22990
rect 8932 22910 8937 22966
rect 8993 22910 9055 22966
rect 9111 22910 9116 22966
rect 8932 22886 9116 22910
rect 8932 22830 8937 22886
rect 8993 22830 9055 22886
rect 9111 22830 9116 22886
rect 8932 22806 9116 22830
rect 8932 22750 8937 22806
rect 8993 22750 9055 22806
rect 9111 22750 9116 22806
rect 8932 22726 9116 22750
rect 8932 22670 8937 22726
rect 8993 22670 9055 22726
rect 9111 22670 9116 22726
rect 8932 22646 9116 22670
rect 8932 22590 8937 22646
rect 8993 22590 9055 22646
rect 9111 22590 9116 22646
rect 8932 22566 9116 22590
rect 8932 22510 8937 22566
rect 8993 22510 9055 22566
rect 9111 22510 9116 22566
rect 8932 22486 9116 22510
rect 8932 22430 8937 22486
rect 8993 22430 9055 22486
rect 9111 22430 9116 22486
rect 8932 22406 9116 22430
rect 8932 22350 8937 22406
rect 8993 22350 9055 22406
rect 9111 22350 9116 22406
rect 8932 22326 9116 22350
rect 8932 22270 8937 22326
rect 8993 22270 9055 22326
rect 9111 22270 9116 22326
rect 8932 22245 9116 22270
rect 8932 22189 8937 22245
rect 8993 22189 9055 22245
rect 9111 22189 9116 22245
rect 8932 22164 9116 22189
rect 8932 22108 8937 22164
rect 8993 22108 9055 22164
rect 9111 22108 9116 22164
rect 8932 22083 9116 22108
rect 8932 22027 8937 22083
rect 8993 22027 9055 22083
rect 9111 22027 9116 22083
rect 8932 22002 9116 22027
rect 8932 21946 8937 22002
rect 8993 21946 9055 22002
rect 9111 21946 9116 22002
rect 8932 21921 9116 21946
rect 8932 21865 8937 21921
rect 8993 21865 9055 21921
rect 9111 21865 9116 21921
rect 8932 21840 9116 21865
rect 8932 21784 8937 21840
rect 8993 21784 9055 21840
rect 9111 21784 9116 21840
rect 8932 21759 9116 21784
rect 8932 21703 8937 21759
rect 8993 21703 9055 21759
rect 9111 21703 9116 21759
rect 8932 21678 9116 21703
rect 8932 21622 8937 21678
rect 8993 21622 9055 21678
rect 9111 21622 9116 21678
rect 8932 21597 9116 21622
rect 8932 21541 8937 21597
rect 8993 21541 9055 21597
rect 9111 21541 9116 21597
rect 8932 21516 9116 21541
rect 8932 21460 8937 21516
rect 8993 21460 9055 21516
rect 9111 21460 9116 21516
rect 8932 21435 9116 21460
rect 8932 21379 8937 21435
rect 8993 21379 9055 21435
rect 9111 21379 9116 21435
rect 8932 21354 9116 21379
rect 8932 21298 8937 21354
rect 8993 21298 9055 21354
rect 9111 21298 9116 21354
rect 8932 21273 9116 21298
rect 8932 21217 8937 21273
rect 8993 21217 9055 21273
rect 9111 21217 9116 21273
rect 8932 21192 9116 21217
rect 8932 21136 8937 21192
rect 8993 21136 9055 21192
rect 9111 21136 9116 21192
rect 8932 19673 9116 21136
rect 8996 19609 9052 19673
rect 8932 19581 9116 19609
rect 8996 19517 9052 19581
rect 8932 19489 9116 19517
rect 8996 19425 9052 19489
rect 8932 19397 9116 19425
rect 8996 19333 9052 19397
rect 8932 19305 9116 19333
rect 8996 19241 9052 19305
rect 8932 19212 9116 19241
rect 8996 19148 9052 19212
rect 8932 19139 9116 19148
rect 9424 26548 9522 27227
rect 9822 27161 10014 29420
rect 10318 32018 10510 34764
rect 11310 39592 11502 39600
rect 11374 39528 11438 39592
rect 11310 39512 11502 39528
rect 11374 39448 11438 39512
rect 11310 39432 11502 39448
rect 11374 39368 11438 39432
rect 11310 39352 11502 39368
rect 11374 39288 11438 39352
rect 11310 39272 11502 39288
rect 11374 39208 11438 39272
rect 11310 39192 11502 39208
rect 11374 39128 11438 39192
rect 11310 39112 11502 39128
rect 11374 39048 11438 39112
rect 11310 39032 11502 39048
rect 11374 38968 11438 39032
rect 11310 38952 11502 38968
rect 11374 38888 11438 38952
rect 11310 38872 11502 38888
rect 11374 38808 11438 38872
rect 11310 38792 11502 38808
rect 11374 38728 11438 38792
rect 11310 38712 11502 38728
rect 11374 38648 11438 38712
rect 11310 38632 11502 38648
rect 11374 38568 11438 38632
rect 11310 38552 11502 38568
rect 11374 38488 11438 38552
rect 11310 38472 11502 38488
rect 11374 38408 11438 38472
rect 11310 38392 11502 38408
rect 11374 38328 11438 38392
rect 11310 38311 11502 38328
rect 11374 38247 11438 38311
rect 11310 38230 11502 38247
rect 11374 38166 11438 38230
rect 11310 38149 11502 38166
rect 11374 38085 11438 38149
rect 11310 38068 11502 38085
rect 11374 38004 11438 38068
rect 11310 37987 11502 38004
rect 11374 37923 11438 37987
rect 11310 37906 11502 37923
rect 11374 37842 11438 37906
rect 11310 37825 11502 37842
rect 11374 37761 11438 37825
rect 11310 37744 11502 37761
rect 11374 37680 11438 37744
rect 11310 37663 11502 37680
rect 11374 37599 11438 37663
rect 11310 37582 11502 37599
rect 11374 37518 11438 37582
rect 11310 37501 11502 37518
rect 11374 37437 11438 37501
rect 11310 37420 11502 37437
rect 11374 37356 11438 37420
rect 11310 37339 11502 37356
rect 11374 37275 11438 37339
rect 11310 37258 11502 37275
rect 11374 37194 11438 37258
rect 11310 37177 11502 37194
rect 11374 37113 11438 37177
rect 11310 37096 11502 37113
rect 11374 37032 11438 37096
rect 11310 37015 11502 37032
rect 11374 36951 11438 37015
rect 11310 36934 11502 36951
rect 11374 36870 11438 36934
rect 11310 36853 11502 36870
rect 11374 36789 11438 36853
rect 11310 36772 11502 36789
rect 11374 36708 11438 36772
rect 11310 36691 11502 36708
rect 11374 36627 11438 36691
rect 11310 36610 11502 36627
rect 11374 36546 11438 36610
rect 11310 36529 11502 36546
rect 11374 36465 11438 36529
rect 11310 36448 11502 36465
rect 11374 36384 11438 36448
rect 11310 36367 11502 36384
rect 11374 36303 11438 36367
rect 11310 36286 11502 36303
rect 11374 36222 11438 36286
rect 11310 36205 11502 36222
rect 11374 36141 11438 36205
rect 11310 36124 11502 36141
rect 11374 36060 11438 36124
rect 11310 36043 11502 36060
rect 11374 35979 11438 36043
rect 11310 35962 11502 35979
rect 11374 35898 11438 35962
rect 11310 35881 11502 35898
rect 11374 35817 11438 35881
rect 11310 35800 11502 35817
rect 11374 35736 11438 35800
rect 11310 35719 11502 35736
rect 11374 35655 11438 35719
rect 11310 35638 11502 35655
rect 11374 35574 11438 35638
rect 11310 35557 11502 35574
rect 11374 35493 11438 35557
rect 11310 35476 11502 35493
rect 11374 35412 11438 35476
rect 11310 35395 11502 35412
rect 11374 35331 11438 35395
rect 11310 35314 11502 35331
rect 11374 35250 11438 35314
rect 11310 35233 11502 35250
rect 11374 35169 11438 35233
rect 11310 35152 11502 35169
rect 11374 35088 11438 35152
rect 11310 35071 11502 35088
rect 11374 35007 11438 35071
rect 11310 34990 11502 35007
rect 11374 34926 11438 34990
rect 11310 34909 11502 34926
rect 11374 34845 11438 34909
rect 11310 34828 11502 34845
rect 11374 34764 11438 34828
rect 10318 31962 10323 32018
rect 10379 31962 10449 32018
rect 10505 31962 10510 32018
rect 10318 31936 10510 31962
rect 10318 31880 10323 31936
rect 10379 31880 10449 31936
rect 10505 31880 10510 31936
rect 10318 31854 10510 31880
rect 10318 31798 10323 31854
rect 10379 31798 10449 31854
rect 10505 31798 10510 31854
rect 10318 31772 10510 31798
rect 10318 31716 10323 31772
rect 10379 31716 10449 31772
rect 10505 31716 10510 31772
rect 10318 31690 10510 31716
rect 10318 31634 10323 31690
rect 10379 31634 10449 31690
rect 10505 31634 10510 31690
rect 10318 31608 10510 31634
rect 10318 31552 10323 31608
rect 10379 31552 10449 31608
rect 10505 31552 10510 31608
rect 10318 31526 10510 31552
rect 10318 31470 10323 31526
rect 10379 31470 10449 31526
rect 10505 31470 10510 31526
rect 10318 31444 10510 31470
rect 10318 31388 10323 31444
rect 10379 31388 10449 31444
rect 10505 31388 10510 31444
rect 10318 31362 10510 31388
rect 10318 31306 10323 31362
rect 10379 31306 10449 31362
rect 10505 31306 10510 31362
rect 10318 31280 10510 31306
rect 10318 31224 10323 31280
rect 10379 31224 10449 31280
rect 10505 31224 10510 31280
rect 10318 31198 10510 31224
rect 10318 31142 10323 31198
rect 10379 31142 10449 31198
rect 10505 31142 10510 31198
rect 10318 31116 10510 31142
rect 10318 31060 10323 31116
rect 10379 31060 10449 31116
rect 10505 31060 10510 31116
rect 10318 31034 10510 31060
rect 10318 30978 10323 31034
rect 10379 30978 10449 31034
rect 10505 30978 10510 31034
rect 10318 30952 10510 30978
rect 10318 30896 10323 30952
rect 10379 30896 10449 30952
rect 10505 30896 10510 30952
rect 10318 30870 10510 30896
rect 10318 30814 10323 30870
rect 10379 30814 10449 30870
rect 10505 30814 10510 30870
rect 10318 30788 10510 30814
rect 10318 30732 10323 30788
rect 10379 30732 10449 30788
rect 10505 30732 10510 30788
rect 10318 30706 10510 30732
rect 10318 30650 10323 30706
rect 10379 30650 10449 30706
rect 10505 30650 10510 30706
rect 10318 30624 10510 30650
rect 10318 30568 10323 30624
rect 10379 30568 10449 30624
rect 10505 30568 10510 30624
rect 10318 30542 10510 30568
rect 10318 30486 10323 30542
rect 10379 30486 10449 30542
rect 10505 30486 10510 30542
rect 10318 30460 10510 30486
rect 10318 30404 10323 30460
rect 10379 30404 10449 30460
rect 10505 30404 10510 30460
rect 10318 30378 10510 30404
rect 10318 30322 10323 30378
rect 10379 30322 10449 30378
rect 10505 30322 10510 30378
rect 10318 30296 10510 30322
rect 10318 30240 10323 30296
rect 10379 30240 10449 30296
rect 10505 30240 10510 30296
rect 10318 30214 10510 30240
rect 10318 30158 10323 30214
rect 10379 30158 10449 30214
rect 10505 30158 10510 30214
rect 10318 30132 10510 30158
rect 10318 30076 10323 30132
rect 10379 30076 10449 30132
rect 10505 30076 10510 30132
rect 10318 30050 10510 30076
rect 10318 29994 10323 30050
rect 10379 29994 10449 30050
rect 10505 29994 10510 30050
rect 10318 29968 10510 29994
rect 10318 29912 10323 29968
rect 10379 29912 10449 29968
rect 10505 29912 10510 29968
rect 10318 29886 10510 29912
rect 10318 29830 10323 29886
rect 10379 29830 10449 29886
rect 10505 29830 10510 29886
rect 10318 29804 10510 29830
rect 10318 29748 10323 29804
rect 10379 29748 10449 29804
rect 10505 29748 10510 29804
rect 10318 29722 10510 29748
rect 10318 29666 10323 29722
rect 10379 29666 10449 29722
rect 10505 29666 10510 29722
rect 10318 29640 10510 29666
rect 10318 29584 10323 29640
rect 10379 29584 10449 29640
rect 10505 29584 10510 29640
rect 10318 29558 10510 29584
rect 10318 29502 10323 29558
rect 10379 29502 10449 29558
rect 10505 29502 10510 29558
rect 10318 29476 10510 29502
rect 10318 29420 10323 29476
rect 10379 29420 10449 29476
rect 10505 29420 10510 29476
rect 10318 29415 10510 29420
rect 10814 34219 11006 34225
rect 10878 34155 10942 34219
rect 10814 34125 11006 34155
rect 10878 34061 10942 34125
rect 10814 34030 11006 34061
rect 10878 33966 10942 34030
rect 10814 33935 11006 33966
rect 10878 33871 10942 33935
rect 10814 33840 11006 33871
rect 10878 33776 10942 33840
rect 10814 33745 11006 33776
rect 10878 33681 10942 33745
rect 10814 32018 11006 33681
rect 10814 31962 10819 32018
rect 10875 31962 10945 32018
rect 11001 31962 11006 32018
rect 10814 31936 11006 31962
rect 10814 31880 10819 31936
rect 10875 31880 10945 31936
rect 11001 31880 11006 31936
rect 10814 31854 11006 31880
rect 10814 31798 10819 31854
rect 10875 31798 10945 31854
rect 11001 31798 11006 31854
rect 10814 31772 11006 31798
rect 10814 31716 10819 31772
rect 10875 31716 10945 31772
rect 11001 31716 11006 31772
rect 10814 31690 11006 31716
rect 10814 31634 10819 31690
rect 10875 31634 10945 31690
rect 11001 31634 11006 31690
rect 10814 31608 11006 31634
rect 10814 31552 10819 31608
rect 10875 31552 10945 31608
rect 11001 31552 11006 31608
rect 10814 31526 11006 31552
rect 10814 31470 10819 31526
rect 10875 31470 10945 31526
rect 11001 31470 11006 31526
rect 10814 31444 11006 31470
rect 10814 31388 10819 31444
rect 10875 31388 10945 31444
rect 11001 31388 11006 31444
rect 10814 31362 11006 31388
rect 10814 31306 10819 31362
rect 10875 31306 10945 31362
rect 11001 31306 11006 31362
rect 10814 31280 11006 31306
rect 10814 31224 10819 31280
rect 10875 31224 10945 31280
rect 11001 31224 11006 31280
rect 10814 31198 11006 31224
rect 10814 31142 10819 31198
rect 10875 31142 10945 31198
rect 11001 31142 11006 31198
rect 10814 31116 11006 31142
rect 10814 31060 10819 31116
rect 10875 31060 10945 31116
rect 11001 31060 11006 31116
rect 10814 31034 11006 31060
rect 10814 30978 10819 31034
rect 10875 30978 10945 31034
rect 11001 30978 11006 31034
rect 10814 30952 11006 30978
rect 10814 30896 10819 30952
rect 10875 30896 10945 30952
rect 11001 30896 11006 30952
rect 10814 30870 11006 30896
rect 10814 30814 10819 30870
rect 10875 30814 10945 30870
rect 11001 30814 11006 30870
rect 10814 30788 11006 30814
rect 10814 30732 10819 30788
rect 10875 30732 10945 30788
rect 11001 30732 11006 30788
rect 10814 30706 11006 30732
rect 10814 30650 10819 30706
rect 10875 30650 10945 30706
rect 11001 30650 11006 30706
rect 10814 30624 11006 30650
rect 10814 30568 10819 30624
rect 10875 30568 10945 30624
rect 11001 30568 11006 30624
rect 10814 30542 11006 30568
rect 10814 30486 10819 30542
rect 10875 30486 10945 30542
rect 11001 30486 11006 30542
rect 10814 30460 11006 30486
rect 10814 30404 10819 30460
rect 10875 30404 10945 30460
rect 11001 30404 11006 30460
rect 10814 30378 11006 30404
rect 10814 30322 10819 30378
rect 10875 30322 10945 30378
rect 11001 30322 11006 30378
rect 10814 30296 11006 30322
rect 10814 30240 10819 30296
rect 10875 30240 10945 30296
rect 11001 30240 11006 30296
rect 10814 30214 11006 30240
rect 10814 30158 10819 30214
rect 10875 30158 10945 30214
rect 11001 30158 11006 30214
rect 10814 30132 11006 30158
rect 10814 30076 10819 30132
rect 10875 30076 10945 30132
rect 11001 30076 11006 30132
rect 10814 30050 11006 30076
rect 10814 29994 10819 30050
rect 10875 29994 10945 30050
rect 11001 29994 11006 30050
rect 10814 29968 11006 29994
rect 10814 29912 10819 29968
rect 10875 29912 10945 29968
rect 11001 29912 11006 29968
rect 10814 29886 11006 29912
rect 10814 29830 10819 29886
rect 10875 29830 10945 29886
rect 11001 29830 11006 29886
rect 10814 29804 11006 29830
rect 10814 29748 10819 29804
rect 10875 29748 10945 29804
rect 11001 29748 11006 29804
rect 10814 29722 11006 29748
rect 10814 29666 10819 29722
rect 10875 29666 10945 29722
rect 11001 29666 11006 29722
rect 10814 29640 11006 29666
rect 10814 29584 10819 29640
rect 10875 29584 10945 29640
rect 11001 29584 11006 29640
rect 10814 29558 11006 29584
rect 10814 29502 10819 29558
rect 10875 29502 10945 29558
rect 11001 29502 11006 29558
rect 10814 29476 11006 29502
rect 10814 29420 10819 29476
rect 10875 29420 10945 29476
rect 11001 29420 11006 29476
tri 10014 27161 10048 27195 sw
rect 10814 27161 11006 29420
rect 11310 32018 11502 34764
rect 12302 39592 12494 39600
rect 12366 39528 12430 39592
rect 12302 39512 12494 39528
rect 12366 39448 12430 39512
rect 12302 39432 12494 39448
rect 12366 39368 12430 39432
rect 12302 39352 12494 39368
rect 12366 39288 12430 39352
rect 12302 39272 12494 39288
rect 12366 39208 12430 39272
rect 12302 39192 12494 39208
rect 12366 39128 12430 39192
rect 12302 39112 12494 39128
rect 12366 39048 12430 39112
rect 12302 39032 12494 39048
rect 12366 38968 12430 39032
rect 12302 38952 12494 38968
rect 12366 38888 12430 38952
rect 12302 38872 12494 38888
rect 12366 38808 12430 38872
rect 12302 38792 12494 38808
rect 12366 38728 12430 38792
rect 12302 38712 12494 38728
rect 12366 38648 12430 38712
rect 12302 38632 12494 38648
rect 12366 38568 12430 38632
rect 12302 38552 12494 38568
rect 12366 38488 12430 38552
rect 12302 38472 12494 38488
rect 12366 38408 12430 38472
rect 12302 38392 12494 38408
rect 12366 38328 12430 38392
rect 12302 38311 12494 38328
rect 12366 38247 12430 38311
rect 12302 38230 12494 38247
rect 12366 38166 12430 38230
rect 12302 38149 12494 38166
rect 12366 38085 12430 38149
rect 12302 38068 12494 38085
rect 12366 38004 12430 38068
rect 12302 37987 12494 38004
rect 12366 37923 12430 37987
rect 12302 37906 12494 37923
rect 12366 37842 12430 37906
rect 12302 37825 12494 37842
rect 12366 37761 12430 37825
rect 12302 37744 12494 37761
rect 12366 37680 12430 37744
rect 12302 37663 12494 37680
rect 12366 37599 12430 37663
rect 12302 37582 12494 37599
rect 12366 37518 12430 37582
rect 12302 37501 12494 37518
rect 12366 37437 12430 37501
rect 12302 37420 12494 37437
rect 12366 37356 12430 37420
rect 12302 37339 12494 37356
rect 12366 37275 12430 37339
rect 12302 37258 12494 37275
rect 12366 37194 12430 37258
rect 12302 37177 12494 37194
rect 12366 37113 12430 37177
rect 12302 37096 12494 37113
rect 12366 37032 12430 37096
rect 12302 37015 12494 37032
rect 12366 36951 12430 37015
rect 12302 36934 12494 36951
rect 12366 36870 12430 36934
rect 12302 36853 12494 36870
rect 12366 36789 12430 36853
rect 12302 36772 12494 36789
rect 12366 36708 12430 36772
rect 12302 36691 12494 36708
rect 12366 36627 12430 36691
rect 12302 36610 12494 36627
rect 12366 36546 12430 36610
rect 12302 36529 12494 36546
rect 12366 36465 12430 36529
rect 12302 36448 12494 36465
rect 12366 36384 12430 36448
rect 12302 36367 12494 36384
rect 12366 36303 12430 36367
rect 12302 36286 12494 36303
rect 12366 36222 12430 36286
rect 12302 36205 12494 36222
rect 12366 36141 12430 36205
rect 12302 36124 12494 36141
rect 12366 36060 12430 36124
rect 12302 36043 12494 36060
rect 12366 35979 12430 36043
rect 12302 35962 12494 35979
rect 12366 35898 12430 35962
rect 12302 35881 12494 35898
rect 12366 35817 12430 35881
rect 12302 35800 12494 35817
rect 12366 35736 12430 35800
rect 12302 35719 12494 35736
rect 12366 35655 12430 35719
rect 12302 35638 12494 35655
rect 12366 35574 12430 35638
rect 12302 35557 12494 35574
rect 12366 35493 12430 35557
rect 12302 35476 12494 35493
rect 12366 35412 12430 35476
rect 12302 35395 12494 35412
rect 12366 35331 12430 35395
rect 12302 35314 12494 35331
rect 12366 35250 12430 35314
rect 12302 35233 12494 35250
rect 12366 35169 12430 35233
rect 12302 35152 12494 35169
rect 12366 35088 12430 35152
rect 12302 35071 12494 35088
rect 12366 35007 12430 35071
rect 12302 34990 12494 35007
rect 12366 34926 12430 34990
rect 12302 34909 12494 34926
rect 12366 34845 12430 34909
rect 12302 34828 12494 34845
rect 12366 34764 12430 34828
rect 11310 31962 11315 32018
rect 11371 31962 11441 32018
rect 11497 31962 11502 32018
rect 11310 31936 11502 31962
rect 11310 31880 11315 31936
rect 11371 31880 11441 31936
rect 11497 31880 11502 31936
rect 11310 31854 11502 31880
rect 11310 31798 11315 31854
rect 11371 31798 11441 31854
rect 11497 31798 11502 31854
rect 11310 31772 11502 31798
rect 11310 31716 11315 31772
rect 11371 31716 11441 31772
rect 11497 31716 11502 31772
rect 11310 31690 11502 31716
rect 11310 31634 11315 31690
rect 11371 31634 11441 31690
rect 11497 31634 11502 31690
rect 11310 31608 11502 31634
rect 11310 31552 11315 31608
rect 11371 31552 11441 31608
rect 11497 31552 11502 31608
rect 11310 31526 11502 31552
rect 11310 31470 11315 31526
rect 11371 31470 11441 31526
rect 11497 31470 11502 31526
rect 11310 31444 11502 31470
rect 11310 31388 11315 31444
rect 11371 31388 11441 31444
rect 11497 31388 11502 31444
rect 11310 31362 11502 31388
rect 11310 31306 11315 31362
rect 11371 31306 11441 31362
rect 11497 31306 11502 31362
rect 11310 31280 11502 31306
rect 11310 31224 11315 31280
rect 11371 31224 11441 31280
rect 11497 31224 11502 31280
rect 11310 31198 11502 31224
rect 11310 31142 11315 31198
rect 11371 31142 11441 31198
rect 11497 31142 11502 31198
rect 11310 31116 11502 31142
rect 11310 31060 11315 31116
rect 11371 31060 11441 31116
rect 11497 31060 11502 31116
rect 11310 31034 11502 31060
rect 11310 30978 11315 31034
rect 11371 30978 11441 31034
rect 11497 30978 11502 31034
rect 11310 30952 11502 30978
rect 11310 30896 11315 30952
rect 11371 30896 11441 30952
rect 11497 30896 11502 30952
rect 11310 30870 11502 30896
rect 11310 30814 11315 30870
rect 11371 30814 11441 30870
rect 11497 30814 11502 30870
rect 11310 30788 11502 30814
rect 11310 30732 11315 30788
rect 11371 30732 11441 30788
rect 11497 30732 11502 30788
rect 11310 30706 11502 30732
rect 11310 30650 11315 30706
rect 11371 30650 11441 30706
rect 11497 30650 11502 30706
rect 11310 30624 11502 30650
rect 11310 30568 11315 30624
rect 11371 30568 11441 30624
rect 11497 30568 11502 30624
rect 11310 30542 11502 30568
rect 11310 30486 11315 30542
rect 11371 30486 11441 30542
rect 11497 30486 11502 30542
rect 11310 30460 11502 30486
rect 11310 30404 11315 30460
rect 11371 30404 11441 30460
rect 11497 30404 11502 30460
rect 11310 30378 11502 30404
rect 11310 30322 11315 30378
rect 11371 30322 11441 30378
rect 11497 30322 11502 30378
rect 11310 30296 11502 30322
rect 11310 30240 11315 30296
rect 11371 30240 11441 30296
rect 11497 30240 11502 30296
rect 11310 30214 11502 30240
rect 11310 30158 11315 30214
rect 11371 30158 11441 30214
rect 11497 30158 11502 30214
rect 11310 30132 11502 30158
rect 11310 30076 11315 30132
rect 11371 30076 11441 30132
rect 11497 30076 11502 30132
rect 11310 30050 11502 30076
rect 11310 29994 11315 30050
rect 11371 29994 11441 30050
rect 11497 29994 11502 30050
rect 11310 29968 11502 29994
rect 11310 29912 11315 29968
rect 11371 29912 11441 29968
rect 11497 29912 11502 29968
rect 11310 29886 11502 29912
rect 11310 29830 11315 29886
rect 11371 29830 11441 29886
rect 11497 29830 11502 29886
rect 11310 29804 11502 29830
rect 11310 29748 11315 29804
rect 11371 29748 11441 29804
rect 11497 29748 11502 29804
rect 11310 29722 11502 29748
rect 11310 29666 11315 29722
rect 11371 29666 11441 29722
rect 11497 29666 11502 29722
rect 11310 29640 11502 29666
rect 11310 29584 11315 29640
rect 11371 29584 11441 29640
rect 11497 29584 11502 29640
rect 11310 29558 11502 29584
rect 11310 29502 11315 29558
rect 11371 29502 11441 29558
rect 11497 29502 11502 29558
rect 11310 29476 11502 29502
rect 11310 29420 11315 29476
rect 11371 29420 11441 29476
rect 11497 29420 11502 29476
rect 11310 29415 11502 29420
rect 11806 34219 11998 34225
rect 11870 34155 11934 34219
rect 11806 34125 11998 34155
rect 11870 34061 11934 34125
rect 11806 34030 11998 34061
rect 11870 33966 11934 34030
rect 11806 33935 11998 33966
rect 11870 33871 11934 33935
rect 11806 33840 11998 33871
rect 11870 33776 11934 33840
rect 11806 33745 11998 33776
rect 11870 33681 11934 33745
rect 11806 32018 11998 33681
rect 11806 31962 11811 32018
rect 11867 31962 11937 32018
rect 11993 31962 11998 32018
rect 11806 31936 11998 31962
rect 11806 31880 11811 31936
rect 11867 31880 11937 31936
rect 11993 31880 11998 31936
rect 11806 31854 11998 31880
rect 11806 31798 11811 31854
rect 11867 31798 11937 31854
rect 11993 31798 11998 31854
rect 11806 31772 11998 31798
rect 11806 31716 11811 31772
rect 11867 31716 11937 31772
rect 11993 31716 11998 31772
rect 11806 31690 11998 31716
rect 11806 31634 11811 31690
rect 11867 31634 11937 31690
rect 11993 31634 11998 31690
rect 11806 31608 11998 31634
rect 11806 31552 11811 31608
rect 11867 31552 11937 31608
rect 11993 31552 11998 31608
rect 11806 31526 11998 31552
rect 11806 31470 11811 31526
rect 11867 31470 11937 31526
rect 11993 31470 11998 31526
rect 11806 31444 11998 31470
rect 11806 31388 11811 31444
rect 11867 31388 11937 31444
rect 11993 31388 11998 31444
rect 11806 31362 11998 31388
rect 11806 31306 11811 31362
rect 11867 31306 11937 31362
rect 11993 31306 11998 31362
rect 11806 31280 11998 31306
rect 11806 31224 11811 31280
rect 11867 31224 11937 31280
rect 11993 31224 11998 31280
rect 11806 31198 11998 31224
rect 11806 31142 11811 31198
rect 11867 31142 11937 31198
rect 11993 31142 11998 31198
rect 11806 31116 11998 31142
rect 11806 31060 11811 31116
rect 11867 31060 11937 31116
rect 11993 31060 11998 31116
rect 11806 31034 11998 31060
rect 11806 30978 11811 31034
rect 11867 30978 11937 31034
rect 11993 30978 11998 31034
rect 11806 30952 11998 30978
rect 11806 30896 11811 30952
rect 11867 30896 11937 30952
rect 11993 30896 11998 30952
rect 11806 30870 11998 30896
rect 11806 30814 11811 30870
rect 11867 30814 11937 30870
rect 11993 30814 11998 30870
rect 11806 30788 11998 30814
rect 11806 30732 11811 30788
rect 11867 30732 11937 30788
rect 11993 30732 11998 30788
rect 11806 30706 11998 30732
rect 11806 30650 11811 30706
rect 11867 30650 11937 30706
rect 11993 30650 11998 30706
rect 11806 30624 11998 30650
rect 11806 30568 11811 30624
rect 11867 30568 11937 30624
rect 11993 30568 11998 30624
rect 11806 30542 11998 30568
rect 11806 30486 11811 30542
rect 11867 30486 11937 30542
rect 11993 30486 11998 30542
rect 11806 30460 11998 30486
rect 11806 30404 11811 30460
rect 11867 30404 11937 30460
rect 11993 30404 11998 30460
rect 11806 30378 11998 30404
rect 11806 30322 11811 30378
rect 11867 30322 11937 30378
rect 11993 30322 11998 30378
rect 11806 30296 11998 30322
rect 11806 30240 11811 30296
rect 11867 30240 11937 30296
rect 11993 30240 11998 30296
rect 11806 30214 11998 30240
rect 11806 30158 11811 30214
rect 11867 30158 11937 30214
rect 11993 30158 11998 30214
rect 11806 30132 11998 30158
rect 11806 30076 11811 30132
rect 11867 30076 11937 30132
rect 11993 30076 11998 30132
rect 11806 30050 11998 30076
rect 11806 29994 11811 30050
rect 11867 29994 11937 30050
rect 11993 29994 11998 30050
rect 11806 29968 11998 29994
rect 11806 29912 11811 29968
rect 11867 29912 11937 29968
rect 11993 29912 11998 29968
rect 11806 29886 11998 29912
rect 11806 29830 11811 29886
rect 11867 29830 11937 29886
rect 11993 29830 11998 29886
rect 11806 29804 11998 29830
rect 11806 29748 11811 29804
rect 11867 29748 11937 29804
rect 11993 29748 11998 29804
rect 11806 29722 11998 29748
rect 11806 29666 11811 29722
rect 11867 29666 11937 29722
rect 11993 29666 11998 29722
rect 11806 29640 11998 29666
rect 11806 29584 11811 29640
rect 11867 29584 11937 29640
rect 11993 29584 11998 29640
rect 11806 29558 11998 29584
rect 11806 29502 11811 29558
rect 11867 29502 11937 29558
rect 11993 29502 11998 29558
rect 11806 29476 11998 29502
rect 11806 29420 11811 29476
rect 11867 29420 11937 29476
rect 11993 29420 11998 29476
tri 11006 27161 11040 27195 sw
rect 11806 27161 11998 29420
rect 12302 32018 12494 34764
rect 13294 39592 13486 39600
rect 13358 39528 13422 39592
rect 13294 39512 13486 39528
rect 13358 39448 13422 39512
rect 13294 39432 13486 39448
rect 13358 39368 13422 39432
rect 13294 39352 13486 39368
rect 13358 39288 13422 39352
rect 13294 39272 13486 39288
rect 13358 39208 13422 39272
rect 13294 39192 13486 39208
rect 13358 39128 13422 39192
rect 13294 39112 13486 39128
rect 13358 39048 13422 39112
rect 13294 39032 13486 39048
rect 13358 38968 13422 39032
rect 13294 38952 13486 38968
rect 13358 38888 13422 38952
rect 13294 38872 13486 38888
rect 13358 38808 13422 38872
rect 13294 38792 13486 38808
rect 13358 38728 13422 38792
rect 13294 38712 13486 38728
rect 13358 38648 13422 38712
rect 13294 38632 13486 38648
rect 13358 38568 13422 38632
rect 13294 38552 13486 38568
rect 13358 38488 13422 38552
rect 13294 38472 13486 38488
rect 13358 38408 13422 38472
rect 13294 38392 13486 38408
rect 13358 38328 13422 38392
rect 13294 38311 13486 38328
rect 13358 38247 13422 38311
rect 13294 38230 13486 38247
rect 13358 38166 13422 38230
rect 13294 38149 13486 38166
rect 13358 38085 13422 38149
rect 13294 38068 13486 38085
rect 13358 38004 13422 38068
rect 13294 37987 13486 38004
rect 13358 37923 13422 37987
rect 13294 37906 13486 37923
rect 13358 37842 13422 37906
rect 13294 37825 13486 37842
rect 13358 37761 13422 37825
rect 13294 37744 13486 37761
rect 13358 37680 13422 37744
rect 13294 37663 13486 37680
rect 13358 37599 13422 37663
rect 13294 37582 13486 37599
rect 13358 37518 13422 37582
rect 13294 37501 13486 37518
rect 13358 37437 13422 37501
rect 13294 37420 13486 37437
rect 13358 37356 13422 37420
rect 13294 37339 13486 37356
rect 13358 37275 13422 37339
rect 13294 37258 13486 37275
rect 13358 37194 13422 37258
rect 13294 37177 13486 37194
rect 13358 37113 13422 37177
rect 13294 37096 13486 37113
rect 13358 37032 13422 37096
rect 13294 37015 13486 37032
rect 13358 36951 13422 37015
rect 13294 36934 13486 36951
rect 13358 36870 13422 36934
rect 13294 36853 13486 36870
rect 13358 36789 13422 36853
rect 13294 36772 13486 36789
rect 13358 36708 13422 36772
rect 13294 36691 13486 36708
rect 13358 36627 13422 36691
rect 13294 36610 13486 36627
rect 13358 36546 13422 36610
rect 13294 36529 13486 36546
rect 13358 36465 13422 36529
rect 13294 36448 13486 36465
rect 13358 36384 13422 36448
rect 13294 36367 13486 36384
rect 13358 36303 13422 36367
rect 13294 36286 13486 36303
rect 13358 36222 13422 36286
rect 13294 36205 13486 36222
rect 13358 36141 13422 36205
rect 13294 36124 13486 36141
rect 13358 36060 13422 36124
rect 13294 36043 13486 36060
rect 13358 35979 13422 36043
rect 13294 35962 13486 35979
rect 13358 35898 13422 35962
rect 13294 35881 13486 35898
rect 13358 35817 13422 35881
rect 13294 35800 13486 35817
rect 13358 35736 13422 35800
rect 13294 35719 13486 35736
rect 13358 35655 13422 35719
rect 13294 35638 13486 35655
rect 13358 35574 13422 35638
rect 13294 35557 13486 35574
rect 13358 35493 13422 35557
rect 13294 35476 13486 35493
rect 13358 35412 13422 35476
rect 13294 35395 13486 35412
rect 13358 35331 13422 35395
rect 13294 35314 13486 35331
rect 13358 35250 13422 35314
rect 13294 35233 13486 35250
rect 13358 35169 13422 35233
rect 13294 35152 13486 35169
rect 13358 35088 13422 35152
rect 13294 35071 13486 35088
rect 13358 35007 13422 35071
rect 13294 34990 13486 35007
rect 13358 34926 13422 34990
rect 13294 34909 13486 34926
rect 13358 34845 13422 34909
rect 13294 34828 13486 34845
rect 13358 34764 13422 34828
rect 12302 31962 12307 32018
rect 12363 31962 12433 32018
rect 12489 31962 12494 32018
rect 12302 31936 12494 31962
rect 12302 31880 12307 31936
rect 12363 31880 12433 31936
rect 12489 31880 12494 31936
rect 12302 31854 12494 31880
rect 12302 31798 12307 31854
rect 12363 31798 12433 31854
rect 12489 31798 12494 31854
rect 12302 31772 12494 31798
rect 12302 31716 12307 31772
rect 12363 31716 12433 31772
rect 12489 31716 12494 31772
rect 12302 31690 12494 31716
rect 12302 31634 12307 31690
rect 12363 31634 12433 31690
rect 12489 31634 12494 31690
rect 12302 31608 12494 31634
rect 12302 31552 12307 31608
rect 12363 31552 12433 31608
rect 12489 31552 12494 31608
rect 12302 31526 12494 31552
rect 12302 31470 12307 31526
rect 12363 31470 12433 31526
rect 12489 31470 12494 31526
rect 12302 31444 12494 31470
rect 12302 31388 12307 31444
rect 12363 31388 12433 31444
rect 12489 31388 12494 31444
rect 12302 31362 12494 31388
rect 12302 31306 12307 31362
rect 12363 31306 12433 31362
rect 12489 31306 12494 31362
rect 12302 31280 12494 31306
rect 12302 31224 12307 31280
rect 12363 31224 12433 31280
rect 12489 31224 12494 31280
rect 12302 31198 12494 31224
rect 12302 31142 12307 31198
rect 12363 31142 12433 31198
rect 12489 31142 12494 31198
rect 12302 31116 12494 31142
rect 12302 31060 12307 31116
rect 12363 31060 12433 31116
rect 12489 31060 12494 31116
rect 12302 31034 12494 31060
rect 12302 30978 12307 31034
rect 12363 30978 12433 31034
rect 12489 30978 12494 31034
rect 12302 30952 12494 30978
rect 12302 30896 12307 30952
rect 12363 30896 12433 30952
rect 12489 30896 12494 30952
rect 12302 30870 12494 30896
rect 12302 30814 12307 30870
rect 12363 30814 12433 30870
rect 12489 30814 12494 30870
rect 12302 30788 12494 30814
rect 12302 30732 12307 30788
rect 12363 30732 12433 30788
rect 12489 30732 12494 30788
rect 12302 30706 12494 30732
rect 12302 30650 12307 30706
rect 12363 30650 12433 30706
rect 12489 30650 12494 30706
rect 12302 30624 12494 30650
rect 12302 30568 12307 30624
rect 12363 30568 12433 30624
rect 12489 30568 12494 30624
rect 12302 30542 12494 30568
rect 12302 30486 12307 30542
rect 12363 30486 12433 30542
rect 12489 30486 12494 30542
rect 12302 30460 12494 30486
rect 12302 30404 12307 30460
rect 12363 30404 12433 30460
rect 12489 30404 12494 30460
rect 12302 30378 12494 30404
rect 12302 30322 12307 30378
rect 12363 30322 12433 30378
rect 12489 30322 12494 30378
rect 12302 30296 12494 30322
rect 12302 30240 12307 30296
rect 12363 30240 12433 30296
rect 12489 30240 12494 30296
rect 12302 30214 12494 30240
rect 12302 30158 12307 30214
rect 12363 30158 12433 30214
rect 12489 30158 12494 30214
rect 12302 30132 12494 30158
rect 12302 30076 12307 30132
rect 12363 30076 12433 30132
rect 12489 30076 12494 30132
rect 12302 30050 12494 30076
rect 12302 29994 12307 30050
rect 12363 29994 12433 30050
rect 12489 29994 12494 30050
rect 12302 29968 12494 29994
rect 12302 29912 12307 29968
rect 12363 29912 12433 29968
rect 12489 29912 12494 29968
rect 12302 29886 12494 29912
rect 12302 29830 12307 29886
rect 12363 29830 12433 29886
rect 12489 29830 12494 29886
rect 12302 29804 12494 29830
rect 12302 29748 12307 29804
rect 12363 29748 12433 29804
rect 12489 29748 12494 29804
rect 12302 29722 12494 29748
rect 12302 29666 12307 29722
rect 12363 29666 12433 29722
rect 12489 29666 12494 29722
rect 12302 29640 12494 29666
rect 12302 29584 12307 29640
rect 12363 29584 12433 29640
rect 12489 29584 12494 29640
rect 12302 29558 12494 29584
rect 12302 29502 12307 29558
rect 12363 29502 12433 29558
rect 12489 29502 12494 29558
rect 12302 29476 12494 29502
rect 12302 29420 12307 29476
rect 12363 29420 12433 29476
rect 12489 29420 12494 29476
rect 12302 29415 12494 29420
rect 12798 33954 12990 33960
rect 12862 33890 12926 33954
rect 12798 33860 12990 33890
rect 12862 33796 12926 33860
rect 12798 33765 12990 33796
rect 12862 33701 12926 33765
rect 12798 33670 12990 33701
rect 12862 33606 12926 33670
rect 12798 33575 12990 33606
rect 12862 33511 12926 33575
rect 12798 33480 12990 33511
rect 12862 33416 12926 33480
rect 12798 32018 12990 33416
rect 12798 31962 12803 32018
rect 12859 31962 12929 32018
rect 12985 31962 12990 32018
rect 12798 31936 12990 31962
rect 12798 31880 12803 31936
rect 12859 31880 12929 31936
rect 12985 31880 12990 31936
rect 12798 31854 12990 31880
rect 12798 31798 12803 31854
rect 12859 31798 12929 31854
rect 12985 31798 12990 31854
rect 12798 31772 12990 31798
rect 12798 31716 12803 31772
rect 12859 31716 12929 31772
rect 12985 31716 12990 31772
rect 12798 31690 12990 31716
rect 12798 31634 12803 31690
rect 12859 31634 12929 31690
rect 12985 31634 12990 31690
rect 12798 31608 12990 31634
rect 12798 31552 12803 31608
rect 12859 31552 12929 31608
rect 12985 31552 12990 31608
rect 12798 31526 12990 31552
rect 12798 31470 12803 31526
rect 12859 31470 12929 31526
rect 12985 31470 12990 31526
rect 12798 31444 12990 31470
rect 12798 31388 12803 31444
rect 12859 31388 12929 31444
rect 12985 31388 12990 31444
rect 12798 31362 12990 31388
rect 12798 31306 12803 31362
rect 12859 31306 12929 31362
rect 12985 31306 12990 31362
rect 12798 31280 12990 31306
rect 12798 31224 12803 31280
rect 12859 31224 12929 31280
rect 12985 31224 12990 31280
rect 12798 31198 12990 31224
rect 12798 31142 12803 31198
rect 12859 31142 12929 31198
rect 12985 31142 12990 31198
rect 12798 31116 12990 31142
rect 12798 31060 12803 31116
rect 12859 31060 12929 31116
rect 12985 31060 12990 31116
rect 12798 31034 12990 31060
rect 12798 30978 12803 31034
rect 12859 30978 12929 31034
rect 12985 30978 12990 31034
rect 12798 30952 12990 30978
rect 12798 30896 12803 30952
rect 12859 30896 12929 30952
rect 12985 30896 12990 30952
rect 12798 30870 12990 30896
rect 12798 30814 12803 30870
rect 12859 30814 12929 30870
rect 12985 30814 12990 30870
rect 12798 30788 12990 30814
rect 12798 30732 12803 30788
rect 12859 30732 12929 30788
rect 12985 30732 12990 30788
rect 12798 30706 12990 30732
rect 12798 30650 12803 30706
rect 12859 30650 12929 30706
rect 12985 30650 12990 30706
rect 12798 30624 12990 30650
rect 12798 30568 12803 30624
rect 12859 30568 12929 30624
rect 12985 30568 12990 30624
rect 12798 30542 12990 30568
rect 12798 30486 12803 30542
rect 12859 30486 12929 30542
rect 12985 30486 12990 30542
rect 12798 30460 12990 30486
rect 12798 30404 12803 30460
rect 12859 30404 12929 30460
rect 12985 30404 12990 30460
rect 12798 30378 12990 30404
rect 12798 30322 12803 30378
rect 12859 30322 12929 30378
rect 12985 30322 12990 30378
rect 12798 30296 12990 30322
rect 12798 30240 12803 30296
rect 12859 30240 12929 30296
rect 12985 30240 12990 30296
rect 12798 30214 12990 30240
rect 12798 30158 12803 30214
rect 12859 30158 12929 30214
rect 12985 30158 12990 30214
rect 12798 30132 12990 30158
rect 12798 30076 12803 30132
rect 12859 30076 12929 30132
rect 12985 30076 12990 30132
rect 12798 30050 12990 30076
rect 12798 29994 12803 30050
rect 12859 29994 12929 30050
rect 12985 29994 12990 30050
rect 12798 29968 12990 29994
rect 12798 29912 12803 29968
rect 12859 29912 12929 29968
rect 12985 29912 12990 29968
rect 12798 29886 12990 29912
rect 12798 29830 12803 29886
rect 12859 29830 12929 29886
rect 12985 29830 12990 29886
rect 12798 29804 12990 29830
rect 12798 29748 12803 29804
rect 12859 29748 12929 29804
rect 12985 29748 12990 29804
rect 12798 29722 12990 29748
rect 12798 29666 12803 29722
rect 12859 29666 12929 29722
rect 12985 29666 12990 29722
rect 12798 29640 12990 29666
rect 12798 29584 12803 29640
rect 12859 29584 12929 29640
rect 12985 29584 12990 29640
rect 12798 29558 12990 29584
rect 12798 29502 12803 29558
rect 12859 29502 12929 29558
rect 12985 29502 12990 29558
rect 12798 29476 12990 29502
rect 12798 29420 12803 29476
rect 12859 29420 12929 29476
rect 12985 29420 12990 29476
tri 11998 27161 12032 27195 sw
rect 12798 27161 12990 29420
rect 13294 32018 13486 34764
rect 14253 39592 14672 39600
rect 14253 39528 14255 39592
rect 14319 39528 14343 39592
rect 14407 39528 14431 39592
rect 14495 39528 14519 39592
rect 14583 39528 14607 39592
rect 14671 39528 14672 39592
rect 14253 39512 14672 39528
rect 14253 39448 14255 39512
rect 14319 39448 14343 39512
rect 14407 39448 14431 39512
rect 14495 39448 14519 39512
rect 14583 39448 14607 39512
rect 14671 39448 14672 39512
rect 14253 39432 14672 39448
rect 14253 39368 14255 39432
rect 14319 39368 14343 39432
rect 14407 39368 14431 39432
rect 14495 39368 14519 39432
rect 14583 39368 14607 39432
rect 14671 39368 14672 39432
rect 14253 39352 14672 39368
rect 14253 39288 14255 39352
rect 14319 39288 14343 39352
rect 14407 39288 14431 39352
rect 14495 39288 14519 39352
rect 14583 39288 14607 39352
rect 14671 39288 14672 39352
rect 14253 39272 14672 39288
rect 14253 39208 14255 39272
rect 14319 39208 14343 39272
rect 14407 39208 14431 39272
rect 14495 39208 14519 39272
rect 14583 39208 14607 39272
rect 14671 39208 14672 39272
rect 14253 39192 14672 39208
rect 14253 39128 14255 39192
rect 14319 39128 14343 39192
rect 14407 39128 14431 39192
rect 14495 39128 14519 39192
rect 14583 39128 14607 39192
rect 14671 39128 14672 39192
rect 14253 39112 14672 39128
rect 14253 39048 14255 39112
rect 14319 39048 14343 39112
rect 14407 39048 14431 39112
rect 14495 39048 14519 39112
rect 14583 39048 14607 39112
rect 14671 39048 14672 39112
rect 14253 39032 14672 39048
rect 14253 38968 14255 39032
rect 14319 38968 14343 39032
rect 14407 38968 14431 39032
rect 14495 38968 14519 39032
rect 14583 38968 14607 39032
rect 14671 38968 14672 39032
rect 14253 38952 14672 38968
rect 14253 38888 14255 38952
rect 14319 38888 14343 38952
rect 14407 38888 14431 38952
rect 14495 38888 14519 38952
rect 14583 38888 14607 38952
rect 14671 38888 14672 38952
rect 14253 38872 14672 38888
rect 14253 38808 14255 38872
rect 14319 38808 14343 38872
rect 14407 38808 14431 38872
rect 14495 38808 14519 38872
rect 14583 38808 14607 38872
rect 14671 38808 14672 38872
rect 14253 38792 14672 38808
rect 14253 38728 14255 38792
rect 14319 38728 14343 38792
rect 14407 38728 14431 38792
rect 14495 38728 14519 38792
rect 14583 38728 14607 38792
rect 14671 38728 14672 38792
rect 14253 38712 14672 38728
rect 14253 38648 14255 38712
rect 14319 38648 14343 38712
rect 14407 38648 14431 38712
rect 14495 38648 14519 38712
rect 14583 38648 14607 38712
rect 14671 38648 14672 38712
rect 14253 38632 14672 38648
rect 14253 38568 14255 38632
rect 14319 38568 14343 38632
rect 14407 38568 14431 38632
rect 14495 38568 14519 38632
rect 14583 38568 14607 38632
rect 14671 38568 14672 38632
rect 14253 38552 14672 38568
rect 14253 38488 14255 38552
rect 14319 38488 14343 38552
rect 14407 38488 14431 38552
rect 14495 38488 14519 38552
rect 14583 38488 14607 38552
rect 14671 38488 14672 38552
rect 14253 38472 14672 38488
rect 14253 38408 14255 38472
rect 14319 38408 14343 38472
rect 14407 38408 14431 38472
rect 14495 38408 14519 38472
rect 14583 38408 14607 38472
rect 14671 38408 14672 38472
rect 14253 38392 14672 38408
rect 14253 38328 14255 38392
rect 14319 38328 14343 38392
rect 14407 38328 14431 38392
rect 14495 38328 14519 38392
rect 14583 38328 14607 38392
rect 14671 38328 14672 38392
rect 14253 38311 14672 38328
rect 14253 38247 14255 38311
rect 14319 38247 14343 38311
rect 14407 38247 14431 38311
rect 14495 38247 14519 38311
rect 14583 38247 14607 38311
rect 14671 38247 14672 38311
rect 14253 38230 14672 38247
rect 14253 38166 14255 38230
rect 14319 38166 14343 38230
rect 14407 38166 14431 38230
rect 14495 38166 14519 38230
rect 14583 38166 14607 38230
rect 14671 38166 14672 38230
rect 14253 38149 14672 38166
rect 14253 38085 14255 38149
rect 14319 38085 14343 38149
rect 14407 38085 14431 38149
rect 14495 38085 14519 38149
rect 14583 38085 14607 38149
rect 14671 38085 14672 38149
rect 14253 38068 14672 38085
rect 14253 38004 14255 38068
rect 14319 38004 14343 38068
rect 14407 38004 14431 38068
rect 14495 38004 14519 38068
rect 14583 38004 14607 38068
rect 14671 38004 14672 38068
rect 14253 37987 14672 38004
rect 14253 37923 14255 37987
rect 14319 37923 14343 37987
rect 14407 37923 14431 37987
rect 14495 37923 14519 37987
rect 14583 37923 14607 37987
rect 14671 37923 14672 37987
rect 14253 37906 14672 37923
rect 14253 37842 14255 37906
rect 14319 37842 14343 37906
rect 14407 37842 14431 37906
rect 14495 37842 14519 37906
rect 14583 37842 14607 37906
rect 14671 37842 14672 37906
rect 14253 37825 14672 37842
rect 14253 37761 14255 37825
rect 14319 37761 14343 37825
rect 14407 37761 14431 37825
rect 14495 37761 14519 37825
rect 14583 37761 14607 37825
rect 14671 37761 14672 37825
rect 14253 37744 14672 37761
rect 14253 37680 14255 37744
rect 14319 37680 14343 37744
rect 14407 37680 14431 37744
rect 14495 37680 14519 37744
rect 14583 37680 14607 37744
rect 14671 37680 14672 37744
rect 14253 37663 14672 37680
rect 14253 37599 14255 37663
rect 14319 37599 14343 37663
rect 14407 37599 14431 37663
rect 14495 37599 14519 37663
rect 14583 37599 14607 37663
rect 14671 37599 14672 37663
rect 14253 37582 14672 37599
rect 14253 37518 14255 37582
rect 14319 37518 14343 37582
rect 14407 37518 14431 37582
rect 14495 37518 14519 37582
rect 14583 37518 14607 37582
rect 14671 37518 14672 37582
rect 14253 37501 14672 37518
rect 14253 37437 14255 37501
rect 14319 37437 14343 37501
rect 14407 37437 14431 37501
rect 14495 37437 14519 37501
rect 14583 37437 14607 37501
rect 14671 37437 14672 37501
rect 14253 37420 14672 37437
rect 14253 37356 14255 37420
rect 14319 37356 14343 37420
rect 14407 37356 14431 37420
rect 14495 37356 14519 37420
rect 14583 37356 14607 37420
rect 14671 37356 14672 37420
rect 14253 37339 14672 37356
rect 14253 37275 14255 37339
rect 14319 37275 14343 37339
rect 14407 37275 14431 37339
rect 14495 37275 14519 37339
rect 14583 37275 14607 37339
rect 14671 37275 14672 37339
rect 14253 37258 14672 37275
rect 14253 37194 14255 37258
rect 14319 37194 14343 37258
rect 14407 37194 14431 37258
rect 14495 37194 14519 37258
rect 14583 37194 14607 37258
rect 14671 37194 14672 37258
rect 14253 37177 14672 37194
rect 14253 37113 14255 37177
rect 14319 37113 14343 37177
rect 14407 37113 14431 37177
rect 14495 37113 14519 37177
rect 14583 37113 14607 37177
rect 14671 37113 14672 37177
rect 14253 37096 14672 37113
rect 14253 37032 14255 37096
rect 14319 37032 14343 37096
rect 14407 37032 14431 37096
rect 14495 37032 14519 37096
rect 14583 37032 14607 37096
rect 14671 37032 14672 37096
rect 14253 37015 14672 37032
rect 14253 36951 14255 37015
rect 14319 36951 14343 37015
rect 14407 36951 14431 37015
rect 14495 36951 14519 37015
rect 14583 36951 14607 37015
rect 14671 36951 14672 37015
rect 14253 36934 14672 36951
rect 14253 36870 14255 36934
rect 14319 36870 14343 36934
rect 14407 36870 14431 36934
rect 14495 36870 14519 36934
rect 14583 36870 14607 36934
rect 14671 36870 14672 36934
rect 14253 36853 14672 36870
rect 14253 36789 14255 36853
rect 14319 36789 14343 36853
rect 14407 36789 14431 36853
rect 14495 36789 14519 36853
rect 14583 36789 14607 36853
rect 14671 36789 14672 36853
rect 14253 36772 14672 36789
rect 14253 36708 14255 36772
rect 14319 36708 14343 36772
rect 14407 36708 14431 36772
rect 14495 36708 14519 36772
rect 14583 36708 14607 36772
rect 14671 36708 14672 36772
rect 14253 36691 14672 36708
rect 14253 36627 14255 36691
rect 14319 36627 14343 36691
rect 14407 36627 14431 36691
rect 14495 36627 14519 36691
rect 14583 36627 14607 36691
rect 14671 36627 14672 36691
rect 14253 36610 14672 36627
rect 14253 36546 14255 36610
rect 14319 36546 14343 36610
rect 14407 36546 14431 36610
rect 14495 36546 14519 36610
rect 14583 36546 14607 36610
rect 14671 36546 14672 36610
rect 14253 36529 14672 36546
rect 14253 36465 14255 36529
rect 14319 36465 14343 36529
rect 14407 36465 14431 36529
rect 14495 36465 14519 36529
rect 14583 36465 14607 36529
rect 14671 36465 14672 36529
rect 14253 36448 14672 36465
rect 14253 36384 14255 36448
rect 14319 36384 14343 36448
rect 14407 36384 14431 36448
rect 14495 36384 14519 36448
rect 14583 36384 14607 36448
rect 14671 36384 14672 36448
rect 14253 36367 14672 36384
rect 14253 36303 14255 36367
rect 14319 36303 14343 36367
rect 14407 36303 14431 36367
rect 14495 36303 14519 36367
rect 14583 36303 14607 36367
rect 14671 36303 14672 36367
rect 14253 36286 14672 36303
rect 14253 36222 14255 36286
rect 14319 36222 14343 36286
rect 14407 36222 14431 36286
rect 14495 36222 14519 36286
rect 14583 36222 14607 36286
rect 14671 36222 14672 36286
rect 14253 36205 14672 36222
rect 14253 36141 14255 36205
rect 14319 36141 14343 36205
rect 14407 36141 14431 36205
rect 14495 36141 14519 36205
rect 14583 36141 14607 36205
rect 14671 36141 14672 36205
rect 14253 36124 14672 36141
rect 14253 36060 14255 36124
rect 14319 36060 14343 36124
rect 14407 36060 14431 36124
rect 14495 36060 14519 36124
rect 14583 36060 14607 36124
rect 14671 36060 14672 36124
rect 14253 36043 14672 36060
rect 14253 35979 14255 36043
rect 14319 35979 14343 36043
rect 14407 35979 14431 36043
rect 14495 35979 14519 36043
rect 14583 35979 14607 36043
rect 14671 35979 14672 36043
rect 14253 35962 14672 35979
rect 14253 35898 14255 35962
rect 14319 35898 14343 35962
rect 14407 35898 14431 35962
rect 14495 35898 14519 35962
rect 14583 35898 14607 35962
rect 14671 35898 14672 35962
rect 14253 35881 14672 35898
rect 14253 35817 14255 35881
rect 14319 35817 14343 35881
rect 14407 35817 14431 35881
rect 14495 35817 14519 35881
rect 14583 35817 14607 35881
rect 14671 35817 14672 35881
rect 14253 35800 14672 35817
rect 14253 35736 14255 35800
rect 14319 35736 14343 35800
rect 14407 35736 14431 35800
rect 14495 35736 14519 35800
rect 14583 35736 14607 35800
rect 14671 35736 14672 35800
rect 14253 35719 14672 35736
rect 14253 35655 14255 35719
rect 14319 35655 14343 35719
rect 14407 35655 14431 35719
rect 14495 35655 14519 35719
rect 14583 35655 14607 35719
rect 14671 35655 14672 35719
rect 14253 35638 14672 35655
rect 14253 35574 14255 35638
rect 14319 35574 14343 35638
rect 14407 35574 14431 35638
rect 14495 35574 14519 35638
rect 14583 35574 14607 35638
rect 14671 35574 14672 35638
rect 14253 35557 14672 35574
rect 14253 35493 14255 35557
rect 14319 35493 14343 35557
rect 14407 35493 14431 35557
rect 14495 35493 14519 35557
rect 14583 35493 14607 35557
rect 14671 35493 14672 35557
rect 14253 35476 14672 35493
rect 14253 35412 14255 35476
rect 14319 35412 14343 35476
rect 14407 35412 14431 35476
rect 14495 35412 14519 35476
rect 14583 35412 14607 35476
rect 14671 35412 14672 35476
rect 14253 35395 14672 35412
rect 14253 35331 14255 35395
rect 14319 35331 14343 35395
rect 14407 35331 14431 35395
rect 14495 35331 14519 35395
rect 14583 35331 14607 35395
rect 14671 35331 14672 35395
rect 14253 35314 14672 35331
rect 14253 35250 14255 35314
rect 14319 35250 14343 35314
rect 14407 35250 14431 35314
rect 14495 35250 14519 35314
rect 14583 35250 14607 35314
rect 14671 35250 14672 35314
rect 14253 35233 14672 35250
rect 14253 35169 14255 35233
rect 14319 35169 14343 35233
rect 14407 35169 14431 35233
rect 14495 35169 14519 35233
rect 14583 35169 14607 35233
rect 14671 35169 14672 35233
rect 14253 35152 14672 35169
rect 14253 35088 14255 35152
rect 14319 35088 14343 35152
rect 14407 35088 14431 35152
rect 14495 35088 14519 35152
rect 14583 35088 14607 35152
rect 14671 35088 14672 35152
rect 14253 35071 14672 35088
rect 14253 35007 14255 35071
rect 14319 35007 14343 35071
rect 14407 35007 14431 35071
rect 14495 35007 14519 35071
rect 14583 35007 14607 35071
rect 14671 35007 14672 35071
rect 14253 34990 14672 35007
rect 14253 34926 14255 34990
rect 14319 34926 14343 34990
rect 14407 34926 14431 34990
rect 14495 34926 14519 34990
rect 14583 34926 14607 34990
rect 14671 34926 14672 34990
rect 14253 34909 14672 34926
rect 14253 34845 14255 34909
rect 14319 34845 14343 34909
rect 14407 34845 14431 34909
rect 14495 34845 14519 34909
rect 14583 34845 14607 34909
rect 14671 34845 14672 34909
rect 14253 34828 14672 34845
rect 14253 34764 14255 34828
rect 14319 34764 14343 34828
rect 14407 34764 14431 34828
rect 14495 34764 14519 34828
rect 14583 34764 14607 34828
rect 14671 34764 14672 34828
rect 13294 31962 13299 32018
rect 13355 31962 13425 32018
rect 13481 31962 13486 32018
rect 13294 31936 13486 31962
rect 13294 31880 13299 31936
rect 13355 31880 13425 31936
rect 13481 31880 13486 31936
rect 13294 31854 13486 31880
rect 13294 31798 13299 31854
rect 13355 31798 13425 31854
rect 13481 31798 13486 31854
rect 13294 31772 13486 31798
rect 13294 31716 13299 31772
rect 13355 31716 13425 31772
rect 13481 31716 13486 31772
rect 13294 31690 13486 31716
rect 13294 31634 13299 31690
rect 13355 31634 13425 31690
rect 13481 31634 13486 31690
rect 13294 31608 13486 31634
rect 13294 31552 13299 31608
rect 13355 31552 13425 31608
rect 13481 31552 13486 31608
rect 13294 31526 13486 31552
rect 13294 31470 13299 31526
rect 13355 31470 13425 31526
rect 13481 31470 13486 31526
rect 13294 31444 13486 31470
rect 13294 31388 13299 31444
rect 13355 31388 13425 31444
rect 13481 31388 13486 31444
rect 13294 31362 13486 31388
rect 13294 31306 13299 31362
rect 13355 31306 13425 31362
rect 13481 31306 13486 31362
rect 13294 31280 13486 31306
rect 13294 31224 13299 31280
rect 13355 31224 13425 31280
rect 13481 31224 13486 31280
rect 13294 31198 13486 31224
rect 13294 31142 13299 31198
rect 13355 31142 13425 31198
rect 13481 31142 13486 31198
rect 13294 31116 13486 31142
rect 13294 31060 13299 31116
rect 13355 31060 13425 31116
rect 13481 31060 13486 31116
rect 13294 31034 13486 31060
rect 13294 30978 13299 31034
rect 13355 30978 13425 31034
rect 13481 30978 13486 31034
rect 13294 30952 13486 30978
rect 13294 30896 13299 30952
rect 13355 30896 13425 30952
rect 13481 30896 13486 30952
rect 13294 30870 13486 30896
rect 13294 30814 13299 30870
rect 13355 30814 13425 30870
rect 13481 30814 13486 30870
rect 13294 30788 13486 30814
rect 13294 30732 13299 30788
rect 13355 30732 13425 30788
rect 13481 30732 13486 30788
rect 13294 30706 13486 30732
rect 13294 30650 13299 30706
rect 13355 30650 13425 30706
rect 13481 30650 13486 30706
rect 13294 30624 13486 30650
rect 13294 30568 13299 30624
rect 13355 30568 13425 30624
rect 13481 30568 13486 30624
rect 13294 30542 13486 30568
rect 13294 30486 13299 30542
rect 13355 30486 13425 30542
rect 13481 30486 13486 30542
rect 13294 30460 13486 30486
rect 13294 30404 13299 30460
rect 13355 30404 13425 30460
rect 13481 30404 13486 30460
rect 13294 30378 13486 30404
rect 13294 30322 13299 30378
rect 13355 30322 13425 30378
rect 13481 30322 13486 30378
rect 13294 30296 13486 30322
rect 13294 30240 13299 30296
rect 13355 30240 13425 30296
rect 13481 30240 13486 30296
rect 13294 30214 13486 30240
rect 13294 30158 13299 30214
rect 13355 30158 13425 30214
rect 13481 30158 13486 30214
rect 13294 30132 13486 30158
rect 13294 30076 13299 30132
rect 13355 30076 13425 30132
rect 13481 30076 13486 30132
rect 13294 30050 13486 30076
rect 13294 29994 13299 30050
rect 13355 29994 13425 30050
rect 13481 29994 13486 30050
rect 13294 29968 13486 29994
rect 13294 29912 13299 29968
rect 13355 29912 13425 29968
rect 13481 29912 13486 29968
rect 13294 29886 13486 29912
rect 13294 29830 13299 29886
rect 13355 29830 13425 29886
rect 13481 29830 13486 29886
rect 13294 29804 13486 29830
rect 13294 29748 13299 29804
rect 13355 29748 13425 29804
rect 13481 29748 13486 29804
rect 13294 29722 13486 29748
rect 13294 29666 13299 29722
rect 13355 29666 13425 29722
rect 13481 29666 13486 29722
rect 13294 29640 13486 29666
rect 13294 29584 13299 29640
rect 13355 29584 13425 29640
rect 13481 29584 13486 29640
rect 13294 29558 13486 29584
rect 13294 29502 13299 29558
rect 13355 29502 13425 29558
rect 13481 29502 13486 29558
rect 13294 29476 13486 29502
rect 13294 29420 13299 29476
rect 13355 29420 13425 29476
rect 13481 29420 13486 29476
rect 13294 29415 13486 29420
rect 13790 32983 13982 32989
rect 13854 32919 13892 32983
rect 13956 32919 13982 32983
rect 13790 32903 13982 32919
rect 13854 32839 13892 32903
rect 13956 32839 13982 32903
rect 13790 32823 13982 32839
rect 13854 32759 13892 32823
rect 13956 32759 13982 32823
rect 13790 32743 13982 32759
rect 13854 32679 13892 32743
rect 13956 32679 13982 32743
rect 13790 32663 13982 32679
rect 13854 32599 13892 32663
rect 13956 32599 13982 32663
rect 13790 32583 13982 32599
rect 13854 32519 13892 32583
rect 13956 32519 13982 32583
rect 13790 32503 13982 32519
rect 13854 32439 13892 32503
rect 13956 32439 13982 32503
rect 13790 32423 13982 32439
rect 13854 32359 13892 32423
rect 13956 32359 13982 32423
rect 13790 32343 13982 32359
rect 13854 32279 13892 32343
rect 13956 32279 13982 32343
rect 13790 32263 13982 32279
rect 13854 32199 13892 32263
rect 13956 32199 13982 32263
rect 13790 32183 13982 32199
rect 13854 32119 13892 32183
rect 13956 32119 13982 32183
rect 13790 32103 13982 32119
rect 13854 32039 13892 32103
rect 13956 32039 13982 32103
rect 13790 32023 13982 32039
rect 13854 31959 13892 32023
rect 13956 32018 13982 32023
rect 13977 31962 13982 32018
rect 13956 31959 13982 31962
rect 13790 31943 13982 31959
rect 13854 31879 13892 31943
rect 13956 31936 13982 31943
rect 13977 31880 13982 31936
rect 13956 31879 13982 31880
rect 13790 31863 13982 31879
rect 13854 31799 13892 31863
rect 13956 31854 13982 31863
rect 13790 31798 13795 31799
rect 13851 31798 13921 31799
rect 13977 31798 13982 31854
rect 13790 31783 13982 31798
rect 13854 31719 13892 31783
rect 13956 31772 13982 31783
rect 13790 31716 13795 31719
rect 13851 31716 13921 31719
rect 13977 31716 13982 31772
rect 13790 31703 13982 31716
rect 13854 31639 13892 31703
rect 13956 31690 13982 31703
rect 13790 31634 13795 31639
rect 13851 31634 13921 31639
rect 13977 31634 13982 31690
rect 13790 31623 13982 31634
rect 13854 31559 13892 31623
rect 13956 31608 13982 31623
rect 13790 31552 13795 31559
rect 13851 31552 13921 31559
rect 13977 31552 13982 31608
rect 13790 31543 13982 31552
rect 13854 31479 13892 31543
rect 13956 31526 13982 31543
rect 13790 31470 13795 31479
rect 13851 31470 13921 31479
rect 13977 31470 13982 31526
rect 13790 31463 13982 31470
rect 13854 31399 13892 31463
rect 13956 31444 13982 31463
rect 13790 31388 13795 31399
rect 13851 31388 13921 31399
rect 13977 31388 13982 31444
rect 13790 31383 13982 31388
rect 13854 31319 13892 31383
rect 13956 31362 13982 31383
rect 13790 31306 13795 31319
rect 13851 31306 13921 31319
rect 13977 31306 13982 31362
rect 13790 31303 13982 31306
rect 13854 31239 13892 31303
rect 13956 31280 13982 31303
rect 13790 31224 13795 31239
rect 13851 31224 13921 31239
rect 13977 31224 13982 31280
rect 13790 31223 13982 31224
rect 13854 31159 13892 31223
rect 13956 31198 13982 31223
rect 13790 31143 13795 31159
rect 13851 31143 13921 31159
rect 13854 31079 13892 31143
rect 13977 31142 13982 31198
rect 13956 31116 13982 31142
rect 13790 31063 13795 31079
rect 13851 31063 13921 31079
rect 13854 30999 13892 31063
rect 13977 31060 13982 31116
rect 13956 31034 13982 31060
rect 13790 30983 13795 30999
rect 13851 30983 13921 30999
rect 13854 30919 13892 30983
rect 13977 30978 13982 31034
rect 13956 30952 13982 30978
rect 13790 30903 13795 30919
rect 13851 30903 13921 30919
rect 13854 30839 13892 30903
rect 13977 30896 13982 30952
rect 13956 30870 13982 30896
rect 13790 30822 13795 30839
rect 13851 30822 13921 30839
rect 13854 30758 13892 30822
rect 13977 30814 13982 30870
rect 13956 30788 13982 30814
rect 13790 30741 13795 30758
rect 13851 30741 13921 30758
rect 13854 30677 13892 30741
rect 13977 30732 13982 30788
rect 13956 30706 13982 30732
rect 13790 30660 13795 30677
rect 13851 30660 13921 30677
rect 13854 30596 13892 30660
rect 13977 30650 13982 30706
rect 13956 30624 13982 30650
rect 13790 30579 13795 30596
rect 13851 30579 13921 30596
rect 13854 30515 13892 30579
rect 13977 30568 13982 30624
rect 13956 30542 13982 30568
rect 13790 30498 13795 30515
rect 13851 30498 13921 30515
rect 13854 30434 13892 30498
rect 13977 30486 13982 30542
rect 13956 30460 13982 30486
rect 13790 30417 13795 30434
rect 13851 30417 13921 30434
rect 13854 30353 13892 30417
rect 13977 30404 13982 30460
rect 13956 30378 13982 30404
rect 13790 30336 13795 30353
rect 13851 30336 13921 30353
rect 13854 30272 13892 30336
rect 13977 30322 13982 30378
rect 13956 30296 13982 30322
rect 13790 30255 13795 30272
rect 13851 30255 13921 30272
rect 13854 30191 13892 30255
rect 13977 30240 13982 30296
rect 13956 30214 13982 30240
rect 13790 30174 13795 30191
rect 13851 30174 13921 30191
rect 13854 30110 13892 30174
rect 13977 30158 13982 30214
rect 13956 30132 13982 30158
rect 13790 30093 13795 30110
rect 13851 30093 13921 30110
rect 13854 30029 13892 30093
rect 13977 30076 13982 30132
rect 13956 30050 13982 30076
rect 13790 30012 13795 30029
rect 13851 30012 13921 30029
rect 13854 29948 13892 30012
rect 13977 29994 13982 30050
rect 13956 29968 13982 29994
rect 13790 29931 13795 29948
rect 13851 29931 13921 29948
rect 13854 29867 13892 29931
rect 13977 29912 13982 29968
rect 13956 29886 13982 29912
rect 13790 29850 13795 29867
rect 13851 29850 13921 29867
rect 13854 29786 13892 29850
rect 13977 29830 13982 29886
rect 13956 29804 13982 29830
rect 13790 29769 13795 29786
rect 13851 29769 13921 29786
rect 13854 29705 13892 29769
rect 13977 29748 13982 29804
rect 13956 29722 13982 29748
rect 13790 29688 13795 29705
rect 13851 29688 13921 29705
rect 13854 29624 13892 29688
rect 13977 29666 13982 29722
rect 13956 29640 13982 29666
rect 13790 29607 13795 29624
rect 13851 29607 13921 29624
rect 13854 29543 13892 29607
rect 13977 29584 13982 29640
rect 13956 29558 13982 29584
rect 13790 29526 13795 29543
rect 13851 29526 13921 29543
rect 13854 29462 13892 29526
rect 13977 29502 13982 29558
rect 13956 29476 13982 29502
rect 13790 29445 13795 29462
rect 13851 29445 13921 29462
rect 13854 29381 13892 29445
rect 13977 29420 13982 29476
rect 13956 29381 13982 29420
rect 13790 29364 13982 29381
rect 13854 29300 13892 29364
rect 13956 29300 13982 29364
rect 13790 29283 13982 29300
rect 13854 29219 13892 29283
rect 13956 29219 13982 29283
rect 13790 29202 13982 29219
rect 13854 29138 13892 29202
rect 13956 29138 13982 29202
rect 13790 29121 13982 29138
rect 13854 29057 13892 29121
rect 13956 29057 13982 29121
rect 14253 32761 14672 34764
rect 14253 32705 14259 32761
rect 14315 32705 14347 32761
rect 14403 32705 14435 32761
rect 14491 32705 14523 32761
rect 14579 32705 14611 32761
rect 14667 32705 14672 32761
rect 14253 32681 14672 32705
rect 14253 32625 14259 32681
rect 14315 32625 14347 32681
rect 14403 32625 14435 32681
rect 14491 32625 14523 32681
rect 14579 32625 14611 32681
rect 14667 32625 14672 32681
rect 14253 32601 14672 32625
rect 14253 32545 14259 32601
rect 14315 32545 14347 32601
rect 14403 32545 14435 32601
rect 14491 32545 14523 32601
rect 14579 32545 14611 32601
rect 14667 32545 14672 32601
rect 14253 32521 14672 32545
rect 14253 32465 14259 32521
rect 14315 32465 14347 32521
rect 14403 32465 14435 32521
rect 14491 32465 14523 32521
rect 14579 32465 14611 32521
rect 14667 32465 14672 32521
rect 14253 32441 14672 32465
rect 14253 32385 14259 32441
rect 14315 32385 14347 32441
rect 14403 32385 14435 32441
rect 14491 32385 14523 32441
rect 14579 32385 14611 32441
rect 14667 32385 14672 32441
rect 14253 32361 14672 32385
rect 14253 32305 14259 32361
rect 14315 32305 14347 32361
rect 14403 32305 14435 32361
rect 14491 32305 14523 32361
rect 14579 32305 14611 32361
rect 14667 32305 14672 32361
rect 14253 32281 14672 32305
rect 14253 32225 14259 32281
rect 14315 32225 14347 32281
rect 14403 32225 14435 32281
rect 14491 32225 14523 32281
rect 14579 32225 14611 32281
rect 14667 32225 14672 32281
rect 14253 32201 14672 32225
rect 14253 32145 14259 32201
rect 14315 32145 14347 32201
rect 14403 32145 14435 32201
rect 14491 32145 14523 32201
rect 14579 32145 14611 32201
rect 14667 32145 14672 32201
rect 14253 32121 14672 32145
rect 14253 32065 14259 32121
rect 14315 32065 14347 32121
rect 14403 32065 14435 32121
rect 14491 32065 14523 32121
rect 14579 32065 14611 32121
rect 14667 32065 14672 32121
rect 14253 32041 14672 32065
rect 14253 31985 14259 32041
rect 14315 31985 14347 32041
rect 14403 31985 14435 32041
rect 14491 31985 14523 32041
rect 14579 31985 14611 32041
rect 14667 31985 14672 32041
rect 14253 31961 14672 31985
rect 14253 31905 14259 31961
rect 14315 31905 14347 31961
rect 14403 31905 14435 31961
rect 14491 31905 14523 31961
rect 14579 31905 14611 31961
rect 14667 31905 14672 31961
rect 14253 31881 14672 31905
rect 14253 31825 14259 31881
rect 14315 31825 14347 31881
rect 14403 31825 14435 31881
rect 14491 31825 14523 31881
rect 14579 31825 14611 31881
rect 14667 31825 14672 31881
rect 14253 31801 14672 31825
rect 14253 31745 14259 31801
rect 14315 31745 14347 31801
rect 14403 31745 14435 31801
rect 14491 31745 14523 31801
rect 14579 31745 14611 31801
rect 14667 31745 14672 31801
rect 14253 31721 14672 31745
rect 14253 31665 14259 31721
rect 14315 31665 14347 31721
rect 14403 31665 14435 31721
rect 14491 31665 14523 31721
rect 14579 31665 14611 31721
rect 14667 31665 14672 31721
rect 14253 31641 14672 31665
rect 14253 31585 14259 31641
rect 14315 31585 14347 31641
rect 14403 31585 14435 31641
rect 14491 31585 14523 31641
rect 14579 31585 14611 31641
rect 14667 31585 14672 31641
rect 14253 31561 14672 31585
rect 14253 31505 14259 31561
rect 14315 31505 14347 31561
rect 14403 31505 14435 31561
rect 14491 31505 14523 31561
rect 14579 31505 14611 31561
rect 14667 31505 14672 31561
rect 14253 31481 14672 31505
rect 14253 31425 14259 31481
rect 14315 31425 14347 31481
rect 14403 31425 14435 31481
rect 14491 31425 14523 31481
rect 14579 31425 14611 31481
rect 14667 31425 14672 31481
rect 14253 31400 14672 31425
rect 14253 31344 14259 31400
rect 14315 31344 14347 31400
rect 14403 31344 14435 31400
rect 14491 31344 14523 31400
rect 14579 31344 14611 31400
rect 14667 31344 14672 31400
rect 14253 31319 14672 31344
rect 14253 31263 14259 31319
rect 14315 31263 14347 31319
rect 14403 31263 14435 31319
rect 14491 31263 14523 31319
rect 14579 31263 14611 31319
rect 14667 31263 14672 31319
rect 14253 31238 14672 31263
rect 14253 31182 14259 31238
rect 14315 31182 14347 31238
rect 14403 31182 14435 31238
rect 14491 31182 14523 31238
rect 14579 31182 14611 31238
rect 14667 31182 14672 31238
rect 14253 31157 14672 31182
rect 14253 31101 14259 31157
rect 14315 31101 14347 31157
rect 14403 31101 14435 31157
rect 14491 31101 14523 31157
rect 14579 31101 14611 31157
rect 14667 31101 14672 31157
rect 14253 31076 14672 31101
rect 14253 31020 14259 31076
rect 14315 31020 14347 31076
rect 14403 31020 14435 31076
rect 14491 31020 14523 31076
rect 14579 31020 14611 31076
rect 14667 31020 14672 31076
rect 14253 30995 14672 31020
rect 14253 30939 14259 30995
rect 14315 30939 14347 30995
rect 14403 30939 14435 30995
rect 14491 30939 14523 30995
rect 14579 30939 14611 30995
rect 14667 30939 14672 30995
rect 14253 30914 14672 30939
rect 14253 30858 14259 30914
rect 14315 30858 14347 30914
rect 14403 30858 14435 30914
rect 14491 30858 14523 30914
rect 14579 30858 14611 30914
rect 14667 30858 14672 30914
rect 14253 30833 14672 30858
rect 14253 30777 14259 30833
rect 14315 30777 14347 30833
rect 14403 30777 14435 30833
rect 14491 30777 14523 30833
rect 14579 30777 14611 30833
rect 14667 30777 14672 30833
rect 14253 30752 14672 30777
rect 14253 30696 14259 30752
rect 14315 30696 14347 30752
rect 14403 30696 14435 30752
rect 14491 30696 14523 30752
rect 14579 30696 14611 30752
rect 14667 30696 14672 30752
rect 14253 30671 14672 30696
rect 14253 30615 14259 30671
rect 14315 30615 14347 30671
rect 14403 30615 14435 30671
rect 14491 30615 14523 30671
rect 14579 30615 14611 30671
rect 14667 30615 14672 30671
rect 14253 30590 14672 30615
rect 14253 30534 14259 30590
rect 14315 30534 14347 30590
rect 14403 30534 14435 30590
rect 14491 30534 14523 30590
rect 14579 30534 14611 30590
rect 14667 30534 14672 30590
rect 14253 30509 14672 30534
rect 14253 30453 14259 30509
rect 14315 30453 14347 30509
rect 14403 30453 14435 30509
rect 14491 30453 14523 30509
rect 14579 30453 14611 30509
rect 14667 30453 14672 30509
rect 14253 30428 14672 30453
rect 14253 30372 14259 30428
rect 14315 30372 14347 30428
rect 14403 30372 14435 30428
rect 14491 30372 14523 30428
rect 14579 30372 14611 30428
rect 14667 30372 14672 30428
rect 14253 30347 14672 30372
rect 14253 30291 14259 30347
rect 14315 30291 14347 30347
rect 14403 30291 14435 30347
rect 14491 30291 14523 30347
rect 14579 30291 14611 30347
rect 14667 30291 14672 30347
rect 14253 30266 14672 30291
rect 14253 30210 14259 30266
rect 14315 30210 14347 30266
rect 14403 30210 14435 30266
rect 14491 30210 14523 30266
rect 14579 30210 14611 30266
rect 14667 30210 14672 30266
rect 14253 30185 14672 30210
rect 14253 30129 14259 30185
rect 14315 30129 14347 30185
rect 14403 30129 14435 30185
rect 14491 30129 14523 30185
rect 14579 30129 14611 30185
rect 14667 30129 14672 30185
rect 14253 30104 14672 30129
rect 14253 30048 14259 30104
rect 14315 30048 14347 30104
rect 14403 30048 14435 30104
rect 14491 30048 14523 30104
rect 14579 30048 14611 30104
rect 14667 30048 14672 30104
rect 14253 30023 14672 30048
rect 14253 29967 14259 30023
rect 14315 29967 14347 30023
rect 14403 29967 14435 30023
rect 14491 29967 14523 30023
rect 14579 29967 14611 30023
rect 14667 29967 14672 30023
rect 14253 29942 14672 29967
rect 14253 29886 14259 29942
rect 14315 29886 14347 29942
rect 14403 29886 14435 29942
rect 14491 29886 14523 29942
rect 14579 29886 14611 29942
rect 14667 29886 14672 29942
rect 14253 29861 14672 29886
rect 14253 29805 14259 29861
rect 14315 29805 14347 29861
rect 14403 29805 14435 29861
rect 14491 29805 14523 29861
rect 14579 29805 14611 29861
rect 14667 29805 14672 29861
rect 14253 29780 14672 29805
rect 14253 29724 14259 29780
rect 14315 29724 14347 29780
rect 14403 29724 14435 29780
rect 14491 29724 14523 29780
rect 14579 29724 14611 29780
rect 14667 29724 14672 29780
rect 14253 29699 14672 29724
rect 14253 29643 14259 29699
rect 14315 29643 14347 29699
rect 14403 29643 14435 29699
rect 14491 29643 14523 29699
rect 14579 29643 14611 29699
rect 14667 29643 14672 29699
rect 14253 29618 14672 29643
rect 14253 29562 14259 29618
rect 14315 29562 14347 29618
rect 14403 29562 14435 29618
rect 14491 29562 14523 29618
rect 14579 29562 14611 29618
rect 14667 29562 14672 29618
rect 14253 29537 14672 29562
rect 14253 29481 14259 29537
rect 14315 29481 14347 29537
rect 14403 29481 14435 29537
rect 14491 29481 14523 29537
rect 14579 29481 14611 29537
rect 14667 29481 14672 29537
rect 14253 29456 14672 29481
rect 14253 29400 14259 29456
rect 14315 29400 14347 29456
rect 14403 29400 14435 29456
rect 14491 29400 14523 29456
rect 14579 29400 14611 29456
rect 14667 29400 14672 29456
rect 14253 29375 14672 29400
rect 14253 29319 14259 29375
rect 14315 29319 14347 29375
rect 14403 29319 14435 29375
rect 14491 29319 14523 29375
rect 14579 29319 14611 29375
rect 14667 29319 14672 29375
rect 14253 29294 14672 29319
rect 14253 29238 14259 29294
rect 14315 29238 14347 29294
rect 14403 29238 14435 29294
rect 14491 29238 14523 29294
rect 14579 29238 14611 29294
rect 14667 29238 14672 29294
rect 14253 29213 14672 29238
rect 14253 29157 14259 29213
rect 14315 29157 14347 29213
rect 14403 29157 14435 29213
rect 14491 29157 14523 29213
rect 14579 29157 14611 29213
rect 14667 29157 14672 29213
rect 14253 29132 14672 29157
rect 14253 29076 14259 29132
rect 14315 29076 14347 29132
rect 14403 29076 14435 29132
rect 14491 29076 14523 29132
rect 14579 29076 14611 29132
rect 14667 29076 14672 29132
rect 14253 29065 14672 29076
rect 13790 29040 13982 29057
rect 13854 28976 13892 29040
rect 13956 28976 13982 29040
rect 13790 28959 13982 28976
rect 13854 28895 13892 28959
rect 13956 28895 13982 28959
rect 13790 28878 13982 28895
rect 13854 28814 13892 28878
rect 13956 28814 13982 28878
rect 13790 28797 13982 28814
rect 13854 28733 13892 28797
rect 13956 28733 13982 28797
rect 13790 28716 13982 28733
rect 13854 28652 13892 28716
rect 13956 28652 13982 28716
rect 13790 28635 13982 28652
rect 13854 28571 13892 28635
rect 13956 28571 13982 28635
rect 13790 28554 13982 28571
rect 13854 28490 13892 28554
rect 13956 28490 13982 28554
rect 13790 28473 13982 28490
rect 13854 28409 13892 28473
rect 13956 28409 13982 28473
rect 13790 28392 13982 28409
rect 13854 28328 13892 28392
rect 13956 28328 13982 28392
rect 13790 28311 13982 28328
rect 13854 28247 13892 28311
rect 13956 28247 13982 28311
rect 13790 28230 13982 28247
rect 13854 28166 13892 28230
rect 13956 28166 13982 28230
rect 13790 28149 13982 28166
rect 13854 28085 13892 28149
rect 13956 28085 13982 28149
rect 13790 28068 13982 28085
rect 13854 28004 13892 28068
rect 13956 28004 13982 28068
rect 13790 27987 13982 28004
rect 13854 27923 13892 27987
rect 13956 27923 13982 27987
rect 13790 27906 13982 27923
rect 13854 27842 13892 27906
rect 13956 27842 13982 27906
rect 13790 27825 13982 27842
rect 13854 27761 13892 27825
rect 13956 27761 13982 27825
rect 13790 27744 13982 27761
rect 13854 27680 13892 27744
rect 13956 27680 13982 27744
rect 13790 27663 13982 27680
rect 13854 27599 13892 27663
rect 13956 27599 13982 27663
rect 13790 27582 13982 27599
rect 13854 27518 13892 27582
rect 13956 27518 13982 27582
rect 13790 27501 13982 27518
rect 13854 27437 13892 27501
rect 13956 27437 13982 27501
rect 13790 27420 13982 27437
rect 13854 27356 13892 27420
rect 13956 27401 13982 27420
rect 14167 28577 14784 28633
rect 14167 28521 14283 28577
rect 14339 28521 14381 28577
rect 14437 28521 14479 28577
rect 14535 28521 14577 28577
rect 14633 28521 14784 28577
rect 14167 28497 14784 28521
rect 14167 28441 14283 28497
rect 14339 28441 14381 28497
rect 14437 28441 14479 28497
rect 14535 28441 14577 28497
rect 14633 28441 14784 28497
rect 14167 28417 14784 28441
rect 14167 28361 14283 28417
rect 14339 28361 14381 28417
rect 14437 28361 14479 28417
rect 14535 28361 14577 28417
rect 14633 28361 14784 28417
rect 14167 28337 14784 28361
rect 14167 28281 14283 28337
rect 14339 28281 14381 28337
rect 14437 28281 14479 28337
rect 14535 28281 14577 28337
rect 14633 28281 14784 28337
rect 14167 28257 14784 28281
rect 14167 28201 14283 28257
rect 14339 28201 14381 28257
rect 14437 28201 14479 28257
rect 14535 28201 14577 28257
rect 14633 28201 14784 28257
rect 14167 28177 14784 28201
rect 14167 28121 14283 28177
rect 14339 28121 14381 28177
rect 14437 28121 14479 28177
rect 14535 28121 14577 28177
rect 14633 28121 14784 28177
rect 14167 28097 14784 28121
rect 14167 28041 14283 28097
rect 14339 28041 14381 28097
rect 14437 28041 14479 28097
rect 14535 28041 14577 28097
rect 14633 28041 14784 28097
rect 14167 28017 14784 28041
rect 14167 27961 14283 28017
rect 14339 27961 14381 28017
rect 14437 27961 14479 28017
rect 14535 27961 14577 28017
rect 14633 27961 14784 28017
rect 14167 27937 14784 27961
rect 14167 27881 14283 27937
rect 14339 27881 14381 27937
rect 14437 27881 14479 27937
rect 14535 27881 14577 27937
rect 14633 27881 14784 27937
rect 14167 27857 14784 27881
rect 14167 27801 14283 27857
rect 14339 27801 14381 27857
rect 14437 27801 14479 27857
rect 14535 27801 14577 27857
rect 14633 27801 14784 27857
rect 14167 27777 14784 27801
rect 14167 27721 14283 27777
rect 14339 27721 14381 27777
rect 14437 27721 14479 27777
rect 14535 27721 14577 27777
rect 14633 27721 14784 27777
rect 14167 27697 14784 27721
rect 14167 27641 14283 27697
rect 14339 27641 14381 27697
rect 14437 27641 14479 27697
rect 14535 27641 14577 27697
rect 14633 27641 14784 27697
rect 14167 27617 14784 27641
rect 14167 27561 14283 27617
rect 14339 27561 14381 27617
rect 14437 27561 14479 27617
rect 14535 27561 14577 27617
rect 14633 27561 14784 27617
rect 14167 27537 14784 27561
rect 14167 27481 14283 27537
rect 14339 27481 14381 27537
rect 14437 27481 14479 27537
rect 14535 27481 14577 27537
rect 14633 27481 14784 27537
rect 14167 27457 14784 27481
tri 13982 27401 13997 27416 sw
rect 14167 27401 14283 27457
rect 14339 27401 14381 27457
rect 14437 27401 14479 27457
rect 14535 27401 14577 27457
rect 14633 27401 14784 27457
rect 13956 27377 13997 27401
tri 13997 27377 14021 27401 sw
rect 14167 27377 14784 27401
rect 13956 27356 14021 27377
rect 13790 27355 14021 27356
tri 14021 27355 14043 27377 sw
rect 13790 27347 14043 27355
rect 13790 27339 13974 27347
rect 13854 27275 13892 27339
rect 13956 27283 13974 27339
rect 14038 27283 14043 27347
rect 13956 27275 14043 27283
rect 13790 27262 14043 27275
rect 13790 27258 13974 27262
tri 13788 27241 13790 27243 se
tri 13764 27217 13788 27241 se
rect 13788 27217 13790 27241
tri 13742 27195 13764 27217 se
rect 13764 27195 13790 27217
tri 12990 27161 13024 27195 sw
tri 13708 27161 13742 27195 se
rect 13742 27194 13790 27195
rect 13854 27194 13892 27258
rect 13956 27198 13974 27258
rect 14038 27198 14043 27262
rect 13956 27194 14043 27198
rect 13742 27177 14043 27194
rect 13742 27161 13790 27177
rect 9822 27137 10048 27161
tri 10048 27137 10072 27161 sw
rect 10814 27137 11040 27161
tri 11040 27137 11064 27161 sw
rect 11806 27137 12032 27161
tri 12032 27137 12056 27161 sw
rect 12798 27137 13024 27161
tri 13024 27137 13048 27161 sw
tri 13684 27137 13708 27161 se
rect 13708 27137 13790 27161
rect 9822 27101 10072 27137
tri 10072 27101 10108 27137 sw
rect 9822 26726 10108 27101
tri 9822 26716 9832 26726 ne
rect 9832 26716 10108 26726
rect 10814 27101 11064 27137
tri 11064 27101 11100 27137 sw
rect 10814 26726 11100 27101
tri 10814 26716 10824 26726 ne
rect 10824 26716 11100 26726
rect 11806 27101 12056 27137
tri 12056 27101 12092 27137 sw
rect 11806 26726 12092 27101
tri 11806 26716 11816 26726 ne
rect 11816 26716 12092 26726
rect 12798 27101 13048 27137
tri 13048 27101 13084 27137 sw
tri 13654 27107 13684 27137 se
rect 13684 27113 13790 27137
rect 13854 27113 13892 27177
rect 13956 27176 14043 27177
rect 13956 27113 13974 27176
rect 13684 27112 13974 27113
rect 14038 27112 14043 27176
rect 13684 27107 14043 27112
tri 13653 27106 13654 27107 se
rect 13654 27106 14043 27107
rect 12798 26726 13084 27101
tri 12798 26716 12808 26726 ne
rect 12808 26716 13084 26726
tri 9832 26660 9888 26716 ne
rect 9888 26660 10108 26716
tri 10824 26660 10880 26716 ne
rect 10880 26660 11100 26716
tri 11816 26660 11872 26716 ne
rect 11872 26660 12092 26716
tri 12808 26660 12864 26716 ne
rect 12864 26660 13084 26716
tri 9888 26657 9891 26660 ne
rect 9891 26657 10108 26660
tri 10880 26657 10883 26660 ne
rect 10883 26657 11100 26660
tri 11872 26657 11875 26660 ne
rect 11875 26657 12092 26660
tri 12864 26657 12867 26660 ne
rect 12867 26657 13084 26660
tri 9891 26632 9916 26657 ne
rect 9916 26632 10108 26657
tri 10883 26632 10908 26657 ne
rect 10908 26632 11100 26657
tri 11875 26632 11900 26657 ne
rect 11900 26632 12092 26657
tri 12867 26632 12892 26657 ne
rect 12892 26632 13084 26657
tri 9916 26624 9924 26632 ne
tri 9522 26548 9526 26552 sw
rect 9424 26492 9526 26548
tri 9526 26492 9582 26548 sw
rect 9424 26458 9582 26492
tri 9582 26458 9616 26492 sw
rect 9424 26176 9616 26458
rect 9424 26120 9429 26176
rect 9485 26120 9555 26176
rect 9611 26120 9616 26176
rect 9424 26081 9616 26120
rect 9424 26025 9429 26081
rect 9485 26025 9555 26081
rect 9611 26025 9616 26081
rect 9424 25986 9616 26025
rect 9424 25930 9429 25986
rect 9485 25930 9555 25986
rect 9611 25930 9616 25986
rect 9424 25891 9616 25930
rect 9424 25835 9429 25891
rect 9485 25835 9555 25891
rect 9611 25835 9616 25891
rect 9424 25795 9616 25835
rect 9424 25739 9429 25795
rect 9485 25739 9555 25795
rect 9611 25739 9616 25795
rect 9424 25699 9616 25739
rect 9424 25643 9429 25699
rect 9485 25643 9555 25699
rect 9611 25643 9616 25699
rect 9424 23686 9616 25643
rect 9424 23630 9433 23686
rect 9489 23630 9551 23686
rect 9607 23630 9616 23686
rect 9424 23606 9616 23630
rect 9424 23550 9433 23606
rect 9489 23550 9551 23606
rect 9607 23550 9616 23606
rect 9424 23526 9616 23550
rect 9424 23470 9433 23526
rect 9489 23470 9551 23526
rect 9607 23470 9616 23526
rect 9424 23446 9616 23470
rect 9424 23390 9433 23446
rect 9489 23390 9551 23446
rect 9607 23390 9616 23446
rect 9424 23366 9616 23390
rect 9424 23310 9433 23366
rect 9489 23310 9551 23366
rect 9607 23310 9616 23366
rect 9424 23286 9616 23310
rect 9424 23230 9433 23286
rect 9489 23230 9551 23286
rect 9607 23230 9616 23286
rect 9424 23206 9616 23230
rect 9424 23150 9433 23206
rect 9489 23150 9551 23206
rect 9607 23150 9616 23206
rect 9424 23126 9616 23150
rect 9424 23070 9433 23126
rect 9489 23070 9551 23126
rect 9607 23070 9616 23126
rect 9424 23046 9616 23070
rect 9424 22990 9433 23046
rect 9489 22990 9551 23046
rect 9607 22990 9616 23046
rect 9424 22966 9616 22990
rect 9424 22910 9433 22966
rect 9489 22910 9551 22966
rect 9607 22910 9616 22966
rect 9424 22886 9616 22910
rect 9424 22830 9433 22886
rect 9489 22830 9551 22886
rect 9607 22830 9616 22886
rect 9424 22806 9616 22830
rect 9424 22750 9433 22806
rect 9489 22750 9551 22806
rect 9607 22750 9616 22806
rect 9424 22726 9616 22750
rect 9424 22670 9433 22726
rect 9489 22670 9551 22726
rect 9607 22670 9616 22726
rect 9424 22646 9616 22670
rect 9424 22590 9433 22646
rect 9489 22590 9551 22646
rect 9607 22590 9616 22646
rect 9424 22566 9616 22590
rect 9424 22510 9433 22566
rect 9489 22510 9551 22566
rect 9607 22510 9616 22566
rect 9424 22486 9616 22510
rect 9424 22430 9433 22486
rect 9489 22430 9551 22486
rect 9607 22430 9616 22486
rect 9424 22406 9616 22430
rect 9424 22350 9433 22406
rect 9489 22350 9551 22406
rect 9607 22350 9616 22406
rect 9424 22326 9616 22350
rect 9424 22270 9433 22326
rect 9489 22270 9551 22326
rect 9607 22270 9616 22326
rect 9424 22245 9616 22270
rect 9424 22189 9433 22245
rect 9489 22189 9551 22245
rect 9607 22189 9616 22245
rect 9424 22164 9616 22189
rect 9424 22108 9433 22164
rect 9489 22108 9551 22164
rect 9607 22108 9616 22164
rect 9424 22083 9616 22108
rect 9424 22027 9433 22083
rect 9489 22027 9551 22083
rect 9607 22027 9616 22083
rect 9424 22002 9616 22027
rect 9424 21946 9433 22002
rect 9489 21946 9551 22002
rect 9607 21946 9616 22002
rect 9424 21921 9616 21946
rect 9424 21865 9433 21921
rect 9489 21865 9551 21921
rect 9607 21865 9616 21921
rect 9424 21840 9616 21865
rect 9424 21784 9433 21840
rect 9489 21784 9551 21840
rect 9607 21784 9616 21840
rect 9424 21759 9616 21784
rect 9424 21703 9433 21759
rect 9489 21703 9551 21759
rect 9607 21703 9616 21759
rect 9424 21678 9616 21703
rect 9424 21622 9433 21678
rect 9489 21622 9551 21678
rect 9607 21622 9616 21678
rect 9424 21597 9616 21622
rect 9424 21541 9433 21597
rect 9489 21541 9551 21597
rect 9607 21541 9616 21597
rect 9424 21516 9616 21541
rect 9424 21460 9433 21516
rect 9489 21460 9551 21516
rect 9607 21460 9616 21516
rect 9424 21435 9616 21460
rect 9424 21379 9433 21435
rect 9489 21379 9551 21435
rect 9607 21379 9616 21435
rect 9424 21354 9616 21379
rect 9424 21298 9433 21354
rect 9489 21298 9551 21354
rect 9607 21298 9616 21354
rect 9424 21273 9616 21298
rect 9424 21217 9433 21273
rect 9489 21217 9551 21273
rect 9607 21217 9616 21273
rect 9424 21192 9616 21217
rect 9424 21136 9433 21192
rect 9489 21136 9551 21192
rect 9607 21136 9616 21192
rect 8496 18528 8560 18592
rect 8432 18512 8624 18528
rect 8496 18448 8560 18512
rect 8432 18432 8624 18448
rect 8496 18368 8560 18432
rect 8432 18352 8624 18368
rect 8496 18288 8560 18352
rect 8432 18272 8624 18288
rect 8496 18208 8560 18272
rect 8432 18192 8624 18208
rect 8496 18128 8560 18192
rect 8432 18112 8624 18128
rect 8496 18048 8560 18112
rect 8432 18032 8624 18048
rect 8496 17968 8560 18032
rect 8432 17952 8624 17968
rect 8496 17888 8560 17952
rect 8432 17872 8624 17888
rect 8496 17808 8560 17872
rect 8432 17792 8624 17808
rect 8496 17728 8560 17792
rect 8432 17712 8624 17728
rect 8496 17648 8560 17712
rect 8432 17632 8624 17648
rect 8496 17568 8560 17632
rect 8432 17552 8624 17568
rect 8496 17488 8560 17552
rect 8432 17472 8624 17488
rect 8496 17408 8560 17472
rect 8432 17392 8624 17408
rect 8496 17328 8560 17392
rect 8432 17312 8624 17328
rect 8496 17248 8560 17312
rect 8432 17232 8624 17248
rect 8496 17168 8560 17232
rect 8432 17152 8624 17168
rect 8496 17088 8560 17152
rect 8432 17072 8624 17088
rect 8496 17008 8560 17072
rect 8432 16992 8624 17008
rect 8496 16928 8560 16992
rect 8432 16912 8624 16928
rect 8496 16848 8560 16912
rect 8432 16832 8624 16848
rect 8496 16768 8560 16832
rect 8432 16752 8624 16768
rect 8496 16688 8560 16752
rect 8432 16672 8624 16688
rect 8496 16608 8560 16672
rect 8432 16592 8624 16608
rect 8496 16528 8560 16592
rect 8432 16512 8624 16528
rect 8496 16448 8560 16512
rect 8432 16432 8624 16448
rect 8496 16368 8560 16432
rect 8432 16351 8624 16368
rect 8496 16287 8560 16351
rect 8432 16270 8624 16287
rect 8496 16206 8560 16270
rect 8432 16189 8624 16206
rect 8496 16125 8560 16189
rect 8432 16108 8624 16125
rect 8496 16044 8560 16108
rect 8432 16027 8624 16044
rect 8496 15963 8560 16027
rect 8432 15946 8624 15963
rect 8496 15882 8560 15946
rect 8432 15865 8624 15882
rect 8496 15801 8560 15865
rect 8432 15784 8624 15801
rect 8496 15720 8560 15784
rect 8432 15703 8624 15720
rect 8496 15639 8560 15703
rect 8432 15622 8624 15639
rect 8496 15558 8560 15622
rect 8432 15541 8624 15558
rect 8496 15477 8560 15541
rect 8432 15460 8624 15477
rect 8496 15396 8560 15460
rect 8432 15379 8624 15396
rect 8496 15315 8560 15379
rect 8432 15298 8624 15315
rect 8496 15234 8560 15298
rect 8432 15217 8624 15234
rect 8496 15153 8560 15217
rect 8432 15136 8624 15153
rect 8496 15072 8560 15136
rect 8432 15055 8624 15072
rect 8496 14991 8560 15055
rect 8432 14974 8624 14991
rect 8496 14910 8560 14974
rect 8432 14893 8624 14910
rect 8496 14829 8560 14893
rect 8432 14812 8624 14829
rect 8496 14748 8560 14812
rect 8432 14731 8624 14748
rect 8496 14667 8560 14731
rect 8432 14650 8624 14667
rect 8496 14586 8560 14650
rect 8432 14569 8624 14586
rect 8496 14505 8560 14569
rect 8432 14488 8624 14505
rect 8496 14424 8560 14488
rect 8432 14407 8624 14424
rect 8496 14343 8560 14407
rect 8432 14326 8624 14343
rect 8496 14262 8560 14326
rect 8432 14245 8624 14262
rect 8496 14181 8560 14245
rect 8432 14164 8624 14181
rect 8496 14100 8560 14164
rect 8432 14083 8624 14100
rect 8496 14019 8560 14083
rect 8432 14002 8624 14019
rect 8496 13938 8560 14002
rect 8432 13921 8624 13938
rect 8496 13857 8560 13921
rect 8432 13840 8624 13857
rect 8496 13776 8560 13840
rect 8432 13759 8624 13776
rect 8496 13695 8560 13759
rect 8432 13678 8624 13695
rect 8496 13614 8560 13678
rect 8432 13607 8624 13614
rect 9424 18592 9616 21136
rect 9924 23686 10108 26632
tri 10908 26624 10916 26632 ne
rect 9924 23630 9929 23686
rect 9985 23630 10047 23686
rect 10103 23630 10108 23686
rect 9924 23606 10108 23630
rect 9924 23550 9929 23606
rect 9985 23550 10047 23606
rect 10103 23550 10108 23606
rect 9924 23526 10108 23550
rect 9924 23470 9929 23526
rect 9985 23470 10047 23526
rect 10103 23470 10108 23526
rect 9924 23446 10108 23470
rect 9924 23390 9929 23446
rect 9985 23390 10047 23446
rect 10103 23390 10108 23446
rect 9924 23366 10108 23390
rect 9924 23310 9929 23366
rect 9985 23310 10047 23366
rect 10103 23310 10108 23366
rect 9924 23286 10108 23310
rect 9924 23230 9929 23286
rect 9985 23230 10047 23286
rect 10103 23230 10108 23286
rect 9924 23206 10108 23230
rect 9924 23150 9929 23206
rect 9985 23150 10047 23206
rect 10103 23150 10108 23206
rect 9924 23126 10108 23150
rect 9924 23070 9929 23126
rect 9985 23070 10047 23126
rect 10103 23070 10108 23126
rect 9924 23046 10108 23070
rect 9924 22990 9929 23046
rect 9985 22990 10047 23046
rect 10103 22990 10108 23046
rect 9924 22966 10108 22990
rect 9924 22910 9929 22966
rect 9985 22910 10047 22966
rect 10103 22910 10108 22966
rect 9924 22886 10108 22910
rect 9924 22830 9929 22886
rect 9985 22830 10047 22886
rect 10103 22830 10108 22886
rect 9924 22806 10108 22830
rect 9924 22750 9929 22806
rect 9985 22750 10047 22806
rect 10103 22750 10108 22806
rect 9924 22726 10108 22750
rect 9924 22670 9929 22726
rect 9985 22670 10047 22726
rect 10103 22670 10108 22726
rect 9924 22646 10108 22670
rect 9924 22590 9929 22646
rect 9985 22590 10047 22646
rect 10103 22590 10108 22646
rect 9924 22566 10108 22590
rect 9924 22510 9929 22566
rect 9985 22510 10047 22566
rect 10103 22510 10108 22566
rect 9924 22486 10108 22510
rect 9924 22430 9929 22486
rect 9985 22430 10047 22486
rect 10103 22430 10108 22486
rect 9924 22406 10108 22430
rect 9924 22350 9929 22406
rect 9985 22350 10047 22406
rect 10103 22350 10108 22406
rect 9924 22326 10108 22350
rect 9924 22270 9929 22326
rect 9985 22270 10047 22326
rect 10103 22270 10108 22326
rect 9924 22245 10108 22270
rect 9924 22189 9929 22245
rect 9985 22189 10047 22245
rect 10103 22189 10108 22245
rect 9924 22164 10108 22189
rect 9924 22108 9929 22164
rect 9985 22108 10047 22164
rect 10103 22108 10108 22164
rect 9924 22083 10108 22108
rect 9924 22027 9929 22083
rect 9985 22027 10047 22083
rect 10103 22027 10108 22083
rect 9924 22002 10108 22027
rect 9924 21946 9929 22002
rect 9985 21946 10047 22002
rect 10103 21946 10108 22002
rect 9924 21921 10108 21946
rect 9924 21865 9929 21921
rect 9985 21865 10047 21921
rect 10103 21865 10108 21921
rect 9924 21840 10108 21865
rect 9924 21784 9929 21840
rect 9985 21784 10047 21840
rect 10103 21784 10108 21840
rect 9924 21759 10108 21784
rect 9924 21703 9929 21759
rect 9985 21703 10047 21759
rect 10103 21703 10108 21759
rect 9924 21678 10108 21703
rect 9924 21622 9929 21678
rect 9985 21622 10047 21678
rect 10103 21622 10108 21678
rect 9924 21597 10108 21622
rect 9924 21541 9929 21597
rect 9985 21541 10047 21597
rect 10103 21541 10108 21597
rect 9924 21516 10108 21541
rect 9924 21460 9929 21516
rect 9985 21460 10047 21516
rect 10103 21460 10108 21516
rect 9924 21435 10108 21460
rect 9924 21379 9929 21435
rect 9985 21379 10047 21435
rect 10103 21379 10108 21435
rect 9924 21354 10108 21379
rect 9924 21298 9929 21354
rect 9985 21298 10047 21354
rect 10103 21298 10108 21354
rect 9924 21273 10108 21298
rect 9924 21217 9929 21273
rect 9985 21217 10047 21273
rect 10103 21217 10108 21273
rect 9924 21192 10108 21217
rect 9924 21136 9929 21192
rect 9985 21136 10047 21192
rect 10103 21136 10108 21192
rect 9924 19673 10108 21136
rect 9988 19609 10044 19673
rect 9924 19581 10108 19609
rect 9988 19517 10044 19581
rect 9924 19489 10108 19517
rect 9988 19425 10044 19489
rect 9924 19397 10108 19425
rect 9988 19333 10044 19397
rect 9924 19305 10108 19333
rect 9988 19241 10044 19305
rect 9924 19212 10108 19241
rect 9988 19148 10044 19212
rect 9924 19139 10108 19148
rect 10416 23686 10608 23721
rect 10416 23630 10425 23686
rect 10481 23630 10543 23686
rect 10599 23630 10608 23686
rect 10416 23606 10608 23630
rect 10416 23550 10425 23606
rect 10481 23550 10543 23606
rect 10599 23550 10608 23606
rect 10416 23526 10608 23550
rect 10416 23470 10425 23526
rect 10481 23470 10543 23526
rect 10599 23470 10608 23526
rect 10416 23446 10608 23470
rect 10416 23390 10425 23446
rect 10481 23390 10543 23446
rect 10599 23390 10608 23446
rect 10416 23366 10608 23390
rect 10416 23310 10425 23366
rect 10481 23310 10543 23366
rect 10599 23310 10608 23366
rect 10416 23286 10608 23310
rect 10416 23230 10425 23286
rect 10481 23230 10543 23286
rect 10599 23230 10608 23286
rect 10416 23206 10608 23230
rect 10416 23150 10425 23206
rect 10481 23150 10543 23206
rect 10599 23150 10608 23206
rect 10416 23126 10608 23150
rect 10416 23070 10425 23126
rect 10481 23070 10543 23126
rect 10599 23070 10608 23126
rect 10416 23046 10608 23070
rect 10416 22990 10425 23046
rect 10481 22990 10543 23046
rect 10599 22990 10608 23046
rect 10416 22966 10608 22990
rect 10416 22910 10425 22966
rect 10481 22910 10543 22966
rect 10599 22910 10608 22966
rect 10416 22886 10608 22910
rect 10416 22830 10425 22886
rect 10481 22830 10543 22886
rect 10599 22830 10608 22886
rect 10416 22806 10608 22830
rect 10416 22750 10425 22806
rect 10481 22750 10543 22806
rect 10599 22750 10608 22806
rect 10416 22726 10608 22750
rect 10416 22670 10425 22726
rect 10481 22670 10543 22726
rect 10599 22670 10608 22726
rect 10416 22646 10608 22670
rect 10416 22590 10425 22646
rect 10481 22590 10543 22646
rect 10599 22590 10608 22646
rect 10416 22566 10608 22590
rect 10416 22510 10425 22566
rect 10481 22510 10543 22566
rect 10599 22510 10608 22566
rect 10416 22486 10608 22510
rect 10416 22430 10425 22486
rect 10481 22430 10543 22486
rect 10599 22430 10608 22486
rect 10416 22406 10608 22430
rect 10416 22350 10425 22406
rect 10481 22350 10543 22406
rect 10599 22350 10608 22406
rect 10416 22326 10608 22350
rect 10416 22270 10425 22326
rect 10481 22270 10543 22326
rect 10599 22270 10608 22326
rect 10416 22245 10608 22270
rect 10416 22189 10425 22245
rect 10481 22189 10543 22245
rect 10599 22189 10608 22245
rect 10416 22164 10608 22189
rect 10416 22108 10425 22164
rect 10481 22108 10543 22164
rect 10599 22108 10608 22164
rect 10416 22083 10608 22108
rect 10416 22027 10425 22083
rect 10481 22027 10543 22083
rect 10599 22027 10608 22083
rect 10416 22002 10608 22027
rect 10416 21946 10425 22002
rect 10481 21946 10543 22002
rect 10599 21946 10608 22002
rect 10416 21921 10608 21946
rect 10416 21865 10425 21921
rect 10481 21865 10543 21921
rect 10599 21865 10608 21921
rect 10416 21840 10608 21865
rect 10416 21784 10425 21840
rect 10481 21784 10543 21840
rect 10599 21784 10608 21840
rect 10416 21759 10608 21784
rect 10416 21703 10425 21759
rect 10481 21703 10543 21759
rect 10599 21703 10608 21759
rect 10416 21678 10608 21703
rect 10416 21622 10425 21678
rect 10481 21622 10543 21678
rect 10599 21622 10608 21678
rect 10416 21597 10608 21622
rect 10416 21541 10425 21597
rect 10481 21541 10543 21597
rect 10599 21541 10608 21597
rect 10416 21516 10608 21541
rect 10416 21460 10425 21516
rect 10481 21460 10543 21516
rect 10599 21460 10608 21516
rect 10416 21435 10608 21460
rect 10416 21379 10425 21435
rect 10481 21379 10543 21435
rect 10599 21379 10608 21435
rect 10416 21354 10608 21379
rect 10416 21298 10425 21354
rect 10481 21298 10543 21354
rect 10599 21298 10608 21354
rect 10416 21273 10608 21298
rect 10416 21217 10425 21273
rect 10481 21217 10543 21273
rect 10599 21217 10608 21273
rect 10416 21192 10608 21217
rect 10416 21136 10425 21192
rect 10481 21136 10543 21192
rect 10599 21136 10608 21192
rect 9488 18528 9552 18592
rect 9424 18512 9616 18528
rect 9488 18448 9552 18512
rect 9424 18432 9616 18448
rect 9488 18368 9552 18432
rect 9424 18352 9616 18368
rect 9488 18288 9552 18352
rect 9424 18272 9616 18288
rect 9488 18208 9552 18272
rect 9424 18192 9616 18208
rect 9488 18128 9552 18192
rect 9424 18112 9616 18128
rect 9488 18048 9552 18112
rect 9424 18032 9616 18048
rect 9488 17968 9552 18032
rect 9424 17952 9616 17968
rect 9488 17888 9552 17952
rect 9424 17872 9616 17888
rect 9488 17808 9552 17872
rect 9424 17792 9616 17808
rect 9488 17728 9552 17792
rect 9424 17712 9616 17728
rect 9488 17648 9552 17712
rect 9424 17632 9616 17648
rect 9488 17568 9552 17632
rect 9424 17552 9616 17568
rect 9488 17488 9552 17552
rect 9424 17472 9616 17488
rect 9488 17408 9552 17472
rect 9424 17392 9616 17408
rect 9488 17328 9552 17392
rect 9424 17312 9616 17328
rect 9488 17248 9552 17312
rect 9424 17232 9616 17248
rect 9488 17168 9552 17232
rect 9424 17152 9616 17168
rect 9488 17088 9552 17152
rect 9424 17072 9616 17088
rect 9488 17008 9552 17072
rect 9424 16992 9616 17008
rect 9488 16928 9552 16992
rect 9424 16912 9616 16928
rect 9488 16848 9552 16912
rect 9424 16832 9616 16848
rect 9488 16768 9552 16832
rect 9424 16752 9616 16768
rect 9488 16688 9552 16752
rect 9424 16672 9616 16688
rect 9488 16608 9552 16672
rect 9424 16592 9616 16608
rect 9488 16528 9552 16592
rect 9424 16512 9616 16528
rect 9488 16448 9552 16512
rect 9424 16432 9616 16448
rect 9488 16368 9552 16432
rect 9424 16351 9616 16368
rect 9488 16287 9552 16351
rect 9424 16270 9616 16287
rect 9488 16206 9552 16270
rect 9424 16189 9616 16206
rect 9488 16125 9552 16189
rect 9424 16108 9616 16125
rect 9488 16044 9552 16108
rect 9424 16027 9616 16044
rect 9488 15963 9552 16027
rect 9424 15946 9616 15963
rect 9488 15882 9552 15946
rect 9424 15865 9616 15882
rect 9488 15801 9552 15865
rect 9424 15784 9616 15801
rect 9488 15720 9552 15784
rect 9424 15703 9616 15720
rect 9488 15639 9552 15703
rect 9424 15622 9616 15639
rect 9488 15558 9552 15622
rect 9424 15541 9616 15558
rect 9488 15477 9552 15541
rect 9424 15460 9616 15477
rect 9488 15396 9552 15460
rect 9424 15379 9616 15396
rect 9488 15315 9552 15379
rect 9424 15298 9616 15315
rect 9488 15234 9552 15298
rect 9424 15217 9616 15234
rect 9488 15153 9552 15217
rect 9424 15136 9616 15153
rect 9488 15072 9552 15136
rect 9424 15055 9616 15072
rect 9488 14991 9552 15055
rect 9424 14974 9616 14991
rect 9488 14910 9552 14974
rect 9424 14893 9616 14910
rect 9488 14829 9552 14893
rect 9424 14812 9616 14829
rect 9488 14748 9552 14812
rect 9424 14731 9616 14748
rect 9488 14667 9552 14731
rect 9424 14650 9616 14667
rect 9488 14586 9552 14650
rect 9424 14569 9616 14586
rect 9488 14505 9552 14569
rect 9424 14488 9616 14505
rect 9488 14424 9552 14488
rect 9424 14407 9616 14424
rect 9488 14343 9552 14407
rect 9424 14326 9616 14343
rect 9488 14262 9552 14326
rect 9424 14245 9616 14262
rect 9488 14181 9552 14245
rect 9424 14164 9616 14181
rect 9488 14100 9552 14164
rect 9424 14083 9616 14100
rect 9488 14019 9552 14083
rect 9424 14002 9616 14019
rect 9488 13938 9552 14002
rect 9424 13921 9616 13938
rect 9488 13857 9552 13921
rect 9424 13840 9616 13857
rect 9488 13776 9552 13840
rect 9424 13759 9616 13776
rect 9488 13695 9552 13759
rect 9424 13678 9616 13695
rect 9488 13614 9552 13678
rect 9424 13607 9616 13614
rect 10416 18592 10608 21136
rect 10916 23686 11100 26632
tri 11900 26624 11908 26632 ne
rect 10916 23630 10921 23686
rect 10977 23630 11039 23686
rect 11095 23630 11100 23686
rect 10916 23606 11100 23630
rect 10916 23550 10921 23606
rect 10977 23550 11039 23606
rect 11095 23550 11100 23606
rect 10916 23526 11100 23550
rect 10916 23470 10921 23526
rect 10977 23470 11039 23526
rect 11095 23470 11100 23526
rect 10916 23446 11100 23470
rect 10916 23390 10921 23446
rect 10977 23390 11039 23446
rect 11095 23390 11100 23446
rect 10916 23366 11100 23390
rect 10916 23310 10921 23366
rect 10977 23310 11039 23366
rect 11095 23310 11100 23366
rect 10916 23286 11100 23310
rect 10916 23230 10921 23286
rect 10977 23230 11039 23286
rect 11095 23230 11100 23286
rect 10916 23206 11100 23230
rect 10916 23150 10921 23206
rect 10977 23150 11039 23206
rect 11095 23150 11100 23206
rect 10916 23126 11100 23150
rect 10916 23070 10921 23126
rect 10977 23070 11039 23126
rect 11095 23070 11100 23126
rect 10916 23046 11100 23070
rect 10916 22990 10921 23046
rect 10977 22990 11039 23046
rect 11095 22990 11100 23046
rect 10916 22966 11100 22990
rect 10916 22910 10921 22966
rect 10977 22910 11039 22966
rect 11095 22910 11100 22966
rect 10916 22886 11100 22910
rect 10916 22830 10921 22886
rect 10977 22830 11039 22886
rect 11095 22830 11100 22886
rect 10916 22806 11100 22830
rect 10916 22750 10921 22806
rect 10977 22750 11039 22806
rect 11095 22750 11100 22806
rect 10916 22726 11100 22750
rect 10916 22670 10921 22726
rect 10977 22670 11039 22726
rect 11095 22670 11100 22726
rect 10916 22646 11100 22670
rect 10916 22590 10921 22646
rect 10977 22590 11039 22646
rect 11095 22590 11100 22646
rect 10916 22566 11100 22590
rect 10916 22510 10921 22566
rect 10977 22510 11039 22566
rect 11095 22510 11100 22566
rect 10916 22486 11100 22510
rect 10916 22430 10921 22486
rect 10977 22430 11039 22486
rect 11095 22430 11100 22486
rect 10916 22406 11100 22430
rect 10916 22350 10921 22406
rect 10977 22350 11039 22406
rect 11095 22350 11100 22406
rect 10916 22326 11100 22350
rect 10916 22270 10921 22326
rect 10977 22270 11039 22326
rect 11095 22270 11100 22326
rect 10916 22245 11100 22270
rect 10916 22189 10921 22245
rect 10977 22189 11039 22245
rect 11095 22189 11100 22245
rect 10916 22164 11100 22189
rect 10916 22108 10921 22164
rect 10977 22108 11039 22164
rect 11095 22108 11100 22164
rect 10916 22083 11100 22108
rect 10916 22027 10921 22083
rect 10977 22027 11039 22083
rect 11095 22027 11100 22083
rect 10916 22002 11100 22027
rect 10916 21946 10921 22002
rect 10977 21946 11039 22002
rect 11095 21946 11100 22002
rect 10916 21921 11100 21946
rect 10916 21865 10921 21921
rect 10977 21865 11039 21921
rect 11095 21865 11100 21921
rect 10916 21840 11100 21865
rect 10916 21784 10921 21840
rect 10977 21784 11039 21840
rect 11095 21784 11100 21840
rect 10916 21759 11100 21784
rect 10916 21703 10921 21759
rect 10977 21703 11039 21759
rect 11095 21703 11100 21759
rect 10916 21678 11100 21703
rect 10916 21622 10921 21678
rect 10977 21622 11039 21678
rect 11095 21622 11100 21678
rect 10916 21597 11100 21622
rect 10916 21541 10921 21597
rect 10977 21541 11039 21597
rect 11095 21541 11100 21597
rect 10916 21516 11100 21541
rect 10916 21460 10921 21516
rect 10977 21460 11039 21516
rect 11095 21460 11100 21516
rect 10916 21435 11100 21460
rect 10916 21379 10921 21435
rect 10977 21379 11039 21435
rect 11095 21379 11100 21435
rect 10916 21354 11100 21379
rect 10916 21298 10921 21354
rect 10977 21298 11039 21354
rect 11095 21298 11100 21354
rect 10916 21273 11100 21298
rect 10916 21217 10921 21273
rect 10977 21217 11039 21273
rect 11095 21217 11100 21273
rect 10916 21192 11100 21217
rect 10916 21136 10921 21192
rect 10977 21136 11039 21192
rect 11095 21136 11100 21192
rect 10916 19673 11100 21136
rect 10980 19609 11036 19673
rect 10916 19581 11100 19609
rect 10980 19517 11036 19581
rect 10916 19489 11100 19517
rect 10980 19425 11036 19489
rect 10916 19397 11100 19425
rect 10980 19333 11036 19397
rect 10916 19305 11100 19333
rect 10980 19241 11036 19305
rect 10916 19212 11100 19241
rect 10980 19148 11036 19212
rect 10916 19139 11100 19148
rect 11408 23686 11600 23721
rect 11408 23630 11417 23686
rect 11473 23630 11535 23686
rect 11591 23630 11600 23686
rect 11408 23606 11600 23630
rect 11408 23550 11417 23606
rect 11473 23550 11535 23606
rect 11591 23550 11600 23606
rect 11408 23526 11600 23550
rect 11408 23470 11417 23526
rect 11473 23470 11535 23526
rect 11591 23470 11600 23526
rect 11408 23446 11600 23470
rect 11408 23390 11417 23446
rect 11473 23390 11535 23446
rect 11591 23390 11600 23446
rect 11408 23366 11600 23390
rect 11408 23310 11417 23366
rect 11473 23310 11535 23366
rect 11591 23310 11600 23366
rect 11408 23286 11600 23310
rect 11408 23230 11417 23286
rect 11473 23230 11535 23286
rect 11591 23230 11600 23286
rect 11408 23206 11600 23230
rect 11408 23150 11417 23206
rect 11473 23150 11535 23206
rect 11591 23150 11600 23206
rect 11408 23126 11600 23150
rect 11408 23070 11417 23126
rect 11473 23070 11535 23126
rect 11591 23070 11600 23126
rect 11408 23046 11600 23070
rect 11408 22990 11417 23046
rect 11473 22990 11535 23046
rect 11591 22990 11600 23046
rect 11408 22966 11600 22990
rect 11408 22910 11417 22966
rect 11473 22910 11535 22966
rect 11591 22910 11600 22966
rect 11408 22886 11600 22910
rect 11408 22830 11417 22886
rect 11473 22830 11535 22886
rect 11591 22830 11600 22886
rect 11408 22806 11600 22830
rect 11408 22750 11417 22806
rect 11473 22750 11535 22806
rect 11591 22750 11600 22806
rect 11408 22726 11600 22750
rect 11408 22670 11417 22726
rect 11473 22670 11535 22726
rect 11591 22670 11600 22726
rect 11408 22646 11600 22670
rect 11408 22590 11417 22646
rect 11473 22590 11535 22646
rect 11591 22590 11600 22646
rect 11408 22566 11600 22590
rect 11408 22510 11417 22566
rect 11473 22510 11535 22566
rect 11591 22510 11600 22566
rect 11408 22486 11600 22510
rect 11408 22430 11417 22486
rect 11473 22430 11535 22486
rect 11591 22430 11600 22486
rect 11408 22406 11600 22430
rect 11408 22350 11417 22406
rect 11473 22350 11535 22406
rect 11591 22350 11600 22406
rect 11408 22326 11600 22350
rect 11408 22270 11417 22326
rect 11473 22270 11535 22326
rect 11591 22270 11600 22326
rect 11408 22245 11600 22270
rect 11408 22189 11417 22245
rect 11473 22189 11535 22245
rect 11591 22189 11600 22245
rect 11408 22164 11600 22189
rect 11408 22108 11417 22164
rect 11473 22108 11535 22164
rect 11591 22108 11600 22164
rect 11408 22083 11600 22108
rect 11408 22027 11417 22083
rect 11473 22027 11535 22083
rect 11591 22027 11600 22083
rect 11408 22002 11600 22027
rect 11408 21946 11417 22002
rect 11473 21946 11535 22002
rect 11591 21946 11600 22002
rect 11408 21921 11600 21946
rect 11408 21865 11417 21921
rect 11473 21865 11535 21921
rect 11591 21865 11600 21921
rect 11408 21840 11600 21865
rect 11408 21784 11417 21840
rect 11473 21784 11535 21840
rect 11591 21784 11600 21840
rect 11408 21759 11600 21784
rect 11408 21703 11417 21759
rect 11473 21703 11535 21759
rect 11591 21703 11600 21759
rect 11408 21678 11600 21703
rect 11408 21622 11417 21678
rect 11473 21622 11535 21678
rect 11591 21622 11600 21678
rect 11408 21597 11600 21622
rect 11408 21541 11417 21597
rect 11473 21541 11535 21597
rect 11591 21541 11600 21597
rect 11408 21516 11600 21541
rect 11408 21460 11417 21516
rect 11473 21460 11535 21516
rect 11591 21460 11600 21516
rect 11408 21435 11600 21460
rect 11408 21379 11417 21435
rect 11473 21379 11535 21435
rect 11591 21379 11600 21435
rect 11408 21354 11600 21379
rect 11408 21298 11417 21354
rect 11473 21298 11535 21354
rect 11591 21298 11600 21354
rect 11408 21273 11600 21298
rect 11408 21217 11417 21273
rect 11473 21217 11535 21273
rect 11591 21217 11600 21273
rect 11408 21192 11600 21217
rect 11408 21136 11417 21192
rect 11473 21136 11535 21192
rect 11591 21136 11600 21192
rect 10480 18528 10544 18592
rect 10416 18512 10608 18528
rect 10480 18448 10544 18512
rect 10416 18432 10608 18448
rect 10480 18368 10544 18432
rect 10416 18352 10608 18368
rect 10480 18288 10544 18352
rect 10416 18272 10608 18288
rect 10480 18208 10544 18272
rect 10416 18192 10608 18208
rect 10480 18128 10544 18192
rect 10416 18112 10608 18128
rect 10480 18048 10544 18112
rect 10416 18032 10608 18048
rect 10480 17968 10544 18032
rect 10416 17952 10608 17968
rect 10480 17888 10544 17952
rect 10416 17872 10608 17888
rect 10480 17808 10544 17872
rect 10416 17792 10608 17808
rect 10480 17728 10544 17792
rect 10416 17712 10608 17728
rect 10480 17648 10544 17712
rect 10416 17632 10608 17648
rect 10480 17568 10544 17632
rect 10416 17552 10608 17568
rect 10480 17488 10544 17552
rect 10416 17472 10608 17488
rect 10480 17408 10544 17472
rect 10416 17392 10608 17408
rect 10480 17328 10544 17392
rect 10416 17312 10608 17328
rect 10480 17248 10544 17312
rect 10416 17232 10608 17248
rect 10480 17168 10544 17232
rect 10416 17152 10608 17168
rect 10480 17088 10544 17152
rect 10416 17072 10608 17088
rect 10480 17008 10544 17072
rect 10416 16992 10608 17008
rect 10480 16928 10544 16992
rect 10416 16912 10608 16928
rect 10480 16848 10544 16912
rect 10416 16832 10608 16848
rect 10480 16768 10544 16832
rect 10416 16752 10608 16768
rect 10480 16688 10544 16752
rect 10416 16672 10608 16688
rect 10480 16608 10544 16672
rect 10416 16592 10608 16608
rect 10480 16528 10544 16592
rect 10416 16512 10608 16528
rect 10480 16448 10544 16512
rect 10416 16432 10608 16448
rect 10480 16368 10544 16432
rect 10416 16351 10608 16368
rect 10480 16287 10544 16351
rect 10416 16270 10608 16287
rect 10480 16206 10544 16270
rect 10416 16189 10608 16206
rect 10480 16125 10544 16189
rect 10416 16108 10608 16125
rect 10480 16044 10544 16108
rect 10416 16027 10608 16044
rect 10480 15963 10544 16027
rect 10416 15946 10608 15963
rect 10480 15882 10544 15946
rect 10416 15865 10608 15882
rect 10480 15801 10544 15865
rect 10416 15784 10608 15801
rect 10480 15720 10544 15784
rect 10416 15703 10608 15720
rect 10480 15639 10544 15703
rect 10416 15622 10608 15639
rect 10480 15558 10544 15622
rect 10416 15541 10608 15558
rect 10480 15477 10544 15541
rect 10416 15460 10608 15477
rect 10480 15396 10544 15460
rect 10416 15379 10608 15396
rect 10480 15315 10544 15379
rect 10416 15298 10608 15315
rect 10480 15234 10544 15298
rect 10416 15217 10608 15234
rect 10480 15153 10544 15217
rect 10416 15136 10608 15153
rect 10480 15072 10544 15136
rect 10416 15055 10608 15072
rect 10480 14991 10544 15055
rect 10416 14974 10608 14991
rect 10480 14910 10544 14974
rect 10416 14893 10608 14910
rect 10480 14829 10544 14893
rect 10416 14812 10608 14829
rect 10480 14748 10544 14812
rect 10416 14731 10608 14748
rect 10480 14667 10544 14731
rect 10416 14650 10608 14667
rect 10480 14586 10544 14650
rect 10416 14569 10608 14586
rect 10480 14505 10544 14569
rect 10416 14488 10608 14505
rect 10480 14424 10544 14488
rect 10416 14407 10608 14424
rect 10480 14343 10544 14407
rect 10416 14326 10608 14343
rect 10480 14262 10544 14326
rect 10416 14245 10608 14262
rect 10480 14181 10544 14245
rect 10416 14164 10608 14181
rect 10480 14100 10544 14164
rect 10416 14083 10608 14100
rect 10480 14019 10544 14083
rect 10416 14002 10608 14019
rect 10480 13938 10544 14002
rect 10416 13921 10608 13938
rect 10480 13857 10544 13921
rect 10416 13840 10608 13857
rect 10480 13776 10544 13840
rect 10416 13759 10608 13776
rect 10480 13695 10544 13759
rect 10416 13678 10608 13695
rect 10480 13614 10544 13678
rect 10416 13607 10608 13614
rect 11408 18592 11600 21136
rect 11908 23686 12092 26632
tri 12892 26624 12900 26632 ne
rect 11908 23630 11913 23686
rect 11969 23630 12031 23686
rect 12087 23630 12092 23686
rect 11908 23606 12092 23630
rect 11908 23550 11913 23606
rect 11969 23550 12031 23606
rect 12087 23550 12092 23606
rect 11908 23526 12092 23550
rect 11908 23470 11913 23526
rect 11969 23470 12031 23526
rect 12087 23470 12092 23526
rect 11908 23446 12092 23470
rect 11908 23390 11913 23446
rect 11969 23390 12031 23446
rect 12087 23390 12092 23446
rect 11908 23366 12092 23390
rect 11908 23310 11913 23366
rect 11969 23310 12031 23366
rect 12087 23310 12092 23366
rect 11908 23286 12092 23310
rect 11908 23230 11913 23286
rect 11969 23230 12031 23286
rect 12087 23230 12092 23286
rect 11908 23206 12092 23230
rect 11908 23150 11913 23206
rect 11969 23150 12031 23206
rect 12087 23150 12092 23206
rect 11908 23126 12092 23150
rect 11908 23070 11913 23126
rect 11969 23070 12031 23126
rect 12087 23070 12092 23126
rect 11908 23046 12092 23070
rect 11908 22990 11913 23046
rect 11969 22990 12031 23046
rect 12087 22990 12092 23046
rect 11908 22966 12092 22990
rect 11908 22910 11913 22966
rect 11969 22910 12031 22966
rect 12087 22910 12092 22966
rect 11908 22886 12092 22910
rect 11908 22830 11913 22886
rect 11969 22830 12031 22886
rect 12087 22830 12092 22886
rect 11908 22806 12092 22830
rect 11908 22750 11913 22806
rect 11969 22750 12031 22806
rect 12087 22750 12092 22806
rect 11908 22726 12092 22750
rect 11908 22670 11913 22726
rect 11969 22670 12031 22726
rect 12087 22670 12092 22726
rect 11908 22646 12092 22670
rect 11908 22590 11913 22646
rect 11969 22590 12031 22646
rect 12087 22590 12092 22646
rect 11908 22566 12092 22590
rect 11908 22510 11913 22566
rect 11969 22510 12031 22566
rect 12087 22510 12092 22566
rect 11908 22486 12092 22510
rect 11908 22430 11913 22486
rect 11969 22430 12031 22486
rect 12087 22430 12092 22486
rect 11908 22406 12092 22430
rect 11908 22350 11913 22406
rect 11969 22350 12031 22406
rect 12087 22350 12092 22406
rect 11908 22326 12092 22350
rect 11908 22270 11913 22326
rect 11969 22270 12031 22326
rect 12087 22270 12092 22326
rect 11908 22245 12092 22270
rect 11908 22189 11913 22245
rect 11969 22189 12031 22245
rect 12087 22189 12092 22245
rect 11908 22164 12092 22189
rect 11908 22108 11913 22164
rect 11969 22108 12031 22164
rect 12087 22108 12092 22164
rect 11908 22083 12092 22108
rect 11908 22027 11913 22083
rect 11969 22027 12031 22083
rect 12087 22027 12092 22083
rect 11908 22002 12092 22027
rect 11908 21946 11913 22002
rect 11969 21946 12031 22002
rect 12087 21946 12092 22002
rect 11908 21921 12092 21946
rect 11908 21865 11913 21921
rect 11969 21865 12031 21921
rect 12087 21865 12092 21921
rect 11908 21840 12092 21865
rect 11908 21784 11913 21840
rect 11969 21784 12031 21840
rect 12087 21784 12092 21840
rect 11908 21759 12092 21784
rect 11908 21703 11913 21759
rect 11969 21703 12031 21759
rect 12087 21703 12092 21759
rect 11908 21678 12092 21703
rect 11908 21622 11913 21678
rect 11969 21622 12031 21678
rect 12087 21622 12092 21678
rect 11908 21597 12092 21622
rect 11908 21541 11913 21597
rect 11969 21541 12031 21597
rect 12087 21541 12092 21597
rect 11908 21516 12092 21541
rect 11908 21460 11913 21516
rect 11969 21460 12031 21516
rect 12087 21460 12092 21516
rect 11908 21435 12092 21460
rect 11908 21379 11913 21435
rect 11969 21379 12031 21435
rect 12087 21379 12092 21435
rect 11908 21354 12092 21379
rect 11908 21298 11913 21354
rect 11969 21298 12031 21354
rect 12087 21298 12092 21354
rect 11908 21273 12092 21298
rect 11908 21217 11913 21273
rect 11969 21217 12031 21273
rect 12087 21217 12092 21273
rect 11908 21192 12092 21217
rect 11908 21136 11913 21192
rect 11969 21136 12031 21192
rect 12087 21136 12092 21192
rect 11908 19673 12092 21136
rect 11972 19609 12028 19673
rect 11908 19581 12092 19609
rect 11972 19517 12028 19581
rect 11908 19489 12092 19517
rect 11972 19425 12028 19489
rect 11908 19397 12092 19425
rect 11972 19333 12028 19397
rect 11908 19305 12092 19333
rect 11972 19241 12028 19305
rect 11908 19212 12092 19241
rect 11972 19148 12028 19212
rect 11908 19139 12092 19148
rect 12400 23686 12592 23721
rect 12400 23630 12409 23686
rect 12465 23630 12527 23686
rect 12583 23630 12592 23686
rect 12400 23606 12592 23630
rect 12400 23550 12409 23606
rect 12465 23550 12527 23606
rect 12583 23550 12592 23606
rect 12400 23526 12592 23550
rect 12400 23470 12409 23526
rect 12465 23470 12527 23526
rect 12583 23470 12592 23526
rect 12400 23446 12592 23470
rect 12400 23390 12409 23446
rect 12465 23390 12527 23446
rect 12583 23390 12592 23446
rect 12400 23366 12592 23390
rect 12400 23310 12409 23366
rect 12465 23310 12527 23366
rect 12583 23310 12592 23366
rect 12400 23286 12592 23310
rect 12400 23230 12409 23286
rect 12465 23230 12527 23286
rect 12583 23230 12592 23286
rect 12400 23206 12592 23230
rect 12400 23150 12409 23206
rect 12465 23150 12527 23206
rect 12583 23150 12592 23206
rect 12400 23126 12592 23150
rect 12400 23070 12409 23126
rect 12465 23070 12527 23126
rect 12583 23070 12592 23126
rect 12400 23046 12592 23070
rect 12400 22990 12409 23046
rect 12465 22990 12527 23046
rect 12583 22990 12592 23046
rect 12400 22966 12592 22990
rect 12400 22910 12409 22966
rect 12465 22910 12527 22966
rect 12583 22910 12592 22966
rect 12400 22886 12592 22910
rect 12400 22830 12409 22886
rect 12465 22830 12527 22886
rect 12583 22830 12592 22886
rect 12400 22806 12592 22830
rect 12400 22750 12409 22806
rect 12465 22750 12527 22806
rect 12583 22750 12592 22806
rect 12400 22726 12592 22750
rect 12400 22670 12409 22726
rect 12465 22670 12527 22726
rect 12583 22670 12592 22726
rect 12400 22646 12592 22670
rect 12400 22590 12409 22646
rect 12465 22590 12527 22646
rect 12583 22590 12592 22646
rect 12400 22566 12592 22590
rect 12400 22510 12409 22566
rect 12465 22510 12527 22566
rect 12583 22510 12592 22566
rect 12400 22486 12592 22510
rect 12400 22430 12409 22486
rect 12465 22430 12527 22486
rect 12583 22430 12592 22486
rect 12400 22406 12592 22430
rect 12400 22350 12409 22406
rect 12465 22350 12527 22406
rect 12583 22350 12592 22406
rect 12400 22326 12592 22350
rect 12400 22270 12409 22326
rect 12465 22270 12527 22326
rect 12583 22270 12592 22326
rect 12400 22245 12592 22270
rect 12400 22189 12409 22245
rect 12465 22189 12527 22245
rect 12583 22189 12592 22245
rect 12400 22164 12592 22189
rect 12400 22108 12409 22164
rect 12465 22108 12527 22164
rect 12583 22108 12592 22164
rect 12400 22083 12592 22108
rect 12400 22027 12409 22083
rect 12465 22027 12527 22083
rect 12583 22027 12592 22083
rect 12400 22002 12592 22027
rect 12400 21946 12409 22002
rect 12465 21946 12527 22002
rect 12583 21946 12592 22002
rect 12400 21921 12592 21946
rect 12400 21865 12409 21921
rect 12465 21865 12527 21921
rect 12583 21865 12592 21921
rect 12400 21840 12592 21865
rect 12400 21784 12409 21840
rect 12465 21784 12527 21840
rect 12583 21784 12592 21840
rect 12400 21759 12592 21784
rect 12400 21703 12409 21759
rect 12465 21703 12527 21759
rect 12583 21703 12592 21759
rect 12400 21678 12592 21703
rect 12400 21622 12409 21678
rect 12465 21622 12527 21678
rect 12583 21622 12592 21678
rect 12400 21597 12592 21622
rect 12400 21541 12409 21597
rect 12465 21541 12527 21597
rect 12583 21541 12592 21597
rect 12400 21516 12592 21541
rect 12400 21460 12409 21516
rect 12465 21460 12527 21516
rect 12583 21460 12592 21516
rect 12400 21435 12592 21460
rect 12400 21379 12409 21435
rect 12465 21379 12527 21435
rect 12583 21379 12592 21435
rect 12400 21354 12592 21379
rect 12400 21298 12409 21354
rect 12465 21298 12527 21354
rect 12583 21298 12592 21354
rect 12400 21273 12592 21298
rect 12400 21217 12409 21273
rect 12465 21217 12527 21273
rect 12583 21217 12592 21273
rect 12400 21192 12592 21217
rect 12400 21136 12409 21192
rect 12465 21136 12527 21192
rect 12583 21136 12592 21192
rect 11472 18528 11536 18592
rect 11408 18512 11600 18528
rect 11472 18448 11536 18512
rect 11408 18432 11600 18448
rect 11472 18368 11536 18432
rect 11408 18352 11600 18368
rect 11472 18288 11536 18352
rect 11408 18272 11600 18288
rect 11472 18208 11536 18272
rect 11408 18192 11600 18208
rect 11472 18128 11536 18192
rect 11408 18112 11600 18128
rect 11472 18048 11536 18112
rect 11408 18032 11600 18048
rect 11472 17968 11536 18032
rect 11408 17952 11600 17968
rect 11472 17888 11536 17952
rect 11408 17872 11600 17888
rect 11472 17808 11536 17872
rect 11408 17792 11600 17808
rect 11472 17728 11536 17792
rect 11408 17712 11600 17728
rect 11472 17648 11536 17712
rect 11408 17632 11600 17648
rect 11472 17568 11536 17632
rect 11408 17552 11600 17568
rect 11472 17488 11536 17552
rect 11408 17472 11600 17488
rect 11472 17408 11536 17472
rect 11408 17392 11600 17408
rect 11472 17328 11536 17392
rect 11408 17312 11600 17328
rect 11472 17248 11536 17312
rect 11408 17232 11600 17248
rect 11472 17168 11536 17232
rect 11408 17152 11600 17168
rect 11472 17088 11536 17152
rect 11408 17072 11600 17088
rect 11472 17008 11536 17072
rect 11408 16992 11600 17008
rect 11472 16928 11536 16992
rect 11408 16912 11600 16928
rect 11472 16848 11536 16912
rect 11408 16832 11600 16848
rect 11472 16768 11536 16832
rect 11408 16752 11600 16768
rect 11472 16688 11536 16752
rect 11408 16672 11600 16688
rect 11472 16608 11536 16672
rect 11408 16592 11600 16608
rect 11472 16528 11536 16592
rect 11408 16512 11600 16528
rect 11472 16448 11536 16512
rect 11408 16432 11600 16448
rect 11472 16368 11536 16432
rect 11408 16351 11600 16368
rect 11472 16287 11536 16351
rect 11408 16270 11600 16287
rect 11472 16206 11536 16270
rect 11408 16189 11600 16206
rect 11472 16125 11536 16189
rect 11408 16108 11600 16125
rect 11472 16044 11536 16108
rect 11408 16027 11600 16044
rect 11472 15963 11536 16027
rect 11408 15946 11600 15963
rect 11472 15882 11536 15946
rect 11408 15865 11600 15882
rect 11472 15801 11536 15865
rect 11408 15784 11600 15801
rect 11472 15720 11536 15784
rect 11408 15703 11600 15720
rect 11472 15639 11536 15703
rect 11408 15622 11600 15639
rect 11472 15558 11536 15622
rect 11408 15541 11600 15558
rect 11472 15477 11536 15541
rect 11408 15460 11600 15477
rect 11472 15396 11536 15460
rect 11408 15379 11600 15396
rect 11472 15315 11536 15379
rect 11408 15298 11600 15315
rect 11472 15234 11536 15298
rect 11408 15217 11600 15234
rect 11472 15153 11536 15217
rect 11408 15136 11600 15153
rect 11472 15072 11536 15136
rect 11408 15055 11600 15072
rect 11472 14991 11536 15055
rect 11408 14974 11600 14991
rect 11472 14910 11536 14974
rect 11408 14893 11600 14910
rect 11472 14829 11536 14893
rect 11408 14812 11600 14829
rect 11472 14748 11536 14812
rect 11408 14731 11600 14748
rect 11472 14667 11536 14731
rect 11408 14650 11600 14667
rect 11472 14586 11536 14650
rect 11408 14569 11600 14586
rect 11472 14505 11536 14569
rect 11408 14488 11600 14505
rect 11472 14424 11536 14488
rect 11408 14407 11600 14424
rect 11472 14343 11536 14407
rect 11408 14326 11600 14343
rect 11472 14262 11536 14326
rect 11408 14245 11600 14262
rect 11472 14181 11536 14245
rect 11408 14164 11600 14181
rect 11472 14100 11536 14164
rect 11408 14083 11600 14100
rect 11472 14019 11536 14083
rect 11408 14002 11600 14019
rect 11472 13938 11536 14002
rect 11408 13921 11600 13938
rect 11472 13857 11536 13921
rect 11408 13840 11600 13857
rect 11472 13776 11536 13840
rect 11408 13759 11600 13776
rect 11472 13695 11536 13759
rect 11408 13678 11600 13695
rect 11472 13614 11536 13678
rect 11408 13607 11600 13614
rect 12400 18592 12592 21136
rect 12900 23686 13084 26632
tri 13646 27099 13653 27106 se
rect 13653 27099 14043 27106
rect 13646 27074 14043 27099
rect 13646 27010 13649 27074
rect 13713 27010 13757 27074
rect 13821 27010 13865 27074
rect 13929 27010 13973 27074
rect 14037 27010 14043 27074
rect 13646 26964 14043 27010
rect 13646 26900 13649 26964
rect 13713 26900 13757 26964
rect 13821 26900 13865 26964
rect 13929 26900 13973 26964
rect 14037 26900 14043 26964
rect 13646 26884 14043 26900
rect 13646 26854 13651 26884
rect 13707 26854 13733 26884
rect 13789 26854 13815 26884
rect 13871 26854 13897 26884
rect 13953 26854 13979 26884
rect 14035 26854 14043 26884
rect 13646 26790 13649 26854
rect 13713 26828 13733 26854
rect 13953 26828 13973 26854
rect 13713 26800 13757 26828
rect 13821 26800 13865 26828
rect 13929 26800 13973 26828
rect 13713 26790 13733 26800
rect 13953 26790 13973 26800
rect 14037 26790 14043 26854
rect 13646 26744 13651 26790
rect 13707 26744 13733 26790
rect 13789 26744 13815 26790
rect 13871 26744 13897 26790
rect 13953 26744 13979 26790
rect 14035 26744 14043 26790
rect 13646 26680 13649 26744
rect 13713 26716 13757 26744
rect 13821 26716 13865 26744
rect 13929 26716 13973 26744
rect 13713 26680 13733 26716
rect 13953 26680 13973 26716
rect 14037 26680 14043 26744
rect 13646 26660 13651 26680
rect 13707 26660 13733 26680
rect 13789 26660 13815 26680
rect 13871 26660 13897 26680
rect 13953 26660 13979 26680
rect 14035 26660 14043 26680
rect 13646 26634 14043 26660
rect 13646 26570 13649 26634
rect 13713 26632 13757 26634
rect 13821 26632 13865 26634
rect 13929 26632 13973 26634
rect 13713 26576 13733 26632
rect 13953 26576 13973 26632
rect 13713 26570 13757 26576
rect 13821 26570 13865 26576
rect 13929 26570 13973 26576
rect 14037 26570 14043 26634
rect 13646 26548 14043 26570
rect 13646 26524 13651 26548
rect 13707 26524 13733 26548
rect 13789 26524 13815 26548
rect 13871 26524 13897 26548
rect 13953 26524 13979 26548
rect 14035 26524 14043 26548
rect 13646 26460 13649 26524
rect 13713 26492 13733 26524
rect 13953 26492 13973 26524
rect 13713 26460 13757 26492
rect 13821 26460 13865 26492
rect 13929 26460 13973 26492
rect 14037 26460 14043 26524
rect 13646 26413 14043 26460
rect 13646 26349 13649 26413
rect 13713 26349 13757 26413
rect 13821 26349 13865 26413
rect 13929 26349 13973 26413
rect 14037 26349 14043 26413
rect 13646 26341 14043 26349
tri 13646 26333 13654 26341 ne
rect 13654 26333 14043 26341
tri 13654 26320 13667 26333 ne
rect 13667 26320 14043 26333
tri 13667 26277 13710 26320 ne
rect 13710 26314 14043 26320
rect 13710 26277 13843 26314
tri 13710 26252 13735 26277 ne
rect 13735 26252 13843 26277
tri 13735 26196 13791 26252 ne
rect 13791 26250 13843 26252
rect 13907 26250 13951 26314
rect 14015 26250 14043 26314
rect 13791 26213 14043 26250
rect 13791 26196 13843 26213
tri 13791 26171 13816 26196 ne
rect 13816 26171 13843 26196
tri 13816 26154 13833 26171 ne
rect 13833 26149 13843 26171
rect 13907 26149 13951 26213
rect 14015 26149 14043 26213
rect 13833 26117 14043 26149
rect 13833 26115 14041 26117
tri 14041 26115 14043 26117 nw
rect 14167 27321 14283 27377
rect 14339 27321 14381 27377
rect 14437 27321 14479 27377
rect 14535 27321 14577 27377
rect 14633 27321 14784 27377
rect 14167 27297 14784 27321
rect 14167 27241 14283 27297
rect 14339 27241 14381 27297
rect 14437 27241 14479 27297
rect 14535 27241 14577 27297
rect 14633 27241 14784 27297
rect 14167 27217 14784 27241
rect 14167 27161 14283 27217
rect 14339 27161 14381 27217
rect 14437 27161 14479 27217
rect 14535 27161 14577 27217
rect 14633 27161 14784 27217
rect 14167 27137 14784 27161
rect 14167 27081 14283 27137
rect 14339 27081 14381 27137
rect 14437 27081 14479 27137
rect 14535 27081 14577 27137
rect 14633 27081 14784 27137
rect 14167 27057 14784 27081
rect 14167 27001 14283 27057
rect 14339 27001 14381 27057
rect 14437 27001 14479 27057
rect 14535 27001 14577 27057
rect 14633 27001 14784 27057
rect 14167 26977 14784 27001
rect 14167 26921 14283 26977
rect 14339 26921 14381 26977
rect 14437 26921 14479 26977
rect 14535 26921 14577 26977
rect 14633 26921 14784 26977
rect 14167 26897 14784 26921
rect 14167 26841 14283 26897
rect 14339 26841 14381 26897
rect 14437 26841 14479 26897
rect 14535 26841 14577 26897
rect 14633 26841 14784 26897
rect 14167 26817 14784 26841
rect 14167 26761 14283 26817
rect 14339 26761 14381 26817
rect 14437 26761 14479 26817
rect 14535 26761 14577 26817
rect 14633 26761 14784 26817
rect 14167 26737 14784 26761
rect 14167 26681 14283 26737
rect 14339 26681 14381 26737
rect 14437 26681 14479 26737
rect 14535 26681 14577 26737
rect 14633 26681 14784 26737
rect 14167 26657 14784 26681
rect 14167 26601 14283 26657
rect 14339 26601 14381 26657
rect 14437 26601 14479 26657
rect 14535 26601 14577 26657
rect 14633 26601 14784 26657
rect 14167 26576 14784 26601
rect 14167 26520 14283 26576
rect 14339 26520 14381 26576
rect 14437 26520 14479 26576
rect 14535 26520 14577 26576
rect 14633 26520 14784 26576
rect 14167 26495 14784 26520
rect 14167 26439 14283 26495
rect 14339 26439 14381 26495
rect 14437 26439 14479 26495
rect 14535 26439 14577 26495
rect 14633 26439 14784 26495
rect 14167 26414 14784 26439
rect 14167 26358 14283 26414
rect 14339 26358 14381 26414
rect 14437 26358 14479 26414
rect 14535 26358 14577 26414
rect 14633 26358 14784 26414
rect 14167 26333 14784 26358
rect 14167 26277 14283 26333
rect 14339 26277 14381 26333
rect 14437 26277 14479 26333
rect 14535 26277 14577 26333
rect 14633 26277 14784 26333
rect 14167 26252 14784 26277
rect 14167 26196 14283 26252
rect 14339 26196 14381 26252
rect 14437 26196 14479 26252
rect 14535 26196 14577 26252
rect 14633 26196 14784 26252
rect 14167 26171 14784 26196
rect 14167 26115 14283 26171
rect 14339 26115 14381 26171
rect 14437 26115 14479 26171
rect 14535 26115 14577 26171
rect 14633 26115 14784 26171
rect 13833 26112 14025 26115
rect 13833 26048 13843 26112
rect 13907 26048 13951 26112
rect 14015 26048 14025 26112
tri 14025 26099 14041 26115 nw
rect 13833 26010 14025 26048
rect 13833 25946 13843 26010
rect 13907 25946 13951 26010
rect 14015 25946 14025 26010
rect 13833 25908 14025 25946
rect 13833 25844 13843 25908
rect 13907 25844 13951 25908
rect 14015 25844 14025 25908
rect 13833 25806 14025 25844
rect 13833 25742 13843 25806
rect 13907 25742 13951 25806
rect 14015 25742 14025 25806
rect 13833 25704 14025 25742
rect 13833 25640 13843 25704
rect 13907 25640 13951 25704
rect 14015 25640 14025 25704
rect 13833 25602 14025 25640
rect 13833 25538 13843 25602
rect 13907 25538 13951 25602
rect 14015 25538 14025 25602
rect 13833 25500 14025 25538
rect 13833 25436 13843 25500
rect 13907 25436 13951 25500
rect 14015 25436 14025 25500
rect 13833 25398 14025 25436
rect 13833 25334 13843 25398
rect 13907 25334 13951 25398
rect 14015 25334 14025 25398
rect 13833 25296 14025 25334
rect 13833 25232 13843 25296
rect 13907 25232 13951 25296
rect 14015 25232 14025 25296
rect 13833 25194 14025 25232
rect 13833 25130 13843 25194
rect 13907 25130 13951 25194
rect 14015 25130 14025 25194
rect 13833 25092 14025 25130
rect 13833 25028 13843 25092
rect 13907 25028 13951 25092
rect 14015 25028 14025 25092
rect 13833 24990 14025 25028
rect 13833 24926 13843 24990
rect 13907 24926 13951 24990
rect 14015 24926 14025 24990
rect 13833 24888 14025 24926
rect 13833 24824 13843 24888
rect 13907 24824 13951 24888
rect 14015 24824 14025 24888
rect 13833 24786 14025 24824
rect 13833 24722 13843 24786
rect 13907 24722 13951 24786
rect 14015 24722 14025 24786
rect 13833 24684 14025 24722
rect 13833 24620 13843 24684
rect 13907 24620 13951 24684
rect 14015 24620 14025 24684
rect 13833 24582 14025 24620
rect 13833 24518 13843 24582
rect 13907 24518 13951 24582
rect 14015 24518 14025 24582
rect 13833 24480 14025 24518
rect 13833 24416 13843 24480
rect 13907 24416 13951 24480
rect 14015 24416 14025 24480
rect 13833 24378 14025 24416
rect 13833 24314 13843 24378
rect 13907 24314 13951 24378
rect 14015 24314 14025 24378
rect 13833 24276 14025 24314
rect 13833 24212 13843 24276
rect 13907 24212 13951 24276
rect 14015 24212 14025 24276
rect 13833 24174 14025 24212
rect 13833 24110 13843 24174
rect 13907 24110 13951 24174
rect 14015 24110 14025 24174
rect 13833 24072 14025 24110
rect 13833 24008 13843 24072
rect 13907 24008 13951 24072
rect 14015 24008 14025 24072
rect 13833 23970 14025 24008
rect 13833 23906 13843 23970
rect 13907 23906 13951 23970
rect 14015 23906 14025 23970
rect 13833 23868 14025 23906
rect 13833 23804 13843 23868
rect 13907 23804 13951 23868
rect 14015 23804 14025 23868
rect 13833 23766 14025 23804
rect 12900 23630 12905 23686
rect 12961 23630 13023 23686
rect 13079 23630 13084 23686
rect 12900 23606 13084 23630
rect 12900 23550 12905 23606
rect 12961 23550 13023 23606
rect 13079 23550 13084 23606
rect 12900 23526 13084 23550
rect 12900 23470 12905 23526
rect 12961 23470 13023 23526
rect 13079 23470 13084 23526
rect 12900 23446 13084 23470
rect 12900 23390 12905 23446
rect 12961 23390 13023 23446
rect 13079 23390 13084 23446
rect 12900 23366 13084 23390
rect 12900 23310 12905 23366
rect 12961 23310 13023 23366
rect 13079 23310 13084 23366
rect 12900 23286 13084 23310
rect 12900 23230 12905 23286
rect 12961 23230 13023 23286
rect 13079 23230 13084 23286
rect 12900 23206 13084 23230
rect 12900 23150 12905 23206
rect 12961 23150 13023 23206
rect 13079 23150 13084 23206
rect 12900 23126 13084 23150
rect 12900 23070 12905 23126
rect 12961 23070 13023 23126
rect 13079 23070 13084 23126
rect 12900 23046 13084 23070
rect 12900 22990 12905 23046
rect 12961 22990 13023 23046
rect 13079 22990 13084 23046
rect 12900 22966 13084 22990
rect 12900 22910 12905 22966
rect 12961 22910 13023 22966
rect 13079 22910 13084 22966
rect 12900 22886 13084 22910
rect 12900 22830 12905 22886
rect 12961 22830 13023 22886
rect 13079 22830 13084 22886
rect 12900 22806 13084 22830
rect 12900 22750 12905 22806
rect 12961 22750 13023 22806
rect 13079 22750 13084 22806
rect 12900 22726 13084 22750
rect 12900 22670 12905 22726
rect 12961 22670 13023 22726
rect 13079 22670 13084 22726
rect 12900 22646 13084 22670
rect 12900 22590 12905 22646
rect 12961 22590 13023 22646
rect 13079 22590 13084 22646
rect 12900 22566 13084 22590
rect 12900 22510 12905 22566
rect 12961 22510 13023 22566
rect 13079 22510 13084 22566
rect 12900 22486 13084 22510
rect 12900 22430 12905 22486
rect 12961 22430 13023 22486
rect 13079 22430 13084 22486
rect 12900 22406 13084 22430
rect 12900 22350 12905 22406
rect 12961 22350 13023 22406
rect 13079 22350 13084 22406
rect 12900 22326 13084 22350
rect 12900 22270 12905 22326
rect 12961 22270 13023 22326
rect 13079 22270 13084 22326
rect 12900 22245 13084 22270
rect 12900 22189 12905 22245
rect 12961 22189 13023 22245
rect 13079 22189 13084 22245
rect 12900 22164 13084 22189
rect 12900 22108 12905 22164
rect 12961 22108 13023 22164
rect 13079 22108 13084 22164
rect 12900 22083 13084 22108
rect 12900 22027 12905 22083
rect 12961 22027 13023 22083
rect 13079 22027 13084 22083
rect 12900 22002 13084 22027
rect 12900 21946 12905 22002
rect 12961 21946 13023 22002
rect 13079 21946 13084 22002
rect 12900 21921 13084 21946
rect 12900 21865 12905 21921
rect 12961 21865 13023 21921
rect 13079 21865 13084 21921
rect 12900 21840 13084 21865
rect 12900 21784 12905 21840
rect 12961 21784 13023 21840
rect 13079 21784 13084 21840
rect 12900 21759 13084 21784
rect 12900 21703 12905 21759
rect 12961 21703 13023 21759
rect 13079 21703 13084 21759
rect 12900 21678 13084 21703
rect 12900 21622 12905 21678
rect 12961 21622 13023 21678
rect 13079 21622 13084 21678
rect 12900 21597 13084 21622
rect 12900 21541 12905 21597
rect 12961 21541 13023 21597
rect 13079 21541 13084 21597
rect 12900 21516 13084 21541
rect 12900 21460 12905 21516
rect 12961 21460 13023 21516
rect 13079 21460 13084 21516
rect 12900 21435 13084 21460
rect 12900 21379 12905 21435
rect 12961 21379 13023 21435
rect 13079 21379 13084 21435
rect 12900 21354 13084 21379
rect 12900 21298 12905 21354
rect 12961 21298 13023 21354
rect 13079 21298 13084 21354
rect 12900 21273 13084 21298
rect 12900 21217 12905 21273
rect 12961 21217 13023 21273
rect 13079 21217 13084 21273
rect 12900 21192 13084 21217
rect 12900 21136 12905 21192
rect 12961 21136 13023 21192
rect 13079 21136 13084 21192
rect 12900 20054 13084 21136
rect 12964 19990 13020 20054
rect 12900 19962 13084 19990
rect 12964 19898 13020 19962
rect 12900 19870 13084 19898
rect 12964 19806 13020 19870
rect 12900 19778 13084 19806
rect 12964 19714 13020 19778
rect 12900 19686 13084 19714
rect 12964 19622 13020 19686
rect 12900 19593 13084 19622
rect 12964 19529 13020 19593
rect 12900 19139 13084 19529
rect 13392 23686 13584 23721
rect 13392 23630 13401 23686
rect 13457 23630 13519 23686
rect 13575 23630 13584 23686
rect 13392 23606 13584 23630
rect 13392 23550 13401 23606
rect 13457 23550 13519 23606
rect 13575 23550 13584 23606
rect 13392 23526 13584 23550
rect 13392 23470 13401 23526
rect 13457 23470 13519 23526
rect 13575 23470 13584 23526
rect 13392 23446 13584 23470
rect 13392 23390 13401 23446
rect 13457 23390 13519 23446
rect 13575 23390 13584 23446
rect 13392 23366 13584 23390
rect 13392 23310 13401 23366
rect 13457 23310 13519 23366
rect 13575 23310 13584 23366
rect 13392 23286 13584 23310
rect 13392 23230 13401 23286
rect 13457 23230 13519 23286
rect 13575 23230 13584 23286
rect 13392 23206 13584 23230
rect 13392 23150 13401 23206
rect 13457 23150 13519 23206
rect 13575 23150 13584 23206
rect 13392 23126 13584 23150
rect 13392 23070 13401 23126
rect 13457 23070 13519 23126
rect 13575 23070 13584 23126
rect 13392 23046 13584 23070
rect 13392 22990 13401 23046
rect 13457 22990 13519 23046
rect 13575 22990 13584 23046
rect 13392 22966 13584 22990
rect 13392 22910 13401 22966
rect 13457 22910 13519 22966
rect 13575 22910 13584 22966
rect 13392 22886 13584 22910
rect 13392 22830 13401 22886
rect 13457 22830 13519 22886
rect 13575 22830 13584 22886
rect 13392 22806 13584 22830
rect 13392 22750 13401 22806
rect 13457 22750 13519 22806
rect 13575 22750 13584 22806
rect 13392 22726 13584 22750
rect 13392 22670 13401 22726
rect 13457 22670 13519 22726
rect 13575 22670 13584 22726
rect 13392 22646 13584 22670
rect 13392 22590 13401 22646
rect 13457 22590 13519 22646
rect 13575 22590 13584 22646
rect 13392 22566 13584 22590
rect 13392 22510 13401 22566
rect 13457 22510 13519 22566
rect 13575 22510 13584 22566
rect 13392 22486 13584 22510
rect 13392 22430 13401 22486
rect 13457 22430 13519 22486
rect 13575 22430 13584 22486
rect 13392 22406 13584 22430
rect 13392 22350 13401 22406
rect 13457 22350 13519 22406
rect 13575 22350 13584 22406
rect 13392 22326 13584 22350
rect 13392 22270 13401 22326
rect 13457 22270 13519 22326
rect 13575 22270 13584 22326
rect 13392 22245 13584 22270
rect 13392 22189 13401 22245
rect 13457 22189 13519 22245
rect 13575 22189 13584 22245
rect 13392 22164 13584 22189
rect 13392 22108 13401 22164
rect 13457 22108 13519 22164
rect 13575 22108 13584 22164
rect 13392 22083 13584 22108
rect 13392 22027 13401 22083
rect 13457 22027 13519 22083
rect 13575 22027 13584 22083
rect 13392 22002 13584 22027
rect 13392 21946 13401 22002
rect 13457 21946 13519 22002
rect 13575 21946 13584 22002
rect 13392 21921 13584 21946
rect 13392 21865 13401 21921
rect 13457 21865 13519 21921
rect 13575 21865 13584 21921
rect 13392 21840 13584 21865
rect 13392 21784 13401 21840
rect 13457 21784 13519 21840
rect 13575 21784 13584 21840
rect 13392 21759 13584 21784
rect 13392 21703 13401 21759
rect 13457 21703 13519 21759
rect 13575 21703 13584 21759
rect 13392 21678 13584 21703
rect 13392 21622 13401 21678
rect 13457 21622 13519 21678
rect 13575 21622 13584 21678
rect 13392 21597 13584 21622
rect 13392 21541 13401 21597
rect 13457 21541 13519 21597
rect 13575 21541 13584 21597
rect 13392 21516 13584 21541
rect 13392 21460 13401 21516
rect 13457 21460 13519 21516
rect 13575 21460 13584 21516
rect 13392 21435 13584 21460
rect 13392 21379 13401 21435
rect 13457 21379 13519 21435
rect 13575 21379 13584 21435
rect 13392 21354 13584 21379
rect 13392 21298 13401 21354
rect 13457 21298 13519 21354
rect 13575 21298 13584 21354
rect 13392 21273 13584 21298
rect 13392 21217 13401 21273
rect 13457 21217 13519 21273
rect 13575 21217 13584 21273
rect 13392 21192 13584 21217
rect 13392 21136 13401 21192
rect 13457 21136 13519 21192
rect 13575 21136 13584 21192
rect 12464 18528 12528 18592
rect 12400 18512 12592 18528
rect 12464 18448 12528 18512
rect 12400 18432 12592 18448
rect 12464 18368 12528 18432
rect 12400 18352 12592 18368
rect 12464 18288 12528 18352
rect 12400 18272 12592 18288
rect 12464 18208 12528 18272
rect 12400 18192 12592 18208
rect 12464 18128 12528 18192
rect 12400 18112 12592 18128
rect 12464 18048 12528 18112
rect 12400 18032 12592 18048
rect 12464 17968 12528 18032
rect 12400 17952 12592 17968
rect 12464 17888 12528 17952
rect 12400 17872 12592 17888
rect 12464 17808 12528 17872
rect 12400 17792 12592 17808
rect 12464 17728 12528 17792
rect 12400 17712 12592 17728
rect 12464 17648 12528 17712
rect 12400 17632 12592 17648
rect 12464 17568 12528 17632
rect 12400 17552 12592 17568
rect 12464 17488 12528 17552
rect 12400 17472 12592 17488
rect 12464 17408 12528 17472
rect 12400 17392 12592 17408
rect 12464 17328 12528 17392
rect 12400 17312 12592 17328
rect 12464 17248 12528 17312
rect 12400 17232 12592 17248
rect 12464 17168 12528 17232
rect 12400 17152 12592 17168
rect 12464 17088 12528 17152
rect 12400 17072 12592 17088
rect 12464 17008 12528 17072
rect 12400 16992 12592 17008
rect 12464 16928 12528 16992
rect 12400 16912 12592 16928
rect 12464 16848 12528 16912
rect 12400 16832 12592 16848
rect 12464 16768 12528 16832
rect 12400 16752 12592 16768
rect 12464 16688 12528 16752
rect 12400 16672 12592 16688
rect 12464 16608 12528 16672
rect 12400 16592 12592 16608
rect 12464 16528 12528 16592
rect 12400 16512 12592 16528
rect 12464 16448 12528 16512
rect 12400 16432 12592 16448
rect 12464 16368 12528 16432
rect 12400 16351 12592 16368
rect 12464 16287 12528 16351
rect 12400 16270 12592 16287
rect 12464 16206 12528 16270
rect 12400 16189 12592 16206
rect 12464 16125 12528 16189
rect 12400 16108 12592 16125
rect 12464 16044 12528 16108
rect 12400 16027 12592 16044
rect 12464 15963 12528 16027
rect 12400 15946 12592 15963
rect 12464 15882 12528 15946
rect 12400 15865 12592 15882
rect 12464 15801 12528 15865
rect 12400 15784 12592 15801
rect 12464 15720 12528 15784
rect 12400 15703 12592 15720
rect 12464 15639 12528 15703
rect 12400 15622 12592 15639
rect 12464 15558 12528 15622
rect 12400 15541 12592 15558
rect 12464 15477 12528 15541
rect 12400 15460 12592 15477
rect 12464 15396 12528 15460
rect 12400 15379 12592 15396
rect 12464 15315 12528 15379
rect 12400 15298 12592 15315
rect 12464 15234 12528 15298
rect 12400 15217 12592 15234
rect 12464 15153 12528 15217
rect 12400 15136 12592 15153
rect 12464 15072 12528 15136
rect 12400 15055 12592 15072
rect 12464 14991 12528 15055
rect 12400 14974 12592 14991
rect 12464 14910 12528 14974
rect 12400 14893 12592 14910
rect 12464 14829 12528 14893
rect 12400 14812 12592 14829
rect 12464 14748 12528 14812
rect 12400 14731 12592 14748
rect 12464 14667 12528 14731
rect 12400 14650 12592 14667
rect 12464 14586 12528 14650
rect 12400 14569 12592 14586
rect 12464 14505 12528 14569
rect 12400 14488 12592 14505
rect 12464 14424 12528 14488
rect 12400 14407 12592 14424
rect 12464 14343 12528 14407
rect 12400 14326 12592 14343
rect 12464 14262 12528 14326
rect 12400 14245 12592 14262
rect 12464 14181 12528 14245
rect 12400 14164 12592 14181
rect 12464 14100 12528 14164
rect 12400 14083 12592 14100
rect 12464 14019 12528 14083
rect 12400 14002 12592 14019
rect 12464 13938 12528 14002
rect 12400 13921 12592 13938
rect 12464 13857 12528 13921
rect 12400 13840 12592 13857
rect 12464 13776 12528 13840
rect 12400 13759 12592 13776
rect 12464 13695 12528 13759
rect 12400 13678 12592 13695
rect 12464 13614 12528 13678
rect 12400 13607 12592 13614
rect 13392 18592 13584 21136
rect 13833 23702 13843 23766
rect 13907 23702 13951 23766
rect 14015 23702 14025 23766
rect 13833 23686 14025 23702
rect 13833 23630 13838 23686
rect 13894 23664 13956 23686
rect 14012 23664 14025 23686
rect 13833 23606 13843 23630
rect 13833 23550 13838 23606
rect 13907 23600 13951 23664
rect 14015 23600 14025 23664
rect 13894 23562 13956 23600
rect 14012 23562 14025 23600
rect 13833 23526 13843 23550
rect 13833 23470 13838 23526
rect 13907 23498 13951 23562
rect 14015 23498 14025 23562
rect 13894 23470 13956 23498
rect 14012 23470 14025 23498
rect 13833 23460 14025 23470
rect 13833 23446 13843 23460
rect 13833 23390 13838 23446
rect 13907 23396 13951 23460
rect 14015 23396 14025 23460
rect 13894 23390 13956 23396
rect 14012 23390 14025 23396
rect 13833 23366 14025 23390
rect 13833 23310 13838 23366
rect 13894 23358 13956 23366
rect 14012 23358 14025 23366
rect 13833 23294 13843 23310
rect 13907 23294 13951 23358
rect 14015 23294 14025 23358
rect 13833 23286 14025 23294
rect 13833 23230 13838 23286
rect 13894 23256 13956 23286
rect 14012 23256 14025 23286
rect 13833 23206 13843 23230
rect 13833 23150 13838 23206
rect 13907 23192 13951 23256
rect 14015 23192 14025 23256
rect 13894 23154 13956 23192
rect 14012 23154 14025 23192
rect 13833 23126 13843 23150
rect 13833 23070 13838 23126
rect 13907 23090 13951 23154
rect 14015 23090 14025 23154
rect 13894 23070 13956 23090
rect 14012 23070 14025 23090
rect 13833 23052 14025 23070
rect 13833 23046 13843 23052
rect 13833 22990 13838 23046
rect 13833 22988 13843 22990
rect 13907 22988 13951 23052
rect 14015 22988 14025 23052
rect 13833 22966 14025 22988
rect 13833 22910 13838 22966
rect 13894 22950 13956 22966
rect 14012 22950 14025 22966
rect 13833 22886 13843 22910
rect 13907 22886 13951 22950
rect 14015 22886 14025 22950
rect 13833 22830 13838 22886
rect 13894 22848 13956 22886
rect 14012 22848 14025 22886
rect 13833 22806 13843 22830
rect 13833 22750 13838 22806
rect 13907 22784 13951 22848
rect 14015 22784 14025 22848
rect 13894 22750 13956 22784
rect 14012 22750 14025 22784
rect 13833 22746 14025 22750
rect 13833 22726 13843 22746
rect 13833 22670 13838 22726
rect 13907 22682 13951 22746
rect 14015 22682 14025 22746
rect 13894 22670 13956 22682
rect 14012 22670 14025 22682
rect 13833 22646 14025 22670
rect 13833 22590 13838 22646
rect 13894 22644 13956 22646
rect 14012 22644 14025 22646
rect 13833 22580 13843 22590
rect 13907 22580 13951 22644
rect 14015 22580 14025 22644
rect 13833 22566 14025 22580
rect 13833 22510 13838 22566
rect 13894 22542 13956 22566
rect 14012 22542 14025 22566
rect 13833 22486 13843 22510
rect 13833 22430 13838 22486
rect 13907 22478 13951 22542
rect 14015 22478 14025 22542
rect 13894 22440 13956 22478
rect 14012 22440 14025 22478
rect 13833 22406 13843 22430
rect 13833 22350 13838 22406
rect 13907 22376 13951 22440
rect 14015 22376 14025 22440
rect 13894 22350 13956 22376
rect 14012 22350 14025 22376
rect 13833 22338 14025 22350
rect 13833 22326 13843 22338
rect 13833 22270 13838 22326
rect 13907 22274 13951 22338
rect 14015 22274 14025 22338
rect 13894 22270 13956 22274
rect 14012 22270 14025 22274
rect 13833 22245 14025 22270
rect 13833 22189 13838 22245
rect 13894 22236 13956 22245
rect 14012 22236 14025 22245
rect 13833 22172 13843 22189
rect 13907 22172 13951 22236
rect 14015 22172 14025 22236
rect 13833 22164 14025 22172
rect 13833 22108 13838 22164
rect 13894 22134 13956 22164
rect 14012 22134 14025 22164
rect 13833 22083 13843 22108
rect 13833 22027 13838 22083
rect 13907 22070 13951 22134
rect 14015 22070 14025 22134
rect 13894 22032 13956 22070
rect 14012 22032 14025 22070
rect 13833 22002 13843 22027
rect 13833 21946 13838 22002
rect 13907 21968 13951 22032
rect 14015 21968 14025 22032
rect 13894 21946 13956 21968
rect 14012 21946 14025 21968
rect 13833 21930 14025 21946
rect 13833 21921 13843 21930
rect 13833 21865 13838 21921
rect 13907 21866 13951 21930
rect 14015 21866 14025 21930
rect 13894 21865 13956 21866
rect 14012 21865 14025 21866
rect 13833 21840 14025 21865
rect 13833 21784 13838 21840
rect 13894 21828 13956 21840
rect 14012 21828 14025 21840
rect 13833 21764 13843 21784
rect 13907 21764 13951 21828
rect 14015 21764 14025 21828
rect 13833 21759 14025 21764
rect 13833 21703 13838 21759
rect 13894 21726 13956 21759
rect 14012 21726 14025 21759
rect 13833 21678 13843 21703
rect 13833 21622 13838 21678
rect 13907 21662 13951 21726
rect 14015 21662 14025 21726
rect 13894 21624 13956 21662
rect 14012 21624 14025 21662
rect 13833 21597 13843 21622
rect 13833 21541 13838 21597
rect 13907 21560 13951 21624
rect 14015 21560 14025 21624
rect 13894 21541 13956 21560
rect 14012 21541 14025 21560
rect 13833 21516 14025 21541
rect 13833 21460 13838 21516
rect 13894 21460 13956 21516
rect 14012 21460 14025 21516
rect 13833 21435 14025 21460
rect 13833 21379 13838 21435
rect 13894 21379 13956 21435
rect 14012 21379 14025 21435
rect 13833 21354 14025 21379
rect 13833 21298 13838 21354
rect 13894 21298 13956 21354
rect 14012 21298 14025 21354
rect 13833 21273 14025 21298
rect 13833 21217 13838 21273
rect 13894 21217 13956 21273
rect 14012 21217 14025 21273
rect 13833 21192 14025 21217
rect 13833 21136 13838 21192
rect 13894 21136 13956 21192
rect 14012 21136 14025 21192
rect 13833 21131 14025 21136
rect 14167 26090 14784 26115
rect 14167 26034 14283 26090
rect 14339 26034 14381 26090
rect 14437 26034 14479 26090
rect 14535 26034 14577 26090
rect 14633 26034 14784 26090
rect 14167 26009 14784 26034
rect 14167 25953 14283 26009
rect 14339 25953 14381 26009
rect 14437 25953 14479 26009
rect 14535 25953 14577 26009
rect 14633 25953 14784 26009
rect 14167 25928 14784 25953
rect 14167 25872 14283 25928
rect 14339 25872 14381 25928
rect 14437 25872 14479 25928
rect 14535 25872 14577 25928
rect 14633 25872 14784 25928
rect 14167 25847 14784 25872
rect 14167 25791 14283 25847
rect 14339 25791 14381 25847
rect 14437 25791 14479 25847
rect 14535 25791 14577 25847
rect 14633 25791 14784 25847
rect 14167 25766 14784 25791
rect 14167 25710 14283 25766
rect 14339 25710 14381 25766
rect 14437 25710 14479 25766
rect 14535 25710 14577 25766
rect 14633 25710 14784 25766
rect 14167 25685 14784 25710
rect 14167 25629 14283 25685
rect 14339 25629 14381 25685
rect 14437 25629 14479 25685
rect 14535 25629 14577 25685
rect 14633 25629 14784 25685
rect 14167 25604 14784 25629
rect 14167 25548 14283 25604
rect 14339 25548 14381 25604
rect 14437 25548 14479 25604
rect 14535 25548 14577 25604
rect 14633 25548 14784 25604
rect 14167 25523 14784 25548
rect 14167 25467 14283 25523
rect 14339 25467 14381 25523
rect 14437 25467 14479 25523
rect 14535 25467 14577 25523
rect 14633 25467 14784 25523
rect 14167 25442 14784 25467
rect 14167 25386 14283 25442
rect 14339 25386 14381 25442
rect 14437 25386 14479 25442
rect 14535 25386 14577 25442
rect 14633 25386 14784 25442
rect 14167 25361 14784 25386
rect 14167 25305 14283 25361
rect 14339 25305 14381 25361
rect 14437 25305 14479 25361
rect 14535 25305 14577 25361
rect 14633 25305 14784 25361
rect 14167 25280 14784 25305
rect 14167 25224 14283 25280
rect 14339 25224 14381 25280
rect 14437 25224 14479 25280
rect 14535 25224 14577 25280
rect 14633 25224 14784 25280
rect 14167 25199 14784 25224
rect 14167 25143 14283 25199
rect 14339 25143 14381 25199
rect 14437 25143 14479 25199
rect 14535 25143 14577 25199
rect 14633 25143 14784 25199
rect 14167 25118 14784 25143
rect 14167 25062 14283 25118
rect 14339 25062 14381 25118
rect 14437 25062 14479 25118
rect 14535 25062 14577 25118
rect 14633 25062 14784 25118
rect 14167 25037 14784 25062
rect 14167 24981 14283 25037
rect 14339 24981 14381 25037
rect 14437 24981 14479 25037
rect 14535 24981 14577 25037
rect 14633 24981 14784 25037
rect 14167 24956 14784 24981
rect 14167 24900 14283 24956
rect 14339 24900 14381 24956
rect 14437 24900 14479 24956
rect 14535 24900 14577 24956
rect 14633 24900 14784 24956
rect 14167 24875 14784 24900
rect 14167 24819 14283 24875
rect 14339 24819 14381 24875
rect 14437 24819 14479 24875
rect 14535 24819 14577 24875
rect 14633 24819 14784 24875
rect 14167 24794 14784 24819
rect 14167 24738 14283 24794
rect 14339 24738 14381 24794
rect 14437 24738 14479 24794
rect 14535 24738 14577 24794
rect 14633 24738 14784 24794
rect 14167 24713 14784 24738
rect 14167 24657 14283 24713
rect 14339 24657 14381 24713
rect 14437 24657 14479 24713
rect 14535 24657 14577 24713
rect 14633 24657 14784 24713
rect 14167 24632 14784 24657
rect 14167 24576 14283 24632
rect 14339 24576 14381 24632
rect 14437 24576 14479 24632
rect 14535 24576 14577 24632
rect 14633 24576 14784 24632
rect 14167 24551 14784 24576
rect 14167 24495 14283 24551
rect 14339 24495 14381 24551
rect 14437 24495 14479 24551
rect 14535 24495 14577 24551
rect 14633 24495 14784 24551
rect 14167 24470 14784 24495
rect 14167 24414 14283 24470
rect 14339 24414 14381 24470
rect 14437 24414 14479 24470
rect 14535 24414 14577 24470
rect 14633 24414 14784 24470
rect 14167 24389 14784 24414
rect 14167 24333 14283 24389
rect 14339 24333 14381 24389
rect 14437 24333 14479 24389
rect 14535 24333 14577 24389
rect 14633 24333 14784 24389
rect 14167 24308 14784 24333
rect 14167 24252 14283 24308
rect 14339 24252 14381 24308
rect 14437 24252 14479 24308
rect 14535 24252 14577 24308
rect 14633 24252 14784 24308
rect 14167 24227 14784 24252
rect 14167 24171 14283 24227
rect 14339 24171 14381 24227
rect 14437 24171 14479 24227
rect 14535 24171 14577 24227
rect 14633 24171 14784 24227
rect 14167 24146 14784 24171
rect 14167 24090 14283 24146
rect 14339 24090 14381 24146
rect 14437 24090 14479 24146
rect 14535 24090 14577 24146
rect 14633 24090 14784 24146
rect 14167 24065 14784 24090
rect 14167 24009 14283 24065
rect 14339 24009 14381 24065
rect 14437 24009 14479 24065
rect 14535 24009 14577 24065
rect 14633 24009 14784 24065
rect 14167 23984 14784 24009
rect 14167 23928 14283 23984
rect 14339 23928 14381 23984
rect 14437 23928 14479 23984
rect 14535 23928 14577 23984
rect 14633 23928 14784 23984
rect 14167 23903 14784 23928
rect 14167 23847 14283 23903
rect 14339 23847 14381 23903
rect 14437 23847 14479 23903
rect 14535 23847 14577 23903
rect 14633 23847 14784 23903
rect 14167 23822 14784 23847
rect 14167 23766 14283 23822
rect 14339 23766 14381 23822
rect 14437 23766 14479 23822
rect 14535 23766 14577 23822
rect 14633 23766 14784 23822
rect 14167 23741 14784 23766
rect 14167 23685 14283 23741
rect 14339 23685 14381 23741
rect 14437 23685 14479 23741
rect 14535 23685 14577 23741
rect 14633 23685 14784 23741
rect 14167 23660 14784 23685
rect 14167 23604 14283 23660
rect 14339 23604 14381 23660
rect 14437 23604 14479 23660
rect 14535 23604 14577 23660
rect 14633 23604 14784 23660
rect 14167 23579 14784 23604
rect 14167 23523 14283 23579
rect 14339 23523 14381 23579
rect 14437 23523 14479 23579
rect 14535 23523 14577 23579
rect 14633 23523 14784 23579
rect 14167 23498 14784 23523
rect 14167 23442 14283 23498
rect 14339 23442 14381 23498
rect 14437 23442 14479 23498
rect 14535 23442 14577 23498
rect 14633 23442 14784 23498
rect 14167 23417 14784 23442
rect 14167 23361 14283 23417
rect 14339 23361 14381 23417
rect 14437 23361 14479 23417
rect 14535 23361 14577 23417
rect 14633 23361 14784 23417
rect 14167 23336 14784 23361
rect 14167 23280 14283 23336
rect 14339 23280 14381 23336
rect 14437 23280 14479 23336
rect 14535 23280 14577 23336
rect 14633 23280 14784 23336
rect 14167 23255 14784 23280
rect 14167 23199 14283 23255
rect 14339 23199 14381 23255
rect 14437 23199 14479 23255
rect 14535 23199 14577 23255
rect 14633 23199 14784 23255
rect 14167 23174 14784 23199
rect 14167 23118 14283 23174
rect 14339 23118 14381 23174
rect 14437 23118 14479 23174
rect 14535 23118 14577 23174
rect 14633 23118 14784 23174
rect 14167 23093 14784 23118
rect 14167 23037 14283 23093
rect 14339 23037 14381 23093
rect 14437 23037 14479 23093
rect 14535 23037 14577 23093
rect 14633 23037 14784 23093
rect 14167 23012 14784 23037
rect 14167 22956 14283 23012
rect 14339 22956 14381 23012
rect 14437 22956 14479 23012
rect 14535 22956 14577 23012
rect 14633 22956 14784 23012
rect 14167 22931 14784 22956
rect 14167 22875 14283 22931
rect 14339 22875 14381 22931
rect 14437 22875 14479 22931
rect 14535 22875 14577 22931
rect 14633 22875 14784 22931
rect 14167 22850 14784 22875
rect 14167 22794 14283 22850
rect 14339 22794 14381 22850
rect 14437 22794 14479 22850
rect 14535 22794 14577 22850
rect 14633 22794 14784 22850
rect 14167 22769 14784 22794
rect 14167 22713 14283 22769
rect 14339 22713 14381 22769
rect 14437 22713 14479 22769
rect 14535 22713 14577 22769
rect 14633 22713 14784 22769
rect 14167 22688 14784 22713
rect 14167 22632 14283 22688
rect 14339 22632 14381 22688
rect 14437 22632 14479 22688
rect 14535 22632 14577 22688
rect 14633 22632 14784 22688
rect 14167 22607 14784 22632
rect 14167 22551 14283 22607
rect 14339 22551 14381 22607
rect 14437 22551 14479 22607
rect 14535 22551 14577 22607
rect 14633 22551 14784 22607
rect 14167 22526 14784 22551
rect 14167 22470 14283 22526
rect 14339 22470 14381 22526
rect 14437 22470 14479 22526
rect 14535 22470 14577 22526
rect 14633 22470 14784 22526
rect 14167 22445 14784 22470
rect 14167 22389 14283 22445
rect 14339 22389 14381 22445
rect 14437 22389 14479 22445
rect 14535 22389 14577 22445
rect 14633 22389 14784 22445
rect 14167 22364 14784 22389
rect 14167 22308 14283 22364
rect 14339 22308 14381 22364
rect 14437 22308 14479 22364
rect 14535 22308 14577 22364
rect 14633 22308 14784 22364
rect 14167 22283 14784 22308
rect 14167 22227 14283 22283
rect 14339 22227 14381 22283
rect 14437 22227 14479 22283
rect 14535 22227 14577 22283
rect 14633 22227 14784 22283
rect 14167 22202 14784 22227
rect 14167 22146 14283 22202
rect 14339 22146 14381 22202
rect 14437 22146 14479 22202
rect 14535 22146 14577 22202
rect 14633 22146 14784 22202
rect 14167 22121 14784 22146
rect 14167 22065 14283 22121
rect 14339 22065 14381 22121
rect 14437 22065 14479 22121
rect 14535 22065 14577 22121
rect 14633 22065 14784 22121
rect 14167 22040 14784 22065
rect 14167 21984 14283 22040
rect 14339 21984 14381 22040
rect 14437 21984 14479 22040
rect 14535 21984 14577 22040
rect 14633 21984 14784 22040
rect 14167 21959 14784 21984
rect 14167 21903 14283 21959
rect 14339 21903 14381 21959
rect 14437 21903 14479 21959
rect 14535 21903 14577 21959
rect 14633 21903 14784 21959
rect 14167 21878 14784 21903
rect 14167 21822 14283 21878
rect 14339 21822 14381 21878
rect 14437 21822 14479 21878
rect 14535 21822 14577 21878
rect 14633 21822 14784 21878
rect 14167 21797 14784 21822
rect 14167 21741 14283 21797
rect 14339 21741 14381 21797
rect 14437 21741 14479 21797
rect 14535 21741 14577 21797
rect 14633 21741 14784 21797
rect 14167 21716 14784 21741
rect 14167 21660 14283 21716
rect 14339 21660 14381 21716
rect 14437 21660 14479 21716
rect 14535 21660 14577 21716
rect 14633 21660 14784 21716
rect 14167 21635 14784 21660
rect 14167 21579 14283 21635
rect 14339 21579 14381 21635
rect 14437 21579 14479 21635
rect 14535 21579 14577 21635
rect 14633 21579 14784 21635
rect 14167 21554 14784 21579
rect 14167 21498 14283 21554
rect 14339 21498 14381 21554
rect 14437 21498 14479 21554
rect 14535 21498 14577 21554
rect 14633 21498 14784 21554
rect 14167 21473 14784 21498
rect 14167 21417 14283 21473
rect 14339 21417 14381 21473
rect 14437 21417 14479 21473
rect 14535 21417 14577 21473
rect 14633 21417 14784 21473
rect 14167 21392 14784 21417
rect 14167 21336 14283 21392
rect 14339 21336 14381 21392
rect 14437 21336 14479 21392
rect 14535 21336 14577 21392
rect 14633 21336 14784 21392
rect 14167 21311 14784 21336
rect 14167 21255 14283 21311
rect 14339 21255 14381 21311
rect 14437 21255 14479 21311
rect 14535 21255 14577 21311
rect 14633 21255 14784 21311
rect 14167 21230 14784 21255
rect 14167 21174 14283 21230
rect 14339 21174 14381 21230
rect 14437 21174 14479 21230
rect 14535 21174 14577 21230
rect 14633 21174 14784 21230
rect 14167 21149 14784 21174
rect 14167 21093 14283 21149
rect 14339 21093 14381 21149
rect 14437 21093 14479 21149
rect 14535 21093 14577 21149
rect 14633 21093 14784 21149
rect 14167 21068 14784 21093
rect 14167 21012 14283 21068
rect 14339 21012 14381 21068
rect 14437 21012 14479 21068
rect 14535 21012 14577 21068
rect 14633 21012 14784 21068
rect 14167 20987 14784 21012
rect 14167 20931 14283 20987
rect 14339 20931 14381 20987
rect 14437 20931 14479 20987
rect 14535 20931 14577 20987
rect 14633 20931 14784 20987
rect 14167 20906 14784 20931
rect 14167 20850 14283 20906
rect 14339 20850 14381 20906
rect 14437 20850 14479 20906
rect 14535 20850 14577 20906
rect 14633 20850 14784 20906
rect 14167 20825 14784 20850
rect 14167 20769 14283 20825
rect 14339 20769 14381 20825
rect 14437 20769 14479 20825
rect 14535 20769 14577 20825
rect 14633 20769 14784 20825
rect 14167 20744 14784 20769
rect 14167 20688 14283 20744
rect 14339 20688 14381 20744
rect 14437 20688 14479 20744
rect 14535 20688 14577 20744
rect 14633 20688 14784 20744
rect 14167 20663 14784 20688
tri 14150 20607 14167 20624 se
rect 14167 20607 14283 20663
rect 14339 20607 14381 20663
rect 14437 20607 14479 20663
rect 14535 20607 14577 20663
rect 14633 20607 14784 20663
tri 14125 20582 14150 20607 se
rect 14150 20582 14784 20607
tri 14069 20526 14125 20582 se
rect 14125 20526 14283 20582
rect 14339 20526 14381 20582
rect 14437 20526 14479 20582
rect 14535 20526 14577 20582
rect 14633 20526 14784 20582
tri 14064 20521 14069 20526 se
rect 14069 20521 14784 20526
rect 13456 18528 13520 18592
rect 13392 18512 13584 18528
rect 13456 18448 13520 18512
rect 13392 18432 13584 18448
rect 13456 18368 13520 18432
rect 13392 18352 13584 18368
rect 13456 18288 13520 18352
rect 13392 18272 13584 18288
rect 13456 18208 13520 18272
rect 13392 18192 13584 18208
rect 13456 18128 13520 18192
rect 13392 18112 13584 18128
rect 13456 18048 13520 18112
rect 13392 18032 13584 18048
rect 13456 17968 13520 18032
rect 13392 17952 13584 17968
rect 13456 17888 13520 17952
rect 13392 17872 13584 17888
rect 13456 17808 13520 17872
rect 13392 17792 13584 17808
rect 13456 17728 13520 17792
rect 13392 17712 13584 17728
rect 13456 17648 13520 17712
rect 13392 17632 13584 17648
rect 13456 17568 13520 17632
rect 13392 17552 13584 17568
rect 13456 17488 13520 17552
rect 13392 17472 13584 17488
rect 13456 17408 13520 17472
rect 13392 17392 13584 17408
rect 13456 17328 13520 17392
rect 13392 17312 13584 17328
rect 13456 17248 13520 17312
rect 13392 17232 13584 17248
rect 13456 17168 13520 17232
rect 13392 17152 13584 17168
rect 13456 17088 13520 17152
rect 13392 17072 13584 17088
rect 13456 17008 13520 17072
rect 13392 16992 13584 17008
rect 13456 16928 13520 16992
rect 13392 16912 13584 16928
rect 13456 16848 13520 16912
rect 13392 16832 13584 16848
rect 13456 16768 13520 16832
rect 13392 16752 13584 16768
rect 13456 16688 13520 16752
rect 13392 16672 13584 16688
rect 13456 16608 13520 16672
rect 13392 16592 13584 16608
rect 13456 16528 13520 16592
rect 13392 16512 13584 16528
rect 13456 16448 13520 16512
rect 13392 16432 13584 16448
rect 13456 16368 13520 16432
rect 13392 16351 13584 16368
rect 13456 16287 13520 16351
rect 13392 16270 13584 16287
rect 13456 16206 13520 16270
rect 13392 16189 13584 16206
rect 13456 16125 13520 16189
rect 13392 16108 13584 16125
rect 13456 16044 13520 16108
rect 13392 16027 13584 16044
rect 13456 15963 13520 16027
rect 13392 15946 13584 15963
rect 13456 15882 13520 15946
rect 13392 15865 13584 15882
rect 13456 15801 13520 15865
rect 13392 15784 13584 15801
rect 13456 15720 13520 15784
rect 13392 15703 13584 15720
rect 13456 15639 13520 15703
rect 13392 15622 13584 15639
rect 13456 15558 13520 15622
rect 13392 15541 13584 15558
rect 13456 15477 13520 15541
rect 13392 15460 13584 15477
rect 13456 15396 13520 15460
rect 13392 15379 13584 15396
rect 13456 15315 13520 15379
rect 13392 15298 13584 15315
rect 13456 15234 13520 15298
rect 13392 15217 13584 15234
rect 13456 15153 13520 15217
rect 13392 15136 13584 15153
rect 13456 15072 13520 15136
rect 13392 15055 13584 15072
rect 13456 14991 13520 15055
rect 13392 14974 13584 14991
rect 13456 14910 13520 14974
rect 13392 14893 13584 14910
rect 13456 14829 13520 14893
rect 13392 14812 13584 14829
rect 13456 14748 13520 14812
rect 13392 14731 13584 14748
rect 13456 14667 13520 14731
rect 13392 14650 13584 14667
rect 13456 14586 13520 14650
rect 13392 14569 13584 14586
rect 13456 14505 13520 14569
rect 13392 14488 13584 14505
rect 13456 14424 13520 14488
rect 13392 14407 13584 14424
rect 13456 14343 13520 14407
rect 13392 14326 13584 14343
rect 13456 14262 13520 14326
rect 13392 14245 13584 14262
rect 13456 14181 13520 14245
rect 13392 14164 13584 14181
rect 13456 14100 13520 14164
rect 13392 14083 13584 14100
rect 13456 14019 13520 14083
rect 13392 14002 13584 14019
rect 13456 13938 13520 14002
rect 13392 13921 13584 13938
rect 13456 13857 13520 13921
rect 13392 13840 13584 13857
rect 13456 13776 13520 13840
rect 13392 13759 13584 13776
rect 13456 13695 13520 13759
rect 13392 13678 13584 13695
rect 13456 13614 13520 13678
rect 13392 13607 13584 13614
tri 13769 20226 14064 20521 se
rect 14064 20226 14784 20521
rect 13769 20131 14784 20226
rect 13769 18590 14555 20131
tri 14555 19902 14784 20131 nw
rect 13769 18526 13777 18590
rect 13841 18526 13863 18590
rect 13927 18526 13949 18590
rect 14013 18526 14035 18590
rect 14099 18526 14121 18590
rect 14185 18526 14207 18590
rect 14271 18526 14293 18590
rect 14357 18526 14379 18590
rect 14443 18526 14465 18590
rect 14529 18526 14555 18590
rect 13769 18510 14555 18526
rect 13769 18446 13777 18510
rect 13841 18446 13863 18510
rect 13927 18446 13949 18510
rect 14013 18446 14035 18510
rect 14099 18446 14121 18510
rect 14185 18446 14207 18510
rect 14271 18446 14293 18510
rect 14357 18446 14379 18510
rect 14443 18446 14465 18510
rect 14529 18446 14555 18510
rect 13769 18430 14555 18446
rect 13769 18366 13777 18430
rect 13841 18366 13863 18430
rect 13927 18366 13949 18430
rect 14013 18366 14035 18430
rect 14099 18366 14121 18430
rect 14185 18366 14207 18430
rect 14271 18366 14293 18430
rect 14357 18366 14379 18430
rect 14443 18366 14465 18430
rect 14529 18366 14555 18430
rect 13769 18350 14555 18366
rect 13769 18286 13777 18350
rect 13841 18286 13863 18350
rect 13927 18286 13949 18350
rect 14013 18286 14035 18350
rect 14099 18286 14121 18350
rect 14185 18286 14207 18350
rect 14271 18286 14293 18350
rect 14357 18286 14379 18350
rect 14443 18286 14465 18350
rect 14529 18286 14555 18350
rect 13769 18270 14555 18286
rect 13769 18206 13777 18270
rect 13841 18206 13863 18270
rect 13927 18206 13949 18270
rect 14013 18206 14035 18270
rect 14099 18206 14121 18270
rect 14185 18206 14207 18270
rect 14271 18206 14293 18270
rect 14357 18206 14379 18270
rect 14443 18206 14465 18270
rect 14529 18206 14555 18270
rect 13769 18190 14555 18206
rect 13769 18126 13777 18190
rect 13841 18126 13863 18190
rect 13927 18126 13949 18190
rect 14013 18126 14035 18190
rect 14099 18126 14121 18190
rect 14185 18126 14207 18190
rect 14271 18126 14293 18190
rect 14357 18126 14379 18190
rect 14443 18126 14465 18190
rect 14529 18126 14555 18190
rect 13769 18110 14555 18126
rect 13769 18046 13777 18110
rect 13841 18046 13863 18110
rect 13927 18046 13949 18110
rect 14013 18046 14035 18110
rect 14099 18046 14121 18110
rect 14185 18046 14207 18110
rect 14271 18046 14293 18110
rect 14357 18046 14379 18110
rect 14443 18046 14465 18110
rect 14529 18046 14555 18110
rect 13769 18030 14555 18046
rect 13769 17966 13777 18030
rect 13841 17966 13863 18030
rect 13927 17966 13949 18030
rect 14013 17966 14035 18030
rect 14099 17966 14121 18030
rect 14185 17966 14207 18030
rect 14271 17966 14293 18030
rect 14357 17966 14379 18030
rect 14443 17966 14465 18030
rect 14529 17966 14555 18030
rect 13769 17950 14555 17966
rect 13769 17886 13777 17950
rect 13841 17886 13863 17950
rect 13927 17886 13949 17950
rect 14013 17886 14035 17950
rect 14099 17886 14121 17950
rect 14185 17886 14207 17950
rect 14271 17886 14293 17950
rect 14357 17886 14379 17950
rect 14443 17886 14465 17950
rect 14529 17886 14555 17950
rect 13769 17870 14555 17886
rect 13769 17806 13777 17870
rect 13841 17806 13863 17870
rect 13927 17806 13949 17870
rect 14013 17806 14035 17870
rect 14099 17806 14121 17870
rect 14185 17806 14207 17870
rect 14271 17806 14293 17870
rect 14357 17806 14379 17870
rect 14443 17806 14465 17870
rect 14529 17806 14555 17870
rect 13769 17790 14555 17806
rect 13769 17726 13777 17790
rect 13841 17726 13863 17790
rect 13927 17726 13949 17790
rect 14013 17726 14035 17790
rect 14099 17726 14121 17790
rect 14185 17726 14207 17790
rect 14271 17726 14293 17790
rect 14357 17726 14379 17790
rect 14443 17726 14465 17790
rect 14529 17726 14555 17790
rect 13769 17710 14555 17726
rect 13769 17646 13777 17710
rect 13841 17646 13863 17710
rect 13927 17646 13949 17710
rect 14013 17646 14035 17710
rect 14099 17646 14121 17710
rect 14185 17646 14207 17710
rect 14271 17646 14293 17710
rect 14357 17646 14379 17710
rect 14443 17646 14465 17710
rect 14529 17646 14555 17710
rect 13769 17630 14555 17646
rect 13769 17566 13777 17630
rect 13841 17566 13863 17630
rect 13927 17566 13949 17630
rect 14013 17566 14035 17630
rect 14099 17566 14121 17630
rect 14185 17566 14207 17630
rect 14271 17566 14293 17630
rect 14357 17566 14379 17630
rect 14443 17566 14465 17630
rect 14529 17566 14555 17630
rect 13769 17550 14555 17566
rect 13769 17486 13777 17550
rect 13841 17486 13863 17550
rect 13927 17486 13949 17550
rect 14013 17486 14035 17550
rect 14099 17486 14121 17550
rect 14185 17486 14207 17550
rect 14271 17486 14293 17550
rect 14357 17486 14379 17550
rect 14443 17486 14465 17550
rect 14529 17486 14555 17550
rect 13769 17470 14555 17486
rect 13769 17406 13777 17470
rect 13841 17406 13863 17470
rect 13927 17406 13949 17470
rect 14013 17406 14035 17470
rect 14099 17406 14121 17470
rect 14185 17406 14207 17470
rect 14271 17406 14293 17470
rect 14357 17406 14379 17470
rect 14443 17406 14465 17470
rect 14529 17406 14555 17470
rect 13769 17390 14555 17406
rect 13769 17326 13777 17390
rect 13841 17326 13863 17390
rect 13927 17326 13949 17390
rect 14013 17326 14035 17390
rect 14099 17326 14121 17390
rect 14185 17326 14207 17390
rect 14271 17326 14293 17390
rect 14357 17326 14379 17390
rect 14443 17326 14465 17390
rect 14529 17326 14555 17390
rect 13769 17310 14555 17326
rect 13769 17246 13777 17310
rect 13841 17246 13863 17310
rect 13927 17246 13949 17310
rect 14013 17246 14035 17310
rect 14099 17246 14121 17310
rect 14185 17246 14207 17310
rect 14271 17246 14293 17310
rect 14357 17246 14379 17310
rect 14443 17246 14465 17310
rect 14529 17246 14555 17310
rect 13769 17230 14555 17246
rect 13769 17166 13777 17230
rect 13841 17166 13863 17230
rect 13927 17166 13949 17230
rect 14013 17166 14035 17230
rect 14099 17166 14121 17230
rect 14185 17166 14207 17230
rect 14271 17166 14293 17230
rect 14357 17166 14379 17230
rect 14443 17166 14465 17230
rect 14529 17166 14555 17230
rect 13769 17150 14555 17166
rect 13769 17086 13777 17150
rect 13841 17086 13863 17150
rect 13927 17086 13949 17150
rect 14013 17086 14035 17150
rect 14099 17086 14121 17150
rect 14185 17086 14207 17150
rect 14271 17086 14293 17150
rect 14357 17086 14379 17150
rect 14443 17086 14465 17150
rect 14529 17086 14555 17150
rect 13769 17070 14555 17086
rect 13769 17006 13777 17070
rect 13841 17006 13863 17070
rect 13927 17006 13949 17070
rect 14013 17006 14035 17070
rect 14099 17006 14121 17070
rect 14185 17006 14207 17070
rect 14271 17006 14293 17070
rect 14357 17006 14379 17070
rect 14443 17006 14465 17070
rect 14529 17006 14555 17070
rect 13769 16990 14555 17006
rect 13769 16926 13777 16990
rect 13841 16926 13863 16990
rect 13927 16926 13949 16990
rect 14013 16926 14035 16990
rect 14099 16926 14121 16990
rect 14185 16926 14207 16990
rect 14271 16926 14293 16990
rect 14357 16926 14379 16990
rect 14443 16926 14465 16990
rect 14529 16926 14555 16990
rect 13769 16910 14555 16926
rect 13769 16846 13777 16910
rect 13841 16846 13863 16910
rect 13927 16846 13949 16910
rect 14013 16846 14035 16910
rect 14099 16846 14121 16910
rect 14185 16846 14207 16910
rect 14271 16846 14293 16910
rect 14357 16846 14379 16910
rect 14443 16846 14465 16910
rect 14529 16846 14555 16910
rect 13769 16830 14555 16846
rect 13769 16766 13777 16830
rect 13841 16766 13863 16830
rect 13927 16766 13949 16830
rect 14013 16766 14035 16830
rect 14099 16766 14121 16830
rect 14185 16766 14207 16830
rect 14271 16766 14293 16830
rect 14357 16766 14379 16830
rect 14443 16766 14465 16830
rect 14529 16766 14555 16830
rect 13769 16750 14555 16766
rect 13769 16686 13777 16750
rect 13841 16686 13863 16750
rect 13927 16686 13949 16750
rect 14013 16686 14035 16750
rect 14099 16686 14121 16750
rect 14185 16686 14207 16750
rect 14271 16686 14293 16750
rect 14357 16686 14379 16750
rect 14443 16686 14465 16750
rect 14529 16686 14555 16750
rect 13769 16670 14555 16686
rect 13769 16606 13777 16670
rect 13841 16606 13863 16670
rect 13927 16606 13949 16670
rect 14013 16606 14035 16670
rect 14099 16606 14121 16670
rect 14185 16606 14207 16670
rect 14271 16606 14293 16670
rect 14357 16606 14379 16670
rect 14443 16606 14465 16670
rect 14529 16606 14555 16670
rect 13769 16590 14555 16606
rect 13769 16526 13777 16590
rect 13841 16526 13863 16590
rect 13927 16526 13949 16590
rect 14013 16526 14035 16590
rect 14099 16526 14121 16590
rect 14185 16526 14207 16590
rect 14271 16526 14293 16590
rect 14357 16526 14379 16590
rect 14443 16526 14465 16590
rect 14529 16526 14555 16590
rect 13769 16510 14555 16526
rect 13769 16446 13777 16510
rect 13841 16446 13863 16510
rect 13927 16446 13949 16510
rect 14013 16446 14035 16510
rect 14099 16446 14121 16510
rect 14185 16446 14207 16510
rect 14271 16446 14293 16510
rect 14357 16446 14379 16510
rect 14443 16446 14465 16510
rect 14529 16446 14555 16510
rect 13769 16430 14555 16446
rect 13769 16366 13777 16430
rect 13841 16366 13863 16430
rect 13927 16366 13949 16430
rect 14013 16366 14035 16430
rect 14099 16366 14121 16430
rect 14185 16366 14207 16430
rect 14271 16366 14293 16430
rect 14357 16366 14379 16430
rect 14443 16366 14465 16430
rect 14529 16366 14555 16430
rect 13769 16350 14555 16366
rect 13769 16286 13777 16350
rect 13841 16286 13863 16350
rect 13927 16286 13949 16350
rect 14013 16286 14035 16350
rect 14099 16286 14121 16350
rect 14185 16286 14207 16350
rect 14271 16286 14293 16350
rect 14357 16286 14379 16350
rect 14443 16286 14465 16350
rect 14529 16286 14555 16350
rect 13769 16270 14555 16286
rect 13769 16206 13777 16270
rect 13841 16206 13863 16270
rect 13927 16206 13949 16270
rect 14013 16206 14035 16270
rect 14099 16206 14121 16270
rect 14185 16206 14207 16270
rect 14271 16206 14293 16270
rect 14357 16206 14379 16270
rect 14443 16206 14465 16270
rect 14529 16206 14555 16270
rect 13769 16190 14555 16206
rect 13769 16126 13777 16190
rect 13841 16126 13863 16190
rect 13927 16126 13949 16190
rect 14013 16126 14035 16190
rect 14099 16126 14121 16190
rect 14185 16126 14207 16190
rect 14271 16126 14293 16190
rect 14357 16126 14379 16190
rect 14443 16126 14465 16190
rect 14529 16126 14555 16190
rect 13769 16110 14555 16126
rect 13769 16046 13777 16110
rect 13841 16046 13863 16110
rect 13927 16046 13949 16110
rect 14013 16046 14035 16110
rect 14099 16046 14121 16110
rect 14185 16046 14207 16110
rect 14271 16046 14293 16110
rect 14357 16046 14379 16110
rect 14443 16046 14465 16110
rect 14529 16046 14555 16110
rect 13769 16030 14555 16046
rect 13769 15966 13777 16030
rect 13841 15966 13863 16030
rect 13927 15966 13949 16030
rect 14013 15966 14035 16030
rect 14099 15966 14121 16030
rect 14185 15966 14207 16030
rect 14271 15966 14293 16030
rect 14357 15966 14379 16030
rect 14443 15966 14465 16030
rect 14529 15966 14555 16030
rect 13769 15950 14555 15966
rect 13769 15886 13777 15950
rect 13841 15886 13863 15950
rect 13927 15886 13949 15950
rect 14013 15886 14035 15950
rect 14099 15886 14121 15950
rect 14185 15886 14207 15950
rect 14271 15886 14293 15950
rect 14357 15886 14379 15950
rect 14443 15886 14465 15950
rect 14529 15886 14555 15950
rect 13769 15870 14555 15886
rect 13769 15806 13777 15870
rect 13841 15806 13863 15870
rect 13927 15806 13949 15870
rect 14013 15806 14035 15870
rect 14099 15806 14121 15870
rect 14185 15806 14207 15870
rect 14271 15806 14293 15870
rect 14357 15806 14379 15870
rect 14443 15806 14465 15870
rect 14529 15806 14555 15870
rect 13769 15790 14555 15806
rect 13769 15726 13777 15790
rect 13841 15726 13863 15790
rect 13927 15726 13949 15790
rect 14013 15726 14035 15790
rect 14099 15726 14121 15790
rect 14185 15726 14207 15790
rect 14271 15726 14293 15790
rect 14357 15726 14379 15790
rect 14443 15726 14465 15790
rect 14529 15726 14555 15790
rect 13769 15710 14555 15726
rect 13769 15646 13777 15710
rect 13841 15646 13863 15710
rect 13927 15646 13949 15710
rect 14013 15646 14035 15710
rect 14099 15646 14121 15710
rect 14185 15646 14207 15710
rect 14271 15646 14293 15710
rect 14357 15646 14379 15710
rect 14443 15646 14465 15710
rect 14529 15646 14555 15710
rect 13769 15630 14555 15646
rect 13769 15566 13777 15630
rect 13841 15566 13863 15630
rect 13927 15566 13949 15630
rect 14013 15566 14035 15630
rect 14099 15566 14121 15630
rect 14185 15566 14207 15630
rect 14271 15566 14293 15630
rect 14357 15566 14379 15630
rect 14443 15566 14465 15630
rect 14529 15566 14555 15630
rect 13769 15550 14555 15566
rect 13769 15486 13777 15550
rect 13841 15486 13863 15550
rect 13927 15486 13949 15550
rect 14013 15486 14035 15550
rect 14099 15486 14121 15550
rect 14185 15486 14207 15550
rect 14271 15486 14293 15550
rect 14357 15486 14379 15550
rect 14443 15486 14465 15550
rect 14529 15486 14555 15550
rect 13769 15470 14555 15486
rect 13769 15406 13777 15470
rect 13841 15406 13863 15470
rect 13927 15406 13949 15470
rect 14013 15406 14035 15470
rect 14099 15406 14121 15470
rect 14185 15406 14207 15470
rect 14271 15406 14293 15470
rect 14357 15406 14379 15470
rect 14443 15406 14465 15470
rect 14529 15406 14555 15470
rect 13769 15390 14555 15406
rect 13769 15326 13777 15390
rect 13841 15326 13863 15390
rect 13927 15326 13949 15390
rect 14013 15326 14035 15390
rect 14099 15326 14121 15390
rect 14185 15326 14207 15390
rect 14271 15326 14293 15390
rect 14357 15326 14379 15390
rect 14443 15326 14465 15390
rect 14529 15326 14555 15390
rect 13769 15310 14555 15326
rect 13769 15246 13777 15310
rect 13841 15246 13863 15310
rect 13927 15246 13949 15310
rect 14013 15246 14035 15310
rect 14099 15246 14121 15310
rect 14185 15246 14207 15310
rect 14271 15246 14293 15310
rect 14357 15246 14379 15310
rect 14443 15246 14465 15310
rect 14529 15246 14555 15310
rect 13769 15230 14555 15246
rect 13769 15166 13777 15230
rect 13841 15166 13863 15230
rect 13927 15166 13949 15230
rect 14013 15166 14035 15230
rect 14099 15166 14121 15230
rect 14185 15166 14207 15230
rect 14271 15166 14293 15230
rect 14357 15166 14379 15230
rect 14443 15166 14465 15230
rect 14529 15166 14555 15230
rect 13769 15149 14555 15166
rect 13769 15085 13777 15149
rect 13841 15085 13863 15149
rect 13927 15085 13949 15149
rect 14013 15085 14035 15149
rect 14099 15085 14121 15149
rect 14185 15085 14207 15149
rect 14271 15085 14293 15149
rect 14357 15085 14379 15149
rect 14443 15085 14465 15149
rect 14529 15085 14555 15149
rect 13769 15068 14555 15085
rect 13769 15004 13777 15068
rect 13841 15004 13863 15068
rect 13927 15004 13949 15068
rect 14013 15004 14035 15068
rect 14099 15004 14121 15068
rect 14185 15004 14207 15068
rect 14271 15004 14293 15068
rect 14357 15004 14379 15068
rect 14443 15004 14465 15068
rect 14529 15004 14555 15068
rect 13769 14987 14555 15004
rect 13769 14923 13777 14987
rect 13841 14923 13863 14987
rect 13927 14923 13949 14987
rect 14013 14923 14035 14987
rect 14099 14923 14121 14987
rect 14185 14923 14207 14987
rect 14271 14923 14293 14987
rect 14357 14923 14379 14987
rect 14443 14923 14465 14987
rect 14529 14923 14555 14987
rect 13769 14906 14555 14923
rect 13769 14842 13777 14906
rect 13841 14842 13863 14906
rect 13927 14842 13949 14906
rect 14013 14842 14035 14906
rect 14099 14842 14121 14906
rect 14185 14842 14207 14906
rect 14271 14842 14293 14906
rect 14357 14842 14379 14906
rect 14443 14842 14465 14906
rect 14529 14842 14555 14906
rect 13769 14825 14555 14842
rect 13769 14761 13777 14825
rect 13841 14761 13863 14825
rect 13927 14761 13949 14825
rect 14013 14761 14035 14825
rect 14099 14761 14121 14825
rect 14185 14761 14207 14825
rect 14271 14761 14293 14825
rect 14357 14761 14379 14825
rect 14443 14761 14465 14825
rect 14529 14761 14555 14825
rect 13769 14744 14555 14761
rect 13769 14680 13777 14744
rect 13841 14680 13863 14744
rect 13927 14680 13949 14744
rect 14013 14680 14035 14744
rect 14099 14680 14121 14744
rect 14185 14680 14207 14744
rect 14271 14680 14293 14744
rect 14357 14680 14379 14744
rect 14443 14680 14465 14744
rect 14529 14680 14555 14744
rect 13769 14663 14555 14680
rect 13769 14599 13777 14663
rect 13841 14599 13863 14663
rect 13927 14599 13949 14663
rect 14013 14599 14035 14663
rect 14099 14599 14121 14663
rect 14185 14599 14207 14663
rect 14271 14599 14293 14663
rect 14357 14599 14379 14663
rect 14443 14599 14465 14663
rect 14529 14599 14555 14663
rect 13769 14582 14555 14599
rect 13769 14518 13777 14582
rect 13841 14518 13863 14582
rect 13927 14518 13949 14582
rect 14013 14518 14035 14582
rect 14099 14518 14121 14582
rect 14185 14518 14207 14582
rect 14271 14518 14293 14582
rect 14357 14518 14379 14582
rect 14443 14518 14465 14582
rect 14529 14518 14555 14582
rect 13769 14501 14555 14518
rect 13769 14437 13777 14501
rect 13841 14437 13863 14501
rect 13927 14437 13949 14501
rect 14013 14437 14035 14501
rect 14099 14437 14121 14501
rect 14185 14437 14207 14501
rect 14271 14437 14293 14501
rect 14357 14437 14379 14501
rect 14443 14437 14465 14501
rect 14529 14437 14555 14501
rect 13769 14420 14555 14437
rect 13769 14356 13777 14420
rect 13841 14356 13863 14420
rect 13927 14356 13949 14420
rect 14013 14356 14035 14420
rect 14099 14356 14121 14420
rect 14185 14356 14207 14420
rect 14271 14356 14293 14420
rect 14357 14356 14379 14420
rect 14443 14356 14465 14420
rect 14529 14356 14555 14420
rect 13769 14339 14555 14356
rect 13769 14275 13777 14339
rect 13841 14275 13863 14339
rect 13927 14275 13949 14339
rect 14013 14275 14035 14339
rect 14099 14275 14121 14339
rect 14185 14275 14207 14339
rect 14271 14275 14293 14339
rect 14357 14275 14379 14339
rect 14443 14275 14465 14339
rect 14529 14275 14555 14339
rect 13769 14258 14555 14275
rect 13769 14194 13777 14258
rect 13841 14194 13863 14258
rect 13927 14194 13949 14258
rect 14013 14194 14035 14258
rect 14099 14194 14121 14258
rect 14185 14194 14207 14258
rect 14271 14194 14293 14258
rect 14357 14194 14379 14258
rect 14443 14194 14465 14258
rect 14529 14194 14555 14258
rect 13769 14177 14555 14194
rect 13769 14113 13777 14177
rect 13841 14113 13863 14177
rect 13927 14113 13949 14177
rect 14013 14113 14035 14177
rect 14099 14113 14121 14177
rect 14185 14113 14207 14177
rect 14271 14113 14293 14177
rect 14357 14113 14379 14177
rect 14443 14113 14465 14177
rect 14529 14113 14555 14177
rect 13769 14096 14555 14113
rect 13769 14032 13777 14096
rect 13841 14032 13863 14096
rect 13927 14032 13949 14096
rect 14013 14032 14035 14096
rect 14099 14032 14121 14096
rect 14185 14032 14207 14096
rect 14271 14032 14293 14096
rect 14357 14032 14379 14096
rect 14443 14032 14465 14096
rect 14529 14032 14555 14096
rect 13769 14015 14555 14032
rect 13769 13951 13777 14015
rect 13841 13951 13863 14015
rect 13927 13951 13949 14015
rect 14013 13951 14035 14015
rect 14099 13951 14121 14015
rect 14185 13951 14207 14015
rect 14271 13951 14293 14015
rect 14357 13951 14379 14015
rect 14443 13951 14465 14015
rect 14529 13951 14555 14015
rect 13769 13934 14555 13951
rect 13769 13870 13777 13934
rect 13841 13870 13863 13934
rect 13927 13870 13949 13934
rect 14013 13870 14035 13934
rect 14099 13870 14121 13934
rect 14185 13870 14207 13934
rect 14271 13870 14293 13934
rect 14357 13870 14379 13934
rect 14443 13870 14465 13934
rect 14529 13870 14555 13934
rect 13769 13853 14555 13870
rect 13769 13789 13777 13853
rect 13841 13789 13863 13853
rect 13927 13789 13949 13853
rect 14013 13789 14035 13853
rect 14099 13789 14121 13853
rect 14185 13789 14207 13853
rect 14271 13789 14293 13853
rect 14357 13789 14379 13853
rect 14443 13789 14465 13853
rect 14529 13789 14555 13853
rect 13769 13772 14555 13789
rect 13769 13708 13777 13772
rect 13841 13708 13863 13772
rect 13927 13708 13949 13772
rect 14013 13708 14035 13772
rect 14099 13708 14121 13772
rect 14185 13708 14207 13772
rect 14271 13708 14293 13772
rect 14357 13708 14379 13772
rect 14443 13708 14465 13772
rect 14529 13708 14555 13772
rect 13769 13691 14555 13708
rect 13769 13627 13777 13691
rect 13841 13627 13863 13691
rect 13927 13627 13949 13691
rect 14013 13627 14035 13691
rect 14099 13627 14121 13691
rect 14185 13627 14207 13691
rect 14271 13627 14293 13691
rect 14357 13627 14379 13691
rect 14443 13627 14465 13691
rect 14529 13627 14555 13691
rect 13769 13607 14555 13627
rect 1982 12398 8124 12887
tri 1982 12130 2250 12398 ne
rect 2250 12130 8124 12398
tri 2250 10485 3895 12130 ne
rect 3895 10485 6479 12130
tri 6479 10485 8124 12130 nw
tri 3895 10213 4167 10485 ne
rect 198 8841 1262 8850
rect 198 8785 203 8841
rect 259 8835 287 8841
rect 343 8835 371 8841
rect 427 8835 454 8841
rect 510 8835 537 8841
rect 593 8835 620 8841
rect 676 8835 703 8841
rect 759 8835 786 8841
rect 842 8835 869 8841
rect 925 8835 952 8841
rect 1008 8835 1035 8841
rect 1091 8835 1118 8841
rect 1174 8835 1201 8841
rect 198 8771 204 8785
rect 268 8771 287 8835
rect 351 8771 370 8835
rect 434 8771 453 8835
rect 517 8771 536 8835
rect 600 8771 618 8835
rect 682 8771 700 8835
rect 764 8771 782 8835
rect 846 8771 864 8835
rect 928 8771 946 8835
rect 1010 8771 1028 8835
rect 1092 8771 1110 8835
rect 1174 8771 1192 8835
rect 1257 8785 1262 8841
rect 1256 8771 1262 8785
rect 198 8755 1262 8771
rect 198 8699 203 8755
rect 259 8751 287 8755
rect 343 8751 371 8755
rect 427 8751 454 8755
rect 510 8751 537 8755
rect 593 8751 620 8755
rect 676 8751 703 8755
rect 759 8751 786 8755
rect 842 8751 869 8755
rect 925 8751 952 8755
rect 1008 8751 1035 8755
rect 1091 8751 1118 8755
rect 1174 8751 1201 8755
rect 198 8687 204 8699
rect 268 8687 287 8751
rect 351 8687 370 8751
rect 434 8687 453 8751
rect 517 8687 536 8751
rect 600 8687 618 8751
rect 682 8687 700 8751
rect 764 8687 782 8751
rect 846 8687 864 8751
rect 928 8687 946 8751
rect 1010 8687 1028 8751
rect 1092 8687 1110 8751
rect 1174 8687 1192 8751
rect 1257 8699 1262 8755
rect 1256 8687 1262 8699
rect 198 8669 1262 8687
rect 198 8613 203 8669
rect 259 8667 287 8669
rect 343 8667 371 8669
rect 427 8667 454 8669
rect 510 8667 537 8669
rect 593 8667 620 8669
rect 676 8667 703 8669
rect 759 8667 786 8669
rect 842 8667 869 8669
rect 925 8667 952 8669
rect 1008 8667 1035 8669
rect 1091 8667 1118 8669
rect 1174 8667 1201 8669
rect 198 8603 204 8613
rect 268 8603 287 8667
rect 351 8603 370 8667
rect 434 8603 453 8667
rect 517 8603 536 8667
rect 600 8603 618 8667
rect 682 8603 700 8667
rect 764 8603 782 8667
rect 846 8603 864 8667
rect 928 8603 946 8667
rect 1010 8603 1028 8667
rect 1092 8603 1110 8667
rect 1174 8603 1192 8667
rect 1257 8613 1262 8669
rect 1256 8603 1262 8613
rect 198 8583 1262 8603
rect 198 8527 203 8583
rect 198 8519 204 8527
rect 268 8519 287 8583
rect 351 8519 370 8583
rect 434 8519 453 8583
rect 517 8519 536 8583
rect 600 8519 618 8583
rect 682 8519 700 8583
rect 764 8519 782 8583
rect 846 8519 864 8583
rect 928 8519 946 8583
rect 1010 8519 1028 8583
rect 1092 8519 1110 8583
rect 1174 8519 1192 8583
rect 1257 8527 1262 8583
rect 1256 8519 1262 8527
rect 198 8499 1262 8519
rect 198 8497 204 8499
rect 198 8441 203 8497
rect 198 8435 204 8441
rect 268 8435 287 8499
rect 351 8435 370 8499
rect 434 8435 453 8499
rect 517 8435 536 8499
rect 600 8435 618 8499
rect 682 8435 700 8499
rect 764 8435 782 8499
rect 846 8435 864 8499
rect 928 8435 946 8499
rect 1010 8435 1028 8499
rect 1092 8435 1110 8499
rect 1174 8435 1192 8499
rect 1256 8497 1262 8499
rect 1257 8441 1262 8497
rect 1256 8435 1262 8441
rect 198 8415 1262 8435
rect 198 8411 204 8415
rect 198 8355 203 8411
rect 198 8351 204 8355
rect 268 8351 287 8415
rect 351 8351 370 8415
rect 434 8351 453 8415
rect 517 8351 536 8415
rect 600 8351 618 8415
rect 682 8351 700 8415
rect 764 8351 782 8415
rect 846 8351 864 8415
rect 928 8351 946 8415
rect 1010 8351 1028 8415
rect 1092 8351 1110 8415
rect 1174 8351 1192 8415
rect 1256 8411 1262 8415
rect 1257 8355 1262 8411
rect 1256 8351 1262 8355
rect 198 8331 1262 8351
rect 198 8325 204 8331
rect 198 8269 203 8325
rect 198 8267 204 8269
rect 268 8267 287 8331
rect 351 8267 370 8331
rect 434 8267 453 8331
rect 517 8267 536 8331
rect 600 8267 618 8331
rect 682 8267 700 8331
rect 764 8267 782 8331
rect 846 8267 864 8331
rect 928 8267 946 8331
rect 1010 8267 1028 8331
rect 1092 8267 1110 8331
rect 1174 8267 1192 8331
rect 1256 8325 1262 8331
rect 1257 8269 1262 8325
rect 1256 8267 1262 8269
rect 198 8247 1262 8267
rect 198 8239 204 8247
rect 198 8183 203 8239
rect 268 8183 287 8247
rect 351 8183 370 8247
rect 434 8183 453 8247
rect 517 8183 536 8247
rect 600 8183 618 8247
rect 682 8183 700 8247
rect 764 8183 782 8247
rect 846 8183 864 8247
rect 928 8183 946 8247
rect 1010 8183 1028 8247
rect 1092 8183 1110 8247
rect 1174 8183 1192 8247
rect 1256 8239 1262 8247
rect 1257 8183 1262 8239
rect 198 8163 1262 8183
rect 198 8153 204 8163
rect 198 8097 203 8153
rect 268 8099 287 8163
rect 351 8099 370 8163
rect 434 8099 453 8163
rect 517 8099 536 8163
rect 600 8099 618 8163
rect 682 8099 700 8163
rect 764 8099 782 8163
rect 846 8099 864 8163
rect 928 8099 946 8163
rect 1010 8099 1028 8163
rect 1092 8099 1110 8163
rect 1174 8099 1192 8163
rect 1256 8153 1262 8163
rect 259 8097 287 8099
rect 343 8097 371 8099
rect 427 8097 454 8099
rect 510 8097 537 8099
rect 593 8097 620 8099
rect 676 8097 703 8099
rect 759 8097 786 8099
rect 842 8097 869 8099
rect 925 8097 952 8099
rect 1008 8097 1035 8099
rect 1091 8097 1118 8099
rect 1174 8097 1201 8099
rect 1257 8097 1262 8153
rect 198 8079 1262 8097
rect 198 8067 204 8079
rect 198 8011 203 8067
rect 268 8015 287 8079
rect 351 8015 370 8079
rect 434 8015 453 8079
rect 517 8015 536 8079
rect 600 8015 618 8079
rect 682 8015 700 8079
rect 764 8015 782 8079
rect 846 8015 864 8079
rect 928 8015 946 8079
rect 1010 8015 1028 8079
rect 1092 8015 1110 8079
rect 1174 8015 1192 8079
rect 1256 8067 1262 8079
rect 259 8011 287 8015
rect 343 8011 371 8015
rect 427 8011 454 8015
rect 510 8011 537 8015
rect 593 8011 620 8015
rect 676 8011 703 8015
rect 759 8011 786 8015
rect 842 8011 869 8015
rect 925 8011 952 8015
rect 1008 8011 1035 8015
rect 1091 8011 1118 8015
rect 1174 8011 1201 8015
rect 1257 8011 1262 8067
rect 198 7995 1262 8011
rect 198 7981 204 7995
rect 198 7925 203 7981
rect 268 7931 287 7995
rect 351 7931 370 7995
rect 434 7931 453 7995
rect 517 7931 536 7995
rect 600 7931 618 7995
rect 682 7931 700 7995
rect 764 7931 782 7995
rect 846 7931 864 7995
rect 928 7931 946 7995
rect 1010 7931 1028 7995
rect 1092 7931 1110 7995
rect 1174 7931 1192 7995
rect 1256 7981 1262 7995
rect 259 7925 287 7931
rect 343 7925 371 7931
rect 427 7925 454 7931
rect 510 7925 537 7931
rect 593 7925 620 7931
rect 676 7925 703 7931
rect 759 7925 786 7931
rect 842 7925 869 7931
rect 925 7925 952 7931
rect 1008 7925 1035 7931
rect 1091 7925 1118 7931
rect 1174 7925 1201 7931
rect 1257 7925 1262 7981
rect 198 7916 1262 7925
rect 4167 6863 6479 10485
rect 8198 8841 9261 8850
rect 8198 8785 8203 8841
rect 8259 8829 8287 8841
rect 8343 8829 8370 8841
rect 8426 8829 8453 8841
rect 8509 8829 8536 8841
rect 8592 8829 8619 8841
rect 8675 8829 8702 8841
rect 8758 8829 8785 8841
rect 8841 8829 8868 8841
rect 8924 8829 8951 8841
rect 9007 8829 9034 8841
rect 9090 8829 9117 8841
rect 9173 8829 9200 8841
rect 8369 8785 8370 8829
rect 8450 8785 8453 8829
rect 8530 8785 8536 8829
rect 8610 8785 8619 8829
rect 8690 8785 8702 8829
rect 8770 8785 8785 8829
rect 8198 8765 8224 8785
rect 8288 8765 8305 8785
rect 8369 8765 8386 8785
rect 8450 8765 8466 8785
rect 8530 8765 8546 8785
rect 8610 8765 8626 8785
rect 8690 8765 8706 8785
rect 8770 8765 8786 8785
rect 8850 8765 8866 8829
rect 8930 8765 8946 8829
rect 9010 8765 9026 8829
rect 9090 8765 9106 8829
rect 9173 8785 9186 8829
rect 9256 8785 9261 8841
rect 9170 8765 9186 8785
rect 9250 8765 9261 8785
rect 8198 8755 9261 8765
rect 8198 8699 8203 8755
rect 8259 8745 8287 8755
rect 8343 8745 8370 8755
rect 8426 8745 8453 8755
rect 8509 8745 8536 8755
rect 8592 8745 8619 8755
rect 8675 8745 8702 8755
rect 8758 8745 8785 8755
rect 8841 8745 8868 8755
rect 8924 8745 8951 8755
rect 9007 8745 9034 8755
rect 9090 8745 9117 8755
rect 9173 8745 9200 8755
rect 8369 8699 8370 8745
rect 8450 8699 8453 8745
rect 8530 8699 8536 8745
rect 8610 8699 8619 8745
rect 8690 8699 8702 8745
rect 8770 8699 8785 8745
rect 8198 8681 8224 8699
rect 8288 8681 8305 8699
rect 8369 8681 8386 8699
rect 8450 8681 8466 8699
rect 8530 8681 8546 8699
rect 8610 8681 8626 8699
rect 8690 8681 8706 8699
rect 8770 8681 8786 8699
rect 8850 8681 8866 8745
rect 8930 8681 8946 8745
rect 9010 8681 9026 8745
rect 9090 8681 9106 8745
rect 9173 8699 9186 8745
rect 9256 8699 9261 8755
rect 9170 8681 9186 8699
rect 9250 8681 9261 8699
rect 8198 8669 9261 8681
rect 8198 8613 8203 8669
rect 8259 8661 8287 8669
rect 8343 8661 8370 8669
rect 8426 8661 8453 8669
rect 8509 8661 8536 8669
rect 8592 8661 8619 8669
rect 8675 8661 8702 8669
rect 8758 8661 8785 8669
rect 8841 8661 8868 8669
rect 8924 8661 8951 8669
rect 9007 8661 9034 8669
rect 9090 8661 9117 8669
rect 9173 8661 9200 8669
rect 8369 8613 8370 8661
rect 8450 8613 8453 8661
rect 8530 8613 8536 8661
rect 8610 8613 8619 8661
rect 8690 8613 8702 8661
rect 8770 8613 8785 8661
rect 8198 8597 8224 8613
rect 8288 8597 8305 8613
rect 8369 8597 8386 8613
rect 8450 8597 8466 8613
rect 8530 8597 8546 8613
rect 8610 8597 8626 8613
rect 8690 8597 8706 8613
rect 8770 8597 8786 8613
rect 8850 8597 8866 8661
rect 8930 8597 8946 8661
rect 9010 8597 9026 8661
rect 9090 8597 9106 8661
rect 9173 8613 9186 8661
rect 9256 8613 9261 8669
rect 9170 8597 9186 8613
rect 9250 8597 9261 8613
rect 8198 8583 9261 8597
rect 8198 8527 8203 8583
rect 8259 8577 8287 8583
rect 8343 8577 8370 8583
rect 8426 8577 8453 8583
rect 8509 8577 8536 8583
rect 8592 8577 8619 8583
rect 8675 8577 8702 8583
rect 8758 8577 8785 8583
rect 8841 8577 8868 8583
rect 8924 8577 8951 8583
rect 9007 8577 9034 8583
rect 9090 8577 9117 8583
rect 9173 8577 9200 8583
rect 8369 8527 8370 8577
rect 8450 8527 8453 8577
rect 8530 8527 8536 8577
rect 8610 8527 8619 8577
rect 8690 8527 8702 8577
rect 8770 8527 8785 8577
rect 8198 8513 8224 8527
rect 8288 8513 8305 8527
rect 8369 8513 8386 8527
rect 8450 8513 8466 8527
rect 8530 8513 8546 8527
rect 8610 8513 8626 8527
rect 8690 8513 8706 8527
rect 8770 8513 8786 8527
rect 8850 8513 8866 8577
rect 8930 8513 8946 8577
rect 9010 8513 9026 8577
rect 9090 8513 9106 8577
rect 9173 8527 9186 8577
rect 9256 8527 9261 8583
rect 9170 8513 9186 8527
rect 9250 8513 9261 8527
rect 8198 8497 9261 8513
rect 8198 8441 8203 8497
rect 8259 8493 8287 8497
rect 8343 8493 8370 8497
rect 8426 8493 8453 8497
rect 8509 8493 8536 8497
rect 8592 8493 8619 8497
rect 8675 8493 8702 8497
rect 8758 8493 8785 8497
rect 8841 8493 8868 8497
rect 8924 8493 8951 8497
rect 9007 8493 9034 8497
rect 9090 8493 9117 8497
rect 9173 8493 9200 8497
rect 8369 8441 8370 8493
rect 8450 8441 8453 8493
rect 8530 8441 8536 8493
rect 8610 8441 8619 8493
rect 8690 8441 8702 8493
rect 8770 8441 8785 8493
rect 8198 8429 8224 8441
rect 8288 8429 8305 8441
rect 8369 8429 8386 8441
rect 8450 8429 8466 8441
rect 8530 8429 8546 8441
rect 8610 8429 8626 8441
rect 8690 8429 8706 8441
rect 8770 8429 8786 8441
rect 8850 8429 8866 8493
rect 8930 8429 8946 8493
rect 9010 8429 9026 8493
rect 9090 8429 9106 8493
rect 9173 8441 9186 8493
rect 9256 8441 9261 8497
rect 9170 8429 9186 8441
rect 9250 8429 9261 8441
rect 8198 8411 9261 8429
rect 8198 8355 8203 8411
rect 8259 8409 8287 8411
rect 8343 8409 8370 8411
rect 8426 8409 8453 8411
rect 8509 8409 8536 8411
rect 8592 8409 8619 8411
rect 8675 8409 8702 8411
rect 8758 8409 8785 8411
rect 8841 8409 8868 8411
rect 8924 8409 8951 8411
rect 9007 8409 9034 8411
rect 9090 8409 9117 8411
rect 9173 8409 9200 8411
rect 8369 8355 8370 8409
rect 8450 8355 8453 8409
rect 8530 8355 8536 8409
rect 8610 8355 8619 8409
rect 8690 8355 8702 8409
rect 8770 8355 8785 8409
rect 8198 8345 8224 8355
rect 8288 8345 8305 8355
rect 8369 8345 8386 8355
rect 8450 8345 8466 8355
rect 8530 8345 8546 8355
rect 8610 8345 8626 8355
rect 8690 8345 8706 8355
rect 8770 8345 8786 8355
rect 8850 8345 8866 8409
rect 8930 8345 8946 8409
rect 9010 8345 9026 8409
rect 9090 8345 9106 8409
rect 9173 8355 9186 8409
rect 9256 8355 9261 8411
rect 9170 8345 9186 8355
rect 9250 8345 9261 8355
rect 8198 8325 9261 8345
rect 8198 8269 8203 8325
rect 8369 8269 8370 8325
rect 8450 8269 8453 8325
rect 8530 8269 8536 8325
rect 8610 8269 8619 8325
rect 8690 8269 8702 8325
rect 8770 8269 8785 8325
rect 8198 8261 8224 8269
rect 8288 8261 8305 8269
rect 8369 8261 8386 8269
rect 8450 8261 8466 8269
rect 8530 8261 8546 8269
rect 8610 8261 8626 8269
rect 8690 8261 8706 8269
rect 8770 8261 8786 8269
rect 8850 8261 8866 8325
rect 8930 8261 8946 8325
rect 9010 8261 9026 8325
rect 9090 8261 9106 8325
rect 9173 8269 9186 8325
rect 9256 8269 9261 8325
rect 9170 8261 9186 8269
rect 9250 8261 9261 8269
rect 8198 8241 9261 8261
rect 8198 8239 8224 8241
rect 8288 8239 8305 8241
rect 8369 8239 8386 8241
rect 8450 8239 8466 8241
rect 8530 8239 8546 8241
rect 8610 8239 8626 8241
rect 8690 8239 8706 8241
rect 8770 8239 8786 8241
rect 8198 8183 8203 8239
rect 8369 8183 8370 8239
rect 8450 8183 8453 8239
rect 8530 8183 8536 8239
rect 8610 8183 8619 8239
rect 8690 8183 8702 8239
rect 8770 8183 8785 8239
rect 8198 8177 8224 8183
rect 8288 8177 8305 8183
rect 8369 8177 8386 8183
rect 8450 8177 8466 8183
rect 8530 8177 8546 8183
rect 8610 8177 8626 8183
rect 8690 8177 8706 8183
rect 8770 8177 8786 8183
rect 8850 8177 8866 8241
rect 8930 8177 8946 8241
rect 9010 8177 9026 8241
rect 9090 8177 9106 8241
rect 9170 8239 9186 8241
rect 9250 8239 9261 8241
rect 9173 8183 9186 8239
rect 9256 8183 9261 8239
rect 9170 8177 9186 8183
rect 9250 8177 9261 8183
rect 8198 8157 9261 8177
rect 8198 8153 8224 8157
rect 8288 8153 8305 8157
rect 8369 8153 8386 8157
rect 8450 8153 8466 8157
rect 8530 8153 8546 8157
rect 8610 8153 8626 8157
rect 8690 8153 8706 8157
rect 8770 8153 8786 8157
rect 8198 8097 8203 8153
rect 8369 8097 8370 8153
rect 8450 8097 8453 8153
rect 8530 8097 8536 8153
rect 8610 8097 8619 8153
rect 8690 8097 8702 8153
rect 8770 8097 8785 8153
rect 8198 8093 8224 8097
rect 8288 8093 8305 8097
rect 8369 8093 8386 8097
rect 8450 8093 8466 8097
rect 8530 8093 8546 8097
rect 8610 8093 8626 8097
rect 8690 8093 8706 8097
rect 8770 8093 8786 8097
rect 8850 8093 8866 8157
rect 8930 8093 8946 8157
rect 9010 8093 9026 8157
rect 9090 8093 9106 8157
rect 9170 8153 9186 8157
rect 9250 8153 9261 8157
rect 9173 8097 9186 8153
rect 9256 8097 9261 8153
rect 9170 8093 9186 8097
rect 9250 8093 9261 8097
rect 8198 8073 9261 8093
rect 8198 8067 8224 8073
rect 8288 8067 8305 8073
rect 8369 8067 8386 8073
rect 8450 8067 8466 8073
rect 8530 8067 8546 8073
rect 8610 8067 8626 8073
rect 8690 8067 8706 8073
rect 8770 8067 8786 8073
rect 8198 8011 8203 8067
rect 8369 8011 8370 8067
rect 8450 8011 8453 8067
rect 8530 8011 8536 8067
rect 8610 8011 8619 8067
rect 8690 8011 8702 8067
rect 8770 8011 8785 8067
rect 8198 8009 8224 8011
rect 8288 8009 8305 8011
rect 8369 8009 8386 8011
rect 8450 8009 8466 8011
rect 8530 8009 8546 8011
rect 8610 8009 8626 8011
rect 8690 8009 8706 8011
rect 8770 8009 8786 8011
rect 8850 8009 8866 8073
rect 8930 8009 8946 8073
rect 9010 8009 9026 8073
rect 9090 8009 9106 8073
rect 9170 8067 9186 8073
rect 9250 8067 9261 8073
rect 9173 8011 9186 8067
rect 9256 8011 9261 8067
rect 9170 8009 9186 8011
rect 9250 8009 9261 8011
rect 8198 7989 9261 8009
rect 8198 7981 8224 7989
rect 8288 7981 8305 7989
rect 8369 7981 8386 7989
rect 8450 7981 8466 7989
rect 8530 7981 8546 7989
rect 8610 7981 8626 7989
rect 8690 7981 8706 7989
rect 8770 7981 8786 7989
rect 8198 7925 8203 7981
rect 8369 7925 8370 7981
rect 8450 7925 8453 7981
rect 8530 7925 8536 7981
rect 8610 7925 8619 7981
rect 8690 7925 8702 7981
rect 8770 7925 8785 7981
rect 8850 7925 8866 7989
rect 8930 7925 8946 7989
rect 9010 7925 9026 7989
rect 9090 7925 9106 7989
rect 9170 7981 9186 7989
rect 9250 7981 9261 7989
rect 9173 7925 9186 7981
rect 9256 7925 9261 7981
rect 8198 7916 9261 7925
tri 4167 6548 4482 6863 ne
rect 4482 6548 6479 6863
tri 6479 6548 7022 7091 sw
tri 4482 4551 6479 6548 ne
rect 6479 4551 7022 6548
tri 6479 4008 7022 4551 ne
tri 7022 4008 9562 6548 sw
tri 7022 3264 7766 4008 ne
rect 7766 3014 9562 4008
rect 7766 0 9562 2834
<< rmetal3 >>
rect 7766 2834 9562 3014
<< via3 >>
rect 462 39528 526 39592
rect 620 39528 684 39592
rect 462 39448 526 39512
rect 620 39448 684 39512
rect 462 39368 526 39432
rect 620 39368 684 39432
rect 462 39288 526 39352
rect 620 39288 684 39352
rect 462 39208 526 39272
rect 620 39208 684 39272
rect 462 39128 526 39192
rect 620 39128 684 39192
rect 462 39048 526 39112
rect 620 39048 684 39112
rect 462 38968 526 39032
rect 620 38968 684 39032
rect 462 38888 526 38952
rect 620 38888 684 38952
rect 462 38808 526 38872
rect 620 38808 684 38872
rect 462 38728 526 38792
rect 620 38728 684 38792
rect 462 38648 526 38712
rect 620 38648 684 38712
rect 462 38568 526 38632
rect 620 38568 684 38632
rect 462 38488 526 38552
rect 620 38488 684 38552
rect 462 38408 526 38472
rect 620 38408 684 38472
rect 462 38328 526 38392
rect 620 38328 684 38392
rect 462 38247 526 38311
rect 620 38247 684 38311
rect 462 38166 526 38230
rect 620 38166 684 38230
rect 462 38085 526 38149
rect 620 38085 684 38149
rect 462 38004 526 38068
rect 620 38004 684 38068
rect 462 37923 526 37987
rect 620 37923 684 37987
rect 462 37842 526 37906
rect 620 37842 684 37906
rect 462 37761 526 37825
rect 620 37761 684 37825
rect 462 37680 526 37744
rect 620 37680 684 37744
rect 462 37599 526 37663
rect 620 37599 684 37663
rect 462 37518 526 37582
rect 620 37518 684 37582
rect 462 37437 526 37501
rect 620 37437 684 37501
rect 462 37356 526 37420
rect 620 37356 684 37420
rect 462 37275 526 37339
rect 620 37275 684 37339
rect 462 37194 526 37258
rect 620 37194 684 37258
rect 462 37113 526 37177
rect 620 37113 684 37177
rect 462 37032 526 37096
rect 620 37032 684 37096
rect 462 36951 526 37015
rect 620 36951 684 37015
rect 462 36870 526 36934
rect 620 36870 684 36934
rect 462 36789 526 36853
rect 620 36789 684 36853
rect 462 36708 526 36772
rect 620 36708 684 36772
rect 462 36627 526 36691
rect 620 36627 684 36691
rect 462 36546 526 36610
rect 620 36546 684 36610
rect 462 36465 526 36529
rect 620 36465 684 36529
rect 462 36384 526 36448
rect 620 36384 684 36448
rect 462 36303 526 36367
rect 620 36303 684 36367
rect 462 36222 526 36286
rect 620 36222 684 36286
rect 462 36141 526 36205
rect 620 36141 684 36205
rect 462 36060 526 36124
rect 620 36060 684 36124
rect 462 35979 526 36043
rect 620 35979 684 36043
rect 462 35898 526 35962
rect 620 35898 684 35962
rect 462 35817 526 35881
rect 620 35817 684 35881
rect 462 35736 526 35800
rect 620 35736 684 35800
rect 462 35655 526 35719
rect 620 35655 684 35719
rect 462 35574 526 35638
rect 620 35574 684 35638
rect 462 35493 526 35557
rect 620 35493 684 35557
rect 462 35412 526 35476
rect 620 35412 684 35476
rect 462 35331 526 35395
rect 620 35331 684 35395
rect 462 35250 526 35314
rect 620 35250 684 35314
rect 462 35169 526 35233
rect 620 35169 684 35233
rect 462 35088 526 35152
rect 620 35088 684 35152
rect 462 35007 526 35071
rect 620 35007 684 35071
rect 462 34926 526 34990
rect 620 34926 684 34990
rect 462 34845 526 34909
rect 620 34845 684 34909
rect 462 34764 526 34828
rect 620 34764 684 34828
rect 1390 39528 1454 39592
rect 1518 39528 1582 39592
rect 1390 39448 1454 39512
rect 1518 39448 1582 39512
rect 1390 39368 1454 39432
rect 1518 39368 1582 39432
rect 1390 39288 1454 39352
rect 1518 39288 1582 39352
rect 1390 39208 1454 39272
rect 1518 39208 1582 39272
rect 1390 39128 1454 39192
rect 1518 39128 1582 39192
rect 1390 39048 1454 39112
rect 1518 39048 1582 39112
rect 1390 38968 1454 39032
rect 1518 38968 1582 39032
rect 1390 38888 1454 38952
rect 1518 38888 1582 38952
rect 1390 38808 1454 38872
rect 1518 38808 1582 38872
rect 1390 38728 1454 38792
rect 1518 38728 1582 38792
rect 1390 38648 1454 38712
rect 1518 38648 1582 38712
rect 1390 38568 1454 38632
rect 1518 38568 1582 38632
rect 1390 38488 1454 38552
rect 1518 38488 1582 38552
rect 1390 38408 1454 38472
rect 1518 38408 1582 38472
rect 1390 38328 1454 38392
rect 1518 38328 1582 38392
rect 1390 38247 1454 38311
rect 1518 38247 1582 38311
rect 1390 38166 1454 38230
rect 1518 38166 1582 38230
rect 1390 38085 1454 38149
rect 1518 38085 1582 38149
rect 1390 38004 1454 38068
rect 1518 38004 1582 38068
rect 1390 37923 1454 37987
rect 1518 37923 1582 37987
rect 1390 37842 1454 37906
rect 1518 37842 1582 37906
rect 1390 37761 1454 37825
rect 1518 37761 1582 37825
rect 1390 37680 1454 37744
rect 1518 37680 1582 37744
rect 1390 37599 1454 37663
rect 1518 37599 1582 37663
rect 1390 37518 1454 37582
rect 1518 37518 1582 37582
rect 1390 37437 1454 37501
rect 1518 37437 1582 37501
rect 1390 37356 1454 37420
rect 1518 37356 1582 37420
rect 1390 37275 1454 37339
rect 1518 37275 1582 37339
rect 1390 37194 1454 37258
rect 1518 37194 1582 37258
rect 1390 37113 1454 37177
rect 1518 37113 1582 37177
rect 1390 37032 1454 37096
rect 1518 37032 1582 37096
rect 1390 36951 1454 37015
rect 1518 36951 1582 37015
rect 1390 36870 1454 36934
rect 1518 36870 1582 36934
rect 1390 36789 1454 36853
rect 1518 36789 1582 36853
rect 1390 36708 1454 36772
rect 1518 36708 1582 36772
rect 1390 36627 1454 36691
rect 1518 36627 1582 36691
rect 1390 36546 1454 36610
rect 1518 36546 1582 36610
rect 1390 36465 1454 36529
rect 1518 36465 1582 36529
rect 1390 36384 1454 36448
rect 1518 36384 1582 36448
rect 1390 36303 1454 36367
rect 1518 36303 1582 36367
rect 1390 36222 1454 36286
rect 1518 36222 1582 36286
rect 1390 36141 1454 36205
rect 1518 36141 1582 36205
rect 1390 36060 1454 36124
rect 1518 36060 1582 36124
rect 1390 35979 1454 36043
rect 1518 35979 1582 36043
rect 1390 35898 1454 35962
rect 1518 35898 1582 35962
rect 1390 35817 1454 35881
rect 1518 35817 1582 35881
rect 1390 35736 1454 35800
rect 1518 35736 1582 35800
rect 1390 35655 1454 35719
rect 1518 35655 1582 35719
rect 1390 35574 1454 35638
rect 1518 35574 1582 35638
rect 1390 35493 1454 35557
rect 1518 35493 1582 35557
rect 1390 35412 1454 35476
rect 1518 35412 1582 35476
rect 1390 35331 1454 35395
rect 1518 35331 1582 35395
rect 1390 35250 1454 35314
rect 1518 35250 1582 35314
rect 1390 35169 1454 35233
rect 1518 35169 1582 35233
rect 1390 35088 1454 35152
rect 1518 35088 1582 35152
rect 1390 35007 1454 35071
rect 1518 35007 1582 35071
rect 1390 34926 1454 34990
rect 1518 34926 1582 34990
rect 1390 34845 1454 34909
rect 1518 34845 1582 34909
rect 1390 34764 1454 34828
rect 1518 34764 1582 34828
rect 862 31962 918 32017
rect 918 31962 926 32017
rect 862 31953 926 31962
rect 990 31962 996 32017
rect 996 31962 1052 32017
rect 1052 31962 1054 32017
rect 990 31953 1054 31962
rect 862 31880 918 31936
rect 918 31880 926 31936
rect 862 31872 926 31880
rect 990 31880 996 31936
rect 996 31880 1052 31936
rect 1052 31880 1054 31936
rect 990 31872 1054 31880
rect 862 31854 926 31855
rect 862 31798 918 31854
rect 918 31798 926 31854
rect 862 31791 926 31798
rect 990 31854 1054 31855
rect 990 31798 996 31854
rect 996 31798 1052 31854
rect 1052 31798 1054 31854
rect 990 31791 1054 31798
rect 862 31772 926 31774
rect 862 31716 918 31772
rect 918 31716 926 31772
rect 862 31710 926 31716
rect 990 31772 1054 31774
rect 990 31716 996 31772
rect 996 31716 1052 31772
rect 1052 31716 1054 31772
rect 990 31710 1054 31716
rect 862 31690 926 31693
rect 862 31634 918 31690
rect 918 31634 926 31690
rect 862 31629 926 31634
rect 990 31690 1054 31693
rect 990 31634 996 31690
rect 996 31634 1052 31690
rect 1052 31634 1054 31690
rect 990 31629 1054 31634
rect 862 31608 926 31612
rect 862 31552 918 31608
rect 918 31552 926 31608
rect 862 31548 926 31552
rect 990 31608 1054 31612
rect 990 31552 996 31608
rect 996 31552 1052 31608
rect 1052 31552 1054 31608
rect 990 31548 1054 31552
rect 862 31526 926 31531
rect 862 31470 918 31526
rect 918 31470 926 31526
rect 862 31467 926 31470
rect 990 31526 1054 31531
rect 990 31470 996 31526
rect 996 31470 1052 31526
rect 1052 31470 1054 31526
rect 990 31467 1054 31470
rect 862 31444 926 31450
rect 862 31388 918 31444
rect 918 31388 926 31444
rect 862 31386 926 31388
rect 990 31444 1054 31450
rect 990 31388 996 31444
rect 996 31388 1052 31444
rect 1052 31388 1054 31444
rect 990 31386 1054 31388
rect 862 31362 926 31369
rect 862 31306 918 31362
rect 918 31306 926 31362
rect 862 31305 926 31306
rect 990 31362 1054 31369
rect 990 31306 996 31362
rect 996 31306 1052 31362
rect 1052 31306 1054 31362
rect 990 31305 1054 31306
rect 862 31280 926 31288
rect 862 31224 918 31280
rect 918 31224 926 31280
rect 990 31280 1054 31288
rect 990 31224 996 31280
rect 996 31224 1052 31280
rect 1052 31224 1054 31280
rect 862 31198 926 31207
rect 862 31143 918 31198
rect 918 31143 926 31198
rect 990 31198 1054 31207
rect 990 31143 996 31198
rect 996 31143 1052 31198
rect 1052 31143 1054 31198
rect 862 31116 926 31125
rect 862 31061 918 31116
rect 918 31061 926 31116
rect 990 31116 1054 31125
rect 990 31061 996 31116
rect 996 31061 1052 31116
rect 1052 31061 1054 31116
rect 862 31034 926 31043
rect 862 30979 918 31034
rect 918 30979 926 31034
rect 990 31034 1054 31043
rect 990 30979 996 31034
rect 996 30979 1052 31034
rect 1052 30979 1054 31034
rect 862 30952 926 30961
rect 862 30897 918 30952
rect 918 30897 926 30952
rect 990 30952 1054 30961
rect 990 30897 996 30952
rect 996 30897 1052 30952
rect 1052 30897 1054 30952
rect 862 30870 926 30879
rect 862 30815 918 30870
rect 918 30815 926 30870
rect 990 30870 1054 30879
rect 990 30815 996 30870
rect 996 30815 1052 30870
rect 1052 30815 1054 30870
rect 862 30788 926 30797
rect 862 30733 918 30788
rect 918 30733 926 30788
rect 990 30788 1054 30797
rect 990 30733 996 30788
rect 996 30733 1052 30788
rect 1052 30733 1054 30788
rect 862 30706 926 30715
rect 862 30651 918 30706
rect 918 30651 926 30706
rect 990 30706 1054 30715
rect 990 30651 996 30706
rect 996 30651 1052 30706
rect 1052 30651 1054 30706
rect 862 30624 926 30633
rect 862 30569 918 30624
rect 918 30569 926 30624
rect 990 30624 1054 30633
rect 990 30569 996 30624
rect 996 30569 1052 30624
rect 1052 30569 1054 30624
rect 862 30542 926 30551
rect 862 30487 918 30542
rect 918 30487 926 30542
rect 990 30542 1054 30551
rect 990 30487 996 30542
rect 996 30487 1052 30542
rect 1052 30487 1054 30542
rect 862 30460 926 30469
rect 862 30405 918 30460
rect 918 30405 926 30460
rect 990 30460 1054 30469
rect 990 30405 996 30460
rect 996 30405 1052 30460
rect 1052 30405 1054 30460
rect 862 30378 926 30387
rect 862 30323 918 30378
rect 918 30323 926 30378
rect 990 30378 1054 30387
rect 990 30323 996 30378
rect 996 30323 1052 30378
rect 1052 30323 1054 30378
rect 862 30296 926 30305
rect 862 30241 918 30296
rect 918 30241 926 30296
rect 990 30296 1054 30305
rect 990 30241 996 30296
rect 996 30241 1052 30296
rect 1052 30241 1054 30296
rect 862 30214 926 30223
rect 862 30159 918 30214
rect 918 30159 926 30214
rect 990 30214 1054 30223
rect 990 30159 996 30214
rect 996 30159 1052 30214
rect 1052 30159 1054 30214
rect 862 30132 926 30141
rect 862 30077 918 30132
rect 918 30077 926 30132
rect 990 30132 1054 30141
rect 990 30077 996 30132
rect 996 30077 1052 30132
rect 1052 30077 1054 30132
rect 862 30050 926 30059
rect 862 29995 918 30050
rect 918 29995 926 30050
rect 990 30050 1054 30059
rect 990 29995 996 30050
rect 996 29995 1052 30050
rect 1052 29995 1054 30050
rect 862 29968 926 29977
rect 862 29913 918 29968
rect 918 29913 926 29968
rect 990 29968 1054 29977
rect 990 29913 996 29968
rect 996 29913 1052 29968
rect 1052 29913 1054 29968
rect 862 29886 926 29895
rect 862 29831 918 29886
rect 918 29831 926 29886
rect 990 29886 1054 29895
rect 990 29831 996 29886
rect 996 29831 1052 29886
rect 1052 29831 1054 29886
rect 862 29804 926 29813
rect 862 29749 918 29804
rect 918 29749 926 29804
rect 990 29804 1054 29813
rect 990 29749 996 29804
rect 996 29749 1052 29804
rect 1052 29749 1054 29804
rect 862 29722 926 29731
rect 862 29667 918 29722
rect 918 29667 926 29722
rect 990 29722 1054 29731
rect 990 29667 996 29722
rect 996 29667 1052 29722
rect 1052 29667 1054 29722
rect 862 29640 926 29649
rect 862 29585 918 29640
rect 918 29585 926 29640
rect 990 29640 1054 29649
rect 990 29585 996 29640
rect 996 29585 1052 29640
rect 1052 29585 1054 29640
rect 862 29558 926 29567
rect 862 29503 918 29558
rect 918 29503 926 29558
rect 990 29558 1054 29567
rect 990 29503 996 29558
rect 996 29503 1052 29558
rect 1052 29503 1054 29558
rect 862 29476 926 29485
rect 862 29421 918 29476
rect 918 29421 926 29476
rect 990 29476 1054 29485
rect 990 29421 996 29476
rect 996 29421 1052 29476
rect 1052 29421 1054 29476
rect 2382 39528 2446 39592
rect 2510 39528 2574 39592
rect 2382 39448 2446 39512
rect 2510 39448 2574 39512
rect 2382 39368 2446 39432
rect 2510 39368 2574 39432
rect 2382 39288 2446 39352
rect 2510 39288 2574 39352
rect 2382 39208 2446 39272
rect 2510 39208 2574 39272
rect 2382 39128 2446 39192
rect 2510 39128 2574 39192
rect 2382 39048 2446 39112
rect 2510 39048 2574 39112
rect 2382 38968 2446 39032
rect 2510 38968 2574 39032
rect 2382 38888 2446 38952
rect 2510 38888 2574 38952
rect 2382 38808 2446 38872
rect 2510 38808 2574 38872
rect 2382 38728 2446 38792
rect 2510 38728 2574 38792
rect 2382 38648 2446 38712
rect 2510 38648 2574 38712
rect 2382 38568 2446 38632
rect 2510 38568 2574 38632
rect 2382 38488 2446 38552
rect 2510 38488 2574 38552
rect 2382 38408 2446 38472
rect 2510 38408 2574 38472
rect 2382 38328 2446 38392
rect 2510 38328 2574 38392
rect 2382 38247 2446 38311
rect 2510 38247 2574 38311
rect 2382 38166 2446 38230
rect 2510 38166 2574 38230
rect 2382 38085 2446 38149
rect 2510 38085 2574 38149
rect 2382 38004 2446 38068
rect 2510 38004 2574 38068
rect 2382 37923 2446 37987
rect 2510 37923 2574 37987
rect 2382 37842 2446 37906
rect 2510 37842 2574 37906
rect 2382 37761 2446 37825
rect 2510 37761 2574 37825
rect 2382 37680 2446 37744
rect 2510 37680 2574 37744
rect 2382 37599 2446 37663
rect 2510 37599 2574 37663
rect 2382 37518 2446 37582
rect 2510 37518 2574 37582
rect 2382 37437 2446 37501
rect 2510 37437 2574 37501
rect 2382 37356 2446 37420
rect 2510 37356 2574 37420
rect 2382 37275 2446 37339
rect 2510 37275 2574 37339
rect 2382 37194 2446 37258
rect 2510 37194 2574 37258
rect 2382 37113 2446 37177
rect 2510 37113 2574 37177
rect 2382 37032 2446 37096
rect 2510 37032 2574 37096
rect 2382 36951 2446 37015
rect 2510 36951 2574 37015
rect 2382 36870 2446 36934
rect 2510 36870 2574 36934
rect 2382 36789 2446 36853
rect 2510 36789 2574 36853
rect 2382 36708 2446 36772
rect 2510 36708 2574 36772
rect 2382 36627 2446 36691
rect 2510 36627 2574 36691
rect 2382 36546 2446 36610
rect 2510 36546 2574 36610
rect 2382 36465 2446 36529
rect 2510 36465 2574 36529
rect 2382 36384 2446 36448
rect 2510 36384 2574 36448
rect 2382 36303 2446 36367
rect 2510 36303 2574 36367
rect 2382 36222 2446 36286
rect 2510 36222 2574 36286
rect 2382 36141 2446 36205
rect 2510 36141 2574 36205
rect 2382 36060 2446 36124
rect 2510 36060 2574 36124
rect 2382 35979 2446 36043
rect 2510 35979 2574 36043
rect 2382 35898 2446 35962
rect 2510 35898 2574 35962
rect 2382 35817 2446 35881
rect 2510 35817 2574 35881
rect 2382 35736 2446 35800
rect 2510 35736 2574 35800
rect 2382 35655 2446 35719
rect 2510 35655 2574 35719
rect 2382 35574 2446 35638
rect 2510 35574 2574 35638
rect 2382 35493 2446 35557
rect 2510 35493 2574 35557
rect 2382 35412 2446 35476
rect 2510 35412 2574 35476
rect 2382 35331 2446 35395
rect 2510 35331 2574 35395
rect 2382 35250 2446 35314
rect 2510 35250 2574 35314
rect 2382 35169 2446 35233
rect 2510 35169 2574 35233
rect 2382 35088 2446 35152
rect 2510 35088 2574 35152
rect 2382 35007 2446 35071
rect 2510 35007 2574 35071
rect 2382 34926 2446 34990
rect 2510 34926 2574 34990
rect 2382 34845 2446 34909
rect 2510 34845 2574 34909
rect 2382 34764 2446 34828
rect 2510 34764 2574 34828
rect 1886 33767 1950 33831
rect 2014 33767 2078 33831
rect 1886 33685 1950 33749
rect 2014 33685 2078 33749
rect 1886 33602 1950 33666
rect 2014 33602 2078 33666
rect 1886 33519 1950 33583
rect 2014 33519 2078 33583
rect 1886 33436 1950 33500
rect 2014 33436 2078 33500
rect 1886 33353 1950 33417
rect 2014 33353 2078 33417
rect 1886 33270 1950 33334
rect 2014 33270 2078 33334
rect 963 28284 1027 28348
rect 1057 28284 1121 28348
rect 1151 28284 1215 28348
rect 1245 28284 1309 28348
rect 1339 28284 1403 28348
rect 1433 28284 1497 28348
rect 963 28204 1027 28268
rect 1057 28204 1121 28268
rect 1151 28204 1215 28268
rect 1245 28204 1309 28268
rect 1339 28204 1403 28268
rect 1433 28204 1497 28268
rect 963 28124 1027 28188
rect 1057 28124 1121 28188
rect 1151 28124 1215 28188
rect 1245 28124 1309 28188
rect 1339 28124 1403 28188
rect 1433 28124 1497 28188
rect 963 28044 1027 28108
rect 1057 28044 1121 28108
rect 1151 28044 1215 28108
rect 1245 28044 1309 28108
rect 1339 28044 1403 28108
rect 1433 28044 1497 28108
rect 963 27964 1027 28028
rect 1057 27964 1121 28028
rect 1151 27964 1215 28028
rect 1245 27964 1309 28028
rect 1339 27964 1403 28028
rect 1433 27964 1497 28028
rect 963 27884 1027 27948
rect 1057 27884 1121 27948
rect 1151 27884 1215 27948
rect 1245 27884 1309 27948
rect 1339 27884 1403 27948
rect 1433 27884 1497 27948
rect 963 27803 1027 27867
rect 1057 27803 1121 27867
rect 1151 27803 1215 27867
rect 1245 27803 1309 27867
rect 1339 27803 1403 27867
rect 1433 27803 1497 27867
rect 963 27722 1027 27786
rect 1057 27722 1121 27786
rect 1151 27722 1215 27786
rect 1245 27722 1309 27786
rect 1339 27722 1403 27786
rect 1433 27722 1497 27786
rect 963 27641 1027 27705
rect 1057 27641 1121 27705
rect 1151 27641 1215 27705
rect 1245 27641 1309 27705
rect 1339 27641 1403 27705
rect 1433 27641 1497 27705
rect 963 27560 1027 27624
rect 1057 27560 1121 27624
rect 1151 27560 1215 27624
rect 1245 27560 1309 27624
rect 1339 27560 1403 27624
rect 1433 27560 1497 27624
rect 963 27479 1027 27543
rect 1057 27479 1121 27543
rect 1151 27479 1215 27543
rect 1245 27479 1309 27543
rect 1339 27479 1403 27543
rect 1433 27479 1497 27543
rect 963 27398 1027 27462
rect 1057 27398 1121 27462
rect 1151 27398 1215 27462
rect 1245 27398 1309 27462
rect 1339 27398 1403 27462
rect 1433 27398 1497 27462
rect 963 27317 1027 27381
rect 1057 27317 1121 27381
rect 1151 27317 1215 27381
rect 1245 27317 1309 27381
rect 1339 27317 1403 27381
rect 1433 27317 1497 27381
rect 963 27236 1027 27300
rect 1057 27236 1121 27300
rect 1151 27236 1215 27300
rect 1245 27236 1309 27300
rect 1339 27236 1403 27300
rect 1433 27236 1497 27300
rect 963 27155 1027 27219
rect 1057 27155 1121 27219
rect 1151 27155 1215 27219
rect 1245 27155 1309 27219
rect 1339 27155 1403 27219
rect 1433 27155 1497 27219
rect 963 27074 1027 27138
rect 1057 27074 1121 27138
rect 1151 27074 1215 27138
rect 1245 27074 1309 27138
rect 1339 27074 1403 27138
rect 1433 27074 1497 27138
rect 963 26993 1027 27057
rect 1057 26993 1121 27057
rect 1151 26993 1215 27057
rect 1245 26993 1309 27057
rect 1339 26993 1403 27057
rect 1433 26993 1497 27057
rect 963 26912 1027 26976
rect 1057 26912 1121 26976
rect 1151 26912 1215 26976
rect 1245 26912 1309 26976
rect 1339 26912 1403 26976
rect 1433 26912 1497 26976
rect 963 26831 1027 26895
rect 1057 26831 1121 26895
rect 1151 26831 1215 26895
rect 1245 26831 1309 26895
rect 1339 26831 1403 26895
rect 1433 26831 1497 26895
rect 3374 39528 3438 39592
rect 3502 39528 3566 39592
rect 3374 39448 3438 39512
rect 3502 39448 3566 39512
rect 3374 39368 3438 39432
rect 3502 39368 3566 39432
rect 3374 39288 3438 39352
rect 3502 39288 3566 39352
rect 3374 39208 3438 39272
rect 3502 39208 3566 39272
rect 3374 39128 3438 39192
rect 3502 39128 3566 39192
rect 3374 39048 3438 39112
rect 3502 39048 3566 39112
rect 3374 38968 3438 39032
rect 3502 38968 3566 39032
rect 3374 38888 3438 38952
rect 3502 38888 3566 38952
rect 3374 38808 3438 38872
rect 3502 38808 3566 38872
rect 3374 38728 3438 38792
rect 3502 38728 3566 38792
rect 3374 38648 3438 38712
rect 3502 38648 3566 38712
rect 3374 38568 3438 38632
rect 3502 38568 3566 38632
rect 3374 38488 3438 38552
rect 3502 38488 3566 38552
rect 3374 38408 3438 38472
rect 3502 38408 3566 38472
rect 3374 38328 3438 38392
rect 3502 38328 3566 38392
rect 3374 38247 3438 38311
rect 3502 38247 3566 38311
rect 3374 38166 3438 38230
rect 3502 38166 3566 38230
rect 3374 38085 3438 38149
rect 3502 38085 3566 38149
rect 3374 38004 3438 38068
rect 3502 38004 3566 38068
rect 3374 37923 3438 37987
rect 3502 37923 3566 37987
rect 3374 37842 3438 37906
rect 3502 37842 3566 37906
rect 3374 37761 3438 37825
rect 3502 37761 3566 37825
rect 3374 37680 3438 37744
rect 3502 37680 3566 37744
rect 3374 37599 3438 37663
rect 3502 37599 3566 37663
rect 3374 37518 3438 37582
rect 3502 37518 3566 37582
rect 3374 37437 3438 37501
rect 3502 37437 3566 37501
rect 3374 37356 3438 37420
rect 3502 37356 3566 37420
rect 3374 37275 3438 37339
rect 3502 37275 3566 37339
rect 3374 37194 3438 37258
rect 3502 37194 3566 37258
rect 3374 37113 3438 37177
rect 3502 37113 3566 37177
rect 3374 37032 3438 37096
rect 3502 37032 3566 37096
rect 3374 36951 3438 37015
rect 3502 36951 3566 37015
rect 3374 36870 3438 36934
rect 3502 36870 3566 36934
rect 3374 36789 3438 36853
rect 3502 36789 3566 36853
rect 3374 36708 3438 36772
rect 3502 36708 3566 36772
rect 3374 36627 3438 36691
rect 3502 36627 3566 36691
rect 3374 36546 3438 36610
rect 3502 36546 3566 36610
rect 3374 36465 3438 36529
rect 3502 36465 3566 36529
rect 3374 36384 3438 36448
rect 3502 36384 3566 36448
rect 3374 36303 3438 36367
rect 3502 36303 3566 36367
rect 3374 36222 3438 36286
rect 3502 36222 3566 36286
rect 3374 36141 3438 36205
rect 3502 36141 3566 36205
rect 3374 36060 3438 36124
rect 3502 36060 3566 36124
rect 3374 35979 3438 36043
rect 3502 35979 3566 36043
rect 3374 35898 3438 35962
rect 3502 35898 3566 35962
rect 3374 35817 3438 35881
rect 3502 35817 3566 35881
rect 3374 35736 3438 35800
rect 3502 35736 3566 35800
rect 3374 35655 3438 35719
rect 3502 35655 3566 35719
rect 3374 35574 3438 35638
rect 3502 35574 3566 35638
rect 3374 35493 3438 35557
rect 3502 35493 3566 35557
rect 3374 35412 3438 35476
rect 3502 35412 3566 35476
rect 3374 35331 3438 35395
rect 3502 35331 3566 35395
rect 3374 35250 3438 35314
rect 3502 35250 3566 35314
rect 3374 35169 3438 35233
rect 3502 35169 3566 35233
rect 3374 35088 3438 35152
rect 3502 35088 3566 35152
rect 3374 35007 3438 35071
rect 3502 35007 3566 35071
rect 3374 34926 3438 34990
rect 3502 34926 3566 34990
rect 3374 34845 3438 34909
rect 3502 34845 3566 34909
rect 3374 34764 3438 34828
rect 3502 34764 3566 34828
rect 2878 34155 2942 34219
rect 3006 34155 3070 34219
rect 2878 34061 2942 34125
rect 3006 34061 3070 34125
rect 2878 33966 2942 34030
rect 3006 33966 3070 34030
rect 2878 33871 2942 33935
rect 3006 33871 3070 33935
rect 2878 33776 2942 33840
rect 3006 33776 3070 33840
rect 2878 33681 2942 33745
rect 3006 33681 3070 33745
rect 4366 39528 4430 39592
rect 4494 39528 4558 39592
rect 4366 39448 4430 39512
rect 4494 39448 4558 39512
rect 4366 39368 4430 39432
rect 4494 39368 4558 39432
rect 4366 39288 4430 39352
rect 4494 39288 4558 39352
rect 4366 39208 4430 39272
rect 4494 39208 4558 39272
rect 4366 39128 4430 39192
rect 4494 39128 4558 39192
rect 4366 39048 4430 39112
rect 4494 39048 4558 39112
rect 4366 38968 4430 39032
rect 4494 38968 4558 39032
rect 4366 38888 4430 38952
rect 4494 38888 4558 38952
rect 4366 38808 4430 38872
rect 4494 38808 4558 38872
rect 4366 38728 4430 38792
rect 4494 38728 4558 38792
rect 4366 38648 4430 38712
rect 4494 38648 4558 38712
rect 4366 38568 4430 38632
rect 4494 38568 4558 38632
rect 4366 38488 4430 38552
rect 4494 38488 4558 38552
rect 4366 38408 4430 38472
rect 4494 38408 4558 38472
rect 4366 38328 4430 38392
rect 4494 38328 4558 38392
rect 4366 38247 4430 38311
rect 4494 38247 4558 38311
rect 4366 38166 4430 38230
rect 4494 38166 4558 38230
rect 4366 38085 4430 38149
rect 4494 38085 4558 38149
rect 4366 38004 4430 38068
rect 4494 38004 4558 38068
rect 4366 37923 4430 37987
rect 4494 37923 4558 37987
rect 4366 37842 4430 37906
rect 4494 37842 4558 37906
rect 4366 37761 4430 37825
rect 4494 37761 4558 37825
rect 4366 37680 4430 37744
rect 4494 37680 4558 37744
rect 4366 37599 4430 37663
rect 4494 37599 4558 37663
rect 4366 37518 4430 37582
rect 4494 37518 4558 37582
rect 4366 37437 4430 37501
rect 4494 37437 4558 37501
rect 4366 37356 4430 37420
rect 4494 37356 4558 37420
rect 4366 37275 4430 37339
rect 4494 37275 4558 37339
rect 4366 37194 4430 37258
rect 4494 37194 4558 37258
rect 4366 37113 4430 37177
rect 4494 37113 4558 37177
rect 4366 37032 4430 37096
rect 4494 37032 4558 37096
rect 4366 36951 4430 37015
rect 4494 36951 4558 37015
rect 4366 36870 4430 36934
rect 4494 36870 4558 36934
rect 4366 36789 4430 36853
rect 4494 36789 4558 36853
rect 4366 36708 4430 36772
rect 4494 36708 4558 36772
rect 4366 36627 4430 36691
rect 4494 36627 4558 36691
rect 4366 36546 4430 36610
rect 4494 36546 4558 36610
rect 4366 36465 4430 36529
rect 4494 36465 4558 36529
rect 4366 36384 4430 36448
rect 4494 36384 4558 36448
rect 4366 36303 4430 36367
rect 4494 36303 4558 36367
rect 4366 36222 4430 36286
rect 4494 36222 4558 36286
rect 4366 36141 4430 36205
rect 4494 36141 4558 36205
rect 4366 36060 4430 36124
rect 4494 36060 4558 36124
rect 4366 35979 4430 36043
rect 4494 35979 4558 36043
rect 4366 35898 4430 35962
rect 4494 35898 4558 35962
rect 4366 35817 4430 35881
rect 4494 35817 4558 35881
rect 4366 35736 4430 35800
rect 4494 35736 4558 35800
rect 4366 35655 4430 35719
rect 4494 35655 4558 35719
rect 4366 35574 4430 35638
rect 4494 35574 4558 35638
rect 4366 35493 4430 35557
rect 4494 35493 4558 35557
rect 4366 35412 4430 35476
rect 4494 35412 4558 35476
rect 4366 35331 4430 35395
rect 4494 35331 4558 35395
rect 4366 35250 4430 35314
rect 4494 35250 4558 35314
rect 4366 35169 4430 35233
rect 4494 35169 4558 35233
rect 4366 35088 4430 35152
rect 4494 35088 4558 35152
rect 4366 35007 4430 35071
rect 4494 35007 4558 35071
rect 4366 34926 4430 34990
rect 4494 34926 4558 34990
rect 4366 34845 4430 34909
rect 4494 34845 4558 34909
rect 4366 34764 4430 34828
rect 4494 34764 4558 34828
rect 3870 34155 3934 34219
rect 3998 34155 4062 34219
rect 3870 34061 3934 34125
rect 3998 34061 4062 34125
rect 3870 33966 3934 34030
rect 3998 33966 4062 34030
rect 3870 33871 3934 33935
rect 3998 33871 4062 33935
rect 3870 33776 3934 33840
rect 3998 33776 4062 33840
rect 3870 33681 3934 33745
rect 3998 33681 4062 33745
rect 963 26750 1027 26814
rect 1057 26750 1121 26814
rect 1151 26750 1215 26814
rect 1245 26750 1309 26814
rect 1339 26750 1403 26814
rect 1433 26750 1497 26814
rect 963 26669 1027 26733
rect 1057 26669 1121 26733
rect 1151 26669 1215 26733
rect 1245 26669 1309 26733
rect 1339 26669 1403 26733
rect 1433 26669 1497 26733
rect 963 26588 1027 26652
rect 1057 26588 1121 26652
rect 1151 26588 1215 26652
rect 1245 26588 1309 26652
rect 1339 26588 1403 26652
rect 1433 26588 1497 26652
rect 963 26507 1027 26571
rect 1057 26507 1121 26571
rect 1151 26507 1215 26571
rect 1245 26507 1309 26571
rect 1339 26507 1403 26571
rect 1433 26507 1497 26571
rect 963 26426 1027 26490
rect 1057 26426 1121 26490
rect 1151 26426 1215 26490
rect 1245 26426 1309 26490
rect 1339 26426 1403 26490
rect 1433 26426 1497 26490
rect 963 26345 1027 26409
rect 1057 26345 1121 26409
rect 1151 26345 1215 26409
rect 1245 26345 1309 26409
rect 1339 26345 1403 26409
rect 1433 26345 1497 26409
rect 963 26264 1027 26328
rect 1057 26264 1121 26328
rect 1151 26264 1215 26328
rect 1245 26264 1309 26328
rect 1339 26264 1403 26328
rect 1433 26264 1497 26328
rect 963 26183 1027 26247
rect 1057 26183 1121 26247
rect 1151 26183 1215 26247
rect 1245 26183 1309 26247
rect 1339 26183 1403 26247
rect 1433 26183 1497 26247
rect 963 26102 1027 26166
rect 1057 26102 1121 26166
rect 1151 26102 1215 26166
rect 1245 26102 1309 26166
rect 1339 26102 1403 26166
rect 1433 26102 1497 26166
rect 963 26021 1027 26085
rect 1057 26021 1121 26085
rect 1151 26021 1215 26085
rect 1245 26021 1309 26085
rect 1339 26021 1403 26085
rect 1433 26021 1497 26085
rect 963 25940 1027 26004
rect 1057 25940 1121 26004
rect 1151 25940 1215 26004
rect 1245 25940 1309 26004
rect 1339 25940 1403 26004
rect 1433 25940 1497 26004
rect 963 25859 1027 25923
rect 1057 25859 1121 25923
rect 1151 25859 1215 25923
rect 1245 25859 1309 25923
rect 1339 25859 1403 25923
rect 1433 25859 1497 25923
rect 963 25778 1027 25842
rect 1057 25778 1121 25842
rect 1151 25778 1215 25842
rect 1245 25778 1309 25842
rect 1339 25778 1403 25842
rect 1433 25778 1497 25842
rect 963 25697 1027 25761
rect 1057 25697 1121 25761
rect 1151 25697 1215 25761
rect 1245 25697 1309 25761
rect 1339 25697 1403 25761
rect 1433 25697 1497 25761
rect 963 25616 1027 25680
rect 1057 25616 1121 25680
rect 1151 25616 1215 25680
rect 1245 25616 1309 25680
rect 1339 25616 1403 25680
rect 1433 25616 1497 25680
rect 963 25535 1027 25599
rect 1057 25535 1121 25599
rect 1151 25535 1215 25599
rect 1245 25535 1309 25599
rect 1339 25535 1403 25599
rect 1433 25535 1497 25599
rect 963 25454 1027 25518
rect 1057 25454 1121 25518
rect 1151 25454 1215 25518
rect 1245 25454 1309 25518
rect 1339 25454 1403 25518
rect 1433 25454 1497 25518
rect 963 25373 1027 25437
rect 1057 25373 1121 25437
rect 1151 25373 1215 25437
rect 1245 25373 1309 25437
rect 1339 25373 1403 25437
rect 1433 25373 1497 25437
rect 963 25292 1027 25356
rect 1057 25292 1121 25356
rect 1151 25292 1215 25356
rect 1245 25292 1309 25356
rect 1339 25292 1403 25356
rect 1433 25292 1497 25356
rect 963 25211 1027 25275
rect 1057 25211 1121 25275
rect 1151 25211 1215 25275
rect 1245 25211 1309 25275
rect 1339 25211 1403 25275
rect 1433 25211 1497 25275
rect 963 25130 1027 25194
rect 1057 25130 1121 25194
rect 1151 25130 1215 25194
rect 1245 25130 1309 25194
rect 1339 25130 1403 25194
rect 1433 25130 1497 25194
rect 963 25049 1027 25113
rect 1057 25049 1121 25113
rect 1151 25049 1215 25113
rect 1245 25049 1309 25113
rect 1339 25049 1403 25113
rect 1433 25049 1497 25113
rect 963 24968 1027 25032
rect 1057 24968 1121 25032
rect 1151 24968 1215 25032
rect 1245 24968 1309 25032
rect 1339 24968 1403 25032
rect 1433 24968 1497 25032
rect 963 24887 1027 24951
rect 1057 24887 1121 24951
rect 1151 24887 1215 24951
rect 1245 24887 1309 24951
rect 1339 24887 1403 24951
rect 1433 24887 1497 24951
rect 1009 23630 1065 23685
rect 1065 23630 1073 23685
rect 1009 23621 1073 23630
rect 1103 23630 1111 23685
rect 1111 23630 1167 23685
rect 1103 23621 1167 23630
rect 1009 23550 1065 23604
rect 1065 23550 1073 23604
rect 1009 23540 1073 23550
rect 1103 23550 1111 23604
rect 1111 23550 1167 23604
rect 1103 23540 1167 23550
rect 1009 23470 1065 23522
rect 1065 23470 1073 23522
rect 1009 23458 1073 23470
rect 1103 23470 1111 23522
rect 1111 23470 1167 23522
rect 1103 23458 1167 23470
rect 1009 23390 1065 23440
rect 1065 23390 1073 23440
rect 1009 23376 1073 23390
rect 1103 23390 1111 23440
rect 1111 23390 1167 23440
rect 1103 23376 1167 23390
rect 1009 23310 1065 23358
rect 1065 23310 1073 23358
rect 1009 23294 1073 23310
rect 1103 23310 1111 23358
rect 1111 23310 1167 23358
rect 1103 23294 1167 23310
rect 1009 23230 1065 23276
rect 1065 23230 1073 23276
rect 1009 23212 1073 23230
rect 1103 23230 1111 23276
rect 1111 23230 1167 23276
rect 1103 23212 1167 23230
rect 1009 23150 1065 23194
rect 1065 23150 1073 23194
rect 1009 23130 1073 23150
rect 1103 23150 1111 23194
rect 1111 23150 1167 23194
rect 1103 23130 1167 23150
rect 1009 23070 1065 23112
rect 1065 23070 1073 23112
rect 1009 23048 1073 23070
rect 1103 23070 1111 23112
rect 1111 23070 1167 23112
rect 1103 23048 1167 23070
rect 1009 22990 1065 23030
rect 1065 22990 1073 23030
rect 1009 22966 1073 22990
rect 1103 22990 1111 23030
rect 1111 22990 1167 23030
rect 1103 22966 1167 22990
rect 1009 22910 1065 22948
rect 1065 22910 1073 22948
rect 1009 22886 1073 22910
rect 1009 22884 1065 22886
rect 1065 22884 1073 22886
rect 1103 22910 1111 22948
rect 1111 22910 1167 22948
rect 1103 22886 1167 22910
rect 1103 22884 1111 22886
rect 1111 22884 1167 22886
rect 1009 22830 1065 22866
rect 1065 22830 1073 22866
rect 1009 22806 1073 22830
rect 1009 22802 1065 22806
rect 1065 22802 1073 22806
rect 1103 22830 1111 22866
rect 1111 22830 1167 22866
rect 1103 22806 1167 22830
rect 1103 22802 1111 22806
rect 1111 22802 1167 22806
rect 1009 22750 1065 22784
rect 1065 22750 1073 22784
rect 1009 22726 1073 22750
rect 1009 22720 1065 22726
rect 1065 22720 1073 22726
rect 1103 22750 1111 22784
rect 1111 22750 1167 22784
rect 1103 22726 1167 22750
rect 1103 22720 1111 22726
rect 1111 22720 1167 22726
rect 1009 22670 1065 22702
rect 1065 22670 1073 22702
rect 1009 22646 1073 22670
rect 1009 22638 1065 22646
rect 1065 22638 1073 22646
rect 1103 22670 1111 22702
rect 1111 22670 1167 22702
rect 1103 22646 1167 22670
rect 1103 22638 1111 22646
rect 1111 22638 1167 22646
rect 1009 22590 1065 22620
rect 1065 22590 1073 22620
rect 1009 22566 1073 22590
rect 1009 22556 1065 22566
rect 1065 22556 1073 22566
rect 1103 22590 1111 22620
rect 1111 22590 1167 22620
rect 1103 22566 1167 22590
rect 1103 22556 1111 22566
rect 1111 22556 1167 22566
rect 1009 22510 1065 22538
rect 1065 22510 1073 22538
rect 1009 22486 1073 22510
rect 1009 22474 1065 22486
rect 1065 22474 1073 22486
rect 1103 22510 1111 22538
rect 1111 22510 1167 22538
rect 1103 22486 1167 22510
rect 1103 22474 1111 22486
rect 1111 22474 1167 22486
rect 1009 22430 1065 22456
rect 1065 22430 1073 22456
rect 1009 22406 1073 22430
rect 1009 22392 1065 22406
rect 1065 22392 1073 22406
rect 1103 22430 1111 22456
rect 1111 22430 1167 22456
rect 1103 22406 1167 22430
rect 1103 22392 1111 22406
rect 1111 22392 1167 22406
rect 1009 22350 1065 22374
rect 1065 22350 1073 22374
rect 1009 22326 1073 22350
rect 1009 22310 1065 22326
rect 1065 22310 1073 22326
rect 1103 22350 1111 22374
rect 1111 22350 1167 22374
rect 1103 22326 1167 22350
rect 1103 22310 1111 22326
rect 1111 22310 1167 22326
rect 1009 22270 1065 22292
rect 1065 22270 1073 22292
rect 1009 22245 1073 22270
rect 1009 22228 1065 22245
rect 1065 22228 1073 22245
rect 1103 22270 1111 22292
rect 1111 22270 1167 22292
rect 1103 22245 1167 22270
rect 1103 22228 1111 22245
rect 1111 22228 1167 22245
rect 1009 22189 1065 22210
rect 1065 22189 1073 22210
rect 1009 22164 1073 22189
rect 1009 22146 1065 22164
rect 1065 22146 1073 22164
rect 1103 22189 1111 22210
rect 1111 22189 1167 22210
rect 1103 22164 1167 22189
rect 1103 22146 1111 22164
rect 1111 22146 1167 22164
rect 1009 22108 1065 22128
rect 1065 22108 1073 22128
rect 1009 22083 1073 22108
rect 1009 22064 1065 22083
rect 1065 22064 1073 22083
rect 1103 22108 1111 22128
rect 1111 22108 1167 22128
rect 1103 22083 1167 22108
rect 1103 22064 1111 22083
rect 1111 22064 1167 22083
rect 1009 22027 1065 22046
rect 1065 22027 1073 22046
rect 1009 22002 1073 22027
rect 1009 21982 1065 22002
rect 1065 21982 1073 22002
rect 1103 22027 1111 22046
rect 1111 22027 1167 22046
rect 1103 22002 1167 22027
rect 1103 21982 1111 22002
rect 1111 21982 1167 22002
rect 1009 21946 1065 21964
rect 1065 21946 1073 21964
rect 1009 21921 1073 21946
rect 1009 21900 1065 21921
rect 1065 21900 1073 21921
rect 1103 21946 1111 21964
rect 1111 21946 1167 21964
rect 1103 21921 1167 21946
rect 1103 21900 1111 21921
rect 1111 21900 1167 21921
rect 1009 21865 1065 21882
rect 1065 21865 1073 21882
rect 1009 21840 1073 21865
rect 1009 21818 1065 21840
rect 1065 21818 1073 21840
rect 1103 21865 1111 21882
rect 1111 21865 1167 21882
rect 1103 21840 1167 21865
rect 1103 21818 1111 21840
rect 1111 21818 1167 21840
rect 1986 19926 2050 19990
rect 2102 19926 2166 19990
rect 456 15484 1160 18588
rect 456 15403 520 15467
rect 536 15403 600 15467
rect 616 15403 680 15467
rect 696 15403 760 15467
rect 776 15403 840 15467
rect 856 15403 920 15467
rect 936 15403 1000 15467
rect 1016 15403 1080 15467
rect 1096 15403 1160 15467
rect 456 15322 520 15386
rect 536 15322 600 15386
rect 616 15322 680 15386
rect 696 15322 760 15386
rect 776 15322 840 15386
rect 856 15322 920 15386
rect 936 15322 1000 15386
rect 1016 15322 1080 15386
rect 1096 15322 1160 15386
rect 456 15241 520 15305
rect 536 15241 600 15305
rect 616 15241 680 15305
rect 696 15241 760 15305
rect 776 15241 840 15305
rect 856 15241 920 15305
rect 936 15241 1000 15305
rect 1016 15241 1080 15305
rect 1096 15241 1160 15305
rect 456 15160 520 15224
rect 536 15160 600 15224
rect 616 15160 680 15224
rect 696 15160 760 15224
rect 776 15160 840 15224
rect 856 15160 920 15224
rect 936 15160 1000 15224
rect 1016 15160 1080 15224
rect 1096 15160 1160 15224
rect 456 15079 520 15143
rect 536 15079 600 15143
rect 616 15079 680 15143
rect 696 15079 760 15143
rect 776 15079 840 15143
rect 856 15079 920 15143
rect 936 15079 1000 15143
rect 1016 15079 1080 15143
rect 1096 15079 1160 15143
rect 456 14998 520 15062
rect 536 14998 600 15062
rect 616 14998 680 15062
rect 696 14998 760 15062
rect 776 14998 840 15062
rect 856 14998 920 15062
rect 936 14998 1000 15062
rect 1016 14998 1080 15062
rect 1096 14998 1160 15062
rect 456 14917 520 14981
rect 536 14917 600 14981
rect 616 14917 680 14981
rect 696 14917 760 14981
rect 776 14917 840 14981
rect 856 14917 920 14981
rect 936 14917 1000 14981
rect 1016 14917 1080 14981
rect 1096 14917 1160 14981
rect 456 14836 520 14900
rect 536 14836 600 14900
rect 616 14836 680 14900
rect 696 14836 760 14900
rect 776 14836 840 14900
rect 856 14836 920 14900
rect 936 14836 1000 14900
rect 1016 14836 1080 14900
rect 1096 14836 1160 14900
rect 456 14755 520 14819
rect 536 14755 600 14819
rect 616 14755 680 14819
rect 696 14755 760 14819
rect 776 14755 840 14819
rect 856 14755 920 14819
rect 936 14755 1000 14819
rect 1016 14755 1080 14819
rect 1096 14755 1160 14819
rect 456 14674 520 14738
rect 536 14674 600 14738
rect 616 14674 680 14738
rect 696 14674 760 14738
rect 776 14674 840 14738
rect 856 14674 920 14738
rect 936 14674 1000 14738
rect 1016 14674 1080 14738
rect 1096 14674 1160 14738
rect 456 14593 520 14657
rect 536 14593 600 14657
rect 616 14593 680 14657
rect 696 14593 760 14657
rect 776 14593 840 14657
rect 856 14593 920 14657
rect 936 14593 1000 14657
rect 1016 14593 1080 14657
rect 1096 14593 1160 14657
rect 456 14512 520 14576
rect 536 14512 600 14576
rect 616 14512 680 14576
rect 696 14512 760 14576
rect 776 14512 840 14576
rect 856 14512 920 14576
rect 936 14512 1000 14576
rect 1016 14512 1080 14576
rect 1096 14512 1160 14576
rect 456 14431 520 14495
rect 536 14431 600 14495
rect 616 14431 680 14495
rect 696 14431 760 14495
rect 776 14431 840 14495
rect 856 14431 920 14495
rect 936 14431 1000 14495
rect 1016 14431 1080 14495
rect 1096 14431 1160 14495
rect 456 14350 520 14414
rect 536 14350 600 14414
rect 616 14350 680 14414
rect 696 14350 760 14414
rect 776 14350 840 14414
rect 856 14350 920 14414
rect 936 14350 1000 14414
rect 1016 14350 1080 14414
rect 1096 14350 1160 14414
rect 456 14269 520 14333
rect 536 14269 600 14333
rect 616 14269 680 14333
rect 696 14269 760 14333
rect 776 14269 840 14333
rect 856 14269 920 14333
rect 936 14269 1000 14333
rect 1016 14269 1080 14333
rect 1096 14269 1160 14333
rect 456 14188 520 14252
rect 536 14188 600 14252
rect 616 14188 680 14252
rect 696 14188 760 14252
rect 776 14188 840 14252
rect 856 14188 920 14252
rect 936 14188 1000 14252
rect 1016 14188 1080 14252
rect 1096 14188 1160 14252
rect 456 14107 520 14171
rect 536 14107 600 14171
rect 616 14107 680 14171
rect 696 14107 760 14171
rect 776 14107 840 14171
rect 856 14107 920 14171
rect 936 14107 1000 14171
rect 1016 14107 1080 14171
rect 1096 14107 1160 14171
rect 456 14026 520 14090
rect 536 14026 600 14090
rect 616 14026 680 14090
rect 696 14026 760 14090
rect 776 14026 840 14090
rect 856 14026 920 14090
rect 936 14026 1000 14090
rect 1016 14026 1080 14090
rect 1096 14026 1160 14090
rect 456 13945 520 14009
rect 536 13945 600 14009
rect 616 13945 680 14009
rect 696 13945 760 14009
rect 776 13945 840 14009
rect 856 13945 920 14009
rect 936 13945 1000 14009
rect 1016 13945 1080 14009
rect 1096 13945 1160 14009
rect 456 13864 520 13928
rect 536 13864 600 13928
rect 616 13864 680 13928
rect 696 13864 760 13928
rect 776 13864 840 13928
rect 856 13864 920 13928
rect 936 13864 1000 13928
rect 1016 13864 1080 13928
rect 1096 13864 1160 13928
rect 456 13783 520 13847
rect 536 13783 600 13847
rect 616 13783 680 13847
rect 696 13783 760 13847
rect 776 13783 840 13847
rect 856 13783 920 13847
rect 936 13783 1000 13847
rect 1016 13783 1080 13847
rect 1096 13783 1160 13847
rect 456 13702 520 13766
rect 536 13702 600 13766
rect 616 13702 680 13766
rect 696 13702 760 13766
rect 776 13702 840 13766
rect 856 13702 920 13766
rect 936 13702 1000 13766
rect 1016 13702 1080 13766
rect 1096 13702 1160 13766
rect 456 13621 520 13685
rect 536 13621 600 13685
rect 616 13621 680 13685
rect 696 13621 760 13685
rect 776 13621 840 13685
rect 856 13621 920 13685
rect 936 13621 1000 13685
rect 1016 13621 1080 13685
rect 1096 13621 1160 13685
rect 1287 18522 1351 18586
rect 1375 18522 1439 18586
rect 1463 18522 1527 18586
rect 1551 18522 1615 18586
rect 1639 18522 1703 18586
rect 1727 18522 1791 18586
rect 1815 18522 1879 18586
rect 1287 18442 1351 18506
rect 1375 18442 1439 18506
rect 1463 18442 1527 18506
rect 1551 18442 1615 18506
rect 1639 18442 1703 18506
rect 1727 18442 1791 18506
rect 1815 18442 1879 18506
rect 1287 18362 1351 18426
rect 1375 18362 1439 18426
rect 1463 18362 1527 18426
rect 1551 18362 1615 18426
rect 1639 18362 1703 18426
rect 1727 18362 1791 18426
rect 1815 18362 1879 18426
rect 1287 18282 1351 18346
rect 1375 18282 1439 18346
rect 1463 18282 1527 18346
rect 1551 18282 1615 18346
rect 1639 18282 1703 18346
rect 1727 18282 1791 18346
rect 1815 18282 1879 18346
rect 1287 18202 1351 18266
rect 1375 18202 1439 18266
rect 1463 18202 1527 18266
rect 1551 18202 1615 18266
rect 1639 18202 1703 18266
rect 1727 18202 1791 18266
rect 1815 18202 1879 18266
rect 1287 18122 1351 18186
rect 1375 18122 1439 18186
rect 1463 18122 1527 18186
rect 1551 18122 1615 18186
rect 1639 18122 1703 18186
rect 1727 18122 1791 18186
rect 1815 18122 1879 18186
rect 1287 18042 1351 18106
rect 1375 18042 1439 18106
rect 1463 18042 1527 18106
rect 1551 18042 1615 18106
rect 1639 18042 1703 18106
rect 1727 18042 1791 18106
rect 1815 18042 1879 18106
rect 1287 17962 1351 18026
rect 1375 17962 1439 18026
rect 1463 17962 1527 18026
rect 1551 17962 1615 18026
rect 1639 17962 1703 18026
rect 1727 17962 1791 18026
rect 1815 17962 1879 18026
rect 1287 17882 1351 17946
rect 1375 17882 1439 17946
rect 1463 17882 1527 17946
rect 1551 17882 1615 17946
rect 1639 17882 1703 17946
rect 1727 17882 1791 17946
rect 1815 17882 1879 17946
rect 1287 17802 1351 17866
rect 1375 17802 1439 17866
rect 1463 17802 1527 17866
rect 1551 17802 1615 17866
rect 1639 17802 1703 17866
rect 1727 17802 1791 17866
rect 1815 17802 1879 17866
rect 1287 17722 1351 17786
rect 1375 17722 1439 17786
rect 1463 17722 1527 17786
rect 1551 17722 1615 17786
rect 1639 17722 1703 17786
rect 1727 17722 1791 17786
rect 1815 17722 1879 17786
rect 1287 17642 1351 17706
rect 1375 17642 1439 17706
rect 1463 17642 1527 17706
rect 1551 17642 1615 17706
rect 1639 17642 1703 17706
rect 1727 17642 1791 17706
rect 1815 17642 1879 17706
rect 1287 17562 1351 17626
rect 1375 17562 1439 17626
rect 1463 17562 1527 17626
rect 1551 17562 1615 17626
rect 1639 17562 1703 17626
rect 1727 17562 1791 17626
rect 1815 17562 1879 17626
rect 1287 17482 1351 17546
rect 1375 17482 1439 17546
rect 1463 17482 1527 17546
rect 1551 17482 1615 17546
rect 1639 17482 1703 17546
rect 1727 17482 1791 17546
rect 1815 17482 1879 17546
rect 1287 17402 1351 17466
rect 1375 17402 1439 17466
rect 1463 17402 1527 17466
rect 1551 17402 1615 17466
rect 1639 17402 1703 17466
rect 1727 17402 1791 17466
rect 1815 17402 1879 17466
rect 1287 17322 1351 17386
rect 1375 17322 1439 17386
rect 1463 17322 1527 17386
rect 1551 17322 1615 17386
rect 1639 17322 1703 17386
rect 1727 17322 1791 17386
rect 1815 17322 1879 17386
rect 1287 17242 1351 17306
rect 1375 17242 1439 17306
rect 1463 17242 1527 17306
rect 1551 17242 1615 17306
rect 1639 17242 1703 17306
rect 1727 17242 1791 17306
rect 1815 17242 1879 17306
rect 1287 17162 1351 17226
rect 1375 17162 1439 17226
rect 1463 17162 1527 17226
rect 1551 17162 1615 17226
rect 1639 17162 1703 17226
rect 1727 17162 1791 17226
rect 1815 17162 1879 17226
rect 1287 17082 1351 17146
rect 1375 17082 1439 17146
rect 1463 17082 1527 17146
rect 1551 17082 1615 17146
rect 1639 17082 1703 17146
rect 1727 17082 1791 17146
rect 1815 17082 1879 17146
rect 1287 17002 1351 17066
rect 1375 17002 1439 17066
rect 1463 17002 1527 17066
rect 1551 17002 1615 17066
rect 1639 17002 1703 17066
rect 1727 17002 1791 17066
rect 1815 17002 1879 17066
rect 1287 16922 1351 16986
rect 1375 16922 1439 16986
rect 1463 16922 1527 16986
rect 1551 16922 1615 16986
rect 1639 16922 1703 16986
rect 1727 16922 1791 16986
rect 1815 16922 1879 16986
rect 1287 16842 1351 16906
rect 1375 16842 1439 16906
rect 1463 16842 1527 16906
rect 1551 16842 1615 16906
rect 1639 16842 1703 16906
rect 1727 16842 1791 16906
rect 1815 16842 1879 16906
rect 1287 16762 1351 16826
rect 1375 16762 1439 16826
rect 1463 16762 1527 16826
rect 1551 16762 1615 16826
rect 1639 16762 1703 16826
rect 1727 16762 1791 16826
rect 1815 16762 1879 16826
rect 1287 16682 1351 16746
rect 1375 16682 1439 16746
rect 1463 16682 1527 16746
rect 1551 16682 1615 16746
rect 1639 16682 1703 16746
rect 1727 16682 1791 16746
rect 1815 16682 1879 16746
rect 1287 16602 1351 16666
rect 1375 16602 1439 16666
rect 1463 16602 1527 16666
rect 1551 16602 1615 16666
rect 1639 16602 1703 16666
rect 1727 16602 1791 16666
rect 1815 16602 1879 16666
rect 1287 16522 1351 16586
rect 1375 16522 1439 16586
rect 1463 16522 1527 16586
rect 1551 16522 1615 16586
rect 1639 16522 1703 16586
rect 1727 16522 1791 16586
rect 1815 16522 1879 16586
rect 1287 16442 1351 16506
rect 1375 16442 1439 16506
rect 1463 16442 1527 16506
rect 1551 16442 1615 16506
rect 1639 16442 1703 16506
rect 1727 16442 1791 16506
rect 1815 16442 1879 16506
rect 1287 16362 1351 16426
rect 1375 16362 1439 16426
rect 1463 16362 1527 16426
rect 1551 16362 1615 16426
rect 1639 16362 1703 16426
rect 1727 16362 1791 16426
rect 1815 16362 1879 16426
rect 1287 16282 1351 16346
rect 1375 16282 1439 16346
rect 1463 16282 1527 16346
rect 1551 16282 1615 16346
rect 1639 16282 1703 16346
rect 1727 16282 1791 16346
rect 1815 16282 1879 16346
rect 1287 16202 1351 16266
rect 1375 16202 1439 16266
rect 1463 16202 1527 16266
rect 1551 16202 1615 16266
rect 1639 16202 1703 16266
rect 1727 16202 1791 16266
rect 1815 16202 1879 16266
rect 1287 16122 1351 16186
rect 1375 16122 1439 16186
rect 1463 16122 1527 16186
rect 1551 16122 1615 16186
rect 1639 16122 1703 16186
rect 1727 16122 1791 16186
rect 1815 16122 1879 16186
rect 1287 16042 1351 16106
rect 1375 16042 1439 16106
rect 1463 16042 1527 16106
rect 1551 16042 1615 16106
rect 1639 16042 1703 16106
rect 1727 16042 1791 16106
rect 1815 16042 1879 16106
rect 1287 15962 1351 16026
rect 1375 15962 1439 16026
rect 1463 15962 1527 16026
rect 1551 15962 1615 16026
rect 1639 15962 1703 16026
rect 1727 15962 1791 16026
rect 1815 15962 1879 16026
rect 1287 15882 1351 15946
rect 1375 15882 1439 15946
rect 1463 15882 1527 15946
rect 1551 15882 1615 15946
rect 1639 15882 1703 15946
rect 1727 15882 1791 15946
rect 1815 15882 1879 15946
rect 1287 15802 1351 15866
rect 1375 15802 1439 15866
rect 1463 15802 1527 15866
rect 1551 15802 1615 15866
rect 1639 15802 1703 15866
rect 1727 15802 1791 15866
rect 1815 15802 1879 15866
rect 1287 15722 1351 15786
rect 1375 15722 1439 15786
rect 1463 15722 1527 15786
rect 1551 15722 1615 15786
rect 1639 15722 1703 15786
rect 1727 15722 1791 15786
rect 1815 15722 1879 15786
rect 1287 15642 1351 15706
rect 1375 15642 1439 15706
rect 1463 15642 1527 15706
rect 1551 15642 1615 15706
rect 1639 15642 1703 15706
rect 1727 15642 1791 15706
rect 1815 15642 1879 15706
rect 1287 15562 1351 15626
rect 1375 15562 1439 15626
rect 1463 15562 1527 15626
rect 1551 15562 1615 15626
rect 1639 15562 1703 15626
rect 1727 15562 1791 15626
rect 1815 15562 1879 15626
rect 1287 15482 1351 15546
rect 1375 15482 1439 15546
rect 1463 15482 1527 15546
rect 1551 15482 1615 15546
rect 1639 15482 1703 15546
rect 1727 15482 1791 15546
rect 1815 15482 1879 15546
rect 1287 15402 1351 15466
rect 1375 15402 1439 15466
rect 1463 15402 1527 15466
rect 1551 15402 1615 15466
rect 1639 15402 1703 15466
rect 1727 15402 1791 15466
rect 1815 15402 1879 15466
rect 1287 15322 1351 15386
rect 1375 15322 1439 15386
rect 1463 15322 1527 15386
rect 1551 15322 1615 15386
rect 1639 15322 1703 15386
rect 1727 15322 1791 15386
rect 1815 15322 1879 15386
rect 1287 15242 1351 15306
rect 1375 15242 1439 15306
rect 1463 15242 1527 15306
rect 1551 15242 1615 15306
rect 1639 15242 1703 15306
rect 1727 15242 1791 15306
rect 1815 15242 1879 15306
rect 1287 15162 1351 15226
rect 1375 15162 1439 15226
rect 1463 15162 1527 15226
rect 1551 15162 1615 15226
rect 1639 15162 1703 15226
rect 1727 15162 1791 15226
rect 1815 15162 1879 15226
rect 1287 15082 1351 15146
rect 1375 15082 1439 15146
rect 1463 15082 1527 15146
rect 1551 15082 1615 15146
rect 1639 15082 1703 15146
rect 1727 15082 1791 15146
rect 1815 15082 1879 15146
rect 1287 15002 1351 15066
rect 1375 15002 1439 15066
rect 1463 15002 1527 15066
rect 1551 15002 1615 15066
rect 1639 15002 1703 15066
rect 1727 15002 1791 15066
rect 1815 15002 1879 15066
rect 1287 14922 1351 14986
rect 1375 14922 1439 14986
rect 1463 14922 1527 14986
rect 1551 14922 1615 14986
rect 1639 14922 1703 14986
rect 1727 14922 1791 14986
rect 1815 14922 1879 14986
rect 1287 14842 1351 14906
rect 1375 14842 1439 14906
rect 1463 14842 1527 14906
rect 1551 14842 1615 14906
rect 1639 14842 1703 14906
rect 1727 14842 1791 14906
rect 1815 14842 1879 14906
rect 1287 14762 1351 14826
rect 1375 14762 1439 14826
rect 1463 14762 1527 14826
rect 1551 14762 1615 14826
rect 1639 14762 1703 14826
rect 1727 14762 1791 14826
rect 1815 14762 1879 14826
rect 1287 14682 1351 14746
rect 1375 14682 1439 14746
rect 1463 14682 1527 14746
rect 1551 14682 1615 14746
rect 1639 14682 1703 14746
rect 1727 14682 1791 14746
rect 1815 14682 1879 14746
rect 1287 14602 1351 14666
rect 1375 14602 1439 14666
rect 1463 14602 1527 14666
rect 1551 14602 1615 14666
rect 1639 14602 1703 14666
rect 1727 14602 1791 14666
rect 1815 14602 1879 14666
rect 1287 14522 1351 14586
rect 1375 14522 1439 14586
rect 1463 14522 1527 14586
rect 1551 14522 1615 14586
rect 1639 14522 1703 14586
rect 1727 14522 1791 14586
rect 1815 14522 1879 14586
rect 1287 14441 1351 14505
rect 1375 14441 1439 14505
rect 1463 14441 1527 14505
rect 1551 14441 1615 14505
rect 1639 14441 1703 14505
rect 1727 14441 1791 14505
rect 1815 14441 1879 14505
rect 1287 14360 1351 14424
rect 1375 14360 1439 14424
rect 1463 14360 1527 14424
rect 1551 14360 1615 14424
rect 1639 14360 1703 14424
rect 1727 14360 1791 14424
rect 1815 14360 1879 14424
rect 1287 14279 1351 14343
rect 1375 14279 1439 14343
rect 1463 14279 1527 14343
rect 1551 14279 1615 14343
rect 1639 14279 1703 14343
rect 1727 14279 1791 14343
rect 1815 14279 1879 14343
rect 1287 14198 1351 14262
rect 1375 14198 1439 14262
rect 1463 14198 1527 14262
rect 1551 14198 1615 14262
rect 1639 14198 1703 14262
rect 1727 14198 1791 14262
rect 1815 14198 1879 14262
rect 1287 14117 1351 14181
rect 1375 14117 1439 14181
rect 1463 14117 1527 14181
rect 1551 14117 1615 14181
rect 1639 14117 1703 14181
rect 1727 14117 1791 14181
rect 1815 14117 1879 14181
rect 1287 14036 1351 14100
rect 1375 14036 1439 14100
rect 1463 14036 1527 14100
rect 1551 14036 1615 14100
rect 1639 14036 1703 14100
rect 1727 14036 1791 14100
rect 1815 14036 1879 14100
rect 1287 13955 1351 14019
rect 1375 13955 1439 14019
rect 1463 13955 1527 14019
rect 1551 13955 1615 14019
rect 1639 13955 1703 14019
rect 1727 13955 1791 14019
rect 1815 13955 1879 14019
rect 1287 13874 1351 13938
rect 1375 13874 1439 13938
rect 1463 13874 1527 13938
rect 1551 13874 1615 13938
rect 1639 13874 1703 13938
rect 1727 13874 1791 13938
rect 1815 13874 1879 13938
rect 1287 13793 1351 13857
rect 1375 13793 1439 13857
rect 1463 13793 1527 13857
rect 1551 13793 1615 13857
rect 1639 13793 1703 13857
rect 1727 13793 1791 13857
rect 1815 13793 1879 13857
rect 1287 13712 1351 13776
rect 1375 13712 1439 13776
rect 1463 13712 1527 13776
rect 1551 13712 1615 13776
rect 1639 13712 1703 13776
rect 1727 13712 1791 13776
rect 1815 13712 1879 13776
rect 1287 13631 1351 13695
rect 1375 13631 1439 13695
rect 1463 13631 1527 13695
rect 1551 13631 1615 13695
rect 1639 13631 1703 13695
rect 1727 13631 1791 13695
rect 1815 13631 1879 13695
rect 1986 19843 2050 19907
rect 2102 19843 2166 19907
rect 1986 19759 2050 19823
rect 2102 19759 2166 19823
rect 1986 19675 2050 19739
rect 2102 19675 2166 19739
rect 1986 19591 2050 19655
rect 2102 19591 2166 19655
rect 1986 19507 2050 19571
rect 2102 19507 2166 19571
rect 1986 19423 2050 19487
rect 2102 19423 2166 19487
rect 2480 18528 2544 18592
rect 2608 18528 2672 18592
rect 2480 18448 2544 18512
rect 2608 18448 2672 18512
rect 2480 18368 2544 18432
rect 2608 18368 2672 18432
rect 2480 18288 2544 18352
rect 2608 18288 2672 18352
rect 2480 18208 2544 18272
rect 2608 18208 2672 18272
rect 2480 18128 2544 18192
rect 2608 18128 2672 18192
rect 2480 18048 2544 18112
rect 2608 18048 2672 18112
rect 2480 17968 2544 18032
rect 2608 17968 2672 18032
rect 2480 17888 2544 17952
rect 2608 17888 2672 17952
rect 2480 17808 2544 17872
rect 2608 17808 2672 17872
rect 2480 17728 2544 17792
rect 2608 17728 2672 17792
rect 2480 17648 2544 17712
rect 2608 17648 2672 17712
rect 2480 17568 2544 17632
rect 2608 17568 2672 17632
rect 2480 17488 2544 17552
rect 2608 17488 2672 17552
rect 2480 17408 2544 17472
rect 2608 17408 2672 17472
rect 2480 17328 2544 17392
rect 2608 17328 2672 17392
rect 2480 17248 2544 17312
rect 2608 17248 2672 17312
rect 2480 17168 2544 17232
rect 2608 17168 2672 17232
rect 2480 17088 2544 17152
rect 2608 17088 2672 17152
rect 2480 17008 2544 17072
rect 2608 17008 2672 17072
rect 2480 16928 2544 16992
rect 2608 16928 2672 16992
rect 2480 16848 2544 16912
rect 2608 16848 2672 16912
rect 2480 16768 2544 16832
rect 2608 16768 2672 16832
rect 2480 16688 2544 16752
rect 2608 16688 2672 16752
rect 2480 16608 2544 16672
rect 2608 16608 2672 16672
rect 2480 16528 2544 16592
rect 2608 16528 2672 16592
rect 2480 16448 2544 16512
rect 2608 16448 2672 16512
rect 2480 16368 2544 16432
rect 2608 16368 2672 16432
rect 2480 16287 2544 16351
rect 2608 16287 2672 16351
rect 2480 16206 2544 16270
rect 2608 16206 2672 16270
rect 2480 16125 2544 16189
rect 2608 16125 2672 16189
rect 2480 16044 2544 16108
rect 2608 16044 2672 16108
rect 2480 15963 2544 16027
rect 2608 15963 2672 16027
rect 2480 15882 2544 15946
rect 2608 15882 2672 15946
rect 2480 15801 2544 15865
rect 2608 15801 2672 15865
rect 2480 15720 2544 15784
rect 2608 15720 2672 15784
rect 2480 15639 2544 15703
rect 2608 15639 2672 15703
rect 2480 15558 2544 15622
rect 2608 15558 2672 15622
rect 2480 15477 2544 15541
rect 2608 15477 2672 15541
rect 2480 15396 2544 15460
rect 2608 15396 2672 15460
rect 2480 15315 2544 15379
rect 2608 15315 2672 15379
rect 2480 15234 2544 15298
rect 2608 15234 2672 15298
rect 2480 15153 2544 15217
rect 2608 15153 2672 15217
rect 2480 15072 2544 15136
rect 2608 15072 2672 15136
rect 2480 14991 2544 15055
rect 2608 14991 2672 15055
rect 2480 14910 2544 14974
rect 2608 14910 2672 14974
rect 2480 14829 2544 14893
rect 2608 14829 2672 14893
rect 2480 14748 2544 14812
rect 2608 14748 2672 14812
rect 2480 14667 2544 14731
rect 2608 14667 2672 14731
rect 2480 14586 2544 14650
rect 2608 14586 2672 14650
rect 2480 14505 2544 14569
rect 2608 14505 2672 14569
rect 2480 14424 2544 14488
rect 2608 14424 2672 14488
rect 2480 14343 2544 14407
rect 2608 14343 2672 14407
rect 2480 14262 2544 14326
rect 2608 14262 2672 14326
rect 2480 14181 2544 14245
rect 2608 14181 2672 14245
rect 2480 14100 2544 14164
rect 2608 14100 2672 14164
rect 2480 14019 2544 14083
rect 2608 14019 2672 14083
rect 2480 13938 2544 14002
rect 2608 13938 2672 14002
rect 2480 13857 2544 13921
rect 2608 13857 2672 13921
rect 2480 13776 2544 13840
rect 2608 13776 2672 13840
rect 2480 13695 2544 13759
rect 2608 13695 2672 13759
rect 2480 13614 2544 13678
rect 2608 13614 2672 13678
rect 2980 19609 3044 19673
rect 3100 19609 3164 19673
rect 2980 19517 3044 19581
rect 3100 19517 3164 19581
rect 2980 19425 3044 19489
rect 3100 19425 3164 19489
rect 2980 19333 3044 19397
rect 3100 19333 3164 19397
rect 2980 19241 3044 19305
rect 3100 19241 3164 19305
rect 2980 19148 3044 19212
rect 3100 19148 3164 19212
rect 5358 39528 5422 39592
rect 5486 39528 5550 39592
rect 5358 39448 5422 39512
rect 5486 39448 5550 39512
rect 5358 39368 5422 39432
rect 5486 39368 5550 39432
rect 5358 39288 5422 39352
rect 5486 39288 5550 39352
rect 5358 39208 5422 39272
rect 5486 39208 5550 39272
rect 5358 39128 5422 39192
rect 5486 39128 5550 39192
rect 5358 39048 5422 39112
rect 5486 39048 5550 39112
rect 5358 38968 5422 39032
rect 5486 38968 5550 39032
rect 5358 38888 5422 38952
rect 5486 38888 5550 38952
rect 5358 38808 5422 38872
rect 5486 38808 5550 38872
rect 5358 38728 5422 38792
rect 5486 38728 5550 38792
rect 5358 38648 5422 38712
rect 5486 38648 5550 38712
rect 5358 38568 5422 38632
rect 5486 38568 5550 38632
rect 5358 38488 5422 38552
rect 5486 38488 5550 38552
rect 5358 38408 5422 38472
rect 5486 38408 5550 38472
rect 5358 38328 5422 38392
rect 5486 38328 5550 38392
rect 5358 38247 5422 38311
rect 5486 38247 5550 38311
rect 5358 38166 5422 38230
rect 5486 38166 5550 38230
rect 5358 38085 5422 38149
rect 5486 38085 5550 38149
rect 5358 38004 5422 38068
rect 5486 38004 5550 38068
rect 5358 37923 5422 37987
rect 5486 37923 5550 37987
rect 5358 37842 5422 37906
rect 5486 37842 5550 37906
rect 5358 37761 5422 37825
rect 5486 37761 5550 37825
rect 5358 37680 5422 37744
rect 5486 37680 5550 37744
rect 5358 37599 5422 37663
rect 5486 37599 5550 37663
rect 5358 37518 5422 37582
rect 5486 37518 5550 37582
rect 5358 37437 5422 37501
rect 5486 37437 5550 37501
rect 5358 37356 5422 37420
rect 5486 37356 5550 37420
rect 5358 37275 5422 37339
rect 5486 37275 5550 37339
rect 5358 37194 5422 37258
rect 5486 37194 5550 37258
rect 5358 37113 5422 37177
rect 5486 37113 5550 37177
rect 5358 37032 5422 37096
rect 5486 37032 5550 37096
rect 5358 36951 5422 37015
rect 5486 36951 5550 37015
rect 5358 36870 5422 36934
rect 5486 36870 5550 36934
rect 5358 36789 5422 36853
rect 5486 36789 5550 36853
rect 5358 36708 5422 36772
rect 5486 36708 5550 36772
rect 5358 36627 5422 36691
rect 5486 36627 5550 36691
rect 5358 36546 5422 36610
rect 5486 36546 5550 36610
rect 5358 36465 5422 36529
rect 5486 36465 5550 36529
rect 5358 36384 5422 36448
rect 5486 36384 5550 36448
rect 5358 36303 5422 36367
rect 5486 36303 5550 36367
rect 5358 36222 5422 36286
rect 5486 36222 5550 36286
rect 5358 36141 5422 36205
rect 5486 36141 5550 36205
rect 5358 36060 5422 36124
rect 5486 36060 5550 36124
rect 5358 35979 5422 36043
rect 5486 35979 5550 36043
rect 5358 35898 5422 35962
rect 5486 35898 5550 35962
rect 5358 35817 5422 35881
rect 5486 35817 5550 35881
rect 5358 35736 5422 35800
rect 5486 35736 5550 35800
rect 5358 35655 5422 35719
rect 5486 35655 5550 35719
rect 5358 35574 5422 35638
rect 5486 35574 5550 35638
rect 5358 35493 5422 35557
rect 5486 35493 5550 35557
rect 5358 35412 5422 35476
rect 5486 35412 5550 35476
rect 5358 35331 5422 35395
rect 5486 35331 5550 35395
rect 5358 35250 5422 35314
rect 5486 35250 5550 35314
rect 5358 35169 5422 35233
rect 5486 35169 5550 35233
rect 5358 35088 5422 35152
rect 5486 35088 5550 35152
rect 5358 35007 5422 35071
rect 5486 35007 5550 35071
rect 5358 34926 5422 34990
rect 5486 34926 5550 34990
rect 5358 34845 5422 34909
rect 5486 34845 5550 34909
rect 5358 34764 5422 34828
rect 5486 34764 5550 34828
rect 4862 34155 4926 34219
rect 4990 34155 5054 34219
rect 4862 34061 4926 34125
rect 4990 34061 5054 34125
rect 4862 33966 4926 34030
rect 4990 33966 5054 34030
rect 4862 33871 4926 33935
rect 4990 33871 5054 33935
rect 4862 33776 4926 33840
rect 4990 33776 5054 33840
rect 4862 33681 4926 33745
rect 4990 33681 5054 33745
rect 3472 18528 3536 18592
rect 3600 18528 3664 18592
rect 3472 18448 3536 18512
rect 3600 18448 3664 18512
rect 3472 18368 3536 18432
rect 3600 18368 3664 18432
rect 3472 18288 3536 18352
rect 3600 18288 3664 18352
rect 3472 18208 3536 18272
rect 3600 18208 3664 18272
rect 3472 18128 3536 18192
rect 3600 18128 3664 18192
rect 3472 18048 3536 18112
rect 3600 18048 3664 18112
rect 3472 17968 3536 18032
rect 3600 17968 3664 18032
rect 3472 17888 3536 17952
rect 3600 17888 3664 17952
rect 3472 17808 3536 17872
rect 3600 17808 3664 17872
rect 3472 17728 3536 17792
rect 3600 17728 3664 17792
rect 3472 17648 3536 17712
rect 3600 17648 3664 17712
rect 3472 17568 3536 17632
rect 3600 17568 3664 17632
rect 3472 17488 3536 17552
rect 3600 17488 3664 17552
rect 3472 17408 3536 17472
rect 3600 17408 3664 17472
rect 3472 17328 3536 17392
rect 3600 17328 3664 17392
rect 3472 17248 3536 17312
rect 3600 17248 3664 17312
rect 3472 17168 3536 17232
rect 3600 17168 3664 17232
rect 3472 17088 3536 17152
rect 3600 17088 3664 17152
rect 3472 17008 3536 17072
rect 3600 17008 3664 17072
rect 3472 16928 3536 16992
rect 3600 16928 3664 16992
rect 3472 16848 3536 16912
rect 3600 16848 3664 16912
rect 3472 16768 3536 16832
rect 3600 16768 3664 16832
rect 3472 16688 3536 16752
rect 3600 16688 3664 16752
rect 3472 16608 3536 16672
rect 3600 16608 3664 16672
rect 3472 16528 3536 16592
rect 3600 16528 3664 16592
rect 3472 16448 3536 16512
rect 3600 16448 3664 16512
rect 3472 16368 3536 16432
rect 3600 16368 3664 16432
rect 3472 16287 3536 16351
rect 3600 16287 3664 16351
rect 3472 16206 3536 16270
rect 3600 16206 3664 16270
rect 3472 16125 3536 16189
rect 3600 16125 3664 16189
rect 3472 16044 3536 16108
rect 3600 16044 3664 16108
rect 3472 15963 3536 16027
rect 3600 15963 3664 16027
rect 3472 15882 3536 15946
rect 3600 15882 3664 15946
rect 3472 15801 3536 15865
rect 3600 15801 3664 15865
rect 3472 15720 3536 15784
rect 3600 15720 3664 15784
rect 3472 15639 3536 15703
rect 3600 15639 3664 15703
rect 3472 15558 3536 15622
rect 3600 15558 3664 15622
rect 3472 15477 3536 15541
rect 3600 15477 3664 15541
rect 3472 15396 3536 15460
rect 3600 15396 3664 15460
rect 3472 15315 3536 15379
rect 3600 15315 3664 15379
rect 3472 15234 3536 15298
rect 3600 15234 3664 15298
rect 3472 15153 3536 15217
rect 3600 15153 3664 15217
rect 3472 15072 3536 15136
rect 3600 15072 3664 15136
rect 3472 14991 3536 15055
rect 3600 14991 3664 15055
rect 3472 14910 3536 14974
rect 3600 14910 3664 14974
rect 3472 14829 3536 14893
rect 3600 14829 3664 14893
rect 3472 14748 3536 14812
rect 3600 14748 3664 14812
rect 3472 14667 3536 14731
rect 3600 14667 3664 14731
rect 3472 14586 3536 14650
rect 3600 14586 3664 14650
rect 3472 14505 3536 14569
rect 3600 14505 3664 14569
rect 3472 14424 3536 14488
rect 3600 14424 3664 14488
rect 3472 14343 3536 14407
rect 3600 14343 3664 14407
rect 3472 14262 3536 14326
rect 3600 14262 3664 14326
rect 3472 14181 3536 14245
rect 3600 14181 3664 14245
rect 3472 14100 3536 14164
rect 3600 14100 3664 14164
rect 3472 14019 3536 14083
rect 3600 14019 3664 14083
rect 3472 13938 3536 14002
rect 3600 13938 3664 14002
rect 3472 13857 3536 13921
rect 3600 13857 3664 13921
rect 3472 13776 3536 13840
rect 3600 13776 3664 13840
rect 3472 13695 3536 13759
rect 3600 13695 3664 13759
rect 3472 13614 3536 13678
rect 3600 13614 3664 13678
rect 3972 19609 4036 19673
rect 4092 19609 4156 19673
rect 3972 19517 4036 19581
rect 4092 19517 4156 19581
rect 3972 19424 4036 19488
rect 4092 19424 4156 19488
rect 3972 19331 4036 19395
rect 4092 19331 4156 19395
rect 3972 19238 4036 19302
rect 4092 19238 4156 19302
rect 3972 19145 4036 19209
rect 4092 19145 4156 19209
rect 6350 39528 6414 39592
rect 6478 39528 6542 39592
rect 6350 39448 6414 39512
rect 6478 39448 6542 39512
rect 6350 39368 6414 39432
rect 6478 39368 6542 39432
rect 6350 39288 6414 39352
rect 6478 39288 6542 39352
rect 6350 39208 6414 39272
rect 6478 39208 6542 39272
rect 6350 39128 6414 39192
rect 6478 39128 6542 39192
rect 6350 39048 6414 39112
rect 6478 39048 6542 39112
rect 6350 38968 6414 39032
rect 6478 38968 6542 39032
rect 6350 38888 6414 38952
rect 6478 38888 6542 38952
rect 6350 38808 6414 38872
rect 6478 38808 6542 38872
rect 6350 38728 6414 38792
rect 6478 38728 6542 38792
rect 6350 38648 6414 38712
rect 6478 38648 6542 38712
rect 6350 38568 6414 38632
rect 6478 38568 6542 38632
rect 6350 38488 6414 38552
rect 6478 38488 6542 38552
rect 6350 38408 6414 38472
rect 6478 38408 6542 38472
rect 6350 38328 6414 38392
rect 6478 38328 6542 38392
rect 6350 38247 6414 38311
rect 6478 38247 6542 38311
rect 6350 38166 6414 38230
rect 6478 38166 6542 38230
rect 6350 38085 6414 38149
rect 6478 38085 6542 38149
rect 6350 38004 6414 38068
rect 6478 38004 6542 38068
rect 6350 37923 6414 37987
rect 6478 37923 6542 37987
rect 6350 37842 6414 37906
rect 6478 37842 6542 37906
rect 6350 37761 6414 37825
rect 6478 37761 6542 37825
rect 6350 37680 6414 37744
rect 6478 37680 6542 37744
rect 6350 37599 6414 37663
rect 6478 37599 6542 37663
rect 6350 37518 6414 37582
rect 6478 37518 6542 37582
rect 6350 37437 6414 37501
rect 6478 37437 6542 37501
rect 6350 37356 6414 37420
rect 6478 37356 6542 37420
rect 6350 37275 6414 37339
rect 6478 37275 6542 37339
rect 6350 37194 6414 37258
rect 6478 37194 6542 37258
rect 6350 37113 6414 37177
rect 6478 37113 6542 37177
rect 6350 37032 6414 37096
rect 6478 37032 6542 37096
rect 6350 36951 6414 37015
rect 6478 36951 6542 37015
rect 6350 36870 6414 36934
rect 6478 36870 6542 36934
rect 6350 36789 6414 36853
rect 6478 36789 6542 36853
rect 6350 36708 6414 36772
rect 6478 36708 6542 36772
rect 6350 36627 6414 36691
rect 6478 36627 6542 36691
rect 6350 36546 6414 36610
rect 6478 36546 6542 36610
rect 6350 36465 6414 36529
rect 6478 36465 6542 36529
rect 6350 36384 6414 36448
rect 6478 36384 6542 36448
rect 6350 36303 6414 36367
rect 6478 36303 6542 36367
rect 6350 36222 6414 36286
rect 6478 36222 6542 36286
rect 6350 36141 6414 36205
rect 6478 36141 6542 36205
rect 6350 36060 6414 36124
rect 6478 36060 6542 36124
rect 6350 35979 6414 36043
rect 6478 35979 6542 36043
rect 6350 35898 6414 35962
rect 6478 35898 6542 35962
rect 6350 35817 6414 35881
rect 6478 35817 6542 35881
rect 6350 35736 6414 35800
rect 6478 35736 6542 35800
rect 6350 35655 6414 35719
rect 6478 35655 6542 35719
rect 6350 35574 6414 35638
rect 6478 35574 6542 35638
rect 6350 35493 6414 35557
rect 6478 35493 6542 35557
rect 6350 35412 6414 35476
rect 6478 35412 6542 35476
rect 6350 35331 6414 35395
rect 6478 35331 6542 35395
rect 6350 35250 6414 35314
rect 6478 35250 6542 35314
rect 6350 35169 6414 35233
rect 6478 35169 6542 35233
rect 6350 35088 6414 35152
rect 6478 35088 6542 35152
rect 6350 35007 6414 35071
rect 6478 35007 6542 35071
rect 6350 34926 6414 34990
rect 6478 34926 6542 34990
rect 6350 34845 6414 34909
rect 6478 34845 6542 34909
rect 6350 34764 6414 34828
rect 6478 34764 6542 34828
rect 5854 34155 5918 34219
rect 5982 34155 6046 34219
rect 5854 34061 5918 34125
rect 5982 34061 6046 34125
rect 5854 33966 5918 34030
rect 5982 33966 6046 34030
rect 5854 33871 5918 33935
rect 5982 33871 6046 33935
rect 5854 33776 5918 33840
rect 5982 33776 6046 33840
rect 5854 33681 5918 33745
rect 5982 33681 6046 33745
rect 4464 18528 4528 18592
rect 4592 18528 4656 18592
rect 4464 18448 4528 18512
rect 4592 18448 4656 18512
rect 4464 18368 4528 18432
rect 4592 18368 4656 18432
rect 4464 18288 4528 18352
rect 4592 18288 4656 18352
rect 4464 18208 4528 18272
rect 4592 18208 4656 18272
rect 4464 18128 4528 18192
rect 4592 18128 4656 18192
rect 4464 18048 4528 18112
rect 4592 18048 4656 18112
rect 4464 17968 4528 18032
rect 4592 17968 4656 18032
rect 4464 17888 4528 17952
rect 4592 17888 4656 17952
rect 4464 17808 4528 17872
rect 4592 17808 4656 17872
rect 4464 17728 4528 17792
rect 4592 17728 4656 17792
rect 4464 17648 4528 17712
rect 4592 17648 4656 17712
rect 4464 17568 4528 17632
rect 4592 17568 4656 17632
rect 4464 17488 4528 17552
rect 4592 17488 4656 17552
rect 4464 17408 4528 17472
rect 4592 17408 4656 17472
rect 4464 17328 4528 17392
rect 4592 17328 4656 17392
rect 4464 17248 4528 17312
rect 4592 17248 4656 17312
rect 4464 17168 4528 17232
rect 4592 17168 4656 17232
rect 4464 17088 4528 17152
rect 4592 17088 4656 17152
rect 4464 17008 4528 17072
rect 4592 17008 4656 17072
rect 4464 16928 4528 16992
rect 4592 16928 4656 16992
rect 4464 16848 4528 16912
rect 4592 16848 4656 16912
rect 4464 16768 4528 16832
rect 4592 16768 4656 16832
rect 4464 16688 4528 16752
rect 4592 16688 4656 16752
rect 4464 16608 4528 16672
rect 4592 16608 4656 16672
rect 4464 16528 4528 16592
rect 4592 16528 4656 16592
rect 4464 16448 4528 16512
rect 4592 16448 4656 16512
rect 4464 16368 4528 16432
rect 4592 16368 4656 16432
rect 4464 16287 4528 16351
rect 4592 16287 4656 16351
rect 4464 16206 4528 16270
rect 4592 16206 4656 16270
rect 4464 16125 4528 16189
rect 4592 16125 4656 16189
rect 4464 16044 4528 16108
rect 4592 16044 4656 16108
rect 4464 15963 4528 16027
rect 4592 15963 4656 16027
rect 4464 15882 4528 15946
rect 4592 15882 4656 15946
rect 4464 15801 4528 15865
rect 4592 15801 4656 15865
rect 4464 15720 4528 15784
rect 4592 15720 4656 15784
rect 4464 15639 4528 15703
rect 4592 15639 4656 15703
rect 4464 15558 4528 15622
rect 4592 15558 4656 15622
rect 4464 15477 4528 15541
rect 4592 15477 4656 15541
rect 4464 15396 4528 15460
rect 4592 15396 4656 15460
rect 4464 15315 4528 15379
rect 4592 15315 4656 15379
rect 4464 15234 4528 15298
rect 4592 15234 4656 15298
rect 4464 15153 4528 15217
rect 4592 15153 4656 15217
rect 4464 15072 4528 15136
rect 4592 15072 4656 15136
rect 4464 14991 4528 15055
rect 4592 14991 4656 15055
rect 4464 14910 4528 14974
rect 4592 14910 4656 14974
rect 4464 14829 4528 14893
rect 4592 14829 4656 14893
rect 4464 14748 4528 14812
rect 4592 14748 4656 14812
rect 4464 14667 4528 14731
rect 4592 14667 4656 14731
rect 4464 14586 4528 14650
rect 4592 14586 4656 14650
rect 4464 14505 4528 14569
rect 4592 14505 4656 14569
rect 4464 14424 4528 14488
rect 4592 14424 4656 14488
rect 4464 14343 4528 14407
rect 4592 14343 4656 14407
rect 4464 14262 4528 14326
rect 4592 14262 4656 14326
rect 4464 14181 4528 14245
rect 4592 14181 4656 14245
rect 4464 14100 4528 14164
rect 4592 14100 4656 14164
rect 4464 14019 4528 14083
rect 4592 14019 4656 14083
rect 4464 13938 4528 14002
rect 4592 13938 4656 14002
rect 4464 13857 4528 13921
rect 4592 13857 4656 13921
rect 4464 13776 4528 13840
rect 4592 13776 4656 13840
rect 4464 13695 4528 13759
rect 4592 13695 4656 13759
rect 4464 13614 4528 13678
rect 4592 13614 4656 13678
rect 4964 19609 5028 19673
rect 5084 19609 5148 19673
rect 4964 19517 5028 19581
rect 5084 19517 5148 19581
rect 4964 19425 5028 19489
rect 5084 19425 5148 19489
rect 4964 19333 5028 19397
rect 5084 19333 5148 19397
rect 4964 19241 5028 19305
rect 5084 19241 5148 19305
rect 4964 19148 5028 19212
rect 5084 19148 5148 19212
rect 7342 39528 7406 39592
rect 7470 39528 7534 39592
rect 7342 39448 7406 39512
rect 7470 39448 7534 39512
rect 7342 39368 7406 39432
rect 7470 39368 7534 39432
rect 7342 39288 7406 39352
rect 7470 39288 7534 39352
rect 7342 39208 7406 39272
rect 7470 39208 7534 39272
rect 7342 39128 7406 39192
rect 7470 39128 7534 39192
rect 7342 39048 7406 39112
rect 7470 39048 7534 39112
rect 7342 38968 7406 39032
rect 7470 38968 7534 39032
rect 7342 38888 7406 38952
rect 7470 38888 7534 38952
rect 7342 38808 7406 38872
rect 7470 38808 7534 38872
rect 7342 38728 7406 38792
rect 7470 38728 7534 38792
rect 7342 38648 7406 38712
rect 7470 38648 7534 38712
rect 7342 38568 7406 38632
rect 7470 38568 7534 38632
rect 7342 38488 7406 38552
rect 7470 38488 7534 38552
rect 7342 38408 7406 38472
rect 7470 38408 7534 38472
rect 7342 38328 7406 38392
rect 7470 38328 7534 38392
rect 7342 38247 7406 38311
rect 7470 38247 7534 38311
rect 7342 38166 7406 38230
rect 7470 38166 7534 38230
rect 7342 38085 7406 38149
rect 7470 38085 7534 38149
rect 7342 38004 7406 38068
rect 7470 38004 7534 38068
rect 7342 37923 7406 37987
rect 7470 37923 7534 37987
rect 7342 37842 7406 37906
rect 7470 37842 7534 37906
rect 7342 37761 7406 37825
rect 7470 37761 7534 37825
rect 7342 37680 7406 37744
rect 7470 37680 7534 37744
rect 7342 37599 7406 37663
rect 7470 37599 7534 37663
rect 7342 37518 7406 37582
rect 7470 37518 7534 37582
rect 7342 37437 7406 37501
rect 7470 37437 7534 37501
rect 7342 37356 7406 37420
rect 7470 37356 7534 37420
rect 7342 37275 7406 37339
rect 7470 37275 7534 37339
rect 7342 37194 7406 37258
rect 7470 37194 7534 37258
rect 7342 37113 7406 37177
rect 7470 37113 7534 37177
rect 7342 37032 7406 37096
rect 7470 37032 7534 37096
rect 7342 36951 7406 37015
rect 7470 36951 7534 37015
rect 7342 36870 7406 36934
rect 7470 36870 7534 36934
rect 7342 36789 7406 36853
rect 7470 36789 7534 36853
rect 7342 36708 7406 36772
rect 7470 36708 7534 36772
rect 7342 36627 7406 36691
rect 7470 36627 7534 36691
rect 7342 36546 7406 36610
rect 7470 36546 7534 36610
rect 7342 36465 7406 36529
rect 7470 36465 7534 36529
rect 7342 36384 7406 36448
rect 7470 36384 7534 36448
rect 7342 36303 7406 36367
rect 7470 36303 7534 36367
rect 7342 36222 7406 36286
rect 7470 36222 7534 36286
rect 7342 36141 7406 36205
rect 7470 36141 7534 36205
rect 7342 36060 7406 36124
rect 7470 36060 7534 36124
rect 7342 35979 7406 36043
rect 7470 35979 7534 36043
rect 7342 35898 7406 35962
rect 7470 35898 7534 35962
rect 7342 35817 7406 35881
rect 7470 35817 7534 35881
rect 7342 35736 7406 35800
rect 7470 35736 7534 35800
rect 7342 35655 7406 35719
rect 7470 35655 7534 35719
rect 7342 35574 7406 35638
rect 7470 35574 7534 35638
rect 7342 35493 7406 35557
rect 7470 35493 7534 35557
rect 7342 35412 7406 35476
rect 7470 35412 7534 35476
rect 7342 35331 7406 35395
rect 7470 35331 7534 35395
rect 7342 35250 7406 35314
rect 7470 35250 7534 35314
rect 7342 35169 7406 35233
rect 7470 35169 7534 35233
rect 7342 35088 7406 35152
rect 7470 35088 7534 35152
rect 7342 35007 7406 35071
rect 7470 35007 7534 35071
rect 7342 34926 7406 34990
rect 7470 34926 7534 34990
rect 7342 34845 7406 34909
rect 7470 34845 7534 34909
rect 7342 34764 7406 34828
rect 7470 34764 7534 34828
rect 6846 34155 6910 34219
rect 6974 34155 7038 34219
rect 6846 34061 6910 34125
rect 6974 34061 7038 34125
rect 6846 33966 6910 34030
rect 6974 33966 7038 34030
rect 6846 33871 6910 33935
rect 6974 33871 7038 33935
rect 6846 33776 6910 33840
rect 6974 33776 7038 33840
rect 6846 33681 6910 33745
rect 6974 33681 7038 33745
rect 5456 18528 5520 18592
rect 5584 18528 5648 18592
rect 5456 18448 5520 18512
rect 5584 18448 5648 18512
rect 5456 18368 5520 18432
rect 5584 18368 5648 18432
rect 5456 18288 5520 18352
rect 5584 18288 5648 18352
rect 5456 18208 5520 18272
rect 5584 18208 5648 18272
rect 5456 18128 5520 18192
rect 5584 18128 5648 18192
rect 5456 18048 5520 18112
rect 5584 18048 5648 18112
rect 5456 17968 5520 18032
rect 5584 17968 5648 18032
rect 5456 17888 5520 17952
rect 5584 17888 5648 17952
rect 5456 17808 5520 17872
rect 5584 17808 5648 17872
rect 5456 17728 5520 17792
rect 5584 17728 5648 17792
rect 5456 17648 5520 17712
rect 5584 17648 5648 17712
rect 5456 17568 5520 17632
rect 5584 17568 5648 17632
rect 5456 17488 5520 17552
rect 5584 17488 5648 17552
rect 5456 17408 5520 17472
rect 5584 17408 5648 17472
rect 5456 17328 5520 17392
rect 5584 17328 5648 17392
rect 5456 17248 5520 17312
rect 5584 17248 5648 17312
rect 5456 17168 5520 17232
rect 5584 17168 5648 17232
rect 5456 17088 5520 17152
rect 5584 17088 5648 17152
rect 5456 17008 5520 17072
rect 5584 17008 5648 17072
rect 5456 16928 5520 16992
rect 5584 16928 5648 16992
rect 5456 16848 5520 16912
rect 5584 16848 5648 16912
rect 5456 16768 5520 16832
rect 5584 16768 5648 16832
rect 5456 16688 5520 16752
rect 5584 16688 5648 16752
rect 5456 16608 5520 16672
rect 5584 16608 5648 16672
rect 5456 16528 5520 16592
rect 5584 16528 5648 16592
rect 5456 16448 5520 16512
rect 5584 16448 5648 16512
rect 5456 16367 5520 16431
rect 5584 16367 5648 16431
rect 5456 16286 5520 16350
rect 5584 16286 5648 16350
rect 5456 16205 5520 16269
rect 5584 16205 5648 16269
rect 5456 16124 5520 16188
rect 5584 16124 5648 16188
rect 5456 16043 5520 16107
rect 5584 16043 5648 16107
rect 5456 15962 5520 16026
rect 5584 15962 5648 16026
rect 5456 15881 5520 15945
rect 5584 15881 5648 15945
rect 5456 15800 5520 15864
rect 5584 15800 5648 15864
rect 5456 15719 5520 15783
rect 5584 15719 5648 15783
rect 5456 15638 5520 15702
rect 5584 15638 5648 15702
rect 5456 15557 5520 15621
rect 5584 15557 5648 15621
rect 5456 15476 5520 15540
rect 5584 15476 5648 15540
rect 5456 15395 5520 15459
rect 5584 15395 5648 15459
rect 5456 15314 5520 15378
rect 5584 15314 5648 15378
rect 5456 15233 5520 15297
rect 5584 15233 5648 15297
rect 5456 15152 5520 15216
rect 5584 15152 5648 15216
rect 5456 15071 5520 15135
rect 5584 15071 5648 15135
rect 5456 14990 5520 15054
rect 5584 14990 5648 15054
rect 5456 14909 5520 14973
rect 5584 14909 5648 14973
rect 5456 14828 5520 14892
rect 5584 14828 5648 14892
rect 5456 14747 5520 14811
rect 5584 14747 5648 14811
rect 5456 14666 5520 14730
rect 5584 14666 5648 14730
rect 5456 14585 5520 14649
rect 5584 14585 5648 14649
rect 5456 14504 5520 14568
rect 5584 14504 5648 14568
rect 5456 14423 5520 14487
rect 5584 14423 5648 14487
rect 5456 14342 5520 14406
rect 5584 14342 5648 14406
rect 5456 14261 5520 14325
rect 5584 14261 5648 14325
rect 5456 14180 5520 14244
rect 5584 14180 5648 14244
rect 5456 14099 5520 14163
rect 5584 14099 5648 14163
rect 5456 14018 5520 14082
rect 5584 14018 5648 14082
rect 5456 13937 5520 14001
rect 5584 13937 5648 14001
rect 5456 13856 5520 13920
rect 5584 13856 5648 13920
rect 5456 13775 5520 13839
rect 5584 13775 5648 13839
rect 5456 13694 5520 13758
rect 5584 13694 5648 13758
rect 5456 13613 5520 13677
rect 5584 13613 5648 13677
rect 5953 19609 6017 19673
rect 6073 19609 6137 19673
rect 5953 19517 6017 19581
rect 6073 19517 6137 19581
rect 5953 19425 6017 19489
rect 6073 19425 6137 19489
rect 5953 19333 6017 19397
rect 6073 19333 6137 19397
rect 5953 19241 6017 19305
rect 6073 19241 6137 19305
rect 5953 19148 6017 19212
rect 6073 19148 6137 19212
rect 8334 39528 8398 39592
rect 8462 39528 8526 39592
rect 8334 39448 8398 39512
rect 8462 39448 8526 39512
rect 8334 39368 8398 39432
rect 8462 39368 8526 39432
rect 8334 39288 8398 39352
rect 8462 39288 8526 39352
rect 8334 39208 8398 39272
rect 8462 39208 8526 39272
rect 8334 39128 8398 39192
rect 8462 39128 8526 39192
rect 8334 39048 8398 39112
rect 8462 39048 8526 39112
rect 8334 38968 8398 39032
rect 8462 38968 8526 39032
rect 8334 38888 8398 38952
rect 8462 38888 8526 38952
rect 8334 38808 8398 38872
rect 8462 38808 8526 38872
rect 8334 38728 8398 38792
rect 8462 38728 8526 38792
rect 8334 38648 8398 38712
rect 8462 38648 8526 38712
rect 8334 38568 8398 38632
rect 8462 38568 8526 38632
rect 8334 38488 8398 38552
rect 8462 38488 8526 38552
rect 8334 38408 8398 38472
rect 8462 38408 8526 38472
rect 8334 38328 8398 38392
rect 8462 38328 8526 38392
rect 8334 38247 8398 38311
rect 8462 38247 8526 38311
rect 8334 38166 8398 38230
rect 8462 38166 8526 38230
rect 8334 38085 8398 38149
rect 8462 38085 8526 38149
rect 8334 38004 8398 38068
rect 8462 38004 8526 38068
rect 8334 37923 8398 37987
rect 8462 37923 8526 37987
rect 8334 37842 8398 37906
rect 8462 37842 8526 37906
rect 8334 37761 8398 37825
rect 8462 37761 8526 37825
rect 8334 37680 8398 37744
rect 8462 37680 8526 37744
rect 8334 37599 8398 37663
rect 8462 37599 8526 37663
rect 8334 37518 8398 37582
rect 8462 37518 8526 37582
rect 8334 37437 8398 37501
rect 8462 37437 8526 37501
rect 8334 37356 8398 37420
rect 8462 37356 8526 37420
rect 8334 37275 8398 37339
rect 8462 37275 8526 37339
rect 8334 37194 8398 37258
rect 8462 37194 8526 37258
rect 8334 37113 8398 37177
rect 8462 37113 8526 37177
rect 8334 37032 8398 37096
rect 8462 37032 8526 37096
rect 8334 36951 8398 37015
rect 8462 36951 8526 37015
rect 8334 36870 8398 36934
rect 8462 36870 8526 36934
rect 8334 36789 8398 36853
rect 8462 36789 8526 36853
rect 8334 36708 8398 36772
rect 8462 36708 8526 36772
rect 8334 36627 8398 36691
rect 8462 36627 8526 36691
rect 8334 36546 8398 36610
rect 8462 36546 8526 36610
rect 8334 36465 8398 36529
rect 8462 36465 8526 36529
rect 8334 36384 8398 36448
rect 8462 36384 8526 36448
rect 8334 36303 8398 36367
rect 8462 36303 8526 36367
rect 8334 36222 8398 36286
rect 8462 36222 8526 36286
rect 8334 36141 8398 36205
rect 8462 36141 8526 36205
rect 8334 36060 8398 36124
rect 8462 36060 8526 36124
rect 8334 35979 8398 36043
rect 8462 35979 8526 36043
rect 8334 35898 8398 35962
rect 8462 35898 8526 35962
rect 8334 35817 8398 35881
rect 8462 35817 8526 35881
rect 8334 35736 8398 35800
rect 8462 35736 8526 35800
rect 8334 35655 8398 35719
rect 8462 35655 8526 35719
rect 8334 35574 8398 35638
rect 8462 35574 8526 35638
rect 8334 35493 8398 35557
rect 8462 35493 8526 35557
rect 8334 35412 8398 35476
rect 8462 35412 8526 35476
rect 8334 35331 8398 35395
rect 8462 35331 8526 35395
rect 8334 35250 8398 35314
rect 8462 35250 8526 35314
rect 8334 35169 8398 35233
rect 8462 35169 8526 35233
rect 8334 35088 8398 35152
rect 8462 35088 8526 35152
rect 8334 35007 8398 35071
rect 8462 35007 8526 35071
rect 8334 34926 8398 34990
rect 8462 34926 8526 34990
rect 8334 34845 8398 34909
rect 8462 34845 8526 34909
rect 8334 34764 8398 34828
rect 8462 34764 8526 34828
rect 7838 34155 7902 34219
rect 7966 34155 8030 34219
rect 7838 34061 7902 34125
rect 7966 34061 8030 34125
rect 7838 33966 7902 34030
rect 7966 33966 8030 34030
rect 7838 33871 7902 33935
rect 7966 33871 8030 33935
rect 7838 33776 7902 33840
rect 7966 33776 8030 33840
rect 7838 33681 7902 33745
rect 7966 33681 8030 33745
rect 6448 18528 6512 18592
rect 6576 18528 6640 18592
rect 6448 18448 6512 18512
rect 6576 18448 6640 18512
rect 6448 18368 6512 18432
rect 6576 18368 6640 18432
rect 6448 18288 6512 18352
rect 6576 18288 6640 18352
rect 6448 18208 6512 18272
rect 6576 18208 6640 18272
rect 6448 18128 6512 18192
rect 6576 18128 6640 18192
rect 6448 18048 6512 18112
rect 6576 18048 6640 18112
rect 6448 17968 6512 18032
rect 6576 17968 6640 18032
rect 6448 17888 6512 17952
rect 6576 17888 6640 17952
rect 6448 17808 6512 17872
rect 6576 17808 6640 17872
rect 6448 17728 6512 17792
rect 6576 17728 6640 17792
rect 6448 17648 6512 17712
rect 6576 17648 6640 17712
rect 6448 17568 6512 17632
rect 6576 17568 6640 17632
rect 6448 17488 6512 17552
rect 6576 17488 6640 17552
rect 6448 17408 6512 17472
rect 6576 17408 6640 17472
rect 6448 17328 6512 17392
rect 6576 17328 6640 17392
rect 6448 17248 6512 17312
rect 6576 17248 6640 17312
rect 6448 17168 6512 17232
rect 6576 17168 6640 17232
rect 6448 17088 6512 17152
rect 6576 17088 6640 17152
rect 6448 17008 6512 17072
rect 6576 17008 6640 17072
rect 6448 16928 6512 16992
rect 6576 16928 6640 16992
rect 6448 16848 6512 16912
rect 6576 16848 6640 16912
rect 6448 16768 6512 16832
rect 6576 16768 6640 16832
rect 6448 16688 6512 16752
rect 6576 16688 6640 16752
rect 6448 16608 6512 16672
rect 6576 16608 6640 16672
rect 6448 16528 6512 16592
rect 6576 16528 6640 16592
rect 6448 16448 6512 16512
rect 6576 16448 6640 16512
rect 6448 16368 6512 16432
rect 6576 16368 6640 16432
rect 6448 16287 6512 16351
rect 6576 16287 6640 16351
rect 6448 16206 6512 16270
rect 6576 16206 6640 16270
rect 6448 16125 6512 16189
rect 6576 16125 6640 16189
rect 6448 16044 6512 16108
rect 6576 16044 6640 16108
rect 6448 15963 6512 16027
rect 6576 15963 6640 16027
rect 6448 15882 6512 15946
rect 6576 15882 6640 15946
rect 6448 15801 6512 15865
rect 6576 15801 6640 15865
rect 6448 15720 6512 15784
rect 6576 15720 6640 15784
rect 6448 15639 6512 15703
rect 6576 15639 6640 15703
rect 6448 15558 6512 15622
rect 6576 15558 6640 15622
rect 6448 15477 6512 15541
rect 6576 15477 6640 15541
rect 6448 15396 6512 15460
rect 6576 15396 6640 15460
rect 6448 15315 6512 15379
rect 6576 15315 6640 15379
rect 6448 15234 6512 15298
rect 6576 15234 6640 15298
rect 6448 15153 6512 15217
rect 6576 15153 6640 15217
rect 6448 15072 6512 15136
rect 6576 15072 6640 15136
rect 6448 14991 6512 15055
rect 6576 14991 6640 15055
rect 6448 14910 6512 14974
rect 6576 14910 6640 14974
rect 6448 14829 6512 14893
rect 6576 14829 6640 14893
rect 6448 14748 6512 14812
rect 6576 14748 6640 14812
rect 6448 14667 6512 14731
rect 6576 14667 6640 14731
rect 6448 14586 6512 14650
rect 6576 14586 6640 14650
rect 6448 14505 6512 14569
rect 6576 14505 6640 14569
rect 6448 14424 6512 14488
rect 6576 14424 6640 14488
rect 6448 14343 6512 14407
rect 6576 14343 6640 14407
rect 6448 14262 6512 14326
rect 6576 14262 6640 14326
rect 6448 14181 6512 14245
rect 6576 14181 6640 14245
rect 6448 14100 6512 14164
rect 6576 14100 6640 14164
rect 6448 14019 6512 14083
rect 6576 14019 6640 14083
rect 6448 13938 6512 14002
rect 6576 13938 6640 14002
rect 6448 13857 6512 13921
rect 6576 13857 6640 13921
rect 6448 13776 6512 13840
rect 6576 13776 6640 13840
rect 6448 13695 6512 13759
rect 6576 13695 6640 13759
rect 6448 13614 6512 13678
rect 6576 13614 6640 13678
rect 6945 19609 7009 19673
rect 7065 19609 7129 19673
rect 6945 19517 7009 19581
rect 7065 19517 7129 19581
rect 6945 19425 7009 19489
rect 7065 19425 7129 19489
rect 6945 19333 7009 19397
rect 7065 19333 7129 19397
rect 6945 19241 7009 19305
rect 7065 19241 7129 19305
rect 6945 19148 7009 19212
rect 7065 19148 7129 19212
rect 9326 39528 9390 39592
rect 9454 39528 9518 39592
rect 9326 39448 9390 39512
rect 9454 39448 9518 39512
rect 9326 39368 9390 39432
rect 9454 39368 9518 39432
rect 9326 39288 9390 39352
rect 9454 39288 9518 39352
rect 9326 39208 9390 39272
rect 9454 39208 9518 39272
rect 9326 39128 9390 39192
rect 9454 39128 9518 39192
rect 9326 39048 9390 39112
rect 9454 39048 9518 39112
rect 9326 38968 9390 39032
rect 9454 38968 9518 39032
rect 9326 38888 9390 38952
rect 9454 38888 9518 38952
rect 9326 38808 9390 38872
rect 9454 38808 9518 38872
rect 9326 38728 9390 38792
rect 9454 38728 9518 38792
rect 9326 38648 9390 38712
rect 9454 38648 9518 38712
rect 9326 38568 9390 38632
rect 9454 38568 9518 38632
rect 9326 38488 9390 38552
rect 9454 38488 9518 38552
rect 9326 38408 9390 38472
rect 9454 38408 9518 38472
rect 9326 38328 9390 38392
rect 9454 38328 9518 38392
rect 9326 38247 9390 38311
rect 9454 38247 9518 38311
rect 9326 38166 9390 38230
rect 9454 38166 9518 38230
rect 9326 38085 9390 38149
rect 9454 38085 9518 38149
rect 9326 38004 9390 38068
rect 9454 38004 9518 38068
rect 9326 37923 9390 37987
rect 9454 37923 9518 37987
rect 9326 37842 9390 37906
rect 9454 37842 9518 37906
rect 9326 37761 9390 37825
rect 9454 37761 9518 37825
rect 9326 37680 9390 37744
rect 9454 37680 9518 37744
rect 9326 37599 9390 37663
rect 9454 37599 9518 37663
rect 9326 37518 9390 37582
rect 9454 37518 9518 37582
rect 9326 37437 9390 37501
rect 9454 37437 9518 37501
rect 9326 37356 9390 37420
rect 9454 37356 9518 37420
rect 9326 37275 9390 37339
rect 9454 37275 9518 37339
rect 9326 37194 9390 37258
rect 9454 37194 9518 37258
rect 9326 37113 9390 37177
rect 9454 37113 9518 37177
rect 9326 37032 9390 37096
rect 9454 37032 9518 37096
rect 9326 36951 9390 37015
rect 9454 36951 9518 37015
rect 9326 36870 9390 36934
rect 9454 36870 9518 36934
rect 9326 36789 9390 36853
rect 9454 36789 9518 36853
rect 9326 36708 9390 36772
rect 9454 36708 9518 36772
rect 9326 36627 9390 36691
rect 9454 36627 9518 36691
rect 9326 36546 9390 36610
rect 9454 36546 9518 36610
rect 9326 36465 9390 36529
rect 9454 36465 9518 36529
rect 9326 36384 9390 36448
rect 9454 36384 9518 36448
rect 9326 36303 9390 36367
rect 9454 36303 9518 36367
rect 9326 36222 9390 36286
rect 9454 36222 9518 36286
rect 9326 36141 9390 36205
rect 9454 36141 9518 36205
rect 9326 36060 9390 36124
rect 9454 36060 9518 36124
rect 9326 35979 9390 36043
rect 9454 35979 9518 36043
rect 9326 35898 9390 35962
rect 9454 35898 9518 35962
rect 9326 35817 9390 35881
rect 9454 35817 9518 35881
rect 9326 35736 9390 35800
rect 9454 35736 9518 35800
rect 9326 35655 9390 35719
rect 9454 35655 9518 35719
rect 9326 35574 9390 35638
rect 9454 35574 9518 35638
rect 9326 35493 9390 35557
rect 9454 35493 9518 35557
rect 9326 35412 9390 35476
rect 9454 35412 9518 35476
rect 9326 35331 9390 35395
rect 9454 35331 9518 35395
rect 9326 35250 9390 35314
rect 9454 35250 9518 35314
rect 9326 35169 9390 35233
rect 9454 35169 9518 35233
rect 9326 35088 9390 35152
rect 9454 35088 9518 35152
rect 9326 35007 9390 35071
rect 9454 35007 9518 35071
rect 9326 34926 9390 34990
rect 9454 34926 9518 34990
rect 9326 34845 9390 34909
rect 9454 34845 9518 34909
rect 9326 34764 9390 34828
rect 9454 34764 9518 34828
rect 8830 34155 8894 34219
rect 8958 34155 9022 34219
rect 8830 34061 8894 34125
rect 8958 34061 9022 34125
rect 8830 33966 8894 34030
rect 8958 33966 9022 34030
rect 8830 33871 8894 33935
rect 8958 33871 9022 33935
rect 8830 33776 8894 33840
rect 8958 33776 9022 33840
rect 8830 33681 8894 33745
rect 8958 33681 9022 33745
rect 7440 18528 7504 18592
rect 7568 18528 7632 18592
rect 7440 18448 7504 18512
rect 7568 18448 7632 18512
rect 7440 18368 7504 18432
rect 7568 18368 7632 18432
rect 7440 18288 7504 18352
rect 7568 18288 7632 18352
rect 7440 18208 7504 18272
rect 7568 18208 7632 18272
rect 7440 18128 7504 18192
rect 7568 18128 7632 18192
rect 7440 18048 7504 18112
rect 7568 18048 7632 18112
rect 7440 17968 7504 18032
rect 7568 17968 7632 18032
rect 7440 17888 7504 17952
rect 7568 17888 7632 17952
rect 7440 17808 7504 17872
rect 7568 17808 7632 17872
rect 7440 17728 7504 17792
rect 7568 17728 7632 17792
rect 7440 17648 7504 17712
rect 7568 17648 7632 17712
rect 7440 17568 7504 17632
rect 7568 17568 7632 17632
rect 7440 17488 7504 17552
rect 7568 17488 7632 17552
rect 7440 17408 7504 17472
rect 7568 17408 7632 17472
rect 7440 17328 7504 17392
rect 7568 17328 7632 17392
rect 7440 17248 7504 17312
rect 7568 17248 7632 17312
rect 7440 17168 7504 17232
rect 7568 17168 7632 17232
rect 7440 17088 7504 17152
rect 7568 17088 7632 17152
rect 7440 17008 7504 17072
rect 7568 17008 7632 17072
rect 7440 16928 7504 16992
rect 7568 16928 7632 16992
rect 7440 16848 7504 16912
rect 7568 16848 7632 16912
rect 7440 16768 7504 16832
rect 7568 16768 7632 16832
rect 7440 16688 7504 16752
rect 7568 16688 7632 16752
rect 7440 16608 7504 16672
rect 7568 16608 7632 16672
rect 7440 16528 7504 16592
rect 7568 16528 7632 16592
rect 7440 16448 7504 16512
rect 7568 16448 7632 16512
rect 7440 16368 7504 16432
rect 7568 16368 7632 16432
rect 7440 16287 7504 16351
rect 7568 16287 7632 16351
rect 7440 16206 7504 16270
rect 7568 16206 7632 16270
rect 7440 16125 7504 16189
rect 7568 16125 7632 16189
rect 7440 16044 7504 16108
rect 7568 16044 7632 16108
rect 7440 15963 7504 16027
rect 7568 15963 7632 16027
rect 7440 15882 7504 15946
rect 7568 15882 7632 15946
rect 7440 15801 7504 15865
rect 7568 15801 7632 15865
rect 7440 15720 7504 15784
rect 7568 15720 7632 15784
rect 7440 15639 7504 15703
rect 7568 15639 7632 15703
rect 7440 15558 7504 15622
rect 7568 15558 7632 15622
rect 7440 15477 7504 15541
rect 7568 15477 7632 15541
rect 7440 15396 7504 15460
rect 7568 15396 7632 15460
rect 7440 15315 7504 15379
rect 7568 15315 7632 15379
rect 7440 15234 7504 15298
rect 7568 15234 7632 15298
rect 7440 15153 7504 15217
rect 7568 15153 7632 15217
rect 7440 15072 7504 15136
rect 7568 15072 7632 15136
rect 7440 14991 7504 15055
rect 7568 14991 7632 15055
rect 7440 14910 7504 14974
rect 7568 14910 7632 14974
rect 7440 14829 7504 14893
rect 7568 14829 7632 14893
rect 7440 14748 7504 14812
rect 7568 14748 7632 14812
rect 7440 14667 7504 14731
rect 7568 14667 7632 14731
rect 7440 14586 7504 14650
rect 7568 14586 7632 14650
rect 7440 14505 7504 14569
rect 7568 14505 7632 14569
rect 7440 14424 7504 14488
rect 7568 14424 7632 14488
rect 7440 14343 7504 14407
rect 7568 14343 7632 14407
rect 7440 14262 7504 14326
rect 7568 14262 7632 14326
rect 7440 14181 7504 14245
rect 7568 14181 7632 14245
rect 7440 14100 7504 14164
rect 7568 14100 7632 14164
rect 7440 14019 7504 14083
rect 7568 14019 7632 14083
rect 7440 13938 7504 14002
rect 7568 13938 7632 14002
rect 7440 13857 7504 13921
rect 7568 13857 7632 13921
rect 7440 13776 7504 13840
rect 7568 13776 7632 13840
rect 7440 13695 7504 13759
rect 7568 13695 7632 13759
rect 7440 13614 7504 13678
rect 7568 13614 7632 13678
rect 7940 19609 8004 19673
rect 8060 19609 8124 19673
rect 7940 19517 8004 19581
rect 8060 19517 8124 19581
rect 7940 19425 8004 19489
rect 8060 19425 8124 19489
rect 7940 19333 8004 19397
rect 8060 19333 8124 19397
rect 7940 19241 8004 19305
rect 8060 19241 8124 19305
rect 7940 19148 8004 19212
rect 8060 19148 8124 19212
rect 10318 39528 10382 39592
rect 10446 39528 10510 39592
rect 10318 39448 10382 39512
rect 10446 39448 10510 39512
rect 10318 39368 10382 39432
rect 10446 39368 10510 39432
rect 10318 39288 10382 39352
rect 10446 39288 10510 39352
rect 10318 39208 10382 39272
rect 10446 39208 10510 39272
rect 10318 39128 10382 39192
rect 10446 39128 10510 39192
rect 10318 39048 10382 39112
rect 10446 39048 10510 39112
rect 10318 38968 10382 39032
rect 10446 38968 10510 39032
rect 10318 38888 10382 38952
rect 10446 38888 10510 38952
rect 10318 38808 10382 38872
rect 10446 38808 10510 38872
rect 10318 38728 10382 38792
rect 10446 38728 10510 38792
rect 10318 38648 10382 38712
rect 10446 38648 10510 38712
rect 10318 38568 10382 38632
rect 10446 38568 10510 38632
rect 10318 38488 10382 38552
rect 10446 38488 10510 38552
rect 10318 38408 10382 38472
rect 10446 38408 10510 38472
rect 10318 38328 10382 38392
rect 10446 38328 10510 38392
rect 10318 38247 10382 38311
rect 10446 38247 10510 38311
rect 10318 38166 10382 38230
rect 10446 38166 10510 38230
rect 10318 38085 10382 38149
rect 10446 38085 10510 38149
rect 10318 38004 10382 38068
rect 10446 38004 10510 38068
rect 10318 37923 10382 37987
rect 10446 37923 10510 37987
rect 10318 37842 10382 37906
rect 10446 37842 10510 37906
rect 10318 37761 10382 37825
rect 10446 37761 10510 37825
rect 10318 37680 10382 37744
rect 10446 37680 10510 37744
rect 10318 37599 10382 37663
rect 10446 37599 10510 37663
rect 10318 37518 10382 37582
rect 10446 37518 10510 37582
rect 10318 37437 10382 37501
rect 10446 37437 10510 37501
rect 10318 37356 10382 37420
rect 10446 37356 10510 37420
rect 10318 37275 10382 37339
rect 10446 37275 10510 37339
rect 10318 37194 10382 37258
rect 10446 37194 10510 37258
rect 10318 37113 10382 37177
rect 10446 37113 10510 37177
rect 10318 37032 10382 37096
rect 10446 37032 10510 37096
rect 10318 36951 10382 37015
rect 10446 36951 10510 37015
rect 10318 36870 10382 36934
rect 10446 36870 10510 36934
rect 10318 36789 10382 36853
rect 10446 36789 10510 36853
rect 10318 36708 10382 36772
rect 10446 36708 10510 36772
rect 10318 36627 10382 36691
rect 10446 36627 10510 36691
rect 10318 36546 10382 36610
rect 10446 36546 10510 36610
rect 10318 36465 10382 36529
rect 10446 36465 10510 36529
rect 10318 36384 10382 36448
rect 10446 36384 10510 36448
rect 10318 36303 10382 36367
rect 10446 36303 10510 36367
rect 10318 36222 10382 36286
rect 10446 36222 10510 36286
rect 10318 36141 10382 36205
rect 10446 36141 10510 36205
rect 10318 36060 10382 36124
rect 10446 36060 10510 36124
rect 10318 35979 10382 36043
rect 10446 35979 10510 36043
rect 10318 35898 10382 35962
rect 10446 35898 10510 35962
rect 10318 35817 10382 35881
rect 10446 35817 10510 35881
rect 10318 35736 10382 35800
rect 10446 35736 10510 35800
rect 10318 35655 10382 35719
rect 10446 35655 10510 35719
rect 10318 35574 10382 35638
rect 10446 35574 10510 35638
rect 10318 35493 10382 35557
rect 10446 35493 10510 35557
rect 10318 35412 10382 35476
rect 10446 35412 10510 35476
rect 10318 35331 10382 35395
rect 10446 35331 10510 35395
rect 10318 35250 10382 35314
rect 10446 35250 10510 35314
rect 10318 35169 10382 35233
rect 10446 35169 10510 35233
rect 10318 35088 10382 35152
rect 10446 35088 10510 35152
rect 10318 35007 10382 35071
rect 10446 35007 10510 35071
rect 10318 34926 10382 34990
rect 10446 34926 10510 34990
rect 10318 34845 10382 34909
rect 10446 34845 10510 34909
rect 10318 34764 10382 34828
rect 10446 34764 10510 34828
rect 9822 34155 9886 34219
rect 9950 34155 10014 34219
rect 9822 34061 9886 34125
rect 9950 34061 10014 34125
rect 9822 33966 9886 34030
rect 9950 33966 10014 34030
rect 9822 33871 9886 33935
rect 9950 33871 10014 33935
rect 9822 33776 9886 33840
rect 9950 33776 10014 33840
rect 9822 33681 9886 33745
rect 9950 33681 10014 33745
rect 8932 19609 8996 19673
rect 9052 19609 9116 19673
rect 8932 19517 8996 19581
rect 9052 19517 9116 19581
rect 8932 19425 8996 19489
rect 9052 19425 9116 19489
rect 8932 19333 8996 19397
rect 9052 19333 9116 19397
rect 8932 19241 8996 19305
rect 9052 19241 9116 19305
rect 8932 19148 8996 19212
rect 9052 19148 9116 19212
rect 11310 39528 11374 39592
rect 11438 39528 11502 39592
rect 11310 39448 11374 39512
rect 11438 39448 11502 39512
rect 11310 39368 11374 39432
rect 11438 39368 11502 39432
rect 11310 39288 11374 39352
rect 11438 39288 11502 39352
rect 11310 39208 11374 39272
rect 11438 39208 11502 39272
rect 11310 39128 11374 39192
rect 11438 39128 11502 39192
rect 11310 39048 11374 39112
rect 11438 39048 11502 39112
rect 11310 38968 11374 39032
rect 11438 38968 11502 39032
rect 11310 38888 11374 38952
rect 11438 38888 11502 38952
rect 11310 38808 11374 38872
rect 11438 38808 11502 38872
rect 11310 38728 11374 38792
rect 11438 38728 11502 38792
rect 11310 38648 11374 38712
rect 11438 38648 11502 38712
rect 11310 38568 11374 38632
rect 11438 38568 11502 38632
rect 11310 38488 11374 38552
rect 11438 38488 11502 38552
rect 11310 38408 11374 38472
rect 11438 38408 11502 38472
rect 11310 38328 11374 38392
rect 11438 38328 11502 38392
rect 11310 38247 11374 38311
rect 11438 38247 11502 38311
rect 11310 38166 11374 38230
rect 11438 38166 11502 38230
rect 11310 38085 11374 38149
rect 11438 38085 11502 38149
rect 11310 38004 11374 38068
rect 11438 38004 11502 38068
rect 11310 37923 11374 37987
rect 11438 37923 11502 37987
rect 11310 37842 11374 37906
rect 11438 37842 11502 37906
rect 11310 37761 11374 37825
rect 11438 37761 11502 37825
rect 11310 37680 11374 37744
rect 11438 37680 11502 37744
rect 11310 37599 11374 37663
rect 11438 37599 11502 37663
rect 11310 37518 11374 37582
rect 11438 37518 11502 37582
rect 11310 37437 11374 37501
rect 11438 37437 11502 37501
rect 11310 37356 11374 37420
rect 11438 37356 11502 37420
rect 11310 37275 11374 37339
rect 11438 37275 11502 37339
rect 11310 37194 11374 37258
rect 11438 37194 11502 37258
rect 11310 37113 11374 37177
rect 11438 37113 11502 37177
rect 11310 37032 11374 37096
rect 11438 37032 11502 37096
rect 11310 36951 11374 37015
rect 11438 36951 11502 37015
rect 11310 36870 11374 36934
rect 11438 36870 11502 36934
rect 11310 36789 11374 36853
rect 11438 36789 11502 36853
rect 11310 36708 11374 36772
rect 11438 36708 11502 36772
rect 11310 36627 11374 36691
rect 11438 36627 11502 36691
rect 11310 36546 11374 36610
rect 11438 36546 11502 36610
rect 11310 36465 11374 36529
rect 11438 36465 11502 36529
rect 11310 36384 11374 36448
rect 11438 36384 11502 36448
rect 11310 36303 11374 36367
rect 11438 36303 11502 36367
rect 11310 36222 11374 36286
rect 11438 36222 11502 36286
rect 11310 36141 11374 36205
rect 11438 36141 11502 36205
rect 11310 36060 11374 36124
rect 11438 36060 11502 36124
rect 11310 35979 11374 36043
rect 11438 35979 11502 36043
rect 11310 35898 11374 35962
rect 11438 35898 11502 35962
rect 11310 35817 11374 35881
rect 11438 35817 11502 35881
rect 11310 35736 11374 35800
rect 11438 35736 11502 35800
rect 11310 35655 11374 35719
rect 11438 35655 11502 35719
rect 11310 35574 11374 35638
rect 11438 35574 11502 35638
rect 11310 35493 11374 35557
rect 11438 35493 11502 35557
rect 11310 35412 11374 35476
rect 11438 35412 11502 35476
rect 11310 35331 11374 35395
rect 11438 35331 11502 35395
rect 11310 35250 11374 35314
rect 11438 35250 11502 35314
rect 11310 35169 11374 35233
rect 11438 35169 11502 35233
rect 11310 35088 11374 35152
rect 11438 35088 11502 35152
rect 11310 35007 11374 35071
rect 11438 35007 11502 35071
rect 11310 34926 11374 34990
rect 11438 34926 11502 34990
rect 11310 34845 11374 34909
rect 11438 34845 11502 34909
rect 11310 34764 11374 34828
rect 11438 34764 11502 34828
rect 10814 34155 10878 34219
rect 10942 34155 11006 34219
rect 10814 34061 10878 34125
rect 10942 34061 11006 34125
rect 10814 33966 10878 34030
rect 10942 33966 11006 34030
rect 10814 33871 10878 33935
rect 10942 33871 11006 33935
rect 10814 33776 10878 33840
rect 10942 33776 11006 33840
rect 10814 33681 10878 33745
rect 10942 33681 11006 33745
rect 12302 39528 12366 39592
rect 12430 39528 12494 39592
rect 12302 39448 12366 39512
rect 12430 39448 12494 39512
rect 12302 39368 12366 39432
rect 12430 39368 12494 39432
rect 12302 39288 12366 39352
rect 12430 39288 12494 39352
rect 12302 39208 12366 39272
rect 12430 39208 12494 39272
rect 12302 39128 12366 39192
rect 12430 39128 12494 39192
rect 12302 39048 12366 39112
rect 12430 39048 12494 39112
rect 12302 38968 12366 39032
rect 12430 38968 12494 39032
rect 12302 38888 12366 38952
rect 12430 38888 12494 38952
rect 12302 38808 12366 38872
rect 12430 38808 12494 38872
rect 12302 38728 12366 38792
rect 12430 38728 12494 38792
rect 12302 38648 12366 38712
rect 12430 38648 12494 38712
rect 12302 38568 12366 38632
rect 12430 38568 12494 38632
rect 12302 38488 12366 38552
rect 12430 38488 12494 38552
rect 12302 38408 12366 38472
rect 12430 38408 12494 38472
rect 12302 38328 12366 38392
rect 12430 38328 12494 38392
rect 12302 38247 12366 38311
rect 12430 38247 12494 38311
rect 12302 38166 12366 38230
rect 12430 38166 12494 38230
rect 12302 38085 12366 38149
rect 12430 38085 12494 38149
rect 12302 38004 12366 38068
rect 12430 38004 12494 38068
rect 12302 37923 12366 37987
rect 12430 37923 12494 37987
rect 12302 37842 12366 37906
rect 12430 37842 12494 37906
rect 12302 37761 12366 37825
rect 12430 37761 12494 37825
rect 12302 37680 12366 37744
rect 12430 37680 12494 37744
rect 12302 37599 12366 37663
rect 12430 37599 12494 37663
rect 12302 37518 12366 37582
rect 12430 37518 12494 37582
rect 12302 37437 12366 37501
rect 12430 37437 12494 37501
rect 12302 37356 12366 37420
rect 12430 37356 12494 37420
rect 12302 37275 12366 37339
rect 12430 37275 12494 37339
rect 12302 37194 12366 37258
rect 12430 37194 12494 37258
rect 12302 37113 12366 37177
rect 12430 37113 12494 37177
rect 12302 37032 12366 37096
rect 12430 37032 12494 37096
rect 12302 36951 12366 37015
rect 12430 36951 12494 37015
rect 12302 36870 12366 36934
rect 12430 36870 12494 36934
rect 12302 36789 12366 36853
rect 12430 36789 12494 36853
rect 12302 36708 12366 36772
rect 12430 36708 12494 36772
rect 12302 36627 12366 36691
rect 12430 36627 12494 36691
rect 12302 36546 12366 36610
rect 12430 36546 12494 36610
rect 12302 36465 12366 36529
rect 12430 36465 12494 36529
rect 12302 36384 12366 36448
rect 12430 36384 12494 36448
rect 12302 36303 12366 36367
rect 12430 36303 12494 36367
rect 12302 36222 12366 36286
rect 12430 36222 12494 36286
rect 12302 36141 12366 36205
rect 12430 36141 12494 36205
rect 12302 36060 12366 36124
rect 12430 36060 12494 36124
rect 12302 35979 12366 36043
rect 12430 35979 12494 36043
rect 12302 35898 12366 35962
rect 12430 35898 12494 35962
rect 12302 35817 12366 35881
rect 12430 35817 12494 35881
rect 12302 35736 12366 35800
rect 12430 35736 12494 35800
rect 12302 35655 12366 35719
rect 12430 35655 12494 35719
rect 12302 35574 12366 35638
rect 12430 35574 12494 35638
rect 12302 35493 12366 35557
rect 12430 35493 12494 35557
rect 12302 35412 12366 35476
rect 12430 35412 12494 35476
rect 12302 35331 12366 35395
rect 12430 35331 12494 35395
rect 12302 35250 12366 35314
rect 12430 35250 12494 35314
rect 12302 35169 12366 35233
rect 12430 35169 12494 35233
rect 12302 35088 12366 35152
rect 12430 35088 12494 35152
rect 12302 35007 12366 35071
rect 12430 35007 12494 35071
rect 12302 34926 12366 34990
rect 12430 34926 12494 34990
rect 12302 34845 12366 34909
rect 12430 34845 12494 34909
rect 12302 34764 12366 34828
rect 12430 34764 12494 34828
rect 11806 34155 11870 34219
rect 11934 34155 11998 34219
rect 11806 34061 11870 34125
rect 11934 34061 11998 34125
rect 11806 33966 11870 34030
rect 11934 33966 11998 34030
rect 11806 33871 11870 33935
rect 11934 33871 11998 33935
rect 11806 33776 11870 33840
rect 11934 33776 11998 33840
rect 11806 33681 11870 33745
rect 11934 33681 11998 33745
rect 13294 39528 13358 39592
rect 13422 39528 13486 39592
rect 13294 39448 13358 39512
rect 13422 39448 13486 39512
rect 13294 39368 13358 39432
rect 13422 39368 13486 39432
rect 13294 39288 13358 39352
rect 13422 39288 13486 39352
rect 13294 39208 13358 39272
rect 13422 39208 13486 39272
rect 13294 39128 13358 39192
rect 13422 39128 13486 39192
rect 13294 39048 13358 39112
rect 13422 39048 13486 39112
rect 13294 38968 13358 39032
rect 13422 38968 13486 39032
rect 13294 38888 13358 38952
rect 13422 38888 13486 38952
rect 13294 38808 13358 38872
rect 13422 38808 13486 38872
rect 13294 38728 13358 38792
rect 13422 38728 13486 38792
rect 13294 38648 13358 38712
rect 13422 38648 13486 38712
rect 13294 38568 13358 38632
rect 13422 38568 13486 38632
rect 13294 38488 13358 38552
rect 13422 38488 13486 38552
rect 13294 38408 13358 38472
rect 13422 38408 13486 38472
rect 13294 38328 13358 38392
rect 13422 38328 13486 38392
rect 13294 38247 13358 38311
rect 13422 38247 13486 38311
rect 13294 38166 13358 38230
rect 13422 38166 13486 38230
rect 13294 38085 13358 38149
rect 13422 38085 13486 38149
rect 13294 38004 13358 38068
rect 13422 38004 13486 38068
rect 13294 37923 13358 37987
rect 13422 37923 13486 37987
rect 13294 37842 13358 37906
rect 13422 37842 13486 37906
rect 13294 37761 13358 37825
rect 13422 37761 13486 37825
rect 13294 37680 13358 37744
rect 13422 37680 13486 37744
rect 13294 37599 13358 37663
rect 13422 37599 13486 37663
rect 13294 37518 13358 37582
rect 13422 37518 13486 37582
rect 13294 37437 13358 37501
rect 13422 37437 13486 37501
rect 13294 37356 13358 37420
rect 13422 37356 13486 37420
rect 13294 37275 13358 37339
rect 13422 37275 13486 37339
rect 13294 37194 13358 37258
rect 13422 37194 13486 37258
rect 13294 37113 13358 37177
rect 13422 37113 13486 37177
rect 13294 37032 13358 37096
rect 13422 37032 13486 37096
rect 13294 36951 13358 37015
rect 13422 36951 13486 37015
rect 13294 36870 13358 36934
rect 13422 36870 13486 36934
rect 13294 36789 13358 36853
rect 13422 36789 13486 36853
rect 13294 36708 13358 36772
rect 13422 36708 13486 36772
rect 13294 36627 13358 36691
rect 13422 36627 13486 36691
rect 13294 36546 13358 36610
rect 13422 36546 13486 36610
rect 13294 36465 13358 36529
rect 13422 36465 13486 36529
rect 13294 36384 13358 36448
rect 13422 36384 13486 36448
rect 13294 36303 13358 36367
rect 13422 36303 13486 36367
rect 13294 36222 13358 36286
rect 13422 36222 13486 36286
rect 13294 36141 13358 36205
rect 13422 36141 13486 36205
rect 13294 36060 13358 36124
rect 13422 36060 13486 36124
rect 13294 35979 13358 36043
rect 13422 35979 13486 36043
rect 13294 35898 13358 35962
rect 13422 35898 13486 35962
rect 13294 35817 13358 35881
rect 13422 35817 13486 35881
rect 13294 35736 13358 35800
rect 13422 35736 13486 35800
rect 13294 35655 13358 35719
rect 13422 35655 13486 35719
rect 13294 35574 13358 35638
rect 13422 35574 13486 35638
rect 13294 35493 13358 35557
rect 13422 35493 13486 35557
rect 13294 35412 13358 35476
rect 13422 35412 13486 35476
rect 13294 35331 13358 35395
rect 13422 35331 13486 35395
rect 13294 35250 13358 35314
rect 13422 35250 13486 35314
rect 13294 35169 13358 35233
rect 13422 35169 13486 35233
rect 13294 35088 13358 35152
rect 13422 35088 13486 35152
rect 13294 35007 13358 35071
rect 13422 35007 13486 35071
rect 13294 34926 13358 34990
rect 13422 34926 13486 34990
rect 13294 34845 13358 34909
rect 13422 34845 13486 34909
rect 13294 34764 13358 34828
rect 13422 34764 13486 34828
rect 12798 33890 12862 33954
rect 12926 33890 12990 33954
rect 12798 33796 12862 33860
rect 12926 33796 12990 33860
rect 12798 33701 12862 33765
rect 12926 33701 12990 33765
rect 12798 33606 12862 33670
rect 12926 33606 12990 33670
rect 12798 33511 12862 33575
rect 12926 33511 12990 33575
rect 12798 33416 12862 33480
rect 12926 33416 12990 33480
rect 14255 39528 14319 39592
rect 14343 39528 14407 39592
rect 14431 39528 14495 39592
rect 14519 39528 14583 39592
rect 14607 39528 14671 39592
rect 14255 39448 14319 39512
rect 14343 39448 14407 39512
rect 14431 39448 14495 39512
rect 14519 39448 14583 39512
rect 14607 39448 14671 39512
rect 14255 39368 14319 39432
rect 14343 39368 14407 39432
rect 14431 39368 14495 39432
rect 14519 39368 14583 39432
rect 14607 39368 14671 39432
rect 14255 39288 14319 39352
rect 14343 39288 14407 39352
rect 14431 39288 14495 39352
rect 14519 39288 14583 39352
rect 14607 39288 14671 39352
rect 14255 39208 14319 39272
rect 14343 39208 14407 39272
rect 14431 39208 14495 39272
rect 14519 39208 14583 39272
rect 14607 39208 14671 39272
rect 14255 39128 14319 39192
rect 14343 39128 14407 39192
rect 14431 39128 14495 39192
rect 14519 39128 14583 39192
rect 14607 39128 14671 39192
rect 14255 39048 14319 39112
rect 14343 39048 14407 39112
rect 14431 39048 14495 39112
rect 14519 39048 14583 39112
rect 14607 39048 14671 39112
rect 14255 38968 14319 39032
rect 14343 38968 14407 39032
rect 14431 38968 14495 39032
rect 14519 38968 14583 39032
rect 14607 38968 14671 39032
rect 14255 38888 14319 38952
rect 14343 38888 14407 38952
rect 14431 38888 14495 38952
rect 14519 38888 14583 38952
rect 14607 38888 14671 38952
rect 14255 38808 14319 38872
rect 14343 38808 14407 38872
rect 14431 38808 14495 38872
rect 14519 38808 14583 38872
rect 14607 38808 14671 38872
rect 14255 38728 14319 38792
rect 14343 38728 14407 38792
rect 14431 38728 14495 38792
rect 14519 38728 14583 38792
rect 14607 38728 14671 38792
rect 14255 38648 14319 38712
rect 14343 38648 14407 38712
rect 14431 38648 14495 38712
rect 14519 38648 14583 38712
rect 14607 38648 14671 38712
rect 14255 38568 14319 38632
rect 14343 38568 14407 38632
rect 14431 38568 14495 38632
rect 14519 38568 14583 38632
rect 14607 38568 14671 38632
rect 14255 38488 14319 38552
rect 14343 38488 14407 38552
rect 14431 38488 14495 38552
rect 14519 38488 14583 38552
rect 14607 38488 14671 38552
rect 14255 38408 14319 38472
rect 14343 38408 14407 38472
rect 14431 38408 14495 38472
rect 14519 38408 14583 38472
rect 14607 38408 14671 38472
rect 14255 38328 14319 38392
rect 14343 38328 14407 38392
rect 14431 38328 14495 38392
rect 14519 38328 14583 38392
rect 14607 38328 14671 38392
rect 14255 38247 14319 38311
rect 14343 38247 14407 38311
rect 14431 38247 14495 38311
rect 14519 38247 14583 38311
rect 14607 38247 14671 38311
rect 14255 38166 14319 38230
rect 14343 38166 14407 38230
rect 14431 38166 14495 38230
rect 14519 38166 14583 38230
rect 14607 38166 14671 38230
rect 14255 38085 14319 38149
rect 14343 38085 14407 38149
rect 14431 38085 14495 38149
rect 14519 38085 14583 38149
rect 14607 38085 14671 38149
rect 14255 38004 14319 38068
rect 14343 38004 14407 38068
rect 14431 38004 14495 38068
rect 14519 38004 14583 38068
rect 14607 38004 14671 38068
rect 14255 37923 14319 37987
rect 14343 37923 14407 37987
rect 14431 37923 14495 37987
rect 14519 37923 14583 37987
rect 14607 37923 14671 37987
rect 14255 37842 14319 37906
rect 14343 37842 14407 37906
rect 14431 37842 14495 37906
rect 14519 37842 14583 37906
rect 14607 37842 14671 37906
rect 14255 37761 14319 37825
rect 14343 37761 14407 37825
rect 14431 37761 14495 37825
rect 14519 37761 14583 37825
rect 14607 37761 14671 37825
rect 14255 37680 14319 37744
rect 14343 37680 14407 37744
rect 14431 37680 14495 37744
rect 14519 37680 14583 37744
rect 14607 37680 14671 37744
rect 14255 37599 14319 37663
rect 14343 37599 14407 37663
rect 14431 37599 14495 37663
rect 14519 37599 14583 37663
rect 14607 37599 14671 37663
rect 14255 37518 14319 37582
rect 14343 37518 14407 37582
rect 14431 37518 14495 37582
rect 14519 37518 14583 37582
rect 14607 37518 14671 37582
rect 14255 37437 14319 37501
rect 14343 37437 14407 37501
rect 14431 37437 14495 37501
rect 14519 37437 14583 37501
rect 14607 37437 14671 37501
rect 14255 37356 14319 37420
rect 14343 37356 14407 37420
rect 14431 37356 14495 37420
rect 14519 37356 14583 37420
rect 14607 37356 14671 37420
rect 14255 37275 14319 37339
rect 14343 37275 14407 37339
rect 14431 37275 14495 37339
rect 14519 37275 14583 37339
rect 14607 37275 14671 37339
rect 14255 37194 14319 37258
rect 14343 37194 14407 37258
rect 14431 37194 14495 37258
rect 14519 37194 14583 37258
rect 14607 37194 14671 37258
rect 14255 37113 14319 37177
rect 14343 37113 14407 37177
rect 14431 37113 14495 37177
rect 14519 37113 14583 37177
rect 14607 37113 14671 37177
rect 14255 37032 14319 37096
rect 14343 37032 14407 37096
rect 14431 37032 14495 37096
rect 14519 37032 14583 37096
rect 14607 37032 14671 37096
rect 14255 36951 14319 37015
rect 14343 36951 14407 37015
rect 14431 36951 14495 37015
rect 14519 36951 14583 37015
rect 14607 36951 14671 37015
rect 14255 36870 14319 36934
rect 14343 36870 14407 36934
rect 14431 36870 14495 36934
rect 14519 36870 14583 36934
rect 14607 36870 14671 36934
rect 14255 36789 14319 36853
rect 14343 36789 14407 36853
rect 14431 36789 14495 36853
rect 14519 36789 14583 36853
rect 14607 36789 14671 36853
rect 14255 36708 14319 36772
rect 14343 36708 14407 36772
rect 14431 36708 14495 36772
rect 14519 36708 14583 36772
rect 14607 36708 14671 36772
rect 14255 36627 14319 36691
rect 14343 36627 14407 36691
rect 14431 36627 14495 36691
rect 14519 36627 14583 36691
rect 14607 36627 14671 36691
rect 14255 36546 14319 36610
rect 14343 36546 14407 36610
rect 14431 36546 14495 36610
rect 14519 36546 14583 36610
rect 14607 36546 14671 36610
rect 14255 36465 14319 36529
rect 14343 36465 14407 36529
rect 14431 36465 14495 36529
rect 14519 36465 14583 36529
rect 14607 36465 14671 36529
rect 14255 36384 14319 36448
rect 14343 36384 14407 36448
rect 14431 36384 14495 36448
rect 14519 36384 14583 36448
rect 14607 36384 14671 36448
rect 14255 36303 14319 36367
rect 14343 36303 14407 36367
rect 14431 36303 14495 36367
rect 14519 36303 14583 36367
rect 14607 36303 14671 36367
rect 14255 36222 14319 36286
rect 14343 36222 14407 36286
rect 14431 36222 14495 36286
rect 14519 36222 14583 36286
rect 14607 36222 14671 36286
rect 14255 36141 14319 36205
rect 14343 36141 14407 36205
rect 14431 36141 14495 36205
rect 14519 36141 14583 36205
rect 14607 36141 14671 36205
rect 14255 36060 14319 36124
rect 14343 36060 14407 36124
rect 14431 36060 14495 36124
rect 14519 36060 14583 36124
rect 14607 36060 14671 36124
rect 14255 35979 14319 36043
rect 14343 35979 14407 36043
rect 14431 35979 14495 36043
rect 14519 35979 14583 36043
rect 14607 35979 14671 36043
rect 14255 35898 14319 35962
rect 14343 35898 14407 35962
rect 14431 35898 14495 35962
rect 14519 35898 14583 35962
rect 14607 35898 14671 35962
rect 14255 35817 14319 35881
rect 14343 35817 14407 35881
rect 14431 35817 14495 35881
rect 14519 35817 14583 35881
rect 14607 35817 14671 35881
rect 14255 35736 14319 35800
rect 14343 35736 14407 35800
rect 14431 35736 14495 35800
rect 14519 35736 14583 35800
rect 14607 35736 14671 35800
rect 14255 35655 14319 35719
rect 14343 35655 14407 35719
rect 14431 35655 14495 35719
rect 14519 35655 14583 35719
rect 14607 35655 14671 35719
rect 14255 35574 14319 35638
rect 14343 35574 14407 35638
rect 14431 35574 14495 35638
rect 14519 35574 14583 35638
rect 14607 35574 14671 35638
rect 14255 35493 14319 35557
rect 14343 35493 14407 35557
rect 14431 35493 14495 35557
rect 14519 35493 14583 35557
rect 14607 35493 14671 35557
rect 14255 35412 14319 35476
rect 14343 35412 14407 35476
rect 14431 35412 14495 35476
rect 14519 35412 14583 35476
rect 14607 35412 14671 35476
rect 14255 35331 14319 35395
rect 14343 35331 14407 35395
rect 14431 35331 14495 35395
rect 14519 35331 14583 35395
rect 14607 35331 14671 35395
rect 14255 35250 14319 35314
rect 14343 35250 14407 35314
rect 14431 35250 14495 35314
rect 14519 35250 14583 35314
rect 14607 35250 14671 35314
rect 14255 35169 14319 35233
rect 14343 35169 14407 35233
rect 14431 35169 14495 35233
rect 14519 35169 14583 35233
rect 14607 35169 14671 35233
rect 14255 35088 14319 35152
rect 14343 35088 14407 35152
rect 14431 35088 14495 35152
rect 14519 35088 14583 35152
rect 14607 35088 14671 35152
rect 14255 35007 14319 35071
rect 14343 35007 14407 35071
rect 14431 35007 14495 35071
rect 14519 35007 14583 35071
rect 14607 35007 14671 35071
rect 14255 34926 14319 34990
rect 14343 34926 14407 34990
rect 14431 34926 14495 34990
rect 14519 34926 14583 34990
rect 14607 34926 14671 34990
rect 14255 34845 14319 34909
rect 14343 34845 14407 34909
rect 14431 34845 14495 34909
rect 14519 34845 14583 34909
rect 14607 34845 14671 34909
rect 14255 34764 14319 34828
rect 14343 34764 14407 34828
rect 14431 34764 14495 34828
rect 14519 34764 14583 34828
rect 14607 34764 14671 34828
rect 13790 32919 13854 32983
rect 13892 32919 13956 32983
rect 13790 32839 13854 32903
rect 13892 32839 13956 32903
rect 13790 32759 13854 32823
rect 13892 32759 13956 32823
rect 13790 32679 13854 32743
rect 13892 32679 13956 32743
rect 13790 32599 13854 32663
rect 13892 32599 13956 32663
rect 13790 32519 13854 32583
rect 13892 32519 13956 32583
rect 13790 32439 13854 32503
rect 13892 32439 13956 32503
rect 13790 32359 13854 32423
rect 13892 32359 13956 32423
rect 13790 32279 13854 32343
rect 13892 32279 13956 32343
rect 13790 32199 13854 32263
rect 13892 32199 13956 32263
rect 13790 32119 13854 32183
rect 13892 32119 13956 32183
rect 13790 32039 13854 32103
rect 13892 32039 13956 32103
rect 13790 32018 13854 32023
rect 13790 31962 13795 32018
rect 13795 31962 13851 32018
rect 13851 31962 13854 32018
rect 13790 31959 13854 31962
rect 13892 32018 13956 32023
rect 13892 31962 13921 32018
rect 13921 31962 13956 32018
rect 13892 31959 13956 31962
rect 13790 31936 13854 31943
rect 13790 31880 13795 31936
rect 13795 31880 13851 31936
rect 13851 31880 13854 31936
rect 13790 31879 13854 31880
rect 13892 31936 13956 31943
rect 13892 31880 13921 31936
rect 13921 31880 13956 31936
rect 13892 31879 13956 31880
rect 13790 31854 13854 31863
rect 13790 31799 13795 31854
rect 13795 31799 13851 31854
rect 13851 31799 13854 31854
rect 13892 31854 13956 31863
rect 13892 31799 13921 31854
rect 13921 31799 13956 31854
rect 13790 31772 13854 31783
rect 13790 31719 13795 31772
rect 13795 31719 13851 31772
rect 13851 31719 13854 31772
rect 13892 31772 13956 31783
rect 13892 31719 13921 31772
rect 13921 31719 13956 31772
rect 13790 31690 13854 31703
rect 13790 31639 13795 31690
rect 13795 31639 13851 31690
rect 13851 31639 13854 31690
rect 13892 31690 13956 31703
rect 13892 31639 13921 31690
rect 13921 31639 13956 31690
rect 13790 31608 13854 31623
rect 13790 31559 13795 31608
rect 13795 31559 13851 31608
rect 13851 31559 13854 31608
rect 13892 31608 13956 31623
rect 13892 31559 13921 31608
rect 13921 31559 13956 31608
rect 13790 31526 13854 31543
rect 13790 31479 13795 31526
rect 13795 31479 13851 31526
rect 13851 31479 13854 31526
rect 13892 31526 13956 31543
rect 13892 31479 13921 31526
rect 13921 31479 13956 31526
rect 13790 31444 13854 31463
rect 13790 31399 13795 31444
rect 13795 31399 13851 31444
rect 13851 31399 13854 31444
rect 13892 31444 13956 31463
rect 13892 31399 13921 31444
rect 13921 31399 13956 31444
rect 13790 31362 13854 31383
rect 13790 31319 13795 31362
rect 13795 31319 13851 31362
rect 13851 31319 13854 31362
rect 13892 31362 13956 31383
rect 13892 31319 13921 31362
rect 13921 31319 13956 31362
rect 13790 31280 13854 31303
rect 13790 31239 13795 31280
rect 13795 31239 13851 31280
rect 13851 31239 13854 31280
rect 13892 31280 13956 31303
rect 13892 31239 13921 31280
rect 13921 31239 13956 31280
rect 13790 31198 13854 31223
rect 13790 31159 13795 31198
rect 13795 31159 13851 31198
rect 13851 31159 13854 31198
rect 13892 31198 13956 31223
rect 13892 31159 13921 31198
rect 13921 31159 13956 31198
rect 13790 31142 13795 31143
rect 13795 31142 13851 31143
rect 13851 31142 13854 31143
rect 13790 31116 13854 31142
rect 13790 31079 13795 31116
rect 13795 31079 13851 31116
rect 13851 31079 13854 31116
rect 13892 31142 13921 31143
rect 13921 31142 13956 31143
rect 13892 31116 13956 31142
rect 13892 31079 13921 31116
rect 13921 31079 13956 31116
rect 13790 31060 13795 31063
rect 13795 31060 13851 31063
rect 13851 31060 13854 31063
rect 13790 31034 13854 31060
rect 13790 30999 13795 31034
rect 13795 30999 13851 31034
rect 13851 30999 13854 31034
rect 13892 31060 13921 31063
rect 13921 31060 13956 31063
rect 13892 31034 13956 31060
rect 13892 30999 13921 31034
rect 13921 30999 13956 31034
rect 13790 30978 13795 30983
rect 13795 30978 13851 30983
rect 13851 30978 13854 30983
rect 13790 30952 13854 30978
rect 13790 30919 13795 30952
rect 13795 30919 13851 30952
rect 13851 30919 13854 30952
rect 13892 30978 13921 30983
rect 13921 30978 13956 30983
rect 13892 30952 13956 30978
rect 13892 30919 13921 30952
rect 13921 30919 13956 30952
rect 13790 30896 13795 30903
rect 13795 30896 13851 30903
rect 13851 30896 13854 30903
rect 13790 30870 13854 30896
rect 13790 30839 13795 30870
rect 13795 30839 13851 30870
rect 13851 30839 13854 30870
rect 13892 30896 13921 30903
rect 13921 30896 13956 30903
rect 13892 30870 13956 30896
rect 13892 30839 13921 30870
rect 13921 30839 13956 30870
rect 13790 30814 13795 30822
rect 13795 30814 13851 30822
rect 13851 30814 13854 30822
rect 13790 30788 13854 30814
rect 13790 30758 13795 30788
rect 13795 30758 13851 30788
rect 13851 30758 13854 30788
rect 13892 30814 13921 30822
rect 13921 30814 13956 30822
rect 13892 30788 13956 30814
rect 13892 30758 13921 30788
rect 13921 30758 13956 30788
rect 13790 30732 13795 30741
rect 13795 30732 13851 30741
rect 13851 30732 13854 30741
rect 13790 30706 13854 30732
rect 13790 30677 13795 30706
rect 13795 30677 13851 30706
rect 13851 30677 13854 30706
rect 13892 30732 13921 30741
rect 13921 30732 13956 30741
rect 13892 30706 13956 30732
rect 13892 30677 13921 30706
rect 13921 30677 13956 30706
rect 13790 30650 13795 30660
rect 13795 30650 13851 30660
rect 13851 30650 13854 30660
rect 13790 30624 13854 30650
rect 13790 30596 13795 30624
rect 13795 30596 13851 30624
rect 13851 30596 13854 30624
rect 13892 30650 13921 30660
rect 13921 30650 13956 30660
rect 13892 30624 13956 30650
rect 13892 30596 13921 30624
rect 13921 30596 13956 30624
rect 13790 30568 13795 30579
rect 13795 30568 13851 30579
rect 13851 30568 13854 30579
rect 13790 30542 13854 30568
rect 13790 30515 13795 30542
rect 13795 30515 13851 30542
rect 13851 30515 13854 30542
rect 13892 30568 13921 30579
rect 13921 30568 13956 30579
rect 13892 30542 13956 30568
rect 13892 30515 13921 30542
rect 13921 30515 13956 30542
rect 13790 30486 13795 30498
rect 13795 30486 13851 30498
rect 13851 30486 13854 30498
rect 13790 30460 13854 30486
rect 13790 30434 13795 30460
rect 13795 30434 13851 30460
rect 13851 30434 13854 30460
rect 13892 30486 13921 30498
rect 13921 30486 13956 30498
rect 13892 30460 13956 30486
rect 13892 30434 13921 30460
rect 13921 30434 13956 30460
rect 13790 30404 13795 30417
rect 13795 30404 13851 30417
rect 13851 30404 13854 30417
rect 13790 30378 13854 30404
rect 13790 30353 13795 30378
rect 13795 30353 13851 30378
rect 13851 30353 13854 30378
rect 13892 30404 13921 30417
rect 13921 30404 13956 30417
rect 13892 30378 13956 30404
rect 13892 30353 13921 30378
rect 13921 30353 13956 30378
rect 13790 30322 13795 30336
rect 13795 30322 13851 30336
rect 13851 30322 13854 30336
rect 13790 30296 13854 30322
rect 13790 30272 13795 30296
rect 13795 30272 13851 30296
rect 13851 30272 13854 30296
rect 13892 30322 13921 30336
rect 13921 30322 13956 30336
rect 13892 30296 13956 30322
rect 13892 30272 13921 30296
rect 13921 30272 13956 30296
rect 13790 30240 13795 30255
rect 13795 30240 13851 30255
rect 13851 30240 13854 30255
rect 13790 30214 13854 30240
rect 13790 30191 13795 30214
rect 13795 30191 13851 30214
rect 13851 30191 13854 30214
rect 13892 30240 13921 30255
rect 13921 30240 13956 30255
rect 13892 30214 13956 30240
rect 13892 30191 13921 30214
rect 13921 30191 13956 30214
rect 13790 30158 13795 30174
rect 13795 30158 13851 30174
rect 13851 30158 13854 30174
rect 13790 30132 13854 30158
rect 13790 30110 13795 30132
rect 13795 30110 13851 30132
rect 13851 30110 13854 30132
rect 13892 30158 13921 30174
rect 13921 30158 13956 30174
rect 13892 30132 13956 30158
rect 13892 30110 13921 30132
rect 13921 30110 13956 30132
rect 13790 30076 13795 30093
rect 13795 30076 13851 30093
rect 13851 30076 13854 30093
rect 13790 30050 13854 30076
rect 13790 30029 13795 30050
rect 13795 30029 13851 30050
rect 13851 30029 13854 30050
rect 13892 30076 13921 30093
rect 13921 30076 13956 30093
rect 13892 30050 13956 30076
rect 13892 30029 13921 30050
rect 13921 30029 13956 30050
rect 13790 29994 13795 30012
rect 13795 29994 13851 30012
rect 13851 29994 13854 30012
rect 13790 29968 13854 29994
rect 13790 29948 13795 29968
rect 13795 29948 13851 29968
rect 13851 29948 13854 29968
rect 13892 29994 13921 30012
rect 13921 29994 13956 30012
rect 13892 29968 13956 29994
rect 13892 29948 13921 29968
rect 13921 29948 13956 29968
rect 13790 29912 13795 29931
rect 13795 29912 13851 29931
rect 13851 29912 13854 29931
rect 13790 29886 13854 29912
rect 13790 29867 13795 29886
rect 13795 29867 13851 29886
rect 13851 29867 13854 29886
rect 13892 29912 13921 29931
rect 13921 29912 13956 29931
rect 13892 29886 13956 29912
rect 13892 29867 13921 29886
rect 13921 29867 13956 29886
rect 13790 29830 13795 29850
rect 13795 29830 13851 29850
rect 13851 29830 13854 29850
rect 13790 29804 13854 29830
rect 13790 29786 13795 29804
rect 13795 29786 13851 29804
rect 13851 29786 13854 29804
rect 13892 29830 13921 29850
rect 13921 29830 13956 29850
rect 13892 29804 13956 29830
rect 13892 29786 13921 29804
rect 13921 29786 13956 29804
rect 13790 29748 13795 29769
rect 13795 29748 13851 29769
rect 13851 29748 13854 29769
rect 13790 29722 13854 29748
rect 13790 29705 13795 29722
rect 13795 29705 13851 29722
rect 13851 29705 13854 29722
rect 13892 29748 13921 29769
rect 13921 29748 13956 29769
rect 13892 29722 13956 29748
rect 13892 29705 13921 29722
rect 13921 29705 13956 29722
rect 13790 29666 13795 29688
rect 13795 29666 13851 29688
rect 13851 29666 13854 29688
rect 13790 29640 13854 29666
rect 13790 29624 13795 29640
rect 13795 29624 13851 29640
rect 13851 29624 13854 29640
rect 13892 29666 13921 29688
rect 13921 29666 13956 29688
rect 13892 29640 13956 29666
rect 13892 29624 13921 29640
rect 13921 29624 13956 29640
rect 13790 29584 13795 29607
rect 13795 29584 13851 29607
rect 13851 29584 13854 29607
rect 13790 29558 13854 29584
rect 13790 29543 13795 29558
rect 13795 29543 13851 29558
rect 13851 29543 13854 29558
rect 13892 29584 13921 29607
rect 13921 29584 13956 29607
rect 13892 29558 13956 29584
rect 13892 29543 13921 29558
rect 13921 29543 13956 29558
rect 13790 29502 13795 29526
rect 13795 29502 13851 29526
rect 13851 29502 13854 29526
rect 13790 29476 13854 29502
rect 13790 29462 13795 29476
rect 13795 29462 13851 29476
rect 13851 29462 13854 29476
rect 13892 29502 13921 29526
rect 13921 29502 13956 29526
rect 13892 29476 13956 29502
rect 13892 29462 13921 29476
rect 13921 29462 13956 29476
rect 13790 29420 13795 29445
rect 13795 29420 13851 29445
rect 13851 29420 13854 29445
rect 13790 29381 13854 29420
rect 13892 29420 13921 29445
rect 13921 29420 13956 29445
rect 13892 29381 13956 29420
rect 13790 29300 13854 29364
rect 13892 29300 13956 29364
rect 13790 29219 13854 29283
rect 13892 29219 13956 29283
rect 13790 29138 13854 29202
rect 13892 29138 13956 29202
rect 13790 29057 13854 29121
rect 13892 29057 13956 29121
rect 13790 28976 13854 29040
rect 13892 28976 13956 29040
rect 13790 28895 13854 28959
rect 13892 28895 13956 28959
rect 13790 28814 13854 28878
rect 13892 28814 13956 28878
rect 13790 28733 13854 28797
rect 13892 28733 13956 28797
rect 13790 28652 13854 28716
rect 13892 28652 13956 28716
rect 13790 28571 13854 28635
rect 13892 28571 13956 28635
rect 13790 28490 13854 28554
rect 13892 28490 13956 28554
rect 13790 28409 13854 28473
rect 13892 28409 13956 28473
rect 13790 28328 13854 28392
rect 13892 28328 13956 28392
rect 13790 28247 13854 28311
rect 13892 28247 13956 28311
rect 13790 28166 13854 28230
rect 13892 28166 13956 28230
rect 13790 28085 13854 28149
rect 13892 28085 13956 28149
rect 13790 28004 13854 28068
rect 13892 28004 13956 28068
rect 13790 27923 13854 27987
rect 13892 27923 13956 27987
rect 13790 27842 13854 27906
rect 13892 27842 13956 27906
rect 13790 27761 13854 27825
rect 13892 27761 13956 27825
rect 13790 27680 13854 27744
rect 13892 27680 13956 27744
rect 13790 27599 13854 27663
rect 13892 27599 13956 27663
rect 13790 27518 13854 27582
rect 13892 27518 13956 27582
rect 13790 27437 13854 27501
rect 13892 27437 13956 27501
rect 13790 27356 13854 27420
rect 13892 27356 13956 27420
rect 13790 27275 13854 27339
rect 13892 27275 13956 27339
rect 13974 27283 14038 27347
rect 13790 27194 13854 27258
rect 13892 27194 13956 27258
rect 13974 27198 14038 27262
rect 13790 27113 13854 27177
rect 13892 27113 13956 27177
rect 13974 27112 14038 27176
rect 8432 18528 8496 18592
rect 8560 18528 8624 18592
rect 8432 18448 8496 18512
rect 8560 18448 8624 18512
rect 8432 18368 8496 18432
rect 8560 18368 8624 18432
rect 8432 18288 8496 18352
rect 8560 18288 8624 18352
rect 8432 18208 8496 18272
rect 8560 18208 8624 18272
rect 8432 18128 8496 18192
rect 8560 18128 8624 18192
rect 8432 18048 8496 18112
rect 8560 18048 8624 18112
rect 8432 17968 8496 18032
rect 8560 17968 8624 18032
rect 8432 17888 8496 17952
rect 8560 17888 8624 17952
rect 8432 17808 8496 17872
rect 8560 17808 8624 17872
rect 8432 17728 8496 17792
rect 8560 17728 8624 17792
rect 8432 17648 8496 17712
rect 8560 17648 8624 17712
rect 8432 17568 8496 17632
rect 8560 17568 8624 17632
rect 8432 17488 8496 17552
rect 8560 17488 8624 17552
rect 8432 17408 8496 17472
rect 8560 17408 8624 17472
rect 8432 17328 8496 17392
rect 8560 17328 8624 17392
rect 8432 17248 8496 17312
rect 8560 17248 8624 17312
rect 8432 17168 8496 17232
rect 8560 17168 8624 17232
rect 8432 17088 8496 17152
rect 8560 17088 8624 17152
rect 8432 17008 8496 17072
rect 8560 17008 8624 17072
rect 8432 16928 8496 16992
rect 8560 16928 8624 16992
rect 8432 16848 8496 16912
rect 8560 16848 8624 16912
rect 8432 16768 8496 16832
rect 8560 16768 8624 16832
rect 8432 16688 8496 16752
rect 8560 16688 8624 16752
rect 8432 16608 8496 16672
rect 8560 16608 8624 16672
rect 8432 16528 8496 16592
rect 8560 16528 8624 16592
rect 8432 16448 8496 16512
rect 8560 16448 8624 16512
rect 8432 16368 8496 16432
rect 8560 16368 8624 16432
rect 8432 16287 8496 16351
rect 8560 16287 8624 16351
rect 8432 16206 8496 16270
rect 8560 16206 8624 16270
rect 8432 16125 8496 16189
rect 8560 16125 8624 16189
rect 8432 16044 8496 16108
rect 8560 16044 8624 16108
rect 8432 15963 8496 16027
rect 8560 15963 8624 16027
rect 8432 15882 8496 15946
rect 8560 15882 8624 15946
rect 8432 15801 8496 15865
rect 8560 15801 8624 15865
rect 8432 15720 8496 15784
rect 8560 15720 8624 15784
rect 8432 15639 8496 15703
rect 8560 15639 8624 15703
rect 8432 15558 8496 15622
rect 8560 15558 8624 15622
rect 8432 15477 8496 15541
rect 8560 15477 8624 15541
rect 8432 15396 8496 15460
rect 8560 15396 8624 15460
rect 8432 15315 8496 15379
rect 8560 15315 8624 15379
rect 8432 15234 8496 15298
rect 8560 15234 8624 15298
rect 8432 15153 8496 15217
rect 8560 15153 8624 15217
rect 8432 15072 8496 15136
rect 8560 15072 8624 15136
rect 8432 14991 8496 15055
rect 8560 14991 8624 15055
rect 8432 14910 8496 14974
rect 8560 14910 8624 14974
rect 8432 14829 8496 14893
rect 8560 14829 8624 14893
rect 8432 14748 8496 14812
rect 8560 14748 8624 14812
rect 8432 14667 8496 14731
rect 8560 14667 8624 14731
rect 8432 14586 8496 14650
rect 8560 14586 8624 14650
rect 8432 14505 8496 14569
rect 8560 14505 8624 14569
rect 8432 14424 8496 14488
rect 8560 14424 8624 14488
rect 8432 14343 8496 14407
rect 8560 14343 8624 14407
rect 8432 14262 8496 14326
rect 8560 14262 8624 14326
rect 8432 14181 8496 14245
rect 8560 14181 8624 14245
rect 8432 14100 8496 14164
rect 8560 14100 8624 14164
rect 8432 14019 8496 14083
rect 8560 14019 8624 14083
rect 8432 13938 8496 14002
rect 8560 13938 8624 14002
rect 8432 13857 8496 13921
rect 8560 13857 8624 13921
rect 8432 13776 8496 13840
rect 8560 13776 8624 13840
rect 8432 13695 8496 13759
rect 8560 13695 8624 13759
rect 8432 13614 8496 13678
rect 8560 13614 8624 13678
rect 9924 19609 9988 19673
rect 10044 19609 10108 19673
rect 9924 19517 9988 19581
rect 10044 19517 10108 19581
rect 9924 19425 9988 19489
rect 10044 19425 10108 19489
rect 9924 19333 9988 19397
rect 10044 19333 10108 19397
rect 9924 19241 9988 19305
rect 10044 19241 10108 19305
rect 9924 19148 9988 19212
rect 10044 19148 10108 19212
rect 9424 18528 9488 18592
rect 9552 18528 9616 18592
rect 9424 18448 9488 18512
rect 9552 18448 9616 18512
rect 9424 18368 9488 18432
rect 9552 18368 9616 18432
rect 9424 18288 9488 18352
rect 9552 18288 9616 18352
rect 9424 18208 9488 18272
rect 9552 18208 9616 18272
rect 9424 18128 9488 18192
rect 9552 18128 9616 18192
rect 9424 18048 9488 18112
rect 9552 18048 9616 18112
rect 9424 17968 9488 18032
rect 9552 17968 9616 18032
rect 9424 17888 9488 17952
rect 9552 17888 9616 17952
rect 9424 17808 9488 17872
rect 9552 17808 9616 17872
rect 9424 17728 9488 17792
rect 9552 17728 9616 17792
rect 9424 17648 9488 17712
rect 9552 17648 9616 17712
rect 9424 17568 9488 17632
rect 9552 17568 9616 17632
rect 9424 17488 9488 17552
rect 9552 17488 9616 17552
rect 9424 17408 9488 17472
rect 9552 17408 9616 17472
rect 9424 17328 9488 17392
rect 9552 17328 9616 17392
rect 9424 17248 9488 17312
rect 9552 17248 9616 17312
rect 9424 17168 9488 17232
rect 9552 17168 9616 17232
rect 9424 17088 9488 17152
rect 9552 17088 9616 17152
rect 9424 17008 9488 17072
rect 9552 17008 9616 17072
rect 9424 16928 9488 16992
rect 9552 16928 9616 16992
rect 9424 16848 9488 16912
rect 9552 16848 9616 16912
rect 9424 16768 9488 16832
rect 9552 16768 9616 16832
rect 9424 16688 9488 16752
rect 9552 16688 9616 16752
rect 9424 16608 9488 16672
rect 9552 16608 9616 16672
rect 9424 16528 9488 16592
rect 9552 16528 9616 16592
rect 9424 16448 9488 16512
rect 9552 16448 9616 16512
rect 9424 16368 9488 16432
rect 9552 16368 9616 16432
rect 9424 16287 9488 16351
rect 9552 16287 9616 16351
rect 9424 16206 9488 16270
rect 9552 16206 9616 16270
rect 9424 16125 9488 16189
rect 9552 16125 9616 16189
rect 9424 16044 9488 16108
rect 9552 16044 9616 16108
rect 9424 15963 9488 16027
rect 9552 15963 9616 16027
rect 9424 15882 9488 15946
rect 9552 15882 9616 15946
rect 9424 15801 9488 15865
rect 9552 15801 9616 15865
rect 9424 15720 9488 15784
rect 9552 15720 9616 15784
rect 9424 15639 9488 15703
rect 9552 15639 9616 15703
rect 9424 15558 9488 15622
rect 9552 15558 9616 15622
rect 9424 15477 9488 15541
rect 9552 15477 9616 15541
rect 9424 15396 9488 15460
rect 9552 15396 9616 15460
rect 9424 15315 9488 15379
rect 9552 15315 9616 15379
rect 9424 15234 9488 15298
rect 9552 15234 9616 15298
rect 9424 15153 9488 15217
rect 9552 15153 9616 15217
rect 9424 15072 9488 15136
rect 9552 15072 9616 15136
rect 9424 14991 9488 15055
rect 9552 14991 9616 15055
rect 9424 14910 9488 14974
rect 9552 14910 9616 14974
rect 9424 14829 9488 14893
rect 9552 14829 9616 14893
rect 9424 14748 9488 14812
rect 9552 14748 9616 14812
rect 9424 14667 9488 14731
rect 9552 14667 9616 14731
rect 9424 14586 9488 14650
rect 9552 14586 9616 14650
rect 9424 14505 9488 14569
rect 9552 14505 9616 14569
rect 9424 14424 9488 14488
rect 9552 14424 9616 14488
rect 9424 14343 9488 14407
rect 9552 14343 9616 14407
rect 9424 14262 9488 14326
rect 9552 14262 9616 14326
rect 9424 14181 9488 14245
rect 9552 14181 9616 14245
rect 9424 14100 9488 14164
rect 9552 14100 9616 14164
rect 9424 14019 9488 14083
rect 9552 14019 9616 14083
rect 9424 13938 9488 14002
rect 9552 13938 9616 14002
rect 9424 13857 9488 13921
rect 9552 13857 9616 13921
rect 9424 13776 9488 13840
rect 9552 13776 9616 13840
rect 9424 13695 9488 13759
rect 9552 13695 9616 13759
rect 9424 13614 9488 13678
rect 9552 13614 9616 13678
rect 10916 19609 10980 19673
rect 11036 19609 11100 19673
rect 10916 19517 10980 19581
rect 11036 19517 11100 19581
rect 10916 19425 10980 19489
rect 11036 19425 11100 19489
rect 10916 19333 10980 19397
rect 11036 19333 11100 19397
rect 10916 19241 10980 19305
rect 11036 19241 11100 19305
rect 10916 19148 10980 19212
rect 11036 19148 11100 19212
rect 10416 18528 10480 18592
rect 10544 18528 10608 18592
rect 10416 18448 10480 18512
rect 10544 18448 10608 18512
rect 10416 18368 10480 18432
rect 10544 18368 10608 18432
rect 10416 18288 10480 18352
rect 10544 18288 10608 18352
rect 10416 18208 10480 18272
rect 10544 18208 10608 18272
rect 10416 18128 10480 18192
rect 10544 18128 10608 18192
rect 10416 18048 10480 18112
rect 10544 18048 10608 18112
rect 10416 17968 10480 18032
rect 10544 17968 10608 18032
rect 10416 17888 10480 17952
rect 10544 17888 10608 17952
rect 10416 17808 10480 17872
rect 10544 17808 10608 17872
rect 10416 17728 10480 17792
rect 10544 17728 10608 17792
rect 10416 17648 10480 17712
rect 10544 17648 10608 17712
rect 10416 17568 10480 17632
rect 10544 17568 10608 17632
rect 10416 17488 10480 17552
rect 10544 17488 10608 17552
rect 10416 17408 10480 17472
rect 10544 17408 10608 17472
rect 10416 17328 10480 17392
rect 10544 17328 10608 17392
rect 10416 17248 10480 17312
rect 10544 17248 10608 17312
rect 10416 17168 10480 17232
rect 10544 17168 10608 17232
rect 10416 17088 10480 17152
rect 10544 17088 10608 17152
rect 10416 17008 10480 17072
rect 10544 17008 10608 17072
rect 10416 16928 10480 16992
rect 10544 16928 10608 16992
rect 10416 16848 10480 16912
rect 10544 16848 10608 16912
rect 10416 16768 10480 16832
rect 10544 16768 10608 16832
rect 10416 16688 10480 16752
rect 10544 16688 10608 16752
rect 10416 16608 10480 16672
rect 10544 16608 10608 16672
rect 10416 16528 10480 16592
rect 10544 16528 10608 16592
rect 10416 16448 10480 16512
rect 10544 16448 10608 16512
rect 10416 16368 10480 16432
rect 10544 16368 10608 16432
rect 10416 16287 10480 16351
rect 10544 16287 10608 16351
rect 10416 16206 10480 16270
rect 10544 16206 10608 16270
rect 10416 16125 10480 16189
rect 10544 16125 10608 16189
rect 10416 16044 10480 16108
rect 10544 16044 10608 16108
rect 10416 15963 10480 16027
rect 10544 15963 10608 16027
rect 10416 15882 10480 15946
rect 10544 15882 10608 15946
rect 10416 15801 10480 15865
rect 10544 15801 10608 15865
rect 10416 15720 10480 15784
rect 10544 15720 10608 15784
rect 10416 15639 10480 15703
rect 10544 15639 10608 15703
rect 10416 15558 10480 15622
rect 10544 15558 10608 15622
rect 10416 15477 10480 15541
rect 10544 15477 10608 15541
rect 10416 15396 10480 15460
rect 10544 15396 10608 15460
rect 10416 15315 10480 15379
rect 10544 15315 10608 15379
rect 10416 15234 10480 15298
rect 10544 15234 10608 15298
rect 10416 15153 10480 15217
rect 10544 15153 10608 15217
rect 10416 15072 10480 15136
rect 10544 15072 10608 15136
rect 10416 14991 10480 15055
rect 10544 14991 10608 15055
rect 10416 14910 10480 14974
rect 10544 14910 10608 14974
rect 10416 14829 10480 14893
rect 10544 14829 10608 14893
rect 10416 14748 10480 14812
rect 10544 14748 10608 14812
rect 10416 14667 10480 14731
rect 10544 14667 10608 14731
rect 10416 14586 10480 14650
rect 10544 14586 10608 14650
rect 10416 14505 10480 14569
rect 10544 14505 10608 14569
rect 10416 14424 10480 14488
rect 10544 14424 10608 14488
rect 10416 14343 10480 14407
rect 10544 14343 10608 14407
rect 10416 14262 10480 14326
rect 10544 14262 10608 14326
rect 10416 14181 10480 14245
rect 10544 14181 10608 14245
rect 10416 14100 10480 14164
rect 10544 14100 10608 14164
rect 10416 14019 10480 14083
rect 10544 14019 10608 14083
rect 10416 13938 10480 14002
rect 10544 13938 10608 14002
rect 10416 13857 10480 13921
rect 10544 13857 10608 13921
rect 10416 13776 10480 13840
rect 10544 13776 10608 13840
rect 10416 13695 10480 13759
rect 10544 13695 10608 13759
rect 10416 13614 10480 13678
rect 10544 13614 10608 13678
rect 11908 19609 11972 19673
rect 12028 19609 12092 19673
rect 11908 19517 11972 19581
rect 12028 19517 12092 19581
rect 11908 19425 11972 19489
rect 12028 19425 12092 19489
rect 11908 19333 11972 19397
rect 12028 19333 12092 19397
rect 11908 19241 11972 19305
rect 12028 19241 12092 19305
rect 11908 19148 11972 19212
rect 12028 19148 12092 19212
rect 11408 18528 11472 18592
rect 11536 18528 11600 18592
rect 11408 18448 11472 18512
rect 11536 18448 11600 18512
rect 11408 18368 11472 18432
rect 11536 18368 11600 18432
rect 11408 18288 11472 18352
rect 11536 18288 11600 18352
rect 11408 18208 11472 18272
rect 11536 18208 11600 18272
rect 11408 18128 11472 18192
rect 11536 18128 11600 18192
rect 11408 18048 11472 18112
rect 11536 18048 11600 18112
rect 11408 17968 11472 18032
rect 11536 17968 11600 18032
rect 11408 17888 11472 17952
rect 11536 17888 11600 17952
rect 11408 17808 11472 17872
rect 11536 17808 11600 17872
rect 11408 17728 11472 17792
rect 11536 17728 11600 17792
rect 11408 17648 11472 17712
rect 11536 17648 11600 17712
rect 11408 17568 11472 17632
rect 11536 17568 11600 17632
rect 11408 17488 11472 17552
rect 11536 17488 11600 17552
rect 11408 17408 11472 17472
rect 11536 17408 11600 17472
rect 11408 17328 11472 17392
rect 11536 17328 11600 17392
rect 11408 17248 11472 17312
rect 11536 17248 11600 17312
rect 11408 17168 11472 17232
rect 11536 17168 11600 17232
rect 11408 17088 11472 17152
rect 11536 17088 11600 17152
rect 11408 17008 11472 17072
rect 11536 17008 11600 17072
rect 11408 16928 11472 16992
rect 11536 16928 11600 16992
rect 11408 16848 11472 16912
rect 11536 16848 11600 16912
rect 11408 16768 11472 16832
rect 11536 16768 11600 16832
rect 11408 16688 11472 16752
rect 11536 16688 11600 16752
rect 11408 16608 11472 16672
rect 11536 16608 11600 16672
rect 11408 16528 11472 16592
rect 11536 16528 11600 16592
rect 11408 16448 11472 16512
rect 11536 16448 11600 16512
rect 11408 16368 11472 16432
rect 11536 16368 11600 16432
rect 11408 16287 11472 16351
rect 11536 16287 11600 16351
rect 11408 16206 11472 16270
rect 11536 16206 11600 16270
rect 11408 16125 11472 16189
rect 11536 16125 11600 16189
rect 11408 16044 11472 16108
rect 11536 16044 11600 16108
rect 11408 15963 11472 16027
rect 11536 15963 11600 16027
rect 11408 15882 11472 15946
rect 11536 15882 11600 15946
rect 11408 15801 11472 15865
rect 11536 15801 11600 15865
rect 11408 15720 11472 15784
rect 11536 15720 11600 15784
rect 11408 15639 11472 15703
rect 11536 15639 11600 15703
rect 11408 15558 11472 15622
rect 11536 15558 11600 15622
rect 11408 15477 11472 15541
rect 11536 15477 11600 15541
rect 11408 15396 11472 15460
rect 11536 15396 11600 15460
rect 11408 15315 11472 15379
rect 11536 15315 11600 15379
rect 11408 15234 11472 15298
rect 11536 15234 11600 15298
rect 11408 15153 11472 15217
rect 11536 15153 11600 15217
rect 11408 15072 11472 15136
rect 11536 15072 11600 15136
rect 11408 14991 11472 15055
rect 11536 14991 11600 15055
rect 11408 14910 11472 14974
rect 11536 14910 11600 14974
rect 11408 14829 11472 14893
rect 11536 14829 11600 14893
rect 11408 14748 11472 14812
rect 11536 14748 11600 14812
rect 11408 14667 11472 14731
rect 11536 14667 11600 14731
rect 11408 14586 11472 14650
rect 11536 14586 11600 14650
rect 11408 14505 11472 14569
rect 11536 14505 11600 14569
rect 11408 14424 11472 14488
rect 11536 14424 11600 14488
rect 11408 14343 11472 14407
rect 11536 14343 11600 14407
rect 11408 14262 11472 14326
rect 11536 14262 11600 14326
rect 11408 14181 11472 14245
rect 11536 14181 11600 14245
rect 11408 14100 11472 14164
rect 11536 14100 11600 14164
rect 11408 14019 11472 14083
rect 11536 14019 11600 14083
rect 11408 13938 11472 14002
rect 11536 13938 11600 14002
rect 11408 13857 11472 13921
rect 11536 13857 11600 13921
rect 11408 13776 11472 13840
rect 11536 13776 11600 13840
rect 11408 13695 11472 13759
rect 11536 13695 11600 13759
rect 11408 13614 11472 13678
rect 11536 13614 11600 13678
rect 13649 27010 13713 27074
rect 13757 27010 13821 27074
rect 13865 27010 13929 27074
rect 13973 27010 14037 27074
rect 13649 26900 13713 26964
rect 13757 26900 13821 26964
rect 13865 26900 13929 26964
rect 13973 26900 14037 26964
rect 13649 26828 13651 26854
rect 13651 26828 13707 26854
rect 13707 26828 13713 26854
rect 13757 26828 13789 26854
rect 13789 26828 13815 26854
rect 13815 26828 13821 26854
rect 13865 26828 13871 26854
rect 13871 26828 13897 26854
rect 13897 26828 13929 26854
rect 13973 26828 13979 26854
rect 13979 26828 14035 26854
rect 14035 26828 14037 26854
rect 13649 26800 13713 26828
rect 13757 26800 13821 26828
rect 13865 26800 13929 26828
rect 13973 26800 14037 26828
rect 13649 26790 13651 26800
rect 13651 26790 13707 26800
rect 13707 26790 13713 26800
rect 13757 26790 13789 26800
rect 13789 26790 13815 26800
rect 13815 26790 13821 26800
rect 13865 26790 13871 26800
rect 13871 26790 13897 26800
rect 13897 26790 13929 26800
rect 13973 26790 13979 26800
rect 13979 26790 14035 26800
rect 14035 26790 14037 26800
rect 13649 26716 13713 26744
rect 13757 26716 13821 26744
rect 13865 26716 13929 26744
rect 13973 26716 14037 26744
rect 13649 26680 13651 26716
rect 13651 26680 13707 26716
rect 13707 26680 13713 26716
rect 13757 26680 13789 26716
rect 13789 26680 13815 26716
rect 13815 26680 13821 26716
rect 13865 26680 13871 26716
rect 13871 26680 13897 26716
rect 13897 26680 13929 26716
rect 13973 26680 13979 26716
rect 13979 26680 14035 26716
rect 14035 26680 14037 26716
rect 13649 26632 13713 26634
rect 13757 26632 13821 26634
rect 13865 26632 13929 26634
rect 13973 26632 14037 26634
rect 13649 26576 13651 26632
rect 13651 26576 13707 26632
rect 13707 26576 13713 26632
rect 13757 26576 13789 26632
rect 13789 26576 13815 26632
rect 13815 26576 13821 26632
rect 13865 26576 13871 26632
rect 13871 26576 13897 26632
rect 13897 26576 13929 26632
rect 13973 26576 13979 26632
rect 13979 26576 14035 26632
rect 14035 26576 14037 26632
rect 13649 26570 13713 26576
rect 13757 26570 13821 26576
rect 13865 26570 13929 26576
rect 13973 26570 14037 26576
rect 13649 26492 13651 26524
rect 13651 26492 13707 26524
rect 13707 26492 13713 26524
rect 13757 26492 13789 26524
rect 13789 26492 13815 26524
rect 13815 26492 13821 26524
rect 13865 26492 13871 26524
rect 13871 26492 13897 26524
rect 13897 26492 13929 26524
rect 13973 26492 13979 26524
rect 13979 26492 14035 26524
rect 14035 26492 14037 26524
rect 13649 26460 13713 26492
rect 13757 26460 13821 26492
rect 13865 26460 13929 26492
rect 13973 26460 14037 26492
rect 13649 26349 13713 26413
rect 13757 26349 13821 26413
rect 13865 26349 13929 26413
rect 13973 26349 14037 26413
rect 13843 26250 13907 26314
rect 13951 26250 14015 26314
rect 13843 26149 13907 26213
rect 13951 26149 14015 26213
rect 13843 26048 13907 26112
rect 13951 26048 14015 26112
rect 13843 25946 13907 26010
rect 13951 25946 14015 26010
rect 13843 25844 13907 25908
rect 13951 25844 14015 25908
rect 13843 25742 13907 25806
rect 13951 25742 14015 25806
rect 13843 25640 13907 25704
rect 13951 25640 14015 25704
rect 13843 25538 13907 25602
rect 13951 25538 14015 25602
rect 13843 25436 13907 25500
rect 13951 25436 14015 25500
rect 13843 25334 13907 25398
rect 13951 25334 14015 25398
rect 13843 25232 13907 25296
rect 13951 25232 14015 25296
rect 13843 25130 13907 25194
rect 13951 25130 14015 25194
rect 13843 25028 13907 25092
rect 13951 25028 14015 25092
rect 13843 24926 13907 24990
rect 13951 24926 14015 24990
rect 13843 24824 13907 24888
rect 13951 24824 14015 24888
rect 13843 24722 13907 24786
rect 13951 24722 14015 24786
rect 13843 24620 13907 24684
rect 13951 24620 14015 24684
rect 13843 24518 13907 24582
rect 13951 24518 14015 24582
rect 13843 24416 13907 24480
rect 13951 24416 14015 24480
rect 13843 24314 13907 24378
rect 13951 24314 14015 24378
rect 13843 24212 13907 24276
rect 13951 24212 14015 24276
rect 13843 24110 13907 24174
rect 13951 24110 14015 24174
rect 13843 24008 13907 24072
rect 13951 24008 14015 24072
rect 13843 23906 13907 23970
rect 13951 23906 14015 23970
rect 13843 23804 13907 23868
rect 13951 23804 14015 23868
rect 12900 19990 12964 20054
rect 13020 19990 13084 20054
rect 12900 19898 12964 19962
rect 13020 19898 13084 19962
rect 12900 19806 12964 19870
rect 13020 19806 13084 19870
rect 12900 19714 12964 19778
rect 13020 19714 13084 19778
rect 12900 19622 12964 19686
rect 13020 19622 13084 19686
rect 12900 19529 12964 19593
rect 13020 19529 13084 19593
rect 12400 18528 12464 18592
rect 12528 18528 12592 18592
rect 12400 18448 12464 18512
rect 12528 18448 12592 18512
rect 12400 18368 12464 18432
rect 12528 18368 12592 18432
rect 12400 18288 12464 18352
rect 12528 18288 12592 18352
rect 12400 18208 12464 18272
rect 12528 18208 12592 18272
rect 12400 18128 12464 18192
rect 12528 18128 12592 18192
rect 12400 18048 12464 18112
rect 12528 18048 12592 18112
rect 12400 17968 12464 18032
rect 12528 17968 12592 18032
rect 12400 17888 12464 17952
rect 12528 17888 12592 17952
rect 12400 17808 12464 17872
rect 12528 17808 12592 17872
rect 12400 17728 12464 17792
rect 12528 17728 12592 17792
rect 12400 17648 12464 17712
rect 12528 17648 12592 17712
rect 12400 17568 12464 17632
rect 12528 17568 12592 17632
rect 12400 17488 12464 17552
rect 12528 17488 12592 17552
rect 12400 17408 12464 17472
rect 12528 17408 12592 17472
rect 12400 17328 12464 17392
rect 12528 17328 12592 17392
rect 12400 17248 12464 17312
rect 12528 17248 12592 17312
rect 12400 17168 12464 17232
rect 12528 17168 12592 17232
rect 12400 17088 12464 17152
rect 12528 17088 12592 17152
rect 12400 17008 12464 17072
rect 12528 17008 12592 17072
rect 12400 16928 12464 16992
rect 12528 16928 12592 16992
rect 12400 16848 12464 16912
rect 12528 16848 12592 16912
rect 12400 16768 12464 16832
rect 12528 16768 12592 16832
rect 12400 16688 12464 16752
rect 12528 16688 12592 16752
rect 12400 16608 12464 16672
rect 12528 16608 12592 16672
rect 12400 16528 12464 16592
rect 12528 16528 12592 16592
rect 12400 16448 12464 16512
rect 12528 16448 12592 16512
rect 12400 16368 12464 16432
rect 12528 16368 12592 16432
rect 12400 16287 12464 16351
rect 12528 16287 12592 16351
rect 12400 16206 12464 16270
rect 12528 16206 12592 16270
rect 12400 16125 12464 16189
rect 12528 16125 12592 16189
rect 12400 16044 12464 16108
rect 12528 16044 12592 16108
rect 12400 15963 12464 16027
rect 12528 15963 12592 16027
rect 12400 15882 12464 15946
rect 12528 15882 12592 15946
rect 12400 15801 12464 15865
rect 12528 15801 12592 15865
rect 12400 15720 12464 15784
rect 12528 15720 12592 15784
rect 12400 15639 12464 15703
rect 12528 15639 12592 15703
rect 12400 15558 12464 15622
rect 12528 15558 12592 15622
rect 12400 15477 12464 15541
rect 12528 15477 12592 15541
rect 12400 15396 12464 15460
rect 12528 15396 12592 15460
rect 12400 15315 12464 15379
rect 12528 15315 12592 15379
rect 12400 15234 12464 15298
rect 12528 15234 12592 15298
rect 12400 15153 12464 15217
rect 12528 15153 12592 15217
rect 12400 15072 12464 15136
rect 12528 15072 12592 15136
rect 12400 14991 12464 15055
rect 12528 14991 12592 15055
rect 12400 14910 12464 14974
rect 12528 14910 12592 14974
rect 12400 14829 12464 14893
rect 12528 14829 12592 14893
rect 12400 14748 12464 14812
rect 12528 14748 12592 14812
rect 12400 14667 12464 14731
rect 12528 14667 12592 14731
rect 12400 14586 12464 14650
rect 12528 14586 12592 14650
rect 12400 14505 12464 14569
rect 12528 14505 12592 14569
rect 12400 14424 12464 14488
rect 12528 14424 12592 14488
rect 12400 14343 12464 14407
rect 12528 14343 12592 14407
rect 12400 14262 12464 14326
rect 12528 14262 12592 14326
rect 12400 14181 12464 14245
rect 12528 14181 12592 14245
rect 12400 14100 12464 14164
rect 12528 14100 12592 14164
rect 12400 14019 12464 14083
rect 12528 14019 12592 14083
rect 12400 13938 12464 14002
rect 12528 13938 12592 14002
rect 12400 13857 12464 13921
rect 12528 13857 12592 13921
rect 12400 13776 12464 13840
rect 12528 13776 12592 13840
rect 12400 13695 12464 13759
rect 12528 13695 12592 13759
rect 12400 13614 12464 13678
rect 12528 13614 12592 13678
rect 13843 23702 13907 23766
rect 13951 23702 14015 23766
rect 13843 23630 13894 23664
rect 13894 23630 13907 23664
rect 13843 23606 13907 23630
rect 13843 23600 13894 23606
rect 13894 23600 13907 23606
rect 13951 23630 13956 23664
rect 13956 23630 14012 23664
rect 14012 23630 14015 23664
rect 13951 23606 14015 23630
rect 13951 23600 13956 23606
rect 13956 23600 14012 23606
rect 14012 23600 14015 23606
rect 13843 23550 13894 23562
rect 13894 23550 13907 23562
rect 13843 23526 13907 23550
rect 13843 23498 13894 23526
rect 13894 23498 13907 23526
rect 13951 23550 13956 23562
rect 13956 23550 14012 23562
rect 14012 23550 14015 23562
rect 13951 23526 14015 23550
rect 13951 23498 13956 23526
rect 13956 23498 14012 23526
rect 14012 23498 14015 23526
rect 13843 23446 13907 23460
rect 13843 23396 13894 23446
rect 13894 23396 13907 23446
rect 13951 23446 14015 23460
rect 13951 23396 13956 23446
rect 13956 23396 14012 23446
rect 14012 23396 14015 23446
rect 13843 23310 13894 23358
rect 13894 23310 13907 23358
rect 13843 23294 13907 23310
rect 13951 23310 13956 23358
rect 13956 23310 14012 23358
rect 14012 23310 14015 23358
rect 13951 23294 14015 23310
rect 13843 23230 13894 23256
rect 13894 23230 13907 23256
rect 13843 23206 13907 23230
rect 13843 23192 13894 23206
rect 13894 23192 13907 23206
rect 13951 23230 13956 23256
rect 13956 23230 14012 23256
rect 14012 23230 14015 23256
rect 13951 23206 14015 23230
rect 13951 23192 13956 23206
rect 13956 23192 14012 23206
rect 14012 23192 14015 23206
rect 13843 23150 13894 23154
rect 13894 23150 13907 23154
rect 13843 23126 13907 23150
rect 13843 23090 13894 23126
rect 13894 23090 13907 23126
rect 13951 23150 13956 23154
rect 13956 23150 14012 23154
rect 14012 23150 14015 23154
rect 13951 23126 14015 23150
rect 13951 23090 13956 23126
rect 13956 23090 14012 23126
rect 14012 23090 14015 23126
rect 13843 23046 13907 23052
rect 13843 22990 13894 23046
rect 13894 22990 13907 23046
rect 13843 22988 13907 22990
rect 13951 23046 14015 23052
rect 13951 22990 13956 23046
rect 13956 22990 14012 23046
rect 14012 22990 14015 23046
rect 13951 22988 14015 22990
rect 13843 22910 13894 22950
rect 13894 22910 13907 22950
rect 13843 22886 13907 22910
rect 13951 22910 13956 22950
rect 13956 22910 14012 22950
rect 14012 22910 14015 22950
rect 13951 22886 14015 22910
rect 13843 22830 13894 22848
rect 13894 22830 13907 22848
rect 13843 22806 13907 22830
rect 13843 22784 13894 22806
rect 13894 22784 13907 22806
rect 13951 22830 13956 22848
rect 13956 22830 14012 22848
rect 14012 22830 14015 22848
rect 13951 22806 14015 22830
rect 13951 22784 13956 22806
rect 13956 22784 14012 22806
rect 14012 22784 14015 22806
rect 13843 22726 13907 22746
rect 13843 22682 13894 22726
rect 13894 22682 13907 22726
rect 13951 22726 14015 22746
rect 13951 22682 13956 22726
rect 13956 22682 14012 22726
rect 14012 22682 14015 22726
rect 13843 22590 13894 22644
rect 13894 22590 13907 22644
rect 13843 22580 13907 22590
rect 13951 22590 13956 22644
rect 13956 22590 14012 22644
rect 14012 22590 14015 22644
rect 13951 22580 14015 22590
rect 13843 22510 13894 22542
rect 13894 22510 13907 22542
rect 13843 22486 13907 22510
rect 13843 22478 13894 22486
rect 13894 22478 13907 22486
rect 13951 22510 13956 22542
rect 13956 22510 14012 22542
rect 14012 22510 14015 22542
rect 13951 22486 14015 22510
rect 13951 22478 13956 22486
rect 13956 22478 14012 22486
rect 14012 22478 14015 22486
rect 13843 22430 13894 22440
rect 13894 22430 13907 22440
rect 13843 22406 13907 22430
rect 13843 22376 13894 22406
rect 13894 22376 13907 22406
rect 13951 22430 13956 22440
rect 13956 22430 14012 22440
rect 14012 22430 14015 22440
rect 13951 22406 14015 22430
rect 13951 22376 13956 22406
rect 13956 22376 14012 22406
rect 14012 22376 14015 22406
rect 13843 22326 13907 22338
rect 13843 22274 13894 22326
rect 13894 22274 13907 22326
rect 13951 22326 14015 22338
rect 13951 22274 13956 22326
rect 13956 22274 14012 22326
rect 14012 22274 14015 22326
rect 13843 22189 13894 22236
rect 13894 22189 13907 22236
rect 13843 22172 13907 22189
rect 13951 22189 13956 22236
rect 13956 22189 14012 22236
rect 14012 22189 14015 22236
rect 13951 22172 14015 22189
rect 13843 22108 13894 22134
rect 13894 22108 13907 22134
rect 13843 22083 13907 22108
rect 13843 22070 13894 22083
rect 13894 22070 13907 22083
rect 13951 22108 13956 22134
rect 13956 22108 14012 22134
rect 14012 22108 14015 22134
rect 13951 22083 14015 22108
rect 13951 22070 13956 22083
rect 13956 22070 14012 22083
rect 14012 22070 14015 22083
rect 13843 22027 13894 22032
rect 13894 22027 13907 22032
rect 13843 22002 13907 22027
rect 13843 21968 13894 22002
rect 13894 21968 13907 22002
rect 13951 22027 13956 22032
rect 13956 22027 14012 22032
rect 14012 22027 14015 22032
rect 13951 22002 14015 22027
rect 13951 21968 13956 22002
rect 13956 21968 14012 22002
rect 14012 21968 14015 22002
rect 13843 21921 13907 21930
rect 13843 21866 13894 21921
rect 13894 21866 13907 21921
rect 13951 21921 14015 21930
rect 13951 21866 13956 21921
rect 13956 21866 14012 21921
rect 14012 21866 14015 21921
rect 13843 21784 13894 21828
rect 13894 21784 13907 21828
rect 13843 21764 13907 21784
rect 13951 21784 13956 21828
rect 13956 21784 14012 21828
rect 14012 21784 14015 21828
rect 13951 21764 14015 21784
rect 13843 21703 13894 21726
rect 13894 21703 13907 21726
rect 13843 21678 13907 21703
rect 13843 21662 13894 21678
rect 13894 21662 13907 21678
rect 13951 21703 13956 21726
rect 13956 21703 14012 21726
rect 14012 21703 14015 21726
rect 13951 21678 14015 21703
rect 13951 21662 13956 21678
rect 13956 21662 14012 21678
rect 14012 21662 14015 21678
rect 13843 21622 13894 21624
rect 13894 21622 13907 21624
rect 13843 21597 13907 21622
rect 13843 21560 13894 21597
rect 13894 21560 13907 21597
rect 13951 21622 13956 21624
rect 13956 21622 14012 21624
rect 14012 21622 14015 21624
rect 13951 21597 14015 21622
rect 13951 21560 13956 21597
rect 13956 21560 14012 21597
rect 14012 21560 14015 21597
rect 13392 18528 13456 18592
rect 13520 18528 13584 18592
rect 13392 18448 13456 18512
rect 13520 18448 13584 18512
rect 13392 18368 13456 18432
rect 13520 18368 13584 18432
rect 13392 18288 13456 18352
rect 13520 18288 13584 18352
rect 13392 18208 13456 18272
rect 13520 18208 13584 18272
rect 13392 18128 13456 18192
rect 13520 18128 13584 18192
rect 13392 18048 13456 18112
rect 13520 18048 13584 18112
rect 13392 17968 13456 18032
rect 13520 17968 13584 18032
rect 13392 17888 13456 17952
rect 13520 17888 13584 17952
rect 13392 17808 13456 17872
rect 13520 17808 13584 17872
rect 13392 17728 13456 17792
rect 13520 17728 13584 17792
rect 13392 17648 13456 17712
rect 13520 17648 13584 17712
rect 13392 17568 13456 17632
rect 13520 17568 13584 17632
rect 13392 17488 13456 17552
rect 13520 17488 13584 17552
rect 13392 17408 13456 17472
rect 13520 17408 13584 17472
rect 13392 17328 13456 17392
rect 13520 17328 13584 17392
rect 13392 17248 13456 17312
rect 13520 17248 13584 17312
rect 13392 17168 13456 17232
rect 13520 17168 13584 17232
rect 13392 17088 13456 17152
rect 13520 17088 13584 17152
rect 13392 17008 13456 17072
rect 13520 17008 13584 17072
rect 13392 16928 13456 16992
rect 13520 16928 13584 16992
rect 13392 16848 13456 16912
rect 13520 16848 13584 16912
rect 13392 16768 13456 16832
rect 13520 16768 13584 16832
rect 13392 16688 13456 16752
rect 13520 16688 13584 16752
rect 13392 16608 13456 16672
rect 13520 16608 13584 16672
rect 13392 16528 13456 16592
rect 13520 16528 13584 16592
rect 13392 16448 13456 16512
rect 13520 16448 13584 16512
rect 13392 16368 13456 16432
rect 13520 16368 13584 16432
rect 13392 16287 13456 16351
rect 13520 16287 13584 16351
rect 13392 16206 13456 16270
rect 13520 16206 13584 16270
rect 13392 16125 13456 16189
rect 13520 16125 13584 16189
rect 13392 16044 13456 16108
rect 13520 16044 13584 16108
rect 13392 15963 13456 16027
rect 13520 15963 13584 16027
rect 13392 15882 13456 15946
rect 13520 15882 13584 15946
rect 13392 15801 13456 15865
rect 13520 15801 13584 15865
rect 13392 15720 13456 15784
rect 13520 15720 13584 15784
rect 13392 15639 13456 15703
rect 13520 15639 13584 15703
rect 13392 15558 13456 15622
rect 13520 15558 13584 15622
rect 13392 15477 13456 15541
rect 13520 15477 13584 15541
rect 13392 15396 13456 15460
rect 13520 15396 13584 15460
rect 13392 15315 13456 15379
rect 13520 15315 13584 15379
rect 13392 15234 13456 15298
rect 13520 15234 13584 15298
rect 13392 15153 13456 15217
rect 13520 15153 13584 15217
rect 13392 15072 13456 15136
rect 13520 15072 13584 15136
rect 13392 14991 13456 15055
rect 13520 14991 13584 15055
rect 13392 14910 13456 14974
rect 13520 14910 13584 14974
rect 13392 14829 13456 14893
rect 13520 14829 13584 14893
rect 13392 14748 13456 14812
rect 13520 14748 13584 14812
rect 13392 14667 13456 14731
rect 13520 14667 13584 14731
rect 13392 14586 13456 14650
rect 13520 14586 13584 14650
rect 13392 14505 13456 14569
rect 13520 14505 13584 14569
rect 13392 14424 13456 14488
rect 13520 14424 13584 14488
rect 13392 14343 13456 14407
rect 13520 14343 13584 14407
rect 13392 14262 13456 14326
rect 13520 14262 13584 14326
rect 13392 14181 13456 14245
rect 13520 14181 13584 14245
rect 13392 14100 13456 14164
rect 13520 14100 13584 14164
rect 13392 14019 13456 14083
rect 13520 14019 13584 14083
rect 13392 13938 13456 14002
rect 13520 13938 13584 14002
rect 13392 13857 13456 13921
rect 13520 13857 13584 13921
rect 13392 13776 13456 13840
rect 13520 13776 13584 13840
rect 13392 13695 13456 13759
rect 13520 13695 13584 13759
rect 13392 13614 13456 13678
rect 13520 13614 13584 13678
rect 13777 18526 13841 18590
rect 13863 18526 13927 18590
rect 13949 18526 14013 18590
rect 14035 18526 14099 18590
rect 14121 18526 14185 18590
rect 14207 18526 14271 18590
rect 14293 18526 14357 18590
rect 14379 18526 14443 18590
rect 14465 18526 14529 18590
rect 13777 18446 13841 18510
rect 13863 18446 13927 18510
rect 13949 18446 14013 18510
rect 14035 18446 14099 18510
rect 14121 18446 14185 18510
rect 14207 18446 14271 18510
rect 14293 18446 14357 18510
rect 14379 18446 14443 18510
rect 14465 18446 14529 18510
rect 13777 18366 13841 18430
rect 13863 18366 13927 18430
rect 13949 18366 14013 18430
rect 14035 18366 14099 18430
rect 14121 18366 14185 18430
rect 14207 18366 14271 18430
rect 14293 18366 14357 18430
rect 14379 18366 14443 18430
rect 14465 18366 14529 18430
rect 13777 18286 13841 18350
rect 13863 18286 13927 18350
rect 13949 18286 14013 18350
rect 14035 18286 14099 18350
rect 14121 18286 14185 18350
rect 14207 18286 14271 18350
rect 14293 18286 14357 18350
rect 14379 18286 14443 18350
rect 14465 18286 14529 18350
rect 13777 18206 13841 18270
rect 13863 18206 13927 18270
rect 13949 18206 14013 18270
rect 14035 18206 14099 18270
rect 14121 18206 14185 18270
rect 14207 18206 14271 18270
rect 14293 18206 14357 18270
rect 14379 18206 14443 18270
rect 14465 18206 14529 18270
rect 13777 18126 13841 18190
rect 13863 18126 13927 18190
rect 13949 18126 14013 18190
rect 14035 18126 14099 18190
rect 14121 18126 14185 18190
rect 14207 18126 14271 18190
rect 14293 18126 14357 18190
rect 14379 18126 14443 18190
rect 14465 18126 14529 18190
rect 13777 18046 13841 18110
rect 13863 18046 13927 18110
rect 13949 18046 14013 18110
rect 14035 18046 14099 18110
rect 14121 18046 14185 18110
rect 14207 18046 14271 18110
rect 14293 18046 14357 18110
rect 14379 18046 14443 18110
rect 14465 18046 14529 18110
rect 13777 17966 13841 18030
rect 13863 17966 13927 18030
rect 13949 17966 14013 18030
rect 14035 17966 14099 18030
rect 14121 17966 14185 18030
rect 14207 17966 14271 18030
rect 14293 17966 14357 18030
rect 14379 17966 14443 18030
rect 14465 17966 14529 18030
rect 13777 17886 13841 17950
rect 13863 17886 13927 17950
rect 13949 17886 14013 17950
rect 14035 17886 14099 17950
rect 14121 17886 14185 17950
rect 14207 17886 14271 17950
rect 14293 17886 14357 17950
rect 14379 17886 14443 17950
rect 14465 17886 14529 17950
rect 13777 17806 13841 17870
rect 13863 17806 13927 17870
rect 13949 17806 14013 17870
rect 14035 17806 14099 17870
rect 14121 17806 14185 17870
rect 14207 17806 14271 17870
rect 14293 17806 14357 17870
rect 14379 17806 14443 17870
rect 14465 17806 14529 17870
rect 13777 17726 13841 17790
rect 13863 17726 13927 17790
rect 13949 17726 14013 17790
rect 14035 17726 14099 17790
rect 14121 17726 14185 17790
rect 14207 17726 14271 17790
rect 14293 17726 14357 17790
rect 14379 17726 14443 17790
rect 14465 17726 14529 17790
rect 13777 17646 13841 17710
rect 13863 17646 13927 17710
rect 13949 17646 14013 17710
rect 14035 17646 14099 17710
rect 14121 17646 14185 17710
rect 14207 17646 14271 17710
rect 14293 17646 14357 17710
rect 14379 17646 14443 17710
rect 14465 17646 14529 17710
rect 13777 17566 13841 17630
rect 13863 17566 13927 17630
rect 13949 17566 14013 17630
rect 14035 17566 14099 17630
rect 14121 17566 14185 17630
rect 14207 17566 14271 17630
rect 14293 17566 14357 17630
rect 14379 17566 14443 17630
rect 14465 17566 14529 17630
rect 13777 17486 13841 17550
rect 13863 17486 13927 17550
rect 13949 17486 14013 17550
rect 14035 17486 14099 17550
rect 14121 17486 14185 17550
rect 14207 17486 14271 17550
rect 14293 17486 14357 17550
rect 14379 17486 14443 17550
rect 14465 17486 14529 17550
rect 13777 17406 13841 17470
rect 13863 17406 13927 17470
rect 13949 17406 14013 17470
rect 14035 17406 14099 17470
rect 14121 17406 14185 17470
rect 14207 17406 14271 17470
rect 14293 17406 14357 17470
rect 14379 17406 14443 17470
rect 14465 17406 14529 17470
rect 13777 17326 13841 17390
rect 13863 17326 13927 17390
rect 13949 17326 14013 17390
rect 14035 17326 14099 17390
rect 14121 17326 14185 17390
rect 14207 17326 14271 17390
rect 14293 17326 14357 17390
rect 14379 17326 14443 17390
rect 14465 17326 14529 17390
rect 13777 17246 13841 17310
rect 13863 17246 13927 17310
rect 13949 17246 14013 17310
rect 14035 17246 14099 17310
rect 14121 17246 14185 17310
rect 14207 17246 14271 17310
rect 14293 17246 14357 17310
rect 14379 17246 14443 17310
rect 14465 17246 14529 17310
rect 13777 17166 13841 17230
rect 13863 17166 13927 17230
rect 13949 17166 14013 17230
rect 14035 17166 14099 17230
rect 14121 17166 14185 17230
rect 14207 17166 14271 17230
rect 14293 17166 14357 17230
rect 14379 17166 14443 17230
rect 14465 17166 14529 17230
rect 13777 17086 13841 17150
rect 13863 17086 13927 17150
rect 13949 17086 14013 17150
rect 14035 17086 14099 17150
rect 14121 17086 14185 17150
rect 14207 17086 14271 17150
rect 14293 17086 14357 17150
rect 14379 17086 14443 17150
rect 14465 17086 14529 17150
rect 13777 17006 13841 17070
rect 13863 17006 13927 17070
rect 13949 17006 14013 17070
rect 14035 17006 14099 17070
rect 14121 17006 14185 17070
rect 14207 17006 14271 17070
rect 14293 17006 14357 17070
rect 14379 17006 14443 17070
rect 14465 17006 14529 17070
rect 13777 16926 13841 16990
rect 13863 16926 13927 16990
rect 13949 16926 14013 16990
rect 14035 16926 14099 16990
rect 14121 16926 14185 16990
rect 14207 16926 14271 16990
rect 14293 16926 14357 16990
rect 14379 16926 14443 16990
rect 14465 16926 14529 16990
rect 13777 16846 13841 16910
rect 13863 16846 13927 16910
rect 13949 16846 14013 16910
rect 14035 16846 14099 16910
rect 14121 16846 14185 16910
rect 14207 16846 14271 16910
rect 14293 16846 14357 16910
rect 14379 16846 14443 16910
rect 14465 16846 14529 16910
rect 13777 16766 13841 16830
rect 13863 16766 13927 16830
rect 13949 16766 14013 16830
rect 14035 16766 14099 16830
rect 14121 16766 14185 16830
rect 14207 16766 14271 16830
rect 14293 16766 14357 16830
rect 14379 16766 14443 16830
rect 14465 16766 14529 16830
rect 13777 16686 13841 16750
rect 13863 16686 13927 16750
rect 13949 16686 14013 16750
rect 14035 16686 14099 16750
rect 14121 16686 14185 16750
rect 14207 16686 14271 16750
rect 14293 16686 14357 16750
rect 14379 16686 14443 16750
rect 14465 16686 14529 16750
rect 13777 16606 13841 16670
rect 13863 16606 13927 16670
rect 13949 16606 14013 16670
rect 14035 16606 14099 16670
rect 14121 16606 14185 16670
rect 14207 16606 14271 16670
rect 14293 16606 14357 16670
rect 14379 16606 14443 16670
rect 14465 16606 14529 16670
rect 13777 16526 13841 16590
rect 13863 16526 13927 16590
rect 13949 16526 14013 16590
rect 14035 16526 14099 16590
rect 14121 16526 14185 16590
rect 14207 16526 14271 16590
rect 14293 16526 14357 16590
rect 14379 16526 14443 16590
rect 14465 16526 14529 16590
rect 13777 16446 13841 16510
rect 13863 16446 13927 16510
rect 13949 16446 14013 16510
rect 14035 16446 14099 16510
rect 14121 16446 14185 16510
rect 14207 16446 14271 16510
rect 14293 16446 14357 16510
rect 14379 16446 14443 16510
rect 14465 16446 14529 16510
rect 13777 16366 13841 16430
rect 13863 16366 13927 16430
rect 13949 16366 14013 16430
rect 14035 16366 14099 16430
rect 14121 16366 14185 16430
rect 14207 16366 14271 16430
rect 14293 16366 14357 16430
rect 14379 16366 14443 16430
rect 14465 16366 14529 16430
rect 13777 16286 13841 16350
rect 13863 16286 13927 16350
rect 13949 16286 14013 16350
rect 14035 16286 14099 16350
rect 14121 16286 14185 16350
rect 14207 16286 14271 16350
rect 14293 16286 14357 16350
rect 14379 16286 14443 16350
rect 14465 16286 14529 16350
rect 13777 16206 13841 16270
rect 13863 16206 13927 16270
rect 13949 16206 14013 16270
rect 14035 16206 14099 16270
rect 14121 16206 14185 16270
rect 14207 16206 14271 16270
rect 14293 16206 14357 16270
rect 14379 16206 14443 16270
rect 14465 16206 14529 16270
rect 13777 16126 13841 16190
rect 13863 16126 13927 16190
rect 13949 16126 14013 16190
rect 14035 16126 14099 16190
rect 14121 16126 14185 16190
rect 14207 16126 14271 16190
rect 14293 16126 14357 16190
rect 14379 16126 14443 16190
rect 14465 16126 14529 16190
rect 13777 16046 13841 16110
rect 13863 16046 13927 16110
rect 13949 16046 14013 16110
rect 14035 16046 14099 16110
rect 14121 16046 14185 16110
rect 14207 16046 14271 16110
rect 14293 16046 14357 16110
rect 14379 16046 14443 16110
rect 14465 16046 14529 16110
rect 13777 15966 13841 16030
rect 13863 15966 13927 16030
rect 13949 15966 14013 16030
rect 14035 15966 14099 16030
rect 14121 15966 14185 16030
rect 14207 15966 14271 16030
rect 14293 15966 14357 16030
rect 14379 15966 14443 16030
rect 14465 15966 14529 16030
rect 13777 15886 13841 15950
rect 13863 15886 13927 15950
rect 13949 15886 14013 15950
rect 14035 15886 14099 15950
rect 14121 15886 14185 15950
rect 14207 15886 14271 15950
rect 14293 15886 14357 15950
rect 14379 15886 14443 15950
rect 14465 15886 14529 15950
rect 13777 15806 13841 15870
rect 13863 15806 13927 15870
rect 13949 15806 14013 15870
rect 14035 15806 14099 15870
rect 14121 15806 14185 15870
rect 14207 15806 14271 15870
rect 14293 15806 14357 15870
rect 14379 15806 14443 15870
rect 14465 15806 14529 15870
rect 13777 15726 13841 15790
rect 13863 15726 13927 15790
rect 13949 15726 14013 15790
rect 14035 15726 14099 15790
rect 14121 15726 14185 15790
rect 14207 15726 14271 15790
rect 14293 15726 14357 15790
rect 14379 15726 14443 15790
rect 14465 15726 14529 15790
rect 13777 15646 13841 15710
rect 13863 15646 13927 15710
rect 13949 15646 14013 15710
rect 14035 15646 14099 15710
rect 14121 15646 14185 15710
rect 14207 15646 14271 15710
rect 14293 15646 14357 15710
rect 14379 15646 14443 15710
rect 14465 15646 14529 15710
rect 13777 15566 13841 15630
rect 13863 15566 13927 15630
rect 13949 15566 14013 15630
rect 14035 15566 14099 15630
rect 14121 15566 14185 15630
rect 14207 15566 14271 15630
rect 14293 15566 14357 15630
rect 14379 15566 14443 15630
rect 14465 15566 14529 15630
rect 13777 15486 13841 15550
rect 13863 15486 13927 15550
rect 13949 15486 14013 15550
rect 14035 15486 14099 15550
rect 14121 15486 14185 15550
rect 14207 15486 14271 15550
rect 14293 15486 14357 15550
rect 14379 15486 14443 15550
rect 14465 15486 14529 15550
rect 13777 15406 13841 15470
rect 13863 15406 13927 15470
rect 13949 15406 14013 15470
rect 14035 15406 14099 15470
rect 14121 15406 14185 15470
rect 14207 15406 14271 15470
rect 14293 15406 14357 15470
rect 14379 15406 14443 15470
rect 14465 15406 14529 15470
rect 13777 15326 13841 15390
rect 13863 15326 13927 15390
rect 13949 15326 14013 15390
rect 14035 15326 14099 15390
rect 14121 15326 14185 15390
rect 14207 15326 14271 15390
rect 14293 15326 14357 15390
rect 14379 15326 14443 15390
rect 14465 15326 14529 15390
rect 13777 15246 13841 15310
rect 13863 15246 13927 15310
rect 13949 15246 14013 15310
rect 14035 15246 14099 15310
rect 14121 15246 14185 15310
rect 14207 15246 14271 15310
rect 14293 15246 14357 15310
rect 14379 15246 14443 15310
rect 14465 15246 14529 15310
rect 13777 15166 13841 15230
rect 13863 15166 13927 15230
rect 13949 15166 14013 15230
rect 14035 15166 14099 15230
rect 14121 15166 14185 15230
rect 14207 15166 14271 15230
rect 14293 15166 14357 15230
rect 14379 15166 14443 15230
rect 14465 15166 14529 15230
rect 13777 15085 13841 15149
rect 13863 15085 13927 15149
rect 13949 15085 14013 15149
rect 14035 15085 14099 15149
rect 14121 15085 14185 15149
rect 14207 15085 14271 15149
rect 14293 15085 14357 15149
rect 14379 15085 14443 15149
rect 14465 15085 14529 15149
rect 13777 15004 13841 15068
rect 13863 15004 13927 15068
rect 13949 15004 14013 15068
rect 14035 15004 14099 15068
rect 14121 15004 14185 15068
rect 14207 15004 14271 15068
rect 14293 15004 14357 15068
rect 14379 15004 14443 15068
rect 14465 15004 14529 15068
rect 13777 14923 13841 14987
rect 13863 14923 13927 14987
rect 13949 14923 14013 14987
rect 14035 14923 14099 14987
rect 14121 14923 14185 14987
rect 14207 14923 14271 14987
rect 14293 14923 14357 14987
rect 14379 14923 14443 14987
rect 14465 14923 14529 14987
rect 13777 14842 13841 14906
rect 13863 14842 13927 14906
rect 13949 14842 14013 14906
rect 14035 14842 14099 14906
rect 14121 14842 14185 14906
rect 14207 14842 14271 14906
rect 14293 14842 14357 14906
rect 14379 14842 14443 14906
rect 14465 14842 14529 14906
rect 13777 14761 13841 14825
rect 13863 14761 13927 14825
rect 13949 14761 14013 14825
rect 14035 14761 14099 14825
rect 14121 14761 14185 14825
rect 14207 14761 14271 14825
rect 14293 14761 14357 14825
rect 14379 14761 14443 14825
rect 14465 14761 14529 14825
rect 13777 14680 13841 14744
rect 13863 14680 13927 14744
rect 13949 14680 14013 14744
rect 14035 14680 14099 14744
rect 14121 14680 14185 14744
rect 14207 14680 14271 14744
rect 14293 14680 14357 14744
rect 14379 14680 14443 14744
rect 14465 14680 14529 14744
rect 13777 14599 13841 14663
rect 13863 14599 13927 14663
rect 13949 14599 14013 14663
rect 14035 14599 14099 14663
rect 14121 14599 14185 14663
rect 14207 14599 14271 14663
rect 14293 14599 14357 14663
rect 14379 14599 14443 14663
rect 14465 14599 14529 14663
rect 13777 14518 13841 14582
rect 13863 14518 13927 14582
rect 13949 14518 14013 14582
rect 14035 14518 14099 14582
rect 14121 14518 14185 14582
rect 14207 14518 14271 14582
rect 14293 14518 14357 14582
rect 14379 14518 14443 14582
rect 14465 14518 14529 14582
rect 13777 14437 13841 14501
rect 13863 14437 13927 14501
rect 13949 14437 14013 14501
rect 14035 14437 14099 14501
rect 14121 14437 14185 14501
rect 14207 14437 14271 14501
rect 14293 14437 14357 14501
rect 14379 14437 14443 14501
rect 14465 14437 14529 14501
rect 13777 14356 13841 14420
rect 13863 14356 13927 14420
rect 13949 14356 14013 14420
rect 14035 14356 14099 14420
rect 14121 14356 14185 14420
rect 14207 14356 14271 14420
rect 14293 14356 14357 14420
rect 14379 14356 14443 14420
rect 14465 14356 14529 14420
rect 13777 14275 13841 14339
rect 13863 14275 13927 14339
rect 13949 14275 14013 14339
rect 14035 14275 14099 14339
rect 14121 14275 14185 14339
rect 14207 14275 14271 14339
rect 14293 14275 14357 14339
rect 14379 14275 14443 14339
rect 14465 14275 14529 14339
rect 13777 14194 13841 14258
rect 13863 14194 13927 14258
rect 13949 14194 14013 14258
rect 14035 14194 14099 14258
rect 14121 14194 14185 14258
rect 14207 14194 14271 14258
rect 14293 14194 14357 14258
rect 14379 14194 14443 14258
rect 14465 14194 14529 14258
rect 13777 14113 13841 14177
rect 13863 14113 13927 14177
rect 13949 14113 14013 14177
rect 14035 14113 14099 14177
rect 14121 14113 14185 14177
rect 14207 14113 14271 14177
rect 14293 14113 14357 14177
rect 14379 14113 14443 14177
rect 14465 14113 14529 14177
rect 13777 14032 13841 14096
rect 13863 14032 13927 14096
rect 13949 14032 14013 14096
rect 14035 14032 14099 14096
rect 14121 14032 14185 14096
rect 14207 14032 14271 14096
rect 14293 14032 14357 14096
rect 14379 14032 14443 14096
rect 14465 14032 14529 14096
rect 13777 13951 13841 14015
rect 13863 13951 13927 14015
rect 13949 13951 14013 14015
rect 14035 13951 14099 14015
rect 14121 13951 14185 14015
rect 14207 13951 14271 14015
rect 14293 13951 14357 14015
rect 14379 13951 14443 14015
rect 14465 13951 14529 14015
rect 13777 13870 13841 13934
rect 13863 13870 13927 13934
rect 13949 13870 14013 13934
rect 14035 13870 14099 13934
rect 14121 13870 14185 13934
rect 14207 13870 14271 13934
rect 14293 13870 14357 13934
rect 14379 13870 14443 13934
rect 14465 13870 14529 13934
rect 13777 13789 13841 13853
rect 13863 13789 13927 13853
rect 13949 13789 14013 13853
rect 14035 13789 14099 13853
rect 14121 13789 14185 13853
rect 14207 13789 14271 13853
rect 14293 13789 14357 13853
rect 14379 13789 14443 13853
rect 14465 13789 14529 13853
rect 13777 13708 13841 13772
rect 13863 13708 13927 13772
rect 13949 13708 14013 13772
rect 14035 13708 14099 13772
rect 14121 13708 14185 13772
rect 14207 13708 14271 13772
rect 14293 13708 14357 13772
rect 14379 13708 14443 13772
rect 14465 13708 14529 13772
rect 13777 13627 13841 13691
rect 13863 13627 13927 13691
rect 13949 13627 14013 13691
rect 14035 13627 14099 13691
rect 14121 13627 14185 13691
rect 14207 13627 14271 13691
rect 14293 13627 14357 13691
rect 14379 13627 14443 13691
rect 14465 13627 14529 13691
rect 204 8785 259 8835
rect 259 8785 268 8835
rect 204 8771 268 8785
rect 287 8785 343 8835
rect 343 8785 351 8835
rect 287 8771 351 8785
rect 370 8785 371 8835
rect 371 8785 427 8835
rect 427 8785 434 8835
rect 370 8771 434 8785
rect 453 8785 454 8835
rect 454 8785 510 8835
rect 510 8785 517 8835
rect 453 8771 517 8785
rect 536 8785 537 8835
rect 537 8785 593 8835
rect 593 8785 600 8835
rect 536 8771 600 8785
rect 618 8785 620 8835
rect 620 8785 676 8835
rect 676 8785 682 8835
rect 618 8771 682 8785
rect 700 8785 703 8835
rect 703 8785 759 8835
rect 759 8785 764 8835
rect 700 8771 764 8785
rect 782 8785 786 8835
rect 786 8785 842 8835
rect 842 8785 846 8835
rect 782 8771 846 8785
rect 864 8785 869 8835
rect 869 8785 925 8835
rect 925 8785 928 8835
rect 864 8771 928 8785
rect 946 8785 952 8835
rect 952 8785 1008 8835
rect 1008 8785 1010 8835
rect 946 8771 1010 8785
rect 1028 8785 1035 8835
rect 1035 8785 1091 8835
rect 1091 8785 1092 8835
rect 1028 8771 1092 8785
rect 1110 8785 1118 8835
rect 1118 8785 1174 8835
rect 1110 8771 1174 8785
rect 1192 8785 1201 8835
rect 1201 8785 1256 8835
rect 1192 8771 1256 8785
rect 204 8699 259 8751
rect 259 8699 268 8751
rect 204 8687 268 8699
rect 287 8699 343 8751
rect 343 8699 351 8751
rect 287 8687 351 8699
rect 370 8699 371 8751
rect 371 8699 427 8751
rect 427 8699 434 8751
rect 370 8687 434 8699
rect 453 8699 454 8751
rect 454 8699 510 8751
rect 510 8699 517 8751
rect 453 8687 517 8699
rect 536 8699 537 8751
rect 537 8699 593 8751
rect 593 8699 600 8751
rect 536 8687 600 8699
rect 618 8699 620 8751
rect 620 8699 676 8751
rect 676 8699 682 8751
rect 618 8687 682 8699
rect 700 8699 703 8751
rect 703 8699 759 8751
rect 759 8699 764 8751
rect 700 8687 764 8699
rect 782 8699 786 8751
rect 786 8699 842 8751
rect 842 8699 846 8751
rect 782 8687 846 8699
rect 864 8699 869 8751
rect 869 8699 925 8751
rect 925 8699 928 8751
rect 864 8687 928 8699
rect 946 8699 952 8751
rect 952 8699 1008 8751
rect 1008 8699 1010 8751
rect 946 8687 1010 8699
rect 1028 8699 1035 8751
rect 1035 8699 1091 8751
rect 1091 8699 1092 8751
rect 1028 8687 1092 8699
rect 1110 8699 1118 8751
rect 1118 8699 1174 8751
rect 1110 8687 1174 8699
rect 1192 8699 1201 8751
rect 1201 8699 1256 8751
rect 1192 8687 1256 8699
rect 204 8613 259 8667
rect 259 8613 268 8667
rect 204 8603 268 8613
rect 287 8613 343 8667
rect 343 8613 351 8667
rect 287 8603 351 8613
rect 370 8613 371 8667
rect 371 8613 427 8667
rect 427 8613 434 8667
rect 370 8603 434 8613
rect 453 8613 454 8667
rect 454 8613 510 8667
rect 510 8613 517 8667
rect 453 8603 517 8613
rect 536 8613 537 8667
rect 537 8613 593 8667
rect 593 8613 600 8667
rect 536 8603 600 8613
rect 618 8613 620 8667
rect 620 8613 676 8667
rect 676 8613 682 8667
rect 618 8603 682 8613
rect 700 8613 703 8667
rect 703 8613 759 8667
rect 759 8613 764 8667
rect 700 8603 764 8613
rect 782 8613 786 8667
rect 786 8613 842 8667
rect 842 8613 846 8667
rect 782 8603 846 8613
rect 864 8613 869 8667
rect 869 8613 925 8667
rect 925 8613 928 8667
rect 864 8603 928 8613
rect 946 8613 952 8667
rect 952 8613 1008 8667
rect 1008 8613 1010 8667
rect 946 8603 1010 8613
rect 1028 8613 1035 8667
rect 1035 8613 1091 8667
rect 1091 8613 1092 8667
rect 1028 8603 1092 8613
rect 1110 8613 1118 8667
rect 1118 8613 1174 8667
rect 1110 8603 1174 8613
rect 1192 8613 1201 8667
rect 1201 8613 1256 8667
rect 1192 8603 1256 8613
rect 204 8527 259 8583
rect 259 8527 268 8583
rect 204 8519 268 8527
rect 287 8527 343 8583
rect 343 8527 351 8583
rect 287 8519 351 8527
rect 370 8527 371 8583
rect 371 8527 427 8583
rect 427 8527 434 8583
rect 370 8519 434 8527
rect 453 8527 454 8583
rect 454 8527 510 8583
rect 510 8527 517 8583
rect 453 8519 517 8527
rect 536 8527 537 8583
rect 537 8527 593 8583
rect 593 8527 600 8583
rect 536 8519 600 8527
rect 618 8527 620 8583
rect 620 8527 676 8583
rect 676 8527 682 8583
rect 618 8519 682 8527
rect 700 8527 703 8583
rect 703 8527 759 8583
rect 759 8527 764 8583
rect 700 8519 764 8527
rect 782 8527 786 8583
rect 786 8527 842 8583
rect 842 8527 846 8583
rect 782 8519 846 8527
rect 864 8527 869 8583
rect 869 8527 925 8583
rect 925 8527 928 8583
rect 864 8519 928 8527
rect 946 8527 952 8583
rect 952 8527 1008 8583
rect 1008 8527 1010 8583
rect 946 8519 1010 8527
rect 1028 8527 1035 8583
rect 1035 8527 1091 8583
rect 1091 8527 1092 8583
rect 1028 8519 1092 8527
rect 1110 8527 1118 8583
rect 1118 8527 1174 8583
rect 1110 8519 1174 8527
rect 1192 8527 1201 8583
rect 1201 8527 1256 8583
rect 1192 8519 1256 8527
rect 204 8497 268 8499
rect 204 8441 259 8497
rect 259 8441 268 8497
rect 204 8435 268 8441
rect 287 8497 351 8499
rect 287 8441 343 8497
rect 343 8441 351 8497
rect 287 8435 351 8441
rect 370 8497 434 8499
rect 370 8441 371 8497
rect 371 8441 427 8497
rect 427 8441 434 8497
rect 370 8435 434 8441
rect 453 8497 517 8499
rect 453 8441 454 8497
rect 454 8441 510 8497
rect 510 8441 517 8497
rect 453 8435 517 8441
rect 536 8497 600 8499
rect 536 8441 537 8497
rect 537 8441 593 8497
rect 593 8441 600 8497
rect 536 8435 600 8441
rect 618 8497 682 8499
rect 618 8441 620 8497
rect 620 8441 676 8497
rect 676 8441 682 8497
rect 618 8435 682 8441
rect 700 8497 764 8499
rect 700 8441 703 8497
rect 703 8441 759 8497
rect 759 8441 764 8497
rect 700 8435 764 8441
rect 782 8497 846 8499
rect 782 8441 786 8497
rect 786 8441 842 8497
rect 842 8441 846 8497
rect 782 8435 846 8441
rect 864 8497 928 8499
rect 864 8441 869 8497
rect 869 8441 925 8497
rect 925 8441 928 8497
rect 864 8435 928 8441
rect 946 8497 1010 8499
rect 946 8441 952 8497
rect 952 8441 1008 8497
rect 1008 8441 1010 8497
rect 946 8435 1010 8441
rect 1028 8497 1092 8499
rect 1028 8441 1035 8497
rect 1035 8441 1091 8497
rect 1091 8441 1092 8497
rect 1028 8435 1092 8441
rect 1110 8497 1174 8499
rect 1110 8441 1118 8497
rect 1118 8441 1174 8497
rect 1110 8435 1174 8441
rect 1192 8497 1256 8499
rect 1192 8441 1201 8497
rect 1201 8441 1256 8497
rect 1192 8435 1256 8441
rect 204 8411 268 8415
rect 204 8355 259 8411
rect 259 8355 268 8411
rect 204 8351 268 8355
rect 287 8411 351 8415
rect 287 8355 343 8411
rect 343 8355 351 8411
rect 287 8351 351 8355
rect 370 8411 434 8415
rect 370 8355 371 8411
rect 371 8355 427 8411
rect 427 8355 434 8411
rect 370 8351 434 8355
rect 453 8411 517 8415
rect 453 8355 454 8411
rect 454 8355 510 8411
rect 510 8355 517 8411
rect 453 8351 517 8355
rect 536 8411 600 8415
rect 536 8355 537 8411
rect 537 8355 593 8411
rect 593 8355 600 8411
rect 536 8351 600 8355
rect 618 8411 682 8415
rect 618 8355 620 8411
rect 620 8355 676 8411
rect 676 8355 682 8411
rect 618 8351 682 8355
rect 700 8411 764 8415
rect 700 8355 703 8411
rect 703 8355 759 8411
rect 759 8355 764 8411
rect 700 8351 764 8355
rect 782 8411 846 8415
rect 782 8355 786 8411
rect 786 8355 842 8411
rect 842 8355 846 8411
rect 782 8351 846 8355
rect 864 8411 928 8415
rect 864 8355 869 8411
rect 869 8355 925 8411
rect 925 8355 928 8411
rect 864 8351 928 8355
rect 946 8411 1010 8415
rect 946 8355 952 8411
rect 952 8355 1008 8411
rect 1008 8355 1010 8411
rect 946 8351 1010 8355
rect 1028 8411 1092 8415
rect 1028 8355 1035 8411
rect 1035 8355 1091 8411
rect 1091 8355 1092 8411
rect 1028 8351 1092 8355
rect 1110 8411 1174 8415
rect 1110 8355 1118 8411
rect 1118 8355 1174 8411
rect 1110 8351 1174 8355
rect 1192 8411 1256 8415
rect 1192 8355 1201 8411
rect 1201 8355 1256 8411
rect 1192 8351 1256 8355
rect 204 8325 268 8331
rect 204 8269 259 8325
rect 259 8269 268 8325
rect 204 8267 268 8269
rect 287 8325 351 8331
rect 287 8269 343 8325
rect 343 8269 351 8325
rect 287 8267 351 8269
rect 370 8325 434 8331
rect 370 8269 371 8325
rect 371 8269 427 8325
rect 427 8269 434 8325
rect 370 8267 434 8269
rect 453 8325 517 8331
rect 453 8269 454 8325
rect 454 8269 510 8325
rect 510 8269 517 8325
rect 453 8267 517 8269
rect 536 8325 600 8331
rect 536 8269 537 8325
rect 537 8269 593 8325
rect 593 8269 600 8325
rect 536 8267 600 8269
rect 618 8325 682 8331
rect 618 8269 620 8325
rect 620 8269 676 8325
rect 676 8269 682 8325
rect 618 8267 682 8269
rect 700 8325 764 8331
rect 700 8269 703 8325
rect 703 8269 759 8325
rect 759 8269 764 8325
rect 700 8267 764 8269
rect 782 8325 846 8331
rect 782 8269 786 8325
rect 786 8269 842 8325
rect 842 8269 846 8325
rect 782 8267 846 8269
rect 864 8325 928 8331
rect 864 8269 869 8325
rect 869 8269 925 8325
rect 925 8269 928 8325
rect 864 8267 928 8269
rect 946 8325 1010 8331
rect 946 8269 952 8325
rect 952 8269 1008 8325
rect 1008 8269 1010 8325
rect 946 8267 1010 8269
rect 1028 8325 1092 8331
rect 1028 8269 1035 8325
rect 1035 8269 1091 8325
rect 1091 8269 1092 8325
rect 1028 8267 1092 8269
rect 1110 8325 1174 8331
rect 1110 8269 1118 8325
rect 1118 8269 1174 8325
rect 1110 8267 1174 8269
rect 1192 8325 1256 8331
rect 1192 8269 1201 8325
rect 1201 8269 1256 8325
rect 1192 8267 1256 8269
rect 204 8239 268 8247
rect 204 8183 259 8239
rect 259 8183 268 8239
rect 287 8239 351 8247
rect 287 8183 343 8239
rect 343 8183 351 8239
rect 370 8239 434 8247
rect 370 8183 371 8239
rect 371 8183 427 8239
rect 427 8183 434 8239
rect 453 8239 517 8247
rect 453 8183 454 8239
rect 454 8183 510 8239
rect 510 8183 517 8239
rect 536 8239 600 8247
rect 536 8183 537 8239
rect 537 8183 593 8239
rect 593 8183 600 8239
rect 618 8239 682 8247
rect 618 8183 620 8239
rect 620 8183 676 8239
rect 676 8183 682 8239
rect 700 8239 764 8247
rect 700 8183 703 8239
rect 703 8183 759 8239
rect 759 8183 764 8239
rect 782 8239 846 8247
rect 782 8183 786 8239
rect 786 8183 842 8239
rect 842 8183 846 8239
rect 864 8239 928 8247
rect 864 8183 869 8239
rect 869 8183 925 8239
rect 925 8183 928 8239
rect 946 8239 1010 8247
rect 946 8183 952 8239
rect 952 8183 1008 8239
rect 1008 8183 1010 8239
rect 1028 8239 1092 8247
rect 1028 8183 1035 8239
rect 1035 8183 1091 8239
rect 1091 8183 1092 8239
rect 1110 8239 1174 8247
rect 1110 8183 1118 8239
rect 1118 8183 1174 8239
rect 1192 8239 1256 8247
rect 1192 8183 1201 8239
rect 1201 8183 1256 8239
rect 204 8153 268 8163
rect 204 8099 259 8153
rect 259 8099 268 8153
rect 287 8153 351 8163
rect 287 8099 343 8153
rect 343 8099 351 8153
rect 370 8153 434 8163
rect 370 8099 371 8153
rect 371 8099 427 8153
rect 427 8099 434 8153
rect 453 8153 517 8163
rect 453 8099 454 8153
rect 454 8099 510 8153
rect 510 8099 517 8153
rect 536 8153 600 8163
rect 536 8099 537 8153
rect 537 8099 593 8153
rect 593 8099 600 8153
rect 618 8153 682 8163
rect 618 8099 620 8153
rect 620 8099 676 8153
rect 676 8099 682 8153
rect 700 8153 764 8163
rect 700 8099 703 8153
rect 703 8099 759 8153
rect 759 8099 764 8153
rect 782 8153 846 8163
rect 782 8099 786 8153
rect 786 8099 842 8153
rect 842 8099 846 8153
rect 864 8153 928 8163
rect 864 8099 869 8153
rect 869 8099 925 8153
rect 925 8099 928 8153
rect 946 8153 1010 8163
rect 946 8099 952 8153
rect 952 8099 1008 8153
rect 1008 8099 1010 8153
rect 1028 8153 1092 8163
rect 1028 8099 1035 8153
rect 1035 8099 1091 8153
rect 1091 8099 1092 8153
rect 1110 8153 1174 8163
rect 1110 8099 1118 8153
rect 1118 8099 1174 8153
rect 1192 8153 1256 8163
rect 1192 8099 1201 8153
rect 1201 8099 1256 8153
rect 204 8067 268 8079
rect 204 8015 259 8067
rect 259 8015 268 8067
rect 287 8067 351 8079
rect 287 8015 343 8067
rect 343 8015 351 8067
rect 370 8067 434 8079
rect 370 8015 371 8067
rect 371 8015 427 8067
rect 427 8015 434 8067
rect 453 8067 517 8079
rect 453 8015 454 8067
rect 454 8015 510 8067
rect 510 8015 517 8067
rect 536 8067 600 8079
rect 536 8015 537 8067
rect 537 8015 593 8067
rect 593 8015 600 8067
rect 618 8067 682 8079
rect 618 8015 620 8067
rect 620 8015 676 8067
rect 676 8015 682 8067
rect 700 8067 764 8079
rect 700 8015 703 8067
rect 703 8015 759 8067
rect 759 8015 764 8067
rect 782 8067 846 8079
rect 782 8015 786 8067
rect 786 8015 842 8067
rect 842 8015 846 8067
rect 864 8067 928 8079
rect 864 8015 869 8067
rect 869 8015 925 8067
rect 925 8015 928 8067
rect 946 8067 1010 8079
rect 946 8015 952 8067
rect 952 8015 1008 8067
rect 1008 8015 1010 8067
rect 1028 8067 1092 8079
rect 1028 8015 1035 8067
rect 1035 8015 1091 8067
rect 1091 8015 1092 8067
rect 1110 8067 1174 8079
rect 1110 8015 1118 8067
rect 1118 8015 1174 8067
rect 1192 8067 1256 8079
rect 1192 8015 1201 8067
rect 1201 8015 1256 8067
rect 204 7981 268 7995
rect 204 7931 259 7981
rect 259 7931 268 7981
rect 287 7981 351 7995
rect 287 7931 343 7981
rect 343 7931 351 7981
rect 370 7981 434 7995
rect 370 7931 371 7981
rect 371 7931 427 7981
rect 427 7931 434 7981
rect 453 7981 517 7995
rect 453 7931 454 7981
rect 454 7931 510 7981
rect 510 7931 517 7981
rect 536 7981 600 7995
rect 536 7931 537 7981
rect 537 7931 593 7981
rect 593 7931 600 7981
rect 618 7981 682 7995
rect 618 7931 620 7981
rect 620 7931 676 7981
rect 676 7931 682 7981
rect 700 7981 764 7995
rect 700 7931 703 7981
rect 703 7931 759 7981
rect 759 7931 764 7981
rect 782 7981 846 7995
rect 782 7931 786 7981
rect 786 7931 842 7981
rect 842 7931 846 7981
rect 864 7981 928 7995
rect 864 7931 869 7981
rect 869 7931 925 7981
rect 925 7931 928 7981
rect 946 7981 1010 7995
rect 946 7931 952 7981
rect 952 7931 1008 7981
rect 1008 7931 1010 7981
rect 1028 7981 1092 7995
rect 1028 7931 1035 7981
rect 1035 7931 1091 7981
rect 1091 7931 1092 7981
rect 1110 7981 1174 7995
rect 1110 7931 1118 7981
rect 1118 7931 1174 7981
rect 1192 7981 1256 7995
rect 1192 7931 1201 7981
rect 1201 7931 1256 7981
rect 8224 8785 8259 8829
rect 8259 8785 8287 8829
rect 8287 8785 8288 8829
rect 8305 8785 8343 8829
rect 8343 8785 8369 8829
rect 8386 8785 8426 8829
rect 8426 8785 8450 8829
rect 8466 8785 8509 8829
rect 8509 8785 8530 8829
rect 8546 8785 8592 8829
rect 8592 8785 8610 8829
rect 8626 8785 8675 8829
rect 8675 8785 8690 8829
rect 8706 8785 8758 8829
rect 8758 8785 8770 8829
rect 8786 8785 8841 8829
rect 8841 8785 8850 8829
rect 8224 8765 8288 8785
rect 8305 8765 8369 8785
rect 8386 8765 8450 8785
rect 8466 8765 8530 8785
rect 8546 8765 8610 8785
rect 8626 8765 8690 8785
rect 8706 8765 8770 8785
rect 8786 8765 8850 8785
rect 8866 8785 8868 8829
rect 8868 8785 8924 8829
rect 8924 8785 8930 8829
rect 8866 8765 8930 8785
rect 8946 8785 8951 8829
rect 8951 8785 9007 8829
rect 9007 8785 9010 8829
rect 8946 8765 9010 8785
rect 9026 8785 9034 8829
rect 9034 8785 9090 8829
rect 9026 8765 9090 8785
rect 9106 8785 9117 8829
rect 9117 8785 9170 8829
rect 9186 8785 9200 8829
rect 9200 8785 9250 8829
rect 9106 8765 9170 8785
rect 9186 8765 9250 8785
rect 8224 8699 8259 8745
rect 8259 8699 8287 8745
rect 8287 8699 8288 8745
rect 8305 8699 8343 8745
rect 8343 8699 8369 8745
rect 8386 8699 8426 8745
rect 8426 8699 8450 8745
rect 8466 8699 8509 8745
rect 8509 8699 8530 8745
rect 8546 8699 8592 8745
rect 8592 8699 8610 8745
rect 8626 8699 8675 8745
rect 8675 8699 8690 8745
rect 8706 8699 8758 8745
rect 8758 8699 8770 8745
rect 8786 8699 8841 8745
rect 8841 8699 8850 8745
rect 8224 8681 8288 8699
rect 8305 8681 8369 8699
rect 8386 8681 8450 8699
rect 8466 8681 8530 8699
rect 8546 8681 8610 8699
rect 8626 8681 8690 8699
rect 8706 8681 8770 8699
rect 8786 8681 8850 8699
rect 8866 8699 8868 8745
rect 8868 8699 8924 8745
rect 8924 8699 8930 8745
rect 8866 8681 8930 8699
rect 8946 8699 8951 8745
rect 8951 8699 9007 8745
rect 9007 8699 9010 8745
rect 8946 8681 9010 8699
rect 9026 8699 9034 8745
rect 9034 8699 9090 8745
rect 9026 8681 9090 8699
rect 9106 8699 9117 8745
rect 9117 8699 9170 8745
rect 9186 8699 9200 8745
rect 9200 8699 9250 8745
rect 9106 8681 9170 8699
rect 9186 8681 9250 8699
rect 8224 8613 8259 8661
rect 8259 8613 8287 8661
rect 8287 8613 8288 8661
rect 8305 8613 8343 8661
rect 8343 8613 8369 8661
rect 8386 8613 8426 8661
rect 8426 8613 8450 8661
rect 8466 8613 8509 8661
rect 8509 8613 8530 8661
rect 8546 8613 8592 8661
rect 8592 8613 8610 8661
rect 8626 8613 8675 8661
rect 8675 8613 8690 8661
rect 8706 8613 8758 8661
rect 8758 8613 8770 8661
rect 8786 8613 8841 8661
rect 8841 8613 8850 8661
rect 8224 8597 8288 8613
rect 8305 8597 8369 8613
rect 8386 8597 8450 8613
rect 8466 8597 8530 8613
rect 8546 8597 8610 8613
rect 8626 8597 8690 8613
rect 8706 8597 8770 8613
rect 8786 8597 8850 8613
rect 8866 8613 8868 8661
rect 8868 8613 8924 8661
rect 8924 8613 8930 8661
rect 8866 8597 8930 8613
rect 8946 8613 8951 8661
rect 8951 8613 9007 8661
rect 9007 8613 9010 8661
rect 8946 8597 9010 8613
rect 9026 8613 9034 8661
rect 9034 8613 9090 8661
rect 9026 8597 9090 8613
rect 9106 8613 9117 8661
rect 9117 8613 9170 8661
rect 9186 8613 9200 8661
rect 9200 8613 9250 8661
rect 9106 8597 9170 8613
rect 9186 8597 9250 8613
rect 8224 8527 8259 8577
rect 8259 8527 8287 8577
rect 8287 8527 8288 8577
rect 8305 8527 8343 8577
rect 8343 8527 8369 8577
rect 8386 8527 8426 8577
rect 8426 8527 8450 8577
rect 8466 8527 8509 8577
rect 8509 8527 8530 8577
rect 8546 8527 8592 8577
rect 8592 8527 8610 8577
rect 8626 8527 8675 8577
rect 8675 8527 8690 8577
rect 8706 8527 8758 8577
rect 8758 8527 8770 8577
rect 8786 8527 8841 8577
rect 8841 8527 8850 8577
rect 8224 8513 8288 8527
rect 8305 8513 8369 8527
rect 8386 8513 8450 8527
rect 8466 8513 8530 8527
rect 8546 8513 8610 8527
rect 8626 8513 8690 8527
rect 8706 8513 8770 8527
rect 8786 8513 8850 8527
rect 8866 8527 8868 8577
rect 8868 8527 8924 8577
rect 8924 8527 8930 8577
rect 8866 8513 8930 8527
rect 8946 8527 8951 8577
rect 8951 8527 9007 8577
rect 9007 8527 9010 8577
rect 8946 8513 9010 8527
rect 9026 8527 9034 8577
rect 9034 8527 9090 8577
rect 9026 8513 9090 8527
rect 9106 8527 9117 8577
rect 9117 8527 9170 8577
rect 9186 8527 9200 8577
rect 9200 8527 9250 8577
rect 9106 8513 9170 8527
rect 9186 8513 9250 8527
rect 8224 8441 8259 8493
rect 8259 8441 8287 8493
rect 8287 8441 8288 8493
rect 8305 8441 8343 8493
rect 8343 8441 8369 8493
rect 8386 8441 8426 8493
rect 8426 8441 8450 8493
rect 8466 8441 8509 8493
rect 8509 8441 8530 8493
rect 8546 8441 8592 8493
rect 8592 8441 8610 8493
rect 8626 8441 8675 8493
rect 8675 8441 8690 8493
rect 8706 8441 8758 8493
rect 8758 8441 8770 8493
rect 8786 8441 8841 8493
rect 8841 8441 8850 8493
rect 8224 8429 8288 8441
rect 8305 8429 8369 8441
rect 8386 8429 8450 8441
rect 8466 8429 8530 8441
rect 8546 8429 8610 8441
rect 8626 8429 8690 8441
rect 8706 8429 8770 8441
rect 8786 8429 8850 8441
rect 8866 8441 8868 8493
rect 8868 8441 8924 8493
rect 8924 8441 8930 8493
rect 8866 8429 8930 8441
rect 8946 8441 8951 8493
rect 8951 8441 9007 8493
rect 9007 8441 9010 8493
rect 8946 8429 9010 8441
rect 9026 8441 9034 8493
rect 9034 8441 9090 8493
rect 9026 8429 9090 8441
rect 9106 8441 9117 8493
rect 9117 8441 9170 8493
rect 9186 8441 9200 8493
rect 9200 8441 9250 8493
rect 9106 8429 9170 8441
rect 9186 8429 9250 8441
rect 8224 8355 8259 8409
rect 8259 8355 8287 8409
rect 8287 8355 8288 8409
rect 8305 8355 8343 8409
rect 8343 8355 8369 8409
rect 8386 8355 8426 8409
rect 8426 8355 8450 8409
rect 8466 8355 8509 8409
rect 8509 8355 8530 8409
rect 8546 8355 8592 8409
rect 8592 8355 8610 8409
rect 8626 8355 8675 8409
rect 8675 8355 8690 8409
rect 8706 8355 8758 8409
rect 8758 8355 8770 8409
rect 8786 8355 8841 8409
rect 8841 8355 8850 8409
rect 8224 8345 8288 8355
rect 8305 8345 8369 8355
rect 8386 8345 8450 8355
rect 8466 8345 8530 8355
rect 8546 8345 8610 8355
rect 8626 8345 8690 8355
rect 8706 8345 8770 8355
rect 8786 8345 8850 8355
rect 8866 8355 8868 8409
rect 8868 8355 8924 8409
rect 8924 8355 8930 8409
rect 8866 8345 8930 8355
rect 8946 8355 8951 8409
rect 8951 8355 9007 8409
rect 9007 8355 9010 8409
rect 8946 8345 9010 8355
rect 9026 8355 9034 8409
rect 9034 8355 9090 8409
rect 9026 8345 9090 8355
rect 9106 8355 9117 8409
rect 9117 8355 9170 8409
rect 9186 8355 9200 8409
rect 9200 8355 9250 8409
rect 9106 8345 9170 8355
rect 9186 8345 9250 8355
rect 8224 8269 8259 8325
rect 8259 8269 8287 8325
rect 8287 8269 8288 8325
rect 8305 8269 8343 8325
rect 8343 8269 8369 8325
rect 8386 8269 8426 8325
rect 8426 8269 8450 8325
rect 8466 8269 8509 8325
rect 8509 8269 8530 8325
rect 8546 8269 8592 8325
rect 8592 8269 8610 8325
rect 8626 8269 8675 8325
rect 8675 8269 8690 8325
rect 8706 8269 8758 8325
rect 8758 8269 8770 8325
rect 8786 8269 8841 8325
rect 8841 8269 8850 8325
rect 8224 8261 8288 8269
rect 8305 8261 8369 8269
rect 8386 8261 8450 8269
rect 8466 8261 8530 8269
rect 8546 8261 8610 8269
rect 8626 8261 8690 8269
rect 8706 8261 8770 8269
rect 8786 8261 8850 8269
rect 8866 8269 8868 8325
rect 8868 8269 8924 8325
rect 8924 8269 8930 8325
rect 8866 8261 8930 8269
rect 8946 8269 8951 8325
rect 8951 8269 9007 8325
rect 9007 8269 9010 8325
rect 8946 8261 9010 8269
rect 9026 8269 9034 8325
rect 9034 8269 9090 8325
rect 9026 8261 9090 8269
rect 9106 8269 9117 8325
rect 9117 8269 9170 8325
rect 9186 8269 9200 8325
rect 9200 8269 9250 8325
rect 9106 8261 9170 8269
rect 9186 8261 9250 8269
rect 8224 8239 8288 8241
rect 8305 8239 8369 8241
rect 8386 8239 8450 8241
rect 8466 8239 8530 8241
rect 8546 8239 8610 8241
rect 8626 8239 8690 8241
rect 8706 8239 8770 8241
rect 8786 8239 8850 8241
rect 8224 8183 8259 8239
rect 8259 8183 8287 8239
rect 8287 8183 8288 8239
rect 8305 8183 8343 8239
rect 8343 8183 8369 8239
rect 8386 8183 8426 8239
rect 8426 8183 8450 8239
rect 8466 8183 8509 8239
rect 8509 8183 8530 8239
rect 8546 8183 8592 8239
rect 8592 8183 8610 8239
rect 8626 8183 8675 8239
rect 8675 8183 8690 8239
rect 8706 8183 8758 8239
rect 8758 8183 8770 8239
rect 8786 8183 8841 8239
rect 8841 8183 8850 8239
rect 8224 8177 8288 8183
rect 8305 8177 8369 8183
rect 8386 8177 8450 8183
rect 8466 8177 8530 8183
rect 8546 8177 8610 8183
rect 8626 8177 8690 8183
rect 8706 8177 8770 8183
rect 8786 8177 8850 8183
rect 8866 8239 8930 8241
rect 8866 8183 8868 8239
rect 8868 8183 8924 8239
rect 8924 8183 8930 8239
rect 8866 8177 8930 8183
rect 8946 8239 9010 8241
rect 8946 8183 8951 8239
rect 8951 8183 9007 8239
rect 9007 8183 9010 8239
rect 8946 8177 9010 8183
rect 9026 8239 9090 8241
rect 9026 8183 9034 8239
rect 9034 8183 9090 8239
rect 9026 8177 9090 8183
rect 9106 8239 9170 8241
rect 9186 8239 9250 8241
rect 9106 8183 9117 8239
rect 9117 8183 9170 8239
rect 9186 8183 9200 8239
rect 9200 8183 9250 8239
rect 9106 8177 9170 8183
rect 9186 8177 9250 8183
rect 8224 8153 8288 8157
rect 8305 8153 8369 8157
rect 8386 8153 8450 8157
rect 8466 8153 8530 8157
rect 8546 8153 8610 8157
rect 8626 8153 8690 8157
rect 8706 8153 8770 8157
rect 8786 8153 8850 8157
rect 8224 8097 8259 8153
rect 8259 8097 8287 8153
rect 8287 8097 8288 8153
rect 8305 8097 8343 8153
rect 8343 8097 8369 8153
rect 8386 8097 8426 8153
rect 8426 8097 8450 8153
rect 8466 8097 8509 8153
rect 8509 8097 8530 8153
rect 8546 8097 8592 8153
rect 8592 8097 8610 8153
rect 8626 8097 8675 8153
rect 8675 8097 8690 8153
rect 8706 8097 8758 8153
rect 8758 8097 8770 8153
rect 8786 8097 8841 8153
rect 8841 8097 8850 8153
rect 8224 8093 8288 8097
rect 8305 8093 8369 8097
rect 8386 8093 8450 8097
rect 8466 8093 8530 8097
rect 8546 8093 8610 8097
rect 8626 8093 8690 8097
rect 8706 8093 8770 8097
rect 8786 8093 8850 8097
rect 8866 8153 8930 8157
rect 8866 8097 8868 8153
rect 8868 8097 8924 8153
rect 8924 8097 8930 8153
rect 8866 8093 8930 8097
rect 8946 8153 9010 8157
rect 8946 8097 8951 8153
rect 8951 8097 9007 8153
rect 9007 8097 9010 8153
rect 8946 8093 9010 8097
rect 9026 8153 9090 8157
rect 9026 8097 9034 8153
rect 9034 8097 9090 8153
rect 9026 8093 9090 8097
rect 9106 8153 9170 8157
rect 9186 8153 9250 8157
rect 9106 8097 9117 8153
rect 9117 8097 9170 8153
rect 9186 8097 9200 8153
rect 9200 8097 9250 8153
rect 9106 8093 9170 8097
rect 9186 8093 9250 8097
rect 8224 8067 8288 8073
rect 8305 8067 8369 8073
rect 8386 8067 8450 8073
rect 8466 8067 8530 8073
rect 8546 8067 8610 8073
rect 8626 8067 8690 8073
rect 8706 8067 8770 8073
rect 8786 8067 8850 8073
rect 8224 8011 8259 8067
rect 8259 8011 8287 8067
rect 8287 8011 8288 8067
rect 8305 8011 8343 8067
rect 8343 8011 8369 8067
rect 8386 8011 8426 8067
rect 8426 8011 8450 8067
rect 8466 8011 8509 8067
rect 8509 8011 8530 8067
rect 8546 8011 8592 8067
rect 8592 8011 8610 8067
rect 8626 8011 8675 8067
rect 8675 8011 8690 8067
rect 8706 8011 8758 8067
rect 8758 8011 8770 8067
rect 8786 8011 8841 8067
rect 8841 8011 8850 8067
rect 8224 8009 8288 8011
rect 8305 8009 8369 8011
rect 8386 8009 8450 8011
rect 8466 8009 8530 8011
rect 8546 8009 8610 8011
rect 8626 8009 8690 8011
rect 8706 8009 8770 8011
rect 8786 8009 8850 8011
rect 8866 8067 8930 8073
rect 8866 8011 8868 8067
rect 8868 8011 8924 8067
rect 8924 8011 8930 8067
rect 8866 8009 8930 8011
rect 8946 8067 9010 8073
rect 8946 8011 8951 8067
rect 8951 8011 9007 8067
rect 9007 8011 9010 8067
rect 8946 8009 9010 8011
rect 9026 8067 9090 8073
rect 9026 8011 9034 8067
rect 9034 8011 9090 8067
rect 9026 8009 9090 8011
rect 9106 8067 9170 8073
rect 9186 8067 9250 8073
rect 9106 8011 9117 8067
rect 9117 8011 9170 8067
rect 9186 8011 9200 8067
rect 9200 8011 9250 8067
rect 9106 8009 9170 8011
rect 9186 8009 9250 8011
rect 8224 7981 8288 7989
rect 8305 7981 8369 7989
rect 8386 7981 8450 7989
rect 8466 7981 8530 7989
rect 8546 7981 8610 7989
rect 8626 7981 8690 7989
rect 8706 7981 8770 7989
rect 8786 7981 8850 7989
rect 8224 7925 8259 7981
rect 8259 7925 8287 7981
rect 8287 7925 8288 7981
rect 8305 7925 8343 7981
rect 8343 7925 8369 7981
rect 8386 7925 8426 7981
rect 8426 7925 8450 7981
rect 8466 7925 8509 7981
rect 8509 7925 8530 7981
rect 8546 7925 8592 7981
rect 8592 7925 8610 7981
rect 8626 7925 8675 7981
rect 8675 7925 8690 7981
rect 8706 7925 8758 7981
rect 8758 7925 8770 7981
rect 8786 7925 8841 7981
rect 8841 7925 8850 7981
rect 8866 7981 8930 7989
rect 8866 7925 8868 7981
rect 8868 7925 8924 7981
rect 8924 7925 8930 7981
rect 8946 7981 9010 7989
rect 8946 7925 8951 7981
rect 8951 7925 9007 7981
rect 9007 7925 9010 7981
rect 9026 7981 9090 7989
rect 9026 7925 9034 7981
rect 9034 7925 9090 7981
rect 9106 7981 9170 7989
rect 9186 7981 9250 7989
rect 9106 7925 9117 7981
rect 9117 7925 9170 7981
rect 9186 7925 9200 7981
rect 9200 7925 9250 7981
<< metal4 >>
rect 0 39592 15000 39600
rect 0 39528 462 39592
rect 526 39528 620 39592
rect 684 39528 1390 39592
rect 1454 39528 1518 39592
rect 1582 39528 2382 39592
rect 2446 39528 2510 39592
rect 2574 39528 3374 39592
rect 3438 39528 3502 39592
rect 3566 39528 4366 39592
rect 4430 39528 4494 39592
rect 4558 39528 5358 39592
rect 5422 39528 5486 39592
rect 5550 39528 6350 39592
rect 6414 39528 6478 39592
rect 6542 39528 7342 39592
rect 7406 39528 7470 39592
rect 7534 39528 8334 39592
rect 8398 39528 8462 39592
rect 8526 39528 9326 39592
rect 9390 39528 9454 39592
rect 9518 39528 10318 39592
rect 10382 39528 10446 39592
rect 10510 39528 11310 39592
rect 11374 39528 11438 39592
rect 11502 39528 12302 39592
rect 12366 39528 12430 39592
rect 12494 39528 13294 39592
rect 13358 39528 13422 39592
rect 13486 39528 14255 39592
rect 14319 39528 14343 39592
rect 14407 39528 14431 39592
rect 14495 39528 14519 39592
rect 14583 39528 14607 39592
rect 14671 39528 15000 39592
rect 0 39512 15000 39528
rect 0 39448 462 39512
rect 526 39448 620 39512
rect 684 39448 1390 39512
rect 1454 39448 1518 39512
rect 1582 39448 2382 39512
rect 2446 39448 2510 39512
rect 2574 39448 3374 39512
rect 3438 39448 3502 39512
rect 3566 39448 4366 39512
rect 4430 39448 4494 39512
rect 4558 39448 5358 39512
rect 5422 39448 5486 39512
rect 5550 39448 6350 39512
rect 6414 39448 6478 39512
rect 6542 39448 7342 39512
rect 7406 39448 7470 39512
rect 7534 39448 8334 39512
rect 8398 39448 8462 39512
rect 8526 39448 9326 39512
rect 9390 39448 9454 39512
rect 9518 39448 10318 39512
rect 10382 39448 10446 39512
rect 10510 39448 11310 39512
rect 11374 39448 11438 39512
rect 11502 39448 12302 39512
rect 12366 39448 12430 39512
rect 12494 39448 13294 39512
rect 13358 39448 13422 39512
rect 13486 39448 14255 39512
rect 14319 39448 14343 39512
rect 14407 39448 14431 39512
rect 14495 39448 14519 39512
rect 14583 39448 14607 39512
rect 14671 39448 15000 39512
rect 0 39432 15000 39448
rect 0 39368 462 39432
rect 526 39368 620 39432
rect 684 39368 1390 39432
rect 1454 39368 1518 39432
rect 1582 39368 2382 39432
rect 2446 39368 2510 39432
rect 2574 39368 3374 39432
rect 3438 39368 3502 39432
rect 3566 39368 4366 39432
rect 4430 39368 4494 39432
rect 4558 39368 5358 39432
rect 5422 39368 5486 39432
rect 5550 39368 6350 39432
rect 6414 39368 6478 39432
rect 6542 39368 7342 39432
rect 7406 39368 7470 39432
rect 7534 39368 8334 39432
rect 8398 39368 8462 39432
rect 8526 39368 9326 39432
rect 9390 39368 9454 39432
rect 9518 39368 10318 39432
rect 10382 39368 10446 39432
rect 10510 39368 11310 39432
rect 11374 39368 11438 39432
rect 11502 39368 12302 39432
rect 12366 39368 12430 39432
rect 12494 39368 13294 39432
rect 13358 39368 13422 39432
rect 13486 39368 14255 39432
rect 14319 39368 14343 39432
rect 14407 39368 14431 39432
rect 14495 39368 14519 39432
rect 14583 39368 14607 39432
rect 14671 39368 15000 39432
rect 0 39352 15000 39368
rect 0 39288 462 39352
rect 526 39288 620 39352
rect 684 39288 1390 39352
rect 1454 39288 1518 39352
rect 1582 39288 2382 39352
rect 2446 39288 2510 39352
rect 2574 39288 3374 39352
rect 3438 39288 3502 39352
rect 3566 39288 4366 39352
rect 4430 39288 4494 39352
rect 4558 39288 5358 39352
rect 5422 39288 5486 39352
rect 5550 39288 6350 39352
rect 6414 39288 6478 39352
rect 6542 39288 7342 39352
rect 7406 39288 7470 39352
rect 7534 39288 8334 39352
rect 8398 39288 8462 39352
rect 8526 39288 9326 39352
rect 9390 39288 9454 39352
rect 9518 39288 10318 39352
rect 10382 39288 10446 39352
rect 10510 39288 11310 39352
rect 11374 39288 11438 39352
rect 11502 39288 12302 39352
rect 12366 39288 12430 39352
rect 12494 39288 13294 39352
rect 13358 39288 13422 39352
rect 13486 39288 14255 39352
rect 14319 39288 14343 39352
rect 14407 39288 14431 39352
rect 14495 39288 14519 39352
rect 14583 39288 14607 39352
rect 14671 39288 15000 39352
rect 0 39272 15000 39288
rect 0 39208 462 39272
rect 526 39208 620 39272
rect 684 39208 1390 39272
rect 1454 39208 1518 39272
rect 1582 39208 2382 39272
rect 2446 39208 2510 39272
rect 2574 39208 3374 39272
rect 3438 39208 3502 39272
rect 3566 39208 4366 39272
rect 4430 39208 4494 39272
rect 4558 39208 5358 39272
rect 5422 39208 5486 39272
rect 5550 39208 6350 39272
rect 6414 39208 6478 39272
rect 6542 39208 7342 39272
rect 7406 39208 7470 39272
rect 7534 39208 8334 39272
rect 8398 39208 8462 39272
rect 8526 39208 9326 39272
rect 9390 39208 9454 39272
rect 9518 39208 10318 39272
rect 10382 39208 10446 39272
rect 10510 39208 11310 39272
rect 11374 39208 11438 39272
rect 11502 39208 12302 39272
rect 12366 39208 12430 39272
rect 12494 39208 13294 39272
rect 13358 39208 13422 39272
rect 13486 39208 14255 39272
rect 14319 39208 14343 39272
rect 14407 39208 14431 39272
rect 14495 39208 14519 39272
rect 14583 39208 14607 39272
rect 14671 39208 15000 39272
rect 0 39192 15000 39208
rect 0 39128 462 39192
rect 526 39128 620 39192
rect 684 39128 1390 39192
rect 1454 39128 1518 39192
rect 1582 39128 2382 39192
rect 2446 39128 2510 39192
rect 2574 39128 3374 39192
rect 3438 39128 3502 39192
rect 3566 39128 4366 39192
rect 4430 39128 4494 39192
rect 4558 39128 5358 39192
rect 5422 39128 5486 39192
rect 5550 39128 6350 39192
rect 6414 39128 6478 39192
rect 6542 39128 7342 39192
rect 7406 39128 7470 39192
rect 7534 39128 8334 39192
rect 8398 39128 8462 39192
rect 8526 39128 9326 39192
rect 9390 39128 9454 39192
rect 9518 39128 10318 39192
rect 10382 39128 10446 39192
rect 10510 39128 11310 39192
rect 11374 39128 11438 39192
rect 11502 39128 12302 39192
rect 12366 39128 12430 39192
rect 12494 39128 13294 39192
rect 13358 39128 13422 39192
rect 13486 39128 14255 39192
rect 14319 39128 14343 39192
rect 14407 39128 14431 39192
rect 14495 39128 14519 39192
rect 14583 39128 14607 39192
rect 14671 39128 15000 39192
rect 0 39112 15000 39128
rect 0 39048 462 39112
rect 526 39048 620 39112
rect 684 39048 1390 39112
rect 1454 39048 1518 39112
rect 1582 39048 2382 39112
rect 2446 39048 2510 39112
rect 2574 39048 3374 39112
rect 3438 39048 3502 39112
rect 3566 39048 4366 39112
rect 4430 39048 4494 39112
rect 4558 39048 5358 39112
rect 5422 39048 5486 39112
rect 5550 39048 6350 39112
rect 6414 39048 6478 39112
rect 6542 39048 7342 39112
rect 7406 39048 7470 39112
rect 7534 39048 8334 39112
rect 8398 39048 8462 39112
rect 8526 39048 9326 39112
rect 9390 39048 9454 39112
rect 9518 39048 10318 39112
rect 10382 39048 10446 39112
rect 10510 39048 11310 39112
rect 11374 39048 11438 39112
rect 11502 39048 12302 39112
rect 12366 39048 12430 39112
rect 12494 39048 13294 39112
rect 13358 39048 13422 39112
rect 13486 39048 14255 39112
rect 14319 39048 14343 39112
rect 14407 39048 14431 39112
rect 14495 39048 14519 39112
rect 14583 39048 14607 39112
rect 14671 39048 15000 39112
rect 0 39032 15000 39048
rect 0 38968 462 39032
rect 526 38968 620 39032
rect 684 38968 1390 39032
rect 1454 38968 1518 39032
rect 1582 38968 2382 39032
rect 2446 38968 2510 39032
rect 2574 38968 3374 39032
rect 3438 38968 3502 39032
rect 3566 38968 4366 39032
rect 4430 38968 4494 39032
rect 4558 38968 5358 39032
rect 5422 38968 5486 39032
rect 5550 38968 6350 39032
rect 6414 38968 6478 39032
rect 6542 38968 7342 39032
rect 7406 38968 7470 39032
rect 7534 38968 8334 39032
rect 8398 38968 8462 39032
rect 8526 38968 9326 39032
rect 9390 38968 9454 39032
rect 9518 38968 10318 39032
rect 10382 38968 10446 39032
rect 10510 38968 11310 39032
rect 11374 38968 11438 39032
rect 11502 38968 12302 39032
rect 12366 38968 12430 39032
rect 12494 38968 13294 39032
rect 13358 38968 13422 39032
rect 13486 38968 14255 39032
rect 14319 38968 14343 39032
rect 14407 38968 14431 39032
rect 14495 38968 14519 39032
rect 14583 38968 14607 39032
rect 14671 38968 15000 39032
rect 0 38952 15000 38968
rect 0 38888 462 38952
rect 526 38888 620 38952
rect 684 38888 1390 38952
rect 1454 38888 1518 38952
rect 1582 38888 2382 38952
rect 2446 38888 2510 38952
rect 2574 38888 3374 38952
rect 3438 38888 3502 38952
rect 3566 38888 4366 38952
rect 4430 38888 4494 38952
rect 4558 38888 5358 38952
rect 5422 38888 5486 38952
rect 5550 38888 6350 38952
rect 6414 38888 6478 38952
rect 6542 38888 7342 38952
rect 7406 38888 7470 38952
rect 7534 38888 8334 38952
rect 8398 38888 8462 38952
rect 8526 38888 9326 38952
rect 9390 38888 9454 38952
rect 9518 38888 10318 38952
rect 10382 38888 10446 38952
rect 10510 38888 11310 38952
rect 11374 38888 11438 38952
rect 11502 38888 12302 38952
rect 12366 38888 12430 38952
rect 12494 38888 13294 38952
rect 13358 38888 13422 38952
rect 13486 38888 14255 38952
rect 14319 38888 14343 38952
rect 14407 38888 14431 38952
rect 14495 38888 14519 38952
rect 14583 38888 14607 38952
rect 14671 38888 15000 38952
rect 0 38872 15000 38888
rect 0 38808 462 38872
rect 526 38808 620 38872
rect 684 38808 1390 38872
rect 1454 38808 1518 38872
rect 1582 38808 2382 38872
rect 2446 38808 2510 38872
rect 2574 38808 3374 38872
rect 3438 38808 3502 38872
rect 3566 38808 4366 38872
rect 4430 38808 4494 38872
rect 4558 38808 5358 38872
rect 5422 38808 5486 38872
rect 5550 38808 6350 38872
rect 6414 38808 6478 38872
rect 6542 38808 7342 38872
rect 7406 38808 7470 38872
rect 7534 38808 8334 38872
rect 8398 38808 8462 38872
rect 8526 38808 9326 38872
rect 9390 38808 9454 38872
rect 9518 38808 10318 38872
rect 10382 38808 10446 38872
rect 10510 38808 11310 38872
rect 11374 38808 11438 38872
rect 11502 38808 12302 38872
rect 12366 38808 12430 38872
rect 12494 38808 13294 38872
rect 13358 38808 13422 38872
rect 13486 38808 14255 38872
rect 14319 38808 14343 38872
rect 14407 38808 14431 38872
rect 14495 38808 14519 38872
rect 14583 38808 14607 38872
rect 14671 38808 15000 38872
rect 0 38792 15000 38808
rect 0 38728 462 38792
rect 526 38728 620 38792
rect 684 38728 1390 38792
rect 1454 38728 1518 38792
rect 1582 38728 2382 38792
rect 2446 38728 2510 38792
rect 2574 38728 3374 38792
rect 3438 38728 3502 38792
rect 3566 38728 4366 38792
rect 4430 38728 4494 38792
rect 4558 38728 5358 38792
rect 5422 38728 5486 38792
rect 5550 38728 6350 38792
rect 6414 38728 6478 38792
rect 6542 38728 7342 38792
rect 7406 38728 7470 38792
rect 7534 38728 8334 38792
rect 8398 38728 8462 38792
rect 8526 38728 9326 38792
rect 9390 38728 9454 38792
rect 9518 38728 10318 38792
rect 10382 38728 10446 38792
rect 10510 38728 11310 38792
rect 11374 38728 11438 38792
rect 11502 38728 12302 38792
rect 12366 38728 12430 38792
rect 12494 38728 13294 38792
rect 13358 38728 13422 38792
rect 13486 38728 14255 38792
rect 14319 38728 14343 38792
rect 14407 38728 14431 38792
rect 14495 38728 14519 38792
rect 14583 38728 14607 38792
rect 14671 38728 15000 38792
rect 0 38712 15000 38728
rect 0 38648 462 38712
rect 526 38648 620 38712
rect 684 38648 1390 38712
rect 1454 38648 1518 38712
rect 1582 38648 2382 38712
rect 2446 38648 2510 38712
rect 2574 38648 3374 38712
rect 3438 38648 3502 38712
rect 3566 38648 4366 38712
rect 4430 38648 4494 38712
rect 4558 38648 5358 38712
rect 5422 38648 5486 38712
rect 5550 38648 6350 38712
rect 6414 38648 6478 38712
rect 6542 38648 7342 38712
rect 7406 38648 7470 38712
rect 7534 38648 8334 38712
rect 8398 38648 8462 38712
rect 8526 38648 9326 38712
rect 9390 38648 9454 38712
rect 9518 38648 10318 38712
rect 10382 38648 10446 38712
rect 10510 38648 11310 38712
rect 11374 38648 11438 38712
rect 11502 38648 12302 38712
rect 12366 38648 12430 38712
rect 12494 38648 13294 38712
rect 13358 38648 13422 38712
rect 13486 38648 14255 38712
rect 14319 38648 14343 38712
rect 14407 38648 14431 38712
rect 14495 38648 14519 38712
rect 14583 38648 14607 38712
rect 14671 38648 15000 38712
rect 0 38632 15000 38648
rect 0 38568 462 38632
rect 526 38568 620 38632
rect 684 38568 1390 38632
rect 1454 38568 1518 38632
rect 1582 38568 2382 38632
rect 2446 38568 2510 38632
rect 2574 38568 3374 38632
rect 3438 38568 3502 38632
rect 3566 38568 4366 38632
rect 4430 38568 4494 38632
rect 4558 38568 5358 38632
rect 5422 38568 5486 38632
rect 5550 38568 6350 38632
rect 6414 38568 6478 38632
rect 6542 38568 7342 38632
rect 7406 38568 7470 38632
rect 7534 38568 8334 38632
rect 8398 38568 8462 38632
rect 8526 38568 9326 38632
rect 9390 38568 9454 38632
rect 9518 38568 10318 38632
rect 10382 38568 10446 38632
rect 10510 38568 11310 38632
rect 11374 38568 11438 38632
rect 11502 38568 12302 38632
rect 12366 38568 12430 38632
rect 12494 38568 13294 38632
rect 13358 38568 13422 38632
rect 13486 38568 14255 38632
rect 14319 38568 14343 38632
rect 14407 38568 14431 38632
rect 14495 38568 14519 38632
rect 14583 38568 14607 38632
rect 14671 38568 15000 38632
rect 0 38552 15000 38568
rect 0 38488 462 38552
rect 526 38488 620 38552
rect 684 38488 1390 38552
rect 1454 38488 1518 38552
rect 1582 38488 2382 38552
rect 2446 38488 2510 38552
rect 2574 38488 3374 38552
rect 3438 38488 3502 38552
rect 3566 38488 4366 38552
rect 4430 38488 4494 38552
rect 4558 38488 5358 38552
rect 5422 38488 5486 38552
rect 5550 38488 6350 38552
rect 6414 38488 6478 38552
rect 6542 38488 7342 38552
rect 7406 38488 7470 38552
rect 7534 38488 8334 38552
rect 8398 38488 8462 38552
rect 8526 38488 9326 38552
rect 9390 38488 9454 38552
rect 9518 38488 10318 38552
rect 10382 38488 10446 38552
rect 10510 38488 11310 38552
rect 11374 38488 11438 38552
rect 11502 38488 12302 38552
rect 12366 38488 12430 38552
rect 12494 38488 13294 38552
rect 13358 38488 13422 38552
rect 13486 38488 14255 38552
rect 14319 38488 14343 38552
rect 14407 38488 14431 38552
rect 14495 38488 14519 38552
rect 14583 38488 14607 38552
rect 14671 38488 15000 38552
rect 0 38472 15000 38488
rect 0 38408 462 38472
rect 526 38408 620 38472
rect 684 38408 1390 38472
rect 1454 38408 1518 38472
rect 1582 38408 2382 38472
rect 2446 38408 2510 38472
rect 2574 38408 3374 38472
rect 3438 38408 3502 38472
rect 3566 38408 4366 38472
rect 4430 38408 4494 38472
rect 4558 38408 5358 38472
rect 5422 38408 5486 38472
rect 5550 38408 6350 38472
rect 6414 38408 6478 38472
rect 6542 38408 7342 38472
rect 7406 38408 7470 38472
rect 7534 38408 8334 38472
rect 8398 38408 8462 38472
rect 8526 38408 9326 38472
rect 9390 38408 9454 38472
rect 9518 38408 10318 38472
rect 10382 38408 10446 38472
rect 10510 38408 11310 38472
rect 11374 38408 11438 38472
rect 11502 38408 12302 38472
rect 12366 38408 12430 38472
rect 12494 38408 13294 38472
rect 13358 38408 13422 38472
rect 13486 38408 14255 38472
rect 14319 38408 14343 38472
rect 14407 38408 14431 38472
rect 14495 38408 14519 38472
rect 14583 38408 14607 38472
rect 14671 38408 15000 38472
rect 0 38392 15000 38408
rect 0 38328 462 38392
rect 526 38328 620 38392
rect 684 38328 1390 38392
rect 1454 38328 1518 38392
rect 1582 38328 2382 38392
rect 2446 38328 2510 38392
rect 2574 38328 3374 38392
rect 3438 38328 3502 38392
rect 3566 38328 4366 38392
rect 4430 38328 4494 38392
rect 4558 38328 5358 38392
rect 5422 38328 5486 38392
rect 5550 38328 6350 38392
rect 6414 38328 6478 38392
rect 6542 38328 7342 38392
rect 7406 38328 7470 38392
rect 7534 38328 8334 38392
rect 8398 38328 8462 38392
rect 8526 38328 9326 38392
rect 9390 38328 9454 38392
rect 9518 38328 10318 38392
rect 10382 38328 10446 38392
rect 10510 38328 11310 38392
rect 11374 38328 11438 38392
rect 11502 38328 12302 38392
rect 12366 38328 12430 38392
rect 12494 38328 13294 38392
rect 13358 38328 13422 38392
rect 13486 38328 14255 38392
rect 14319 38328 14343 38392
rect 14407 38328 14431 38392
rect 14495 38328 14519 38392
rect 14583 38328 14607 38392
rect 14671 38328 15000 38392
rect 0 38311 15000 38328
rect 0 38247 462 38311
rect 526 38247 620 38311
rect 684 38247 1390 38311
rect 1454 38247 1518 38311
rect 1582 38247 2382 38311
rect 2446 38247 2510 38311
rect 2574 38247 3374 38311
rect 3438 38247 3502 38311
rect 3566 38247 4366 38311
rect 4430 38247 4494 38311
rect 4558 38247 5358 38311
rect 5422 38247 5486 38311
rect 5550 38247 6350 38311
rect 6414 38247 6478 38311
rect 6542 38247 7342 38311
rect 7406 38247 7470 38311
rect 7534 38247 8334 38311
rect 8398 38247 8462 38311
rect 8526 38247 9326 38311
rect 9390 38247 9454 38311
rect 9518 38247 10318 38311
rect 10382 38247 10446 38311
rect 10510 38247 11310 38311
rect 11374 38247 11438 38311
rect 11502 38247 12302 38311
rect 12366 38247 12430 38311
rect 12494 38247 13294 38311
rect 13358 38247 13422 38311
rect 13486 38247 14255 38311
rect 14319 38247 14343 38311
rect 14407 38247 14431 38311
rect 14495 38247 14519 38311
rect 14583 38247 14607 38311
rect 14671 38247 15000 38311
rect 0 38230 15000 38247
rect 0 38166 462 38230
rect 526 38166 620 38230
rect 684 38166 1390 38230
rect 1454 38166 1518 38230
rect 1582 38166 2382 38230
rect 2446 38166 2510 38230
rect 2574 38166 3374 38230
rect 3438 38166 3502 38230
rect 3566 38166 4366 38230
rect 4430 38166 4494 38230
rect 4558 38166 5358 38230
rect 5422 38166 5486 38230
rect 5550 38166 6350 38230
rect 6414 38166 6478 38230
rect 6542 38166 7342 38230
rect 7406 38166 7470 38230
rect 7534 38166 8334 38230
rect 8398 38166 8462 38230
rect 8526 38166 9326 38230
rect 9390 38166 9454 38230
rect 9518 38166 10318 38230
rect 10382 38166 10446 38230
rect 10510 38166 11310 38230
rect 11374 38166 11438 38230
rect 11502 38166 12302 38230
rect 12366 38166 12430 38230
rect 12494 38166 13294 38230
rect 13358 38166 13422 38230
rect 13486 38166 14255 38230
rect 14319 38166 14343 38230
rect 14407 38166 14431 38230
rect 14495 38166 14519 38230
rect 14583 38166 14607 38230
rect 14671 38166 15000 38230
rect 0 38149 15000 38166
rect 0 38085 462 38149
rect 526 38085 620 38149
rect 684 38085 1390 38149
rect 1454 38085 1518 38149
rect 1582 38085 2382 38149
rect 2446 38085 2510 38149
rect 2574 38085 3374 38149
rect 3438 38085 3502 38149
rect 3566 38085 4366 38149
rect 4430 38085 4494 38149
rect 4558 38085 5358 38149
rect 5422 38085 5486 38149
rect 5550 38085 6350 38149
rect 6414 38085 6478 38149
rect 6542 38085 7342 38149
rect 7406 38085 7470 38149
rect 7534 38085 8334 38149
rect 8398 38085 8462 38149
rect 8526 38085 9326 38149
rect 9390 38085 9454 38149
rect 9518 38085 10318 38149
rect 10382 38085 10446 38149
rect 10510 38085 11310 38149
rect 11374 38085 11438 38149
rect 11502 38085 12302 38149
rect 12366 38085 12430 38149
rect 12494 38085 13294 38149
rect 13358 38085 13422 38149
rect 13486 38085 14255 38149
rect 14319 38085 14343 38149
rect 14407 38085 14431 38149
rect 14495 38085 14519 38149
rect 14583 38085 14607 38149
rect 14671 38085 15000 38149
rect 0 38068 15000 38085
rect 0 38004 462 38068
rect 526 38004 620 38068
rect 684 38004 1390 38068
rect 1454 38004 1518 38068
rect 1582 38004 2382 38068
rect 2446 38004 2510 38068
rect 2574 38004 3374 38068
rect 3438 38004 3502 38068
rect 3566 38004 4366 38068
rect 4430 38004 4494 38068
rect 4558 38004 5358 38068
rect 5422 38004 5486 38068
rect 5550 38004 6350 38068
rect 6414 38004 6478 38068
rect 6542 38004 7342 38068
rect 7406 38004 7470 38068
rect 7534 38004 8334 38068
rect 8398 38004 8462 38068
rect 8526 38004 9326 38068
rect 9390 38004 9454 38068
rect 9518 38004 10318 38068
rect 10382 38004 10446 38068
rect 10510 38004 11310 38068
rect 11374 38004 11438 38068
rect 11502 38004 12302 38068
rect 12366 38004 12430 38068
rect 12494 38004 13294 38068
rect 13358 38004 13422 38068
rect 13486 38004 14255 38068
rect 14319 38004 14343 38068
rect 14407 38004 14431 38068
rect 14495 38004 14519 38068
rect 14583 38004 14607 38068
rect 14671 38004 15000 38068
rect 0 37987 15000 38004
rect 0 37923 462 37987
rect 526 37923 620 37987
rect 684 37923 1390 37987
rect 1454 37923 1518 37987
rect 1582 37923 2382 37987
rect 2446 37923 2510 37987
rect 2574 37923 3374 37987
rect 3438 37923 3502 37987
rect 3566 37923 4366 37987
rect 4430 37923 4494 37987
rect 4558 37923 5358 37987
rect 5422 37923 5486 37987
rect 5550 37923 6350 37987
rect 6414 37923 6478 37987
rect 6542 37923 7342 37987
rect 7406 37923 7470 37987
rect 7534 37923 8334 37987
rect 8398 37923 8462 37987
rect 8526 37923 9326 37987
rect 9390 37923 9454 37987
rect 9518 37923 10318 37987
rect 10382 37923 10446 37987
rect 10510 37923 11310 37987
rect 11374 37923 11438 37987
rect 11502 37923 12302 37987
rect 12366 37923 12430 37987
rect 12494 37923 13294 37987
rect 13358 37923 13422 37987
rect 13486 37923 14255 37987
rect 14319 37923 14343 37987
rect 14407 37923 14431 37987
rect 14495 37923 14519 37987
rect 14583 37923 14607 37987
rect 14671 37923 15000 37987
rect 0 37906 15000 37923
rect 0 37842 462 37906
rect 526 37842 620 37906
rect 684 37842 1390 37906
rect 1454 37842 1518 37906
rect 1582 37842 2382 37906
rect 2446 37842 2510 37906
rect 2574 37842 3374 37906
rect 3438 37842 3502 37906
rect 3566 37842 4366 37906
rect 4430 37842 4494 37906
rect 4558 37842 5358 37906
rect 5422 37842 5486 37906
rect 5550 37842 6350 37906
rect 6414 37842 6478 37906
rect 6542 37842 7342 37906
rect 7406 37842 7470 37906
rect 7534 37842 8334 37906
rect 8398 37842 8462 37906
rect 8526 37842 9326 37906
rect 9390 37842 9454 37906
rect 9518 37842 10318 37906
rect 10382 37842 10446 37906
rect 10510 37842 11310 37906
rect 11374 37842 11438 37906
rect 11502 37842 12302 37906
rect 12366 37842 12430 37906
rect 12494 37842 13294 37906
rect 13358 37842 13422 37906
rect 13486 37842 14255 37906
rect 14319 37842 14343 37906
rect 14407 37842 14431 37906
rect 14495 37842 14519 37906
rect 14583 37842 14607 37906
rect 14671 37842 15000 37906
rect 0 37825 15000 37842
rect 0 37761 462 37825
rect 526 37761 620 37825
rect 684 37761 1390 37825
rect 1454 37761 1518 37825
rect 1582 37761 2382 37825
rect 2446 37761 2510 37825
rect 2574 37761 3374 37825
rect 3438 37761 3502 37825
rect 3566 37761 4366 37825
rect 4430 37761 4494 37825
rect 4558 37761 5358 37825
rect 5422 37761 5486 37825
rect 5550 37761 6350 37825
rect 6414 37761 6478 37825
rect 6542 37761 7342 37825
rect 7406 37761 7470 37825
rect 7534 37761 8334 37825
rect 8398 37761 8462 37825
rect 8526 37761 9326 37825
rect 9390 37761 9454 37825
rect 9518 37761 10318 37825
rect 10382 37761 10446 37825
rect 10510 37761 11310 37825
rect 11374 37761 11438 37825
rect 11502 37761 12302 37825
rect 12366 37761 12430 37825
rect 12494 37761 13294 37825
rect 13358 37761 13422 37825
rect 13486 37761 14255 37825
rect 14319 37761 14343 37825
rect 14407 37761 14431 37825
rect 14495 37761 14519 37825
rect 14583 37761 14607 37825
rect 14671 37761 15000 37825
rect 0 37744 15000 37761
rect 0 37680 462 37744
rect 526 37680 620 37744
rect 684 37680 1390 37744
rect 1454 37680 1518 37744
rect 1582 37680 2382 37744
rect 2446 37680 2510 37744
rect 2574 37680 3374 37744
rect 3438 37680 3502 37744
rect 3566 37680 4366 37744
rect 4430 37680 4494 37744
rect 4558 37680 5358 37744
rect 5422 37680 5486 37744
rect 5550 37680 6350 37744
rect 6414 37680 6478 37744
rect 6542 37680 7342 37744
rect 7406 37680 7470 37744
rect 7534 37680 8334 37744
rect 8398 37680 8462 37744
rect 8526 37680 9326 37744
rect 9390 37680 9454 37744
rect 9518 37680 10318 37744
rect 10382 37680 10446 37744
rect 10510 37680 11310 37744
rect 11374 37680 11438 37744
rect 11502 37680 12302 37744
rect 12366 37680 12430 37744
rect 12494 37680 13294 37744
rect 13358 37680 13422 37744
rect 13486 37680 14255 37744
rect 14319 37680 14343 37744
rect 14407 37680 14431 37744
rect 14495 37680 14519 37744
rect 14583 37680 14607 37744
rect 14671 37680 15000 37744
rect 0 37663 15000 37680
rect 0 37599 462 37663
rect 526 37599 620 37663
rect 684 37599 1390 37663
rect 1454 37599 1518 37663
rect 1582 37599 2382 37663
rect 2446 37599 2510 37663
rect 2574 37599 3374 37663
rect 3438 37599 3502 37663
rect 3566 37599 4366 37663
rect 4430 37599 4494 37663
rect 4558 37599 5358 37663
rect 5422 37599 5486 37663
rect 5550 37599 6350 37663
rect 6414 37599 6478 37663
rect 6542 37599 7342 37663
rect 7406 37599 7470 37663
rect 7534 37599 8334 37663
rect 8398 37599 8462 37663
rect 8526 37599 9326 37663
rect 9390 37599 9454 37663
rect 9518 37599 10318 37663
rect 10382 37599 10446 37663
rect 10510 37599 11310 37663
rect 11374 37599 11438 37663
rect 11502 37599 12302 37663
rect 12366 37599 12430 37663
rect 12494 37599 13294 37663
rect 13358 37599 13422 37663
rect 13486 37599 14255 37663
rect 14319 37599 14343 37663
rect 14407 37599 14431 37663
rect 14495 37599 14519 37663
rect 14583 37599 14607 37663
rect 14671 37599 15000 37663
rect 0 37582 15000 37599
rect 0 37518 462 37582
rect 526 37518 620 37582
rect 684 37518 1390 37582
rect 1454 37518 1518 37582
rect 1582 37518 2382 37582
rect 2446 37518 2510 37582
rect 2574 37518 3374 37582
rect 3438 37518 3502 37582
rect 3566 37518 4366 37582
rect 4430 37518 4494 37582
rect 4558 37518 5358 37582
rect 5422 37518 5486 37582
rect 5550 37518 6350 37582
rect 6414 37518 6478 37582
rect 6542 37518 7342 37582
rect 7406 37518 7470 37582
rect 7534 37518 8334 37582
rect 8398 37518 8462 37582
rect 8526 37518 9326 37582
rect 9390 37518 9454 37582
rect 9518 37518 10318 37582
rect 10382 37518 10446 37582
rect 10510 37518 11310 37582
rect 11374 37518 11438 37582
rect 11502 37518 12302 37582
rect 12366 37518 12430 37582
rect 12494 37518 13294 37582
rect 13358 37518 13422 37582
rect 13486 37518 14255 37582
rect 14319 37518 14343 37582
rect 14407 37518 14431 37582
rect 14495 37518 14519 37582
rect 14583 37518 14607 37582
rect 14671 37518 15000 37582
rect 0 37501 15000 37518
rect 0 37437 462 37501
rect 526 37437 620 37501
rect 684 37437 1390 37501
rect 1454 37437 1518 37501
rect 1582 37437 2382 37501
rect 2446 37437 2510 37501
rect 2574 37437 3374 37501
rect 3438 37437 3502 37501
rect 3566 37437 4366 37501
rect 4430 37437 4494 37501
rect 4558 37437 5358 37501
rect 5422 37437 5486 37501
rect 5550 37437 6350 37501
rect 6414 37437 6478 37501
rect 6542 37437 7342 37501
rect 7406 37437 7470 37501
rect 7534 37437 8334 37501
rect 8398 37437 8462 37501
rect 8526 37437 9326 37501
rect 9390 37437 9454 37501
rect 9518 37437 10318 37501
rect 10382 37437 10446 37501
rect 10510 37437 11310 37501
rect 11374 37437 11438 37501
rect 11502 37437 12302 37501
rect 12366 37437 12430 37501
rect 12494 37437 13294 37501
rect 13358 37437 13422 37501
rect 13486 37437 14255 37501
rect 14319 37437 14343 37501
rect 14407 37437 14431 37501
rect 14495 37437 14519 37501
rect 14583 37437 14607 37501
rect 14671 37437 15000 37501
rect 0 37420 15000 37437
rect 0 37356 462 37420
rect 526 37356 620 37420
rect 684 37356 1390 37420
rect 1454 37356 1518 37420
rect 1582 37356 2382 37420
rect 2446 37356 2510 37420
rect 2574 37356 3374 37420
rect 3438 37356 3502 37420
rect 3566 37356 4366 37420
rect 4430 37356 4494 37420
rect 4558 37356 5358 37420
rect 5422 37356 5486 37420
rect 5550 37356 6350 37420
rect 6414 37356 6478 37420
rect 6542 37356 7342 37420
rect 7406 37356 7470 37420
rect 7534 37356 8334 37420
rect 8398 37356 8462 37420
rect 8526 37356 9326 37420
rect 9390 37356 9454 37420
rect 9518 37356 10318 37420
rect 10382 37356 10446 37420
rect 10510 37356 11310 37420
rect 11374 37356 11438 37420
rect 11502 37356 12302 37420
rect 12366 37356 12430 37420
rect 12494 37356 13294 37420
rect 13358 37356 13422 37420
rect 13486 37356 14255 37420
rect 14319 37356 14343 37420
rect 14407 37356 14431 37420
rect 14495 37356 14519 37420
rect 14583 37356 14607 37420
rect 14671 37356 15000 37420
rect 0 37339 15000 37356
rect 0 37275 462 37339
rect 526 37275 620 37339
rect 684 37275 1390 37339
rect 1454 37275 1518 37339
rect 1582 37275 2382 37339
rect 2446 37275 2510 37339
rect 2574 37275 3374 37339
rect 3438 37275 3502 37339
rect 3566 37275 4366 37339
rect 4430 37275 4494 37339
rect 4558 37275 5358 37339
rect 5422 37275 5486 37339
rect 5550 37275 6350 37339
rect 6414 37275 6478 37339
rect 6542 37275 7342 37339
rect 7406 37275 7470 37339
rect 7534 37275 8334 37339
rect 8398 37275 8462 37339
rect 8526 37275 9326 37339
rect 9390 37275 9454 37339
rect 9518 37275 10318 37339
rect 10382 37275 10446 37339
rect 10510 37275 11310 37339
rect 11374 37275 11438 37339
rect 11502 37275 12302 37339
rect 12366 37275 12430 37339
rect 12494 37275 13294 37339
rect 13358 37275 13422 37339
rect 13486 37275 14255 37339
rect 14319 37275 14343 37339
rect 14407 37275 14431 37339
rect 14495 37275 14519 37339
rect 14583 37275 14607 37339
rect 14671 37275 15000 37339
rect 0 37258 15000 37275
rect 0 37194 462 37258
rect 526 37194 620 37258
rect 684 37194 1390 37258
rect 1454 37194 1518 37258
rect 1582 37194 2382 37258
rect 2446 37194 2510 37258
rect 2574 37194 3374 37258
rect 3438 37194 3502 37258
rect 3566 37194 4366 37258
rect 4430 37194 4494 37258
rect 4558 37194 5358 37258
rect 5422 37194 5486 37258
rect 5550 37194 6350 37258
rect 6414 37194 6478 37258
rect 6542 37194 7342 37258
rect 7406 37194 7470 37258
rect 7534 37194 8334 37258
rect 8398 37194 8462 37258
rect 8526 37194 9326 37258
rect 9390 37194 9454 37258
rect 9518 37194 10318 37258
rect 10382 37194 10446 37258
rect 10510 37194 11310 37258
rect 11374 37194 11438 37258
rect 11502 37194 12302 37258
rect 12366 37194 12430 37258
rect 12494 37194 13294 37258
rect 13358 37194 13422 37258
rect 13486 37194 14255 37258
rect 14319 37194 14343 37258
rect 14407 37194 14431 37258
rect 14495 37194 14519 37258
rect 14583 37194 14607 37258
rect 14671 37194 15000 37258
rect 0 37177 15000 37194
rect 0 37113 462 37177
rect 526 37113 620 37177
rect 684 37113 1390 37177
rect 1454 37113 1518 37177
rect 1582 37113 2382 37177
rect 2446 37113 2510 37177
rect 2574 37113 3374 37177
rect 3438 37113 3502 37177
rect 3566 37113 4366 37177
rect 4430 37113 4494 37177
rect 4558 37113 5358 37177
rect 5422 37113 5486 37177
rect 5550 37113 6350 37177
rect 6414 37113 6478 37177
rect 6542 37113 7342 37177
rect 7406 37113 7470 37177
rect 7534 37113 8334 37177
rect 8398 37113 8462 37177
rect 8526 37113 9326 37177
rect 9390 37113 9454 37177
rect 9518 37113 10318 37177
rect 10382 37113 10446 37177
rect 10510 37113 11310 37177
rect 11374 37113 11438 37177
rect 11502 37113 12302 37177
rect 12366 37113 12430 37177
rect 12494 37113 13294 37177
rect 13358 37113 13422 37177
rect 13486 37113 14255 37177
rect 14319 37113 14343 37177
rect 14407 37113 14431 37177
rect 14495 37113 14519 37177
rect 14583 37113 14607 37177
rect 14671 37113 15000 37177
rect 0 37096 15000 37113
rect 0 37032 462 37096
rect 526 37032 620 37096
rect 684 37032 1390 37096
rect 1454 37032 1518 37096
rect 1582 37032 2382 37096
rect 2446 37032 2510 37096
rect 2574 37032 3374 37096
rect 3438 37032 3502 37096
rect 3566 37032 4366 37096
rect 4430 37032 4494 37096
rect 4558 37032 5358 37096
rect 5422 37032 5486 37096
rect 5550 37032 6350 37096
rect 6414 37032 6478 37096
rect 6542 37032 7342 37096
rect 7406 37032 7470 37096
rect 7534 37032 8334 37096
rect 8398 37032 8462 37096
rect 8526 37032 9326 37096
rect 9390 37032 9454 37096
rect 9518 37032 10318 37096
rect 10382 37032 10446 37096
rect 10510 37032 11310 37096
rect 11374 37032 11438 37096
rect 11502 37032 12302 37096
rect 12366 37032 12430 37096
rect 12494 37032 13294 37096
rect 13358 37032 13422 37096
rect 13486 37032 14255 37096
rect 14319 37032 14343 37096
rect 14407 37032 14431 37096
rect 14495 37032 14519 37096
rect 14583 37032 14607 37096
rect 14671 37032 15000 37096
rect 0 37015 15000 37032
rect 0 36951 462 37015
rect 526 36951 620 37015
rect 684 36951 1390 37015
rect 1454 36951 1518 37015
rect 1582 36951 2382 37015
rect 2446 36951 2510 37015
rect 2574 36951 3374 37015
rect 3438 36951 3502 37015
rect 3566 36951 4366 37015
rect 4430 36951 4494 37015
rect 4558 36951 5358 37015
rect 5422 36951 5486 37015
rect 5550 36951 6350 37015
rect 6414 36951 6478 37015
rect 6542 36951 7342 37015
rect 7406 36951 7470 37015
rect 7534 36951 8334 37015
rect 8398 36951 8462 37015
rect 8526 36951 9326 37015
rect 9390 36951 9454 37015
rect 9518 36951 10318 37015
rect 10382 36951 10446 37015
rect 10510 36951 11310 37015
rect 11374 36951 11438 37015
rect 11502 36951 12302 37015
rect 12366 36951 12430 37015
rect 12494 36951 13294 37015
rect 13358 36951 13422 37015
rect 13486 36951 14255 37015
rect 14319 36951 14343 37015
rect 14407 36951 14431 37015
rect 14495 36951 14519 37015
rect 14583 36951 14607 37015
rect 14671 36951 15000 37015
rect 0 36934 15000 36951
rect 0 36870 462 36934
rect 526 36870 620 36934
rect 684 36870 1390 36934
rect 1454 36870 1518 36934
rect 1582 36870 2382 36934
rect 2446 36870 2510 36934
rect 2574 36870 3374 36934
rect 3438 36870 3502 36934
rect 3566 36870 4366 36934
rect 4430 36870 4494 36934
rect 4558 36870 5358 36934
rect 5422 36870 5486 36934
rect 5550 36870 6350 36934
rect 6414 36870 6478 36934
rect 6542 36870 7342 36934
rect 7406 36870 7470 36934
rect 7534 36870 8334 36934
rect 8398 36870 8462 36934
rect 8526 36870 9326 36934
rect 9390 36870 9454 36934
rect 9518 36870 10318 36934
rect 10382 36870 10446 36934
rect 10510 36870 11310 36934
rect 11374 36870 11438 36934
rect 11502 36870 12302 36934
rect 12366 36870 12430 36934
rect 12494 36870 13294 36934
rect 13358 36870 13422 36934
rect 13486 36870 14255 36934
rect 14319 36870 14343 36934
rect 14407 36870 14431 36934
rect 14495 36870 14519 36934
rect 14583 36870 14607 36934
rect 14671 36870 15000 36934
rect 0 36853 15000 36870
rect 0 36789 462 36853
rect 526 36789 620 36853
rect 684 36789 1390 36853
rect 1454 36789 1518 36853
rect 1582 36789 2382 36853
rect 2446 36789 2510 36853
rect 2574 36789 3374 36853
rect 3438 36789 3502 36853
rect 3566 36789 4366 36853
rect 4430 36789 4494 36853
rect 4558 36789 5358 36853
rect 5422 36789 5486 36853
rect 5550 36789 6350 36853
rect 6414 36789 6478 36853
rect 6542 36789 7342 36853
rect 7406 36789 7470 36853
rect 7534 36789 8334 36853
rect 8398 36789 8462 36853
rect 8526 36789 9326 36853
rect 9390 36789 9454 36853
rect 9518 36789 10318 36853
rect 10382 36789 10446 36853
rect 10510 36789 11310 36853
rect 11374 36789 11438 36853
rect 11502 36789 12302 36853
rect 12366 36789 12430 36853
rect 12494 36789 13294 36853
rect 13358 36789 13422 36853
rect 13486 36789 14255 36853
rect 14319 36789 14343 36853
rect 14407 36789 14431 36853
rect 14495 36789 14519 36853
rect 14583 36789 14607 36853
rect 14671 36789 15000 36853
rect 0 36772 15000 36789
rect 0 36708 462 36772
rect 526 36708 620 36772
rect 684 36708 1390 36772
rect 1454 36708 1518 36772
rect 1582 36708 2382 36772
rect 2446 36708 2510 36772
rect 2574 36708 3374 36772
rect 3438 36708 3502 36772
rect 3566 36708 4366 36772
rect 4430 36708 4494 36772
rect 4558 36708 5358 36772
rect 5422 36708 5486 36772
rect 5550 36708 6350 36772
rect 6414 36708 6478 36772
rect 6542 36708 7342 36772
rect 7406 36708 7470 36772
rect 7534 36708 8334 36772
rect 8398 36708 8462 36772
rect 8526 36708 9326 36772
rect 9390 36708 9454 36772
rect 9518 36708 10318 36772
rect 10382 36708 10446 36772
rect 10510 36708 11310 36772
rect 11374 36708 11438 36772
rect 11502 36708 12302 36772
rect 12366 36708 12430 36772
rect 12494 36708 13294 36772
rect 13358 36708 13422 36772
rect 13486 36708 14255 36772
rect 14319 36708 14343 36772
rect 14407 36708 14431 36772
rect 14495 36708 14519 36772
rect 14583 36708 14607 36772
rect 14671 36708 15000 36772
rect 0 36691 15000 36708
rect 0 36627 462 36691
rect 526 36627 620 36691
rect 684 36627 1390 36691
rect 1454 36627 1518 36691
rect 1582 36627 2382 36691
rect 2446 36627 2510 36691
rect 2574 36627 3374 36691
rect 3438 36627 3502 36691
rect 3566 36627 4366 36691
rect 4430 36627 4494 36691
rect 4558 36627 5358 36691
rect 5422 36627 5486 36691
rect 5550 36627 6350 36691
rect 6414 36627 6478 36691
rect 6542 36627 7342 36691
rect 7406 36627 7470 36691
rect 7534 36627 8334 36691
rect 8398 36627 8462 36691
rect 8526 36627 9326 36691
rect 9390 36627 9454 36691
rect 9518 36627 10318 36691
rect 10382 36627 10446 36691
rect 10510 36627 11310 36691
rect 11374 36627 11438 36691
rect 11502 36627 12302 36691
rect 12366 36627 12430 36691
rect 12494 36627 13294 36691
rect 13358 36627 13422 36691
rect 13486 36627 14255 36691
rect 14319 36627 14343 36691
rect 14407 36627 14431 36691
rect 14495 36627 14519 36691
rect 14583 36627 14607 36691
rect 14671 36627 15000 36691
rect 0 36610 15000 36627
rect 0 36546 462 36610
rect 526 36546 620 36610
rect 684 36546 1390 36610
rect 1454 36546 1518 36610
rect 1582 36546 2382 36610
rect 2446 36546 2510 36610
rect 2574 36546 3374 36610
rect 3438 36546 3502 36610
rect 3566 36546 4366 36610
rect 4430 36546 4494 36610
rect 4558 36546 5358 36610
rect 5422 36546 5486 36610
rect 5550 36546 6350 36610
rect 6414 36546 6478 36610
rect 6542 36546 7342 36610
rect 7406 36546 7470 36610
rect 7534 36546 8334 36610
rect 8398 36546 8462 36610
rect 8526 36546 9326 36610
rect 9390 36546 9454 36610
rect 9518 36546 10318 36610
rect 10382 36546 10446 36610
rect 10510 36546 11310 36610
rect 11374 36546 11438 36610
rect 11502 36546 12302 36610
rect 12366 36546 12430 36610
rect 12494 36546 13294 36610
rect 13358 36546 13422 36610
rect 13486 36546 14255 36610
rect 14319 36546 14343 36610
rect 14407 36546 14431 36610
rect 14495 36546 14519 36610
rect 14583 36546 14607 36610
rect 14671 36546 15000 36610
rect 0 36529 15000 36546
rect 0 36465 462 36529
rect 526 36465 620 36529
rect 684 36465 1390 36529
rect 1454 36465 1518 36529
rect 1582 36465 2382 36529
rect 2446 36465 2510 36529
rect 2574 36465 3374 36529
rect 3438 36465 3502 36529
rect 3566 36465 4366 36529
rect 4430 36465 4494 36529
rect 4558 36465 5358 36529
rect 5422 36465 5486 36529
rect 5550 36465 6350 36529
rect 6414 36465 6478 36529
rect 6542 36465 7342 36529
rect 7406 36465 7470 36529
rect 7534 36465 8334 36529
rect 8398 36465 8462 36529
rect 8526 36465 9326 36529
rect 9390 36465 9454 36529
rect 9518 36465 10318 36529
rect 10382 36465 10446 36529
rect 10510 36465 11310 36529
rect 11374 36465 11438 36529
rect 11502 36465 12302 36529
rect 12366 36465 12430 36529
rect 12494 36465 13294 36529
rect 13358 36465 13422 36529
rect 13486 36465 14255 36529
rect 14319 36465 14343 36529
rect 14407 36465 14431 36529
rect 14495 36465 14519 36529
rect 14583 36465 14607 36529
rect 14671 36465 15000 36529
rect 0 36448 15000 36465
rect 0 36384 462 36448
rect 526 36384 620 36448
rect 684 36384 1390 36448
rect 1454 36384 1518 36448
rect 1582 36384 2382 36448
rect 2446 36384 2510 36448
rect 2574 36384 3374 36448
rect 3438 36384 3502 36448
rect 3566 36384 4366 36448
rect 4430 36384 4494 36448
rect 4558 36384 5358 36448
rect 5422 36384 5486 36448
rect 5550 36384 6350 36448
rect 6414 36384 6478 36448
rect 6542 36384 7342 36448
rect 7406 36384 7470 36448
rect 7534 36384 8334 36448
rect 8398 36384 8462 36448
rect 8526 36384 9326 36448
rect 9390 36384 9454 36448
rect 9518 36384 10318 36448
rect 10382 36384 10446 36448
rect 10510 36384 11310 36448
rect 11374 36384 11438 36448
rect 11502 36384 12302 36448
rect 12366 36384 12430 36448
rect 12494 36384 13294 36448
rect 13358 36384 13422 36448
rect 13486 36384 14255 36448
rect 14319 36384 14343 36448
rect 14407 36384 14431 36448
rect 14495 36384 14519 36448
rect 14583 36384 14607 36448
rect 14671 36384 15000 36448
rect 0 36367 15000 36384
rect 0 36303 462 36367
rect 526 36303 620 36367
rect 684 36303 1390 36367
rect 1454 36303 1518 36367
rect 1582 36303 2382 36367
rect 2446 36303 2510 36367
rect 2574 36303 3374 36367
rect 3438 36303 3502 36367
rect 3566 36303 4366 36367
rect 4430 36303 4494 36367
rect 4558 36303 5358 36367
rect 5422 36303 5486 36367
rect 5550 36303 6350 36367
rect 6414 36303 6478 36367
rect 6542 36303 7342 36367
rect 7406 36303 7470 36367
rect 7534 36303 8334 36367
rect 8398 36303 8462 36367
rect 8526 36303 9326 36367
rect 9390 36303 9454 36367
rect 9518 36303 10318 36367
rect 10382 36303 10446 36367
rect 10510 36303 11310 36367
rect 11374 36303 11438 36367
rect 11502 36303 12302 36367
rect 12366 36303 12430 36367
rect 12494 36303 13294 36367
rect 13358 36303 13422 36367
rect 13486 36303 14255 36367
rect 14319 36303 14343 36367
rect 14407 36303 14431 36367
rect 14495 36303 14519 36367
rect 14583 36303 14607 36367
rect 14671 36303 15000 36367
rect 0 36286 15000 36303
rect 0 36222 462 36286
rect 526 36222 620 36286
rect 684 36222 1390 36286
rect 1454 36222 1518 36286
rect 1582 36222 2382 36286
rect 2446 36222 2510 36286
rect 2574 36222 3374 36286
rect 3438 36222 3502 36286
rect 3566 36222 4366 36286
rect 4430 36222 4494 36286
rect 4558 36222 5358 36286
rect 5422 36222 5486 36286
rect 5550 36222 6350 36286
rect 6414 36222 6478 36286
rect 6542 36222 7342 36286
rect 7406 36222 7470 36286
rect 7534 36222 8334 36286
rect 8398 36222 8462 36286
rect 8526 36222 9326 36286
rect 9390 36222 9454 36286
rect 9518 36222 10318 36286
rect 10382 36222 10446 36286
rect 10510 36222 11310 36286
rect 11374 36222 11438 36286
rect 11502 36222 12302 36286
rect 12366 36222 12430 36286
rect 12494 36222 13294 36286
rect 13358 36222 13422 36286
rect 13486 36222 14255 36286
rect 14319 36222 14343 36286
rect 14407 36222 14431 36286
rect 14495 36222 14519 36286
rect 14583 36222 14607 36286
rect 14671 36222 15000 36286
rect 0 36205 15000 36222
rect 0 36141 462 36205
rect 526 36141 620 36205
rect 684 36141 1390 36205
rect 1454 36141 1518 36205
rect 1582 36141 2382 36205
rect 2446 36141 2510 36205
rect 2574 36141 3374 36205
rect 3438 36141 3502 36205
rect 3566 36141 4366 36205
rect 4430 36141 4494 36205
rect 4558 36141 5358 36205
rect 5422 36141 5486 36205
rect 5550 36141 6350 36205
rect 6414 36141 6478 36205
rect 6542 36141 7342 36205
rect 7406 36141 7470 36205
rect 7534 36141 8334 36205
rect 8398 36141 8462 36205
rect 8526 36141 9326 36205
rect 9390 36141 9454 36205
rect 9518 36141 10318 36205
rect 10382 36141 10446 36205
rect 10510 36141 11310 36205
rect 11374 36141 11438 36205
rect 11502 36141 12302 36205
rect 12366 36141 12430 36205
rect 12494 36141 13294 36205
rect 13358 36141 13422 36205
rect 13486 36141 14255 36205
rect 14319 36141 14343 36205
rect 14407 36141 14431 36205
rect 14495 36141 14519 36205
rect 14583 36141 14607 36205
rect 14671 36141 15000 36205
rect 0 36124 15000 36141
rect 0 36060 462 36124
rect 526 36060 620 36124
rect 684 36060 1390 36124
rect 1454 36060 1518 36124
rect 1582 36060 2382 36124
rect 2446 36060 2510 36124
rect 2574 36060 3374 36124
rect 3438 36060 3502 36124
rect 3566 36060 4366 36124
rect 4430 36060 4494 36124
rect 4558 36060 5358 36124
rect 5422 36060 5486 36124
rect 5550 36060 6350 36124
rect 6414 36060 6478 36124
rect 6542 36060 7342 36124
rect 7406 36060 7470 36124
rect 7534 36060 8334 36124
rect 8398 36060 8462 36124
rect 8526 36060 9326 36124
rect 9390 36060 9454 36124
rect 9518 36060 10318 36124
rect 10382 36060 10446 36124
rect 10510 36060 11310 36124
rect 11374 36060 11438 36124
rect 11502 36060 12302 36124
rect 12366 36060 12430 36124
rect 12494 36060 13294 36124
rect 13358 36060 13422 36124
rect 13486 36060 14255 36124
rect 14319 36060 14343 36124
rect 14407 36060 14431 36124
rect 14495 36060 14519 36124
rect 14583 36060 14607 36124
rect 14671 36060 15000 36124
rect 0 36043 15000 36060
rect 0 35979 462 36043
rect 526 35979 620 36043
rect 684 35979 1390 36043
rect 1454 35979 1518 36043
rect 1582 35979 2382 36043
rect 2446 35979 2510 36043
rect 2574 35979 3374 36043
rect 3438 35979 3502 36043
rect 3566 35979 4366 36043
rect 4430 35979 4494 36043
rect 4558 35979 5358 36043
rect 5422 35979 5486 36043
rect 5550 35979 6350 36043
rect 6414 35979 6478 36043
rect 6542 35979 7342 36043
rect 7406 35979 7470 36043
rect 7534 35979 8334 36043
rect 8398 35979 8462 36043
rect 8526 35979 9326 36043
rect 9390 35979 9454 36043
rect 9518 35979 10318 36043
rect 10382 35979 10446 36043
rect 10510 35979 11310 36043
rect 11374 35979 11438 36043
rect 11502 35979 12302 36043
rect 12366 35979 12430 36043
rect 12494 35979 13294 36043
rect 13358 35979 13422 36043
rect 13486 35979 14255 36043
rect 14319 35979 14343 36043
rect 14407 35979 14431 36043
rect 14495 35979 14519 36043
rect 14583 35979 14607 36043
rect 14671 35979 15000 36043
rect 0 35962 15000 35979
rect 0 35898 462 35962
rect 526 35898 620 35962
rect 684 35898 1390 35962
rect 1454 35898 1518 35962
rect 1582 35898 2382 35962
rect 2446 35898 2510 35962
rect 2574 35898 3374 35962
rect 3438 35898 3502 35962
rect 3566 35898 4366 35962
rect 4430 35898 4494 35962
rect 4558 35898 5358 35962
rect 5422 35898 5486 35962
rect 5550 35898 6350 35962
rect 6414 35898 6478 35962
rect 6542 35898 7342 35962
rect 7406 35898 7470 35962
rect 7534 35898 8334 35962
rect 8398 35898 8462 35962
rect 8526 35898 9326 35962
rect 9390 35898 9454 35962
rect 9518 35898 10318 35962
rect 10382 35898 10446 35962
rect 10510 35898 11310 35962
rect 11374 35898 11438 35962
rect 11502 35898 12302 35962
rect 12366 35898 12430 35962
rect 12494 35898 13294 35962
rect 13358 35898 13422 35962
rect 13486 35898 14255 35962
rect 14319 35898 14343 35962
rect 14407 35898 14431 35962
rect 14495 35898 14519 35962
rect 14583 35898 14607 35962
rect 14671 35898 15000 35962
rect 0 35881 15000 35898
rect 0 35817 462 35881
rect 526 35817 620 35881
rect 684 35817 1390 35881
rect 1454 35817 1518 35881
rect 1582 35817 2382 35881
rect 2446 35817 2510 35881
rect 2574 35817 3374 35881
rect 3438 35817 3502 35881
rect 3566 35817 4366 35881
rect 4430 35817 4494 35881
rect 4558 35817 5358 35881
rect 5422 35817 5486 35881
rect 5550 35817 6350 35881
rect 6414 35817 6478 35881
rect 6542 35817 7342 35881
rect 7406 35817 7470 35881
rect 7534 35817 8334 35881
rect 8398 35817 8462 35881
rect 8526 35817 9326 35881
rect 9390 35817 9454 35881
rect 9518 35817 10318 35881
rect 10382 35817 10446 35881
rect 10510 35817 11310 35881
rect 11374 35817 11438 35881
rect 11502 35817 12302 35881
rect 12366 35817 12430 35881
rect 12494 35817 13294 35881
rect 13358 35817 13422 35881
rect 13486 35817 14255 35881
rect 14319 35817 14343 35881
rect 14407 35817 14431 35881
rect 14495 35817 14519 35881
rect 14583 35817 14607 35881
rect 14671 35817 15000 35881
rect 0 35800 15000 35817
rect 0 35736 462 35800
rect 526 35736 620 35800
rect 684 35736 1390 35800
rect 1454 35736 1518 35800
rect 1582 35736 2382 35800
rect 2446 35736 2510 35800
rect 2574 35736 3374 35800
rect 3438 35736 3502 35800
rect 3566 35736 4366 35800
rect 4430 35736 4494 35800
rect 4558 35736 5358 35800
rect 5422 35736 5486 35800
rect 5550 35736 6350 35800
rect 6414 35736 6478 35800
rect 6542 35736 7342 35800
rect 7406 35736 7470 35800
rect 7534 35736 8334 35800
rect 8398 35736 8462 35800
rect 8526 35736 9326 35800
rect 9390 35736 9454 35800
rect 9518 35736 10318 35800
rect 10382 35736 10446 35800
rect 10510 35736 11310 35800
rect 11374 35736 11438 35800
rect 11502 35736 12302 35800
rect 12366 35736 12430 35800
rect 12494 35736 13294 35800
rect 13358 35736 13422 35800
rect 13486 35736 14255 35800
rect 14319 35736 14343 35800
rect 14407 35736 14431 35800
rect 14495 35736 14519 35800
rect 14583 35736 14607 35800
rect 14671 35736 15000 35800
rect 0 35719 15000 35736
rect 0 35655 462 35719
rect 526 35655 620 35719
rect 684 35655 1390 35719
rect 1454 35655 1518 35719
rect 1582 35655 2382 35719
rect 2446 35655 2510 35719
rect 2574 35655 3374 35719
rect 3438 35655 3502 35719
rect 3566 35655 4366 35719
rect 4430 35655 4494 35719
rect 4558 35655 5358 35719
rect 5422 35655 5486 35719
rect 5550 35655 6350 35719
rect 6414 35655 6478 35719
rect 6542 35655 7342 35719
rect 7406 35655 7470 35719
rect 7534 35655 8334 35719
rect 8398 35655 8462 35719
rect 8526 35655 9326 35719
rect 9390 35655 9454 35719
rect 9518 35655 10318 35719
rect 10382 35655 10446 35719
rect 10510 35655 11310 35719
rect 11374 35655 11438 35719
rect 11502 35655 12302 35719
rect 12366 35655 12430 35719
rect 12494 35655 13294 35719
rect 13358 35655 13422 35719
rect 13486 35655 14255 35719
rect 14319 35655 14343 35719
rect 14407 35655 14431 35719
rect 14495 35655 14519 35719
rect 14583 35655 14607 35719
rect 14671 35655 15000 35719
rect 0 35638 15000 35655
rect 0 35574 462 35638
rect 526 35574 620 35638
rect 684 35574 1390 35638
rect 1454 35574 1518 35638
rect 1582 35574 2382 35638
rect 2446 35574 2510 35638
rect 2574 35574 3374 35638
rect 3438 35574 3502 35638
rect 3566 35574 4366 35638
rect 4430 35574 4494 35638
rect 4558 35574 5358 35638
rect 5422 35574 5486 35638
rect 5550 35574 6350 35638
rect 6414 35574 6478 35638
rect 6542 35574 7342 35638
rect 7406 35574 7470 35638
rect 7534 35574 8334 35638
rect 8398 35574 8462 35638
rect 8526 35574 9326 35638
rect 9390 35574 9454 35638
rect 9518 35574 10318 35638
rect 10382 35574 10446 35638
rect 10510 35574 11310 35638
rect 11374 35574 11438 35638
rect 11502 35574 12302 35638
rect 12366 35574 12430 35638
rect 12494 35574 13294 35638
rect 13358 35574 13422 35638
rect 13486 35574 14255 35638
rect 14319 35574 14343 35638
rect 14407 35574 14431 35638
rect 14495 35574 14519 35638
rect 14583 35574 14607 35638
rect 14671 35574 15000 35638
rect 0 35557 15000 35574
rect 0 35493 462 35557
rect 526 35493 620 35557
rect 684 35493 1390 35557
rect 1454 35493 1518 35557
rect 1582 35493 2382 35557
rect 2446 35493 2510 35557
rect 2574 35493 3374 35557
rect 3438 35493 3502 35557
rect 3566 35493 4366 35557
rect 4430 35493 4494 35557
rect 4558 35493 5358 35557
rect 5422 35493 5486 35557
rect 5550 35493 6350 35557
rect 6414 35493 6478 35557
rect 6542 35493 7342 35557
rect 7406 35493 7470 35557
rect 7534 35493 8334 35557
rect 8398 35493 8462 35557
rect 8526 35493 9326 35557
rect 9390 35493 9454 35557
rect 9518 35493 10318 35557
rect 10382 35493 10446 35557
rect 10510 35493 11310 35557
rect 11374 35493 11438 35557
rect 11502 35493 12302 35557
rect 12366 35493 12430 35557
rect 12494 35493 13294 35557
rect 13358 35493 13422 35557
rect 13486 35493 14255 35557
rect 14319 35493 14343 35557
rect 14407 35493 14431 35557
rect 14495 35493 14519 35557
rect 14583 35493 14607 35557
rect 14671 35493 15000 35557
rect 0 35476 15000 35493
rect 0 35412 462 35476
rect 526 35412 620 35476
rect 684 35412 1390 35476
rect 1454 35412 1518 35476
rect 1582 35412 2382 35476
rect 2446 35412 2510 35476
rect 2574 35412 3374 35476
rect 3438 35412 3502 35476
rect 3566 35412 4366 35476
rect 4430 35412 4494 35476
rect 4558 35412 5358 35476
rect 5422 35412 5486 35476
rect 5550 35412 6350 35476
rect 6414 35412 6478 35476
rect 6542 35412 7342 35476
rect 7406 35412 7470 35476
rect 7534 35412 8334 35476
rect 8398 35412 8462 35476
rect 8526 35412 9326 35476
rect 9390 35412 9454 35476
rect 9518 35412 10318 35476
rect 10382 35412 10446 35476
rect 10510 35412 11310 35476
rect 11374 35412 11438 35476
rect 11502 35412 12302 35476
rect 12366 35412 12430 35476
rect 12494 35412 13294 35476
rect 13358 35412 13422 35476
rect 13486 35412 14255 35476
rect 14319 35412 14343 35476
rect 14407 35412 14431 35476
rect 14495 35412 14519 35476
rect 14583 35412 14607 35476
rect 14671 35412 15000 35476
rect 0 35395 15000 35412
rect 0 35331 462 35395
rect 526 35331 620 35395
rect 684 35331 1390 35395
rect 1454 35331 1518 35395
rect 1582 35331 2382 35395
rect 2446 35331 2510 35395
rect 2574 35331 3374 35395
rect 3438 35331 3502 35395
rect 3566 35331 4366 35395
rect 4430 35331 4494 35395
rect 4558 35331 5358 35395
rect 5422 35331 5486 35395
rect 5550 35331 6350 35395
rect 6414 35331 6478 35395
rect 6542 35331 7342 35395
rect 7406 35331 7470 35395
rect 7534 35331 8334 35395
rect 8398 35331 8462 35395
rect 8526 35331 9326 35395
rect 9390 35331 9454 35395
rect 9518 35331 10318 35395
rect 10382 35331 10446 35395
rect 10510 35331 11310 35395
rect 11374 35331 11438 35395
rect 11502 35331 12302 35395
rect 12366 35331 12430 35395
rect 12494 35331 13294 35395
rect 13358 35331 13422 35395
rect 13486 35331 14255 35395
rect 14319 35331 14343 35395
rect 14407 35331 14431 35395
rect 14495 35331 14519 35395
rect 14583 35331 14607 35395
rect 14671 35331 15000 35395
rect 0 35314 15000 35331
rect 0 35250 462 35314
rect 526 35250 620 35314
rect 684 35250 1390 35314
rect 1454 35250 1518 35314
rect 1582 35250 2382 35314
rect 2446 35250 2510 35314
rect 2574 35250 3374 35314
rect 3438 35250 3502 35314
rect 3566 35250 4366 35314
rect 4430 35250 4494 35314
rect 4558 35250 5358 35314
rect 5422 35250 5486 35314
rect 5550 35250 6350 35314
rect 6414 35250 6478 35314
rect 6542 35250 7342 35314
rect 7406 35250 7470 35314
rect 7534 35250 8334 35314
rect 8398 35250 8462 35314
rect 8526 35250 9326 35314
rect 9390 35250 9454 35314
rect 9518 35250 10318 35314
rect 10382 35250 10446 35314
rect 10510 35250 11310 35314
rect 11374 35250 11438 35314
rect 11502 35250 12302 35314
rect 12366 35250 12430 35314
rect 12494 35250 13294 35314
rect 13358 35250 13422 35314
rect 13486 35250 14255 35314
rect 14319 35250 14343 35314
rect 14407 35250 14431 35314
rect 14495 35250 14519 35314
rect 14583 35250 14607 35314
rect 14671 35250 15000 35314
rect 0 35233 15000 35250
rect 0 35169 462 35233
rect 526 35169 620 35233
rect 684 35169 1390 35233
rect 1454 35169 1518 35233
rect 1582 35169 2382 35233
rect 2446 35169 2510 35233
rect 2574 35169 3374 35233
rect 3438 35169 3502 35233
rect 3566 35169 4366 35233
rect 4430 35169 4494 35233
rect 4558 35169 5358 35233
rect 5422 35169 5486 35233
rect 5550 35169 6350 35233
rect 6414 35169 6478 35233
rect 6542 35169 7342 35233
rect 7406 35169 7470 35233
rect 7534 35169 8334 35233
rect 8398 35169 8462 35233
rect 8526 35169 9326 35233
rect 9390 35169 9454 35233
rect 9518 35169 10318 35233
rect 10382 35169 10446 35233
rect 10510 35169 11310 35233
rect 11374 35169 11438 35233
rect 11502 35169 12302 35233
rect 12366 35169 12430 35233
rect 12494 35169 13294 35233
rect 13358 35169 13422 35233
rect 13486 35169 14255 35233
rect 14319 35169 14343 35233
rect 14407 35169 14431 35233
rect 14495 35169 14519 35233
rect 14583 35169 14607 35233
rect 14671 35169 15000 35233
rect 0 35152 15000 35169
rect 0 35088 462 35152
rect 526 35088 620 35152
rect 684 35088 1390 35152
rect 1454 35088 1518 35152
rect 1582 35088 2382 35152
rect 2446 35088 2510 35152
rect 2574 35088 3374 35152
rect 3438 35088 3502 35152
rect 3566 35088 4366 35152
rect 4430 35088 4494 35152
rect 4558 35088 5358 35152
rect 5422 35088 5486 35152
rect 5550 35088 6350 35152
rect 6414 35088 6478 35152
rect 6542 35088 7342 35152
rect 7406 35088 7470 35152
rect 7534 35088 8334 35152
rect 8398 35088 8462 35152
rect 8526 35088 9326 35152
rect 9390 35088 9454 35152
rect 9518 35088 10318 35152
rect 10382 35088 10446 35152
rect 10510 35088 11310 35152
rect 11374 35088 11438 35152
rect 11502 35088 12302 35152
rect 12366 35088 12430 35152
rect 12494 35088 13294 35152
rect 13358 35088 13422 35152
rect 13486 35088 14255 35152
rect 14319 35088 14343 35152
rect 14407 35088 14431 35152
rect 14495 35088 14519 35152
rect 14583 35088 14607 35152
rect 14671 35088 15000 35152
rect 0 35071 15000 35088
rect 0 35007 462 35071
rect 526 35007 620 35071
rect 684 35007 1390 35071
rect 1454 35007 1518 35071
rect 1582 35007 2382 35071
rect 2446 35007 2510 35071
rect 2574 35007 3374 35071
rect 3438 35007 3502 35071
rect 3566 35007 4366 35071
rect 4430 35007 4494 35071
rect 4558 35007 5358 35071
rect 5422 35007 5486 35071
rect 5550 35007 6350 35071
rect 6414 35007 6478 35071
rect 6542 35007 7342 35071
rect 7406 35007 7470 35071
rect 7534 35007 8334 35071
rect 8398 35007 8462 35071
rect 8526 35007 9326 35071
rect 9390 35007 9454 35071
rect 9518 35007 10318 35071
rect 10382 35007 10446 35071
rect 10510 35007 11310 35071
rect 11374 35007 11438 35071
rect 11502 35007 12302 35071
rect 12366 35007 12430 35071
rect 12494 35007 13294 35071
rect 13358 35007 13422 35071
rect 13486 35007 14255 35071
rect 14319 35007 14343 35071
rect 14407 35007 14431 35071
rect 14495 35007 14519 35071
rect 14583 35007 14607 35071
rect 14671 35007 15000 35071
rect 0 34990 15000 35007
rect 0 34926 462 34990
rect 526 34926 620 34990
rect 684 34926 1390 34990
rect 1454 34926 1518 34990
rect 1582 34926 2382 34990
rect 2446 34926 2510 34990
rect 2574 34926 3374 34990
rect 3438 34926 3502 34990
rect 3566 34926 4366 34990
rect 4430 34926 4494 34990
rect 4558 34926 5358 34990
rect 5422 34926 5486 34990
rect 5550 34926 6350 34990
rect 6414 34926 6478 34990
rect 6542 34926 7342 34990
rect 7406 34926 7470 34990
rect 7534 34926 8334 34990
rect 8398 34926 8462 34990
rect 8526 34926 9326 34990
rect 9390 34926 9454 34990
rect 9518 34926 10318 34990
rect 10382 34926 10446 34990
rect 10510 34926 11310 34990
rect 11374 34926 11438 34990
rect 11502 34926 12302 34990
rect 12366 34926 12430 34990
rect 12494 34926 13294 34990
rect 13358 34926 13422 34990
rect 13486 34926 14255 34990
rect 14319 34926 14343 34990
rect 14407 34926 14431 34990
rect 14495 34926 14519 34990
rect 14583 34926 14607 34990
rect 14671 34926 15000 34990
rect 0 34909 15000 34926
rect 0 34845 462 34909
rect 526 34845 620 34909
rect 684 34845 1390 34909
rect 1454 34845 1518 34909
rect 1582 34845 2382 34909
rect 2446 34845 2510 34909
rect 2574 34845 3374 34909
rect 3438 34845 3502 34909
rect 3566 34845 4366 34909
rect 4430 34845 4494 34909
rect 4558 34845 5358 34909
rect 5422 34845 5486 34909
rect 5550 34845 6350 34909
rect 6414 34845 6478 34909
rect 6542 34845 7342 34909
rect 7406 34845 7470 34909
rect 7534 34845 8334 34909
rect 8398 34845 8462 34909
rect 8526 34845 9326 34909
rect 9390 34845 9454 34909
rect 9518 34845 10318 34909
rect 10382 34845 10446 34909
rect 10510 34845 11310 34909
rect 11374 34845 11438 34909
rect 11502 34845 12302 34909
rect 12366 34845 12430 34909
rect 12494 34845 13294 34909
rect 13358 34845 13422 34909
rect 13486 34845 14255 34909
rect 14319 34845 14343 34909
rect 14407 34845 14431 34909
rect 14495 34845 14519 34909
rect 14583 34845 14607 34909
rect 14671 34845 15000 34909
rect 0 34828 15000 34845
rect 0 34764 462 34828
rect 526 34764 620 34828
rect 684 34764 1390 34828
rect 1454 34764 1518 34828
rect 1582 34764 2382 34828
rect 2446 34764 2510 34828
rect 2574 34764 3374 34828
rect 3438 34764 3502 34828
rect 3566 34764 4366 34828
rect 4430 34764 4494 34828
rect 4558 34764 5358 34828
rect 5422 34764 5486 34828
rect 5550 34764 6350 34828
rect 6414 34764 6478 34828
rect 6542 34764 7342 34828
rect 7406 34764 7470 34828
rect 7534 34764 8334 34828
rect 8398 34764 8462 34828
rect 8526 34764 9326 34828
rect 9390 34764 9454 34828
rect 9518 34764 10318 34828
rect 10382 34764 10446 34828
rect 10510 34764 11310 34828
rect 11374 34764 11438 34828
rect 11502 34764 12302 34828
rect 12366 34764 12430 34828
rect 12494 34764 13294 34828
rect 13358 34764 13422 34828
rect 13486 34764 14255 34828
rect 14319 34764 14343 34828
rect 14407 34764 14431 34828
rect 14495 34764 14519 34828
rect 14583 34764 14607 34828
rect 14671 34764 15000 34828
rect 0 34757 15000 34764
rect 2877 34219 3071 34220
rect 2877 34155 2878 34219
rect 2942 34155 3006 34219
rect 3070 34155 3071 34219
rect 2877 34125 3071 34155
rect 2877 34061 2878 34125
rect 2942 34061 3006 34125
rect 3070 34061 3071 34125
rect 2877 34030 3071 34061
rect 2877 33966 2878 34030
rect 2942 33966 3006 34030
rect 3070 33966 3071 34030
rect 2877 33935 3071 33966
rect 2877 33871 2878 33935
rect 2942 33871 3006 33935
rect 3070 33871 3071 33935
rect 2877 33840 3071 33871
rect 1885 33831 2079 33832
rect 1885 33767 1886 33831
rect 1950 33767 2014 33831
rect 2078 33767 2079 33831
rect 1885 33749 2079 33767
rect 1885 33685 1886 33749
rect 1950 33685 2014 33749
rect 2078 33685 2079 33749
rect 1885 33666 2079 33685
rect 2877 33776 2878 33840
rect 2942 33776 3006 33840
rect 3070 33776 3071 33840
rect 2877 33745 3071 33776
rect 2877 33681 2878 33745
rect 2942 33681 3006 33745
rect 3070 33681 3071 33745
rect 2877 33680 3071 33681
rect 3869 34219 4063 34220
rect 3869 34155 3870 34219
rect 3934 34155 3998 34219
rect 4062 34155 4063 34219
rect 3869 34125 4063 34155
rect 3869 34061 3870 34125
rect 3934 34061 3998 34125
rect 4062 34061 4063 34125
rect 3869 34030 4063 34061
rect 3869 33966 3870 34030
rect 3934 33966 3998 34030
rect 4062 33966 4063 34030
rect 3869 33935 4063 33966
rect 3869 33871 3870 33935
rect 3934 33871 3998 33935
rect 4062 33871 4063 33935
rect 3869 33840 4063 33871
rect 3869 33776 3870 33840
rect 3934 33776 3998 33840
rect 4062 33776 4063 33840
rect 3869 33745 4063 33776
rect 3869 33681 3870 33745
rect 3934 33681 3998 33745
rect 4062 33681 4063 33745
rect 3869 33680 4063 33681
rect 4861 34219 5055 34220
rect 4861 34155 4862 34219
rect 4926 34155 4990 34219
rect 5054 34155 5055 34219
rect 4861 34125 5055 34155
rect 4861 34061 4862 34125
rect 4926 34061 4990 34125
rect 5054 34061 5055 34125
rect 4861 34030 5055 34061
rect 4861 33966 4862 34030
rect 4926 33966 4990 34030
rect 5054 33966 5055 34030
rect 4861 33935 5055 33966
rect 4861 33871 4862 33935
rect 4926 33871 4990 33935
rect 5054 33871 5055 33935
rect 4861 33840 5055 33871
rect 4861 33776 4862 33840
rect 4926 33776 4990 33840
rect 5054 33776 5055 33840
rect 4861 33745 5055 33776
rect 4861 33681 4862 33745
rect 4926 33681 4990 33745
rect 5054 33681 5055 33745
rect 4861 33680 5055 33681
rect 5853 34219 6047 34220
rect 5853 34155 5854 34219
rect 5918 34155 5982 34219
rect 6046 34155 6047 34219
rect 5853 34125 6047 34155
rect 5853 34061 5854 34125
rect 5918 34061 5982 34125
rect 6046 34061 6047 34125
rect 5853 34030 6047 34061
rect 5853 33966 5854 34030
rect 5918 33966 5982 34030
rect 6046 33966 6047 34030
rect 5853 33935 6047 33966
rect 5853 33871 5854 33935
rect 5918 33871 5982 33935
rect 6046 33871 6047 33935
rect 5853 33840 6047 33871
rect 5853 33776 5854 33840
rect 5918 33776 5982 33840
rect 6046 33776 6047 33840
rect 5853 33745 6047 33776
rect 5853 33681 5854 33745
rect 5918 33681 5982 33745
rect 6046 33681 6047 33745
rect 5853 33680 6047 33681
rect 6845 34219 7039 34220
rect 6845 34155 6846 34219
rect 6910 34155 6974 34219
rect 7038 34155 7039 34219
rect 6845 34125 7039 34155
rect 6845 34061 6846 34125
rect 6910 34061 6974 34125
rect 7038 34061 7039 34125
rect 6845 34030 7039 34061
rect 6845 33966 6846 34030
rect 6910 33966 6974 34030
rect 7038 33966 7039 34030
rect 6845 33935 7039 33966
rect 6845 33871 6846 33935
rect 6910 33871 6974 33935
rect 7038 33871 7039 33935
rect 6845 33840 7039 33871
rect 6845 33776 6846 33840
rect 6910 33776 6974 33840
rect 7038 33776 7039 33840
rect 6845 33745 7039 33776
rect 6845 33681 6846 33745
rect 6910 33681 6974 33745
rect 7038 33681 7039 33745
rect 6845 33680 7039 33681
rect 7837 34219 8031 34220
rect 7837 34155 7838 34219
rect 7902 34155 7966 34219
rect 8030 34155 8031 34219
rect 7837 34125 8031 34155
rect 7837 34061 7838 34125
rect 7902 34061 7966 34125
rect 8030 34061 8031 34125
rect 7837 34030 8031 34061
rect 7837 33966 7838 34030
rect 7902 33966 7966 34030
rect 8030 33966 8031 34030
rect 7837 33935 8031 33966
rect 7837 33871 7838 33935
rect 7902 33871 7966 33935
rect 8030 33871 8031 33935
rect 7837 33840 8031 33871
rect 7837 33776 7838 33840
rect 7902 33776 7966 33840
rect 8030 33776 8031 33840
rect 7837 33745 8031 33776
rect 7837 33681 7838 33745
rect 7902 33681 7966 33745
rect 8030 33681 8031 33745
rect 7837 33680 8031 33681
rect 8829 34219 9023 34220
rect 8829 34155 8830 34219
rect 8894 34155 8958 34219
rect 9022 34155 9023 34219
rect 8829 34125 9023 34155
rect 8829 34061 8830 34125
rect 8894 34061 8958 34125
rect 9022 34061 9023 34125
rect 8829 34030 9023 34061
rect 8829 33966 8830 34030
rect 8894 33966 8958 34030
rect 9022 33966 9023 34030
rect 8829 33935 9023 33966
rect 8829 33871 8830 33935
rect 8894 33871 8958 33935
rect 9022 33871 9023 33935
rect 8829 33840 9023 33871
rect 8829 33776 8830 33840
rect 8894 33776 8958 33840
rect 9022 33776 9023 33840
rect 8829 33745 9023 33776
rect 8829 33681 8830 33745
rect 8894 33681 8958 33745
rect 9022 33681 9023 33745
rect 8829 33680 9023 33681
rect 9821 34219 10015 34220
rect 9821 34155 9822 34219
rect 9886 34155 9950 34219
rect 10014 34155 10015 34219
rect 9821 34125 10015 34155
rect 9821 34061 9822 34125
rect 9886 34061 9950 34125
rect 10014 34061 10015 34125
rect 9821 34030 10015 34061
rect 9821 33966 9822 34030
rect 9886 33966 9950 34030
rect 10014 33966 10015 34030
rect 9821 33935 10015 33966
rect 9821 33871 9822 33935
rect 9886 33871 9950 33935
rect 10014 33871 10015 33935
rect 9821 33840 10015 33871
rect 9821 33776 9822 33840
rect 9886 33776 9950 33840
rect 10014 33776 10015 33840
rect 9821 33745 10015 33776
rect 9821 33681 9822 33745
rect 9886 33681 9950 33745
rect 10014 33681 10015 33745
rect 9821 33680 10015 33681
rect 10813 34219 11007 34220
rect 10813 34155 10814 34219
rect 10878 34155 10942 34219
rect 11006 34155 11007 34219
rect 10813 34125 11007 34155
rect 10813 34061 10814 34125
rect 10878 34061 10942 34125
rect 11006 34061 11007 34125
rect 10813 34030 11007 34061
rect 10813 33966 10814 34030
rect 10878 33966 10942 34030
rect 11006 33966 11007 34030
rect 10813 33935 11007 33966
rect 10813 33871 10814 33935
rect 10878 33871 10942 33935
rect 11006 33871 11007 33935
rect 10813 33840 11007 33871
rect 10813 33776 10814 33840
rect 10878 33776 10942 33840
rect 11006 33776 11007 33840
rect 10813 33745 11007 33776
rect 10813 33681 10814 33745
rect 10878 33681 10942 33745
rect 11006 33681 11007 33745
rect 10813 33680 11007 33681
rect 11805 34219 11999 34220
rect 11805 34155 11806 34219
rect 11870 34155 11934 34219
rect 11998 34155 11999 34219
rect 11805 34125 11999 34155
rect 11805 34061 11806 34125
rect 11870 34061 11934 34125
rect 11998 34061 11999 34125
rect 11805 34030 11999 34061
rect 11805 33966 11806 34030
rect 11870 33966 11934 34030
rect 11998 33966 11999 34030
rect 11805 33935 11999 33966
rect 11805 33871 11806 33935
rect 11870 33871 11934 33935
rect 11998 33871 11999 33935
rect 11805 33840 11999 33871
rect 11805 33776 11806 33840
rect 11870 33776 11934 33840
rect 11998 33776 11999 33840
rect 11805 33745 11999 33776
rect 11805 33681 11806 33745
rect 11870 33681 11934 33745
rect 11998 33681 11999 33745
rect 11805 33680 11999 33681
rect 12797 33954 12991 33955
rect 12797 33890 12798 33954
rect 12862 33890 12926 33954
rect 12990 33890 12991 33954
rect 12797 33860 12991 33890
rect 12797 33796 12798 33860
rect 12862 33796 12926 33860
rect 12990 33796 12991 33860
rect 12797 33765 12991 33796
rect 12797 33701 12798 33765
rect 12862 33701 12926 33765
rect 12990 33701 12991 33765
rect 1885 33602 1886 33666
rect 1950 33602 2014 33666
rect 2078 33602 2079 33666
rect 1885 33583 2079 33602
rect 1885 33519 1886 33583
rect 1950 33519 2014 33583
rect 2078 33519 2079 33583
rect 1885 33500 2079 33519
rect 1885 33436 1886 33500
rect 1950 33436 2014 33500
rect 2078 33436 2079 33500
rect 1885 33417 2079 33436
rect 1885 33353 1886 33417
rect 1950 33353 2014 33417
rect 2078 33353 2079 33417
rect 12797 33670 12991 33701
rect 12797 33606 12798 33670
rect 12862 33606 12926 33670
rect 12990 33606 12991 33670
rect 12797 33575 12991 33606
rect 12797 33511 12798 33575
rect 12862 33511 12926 33575
rect 12990 33511 12991 33575
rect 12797 33480 12991 33511
rect 12797 33416 12798 33480
rect 12862 33416 12926 33480
rect 12990 33416 12991 33480
rect 12797 33415 12991 33416
rect 1885 33334 2079 33353
rect 1885 33270 1886 33334
rect 1950 33270 2014 33334
rect 2078 33270 2079 33334
rect 1885 33269 2079 33270
rect 13789 32983 13957 32984
rect 13789 32919 13790 32983
rect 13854 32919 13892 32983
rect 13956 32919 13957 32983
rect 13789 32903 13957 32919
rect 13789 32839 13790 32903
rect 13854 32839 13892 32903
rect 13956 32839 13957 32903
rect 13789 32823 13957 32839
rect 13789 32759 13790 32823
rect 13854 32759 13892 32823
rect 13956 32759 13957 32823
rect 13789 32743 13957 32759
rect 13789 32679 13790 32743
rect 13854 32679 13892 32743
rect 13956 32679 13957 32743
rect 13789 32663 13957 32679
rect 13789 32599 13790 32663
rect 13854 32599 13892 32663
rect 13956 32599 13957 32663
rect 13789 32583 13957 32599
rect 13789 32519 13790 32583
rect 13854 32519 13892 32583
rect 13956 32519 13957 32583
rect 13789 32503 13957 32519
rect 13789 32439 13790 32503
rect 13854 32439 13892 32503
rect 13956 32439 13957 32503
rect 13789 32423 13957 32439
tri 1024 32359 1079 32414 se
tri 1008 32343 1024 32359 se
rect 1024 32343 1079 32359
tri 944 32279 1008 32343 se
rect 1008 32279 1079 32343
tri 928 32263 944 32279 se
rect 944 32263 1079 32279
tri 864 32199 928 32263 se
rect 928 32199 1079 32263
tri 848 32183 864 32199 se
rect 864 32183 1079 32199
tri 784 32119 848 32183 se
rect 848 32119 1079 32183
tri 768 32103 784 32119 se
rect 784 32103 1079 32119
tri 706 32041 768 32103 se
rect 768 32041 1079 32103
rect 706 32017 1079 32041
rect 706 31953 862 32017
rect 926 31953 990 32017
rect 1054 31953 1079 32017
rect 706 31936 1079 31953
rect 706 31872 862 31936
rect 926 31872 990 31936
rect 1054 31872 1079 31936
rect 706 31855 1079 31872
rect 706 31791 862 31855
rect 926 31791 990 31855
rect 1054 31791 1079 31855
rect 706 31774 1079 31791
rect 706 31710 862 31774
rect 926 31710 990 31774
rect 1054 31710 1079 31774
rect 706 31693 1079 31710
rect 706 31629 862 31693
rect 926 31629 990 31693
rect 1054 31629 1079 31693
rect 706 31612 1079 31629
rect 706 31548 862 31612
rect 926 31548 990 31612
rect 1054 31548 1079 31612
rect 706 31531 1079 31548
rect 706 31467 862 31531
rect 926 31467 990 31531
rect 1054 31467 1079 31531
rect 706 31450 1079 31467
rect 706 31386 862 31450
rect 926 31386 990 31450
rect 1054 31386 1079 31450
rect 706 31369 1079 31386
rect 706 31305 862 31369
rect 926 31305 990 31369
rect 1054 31305 1079 31369
rect 706 31288 1079 31305
rect 706 31224 862 31288
rect 926 31224 990 31288
rect 1054 31224 1079 31288
rect 706 31207 1079 31224
rect 706 31143 862 31207
rect 926 31143 990 31207
rect 1054 31143 1079 31207
rect 706 31125 1079 31143
rect 706 31061 862 31125
rect 926 31061 990 31125
rect 1054 31061 1079 31125
rect 706 31043 1079 31061
rect 706 30979 862 31043
rect 926 30979 990 31043
rect 1054 30979 1079 31043
rect 706 30961 1079 30979
rect 706 30897 862 30961
rect 926 30897 990 30961
rect 1054 30897 1079 30961
rect 706 30879 1079 30897
rect 706 30815 862 30879
rect 926 30815 990 30879
rect 1054 30815 1079 30879
rect 706 30797 1079 30815
rect 706 30733 862 30797
rect 926 30733 990 30797
rect 1054 30733 1079 30797
rect 706 30715 1079 30733
rect 706 30651 862 30715
rect 926 30651 990 30715
rect 1054 30651 1079 30715
rect 706 30633 1079 30651
rect 706 30569 862 30633
rect 926 30569 990 30633
rect 1054 30569 1079 30633
rect 706 30551 1079 30569
rect 706 30487 862 30551
rect 926 30487 990 30551
rect 1054 30487 1079 30551
rect 706 30469 1079 30487
rect 706 30405 862 30469
rect 926 30405 990 30469
rect 1054 30405 1079 30469
rect 706 30387 1079 30405
rect 706 30323 862 30387
rect 926 30323 990 30387
rect 1054 30323 1079 30387
rect 706 30305 1079 30323
rect 706 30241 862 30305
rect 926 30241 990 30305
rect 1054 30241 1079 30305
rect 706 30223 1079 30241
rect 706 30159 862 30223
rect 926 30159 990 30223
rect 1054 30159 1079 30223
rect 706 30141 1079 30159
rect 706 30077 862 30141
rect 926 30077 990 30141
rect 1054 30077 1079 30141
rect 706 30059 1079 30077
rect 706 29995 862 30059
rect 926 29995 990 30059
rect 1054 29995 1079 30059
rect 706 29977 1079 29995
rect 706 29913 862 29977
rect 926 29913 990 29977
rect 1054 29913 1079 29977
rect 706 29895 1079 29913
rect 706 29831 862 29895
rect 926 29831 990 29895
rect 1054 29831 1079 29895
rect 706 29813 1079 29831
rect 706 29749 862 29813
rect 926 29749 990 29813
rect 1054 29749 1079 29813
rect 706 29731 1079 29749
rect 706 29667 862 29731
rect 926 29667 990 29731
rect 1054 29667 1079 29731
rect 706 29649 1079 29667
rect 706 29585 862 29649
rect 926 29585 990 29649
rect 1054 29585 1079 29649
rect 706 29567 1079 29585
rect 706 29503 862 29567
rect 926 29503 990 29567
rect 1054 29503 1079 29567
rect 706 29485 1079 29503
rect 706 29421 862 29485
rect 926 29421 990 29485
rect 1054 29421 1079 29485
rect 706 29367 1079 29421
tri 706 29364 709 29367 ne
rect 709 29364 1079 29367
tri 709 29300 773 29364 ne
rect 773 29300 1079 29364
tri 773 29283 790 29300 ne
rect 790 29283 1079 29300
tri 790 29219 854 29283 ne
rect 854 29219 1079 29283
tri 854 29202 871 29219 ne
rect 871 29202 1079 29219
tri 871 29138 935 29202 ne
rect 935 29138 1079 29202
tri 935 29121 952 29138 ne
rect 952 29121 1079 29138
tri 952 29057 1016 29121 ne
rect 1016 29057 1079 29121
tri 1016 29040 1033 29057 ne
rect 1033 29040 1079 29057
tri 1033 28994 1079 29040 ne
rect 13789 32359 13790 32423
rect 13854 32359 13892 32423
rect 13956 32359 13957 32423
rect 13789 32343 13957 32359
rect 13789 32279 13790 32343
rect 13854 32279 13892 32343
rect 13956 32279 13957 32343
rect 13789 32263 13957 32279
rect 13789 32199 13790 32263
rect 13854 32199 13892 32263
rect 13956 32199 13957 32263
rect 13789 32183 13957 32199
rect 13789 32119 13790 32183
rect 13854 32119 13892 32183
rect 13956 32119 13957 32183
rect 13789 32103 13957 32119
rect 13789 32039 13790 32103
rect 13854 32039 13892 32103
rect 13956 32039 13957 32103
rect 13789 32023 13957 32039
rect 13789 31959 13790 32023
rect 13854 31959 13892 32023
rect 13956 31959 13957 32023
rect 13789 31943 13957 31959
rect 13789 31879 13790 31943
rect 13854 31879 13892 31943
rect 13956 31879 13957 31943
rect 13789 31863 13957 31879
rect 13789 31799 13790 31863
rect 13854 31799 13892 31863
rect 13956 31799 13957 31863
rect 13789 31783 13957 31799
rect 13789 31719 13790 31783
rect 13854 31719 13892 31783
rect 13956 31719 13957 31783
rect 13789 31703 13957 31719
rect 13789 31639 13790 31703
rect 13854 31639 13892 31703
rect 13956 31639 13957 31703
rect 13789 31623 13957 31639
rect 13789 31559 13790 31623
rect 13854 31559 13892 31623
rect 13956 31559 13957 31623
rect 13789 31543 13957 31559
rect 13789 31479 13790 31543
rect 13854 31479 13892 31543
rect 13956 31479 13957 31543
rect 13789 31463 13957 31479
rect 13789 31399 13790 31463
rect 13854 31399 13892 31463
rect 13956 31399 13957 31463
rect 13789 31383 13957 31399
rect 13789 31319 13790 31383
rect 13854 31319 13892 31383
rect 13956 31319 13957 31383
rect 13789 31303 13957 31319
rect 13789 31239 13790 31303
rect 13854 31239 13892 31303
rect 13956 31239 13957 31303
rect 13789 31223 13957 31239
rect 13789 31159 13790 31223
rect 13854 31159 13892 31223
rect 13956 31159 13957 31223
rect 13789 31143 13957 31159
rect 13789 31079 13790 31143
rect 13854 31079 13892 31143
rect 13956 31079 13957 31143
rect 13789 31063 13957 31079
rect 13789 30999 13790 31063
rect 13854 30999 13892 31063
rect 13956 30999 13957 31063
rect 13789 30983 13957 30999
rect 13789 30919 13790 30983
rect 13854 30919 13892 30983
rect 13956 30919 13957 30983
rect 13789 30903 13957 30919
rect 13789 30839 13790 30903
rect 13854 30839 13892 30903
rect 13956 30839 13957 30903
rect 13789 30822 13957 30839
rect 13789 30758 13790 30822
rect 13854 30758 13892 30822
rect 13956 30758 13957 30822
rect 13789 30741 13957 30758
rect 13789 30677 13790 30741
rect 13854 30677 13892 30741
rect 13956 30677 13957 30741
rect 13789 30660 13957 30677
rect 13789 30596 13790 30660
rect 13854 30596 13892 30660
rect 13956 30596 13957 30660
rect 13789 30579 13957 30596
rect 13789 30515 13790 30579
rect 13854 30515 13892 30579
rect 13956 30515 13957 30579
rect 13789 30498 13957 30515
rect 13789 30434 13790 30498
rect 13854 30434 13892 30498
rect 13956 30434 13957 30498
rect 13789 30417 13957 30434
rect 13789 30353 13790 30417
rect 13854 30353 13892 30417
rect 13956 30353 13957 30417
rect 13789 30336 13957 30353
rect 13789 30272 13790 30336
rect 13854 30272 13892 30336
rect 13956 30272 13957 30336
rect 13789 30255 13957 30272
rect 13789 30191 13790 30255
rect 13854 30191 13892 30255
rect 13956 30191 13957 30255
rect 13789 30174 13957 30191
rect 13789 30110 13790 30174
rect 13854 30110 13892 30174
rect 13956 30110 13957 30174
rect 13789 30093 13957 30110
rect 13789 30029 13790 30093
rect 13854 30029 13892 30093
rect 13956 30029 13957 30093
rect 13789 30012 13957 30029
rect 13789 29948 13790 30012
rect 13854 29948 13892 30012
rect 13956 29948 13957 30012
rect 13789 29931 13957 29948
rect 13789 29867 13790 29931
rect 13854 29867 13892 29931
rect 13956 29867 13957 29931
rect 13789 29850 13957 29867
rect 13789 29786 13790 29850
rect 13854 29786 13892 29850
rect 13956 29786 13957 29850
rect 13789 29769 13957 29786
rect 13789 29705 13790 29769
rect 13854 29705 13892 29769
rect 13956 29705 13957 29769
rect 13789 29688 13957 29705
rect 13789 29624 13790 29688
rect 13854 29624 13892 29688
rect 13956 29624 13957 29688
rect 13789 29607 13957 29624
rect 13789 29543 13790 29607
rect 13854 29543 13892 29607
rect 13956 29543 13957 29607
rect 13789 29526 13957 29543
rect 13789 29462 13790 29526
rect 13854 29462 13892 29526
rect 13956 29462 13957 29526
rect 13789 29445 13957 29462
rect 13789 29381 13790 29445
rect 13854 29381 13892 29445
rect 13956 29381 13957 29445
rect 13789 29364 13957 29381
rect 13789 29300 13790 29364
rect 13854 29300 13892 29364
rect 13956 29300 13957 29364
rect 13789 29283 13957 29300
rect 13789 29219 13790 29283
rect 13854 29219 13892 29283
rect 13956 29219 13957 29283
rect 13789 29202 13957 29219
rect 13789 29138 13790 29202
rect 13854 29138 13892 29202
rect 13956 29138 13957 29202
rect 13789 29121 13957 29138
rect 13789 29057 13790 29121
rect 13854 29057 13892 29121
rect 13956 29057 13957 29121
rect 13789 29040 13957 29057
rect 13789 28976 13790 29040
rect 13854 28976 13892 29040
rect 13956 28976 13957 29040
rect 13789 28959 13957 28976
rect 13789 28895 13790 28959
rect 13854 28895 13892 28959
rect 13956 28895 13957 28959
rect 13789 28878 13957 28895
rect 13789 28814 13790 28878
rect 13854 28814 13892 28878
rect 13956 28814 13957 28878
rect 13789 28797 13957 28814
rect 13789 28733 13790 28797
rect 13854 28733 13892 28797
rect 13956 28733 13957 28797
rect 13789 28716 13957 28733
rect 13789 28652 13790 28716
rect 13854 28652 13892 28716
rect 13956 28652 13957 28716
rect 13789 28635 13957 28652
rect 13789 28571 13790 28635
rect 13854 28571 13892 28635
rect 13956 28571 13957 28635
rect 13789 28554 13957 28571
rect 13789 28490 13790 28554
rect 13854 28490 13892 28554
rect 13956 28490 13957 28554
rect 13789 28473 13957 28490
rect 13789 28409 13790 28473
rect 13854 28409 13892 28473
rect 13956 28409 13957 28473
rect 13789 28392 13957 28409
rect 960 28348 1500 28349
rect 960 28284 963 28348
rect 1027 28284 1057 28348
rect 1121 28284 1151 28348
rect 1215 28284 1245 28348
rect 1309 28284 1339 28348
rect 1403 28284 1433 28348
rect 1497 28284 1500 28348
rect 960 28268 1500 28284
rect 960 28204 963 28268
rect 1027 28204 1057 28268
rect 1121 28204 1151 28268
rect 1215 28204 1245 28268
rect 1309 28204 1339 28268
rect 1403 28204 1433 28268
rect 1497 28204 1500 28268
rect 960 28188 1500 28204
rect 960 28124 963 28188
rect 1027 28124 1057 28188
rect 1121 28124 1151 28188
rect 1215 28124 1245 28188
rect 1309 28124 1339 28188
rect 1403 28124 1433 28188
rect 1497 28124 1500 28188
rect 960 28108 1500 28124
rect 960 28044 963 28108
rect 1027 28044 1057 28108
rect 1121 28044 1151 28108
rect 1215 28044 1245 28108
rect 1309 28044 1339 28108
rect 1403 28044 1433 28108
rect 1497 28044 1500 28108
rect 960 28028 1500 28044
rect 960 27964 963 28028
rect 1027 27964 1057 28028
rect 1121 27964 1151 28028
rect 1215 27964 1245 28028
rect 1309 27964 1339 28028
rect 1403 27964 1433 28028
rect 1497 27964 1500 28028
rect 960 27948 1500 27964
rect 960 27884 963 27948
rect 1027 27884 1057 27948
rect 1121 27884 1151 27948
rect 1215 27884 1245 27948
rect 1309 27884 1339 27948
rect 1403 27884 1433 27948
rect 1497 27884 1500 27948
rect 960 27867 1500 27884
rect 960 27803 963 27867
rect 1027 27803 1057 27867
rect 1121 27803 1151 27867
rect 1215 27803 1245 27867
rect 1309 27803 1339 27867
rect 1403 27803 1433 27867
rect 1497 27803 1500 27867
rect 960 27786 1500 27803
rect 960 27722 963 27786
rect 1027 27722 1057 27786
rect 1121 27722 1151 27786
rect 1215 27722 1245 27786
rect 1309 27722 1339 27786
rect 1403 27722 1433 27786
rect 1497 27722 1500 27786
rect 960 27705 1500 27722
rect 960 27641 963 27705
rect 1027 27641 1057 27705
rect 1121 27641 1151 27705
rect 1215 27641 1245 27705
rect 1309 27641 1339 27705
rect 1403 27641 1433 27705
rect 1497 27641 1500 27705
rect 960 27624 1500 27641
rect 960 27560 963 27624
rect 1027 27560 1057 27624
rect 1121 27560 1151 27624
rect 1215 27560 1245 27624
rect 1309 27560 1339 27624
rect 1403 27560 1433 27624
rect 1497 27560 1500 27624
rect 960 27543 1500 27560
rect 960 27479 963 27543
rect 1027 27479 1057 27543
rect 1121 27479 1151 27543
rect 1215 27479 1245 27543
rect 1309 27479 1339 27543
rect 1403 27479 1433 27543
rect 1497 27479 1500 27543
rect 960 27462 1500 27479
rect 960 27398 963 27462
rect 1027 27398 1057 27462
rect 1121 27398 1151 27462
rect 1215 27398 1245 27462
rect 1309 27398 1339 27462
rect 1403 27398 1433 27462
rect 1497 27398 1500 27462
rect 960 27381 1500 27398
rect 960 27317 963 27381
rect 1027 27317 1057 27381
rect 1121 27317 1151 27381
rect 1215 27317 1245 27381
rect 1309 27317 1339 27381
rect 1403 27317 1433 27381
rect 1497 27317 1500 27381
rect 960 27300 1500 27317
rect 960 27236 963 27300
rect 1027 27236 1057 27300
rect 1121 27236 1151 27300
rect 1215 27236 1245 27300
rect 1309 27236 1339 27300
rect 1403 27236 1433 27300
rect 1497 27236 1500 27300
rect 960 27219 1500 27236
rect 960 27155 963 27219
rect 1027 27155 1057 27219
rect 1121 27155 1151 27219
rect 1215 27155 1245 27219
rect 1309 27155 1339 27219
rect 1403 27155 1433 27219
rect 1497 27155 1500 27219
rect 960 27138 1500 27155
rect 960 27074 963 27138
rect 1027 27074 1057 27138
rect 1121 27074 1151 27138
rect 1215 27074 1245 27138
rect 1309 27074 1339 27138
rect 1403 27074 1433 27138
rect 1497 27074 1500 27138
rect 13789 28328 13790 28392
rect 13854 28328 13892 28392
rect 13956 28328 13957 28392
rect 13789 28311 13957 28328
rect 13789 28247 13790 28311
rect 13854 28247 13892 28311
rect 13956 28247 13957 28311
rect 13789 28230 13957 28247
rect 13789 28166 13790 28230
rect 13854 28166 13892 28230
rect 13956 28166 13957 28230
rect 13789 28149 13957 28166
rect 13789 28085 13790 28149
rect 13854 28085 13892 28149
rect 13956 28085 13957 28149
rect 13789 28068 13957 28085
rect 13789 28004 13790 28068
rect 13854 28004 13892 28068
rect 13956 28004 13957 28068
rect 13789 27987 13957 28004
rect 13789 27923 13790 27987
rect 13854 27923 13892 27987
rect 13956 27923 13957 27987
rect 13789 27906 13957 27923
rect 13789 27842 13790 27906
rect 13854 27842 13892 27906
rect 13956 27842 13957 27906
rect 13789 27825 13957 27842
rect 13789 27761 13790 27825
rect 13854 27761 13892 27825
rect 13956 27761 13957 27825
rect 13789 27744 13957 27761
rect 13789 27680 13790 27744
rect 13854 27680 13892 27744
rect 13956 27680 13957 27744
rect 13789 27663 13957 27680
rect 13789 27599 13790 27663
rect 13854 27599 13892 27663
rect 13956 27599 13957 27663
rect 13789 27582 13957 27599
rect 13789 27518 13790 27582
rect 13854 27518 13892 27582
rect 13956 27518 13957 27582
rect 13789 27501 13957 27518
rect 13789 27437 13790 27501
rect 13854 27437 13892 27501
rect 13956 27437 13957 27501
rect 13789 27420 13957 27437
rect 13789 27356 13790 27420
rect 13854 27356 13892 27420
rect 13956 27356 13957 27420
rect 13789 27339 13957 27356
rect 13789 27275 13790 27339
rect 13854 27275 13892 27339
rect 13956 27275 13957 27339
rect 13789 27258 13957 27275
rect 13789 27194 13790 27258
rect 13854 27194 13892 27258
rect 13956 27194 13957 27258
rect 13789 27177 13957 27194
rect 13789 27113 13790 27177
rect 13854 27113 13892 27177
rect 13956 27113 13957 27177
rect 13789 27112 13957 27113
rect 13973 27347 14039 27348
rect 13973 27283 13974 27347
rect 14038 27283 14039 27347
rect 13973 27262 14039 27283
rect 13973 27198 13974 27262
rect 14038 27198 14039 27262
rect 13973 27176 14039 27198
rect 13973 27112 13974 27176
rect 14038 27112 14039 27176
rect 13973 27111 14039 27112
rect 960 27057 1500 27074
rect 960 26993 963 27057
rect 1027 26993 1057 27057
rect 1121 26993 1151 27057
rect 1215 26993 1245 27057
rect 1309 26993 1339 27057
rect 1403 26993 1433 27057
rect 1497 26993 1500 27057
rect 960 26976 1500 26993
rect 960 26912 963 26976
rect 1027 26912 1057 26976
rect 1121 26912 1151 26976
rect 1215 26912 1245 26976
rect 1309 26912 1339 26976
rect 1403 26912 1433 26976
rect 1497 26912 1500 26976
rect 960 26895 1500 26912
rect 960 26831 963 26895
rect 1027 26831 1057 26895
rect 1121 26831 1151 26895
rect 1215 26831 1245 26895
rect 1309 26831 1339 26895
rect 1403 26831 1433 26895
rect 1497 26831 1500 26895
rect 960 26814 1500 26831
rect 960 26750 963 26814
rect 1027 26750 1057 26814
rect 1121 26750 1151 26814
rect 1215 26750 1245 26814
rect 1309 26750 1339 26814
rect 1403 26750 1433 26814
rect 1497 26750 1500 26814
rect 960 26733 1500 26750
rect 960 26669 963 26733
rect 1027 26669 1057 26733
rect 1121 26669 1151 26733
rect 1215 26669 1245 26733
rect 1309 26669 1339 26733
rect 1403 26669 1433 26733
rect 1497 26669 1500 26733
rect 960 26652 1500 26669
rect 960 26588 963 26652
rect 1027 26588 1057 26652
rect 1121 26588 1151 26652
rect 1215 26588 1245 26652
rect 1309 26588 1339 26652
rect 1403 26588 1433 26652
rect 1497 26588 1500 26652
rect 960 26571 1500 26588
rect 960 26507 963 26571
rect 1027 26507 1057 26571
rect 1121 26507 1151 26571
rect 1215 26507 1245 26571
rect 1309 26507 1339 26571
rect 1403 26507 1433 26571
rect 1497 26507 1500 26571
rect 960 26490 1500 26507
rect 960 26426 963 26490
rect 1027 26426 1057 26490
rect 1121 26426 1151 26490
rect 1215 26426 1245 26490
rect 1309 26426 1339 26490
rect 1403 26426 1433 26490
rect 1497 26426 1500 26490
rect 960 26409 1500 26426
rect 960 26345 963 26409
rect 1027 26345 1057 26409
rect 1121 26345 1151 26409
rect 1215 26345 1245 26409
rect 1309 26345 1339 26409
rect 1403 26345 1433 26409
rect 1497 26345 1500 26409
rect 13646 27074 14040 27075
rect 13646 27010 13649 27074
rect 13713 27010 13757 27074
rect 13821 27010 13865 27074
rect 13929 27010 13973 27074
rect 14037 27010 14040 27074
rect 13646 26964 14040 27010
rect 13646 26900 13649 26964
rect 13713 26900 13757 26964
rect 13821 26900 13865 26964
rect 13929 26900 13973 26964
rect 14037 26900 14040 26964
rect 13646 26854 14040 26900
rect 13646 26790 13649 26854
rect 13713 26790 13757 26854
rect 13821 26790 13865 26854
rect 13929 26790 13973 26854
rect 14037 26790 14040 26854
rect 13646 26744 14040 26790
rect 13646 26680 13649 26744
rect 13713 26680 13757 26744
rect 13821 26680 13865 26744
rect 13929 26680 13973 26744
rect 14037 26680 14040 26744
rect 13646 26634 14040 26680
rect 13646 26570 13649 26634
rect 13713 26570 13757 26634
rect 13821 26570 13865 26634
rect 13929 26570 13973 26634
rect 14037 26570 14040 26634
rect 13646 26524 14040 26570
rect 13646 26460 13649 26524
rect 13713 26460 13757 26524
rect 13821 26460 13865 26524
rect 13929 26460 13973 26524
rect 14037 26460 14040 26524
rect 13646 26413 14040 26460
rect 13646 26349 13649 26413
rect 13713 26349 13757 26413
rect 13821 26349 13865 26413
rect 13929 26349 13973 26413
rect 14037 26349 14040 26413
rect 13646 26348 14040 26349
rect 960 26328 1500 26345
rect 960 26264 963 26328
rect 1027 26264 1057 26328
rect 1121 26264 1151 26328
rect 1215 26264 1245 26328
rect 1309 26264 1339 26328
rect 1403 26264 1433 26328
rect 1497 26264 1500 26328
rect 960 26247 1500 26264
rect 960 26183 963 26247
rect 1027 26183 1057 26247
rect 1121 26183 1151 26247
rect 1215 26183 1245 26247
rect 1309 26183 1339 26247
rect 1403 26183 1433 26247
rect 1497 26183 1500 26247
rect 960 26166 1500 26183
rect 960 26102 963 26166
rect 1027 26102 1057 26166
rect 1121 26102 1151 26166
rect 1215 26102 1245 26166
rect 1309 26102 1339 26166
rect 1403 26102 1433 26166
rect 1497 26102 1500 26166
rect 960 26085 1500 26102
rect 960 26021 963 26085
rect 1027 26021 1057 26085
rect 1121 26021 1151 26085
rect 1215 26021 1245 26085
rect 1309 26021 1339 26085
rect 1403 26021 1433 26085
rect 1497 26021 1500 26085
rect 960 26004 1500 26021
rect 960 25940 963 26004
rect 1027 25940 1057 26004
rect 1121 25940 1151 26004
rect 1215 25940 1245 26004
rect 1309 25940 1339 26004
rect 1403 25940 1433 26004
rect 1497 25940 1500 26004
rect 960 25923 1500 25940
rect 960 25859 963 25923
rect 1027 25859 1057 25923
rect 1121 25859 1151 25923
rect 1215 25859 1245 25923
rect 1309 25859 1339 25923
rect 1403 25859 1433 25923
rect 1497 25859 1500 25923
rect 960 25842 1500 25859
rect 960 25778 963 25842
rect 1027 25778 1057 25842
rect 1121 25778 1151 25842
rect 1215 25778 1245 25842
rect 1309 25778 1339 25842
rect 1403 25778 1433 25842
rect 1497 25778 1500 25842
rect 960 25761 1500 25778
rect 960 25697 963 25761
rect 1027 25697 1057 25761
rect 1121 25697 1151 25761
rect 1215 25697 1245 25761
rect 1309 25697 1339 25761
rect 1403 25697 1433 25761
rect 1497 25697 1500 25761
rect 960 25680 1500 25697
rect 960 25616 963 25680
rect 1027 25616 1057 25680
rect 1121 25616 1151 25680
rect 1215 25616 1245 25680
rect 1309 25616 1339 25680
rect 1403 25616 1433 25680
rect 1497 25616 1500 25680
rect 960 25599 1500 25616
rect 960 25535 963 25599
rect 1027 25535 1057 25599
rect 1121 25535 1151 25599
rect 1215 25535 1245 25599
rect 1309 25535 1339 25599
rect 1403 25535 1433 25599
rect 1497 25535 1500 25599
rect 960 25518 1500 25535
rect 960 25454 963 25518
rect 1027 25454 1057 25518
rect 1121 25454 1151 25518
rect 1215 25454 1245 25518
rect 1309 25454 1339 25518
rect 1403 25454 1433 25518
rect 1497 25454 1500 25518
rect 960 25437 1500 25454
rect 960 25373 963 25437
rect 1027 25373 1057 25437
rect 1121 25373 1151 25437
rect 1215 25373 1245 25437
rect 1309 25373 1339 25437
rect 1403 25373 1433 25437
rect 1497 25373 1500 25437
rect 960 25356 1500 25373
rect 960 25292 963 25356
rect 1027 25292 1057 25356
rect 1121 25292 1151 25356
rect 1215 25292 1245 25356
rect 1309 25292 1339 25356
rect 1403 25292 1433 25356
rect 1497 25292 1500 25356
rect 960 25275 1500 25292
rect 960 25211 963 25275
rect 1027 25211 1057 25275
rect 1121 25211 1151 25275
rect 1215 25211 1245 25275
rect 1309 25211 1339 25275
rect 1403 25211 1433 25275
rect 1497 25211 1500 25275
rect 960 25194 1500 25211
rect 960 25130 963 25194
rect 1027 25130 1057 25194
rect 1121 25130 1151 25194
rect 1215 25130 1245 25194
rect 1309 25130 1339 25194
rect 1403 25130 1433 25194
rect 1497 25130 1500 25194
rect 960 25113 1500 25130
rect 960 25049 963 25113
rect 1027 25049 1057 25113
rect 1121 25049 1151 25113
rect 1215 25049 1245 25113
rect 1309 25049 1339 25113
rect 1403 25049 1433 25113
rect 1497 25049 1500 25113
rect 960 25032 1500 25049
rect 960 24968 963 25032
rect 1027 24968 1057 25032
rect 1121 24968 1151 25032
rect 1215 24968 1245 25032
rect 1309 24968 1339 25032
rect 1403 24968 1433 25032
rect 1497 24968 1500 25032
rect 960 24951 1500 24968
rect 960 24887 963 24951
rect 1027 24887 1057 24951
rect 1121 24887 1151 24951
rect 1215 24887 1245 24951
rect 1309 24887 1339 24951
rect 1403 24887 1433 24951
rect 1497 24887 1500 24951
rect 960 24886 1500 24887
rect 13842 26314 14016 26315
rect 13842 26250 13843 26314
rect 13907 26250 13951 26314
rect 14015 26250 14016 26314
rect 13842 26213 14016 26250
rect 13842 26149 13843 26213
rect 13907 26149 13951 26213
rect 14015 26149 14016 26213
rect 13842 26112 14016 26149
rect 13842 26048 13843 26112
rect 13907 26048 13951 26112
rect 14015 26048 14016 26112
rect 13842 26010 14016 26048
rect 13842 25946 13843 26010
rect 13907 25946 13951 26010
rect 14015 25946 14016 26010
rect 13842 25908 14016 25946
rect 13842 25844 13843 25908
rect 13907 25844 13951 25908
rect 14015 25844 14016 25908
rect 13842 25806 14016 25844
rect 13842 25742 13843 25806
rect 13907 25742 13951 25806
rect 14015 25742 14016 25806
rect 13842 25704 14016 25742
rect 13842 25640 13843 25704
rect 13907 25640 13951 25704
rect 14015 25640 14016 25704
rect 13842 25602 14016 25640
rect 13842 25538 13843 25602
rect 13907 25538 13951 25602
rect 14015 25538 14016 25602
rect 13842 25500 14016 25538
rect 13842 25436 13843 25500
rect 13907 25436 13951 25500
rect 14015 25436 14016 25500
rect 13842 25398 14016 25436
rect 13842 25334 13843 25398
rect 13907 25334 13951 25398
rect 14015 25334 14016 25398
rect 13842 25296 14016 25334
rect 13842 25232 13843 25296
rect 13907 25232 13951 25296
rect 14015 25232 14016 25296
rect 13842 25194 14016 25232
rect 13842 25130 13843 25194
rect 13907 25130 13951 25194
rect 14015 25130 14016 25194
rect 13842 25092 14016 25130
rect 13842 25028 13843 25092
rect 13907 25028 13951 25092
rect 14015 25028 14016 25092
rect 13842 24990 14016 25028
rect 13842 24926 13843 24990
rect 13907 24926 13951 24990
rect 14015 24926 14016 24990
rect 13842 24888 14016 24926
rect 13842 24824 13843 24888
rect 13907 24824 13951 24888
rect 14015 24824 14016 24888
rect 13842 24786 14016 24824
rect 13842 24722 13843 24786
rect 13907 24722 13951 24786
rect 14015 24722 14016 24786
rect 13842 24684 14016 24722
rect 13842 24620 13843 24684
rect 13907 24620 13951 24684
rect 14015 24620 14016 24684
rect 13842 24582 14016 24620
rect 13842 24518 13843 24582
rect 13907 24518 13951 24582
rect 14015 24518 14016 24582
rect 13842 24480 14016 24518
rect 13842 24416 13843 24480
rect 13907 24416 13951 24480
rect 14015 24416 14016 24480
rect 13842 24378 14016 24416
rect 13842 24314 13843 24378
rect 13907 24314 13951 24378
rect 14015 24314 14016 24378
rect 13842 24276 14016 24314
rect 13842 24212 13843 24276
rect 13907 24212 13951 24276
rect 14015 24212 14016 24276
rect 13842 24174 14016 24212
rect 13842 24110 13843 24174
rect 13907 24110 13951 24174
rect 14015 24110 14016 24174
rect 13842 24072 14016 24110
rect 13842 24008 13843 24072
rect 13907 24008 13951 24072
rect 14015 24008 14016 24072
rect 13842 23970 14016 24008
rect 13842 23906 13843 23970
rect 13907 23906 13951 23970
rect 14015 23906 14016 23970
rect 13842 23868 14016 23906
rect 13842 23804 13843 23868
rect 13907 23804 13951 23868
rect 14015 23804 14016 23868
rect 13842 23766 14016 23804
tri 1034 23702 1079 23747 se
tri 1018 23686 1034 23702 se
rect 1034 23686 1079 23702
rect 13842 23702 13843 23766
rect 13907 23702 13951 23766
rect 14015 23702 14016 23766
rect 1008 23685 1168 23686
tri 953 23621 1008 23676 se
rect 1008 23621 1009 23685
rect 1073 23621 1103 23685
rect 1167 23621 1168 23685
tri 936 23604 953 23621 se
rect 953 23604 1168 23621
tri 872 23540 936 23604 se
rect 936 23540 1009 23604
rect 1073 23540 1103 23604
rect 1167 23540 1168 23604
tri 854 23522 872 23540 se
rect 872 23522 1168 23540
tri 790 23458 854 23522 se
rect 854 23458 1009 23522
rect 1073 23458 1103 23522
rect 1167 23458 1168 23522
tri 772 23440 790 23458 se
rect 790 23440 1168 23458
tri 708 23376 772 23440 se
rect 772 23376 1009 23440
rect 1073 23376 1103 23440
rect 1167 23376 1168 23440
tri 700 23368 708 23376 se
rect 708 23368 1168 23376
rect 700 23358 1168 23368
rect 700 23294 1009 23358
rect 1073 23294 1103 23358
rect 1167 23294 1168 23358
rect 700 23276 1168 23294
rect 700 23212 1009 23276
rect 1073 23212 1103 23276
rect 1167 23212 1168 23276
rect 700 23194 1168 23212
rect 700 23130 1009 23194
rect 1073 23130 1103 23194
rect 1167 23130 1168 23194
rect 700 23112 1168 23130
rect 700 23048 1009 23112
rect 1073 23048 1103 23112
rect 1167 23048 1168 23112
rect 700 23030 1168 23048
rect 700 22966 1009 23030
rect 1073 22966 1103 23030
rect 1167 22966 1168 23030
rect 700 22948 1168 22966
rect 700 22884 1009 22948
rect 1073 22884 1103 22948
rect 1167 22884 1168 22948
rect 700 22866 1168 22884
rect 700 22802 1009 22866
rect 1073 22802 1103 22866
rect 1167 22802 1168 22866
rect 700 22784 1168 22802
rect 700 22720 1009 22784
rect 1073 22720 1103 22784
rect 1167 22720 1168 22784
rect 700 22702 1168 22720
rect 700 22638 1009 22702
rect 1073 22638 1103 22702
rect 1167 22638 1168 22702
rect 700 22620 1168 22638
rect 700 22556 1009 22620
rect 1073 22556 1103 22620
rect 1167 22556 1168 22620
rect 700 22538 1168 22556
rect 700 22474 1009 22538
rect 1073 22474 1103 22538
rect 1167 22474 1168 22538
rect 700 22456 1168 22474
rect 700 22392 1009 22456
rect 1073 22392 1103 22456
rect 1167 22392 1168 22456
rect 700 22374 1168 22392
rect 700 22310 1009 22374
rect 1073 22310 1103 22374
rect 1167 22310 1168 22374
rect 700 22292 1168 22310
rect 700 22228 1009 22292
rect 1073 22228 1103 22292
rect 1167 22228 1168 22292
rect 700 22210 1168 22228
rect 700 22146 1009 22210
rect 1073 22146 1103 22210
rect 1167 22146 1168 22210
rect 700 22128 1168 22146
rect 700 22064 1009 22128
rect 1073 22064 1103 22128
rect 1167 22064 1168 22128
rect 700 22046 1168 22064
rect 700 21982 1009 22046
rect 1073 21982 1103 22046
rect 1167 21982 1168 22046
rect 700 21964 1168 21982
rect 700 21900 1009 21964
rect 1073 21900 1103 21964
rect 1167 21900 1168 21964
rect 700 21882 1168 21900
rect 700 21818 1009 21882
rect 1073 21818 1103 21882
rect 1167 21818 1168 21882
rect 700 21817 1168 21818
rect 13842 23664 14016 23702
rect 13842 23600 13843 23664
rect 13907 23600 13951 23664
rect 14015 23600 14016 23664
rect 13842 23562 14016 23600
rect 13842 23498 13843 23562
rect 13907 23498 13951 23562
rect 14015 23498 14016 23562
rect 13842 23460 14016 23498
rect 13842 23396 13843 23460
rect 13907 23396 13951 23460
rect 14015 23396 14016 23460
rect 13842 23358 14016 23396
rect 13842 23294 13843 23358
rect 13907 23294 13951 23358
rect 14015 23294 14016 23358
rect 13842 23256 14016 23294
rect 13842 23192 13843 23256
rect 13907 23192 13951 23256
rect 14015 23192 14016 23256
rect 13842 23154 14016 23192
rect 13842 23090 13843 23154
rect 13907 23090 13951 23154
rect 14015 23090 14016 23154
rect 13842 23052 14016 23090
rect 13842 22988 13843 23052
rect 13907 22988 13951 23052
rect 14015 22988 14016 23052
rect 13842 22950 14016 22988
rect 13842 22886 13843 22950
rect 13907 22886 13951 22950
rect 14015 22886 14016 22950
rect 13842 22848 14016 22886
rect 13842 22784 13843 22848
rect 13907 22784 13951 22848
rect 14015 22784 14016 22848
rect 13842 22746 14016 22784
rect 13842 22682 13843 22746
rect 13907 22682 13951 22746
rect 14015 22682 14016 22746
rect 13842 22644 14016 22682
rect 13842 22580 13843 22644
rect 13907 22580 13951 22644
rect 14015 22580 14016 22644
rect 13842 22542 14016 22580
rect 13842 22478 13843 22542
rect 13907 22478 13951 22542
rect 14015 22478 14016 22542
rect 13842 22440 14016 22478
rect 13842 22376 13843 22440
rect 13907 22376 13951 22440
rect 14015 22376 14016 22440
rect 13842 22338 14016 22376
rect 13842 22274 13843 22338
rect 13907 22274 13951 22338
rect 14015 22274 14016 22338
rect 13842 22236 14016 22274
rect 13842 22172 13843 22236
rect 13907 22172 13951 22236
rect 14015 22172 14016 22236
rect 13842 22134 14016 22172
rect 13842 22070 13843 22134
rect 13907 22070 13951 22134
rect 14015 22070 14016 22134
rect 13842 22032 14016 22070
rect 13842 21968 13843 22032
rect 13907 21968 13951 22032
rect 14015 21968 14016 22032
rect 13842 21930 14016 21968
rect 13842 21866 13843 21930
rect 13907 21866 13951 21930
rect 14015 21866 14016 21930
rect 13842 21828 14016 21866
rect 700 20706 1079 21817
rect 13842 21764 13843 21828
rect 13907 21764 13951 21828
rect 14015 21764 14016 21828
rect 13842 21726 14016 21764
rect 13842 21662 13843 21726
rect 13907 21662 13951 21726
rect 14015 21662 14016 21726
rect 13842 21624 14016 21662
rect 13842 21560 13843 21624
rect 13907 21560 13951 21624
rect 14015 21560 14016 21624
rect 13842 21559 14016 21560
tri 700 20327 1079 20706 ne
rect 12899 20054 13085 20055
rect 1985 19990 2167 19991
rect 1985 19926 1986 19990
rect 2050 19926 2102 19990
rect 2166 19926 2167 19990
rect 1985 19907 2167 19926
rect 1985 19843 1986 19907
rect 2050 19843 2102 19907
rect 2166 19843 2167 19907
rect 1985 19823 2167 19843
rect 1985 19759 1986 19823
rect 2050 19759 2102 19823
rect 2166 19759 2167 19823
rect 1985 19739 2167 19759
rect 1985 19675 1986 19739
rect 2050 19675 2102 19739
rect 2166 19675 2167 19739
rect 1985 19655 2167 19675
rect 12899 19990 12900 20054
rect 12964 19990 13020 20054
rect 13084 19990 13085 20054
rect 12899 19962 13085 19990
rect 12899 19898 12900 19962
rect 12964 19898 13020 19962
rect 13084 19898 13085 19962
rect 12899 19870 13085 19898
rect 12899 19806 12900 19870
rect 12964 19806 13020 19870
rect 13084 19806 13085 19870
rect 12899 19778 13085 19806
rect 12899 19714 12900 19778
rect 12964 19714 13020 19778
rect 13084 19714 13085 19778
rect 12899 19686 13085 19714
rect 1985 19591 1986 19655
rect 2050 19591 2102 19655
rect 2166 19591 2167 19655
rect 1985 19571 2167 19591
rect 1985 19507 1986 19571
rect 2050 19507 2102 19571
rect 2166 19507 2167 19571
rect 1985 19487 2167 19507
rect 1985 19423 1986 19487
rect 2050 19423 2102 19487
rect 2166 19423 2167 19487
rect 1985 19422 2167 19423
rect 2979 19673 3165 19674
rect 2979 19609 2980 19673
rect 3044 19609 3100 19673
rect 3164 19609 3165 19673
rect 2979 19581 3165 19609
rect 2979 19517 2980 19581
rect 3044 19517 3100 19581
rect 3164 19517 3165 19581
rect 2979 19489 3165 19517
rect 2979 19425 2980 19489
rect 3044 19425 3100 19489
rect 3164 19425 3165 19489
rect 2979 19397 3165 19425
rect 2979 19333 2980 19397
rect 3044 19333 3100 19397
rect 3164 19333 3165 19397
rect 2979 19305 3165 19333
rect 2979 19241 2980 19305
rect 3044 19241 3100 19305
rect 3164 19241 3165 19305
rect 2979 19212 3165 19241
rect 2979 19148 2980 19212
rect 3044 19148 3100 19212
rect 3164 19148 3165 19212
rect 2979 19147 3165 19148
rect 3971 19673 4157 19674
rect 3971 19609 3972 19673
rect 4036 19609 4092 19673
rect 4156 19609 4157 19673
rect 3971 19581 4157 19609
rect 3971 19517 3972 19581
rect 4036 19517 4092 19581
rect 4156 19517 4157 19581
rect 3971 19488 4157 19517
rect 3971 19424 3972 19488
rect 4036 19424 4092 19488
rect 4156 19424 4157 19488
rect 3971 19395 4157 19424
rect 3971 19331 3972 19395
rect 4036 19331 4092 19395
rect 4156 19331 4157 19395
rect 3971 19302 4157 19331
rect 3971 19238 3972 19302
rect 4036 19238 4092 19302
rect 4156 19238 4157 19302
rect 3971 19209 4157 19238
rect 3971 19145 3972 19209
rect 4036 19145 4092 19209
rect 4156 19145 4157 19209
rect 4963 19673 5149 19674
rect 4963 19609 4964 19673
rect 5028 19609 5084 19673
rect 5148 19609 5149 19673
rect 4963 19581 5149 19609
rect 4963 19517 4964 19581
rect 5028 19517 5084 19581
rect 5148 19517 5149 19581
rect 4963 19489 5149 19517
rect 4963 19425 4964 19489
rect 5028 19425 5084 19489
rect 5148 19425 5149 19489
rect 4963 19397 5149 19425
rect 4963 19333 4964 19397
rect 5028 19333 5084 19397
rect 5148 19333 5149 19397
rect 4963 19305 5149 19333
rect 4963 19241 4964 19305
rect 5028 19241 5084 19305
rect 5148 19241 5149 19305
rect 4963 19212 5149 19241
rect 4963 19148 4964 19212
rect 5028 19148 5084 19212
rect 5148 19148 5149 19212
rect 4963 19147 5149 19148
rect 5952 19673 6138 19674
rect 5952 19609 5953 19673
rect 6017 19609 6073 19673
rect 6137 19609 6138 19673
rect 5952 19581 6138 19609
rect 5952 19517 5953 19581
rect 6017 19517 6073 19581
rect 6137 19517 6138 19581
rect 5952 19489 6138 19517
rect 5952 19425 5953 19489
rect 6017 19425 6073 19489
rect 6137 19425 6138 19489
rect 5952 19397 6138 19425
rect 5952 19333 5953 19397
rect 6017 19333 6073 19397
rect 6137 19333 6138 19397
rect 5952 19305 6138 19333
rect 5952 19241 5953 19305
rect 6017 19241 6073 19305
rect 6137 19241 6138 19305
rect 5952 19212 6138 19241
rect 5952 19148 5953 19212
rect 6017 19148 6073 19212
rect 6137 19148 6138 19212
rect 5952 19147 6138 19148
rect 6944 19673 7130 19674
rect 6944 19609 6945 19673
rect 7009 19609 7065 19673
rect 7129 19609 7130 19673
rect 6944 19581 7130 19609
rect 6944 19517 6945 19581
rect 7009 19517 7065 19581
rect 7129 19517 7130 19581
rect 6944 19489 7130 19517
rect 6944 19425 6945 19489
rect 7009 19425 7065 19489
rect 7129 19425 7130 19489
rect 6944 19397 7130 19425
rect 6944 19333 6945 19397
rect 7009 19333 7065 19397
rect 7129 19333 7130 19397
rect 6944 19305 7130 19333
rect 6944 19241 6945 19305
rect 7009 19241 7065 19305
rect 7129 19241 7130 19305
rect 6944 19212 7130 19241
rect 6944 19148 6945 19212
rect 7009 19148 7065 19212
rect 7129 19148 7130 19212
rect 6944 19147 7130 19148
rect 7939 19673 8125 19674
rect 7939 19609 7940 19673
rect 8004 19609 8060 19673
rect 8124 19609 8125 19673
rect 7939 19581 8125 19609
rect 7939 19517 7940 19581
rect 8004 19517 8060 19581
rect 8124 19517 8125 19581
rect 7939 19489 8125 19517
rect 7939 19425 7940 19489
rect 8004 19425 8060 19489
rect 8124 19425 8125 19489
rect 7939 19397 8125 19425
rect 7939 19333 7940 19397
rect 8004 19333 8060 19397
rect 8124 19333 8125 19397
rect 7939 19305 8125 19333
rect 7939 19241 7940 19305
rect 8004 19241 8060 19305
rect 8124 19241 8125 19305
rect 7939 19212 8125 19241
rect 7939 19148 7940 19212
rect 8004 19148 8060 19212
rect 8124 19148 8125 19212
rect 7939 19147 8125 19148
rect 8931 19673 9117 19674
rect 8931 19609 8932 19673
rect 8996 19609 9052 19673
rect 9116 19609 9117 19673
rect 8931 19581 9117 19609
rect 8931 19517 8932 19581
rect 8996 19517 9052 19581
rect 9116 19517 9117 19581
rect 8931 19489 9117 19517
rect 8931 19425 8932 19489
rect 8996 19425 9052 19489
rect 9116 19425 9117 19489
rect 8931 19397 9117 19425
rect 8931 19333 8932 19397
rect 8996 19333 9052 19397
rect 9116 19333 9117 19397
rect 8931 19305 9117 19333
rect 8931 19241 8932 19305
rect 8996 19241 9052 19305
rect 9116 19241 9117 19305
rect 8931 19212 9117 19241
rect 8931 19148 8932 19212
rect 8996 19148 9052 19212
rect 9116 19148 9117 19212
rect 8931 19147 9117 19148
rect 9923 19673 10109 19674
rect 9923 19609 9924 19673
rect 9988 19609 10044 19673
rect 10108 19609 10109 19673
rect 9923 19581 10109 19609
rect 9923 19517 9924 19581
rect 9988 19517 10044 19581
rect 10108 19517 10109 19581
rect 9923 19489 10109 19517
rect 9923 19425 9924 19489
rect 9988 19425 10044 19489
rect 10108 19425 10109 19489
rect 9923 19397 10109 19425
rect 9923 19333 9924 19397
rect 9988 19333 10044 19397
rect 10108 19333 10109 19397
rect 9923 19305 10109 19333
rect 9923 19241 9924 19305
rect 9988 19241 10044 19305
rect 10108 19241 10109 19305
rect 9923 19212 10109 19241
rect 9923 19148 9924 19212
rect 9988 19148 10044 19212
rect 10108 19148 10109 19212
rect 9923 19147 10109 19148
rect 10915 19673 11101 19674
rect 10915 19609 10916 19673
rect 10980 19609 11036 19673
rect 11100 19609 11101 19673
rect 10915 19581 11101 19609
rect 10915 19517 10916 19581
rect 10980 19517 11036 19581
rect 11100 19517 11101 19581
rect 10915 19489 11101 19517
rect 10915 19425 10916 19489
rect 10980 19425 11036 19489
rect 11100 19425 11101 19489
rect 10915 19397 11101 19425
rect 10915 19333 10916 19397
rect 10980 19333 11036 19397
rect 11100 19333 11101 19397
rect 10915 19305 11101 19333
rect 10915 19241 10916 19305
rect 10980 19241 11036 19305
rect 11100 19241 11101 19305
rect 10915 19212 11101 19241
rect 10915 19148 10916 19212
rect 10980 19148 11036 19212
rect 11100 19148 11101 19212
rect 10915 19147 11101 19148
rect 11907 19673 12093 19674
rect 11907 19609 11908 19673
rect 11972 19609 12028 19673
rect 12092 19609 12093 19673
rect 11907 19581 12093 19609
rect 11907 19517 11908 19581
rect 11972 19517 12028 19581
rect 12092 19517 12093 19581
rect 12899 19622 12900 19686
rect 12964 19622 13020 19686
rect 13084 19622 13085 19686
rect 12899 19593 13085 19622
rect 12899 19529 12900 19593
rect 12964 19529 13020 19593
rect 13084 19529 13085 19593
rect 12899 19528 13085 19529
rect 11907 19489 12093 19517
rect 11907 19425 11908 19489
rect 11972 19425 12028 19489
rect 12092 19425 12093 19489
rect 11907 19397 12093 19425
rect 11907 19333 11908 19397
rect 11972 19333 12028 19397
rect 12092 19333 12093 19397
rect 11907 19305 12093 19333
rect 11907 19241 11908 19305
rect 11972 19241 12028 19305
rect 12092 19241 12093 19305
rect 11907 19212 12093 19241
rect 11907 19148 11908 19212
rect 11972 19148 12028 19212
rect 12092 19148 12093 19212
rect 11907 19147 12093 19148
rect 3971 19144 4157 19145
rect 0 18592 15000 18600
rect 0 18588 2480 18592
rect 0 15484 456 18588
rect 1160 18586 2480 18588
rect 1160 18522 1287 18586
rect 1351 18522 1375 18586
rect 1439 18522 1463 18586
rect 1527 18522 1551 18586
rect 1615 18522 1639 18586
rect 1703 18522 1727 18586
rect 1791 18522 1815 18586
rect 1879 18528 2480 18586
rect 2544 18528 2608 18592
rect 2672 18528 3472 18592
rect 3536 18528 3600 18592
rect 3664 18528 4464 18592
rect 4528 18528 4592 18592
rect 4656 18528 5456 18592
rect 5520 18528 5584 18592
rect 5648 18528 6448 18592
rect 6512 18528 6576 18592
rect 6640 18528 7440 18592
rect 7504 18528 7568 18592
rect 7632 18528 8432 18592
rect 8496 18528 8560 18592
rect 8624 18528 9424 18592
rect 9488 18528 9552 18592
rect 9616 18528 10416 18592
rect 10480 18528 10544 18592
rect 10608 18528 11408 18592
rect 11472 18528 11536 18592
rect 11600 18528 12400 18592
rect 12464 18528 12528 18592
rect 12592 18528 13392 18592
rect 13456 18528 13520 18592
rect 13584 18590 15000 18592
rect 13584 18528 13777 18590
rect 1879 18526 13777 18528
rect 13841 18526 13863 18590
rect 13927 18526 13949 18590
rect 14013 18526 14035 18590
rect 14099 18526 14121 18590
rect 14185 18526 14207 18590
rect 14271 18526 14293 18590
rect 14357 18526 14379 18590
rect 14443 18526 14465 18590
rect 14529 18526 15000 18590
rect 1879 18522 15000 18526
rect 1160 18512 15000 18522
rect 1160 18506 2480 18512
rect 1160 18442 1287 18506
rect 1351 18442 1375 18506
rect 1439 18442 1463 18506
rect 1527 18442 1551 18506
rect 1615 18442 1639 18506
rect 1703 18442 1727 18506
rect 1791 18442 1815 18506
rect 1879 18448 2480 18506
rect 2544 18448 2608 18512
rect 2672 18448 3472 18512
rect 3536 18448 3600 18512
rect 3664 18448 4464 18512
rect 4528 18448 4592 18512
rect 4656 18448 5456 18512
rect 5520 18448 5584 18512
rect 5648 18448 6448 18512
rect 6512 18448 6576 18512
rect 6640 18448 7440 18512
rect 7504 18448 7568 18512
rect 7632 18448 8432 18512
rect 8496 18448 8560 18512
rect 8624 18448 9424 18512
rect 9488 18448 9552 18512
rect 9616 18448 10416 18512
rect 10480 18448 10544 18512
rect 10608 18448 11408 18512
rect 11472 18448 11536 18512
rect 11600 18448 12400 18512
rect 12464 18448 12528 18512
rect 12592 18448 13392 18512
rect 13456 18448 13520 18512
rect 13584 18510 15000 18512
rect 13584 18448 13777 18510
rect 1879 18446 13777 18448
rect 13841 18446 13863 18510
rect 13927 18446 13949 18510
rect 14013 18446 14035 18510
rect 14099 18446 14121 18510
rect 14185 18446 14207 18510
rect 14271 18446 14293 18510
rect 14357 18446 14379 18510
rect 14443 18446 14465 18510
rect 14529 18446 15000 18510
rect 1879 18442 15000 18446
rect 1160 18432 15000 18442
rect 1160 18426 2480 18432
rect 1160 18362 1287 18426
rect 1351 18362 1375 18426
rect 1439 18362 1463 18426
rect 1527 18362 1551 18426
rect 1615 18362 1639 18426
rect 1703 18362 1727 18426
rect 1791 18362 1815 18426
rect 1879 18368 2480 18426
rect 2544 18368 2608 18432
rect 2672 18368 3472 18432
rect 3536 18368 3600 18432
rect 3664 18368 4464 18432
rect 4528 18368 4592 18432
rect 4656 18368 5456 18432
rect 5520 18368 5584 18432
rect 5648 18368 6448 18432
rect 6512 18368 6576 18432
rect 6640 18368 7440 18432
rect 7504 18368 7568 18432
rect 7632 18368 8432 18432
rect 8496 18368 8560 18432
rect 8624 18368 9424 18432
rect 9488 18368 9552 18432
rect 9616 18368 10416 18432
rect 10480 18368 10544 18432
rect 10608 18368 11408 18432
rect 11472 18368 11536 18432
rect 11600 18368 12400 18432
rect 12464 18368 12528 18432
rect 12592 18368 13392 18432
rect 13456 18368 13520 18432
rect 13584 18430 15000 18432
rect 13584 18368 13777 18430
rect 1879 18366 13777 18368
rect 13841 18366 13863 18430
rect 13927 18366 13949 18430
rect 14013 18366 14035 18430
rect 14099 18366 14121 18430
rect 14185 18366 14207 18430
rect 14271 18366 14293 18430
rect 14357 18366 14379 18430
rect 14443 18366 14465 18430
rect 14529 18366 15000 18430
rect 1879 18362 15000 18366
rect 1160 18352 15000 18362
rect 1160 18346 2480 18352
rect 1160 18282 1287 18346
rect 1351 18282 1375 18346
rect 1439 18282 1463 18346
rect 1527 18282 1551 18346
rect 1615 18282 1639 18346
rect 1703 18282 1727 18346
rect 1791 18282 1815 18346
rect 1879 18288 2480 18346
rect 2544 18288 2608 18352
rect 2672 18288 3472 18352
rect 3536 18288 3600 18352
rect 3664 18288 4464 18352
rect 4528 18288 4592 18352
rect 4656 18288 5456 18352
rect 5520 18288 5584 18352
rect 5648 18288 6448 18352
rect 6512 18288 6576 18352
rect 6640 18288 7440 18352
rect 7504 18288 7568 18352
rect 7632 18288 8432 18352
rect 8496 18288 8560 18352
rect 8624 18288 9424 18352
rect 9488 18288 9552 18352
rect 9616 18288 10416 18352
rect 10480 18288 10544 18352
rect 10608 18288 11408 18352
rect 11472 18288 11536 18352
rect 11600 18288 12400 18352
rect 12464 18288 12528 18352
rect 12592 18288 13392 18352
rect 13456 18288 13520 18352
rect 13584 18350 15000 18352
rect 13584 18288 13777 18350
rect 1879 18286 13777 18288
rect 13841 18286 13863 18350
rect 13927 18286 13949 18350
rect 14013 18286 14035 18350
rect 14099 18286 14121 18350
rect 14185 18286 14207 18350
rect 14271 18286 14293 18350
rect 14357 18286 14379 18350
rect 14443 18286 14465 18350
rect 14529 18286 15000 18350
rect 1879 18282 15000 18286
rect 1160 18272 15000 18282
rect 1160 18266 2480 18272
rect 1160 18202 1287 18266
rect 1351 18202 1375 18266
rect 1439 18202 1463 18266
rect 1527 18202 1551 18266
rect 1615 18202 1639 18266
rect 1703 18202 1727 18266
rect 1791 18202 1815 18266
rect 1879 18208 2480 18266
rect 2544 18208 2608 18272
rect 2672 18208 3472 18272
rect 3536 18208 3600 18272
rect 3664 18208 4464 18272
rect 4528 18208 4592 18272
rect 4656 18208 5456 18272
rect 5520 18208 5584 18272
rect 5648 18208 6448 18272
rect 6512 18208 6576 18272
rect 6640 18208 7440 18272
rect 7504 18208 7568 18272
rect 7632 18208 8432 18272
rect 8496 18208 8560 18272
rect 8624 18208 9424 18272
rect 9488 18208 9552 18272
rect 9616 18208 10416 18272
rect 10480 18208 10544 18272
rect 10608 18208 11408 18272
rect 11472 18208 11536 18272
rect 11600 18208 12400 18272
rect 12464 18208 12528 18272
rect 12592 18208 13392 18272
rect 13456 18208 13520 18272
rect 13584 18270 15000 18272
rect 13584 18208 13777 18270
rect 1879 18206 13777 18208
rect 13841 18206 13863 18270
rect 13927 18206 13949 18270
rect 14013 18206 14035 18270
rect 14099 18206 14121 18270
rect 14185 18206 14207 18270
rect 14271 18206 14293 18270
rect 14357 18206 14379 18270
rect 14443 18206 14465 18270
rect 14529 18206 15000 18270
rect 1879 18202 15000 18206
rect 1160 18192 15000 18202
rect 1160 18186 2480 18192
rect 1160 18122 1287 18186
rect 1351 18122 1375 18186
rect 1439 18122 1463 18186
rect 1527 18122 1551 18186
rect 1615 18122 1639 18186
rect 1703 18122 1727 18186
rect 1791 18122 1815 18186
rect 1879 18128 2480 18186
rect 2544 18128 2608 18192
rect 2672 18128 3472 18192
rect 3536 18128 3600 18192
rect 3664 18128 4464 18192
rect 4528 18128 4592 18192
rect 4656 18128 5456 18192
rect 5520 18128 5584 18192
rect 5648 18128 6448 18192
rect 6512 18128 6576 18192
rect 6640 18128 7440 18192
rect 7504 18128 7568 18192
rect 7632 18128 8432 18192
rect 8496 18128 8560 18192
rect 8624 18128 9424 18192
rect 9488 18128 9552 18192
rect 9616 18128 10416 18192
rect 10480 18128 10544 18192
rect 10608 18128 11408 18192
rect 11472 18128 11536 18192
rect 11600 18128 12400 18192
rect 12464 18128 12528 18192
rect 12592 18128 13392 18192
rect 13456 18128 13520 18192
rect 13584 18190 15000 18192
rect 13584 18128 13777 18190
rect 1879 18126 13777 18128
rect 13841 18126 13863 18190
rect 13927 18126 13949 18190
rect 14013 18126 14035 18190
rect 14099 18126 14121 18190
rect 14185 18126 14207 18190
rect 14271 18126 14293 18190
rect 14357 18126 14379 18190
rect 14443 18126 14465 18190
rect 14529 18126 15000 18190
rect 1879 18122 15000 18126
rect 1160 18112 15000 18122
rect 1160 18106 2480 18112
rect 1160 18042 1287 18106
rect 1351 18042 1375 18106
rect 1439 18042 1463 18106
rect 1527 18042 1551 18106
rect 1615 18042 1639 18106
rect 1703 18042 1727 18106
rect 1791 18042 1815 18106
rect 1879 18048 2480 18106
rect 2544 18048 2608 18112
rect 2672 18048 3472 18112
rect 3536 18048 3600 18112
rect 3664 18048 4464 18112
rect 4528 18048 4592 18112
rect 4656 18048 5456 18112
rect 5520 18048 5584 18112
rect 5648 18048 6448 18112
rect 6512 18048 6576 18112
rect 6640 18048 7440 18112
rect 7504 18048 7568 18112
rect 7632 18048 8432 18112
rect 8496 18048 8560 18112
rect 8624 18048 9424 18112
rect 9488 18048 9552 18112
rect 9616 18048 10416 18112
rect 10480 18048 10544 18112
rect 10608 18048 11408 18112
rect 11472 18048 11536 18112
rect 11600 18048 12400 18112
rect 12464 18048 12528 18112
rect 12592 18048 13392 18112
rect 13456 18048 13520 18112
rect 13584 18110 15000 18112
rect 13584 18048 13777 18110
rect 1879 18046 13777 18048
rect 13841 18046 13863 18110
rect 13927 18046 13949 18110
rect 14013 18046 14035 18110
rect 14099 18046 14121 18110
rect 14185 18046 14207 18110
rect 14271 18046 14293 18110
rect 14357 18046 14379 18110
rect 14443 18046 14465 18110
rect 14529 18046 15000 18110
rect 1879 18042 15000 18046
rect 1160 18032 15000 18042
rect 1160 18026 2480 18032
rect 1160 17962 1287 18026
rect 1351 17962 1375 18026
rect 1439 17962 1463 18026
rect 1527 17962 1551 18026
rect 1615 17962 1639 18026
rect 1703 17962 1727 18026
rect 1791 17962 1815 18026
rect 1879 17968 2480 18026
rect 2544 17968 2608 18032
rect 2672 17968 3472 18032
rect 3536 17968 3600 18032
rect 3664 17968 4464 18032
rect 4528 17968 4592 18032
rect 4656 17968 5456 18032
rect 5520 17968 5584 18032
rect 5648 17968 6448 18032
rect 6512 17968 6576 18032
rect 6640 17968 7440 18032
rect 7504 17968 7568 18032
rect 7632 17968 8432 18032
rect 8496 17968 8560 18032
rect 8624 17968 9424 18032
rect 9488 17968 9552 18032
rect 9616 17968 10416 18032
rect 10480 17968 10544 18032
rect 10608 17968 11408 18032
rect 11472 17968 11536 18032
rect 11600 17968 12400 18032
rect 12464 17968 12528 18032
rect 12592 17968 13392 18032
rect 13456 17968 13520 18032
rect 13584 18030 15000 18032
rect 13584 17968 13777 18030
rect 1879 17966 13777 17968
rect 13841 17966 13863 18030
rect 13927 17966 13949 18030
rect 14013 17966 14035 18030
rect 14099 17966 14121 18030
rect 14185 17966 14207 18030
rect 14271 17966 14293 18030
rect 14357 17966 14379 18030
rect 14443 17966 14465 18030
rect 14529 17966 15000 18030
rect 1879 17962 15000 17966
rect 1160 17952 15000 17962
rect 1160 17946 2480 17952
rect 1160 17882 1287 17946
rect 1351 17882 1375 17946
rect 1439 17882 1463 17946
rect 1527 17882 1551 17946
rect 1615 17882 1639 17946
rect 1703 17882 1727 17946
rect 1791 17882 1815 17946
rect 1879 17888 2480 17946
rect 2544 17888 2608 17952
rect 2672 17888 3472 17952
rect 3536 17888 3600 17952
rect 3664 17888 4464 17952
rect 4528 17888 4592 17952
rect 4656 17888 5456 17952
rect 5520 17888 5584 17952
rect 5648 17888 6448 17952
rect 6512 17888 6576 17952
rect 6640 17888 7440 17952
rect 7504 17888 7568 17952
rect 7632 17888 8432 17952
rect 8496 17888 8560 17952
rect 8624 17888 9424 17952
rect 9488 17888 9552 17952
rect 9616 17888 10416 17952
rect 10480 17888 10544 17952
rect 10608 17888 11408 17952
rect 11472 17888 11536 17952
rect 11600 17888 12400 17952
rect 12464 17888 12528 17952
rect 12592 17888 13392 17952
rect 13456 17888 13520 17952
rect 13584 17950 15000 17952
rect 13584 17888 13777 17950
rect 1879 17886 13777 17888
rect 13841 17886 13863 17950
rect 13927 17886 13949 17950
rect 14013 17886 14035 17950
rect 14099 17886 14121 17950
rect 14185 17886 14207 17950
rect 14271 17886 14293 17950
rect 14357 17886 14379 17950
rect 14443 17886 14465 17950
rect 14529 17886 15000 17950
rect 1879 17882 15000 17886
rect 1160 17872 15000 17882
rect 1160 17866 2480 17872
rect 1160 17802 1287 17866
rect 1351 17802 1375 17866
rect 1439 17802 1463 17866
rect 1527 17802 1551 17866
rect 1615 17802 1639 17866
rect 1703 17802 1727 17866
rect 1791 17802 1815 17866
rect 1879 17808 2480 17866
rect 2544 17808 2608 17872
rect 2672 17808 3472 17872
rect 3536 17808 3600 17872
rect 3664 17808 4464 17872
rect 4528 17808 4592 17872
rect 4656 17808 5456 17872
rect 5520 17808 5584 17872
rect 5648 17808 6448 17872
rect 6512 17808 6576 17872
rect 6640 17808 7440 17872
rect 7504 17808 7568 17872
rect 7632 17808 8432 17872
rect 8496 17808 8560 17872
rect 8624 17808 9424 17872
rect 9488 17808 9552 17872
rect 9616 17808 10416 17872
rect 10480 17808 10544 17872
rect 10608 17808 11408 17872
rect 11472 17808 11536 17872
rect 11600 17808 12400 17872
rect 12464 17808 12528 17872
rect 12592 17808 13392 17872
rect 13456 17808 13520 17872
rect 13584 17870 15000 17872
rect 13584 17808 13777 17870
rect 1879 17806 13777 17808
rect 13841 17806 13863 17870
rect 13927 17806 13949 17870
rect 14013 17806 14035 17870
rect 14099 17806 14121 17870
rect 14185 17806 14207 17870
rect 14271 17806 14293 17870
rect 14357 17806 14379 17870
rect 14443 17806 14465 17870
rect 14529 17806 15000 17870
rect 1879 17802 15000 17806
rect 1160 17792 15000 17802
rect 1160 17786 2480 17792
rect 1160 17722 1287 17786
rect 1351 17722 1375 17786
rect 1439 17722 1463 17786
rect 1527 17722 1551 17786
rect 1615 17722 1639 17786
rect 1703 17722 1727 17786
rect 1791 17722 1815 17786
rect 1879 17728 2480 17786
rect 2544 17728 2608 17792
rect 2672 17728 3472 17792
rect 3536 17728 3600 17792
rect 3664 17728 4464 17792
rect 4528 17728 4592 17792
rect 4656 17728 5456 17792
rect 5520 17728 5584 17792
rect 5648 17728 6448 17792
rect 6512 17728 6576 17792
rect 6640 17728 7440 17792
rect 7504 17728 7568 17792
rect 7632 17728 8432 17792
rect 8496 17728 8560 17792
rect 8624 17728 9424 17792
rect 9488 17728 9552 17792
rect 9616 17728 10416 17792
rect 10480 17728 10544 17792
rect 10608 17728 11408 17792
rect 11472 17728 11536 17792
rect 11600 17728 12400 17792
rect 12464 17728 12528 17792
rect 12592 17728 13392 17792
rect 13456 17728 13520 17792
rect 13584 17790 15000 17792
rect 13584 17728 13777 17790
rect 1879 17726 13777 17728
rect 13841 17726 13863 17790
rect 13927 17726 13949 17790
rect 14013 17726 14035 17790
rect 14099 17726 14121 17790
rect 14185 17726 14207 17790
rect 14271 17726 14293 17790
rect 14357 17726 14379 17790
rect 14443 17726 14465 17790
rect 14529 17726 15000 17790
rect 1879 17722 15000 17726
rect 1160 17712 15000 17722
rect 1160 17706 2480 17712
rect 1160 17642 1287 17706
rect 1351 17642 1375 17706
rect 1439 17642 1463 17706
rect 1527 17642 1551 17706
rect 1615 17642 1639 17706
rect 1703 17642 1727 17706
rect 1791 17642 1815 17706
rect 1879 17648 2480 17706
rect 2544 17648 2608 17712
rect 2672 17648 3472 17712
rect 3536 17648 3600 17712
rect 3664 17648 4464 17712
rect 4528 17648 4592 17712
rect 4656 17648 5456 17712
rect 5520 17648 5584 17712
rect 5648 17648 6448 17712
rect 6512 17648 6576 17712
rect 6640 17648 7440 17712
rect 7504 17648 7568 17712
rect 7632 17648 8432 17712
rect 8496 17648 8560 17712
rect 8624 17648 9424 17712
rect 9488 17648 9552 17712
rect 9616 17648 10416 17712
rect 10480 17648 10544 17712
rect 10608 17648 11408 17712
rect 11472 17648 11536 17712
rect 11600 17648 12400 17712
rect 12464 17648 12528 17712
rect 12592 17648 13392 17712
rect 13456 17648 13520 17712
rect 13584 17710 15000 17712
rect 13584 17648 13777 17710
rect 1879 17646 13777 17648
rect 13841 17646 13863 17710
rect 13927 17646 13949 17710
rect 14013 17646 14035 17710
rect 14099 17646 14121 17710
rect 14185 17646 14207 17710
rect 14271 17646 14293 17710
rect 14357 17646 14379 17710
rect 14443 17646 14465 17710
rect 14529 17646 15000 17710
rect 1879 17642 15000 17646
rect 1160 17632 15000 17642
rect 1160 17626 2480 17632
rect 1160 17562 1287 17626
rect 1351 17562 1375 17626
rect 1439 17562 1463 17626
rect 1527 17562 1551 17626
rect 1615 17562 1639 17626
rect 1703 17562 1727 17626
rect 1791 17562 1815 17626
rect 1879 17568 2480 17626
rect 2544 17568 2608 17632
rect 2672 17568 3472 17632
rect 3536 17568 3600 17632
rect 3664 17568 4464 17632
rect 4528 17568 4592 17632
rect 4656 17568 5456 17632
rect 5520 17568 5584 17632
rect 5648 17568 6448 17632
rect 6512 17568 6576 17632
rect 6640 17568 7440 17632
rect 7504 17568 7568 17632
rect 7632 17568 8432 17632
rect 8496 17568 8560 17632
rect 8624 17568 9424 17632
rect 9488 17568 9552 17632
rect 9616 17568 10416 17632
rect 10480 17568 10544 17632
rect 10608 17568 11408 17632
rect 11472 17568 11536 17632
rect 11600 17568 12400 17632
rect 12464 17568 12528 17632
rect 12592 17568 13392 17632
rect 13456 17568 13520 17632
rect 13584 17630 15000 17632
rect 13584 17568 13777 17630
rect 1879 17566 13777 17568
rect 13841 17566 13863 17630
rect 13927 17566 13949 17630
rect 14013 17566 14035 17630
rect 14099 17566 14121 17630
rect 14185 17566 14207 17630
rect 14271 17566 14293 17630
rect 14357 17566 14379 17630
rect 14443 17566 14465 17630
rect 14529 17566 15000 17630
rect 1879 17562 15000 17566
rect 1160 17552 15000 17562
rect 1160 17546 2480 17552
rect 1160 17482 1287 17546
rect 1351 17482 1375 17546
rect 1439 17482 1463 17546
rect 1527 17482 1551 17546
rect 1615 17482 1639 17546
rect 1703 17482 1727 17546
rect 1791 17482 1815 17546
rect 1879 17488 2480 17546
rect 2544 17488 2608 17552
rect 2672 17488 3472 17552
rect 3536 17488 3600 17552
rect 3664 17488 4464 17552
rect 4528 17488 4592 17552
rect 4656 17488 5456 17552
rect 5520 17488 5584 17552
rect 5648 17488 6448 17552
rect 6512 17488 6576 17552
rect 6640 17488 7440 17552
rect 7504 17488 7568 17552
rect 7632 17488 8432 17552
rect 8496 17488 8560 17552
rect 8624 17488 9424 17552
rect 9488 17488 9552 17552
rect 9616 17488 10416 17552
rect 10480 17488 10544 17552
rect 10608 17488 11408 17552
rect 11472 17488 11536 17552
rect 11600 17488 12400 17552
rect 12464 17488 12528 17552
rect 12592 17488 13392 17552
rect 13456 17488 13520 17552
rect 13584 17550 15000 17552
rect 13584 17488 13777 17550
rect 1879 17486 13777 17488
rect 13841 17486 13863 17550
rect 13927 17486 13949 17550
rect 14013 17486 14035 17550
rect 14099 17486 14121 17550
rect 14185 17486 14207 17550
rect 14271 17486 14293 17550
rect 14357 17486 14379 17550
rect 14443 17486 14465 17550
rect 14529 17486 15000 17550
rect 1879 17482 15000 17486
rect 1160 17472 15000 17482
rect 1160 17466 2480 17472
rect 1160 17402 1287 17466
rect 1351 17402 1375 17466
rect 1439 17402 1463 17466
rect 1527 17402 1551 17466
rect 1615 17402 1639 17466
rect 1703 17402 1727 17466
rect 1791 17402 1815 17466
rect 1879 17408 2480 17466
rect 2544 17408 2608 17472
rect 2672 17408 3472 17472
rect 3536 17408 3600 17472
rect 3664 17408 4464 17472
rect 4528 17408 4592 17472
rect 4656 17408 5456 17472
rect 5520 17408 5584 17472
rect 5648 17408 6448 17472
rect 6512 17408 6576 17472
rect 6640 17408 7440 17472
rect 7504 17408 7568 17472
rect 7632 17408 8432 17472
rect 8496 17408 8560 17472
rect 8624 17408 9424 17472
rect 9488 17408 9552 17472
rect 9616 17408 10416 17472
rect 10480 17408 10544 17472
rect 10608 17408 11408 17472
rect 11472 17408 11536 17472
rect 11600 17408 12400 17472
rect 12464 17408 12528 17472
rect 12592 17408 13392 17472
rect 13456 17408 13520 17472
rect 13584 17470 15000 17472
rect 13584 17408 13777 17470
rect 1879 17406 13777 17408
rect 13841 17406 13863 17470
rect 13927 17406 13949 17470
rect 14013 17406 14035 17470
rect 14099 17406 14121 17470
rect 14185 17406 14207 17470
rect 14271 17406 14293 17470
rect 14357 17406 14379 17470
rect 14443 17406 14465 17470
rect 14529 17406 15000 17470
rect 1879 17402 15000 17406
rect 1160 17392 15000 17402
rect 1160 17386 2480 17392
rect 1160 17322 1287 17386
rect 1351 17322 1375 17386
rect 1439 17322 1463 17386
rect 1527 17322 1551 17386
rect 1615 17322 1639 17386
rect 1703 17322 1727 17386
rect 1791 17322 1815 17386
rect 1879 17328 2480 17386
rect 2544 17328 2608 17392
rect 2672 17328 3472 17392
rect 3536 17328 3600 17392
rect 3664 17328 4464 17392
rect 4528 17328 4592 17392
rect 4656 17328 5456 17392
rect 5520 17328 5584 17392
rect 5648 17328 6448 17392
rect 6512 17328 6576 17392
rect 6640 17328 7440 17392
rect 7504 17328 7568 17392
rect 7632 17328 8432 17392
rect 8496 17328 8560 17392
rect 8624 17328 9424 17392
rect 9488 17328 9552 17392
rect 9616 17328 10416 17392
rect 10480 17328 10544 17392
rect 10608 17328 11408 17392
rect 11472 17328 11536 17392
rect 11600 17328 12400 17392
rect 12464 17328 12528 17392
rect 12592 17328 13392 17392
rect 13456 17328 13520 17392
rect 13584 17390 15000 17392
rect 13584 17328 13777 17390
rect 1879 17326 13777 17328
rect 13841 17326 13863 17390
rect 13927 17326 13949 17390
rect 14013 17326 14035 17390
rect 14099 17326 14121 17390
rect 14185 17326 14207 17390
rect 14271 17326 14293 17390
rect 14357 17326 14379 17390
rect 14443 17326 14465 17390
rect 14529 17326 15000 17390
rect 1879 17322 15000 17326
rect 1160 17312 15000 17322
rect 1160 17306 2480 17312
rect 1160 17242 1287 17306
rect 1351 17242 1375 17306
rect 1439 17242 1463 17306
rect 1527 17242 1551 17306
rect 1615 17242 1639 17306
rect 1703 17242 1727 17306
rect 1791 17242 1815 17306
rect 1879 17248 2480 17306
rect 2544 17248 2608 17312
rect 2672 17248 3472 17312
rect 3536 17248 3600 17312
rect 3664 17248 4464 17312
rect 4528 17248 4592 17312
rect 4656 17248 5456 17312
rect 5520 17248 5584 17312
rect 5648 17248 6448 17312
rect 6512 17248 6576 17312
rect 6640 17248 7440 17312
rect 7504 17248 7568 17312
rect 7632 17248 8432 17312
rect 8496 17248 8560 17312
rect 8624 17248 9424 17312
rect 9488 17248 9552 17312
rect 9616 17248 10416 17312
rect 10480 17248 10544 17312
rect 10608 17248 11408 17312
rect 11472 17248 11536 17312
rect 11600 17248 12400 17312
rect 12464 17248 12528 17312
rect 12592 17248 13392 17312
rect 13456 17248 13520 17312
rect 13584 17310 15000 17312
rect 13584 17248 13777 17310
rect 1879 17246 13777 17248
rect 13841 17246 13863 17310
rect 13927 17246 13949 17310
rect 14013 17246 14035 17310
rect 14099 17246 14121 17310
rect 14185 17246 14207 17310
rect 14271 17246 14293 17310
rect 14357 17246 14379 17310
rect 14443 17246 14465 17310
rect 14529 17246 15000 17310
rect 1879 17242 15000 17246
rect 1160 17232 15000 17242
rect 1160 17226 2480 17232
rect 1160 17162 1287 17226
rect 1351 17162 1375 17226
rect 1439 17162 1463 17226
rect 1527 17162 1551 17226
rect 1615 17162 1639 17226
rect 1703 17162 1727 17226
rect 1791 17162 1815 17226
rect 1879 17168 2480 17226
rect 2544 17168 2608 17232
rect 2672 17168 3472 17232
rect 3536 17168 3600 17232
rect 3664 17168 4464 17232
rect 4528 17168 4592 17232
rect 4656 17168 5456 17232
rect 5520 17168 5584 17232
rect 5648 17168 6448 17232
rect 6512 17168 6576 17232
rect 6640 17168 7440 17232
rect 7504 17168 7568 17232
rect 7632 17168 8432 17232
rect 8496 17168 8560 17232
rect 8624 17168 9424 17232
rect 9488 17168 9552 17232
rect 9616 17168 10416 17232
rect 10480 17168 10544 17232
rect 10608 17168 11408 17232
rect 11472 17168 11536 17232
rect 11600 17168 12400 17232
rect 12464 17168 12528 17232
rect 12592 17168 13392 17232
rect 13456 17168 13520 17232
rect 13584 17230 15000 17232
rect 13584 17168 13777 17230
rect 1879 17166 13777 17168
rect 13841 17166 13863 17230
rect 13927 17166 13949 17230
rect 14013 17166 14035 17230
rect 14099 17166 14121 17230
rect 14185 17166 14207 17230
rect 14271 17166 14293 17230
rect 14357 17166 14379 17230
rect 14443 17166 14465 17230
rect 14529 17166 15000 17230
rect 1879 17162 15000 17166
rect 1160 17152 15000 17162
rect 1160 17146 2480 17152
rect 1160 17082 1287 17146
rect 1351 17082 1375 17146
rect 1439 17082 1463 17146
rect 1527 17082 1551 17146
rect 1615 17082 1639 17146
rect 1703 17082 1727 17146
rect 1791 17082 1815 17146
rect 1879 17088 2480 17146
rect 2544 17088 2608 17152
rect 2672 17088 3472 17152
rect 3536 17088 3600 17152
rect 3664 17088 4464 17152
rect 4528 17088 4592 17152
rect 4656 17088 5456 17152
rect 5520 17088 5584 17152
rect 5648 17088 6448 17152
rect 6512 17088 6576 17152
rect 6640 17088 7440 17152
rect 7504 17088 7568 17152
rect 7632 17088 8432 17152
rect 8496 17088 8560 17152
rect 8624 17088 9424 17152
rect 9488 17088 9552 17152
rect 9616 17088 10416 17152
rect 10480 17088 10544 17152
rect 10608 17088 11408 17152
rect 11472 17088 11536 17152
rect 11600 17088 12400 17152
rect 12464 17088 12528 17152
rect 12592 17088 13392 17152
rect 13456 17088 13520 17152
rect 13584 17150 15000 17152
rect 13584 17088 13777 17150
rect 1879 17086 13777 17088
rect 13841 17086 13863 17150
rect 13927 17086 13949 17150
rect 14013 17086 14035 17150
rect 14099 17086 14121 17150
rect 14185 17086 14207 17150
rect 14271 17086 14293 17150
rect 14357 17086 14379 17150
rect 14443 17086 14465 17150
rect 14529 17086 15000 17150
rect 1879 17082 15000 17086
rect 1160 17072 15000 17082
rect 1160 17066 2480 17072
rect 1160 17002 1287 17066
rect 1351 17002 1375 17066
rect 1439 17002 1463 17066
rect 1527 17002 1551 17066
rect 1615 17002 1639 17066
rect 1703 17002 1727 17066
rect 1791 17002 1815 17066
rect 1879 17008 2480 17066
rect 2544 17008 2608 17072
rect 2672 17008 3472 17072
rect 3536 17008 3600 17072
rect 3664 17008 4464 17072
rect 4528 17008 4592 17072
rect 4656 17008 5456 17072
rect 5520 17008 5584 17072
rect 5648 17008 6448 17072
rect 6512 17008 6576 17072
rect 6640 17008 7440 17072
rect 7504 17008 7568 17072
rect 7632 17008 8432 17072
rect 8496 17008 8560 17072
rect 8624 17008 9424 17072
rect 9488 17008 9552 17072
rect 9616 17008 10416 17072
rect 10480 17008 10544 17072
rect 10608 17008 11408 17072
rect 11472 17008 11536 17072
rect 11600 17008 12400 17072
rect 12464 17008 12528 17072
rect 12592 17008 13392 17072
rect 13456 17008 13520 17072
rect 13584 17070 15000 17072
rect 13584 17008 13777 17070
rect 1879 17006 13777 17008
rect 13841 17006 13863 17070
rect 13927 17006 13949 17070
rect 14013 17006 14035 17070
rect 14099 17006 14121 17070
rect 14185 17006 14207 17070
rect 14271 17006 14293 17070
rect 14357 17006 14379 17070
rect 14443 17006 14465 17070
rect 14529 17006 15000 17070
rect 1879 17002 15000 17006
rect 1160 16992 15000 17002
rect 1160 16986 2480 16992
rect 1160 16922 1287 16986
rect 1351 16922 1375 16986
rect 1439 16922 1463 16986
rect 1527 16922 1551 16986
rect 1615 16922 1639 16986
rect 1703 16922 1727 16986
rect 1791 16922 1815 16986
rect 1879 16928 2480 16986
rect 2544 16928 2608 16992
rect 2672 16928 3472 16992
rect 3536 16928 3600 16992
rect 3664 16928 4464 16992
rect 4528 16928 4592 16992
rect 4656 16928 5456 16992
rect 5520 16928 5584 16992
rect 5648 16928 6448 16992
rect 6512 16928 6576 16992
rect 6640 16928 7440 16992
rect 7504 16928 7568 16992
rect 7632 16928 8432 16992
rect 8496 16928 8560 16992
rect 8624 16928 9424 16992
rect 9488 16928 9552 16992
rect 9616 16928 10416 16992
rect 10480 16928 10544 16992
rect 10608 16928 11408 16992
rect 11472 16928 11536 16992
rect 11600 16928 12400 16992
rect 12464 16928 12528 16992
rect 12592 16928 13392 16992
rect 13456 16928 13520 16992
rect 13584 16990 15000 16992
rect 13584 16928 13777 16990
rect 1879 16926 13777 16928
rect 13841 16926 13863 16990
rect 13927 16926 13949 16990
rect 14013 16926 14035 16990
rect 14099 16926 14121 16990
rect 14185 16926 14207 16990
rect 14271 16926 14293 16990
rect 14357 16926 14379 16990
rect 14443 16926 14465 16990
rect 14529 16926 15000 16990
rect 1879 16922 15000 16926
rect 1160 16912 15000 16922
rect 1160 16906 2480 16912
rect 1160 16842 1287 16906
rect 1351 16842 1375 16906
rect 1439 16842 1463 16906
rect 1527 16842 1551 16906
rect 1615 16842 1639 16906
rect 1703 16842 1727 16906
rect 1791 16842 1815 16906
rect 1879 16848 2480 16906
rect 2544 16848 2608 16912
rect 2672 16848 3472 16912
rect 3536 16848 3600 16912
rect 3664 16848 4464 16912
rect 4528 16848 4592 16912
rect 4656 16848 5456 16912
rect 5520 16848 5584 16912
rect 5648 16848 6448 16912
rect 6512 16848 6576 16912
rect 6640 16848 7440 16912
rect 7504 16848 7568 16912
rect 7632 16848 8432 16912
rect 8496 16848 8560 16912
rect 8624 16848 9424 16912
rect 9488 16848 9552 16912
rect 9616 16848 10416 16912
rect 10480 16848 10544 16912
rect 10608 16848 11408 16912
rect 11472 16848 11536 16912
rect 11600 16848 12400 16912
rect 12464 16848 12528 16912
rect 12592 16848 13392 16912
rect 13456 16848 13520 16912
rect 13584 16910 15000 16912
rect 13584 16848 13777 16910
rect 1879 16846 13777 16848
rect 13841 16846 13863 16910
rect 13927 16846 13949 16910
rect 14013 16846 14035 16910
rect 14099 16846 14121 16910
rect 14185 16846 14207 16910
rect 14271 16846 14293 16910
rect 14357 16846 14379 16910
rect 14443 16846 14465 16910
rect 14529 16846 15000 16910
rect 1879 16842 15000 16846
rect 1160 16832 15000 16842
rect 1160 16826 2480 16832
rect 1160 16762 1287 16826
rect 1351 16762 1375 16826
rect 1439 16762 1463 16826
rect 1527 16762 1551 16826
rect 1615 16762 1639 16826
rect 1703 16762 1727 16826
rect 1791 16762 1815 16826
rect 1879 16768 2480 16826
rect 2544 16768 2608 16832
rect 2672 16768 3472 16832
rect 3536 16768 3600 16832
rect 3664 16768 4464 16832
rect 4528 16768 4592 16832
rect 4656 16768 5456 16832
rect 5520 16768 5584 16832
rect 5648 16768 6448 16832
rect 6512 16768 6576 16832
rect 6640 16768 7440 16832
rect 7504 16768 7568 16832
rect 7632 16768 8432 16832
rect 8496 16768 8560 16832
rect 8624 16768 9424 16832
rect 9488 16768 9552 16832
rect 9616 16768 10416 16832
rect 10480 16768 10544 16832
rect 10608 16768 11408 16832
rect 11472 16768 11536 16832
rect 11600 16768 12400 16832
rect 12464 16768 12528 16832
rect 12592 16768 13392 16832
rect 13456 16768 13520 16832
rect 13584 16830 15000 16832
rect 13584 16768 13777 16830
rect 1879 16766 13777 16768
rect 13841 16766 13863 16830
rect 13927 16766 13949 16830
rect 14013 16766 14035 16830
rect 14099 16766 14121 16830
rect 14185 16766 14207 16830
rect 14271 16766 14293 16830
rect 14357 16766 14379 16830
rect 14443 16766 14465 16830
rect 14529 16766 15000 16830
rect 1879 16762 15000 16766
rect 1160 16752 15000 16762
rect 1160 16746 2480 16752
rect 1160 16682 1287 16746
rect 1351 16682 1375 16746
rect 1439 16682 1463 16746
rect 1527 16682 1551 16746
rect 1615 16682 1639 16746
rect 1703 16682 1727 16746
rect 1791 16682 1815 16746
rect 1879 16688 2480 16746
rect 2544 16688 2608 16752
rect 2672 16688 3472 16752
rect 3536 16688 3600 16752
rect 3664 16688 4464 16752
rect 4528 16688 4592 16752
rect 4656 16688 5456 16752
rect 5520 16688 5584 16752
rect 5648 16688 6448 16752
rect 6512 16688 6576 16752
rect 6640 16688 7440 16752
rect 7504 16688 7568 16752
rect 7632 16688 8432 16752
rect 8496 16688 8560 16752
rect 8624 16688 9424 16752
rect 9488 16688 9552 16752
rect 9616 16688 10416 16752
rect 10480 16688 10544 16752
rect 10608 16688 11408 16752
rect 11472 16688 11536 16752
rect 11600 16688 12400 16752
rect 12464 16688 12528 16752
rect 12592 16688 13392 16752
rect 13456 16688 13520 16752
rect 13584 16750 15000 16752
rect 13584 16688 13777 16750
rect 1879 16686 13777 16688
rect 13841 16686 13863 16750
rect 13927 16686 13949 16750
rect 14013 16686 14035 16750
rect 14099 16686 14121 16750
rect 14185 16686 14207 16750
rect 14271 16686 14293 16750
rect 14357 16686 14379 16750
rect 14443 16686 14465 16750
rect 14529 16686 15000 16750
rect 1879 16682 15000 16686
rect 1160 16672 15000 16682
rect 1160 16666 2480 16672
rect 1160 16602 1287 16666
rect 1351 16602 1375 16666
rect 1439 16602 1463 16666
rect 1527 16602 1551 16666
rect 1615 16602 1639 16666
rect 1703 16602 1727 16666
rect 1791 16602 1815 16666
rect 1879 16608 2480 16666
rect 2544 16608 2608 16672
rect 2672 16608 3472 16672
rect 3536 16608 3600 16672
rect 3664 16608 4464 16672
rect 4528 16608 4592 16672
rect 4656 16608 5456 16672
rect 5520 16608 5584 16672
rect 5648 16608 6448 16672
rect 6512 16608 6576 16672
rect 6640 16608 7440 16672
rect 7504 16608 7568 16672
rect 7632 16608 8432 16672
rect 8496 16608 8560 16672
rect 8624 16608 9424 16672
rect 9488 16608 9552 16672
rect 9616 16608 10416 16672
rect 10480 16608 10544 16672
rect 10608 16608 11408 16672
rect 11472 16608 11536 16672
rect 11600 16608 12400 16672
rect 12464 16608 12528 16672
rect 12592 16608 13392 16672
rect 13456 16608 13520 16672
rect 13584 16670 15000 16672
rect 13584 16608 13777 16670
rect 1879 16606 13777 16608
rect 13841 16606 13863 16670
rect 13927 16606 13949 16670
rect 14013 16606 14035 16670
rect 14099 16606 14121 16670
rect 14185 16606 14207 16670
rect 14271 16606 14293 16670
rect 14357 16606 14379 16670
rect 14443 16606 14465 16670
rect 14529 16606 15000 16670
rect 1879 16602 15000 16606
rect 1160 16592 15000 16602
rect 1160 16586 2480 16592
rect 1160 16522 1287 16586
rect 1351 16522 1375 16586
rect 1439 16522 1463 16586
rect 1527 16522 1551 16586
rect 1615 16522 1639 16586
rect 1703 16522 1727 16586
rect 1791 16522 1815 16586
rect 1879 16528 2480 16586
rect 2544 16528 2608 16592
rect 2672 16528 3472 16592
rect 3536 16528 3600 16592
rect 3664 16528 4464 16592
rect 4528 16528 4592 16592
rect 4656 16528 5456 16592
rect 5520 16528 5584 16592
rect 5648 16528 6448 16592
rect 6512 16528 6576 16592
rect 6640 16528 7440 16592
rect 7504 16528 7568 16592
rect 7632 16528 8432 16592
rect 8496 16528 8560 16592
rect 8624 16528 9424 16592
rect 9488 16528 9552 16592
rect 9616 16528 10416 16592
rect 10480 16528 10544 16592
rect 10608 16528 11408 16592
rect 11472 16528 11536 16592
rect 11600 16528 12400 16592
rect 12464 16528 12528 16592
rect 12592 16528 13392 16592
rect 13456 16528 13520 16592
rect 13584 16590 15000 16592
rect 13584 16528 13777 16590
rect 1879 16526 13777 16528
rect 13841 16526 13863 16590
rect 13927 16526 13949 16590
rect 14013 16526 14035 16590
rect 14099 16526 14121 16590
rect 14185 16526 14207 16590
rect 14271 16526 14293 16590
rect 14357 16526 14379 16590
rect 14443 16526 14465 16590
rect 14529 16526 15000 16590
rect 1879 16522 15000 16526
rect 1160 16512 15000 16522
rect 1160 16506 2480 16512
rect 1160 16442 1287 16506
rect 1351 16442 1375 16506
rect 1439 16442 1463 16506
rect 1527 16442 1551 16506
rect 1615 16442 1639 16506
rect 1703 16442 1727 16506
rect 1791 16442 1815 16506
rect 1879 16448 2480 16506
rect 2544 16448 2608 16512
rect 2672 16448 3472 16512
rect 3536 16448 3600 16512
rect 3664 16448 4464 16512
rect 4528 16448 4592 16512
rect 4656 16448 5456 16512
rect 5520 16448 5584 16512
rect 5648 16448 6448 16512
rect 6512 16448 6576 16512
rect 6640 16448 7440 16512
rect 7504 16448 7568 16512
rect 7632 16448 8432 16512
rect 8496 16448 8560 16512
rect 8624 16448 9424 16512
rect 9488 16448 9552 16512
rect 9616 16448 10416 16512
rect 10480 16448 10544 16512
rect 10608 16448 11408 16512
rect 11472 16448 11536 16512
rect 11600 16448 12400 16512
rect 12464 16448 12528 16512
rect 12592 16448 13392 16512
rect 13456 16448 13520 16512
rect 13584 16510 15000 16512
rect 13584 16448 13777 16510
rect 1879 16446 13777 16448
rect 13841 16446 13863 16510
rect 13927 16446 13949 16510
rect 14013 16446 14035 16510
rect 14099 16446 14121 16510
rect 14185 16446 14207 16510
rect 14271 16446 14293 16510
rect 14357 16446 14379 16510
rect 14443 16446 14465 16510
rect 14529 16446 15000 16510
rect 1879 16442 15000 16446
rect 1160 16432 15000 16442
rect 1160 16426 2480 16432
rect 1160 16362 1287 16426
rect 1351 16362 1375 16426
rect 1439 16362 1463 16426
rect 1527 16362 1551 16426
rect 1615 16362 1639 16426
rect 1703 16362 1727 16426
rect 1791 16362 1815 16426
rect 1879 16368 2480 16426
rect 2544 16368 2608 16432
rect 2672 16368 3472 16432
rect 3536 16368 3600 16432
rect 3664 16368 4464 16432
rect 4528 16368 4592 16432
rect 4656 16431 6448 16432
rect 4656 16368 5456 16431
rect 1879 16367 5456 16368
rect 5520 16367 5584 16431
rect 5648 16368 6448 16431
rect 6512 16368 6576 16432
rect 6640 16368 7440 16432
rect 7504 16368 7568 16432
rect 7632 16368 8432 16432
rect 8496 16368 8560 16432
rect 8624 16368 9424 16432
rect 9488 16368 9552 16432
rect 9616 16368 10416 16432
rect 10480 16368 10544 16432
rect 10608 16368 11408 16432
rect 11472 16368 11536 16432
rect 11600 16368 12400 16432
rect 12464 16368 12528 16432
rect 12592 16368 13392 16432
rect 13456 16368 13520 16432
rect 13584 16430 15000 16432
rect 13584 16368 13777 16430
rect 5648 16367 13777 16368
rect 1879 16366 13777 16367
rect 13841 16366 13863 16430
rect 13927 16366 13949 16430
rect 14013 16366 14035 16430
rect 14099 16366 14121 16430
rect 14185 16366 14207 16430
rect 14271 16366 14293 16430
rect 14357 16366 14379 16430
rect 14443 16366 14465 16430
rect 14529 16366 15000 16430
rect 1879 16362 15000 16366
rect 1160 16351 15000 16362
rect 1160 16346 2480 16351
rect 1160 16282 1287 16346
rect 1351 16282 1375 16346
rect 1439 16282 1463 16346
rect 1527 16282 1551 16346
rect 1615 16282 1639 16346
rect 1703 16282 1727 16346
rect 1791 16282 1815 16346
rect 1879 16287 2480 16346
rect 2544 16287 2608 16351
rect 2672 16287 3472 16351
rect 3536 16287 3600 16351
rect 3664 16287 4464 16351
rect 4528 16287 4592 16351
rect 4656 16350 6448 16351
rect 4656 16287 5456 16350
rect 1879 16286 5456 16287
rect 5520 16286 5584 16350
rect 5648 16287 6448 16350
rect 6512 16287 6576 16351
rect 6640 16287 7440 16351
rect 7504 16287 7568 16351
rect 7632 16287 8432 16351
rect 8496 16287 8560 16351
rect 8624 16287 9424 16351
rect 9488 16287 9552 16351
rect 9616 16287 10416 16351
rect 10480 16287 10544 16351
rect 10608 16287 11408 16351
rect 11472 16287 11536 16351
rect 11600 16287 12400 16351
rect 12464 16287 12528 16351
rect 12592 16287 13392 16351
rect 13456 16287 13520 16351
rect 13584 16350 15000 16351
rect 13584 16287 13777 16350
rect 5648 16286 13777 16287
rect 13841 16286 13863 16350
rect 13927 16286 13949 16350
rect 14013 16286 14035 16350
rect 14099 16286 14121 16350
rect 14185 16286 14207 16350
rect 14271 16286 14293 16350
rect 14357 16286 14379 16350
rect 14443 16286 14465 16350
rect 14529 16286 15000 16350
rect 1879 16282 15000 16286
rect 1160 16270 15000 16282
rect 1160 16266 2480 16270
rect 1160 16202 1287 16266
rect 1351 16202 1375 16266
rect 1439 16202 1463 16266
rect 1527 16202 1551 16266
rect 1615 16202 1639 16266
rect 1703 16202 1727 16266
rect 1791 16202 1815 16266
rect 1879 16206 2480 16266
rect 2544 16206 2608 16270
rect 2672 16206 3472 16270
rect 3536 16206 3600 16270
rect 3664 16206 4464 16270
rect 4528 16206 4592 16270
rect 4656 16269 6448 16270
rect 4656 16206 5456 16269
rect 1879 16205 5456 16206
rect 5520 16205 5584 16269
rect 5648 16206 6448 16269
rect 6512 16206 6576 16270
rect 6640 16206 7440 16270
rect 7504 16206 7568 16270
rect 7632 16206 8432 16270
rect 8496 16206 8560 16270
rect 8624 16206 9424 16270
rect 9488 16206 9552 16270
rect 9616 16206 10416 16270
rect 10480 16206 10544 16270
rect 10608 16206 11408 16270
rect 11472 16206 11536 16270
rect 11600 16206 12400 16270
rect 12464 16206 12528 16270
rect 12592 16206 13392 16270
rect 13456 16206 13520 16270
rect 13584 16206 13777 16270
rect 13841 16206 13863 16270
rect 13927 16206 13949 16270
rect 14013 16206 14035 16270
rect 14099 16206 14121 16270
rect 14185 16206 14207 16270
rect 14271 16206 14293 16270
rect 14357 16206 14379 16270
rect 14443 16206 14465 16270
rect 14529 16206 15000 16270
rect 5648 16205 15000 16206
rect 1879 16202 15000 16205
rect 1160 16190 15000 16202
rect 1160 16189 13777 16190
rect 1160 16186 2480 16189
rect 1160 16122 1287 16186
rect 1351 16122 1375 16186
rect 1439 16122 1463 16186
rect 1527 16122 1551 16186
rect 1615 16122 1639 16186
rect 1703 16122 1727 16186
rect 1791 16122 1815 16186
rect 1879 16125 2480 16186
rect 2544 16125 2608 16189
rect 2672 16125 3472 16189
rect 3536 16125 3600 16189
rect 3664 16125 4464 16189
rect 4528 16125 4592 16189
rect 4656 16188 6448 16189
rect 4656 16125 5456 16188
rect 1879 16124 5456 16125
rect 5520 16124 5584 16188
rect 5648 16125 6448 16188
rect 6512 16125 6576 16189
rect 6640 16125 7440 16189
rect 7504 16125 7568 16189
rect 7632 16125 8432 16189
rect 8496 16125 8560 16189
rect 8624 16125 9424 16189
rect 9488 16125 9552 16189
rect 9616 16125 10416 16189
rect 10480 16125 10544 16189
rect 10608 16125 11408 16189
rect 11472 16125 11536 16189
rect 11600 16125 12400 16189
rect 12464 16125 12528 16189
rect 12592 16125 13392 16189
rect 13456 16125 13520 16189
rect 13584 16126 13777 16189
rect 13841 16126 13863 16190
rect 13927 16126 13949 16190
rect 14013 16126 14035 16190
rect 14099 16126 14121 16190
rect 14185 16126 14207 16190
rect 14271 16126 14293 16190
rect 14357 16126 14379 16190
rect 14443 16126 14465 16190
rect 14529 16126 15000 16190
rect 13584 16125 15000 16126
rect 5648 16124 15000 16125
rect 1879 16122 15000 16124
rect 1160 16110 15000 16122
rect 1160 16108 13777 16110
rect 1160 16106 2480 16108
rect 1160 16042 1287 16106
rect 1351 16042 1375 16106
rect 1439 16042 1463 16106
rect 1527 16042 1551 16106
rect 1615 16042 1639 16106
rect 1703 16042 1727 16106
rect 1791 16042 1815 16106
rect 1879 16044 2480 16106
rect 2544 16044 2608 16108
rect 2672 16044 3472 16108
rect 3536 16044 3600 16108
rect 3664 16044 4464 16108
rect 4528 16044 4592 16108
rect 4656 16107 6448 16108
rect 4656 16044 5456 16107
rect 1879 16043 5456 16044
rect 5520 16043 5584 16107
rect 5648 16044 6448 16107
rect 6512 16044 6576 16108
rect 6640 16044 7440 16108
rect 7504 16044 7568 16108
rect 7632 16044 8432 16108
rect 8496 16044 8560 16108
rect 8624 16044 9424 16108
rect 9488 16044 9552 16108
rect 9616 16044 10416 16108
rect 10480 16044 10544 16108
rect 10608 16044 11408 16108
rect 11472 16044 11536 16108
rect 11600 16044 12400 16108
rect 12464 16044 12528 16108
rect 12592 16044 13392 16108
rect 13456 16044 13520 16108
rect 13584 16046 13777 16108
rect 13841 16046 13863 16110
rect 13927 16046 13949 16110
rect 14013 16046 14035 16110
rect 14099 16046 14121 16110
rect 14185 16046 14207 16110
rect 14271 16046 14293 16110
rect 14357 16046 14379 16110
rect 14443 16046 14465 16110
rect 14529 16046 15000 16110
rect 13584 16044 15000 16046
rect 5648 16043 15000 16044
rect 1879 16042 15000 16043
rect 1160 16030 15000 16042
rect 1160 16027 13777 16030
rect 1160 16026 2480 16027
rect 1160 15962 1287 16026
rect 1351 15962 1375 16026
rect 1439 15962 1463 16026
rect 1527 15962 1551 16026
rect 1615 15962 1639 16026
rect 1703 15962 1727 16026
rect 1791 15962 1815 16026
rect 1879 15963 2480 16026
rect 2544 15963 2608 16027
rect 2672 15963 3472 16027
rect 3536 15963 3600 16027
rect 3664 15963 4464 16027
rect 4528 15963 4592 16027
rect 4656 16026 6448 16027
rect 4656 15963 5456 16026
rect 1879 15962 5456 15963
rect 5520 15962 5584 16026
rect 5648 15963 6448 16026
rect 6512 15963 6576 16027
rect 6640 15963 7440 16027
rect 7504 15963 7568 16027
rect 7632 15963 8432 16027
rect 8496 15963 8560 16027
rect 8624 15963 9424 16027
rect 9488 15963 9552 16027
rect 9616 15963 10416 16027
rect 10480 15963 10544 16027
rect 10608 15963 11408 16027
rect 11472 15963 11536 16027
rect 11600 15963 12400 16027
rect 12464 15963 12528 16027
rect 12592 15963 13392 16027
rect 13456 15963 13520 16027
rect 13584 15966 13777 16027
rect 13841 15966 13863 16030
rect 13927 15966 13949 16030
rect 14013 15966 14035 16030
rect 14099 15966 14121 16030
rect 14185 15966 14207 16030
rect 14271 15966 14293 16030
rect 14357 15966 14379 16030
rect 14443 15966 14465 16030
rect 14529 15966 15000 16030
rect 13584 15963 15000 15966
rect 5648 15962 15000 15963
rect 1160 15950 15000 15962
rect 1160 15946 13777 15950
rect 1160 15882 1287 15946
rect 1351 15882 1375 15946
rect 1439 15882 1463 15946
rect 1527 15882 1551 15946
rect 1615 15882 1639 15946
rect 1703 15882 1727 15946
rect 1791 15882 1815 15946
rect 1879 15882 2480 15946
rect 2544 15882 2608 15946
rect 2672 15882 3472 15946
rect 3536 15882 3600 15946
rect 3664 15882 4464 15946
rect 4528 15882 4592 15946
rect 4656 15945 6448 15946
rect 4656 15882 5456 15945
rect 1160 15881 5456 15882
rect 5520 15881 5584 15945
rect 5648 15882 6448 15945
rect 6512 15882 6576 15946
rect 6640 15882 7440 15946
rect 7504 15882 7568 15946
rect 7632 15882 8432 15946
rect 8496 15882 8560 15946
rect 8624 15882 9424 15946
rect 9488 15882 9552 15946
rect 9616 15882 10416 15946
rect 10480 15882 10544 15946
rect 10608 15882 11408 15946
rect 11472 15882 11536 15946
rect 11600 15882 12400 15946
rect 12464 15882 12528 15946
rect 12592 15882 13392 15946
rect 13456 15882 13520 15946
rect 13584 15886 13777 15946
rect 13841 15886 13863 15950
rect 13927 15886 13949 15950
rect 14013 15886 14035 15950
rect 14099 15886 14121 15950
rect 14185 15886 14207 15950
rect 14271 15886 14293 15950
rect 14357 15886 14379 15950
rect 14443 15886 14465 15950
rect 14529 15886 15000 15950
rect 13584 15882 15000 15886
rect 5648 15881 15000 15882
rect 1160 15870 15000 15881
rect 1160 15866 13777 15870
rect 1160 15802 1287 15866
rect 1351 15802 1375 15866
rect 1439 15802 1463 15866
rect 1527 15802 1551 15866
rect 1615 15802 1639 15866
rect 1703 15802 1727 15866
rect 1791 15802 1815 15866
rect 1879 15865 13777 15866
rect 1879 15802 2480 15865
rect 1160 15801 2480 15802
rect 2544 15801 2608 15865
rect 2672 15801 3472 15865
rect 3536 15801 3600 15865
rect 3664 15801 4464 15865
rect 4528 15801 4592 15865
rect 4656 15864 6448 15865
rect 4656 15801 5456 15864
rect 1160 15800 5456 15801
rect 5520 15800 5584 15864
rect 5648 15801 6448 15864
rect 6512 15801 6576 15865
rect 6640 15801 7440 15865
rect 7504 15801 7568 15865
rect 7632 15801 8432 15865
rect 8496 15801 8560 15865
rect 8624 15801 9424 15865
rect 9488 15801 9552 15865
rect 9616 15801 10416 15865
rect 10480 15801 10544 15865
rect 10608 15801 11408 15865
rect 11472 15801 11536 15865
rect 11600 15801 12400 15865
rect 12464 15801 12528 15865
rect 12592 15801 13392 15865
rect 13456 15801 13520 15865
rect 13584 15806 13777 15865
rect 13841 15806 13863 15870
rect 13927 15806 13949 15870
rect 14013 15806 14035 15870
rect 14099 15806 14121 15870
rect 14185 15806 14207 15870
rect 14271 15806 14293 15870
rect 14357 15806 14379 15870
rect 14443 15806 14465 15870
rect 14529 15806 15000 15870
rect 13584 15801 15000 15806
rect 5648 15800 15000 15801
rect 1160 15790 15000 15800
rect 1160 15786 13777 15790
rect 1160 15722 1287 15786
rect 1351 15722 1375 15786
rect 1439 15722 1463 15786
rect 1527 15722 1551 15786
rect 1615 15722 1639 15786
rect 1703 15722 1727 15786
rect 1791 15722 1815 15786
rect 1879 15784 13777 15786
rect 1879 15722 2480 15784
rect 1160 15720 2480 15722
rect 2544 15720 2608 15784
rect 2672 15720 3472 15784
rect 3536 15720 3600 15784
rect 3664 15720 4464 15784
rect 4528 15720 4592 15784
rect 4656 15783 6448 15784
rect 4656 15720 5456 15783
rect 1160 15719 5456 15720
rect 5520 15719 5584 15783
rect 5648 15720 6448 15783
rect 6512 15720 6576 15784
rect 6640 15720 7440 15784
rect 7504 15720 7568 15784
rect 7632 15720 8432 15784
rect 8496 15720 8560 15784
rect 8624 15720 9424 15784
rect 9488 15720 9552 15784
rect 9616 15720 10416 15784
rect 10480 15720 10544 15784
rect 10608 15720 11408 15784
rect 11472 15720 11536 15784
rect 11600 15720 12400 15784
rect 12464 15720 12528 15784
rect 12592 15720 13392 15784
rect 13456 15720 13520 15784
rect 13584 15726 13777 15784
rect 13841 15726 13863 15790
rect 13927 15726 13949 15790
rect 14013 15726 14035 15790
rect 14099 15726 14121 15790
rect 14185 15726 14207 15790
rect 14271 15726 14293 15790
rect 14357 15726 14379 15790
rect 14443 15726 14465 15790
rect 14529 15726 15000 15790
rect 13584 15720 15000 15726
rect 5648 15719 15000 15720
rect 1160 15710 15000 15719
rect 1160 15706 13777 15710
rect 1160 15642 1287 15706
rect 1351 15642 1375 15706
rect 1439 15642 1463 15706
rect 1527 15642 1551 15706
rect 1615 15642 1639 15706
rect 1703 15642 1727 15706
rect 1791 15642 1815 15706
rect 1879 15703 13777 15706
rect 1879 15642 2480 15703
rect 1160 15639 2480 15642
rect 2544 15639 2608 15703
rect 2672 15639 3472 15703
rect 3536 15639 3600 15703
rect 3664 15639 4464 15703
rect 4528 15639 4592 15703
rect 4656 15702 6448 15703
rect 4656 15639 5456 15702
rect 1160 15638 5456 15639
rect 5520 15638 5584 15702
rect 5648 15639 6448 15702
rect 6512 15639 6576 15703
rect 6640 15639 7440 15703
rect 7504 15639 7568 15703
rect 7632 15639 8432 15703
rect 8496 15639 8560 15703
rect 8624 15639 9424 15703
rect 9488 15639 9552 15703
rect 9616 15639 10416 15703
rect 10480 15639 10544 15703
rect 10608 15639 11408 15703
rect 11472 15639 11536 15703
rect 11600 15639 12400 15703
rect 12464 15639 12528 15703
rect 12592 15639 13392 15703
rect 13456 15639 13520 15703
rect 13584 15646 13777 15703
rect 13841 15646 13863 15710
rect 13927 15646 13949 15710
rect 14013 15646 14035 15710
rect 14099 15646 14121 15710
rect 14185 15646 14207 15710
rect 14271 15646 14293 15710
rect 14357 15646 14379 15710
rect 14443 15646 14465 15710
rect 14529 15646 15000 15710
rect 13584 15639 15000 15646
rect 5648 15638 15000 15639
rect 1160 15630 15000 15638
rect 1160 15626 13777 15630
rect 1160 15562 1287 15626
rect 1351 15562 1375 15626
rect 1439 15562 1463 15626
rect 1527 15562 1551 15626
rect 1615 15562 1639 15626
rect 1703 15562 1727 15626
rect 1791 15562 1815 15626
rect 1879 15622 13777 15626
rect 1879 15562 2480 15622
rect 1160 15558 2480 15562
rect 2544 15558 2608 15622
rect 2672 15558 3472 15622
rect 3536 15558 3600 15622
rect 3664 15558 4464 15622
rect 4528 15558 4592 15622
rect 4656 15621 6448 15622
rect 4656 15558 5456 15621
rect 1160 15557 5456 15558
rect 5520 15557 5584 15621
rect 5648 15558 6448 15621
rect 6512 15558 6576 15622
rect 6640 15558 7440 15622
rect 7504 15558 7568 15622
rect 7632 15558 8432 15622
rect 8496 15558 8560 15622
rect 8624 15558 9424 15622
rect 9488 15558 9552 15622
rect 9616 15558 10416 15622
rect 10480 15558 10544 15622
rect 10608 15558 11408 15622
rect 11472 15558 11536 15622
rect 11600 15558 12400 15622
rect 12464 15558 12528 15622
rect 12592 15558 13392 15622
rect 13456 15558 13520 15622
rect 13584 15566 13777 15622
rect 13841 15566 13863 15630
rect 13927 15566 13949 15630
rect 14013 15566 14035 15630
rect 14099 15566 14121 15630
rect 14185 15566 14207 15630
rect 14271 15566 14293 15630
rect 14357 15566 14379 15630
rect 14443 15566 14465 15630
rect 14529 15566 15000 15630
rect 13584 15558 15000 15566
rect 5648 15557 15000 15558
rect 1160 15550 15000 15557
rect 1160 15546 13777 15550
rect 1160 15484 1287 15546
rect 0 15482 1287 15484
rect 1351 15482 1375 15546
rect 1439 15482 1463 15546
rect 1527 15482 1551 15546
rect 1615 15482 1639 15546
rect 1703 15482 1727 15546
rect 1791 15482 1815 15546
rect 1879 15541 13777 15546
rect 1879 15482 2480 15541
rect 0 15477 2480 15482
rect 2544 15477 2608 15541
rect 2672 15477 3472 15541
rect 3536 15477 3600 15541
rect 3664 15477 4464 15541
rect 4528 15477 4592 15541
rect 4656 15540 6448 15541
rect 4656 15477 5456 15540
rect 0 15476 5456 15477
rect 5520 15476 5584 15540
rect 5648 15477 6448 15540
rect 6512 15477 6576 15541
rect 6640 15477 7440 15541
rect 7504 15477 7568 15541
rect 7632 15477 8432 15541
rect 8496 15477 8560 15541
rect 8624 15477 9424 15541
rect 9488 15477 9552 15541
rect 9616 15477 10416 15541
rect 10480 15477 10544 15541
rect 10608 15477 11408 15541
rect 11472 15477 11536 15541
rect 11600 15477 12400 15541
rect 12464 15477 12528 15541
rect 12592 15477 13392 15541
rect 13456 15477 13520 15541
rect 13584 15486 13777 15541
rect 13841 15486 13863 15550
rect 13927 15486 13949 15550
rect 14013 15486 14035 15550
rect 14099 15486 14121 15550
rect 14185 15486 14207 15550
rect 14271 15486 14293 15550
rect 14357 15486 14379 15550
rect 14443 15486 14465 15550
rect 14529 15486 15000 15550
rect 13584 15477 15000 15486
rect 5648 15476 15000 15477
rect 0 15470 15000 15476
rect 0 15467 13777 15470
rect 0 15403 456 15467
rect 520 15403 536 15467
rect 600 15403 616 15467
rect 680 15403 696 15467
rect 760 15403 776 15467
rect 840 15403 856 15467
rect 920 15403 936 15467
rect 1000 15403 1016 15467
rect 1080 15403 1096 15467
rect 1160 15466 13777 15467
rect 1160 15403 1287 15466
rect 0 15402 1287 15403
rect 1351 15402 1375 15466
rect 1439 15402 1463 15466
rect 1527 15402 1551 15466
rect 1615 15402 1639 15466
rect 1703 15402 1727 15466
rect 1791 15402 1815 15466
rect 1879 15460 13777 15466
rect 1879 15402 2480 15460
rect 0 15396 2480 15402
rect 2544 15396 2608 15460
rect 2672 15396 3472 15460
rect 3536 15396 3600 15460
rect 3664 15396 4464 15460
rect 4528 15396 4592 15460
rect 4656 15459 6448 15460
rect 4656 15396 5456 15459
rect 0 15395 5456 15396
rect 5520 15395 5584 15459
rect 5648 15396 6448 15459
rect 6512 15396 6576 15460
rect 6640 15396 7440 15460
rect 7504 15396 7568 15460
rect 7632 15396 8432 15460
rect 8496 15396 8560 15460
rect 8624 15396 9424 15460
rect 9488 15396 9552 15460
rect 9616 15396 10416 15460
rect 10480 15396 10544 15460
rect 10608 15396 11408 15460
rect 11472 15396 11536 15460
rect 11600 15396 12400 15460
rect 12464 15396 12528 15460
rect 12592 15396 13392 15460
rect 13456 15396 13520 15460
rect 13584 15406 13777 15460
rect 13841 15406 13863 15470
rect 13927 15406 13949 15470
rect 14013 15406 14035 15470
rect 14099 15406 14121 15470
rect 14185 15406 14207 15470
rect 14271 15406 14293 15470
rect 14357 15406 14379 15470
rect 14443 15406 14465 15470
rect 14529 15406 15000 15470
rect 13584 15396 15000 15406
rect 5648 15395 15000 15396
rect 0 15390 15000 15395
rect 0 15386 13777 15390
rect 0 15322 456 15386
rect 520 15322 536 15386
rect 600 15322 616 15386
rect 680 15322 696 15386
rect 760 15322 776 15386
rect 840 15322 856 15386
rect 920 15322 936 15386
rect 1000 15322 1016 15386
rect 1080 15322 1096 15386
rect 1160 15322 1287 15386
rect 1351 15322 1375 15386
rect 1439 15322 1463 15386
rect 1527 15322 1551 15386
rect 1615 15322 1639 15386
rect 1703 15322 1727 15386
rect 1791 15322 1815 15386
rect 1879 15379 13777 15386
rect 1879 15322 2480 15379
rect 0 15315 2480 15322
rect 2544 15315 2608 15379
rect 2672 15315 3472 15379
rect 3536 15315 3600 15379
rect 3664 15315 4464 15379
rect 4528 15315 4592 15379
rect 4656 15378 6448 15379
rect 4656 15315 5456 15378
rect 0 15314 5456 15315
rect 5520 15314 5584 15378
rect 5648 15315 6448 15378
rect 6512 15315 6576 15379
rect 6640 15315 7440 15379
rect 7504 15315 7568 15379
rect 7632 15315 8432 15379
rect 8496 15315 8560 15379
rect 8624 15315 9424 15379
rect 9488 15315 9552 15379
rect 9616 15315 10416 15379
rect 10480 15315 10544 15379
rect 10608 15315 11408 15379
rect 11472 15315 11536 15379
rect 11600 15315 12400 15379
rect 12464 15315 12528 15379
rect 12592 15315 13392 15379
rect 13456 15315 13520 15379
rect 13584 15326 13777 15379
rect 13841 15326 13863 15390
rect 13927 15326 13949 15390
rect 14013 15326 14035 15390
rect 14099 15326 14121 15390
rect 14185 15326 14207 15390
rect 14271 15326 14293 15390
rect 14357 15326 14379 15390
rect 14443 15326 14465 15390
rect 14529 15326 15000 15390
rect 13584 15315 15000 15326
rect 5648 15314 15000 15315
rect 0 15310 15000 15314
rect 0 15306 13777 15310
rect 0 15305 1287 15306
rect 0 15241 456 15305
rect 520 15241 536 15305
rect 600 15241 616 15305
rect 680 15241 696 15305
rect 760 15241 776 15305
rect 840 15241 856 15305
rect 920 15241 936 15305
rect 1000 15241 1016 15305
rect 1080 15241 1096 15305
rect 1160 15242 1287 15305
rect 1351 15242 1375 15306
rect 1439 15242 1463 15306
rect 1527 15242 1551 15306
rect 1615 15242 1639 15306
rect 1703 15242 1727 15306
rect 1791 15242 1815 15306
rect 1879 15298 13777 15306
rect 1879 15242 2480 15298
rect 1160 15241 2480 15242
rect 0 15234 2480 15241
rect 2544 15234 2608 15298
rect 2672 15234 3472 15298
rect 3536 15234 3600 15298
rect 3664 15234 4464 15298
rect 4528 15234 4592 15298
rect 4656 15297 6448 15298
rect 4656 15234 5456 15297
rect 0 15233 5456 15234
rect 5520 15233 5584 15297
rect 5648 15234 6448 15297
rect 6512 15234 6576 15298
rect 6640 15234 7440 15298
rect 7504 15234 7568 15298
rect 7632 15234 8432 15298
rect 8496 15234 8560 15298
rect 8624 15234 9424 15298
rect 9488 15234 9552 15298
rect 9616 15234 10416 15298
rect 10480 15234 10544 15298
rect 10608 15234 11408 15298
rect 11472 15234 11536 15298
rect 11600 15234 12400 15298
rect 12464 15234 12528 15298
rect 12592 15234 13392 15298
rect 13456 15234 13520 15298
rect 13584 15246 13777 15298
rect 13841 15246 13863 15310
rect 13927 15246 13949 15310
rect 14013 15246 14035 15310
rect 14099 15246 14121 15310
rect 14185 15246 14207 15310
rect 14271 15246 14293 15310
rect 14357 15246 14379 15310
rect 14443 15246 14465 15310
rect 14529 15246 15000 15310
rect 13584 15234 15000 15246
rect 5648 15233 15000 15234
rect 0 15230 15000 15233
rect 0 15226 13777 15230
rect 0 15224 1287 15226
rect 0 15160 456 15224
rect 520 15160 536 15224
rect 600 15160 616 15224
rect 680 15160 696 15224
rect 760 15160 776 15224
rect 840 15160 856 15224
rect 920 15160 936 15224
rect 1000 15160 1016 15224
rect 1080 15160 1096 15224
rect 1160 15162 1287 15224
rect 1351 15162 1375 15226
rect 1439 15162 1463 15226
rect 1527 15162 1551 15226
rect 1615 15162 1639 15226
rect 1703 15162 1727 15226
rect 1791 15162 1815 15226
rect 1879 15217 13777 15226
rect 1879 15162 2480 15217
rect 1160 15160 2480 15162
rect 0 15153 2480 15160
rect 2544 15153 2608 15217
rect 2672 15153 3472 15217
rect 3536 15153 3600 15217
rect 3664 15153 4464 15217
rect 4528 15153 4592 15217
rect 4656 15216 6448 15217
rect 4656 15153 5456 15216
rect 0 15152 5456 15153
rect 5520 15152 5584 15216
rect 5648 15153 6448 15216
rect 6512 15153 6576 15217
rect 6640 15153 7440 15217
rect 7504 15153 7568 15217
rect 7632 15153 8432 15217
rect 8496 15153 8560 15217
rect 8624 15153 9424 15217
rect 9488 15153 9552 15217
rect 9616 15153 10416 15217
rect 10480 15153 10544 15217
rect 10608 15153 11408 15217
rect 11472 15153 11536 15217
rect 11600 15153 12400 15217
rect 12464 15153 12528 15217
rect 12592 15153 13392 15217
rect 13456 15153 13520 15217
rect 13584 15166 13777 15217
rect 13841 15166 13863 15230
rect 13927 15166 13949 15230
rect 14013 15166 14035 15230
rect 14099 15166 14121 15230
rect 14185 15166 14207 15230
rect 14271 15166 14293 15230
rect 14357 15166 14379 15230
rect 14443 15166 14465 15230
rect 14529 15166 15000 15230
rect 13584 15153 15000 15166
rect 5648 15152 15000 15153
rect 0 15149 15000 15152
rect 0 15146 13777 15149
rect 0 15143 1287 15146
rect 0 15079 456 15143
rect 520 15079 536 15143
rect 600 15079 616 15143
rect 680 15079 696 15143
rect 760 15079 776 15143
rect 840 15079 856 15143
rect 920 15079 936 15143
rect 1000 15079 1016 15143
rect 1080 15079 1096 15143
rect 1160 15082 1287 15143
rect 1351 15082 1375 15146
rect 1439 15082 1463 15146
rect 1527 15082 1551 15146
rect 1615 15082 1639 15146
rect 1703 15082 1727 15146
rect 1791 15082 1815 15146
rect 1879 15136 13777 15146
rect 1879 15082 2480 15136
rect 1160 15079 2480 15082
rect 0 15072 2480 15079
rect 2544 15072 2608 15136
rect 2672 15072 3472 15136
rect 3536 15072 3600 15136
rect 3664 15072 4464 15136
rect 4528 15072 4592 15136
rect 4656 15135 6448 15136
rect 4656 15072 5456 15135
rect 0 15071 5456 15072
rect 5520 15071 5584 15135
rect 5648 15072 6448 15135
rect 6512 15072 6576 15136
rect 6640 15072 7440 15136
rect 7504 15072 7568 15136
rect 7632 15072 8432 15136
rect 8496 15072 8560 15136
rect 8624 15072 9424 15136
rect 9488 15072 9552 15136
rect 9616 15072 10416 15136
rect 10480 15072 10544 15136
rect 10608 15072 11408 15136
rect 11472 15072 11536 15136
rect 11600 15072 12400 15136
rect 12464 15072 12528 15136
rect 12592 15072 13392 15136
rect 13456 15072 13520 15136
rect 13584 15085 13777 15136
rect 13841 15085 13863 15149
rect 13927 15085 13949 15149
rect 14013 15085 14035 15149
rect 14099 15085 14121 15149
rect 14185 15085 14207 15149
rect 14271 15085 14293 15149
rect 14357 15085 14379 15149
rect 14443 15085 14465 15149
rect 14529 15085 15000 15149
rect 13584 15072 15000 15085
rect 5648 15071 15000 15072
rect 0 15068 15000 15071
rect 0 15066 13777 15068
rect 0 15062 1287 15066
rect 0 14998 456 15062
rect 520 14998 536 15062
rect 600 14998 616 15062
rect 680 14998 696 15062
rect 760 14998 776 15062
rect 840 14998 856 15062
rect 920 14998 936 15062
rect 1000 14998 1016 15062
rect 1080 14998 1096 15062
rect 1160 15002 1287 15062
rect 1351 15002 1375 15066
rect 1439 15002 1463 15066
rect 1527 15002 1551 15066
rect 1615 15002 1639 15066
rect 1703 15002 1727 15066
rect 1791 15002 1815 15066
rect 1879 15055 13777 15066
rect 1879 15002 2480 15055
rect 1160 14998 2480 15002
rect 0 14991 2480 14998
rect 2544 14991 2608 15055
rect 2672 14991 3472 15055
rect 3536 14991 3600 15055
rect 3664 14991 4464 15055
rect 4528 14991 4592 15055
rect 4656 15054 6448 15055
rect 4656 14991 5456 15054
rect 0 14990 5456 14991
rect 5520 14990 5584 15054
rect 5648 14991 6448 15054
rect 6512 14991 6576 15055
rect 6640 14991 7440 15055
rect 7504 14991 7568 15055
rect 7632 14991 8432 15055
rect 8496 14991 8560 15055
rect 8624 14991 9424 15055
rect 9488 14991 9552 15055
rect 9616 14991 10416 15055
rect 10480 14991 10544 15055
rect 10608 14991 11408 15055
rect 11472 14991 11536 15055
rect 11600 14991 12400 15055
rect 12464 14991 12528 15055
rect 12592 14991 13392 15055
rect 13456 14991 13520 15055
rect 13584 15004 13777 15055
rect 13841 15004 13863 15068
rect 13927 15004 13949 15068
rect 14013 15004 14035 15068
rect 14099 15004 14121 15068
rect 14185 15004 14207 15068
rect 14271 15004 14293 15068
rect 14357 15004 14379 15068
rect 14443 15004 14465 15068
rect 14529 15004 15000 15068
rect 13584 14991 15000 15004
rect 5648 14990 15000 14991
rect 0 14987 15000 14990
rect 0 14986 13777 14987
rect 0 14981 1287 14986
rect 0 14917 456 14981
rect 520 14917 536 14981
rect 600 14917 616 14981
rect 680 14917 696 14981
rect 760 14917 776 14981
rect 840 14917 856 14981
rect 920 14917 936 14981
rect 1000 14917 1016 14981
rect 1080 14917 1096 14981
rect 1160 14922 1287 14981
rect 1351 14922 1375 14986
rect 1439 14922 1463 14986
rect 1527 14922 1551 14986
rect 1615 14922 1639 14986
rect 1703 14922 1727 14986
rect 1791 14922 1815 14986
rect 1879 14974 13777 14986
rect 1879 14922 2480 14974
rect 1160 14917 2480 14922
rect 0 14910 2480 14917
rect 2544 14910 2608 14974
rect 2672 14910 3472 14974
rect 3536 14910 3600 14974
rect 3664 14910 4464 14974
rect 4528 14910 4592 14974
rect 4656 14973 6448 14974
rect 4656 14910 5456 14973
rect 0 14909 5456 14910
rect 5520 14909 5584 14973
rect 5648 14910 6448 14973
rect 6512 14910 6576 14974
rect 6640 14910 7440 14974
rect 7504 14910 7568 14974
rect 7632 14910 8432 14974
rect 8496 14910 8560 14974
rect 8624 14910 9424 14974
rect 9488 14910 9552 14974
rect 9616 14910 10416 14974
rect 10480 14910 10544 14974
rect 10608 14910 11408 14974
rect 11472 14910 11536 14974
rect 11600 14910 12400 14974
rect 12464 14910 12528 14974
rect 12592 14910 13392 14974
rect 13456 14910 13520 14974
rect 13584 14923 13777 14974
rect 13841 14923 13863 14987
rect 13927 14923 13949 14987
rect 14013 14923 14035 14987
rect 14099 14923 14121 14987
rect 14185 14923 14207 14987
rect 14271 14923 14293 14987
rect 14357 14923 14379 14987
rect 14443 14923 14465 14987
rect 14529 14923 15000 14987
rect 13584 14910 15000 14923
rect 5648 14909 15000 14910
rect 0 14906 15000 14909
rect 0 14900 1287 14906
rect 0 14836 456 14900
rect 520 14836 536 14900
rect 600 14836 616 14900
rect 680 14836 696 14900
rect 760 14836 776 14900
rect 840 14836 856 14900
rect 920 14836 936 14900
rect 1000 14836 1016 14900
rect 1080 14836 1096 14900
rect 1160 14842 1287 14900
rect 1351 14842 1375 14906
rect 1439 14842 1463 14906
rect 1527 14842 1551 14906
rect 1615 14842 1639 14906
rect 1703 14842 1727 14906
rect 1791 14842 1815 14906
rect 1879 14893 13777 14906
rect 1879 14842 2480 14893
rect 1160 14836 2480 14842
rect 0 14829 2480 14836
rect 2544 14829 2608 14893
rect 2672 14829 3472 14893
rect 3536 14829 3600 14893
rect 3664 14829 4464 14893
rect 4528 14829 4592 14893
rect 4656 14892 6448 14893
rect 4656 14829 5456 14892
rect 0 14828 5456 14829
rect 5520 14828 5584 14892
rect 5648 14829 6448 14892
rect 6512 14829 6576 14893
rect 6640 14829 7440 14893
rect 7504 14829 7568 14893
rect 7632 14829 8432 14893
rect 8496 14829 8560 14893
rect 8624 14829 9424 14893
rect 9488 14829 9552 14893
rect 9616 14829 10416 14893
rect 10480 14829 10544 14893
rect 10608 14829 11408 14893
rect 11472 14829 11536 14893
rect 11600 14829 12400 14893
rect 12464 14829 12528 14893
rect 12592 14829 13392 14893
rect 13456 14829 13520 14893
rect 13584 14842 13777 14893
rect 13841 14842 13863 14906
rect 13927 14842 13949 14906
rect 14013 14842 14035 14906
rect 14099 14842 14121 14906
rect 14185 14842 14207 14906
rect 14271 14842 14293 14906
rect 14357 14842 14379 14906
rect 14443 14842 14465 14906
rect 14529 14842 15000 14906
rect 13584 14829 15000 14842
rect 5648 14828 15000 14829
rect 0 14826 15000 14828
rect 0 14819 1287 14826
rect 0 14755 456 14819
rect 520 14755 536 14819
rect 600 14755 616 14819
rect 680 14755 696 14819
rect 760 14755 776 14819
rect 840 14755 856 14819
rect 920 14755 936 14819
rect 1000 14755 1016 14819
rect 1080 14755 1096 14819
rect 1160 14762 1287 14819
rect 1351 14762 1375 14826
rect 1439 14762 1463 14826
rect 1527 14762 1551 14826
rect 1615 14762 1639 14826
rect 1703 14762 1727 14826
rect 1791 14762 1815 14826
rect 1879 14825 15000 14826
rect 1879 14812 13777 14825
rect 1879 14762 2480 14812
rect 1160 14755 2480 14762
rect 0 14748 2480 14755
rect 2544 14748 2608 14812
rect 2672 14748 3472 14812
rect 3536 14748 3600 14812
rect 3664 14748 4464 14812
rect 4528 14748 4592 14812
rect 4656 14811 6448 14812
rect 4656 14748 5456 14811
rect 0 14747 5456 14748
rect 5520 14747 5584 14811
rect 5648 14748 6448 14811
rect 6512 14748 6576 14812
rect 6640 14748 7440 14812
rect 7504 14748 7568 14812
rect 7632 14748 8432 14812
rect 8496 14748 8560 14812
rect 8624 14748 9424 14812
rect 9488 14748 9552 14812
rect 9616 14748 10416 14812
rect 10480 14748 10544 14812
rect 10608 14748 11408 14812
rect 11472 14748 11536 14812
rect 11600 14748 12400 14812
rect 12464 14748 12528 14812
rect 12592 14748 13392 14812
rect 13456 14748 13520 14812
rect 13584 14761 13777 14812
rect 13841 14761 13863 14825
rect 13927 14761 13949 14825
rect 14013 14761 14035 14825
rect 14099 14761 14121 14825
rect 14185 14761 14207 14825
rect 14271 14761 14293 14825
rect 14357 14761 14379 14825
rect 14443 14761 14465 14825
rect 14529 14761 15000 14825
rect 13584 14748 15000 14761
rect 5648 14747 15000 14748
rect 0 14746 15000 14747
rect 0 14738 1287 14746
rect 0 14674 456 14738
rect 520 14674 536 14738
rect 600 14674 616 14738
rect 680 14674 696 14738
rect 760 14674 776 14738
rect 840 14674 856 14738
rect 920 14674 936 14738
rect 1000 14674 1016 14738
rect 1080 14674 1096 14738
rect 1160 14682 1287 14738
rect 1351 14682 1375 14746
rect 1439 14682 1463 14746
rect 1527 14682 1551 14746
rect 1615 14682 1639 14746
rect 1703 14682 1727 14746
rect 1791 14682 1815 14746
rect 1879 14744 15000 14746
rect 1879 14731 13777 14744
rect 1879 14682 2480 14731
rect 1160 14674 2480 14682
rect 0 14667 2480 14674
rect 2544 14667 2608 14731
rect 2672 14667 3472 14731
rect 3536 14667 3600 14731
rect 3664 14667 4464 14731
rect 4528 14667 4592 14731
rect 4656 14730 6448 14731
rect 4656 14667 5456 14730
rect 0 14666 5456 14667
rect 5520 14666 5584 14730
rect 5648 14667 6448 14730
rect 6512 14667 6576 14731
rect 6640 14667 7440 14731
rect 7504 14667 7568 14731
rect 7632 14667 8432 14731
rect 8496 14667 8560 14731
rect 8624 14667 9424 14731
rect 9488 14667 9552 14731
rect 9616 14667 10416 14731
rect 10480 14667 10544 14731
rect 10608 14667 11408 14731
rect 11472 14667 11536 14731
rect 11600 14667 12400 14731
rect 12464 14667 12528 14731
rect 12592 14667 13392 14731
rect 13456 14667 13520 14731
rect 13584 14680 13777 14731
rect 13841 14680 13863 14744
rect 13927 14680 13949 14744
rect 14013 14680 14035 14744
rect 14099 14680 14121 14744
rect 14185 14680 14207 14744
rect 14271 14680 14293 14744
rect 14357 14680 14379 14744
rect 14443 14680 14465 14744
rect 14529 14680 15000 14744
rect 13584 14667 15000 14680
rect 5648 14666 15000 14667
rect 0 14657 1287 14666
rect 0 14593 456 14657
rect 520 14593 536 14657
rect 600 14593 616 14657
rect 680 14593 696 14657
rect 760 14593 776 14657
rect 840 14593 856 14657
rect 920 14593 936 14657
rect 1000 14593 1016 14657
rect 1080 14593 1096 14657
rect 1160 14602 1287 14657
rect 1351 14602 1375 14666
rect 1439 14602 1463 14666
rect 1527 14602 1551 14666
rect 1615 14602 1639 14666
rect 1703 14602 1727 14666
rect 1791 14602 1815 14666
rect 1879 14663 15000 14666
rect 1879 14650 13777 14663
rect 1879 14602 2480 14650
rect 1160 14593 2480 14602
rect 0 14586 2480 14593
rect 2544 14586 2608 14650
rect 2672 14586 3472 14650
rect 3536 14586 3600 14650
rect 3664 14586 4464 14650
rect 4528 14586 4592 14650
rect 4656 14649 6448 14650
rect 4656 14586 5456 14649
rect 0 14576 1287 14586
rect 0 14512 456 14576
rect 520 14512 536 14576
rect 600 14512 616 14576
rect 680 14512 696 14576
rect 760 14512 776 14576
rect 840 14512 856 14576
rect 920 14512 936 14576
rect 1000 14512 1016 14576
rect 1080 14512 1096 14576
rect 1160 14522 1287 14576
rect 1351 14522 1375 14586
rect 1439 14522 1463 14586
rect 1527 14522 1551 14586
rect 1615 14522 1639 14586
rect 1703 14522 1727 14586
rect 1791 14522 1815 14586
rect 1879 14585 5456 14586
rect 5520 14585 5584 14649
rect 5648 14586 6448 14649
rect 6512 14586 6576 14650
rect 6640 14586 7440 14650
rect 7504 14586 7568 14650
rect 7632 14586 8432 14650
rect 8496 14586 8560 14650
rect 8624 14586 9424 14650
rect 9488 14586 9552 14650
rect 9616 14586 10416 14650
rect 10480 14586 10544 14650
rect 10608 14586 11408 14650
rect 11472 14586 11536 14650
rect 11600 14586 12400 14650
rect 12464 14586 12528 14650
rect 12592 14586 13392 14650
rect 13456 14586 13520 14650
rect 13584 14599 13777 14650
rect 13841 14599 13863 14663
rect 13927 14599 13949 14663
rect 14013 14599 14035 14663
rect 14099 14599 14121 14663
rect 14185 14599 14207 14663
rect 14271 14599 14293 14663
rect 14357 14599 14379 14663
rect 14443 14599 14465 14663
rect 14529 14599 15000 14663
rect 13584 14586 15000 14599
rect 5648 14585 15000 14586
rect 1879 14582 15000 14585
rect 1879 14569 13777 14582
rect 1879 14522 2480 14569
rect 1160 14512 2480 14522
rect 0 14505 2480 14512
rect 2544 14505 2608 14569
rect 2672 14505 3472 14569
rect 3536 14505 3600 14569
rect 3664 14505 4464 14569
rect 4528 14505 4592 14569
rect 4656 14568 6448 14569
rect 4656 14505 5456 14568
rect 0 14495 1287 14505
rect 0 14431 456 14495
rect 520 14431 536 14495
rect 600 14431 616 14495
rect 680 14431 696 14495
rect 760 14431 776 14495
rect 840 14431 856 14495
rect 920 14431 936 14495
rect 1000 14431 1016 14495
rect 1080 14431 1096 14495
rect 1160 14441 1287 14495
rect 1351 14441 1375 14505
rect 1439 14441 1463 14505
rect 1527 14441 1551 14505
rect 1615 14441 1639 14505
rect 1703 14441 1727 14505
rect 1791 14441 1815 14505
rect 1879 14504 5456 14505
rect 5520 14504 5584 14568
rect 5648 14505 6448 14568
rect 6512 14505 6576 14569
rect 6640 14505 7440 14569
rect 7504 14505 7568 14569
rect 7632 14505 8432 14569
rect 8496 14505 8560 14569
rect 8624 14505 9424 14569
rect 9488 14505 9552 14569
rect 9616 14505 10416 14569
rect 10480 14505 10544 14569
rect 10608 14505 11408 14569
rect 11472 14505 11536 14569
rect 11600 14505 12400 14569
rect 12464 14505 12528 14569
rect 12592 14505 13392 14569
rect 13456 14505 13520 14569
rect 13584 14518 13777 14569
rect 13841 14518 13863 14582
rect 13927 14518 13949 14582
rect 14013 14518 14035 14582
rect 14099 14518 14121 14582
rect 14185 14518 14207 14582
rect 14271 14518 14293 14582
rect 14357 14518 14379 14582
rect 14443 14518 14465 14582
rect 14529 14518 15000 14582
rect 13584 14505 15000 14518
rect 5648 14504 15000 14505
rect 1879 14501 15000 14504
rect 1879 14488 13777 14501
rect 1879 14441 2480 14488
rect 1160 14431 2480 14441
rect 0 14424 2480 14431
rect 2544 14424 2608 14488
rect 2672 14424 3472 14488
rect 3536 14424 3600 14488
rect 3664 14424 4464 14488
rect 4528 14424 4592 14488
rect 4656 14487 6448 14488
rect 4656 14424 5456 14487
rect 0 14414 1287 14424
rect 0 14350 456 14414
rect 520 14350 536 14414
rect 600 14350 616 14414
rect 680 14350 696 14414
rect 760 14350 776 14414
rect 840 14350 856 14414
rect 920 14350 936 14414
rect 1000 14350 1016 14414
rect 1080 14350 1096 14414
rect 1160 14360 1287 14414
rect 1351 14360 1375 14424
rect 1439 14360 1463 14424
rect 1527 14360 1551 14424
rect 1615 14360 1639 14424
rect 1703 14360 1727 14424
rect 1791 14360 1815 14424
rect 1879 14423 5456 14424
rect 5520 14423 5584 14487
rect 5648 14424 6448 14487
rect 6512 14424 6576 14488
rect 6640 14424 7440 14488
rect 7504 14424 7568 14488
rect 7632 14424 8432 14488
rect 8496 14424 8560 14488
rect 8624 14424 9424 14488
rect 9488 14424 9552 14488
rect 9616 14424 10416 14488
rect 10480 14424 10544 14488
rect 10608 14424 11408 14488
rect 11472 14424 11536 14488
rect 11600 14424 12400 14488
rect 12464 14424 12528 14488
rect 12592 14424 13392 14488
rect 13456 14424 13520 14488
rect 13584 14437 13777 14488
rect 13841 14437 13863 14501
rect 13927 14437 13949 14501
rect 14013 14437 14035 14501
rect 14099 14437 14121 14501
rect 14185 14437 14207 14501
rect 14271 14437 14293 14501
rect 14357 14437 14379 14501
rect 14443 14437 14465 14501
rect 14529 14437 15000 14501
rect 13584 14424 15000 14437
rect 5648 14423 15000 14424
rect 1879 14420 15000 14423
rect 1879 14407 13777 14420
rect 1879 14360 2480 14407
rect 1160 14350 2480 14360
rect 0 14343 2480 14350
rect 2544 14343 2608 14407
rect 2672 14343 3472 14407
rect 3536 14343 3600 14407
rect 3664 14343 4464 14407
rect 4528 14343 4592 14407
rect 4656 14406 6448 14407
rect 4656 14343 5456 14406
rect 0 14333 1287 14343
rect 0 14269 456 14333
rect 520 14269 536 14333
rect 600 14269 616 14333
rect 680 14269 696 14333
rect 760 14269 776 14333
rect 840 14269 856 14333
rect 920 14269 936 14333
rect 1000 14269 1016 14333
rect 1080 14269 1096 14333
rect 1160 14279 1287 14333
rect 1351 14279 1375 14343
rect 1439 14279 1463 14343
rect 1527 14279 1551 14343
rect 1615 14279 1639 14343
rect 1703 14279 1727 14343
rect 1791 14279 1815 14343
rect 1879 14342 5456 14343
rect 5520 14342 5584 14406
rect 5648 14343 6448 14406
rect 6512 14343 6576 14407
rect 6640 14343 7440 14407
rect 7504 14343 7568 14407
rect 7632 14343 8432 14407
rect 8496 14343 8560 14407
rect 8624 14343 9424 14407
rect 9488 14343 9552 14407
rect 9616 14343 10416 14407
rect 10480 14343 10544 14407
rect 10608 14343 11408 14407
rect 11472 14343 11536 14407
rect 11600 14343 12400 14407
rect 12464 14343 12528 14407
rect 12592 14343 13392 14407
rect 13456 14343 13520 14407
rect 13584 14356 13777 14407
rect 13841 14356 13863 14420
rect 13927 14356 13949 14420
rect 14013 14356 14035 14420
rect 14099 14356 14121 14420
rect 14185 14356 14207 14420
rect 14271 14356 14293 14420
rect 14357 14356 14379 14420
rect 14443 14356 14465 14420
rect 14529 14356 15000 14420
rect 13584 14343 15000 14356
rect 5648 14342 15000 14343
rect 1879 14339 15000 14342
rect 1879 14326 13777 14339
rect 1879 14279 2480 14326
rect 1160 14269 2480 14279
rect 0 14262 2480 14269
rect 2544 14262 2608 14326
rect 2672 14262 3472 14326
rect 3536 14262 3600 14326
rect 3664 14262 4464 14326
rect 4528 14262 4592 14326
rect 4656 14325 6448 14326
rect 4656 14262 5456 14325
rect 0 14252 1287 14262
rect 0 14188 456 14252
rect 520 14188 536 14252
rect 600 14188 616 14252
rect 680 14188 696 14252
rect 760 14188 776 14252
rect 840 14188 856 14252
rect 920 14188 936 14252
rect 1000 14188 1016 14252
rect 1080 14188 1096 14252
rect 1160 14198 1287 14252
rect 1351 14198 1375 14262
rect 1439 14198 1463 14262
rect 1527 14198 1551 14262
rect 1615 14198 1639 14262
rect 1703 14198 1727 14262
rect 1791 14198 1815 14262
rect 1879 14261 5456 14262
rect 5520 14261 5584 14325
rect 5648 14262 6448 14325
rect 6512 14262 6576 14326
rect 6640 14262 7440 14326
rect 7504 14262 7568 14326
rect 7632 14262 8432 14326
rect 8496 14262 8560 14326
rect 8624 14262 9424 14326
rect 9488 14262 9552 14326
rect 9616 14262 10416 14326
rect 10480 14262 10544 14326
rect 10608 14262 11408 14326
rect 11472 14262 11536 14326
rect 11600 14262 12400 14326
rect 12464 14262 12528 14326
rect 12592 14262 13392 14326
rect 13456 14262 13520 14326
rect 13584 14275 13777 14326
rect 13841 14275 13863 14339
rect 13927 14275 13949 14339
rect 14013 14275 14035 14339
rect 14099 14275 14121 14339
rect 14185 14275 14207 14339
rect 14271 14275 14293 14339
rect 14357 14275 14379 14339
rect 14443 14275 14465 14339
rect 14529 14275 15000 14339
rect 13584 14262 15000 14275
rect 5648 14261 15000 14262
rect 1879 14258 15000 14261
rect 1879 14245 13777 14258
rect 1879 14198 2480 14245
rect 1160 14188 2480 14198
rect 0 14181 2480 14188
rect 2544 14181 2608 14245
rect 2672 14181 3472 14245
rect 3536 14181 3600 14245
rect 3664 14181 4464 14245
rect 4528 14181 4592 14245
rect 4656 14244 6448 14245
rect 4656 14181 5456 14244
rect 0 14171 1287 14181
rect 0 14107 456 14171
rect 520 14107 536 14171
rect 600 14107 616 14171
rect 680 14107 696 14171
rect 760 14107 776 14171
rect 840 14107 856 14171
rect 920 14107 936 14171
rect 1000 14107 1016 14171
rect 1080 14107 1096 14171
rect 1160 14117 1287 14171
rect 1351 14117 1375 14181
rect 1439 14117 1463 14181
rect 1527 14117 1551 14181
rect 1615 14117 1639 14181
rect 1703 14117 1727 14181
rect 1791 14117 1815 14181
rect 1879 14180 5456 14181
rect 5520 14180 5584 14244
rect 5648 14181 6448 14244
rect 6512 14181 6576 14245
rect 6640 14181 7440 14245
rect 7504 14181 7568 14245
rect 7632 14181 8432 14245
rect 8496 14181 8560 14245
rect 8624 14181 9424 14245
rect 9488 14181 9552 14245
rect 9616 14181 10416 14245
rect 10480 14181 10544 14245
rect 10608 14181 11408 14245
rect 11472 14181 11536 14245
rect 11600 14181 12400 14245
rect 12464 14181 12528 14245
rect 12592 14181 13392 14245
rect 13456 14181 13520 14245
rect 13584 14194 13777 14245
rect 13841 14194 13863 14258
rect 13927 14194 13949 14258
rect 14013 14194 14035 14258
rect 14099 14194 14121 14258
rect 14185 14194 14207 14258
rect 14271 14194 14293 14258
rect 14357 14194 14379 14258
rect 14443 14194 14465 14258
rect 14529 14194 15000 14258
rect 13584 14181 15000 14194
rect 5648 14180 15000 14181
rect 1879 14177 15000 14180
rect 1879 14164 13777 14177
rect 1879 14117 2480 14164
rect 1160 14107 2480 14117
rect 0 14100 2480 14107
rect 2544 14100 2608 14164
rect 2672 14100 3472 14164
rect 3536 14100 3600 14164
rect 3664 14100 4464 14164
rect 4528 14100 4592 14164
rect 4656 14163 6448 14164
rect 4656 14100 5456 14163
rect 0 14090 1287 14100
rect 0 14026 456 14090
rect 520 14026 536 14090
rect 600 14026 616 14090
rect 680 14026 696 14090
rect 760 14026 776 14090
rect 840 14026 856 14090
rect 920 14026 936 14090
rect 1000 14026 1016 14090
rect 1080 14026 1096 14090
rect 1160 14036 1287 14090
rect 1351 14036 1375 14100
rect 1439 14036 1463 14100
rect 1527 14036 1551 14100
rect 1615 14036 1639 14100
rect 1703 14036 1727 14100
rect 1791 14036 1815 14100
rect 1879 14099 5456 14100
rect 5520 14099 5584 14163
rect 5648 14100 6448 14163
rect 6512 14100 6576 14164
rect 6640 14100 7440 14164
rect 7504 14100 7568 14164
rect 7632 14100 8432 14164
rect 8496 14100 8560 14164
rect 8624 14100 9424 14164
rect 9488 14100 9552 14164
rect 9616 14100 10416 14164
rect 10480 14100 10544 14164
rect 10608 14100 11408 14164
rect 11472 14100 11536 14164
rect 11600 14100 12400 14164
rect 12464 14100 12528 14164
rect 12592 14100 13392 14164
rect 13456 14100 13520 14164
rect 13584 14113 13777 14164
rect 13841 14113 13863 14177
rect 13927 14113 13949 14177
rect 14013 14113 14035 14177
rect 14099 14113 14121 14177
rect 14185 14113 14207 14177
rect 14271 14113 14293 14177
rect 14357 14113 14379 14177
rect 14443 14113 14465 14177
rect 14529 14113 15000 14177
rect 13584 14100 15000 14113
rect 5648 14099 15000 14100
rect 1879 14096 15000 14099
rect 1879 14083 13777 14096
rect 1879 14036 2480 14083
rect 1160 14026 2480 14036
rect 0 14019 2480 14026
rect 2544 14019 2608 14083
rect 2672 14019 3472 14083
rect 3536 14019 3600 14083
rect 3664 14019 4464 14083
rect 4528 14019 4592 14083
rect 4656 14082 6448 14083
rect 4656 14019 5456 14082
rect 0 14009 1287 14019
rect 0 13945 456 14009
rect 520 13945 536 14009
rect 600 13945 616 14009
rect 680 13945 696 14009
rect 760 13945 776 14009
rect 840 13945 856 14009
rect 920 13945 936 14009
rect 1000 13945 1016 14009
rect 1080 13945 1096 14009
rect 1160 13955 1287 14009
rect 1351 13955 1375 14019
rect 1439 13955 1463 14019
rect 1527 13955 1551 14019
rect 1615 13955 1639 14019
rect 1703 13955 1727 14019
rect 1791 13955 1815 14019
rect 1879 14018 5456 14019
rect 5520 14018 5584 14082
rect 5648 14019 6448 14082
rect 6512 14019 6576 14083
rect 6640 14019 7440 14083
rect 7504 14019 7568 14083
rect 7632 14019 8432 14083
rect 8496 14019 8560 14083
rect 8624 14019 9424 14083
rect 9488 14019 9552 14083
rect 9616 14019 10416 14083
rect 10480 14019 10544 14083
rect 10608 14019 11408 14083
rect 11472 14019 11536 14083
rect 11600 14019 12400 14083
rect 12464 14019 12528 14083
rect 12592 14019 13392 14083
rect 13456 14019 13520 14083
rect 13584 14032 13777 14083
rect 13841 14032 13863 14096
rect 13927 14032 13949 14096
rect 14013 14032 14035 14096
rect 14099 14032 14121 14096
rect 14185 14032 14207 14096
rect 14271 14032 14293 14096
rect 14357 14032 14379 14096
rect 14443 14032 14465 14096
rect 14529 14032 15000 14096
rect 13584 14019 15000 14032
rect 5648 14018 15000 14019
rect 1879 14015 15000 14018
rect 1879 14002 13777 14015
rect 1879 13955 2480 14002
rect 1160 13945 2480 13955
rect 0 13938 2480 13945
rect 2544 13938 2608 14002
rect 2672 13938 3472 14002
rect 3536 13938 3600 14002
rect 3664 13938 4464 14002
rect 4528 13938 4592 14002
rect 4656 14001 6448 14002
rect 4656 13938 5456 14001
rect 0 13928 1287 13938
rect 0 13864 456 13928
rect 520 13864 536 13928
rect 600 13864 616 13928
rect 680 13864 696 13928
rect 760 13864 776 13928
rect 840 13864 856 13928
rect 920 13864 936 13928
rect 1000 13864 1016 13928
rect 1080 13864 1096 13928
rect 1160 13874 1287 13928
rect 1351 13874 1375 13938
rect 1439 13874 1463 13938
rect 1527 13874 1551 13938
rect 1615 13874 1639 13938
rect 1703 13874 1727 13938
rect 1791 13874 1815 13938
rect 1879 13937 5456 13938
rect 5520 13937 5584 14001
rect 5648 13938 6448 14001
rect 6512 13938 6576 14002
rect 6640 13938 7440 14002
rect 7504 13938 7568 14002
rect 7632 13938 8432 14002
rect 8496 13938 8560 14002
rect 8624 13938 9424 14002
rect 9488 13938 9552 14002
rect 9616 13938 10416 14002
rect 10480 13938 10544 14002
rect 10608 13938 11408 14002
rect 11472 13938 11536 14002
rect 11600 13938 12400 14002
rect 12464 13938 12528 14002
rect 12592 13938 13392 14002
rect 13456 13938 13520 14002
rect 13584 13951 13777 14002
rect 13841 13951 13863 14015
rect 13927 13951 13949 14015
rect 14013 13951 14035 14015
rect 14099 13951 14121 14015
rect 14185 13951 14207 14015
rect 14271 13951 14293 14015
rect 14357 13951 14379 14015
rect 14443 13951 14465 14015
rect 14529 13951 15000 14015
rect 13584 13938 15000 13951
rect 5648 13937 15000 13938
rect 1879 13934 15000 13937
rect 1879 13921 13777 13934
rect 1879 13874 2480 13921
rect 1160 13864 2480 13874
rect 0 13857 2480 13864
rect 2544 13857 2608 13921
rect 2672 13857 3472 13921
rect 3536 13857 3600 13921
rect 3664 13857 4464 13921
rect 4528 13857 4592 13921
rect 4656 13920 6448 13921
rect 4656 13857 5456 13920
rect 0 13847 1287 13857
rect 0 13783 456 13847
rect 520 13783 536 13847
rect 600 13783 616 13847
rect 680 13783 696 13847
rect 760 13783 776 13847
rect 840 13783 856 13847
rect 920 13783 936 13847
rect 1000 13783 1016 13847
rect 1080 13783 1096 13847
rect 1160 13793 1287 13847
rect 1351 13793 1375 13857
rect 1439 13793 1463 13857
rect 1527 13793 1551 13857
rect 1615 13793 1639 13857
rect 1703 13793 1727 13857
rect 1791 13793 1815 13857
rect 1879 13856 5456 13857
rect 5520 13856 5584 13920
rect 5648 13857 6448 13920
rect 6512 13857 6576 13921
rect 6640 13857 7440 13921
rect 7504 13857 7568 13921
rect 7632 13857 8432 13921
rect 8496 13857 8560 13921
rect 8624 13857 9424 13921
rect 9488 13857 9552 13921
rect 9616 13857 10416 13921
rect 10480 13857 10544 13921
rect 10608 13857 11408 13921
rect 11472 13857 11536 13921
rect 11600 13857 12400 13921
rect 12464 13857 12528 13921
rect 12592 13857 13392 13921
rect 13456 13857 13520 13921
rect 13584 13870 13777 13921
rect 13841 13870 13863 13934
rect 13927 13870 13949 13934
rect 14013 13870 14035 13934
rect 14099 13870 14121 13934
rect 14185 13870 14207 13934
rect 14271 13870 14293 13934
rect 14357 13870 14379 13934
rect 14443 13870 14465 13934
rect 14529 13870 15000 13934
rect 13584 13857 15000 13870
rect 5648 13856 15000 13857
rect 1879 13853 15000 13856
rect 1879 13840 13777 13853
rect 1879 13793 2480 13840
rect 1160 13783 2480 13793
rect 0 13776 2480 13783
rect 2544 13776 2608 13840
rect 2672 13776 3472 13840
rect 3536 13776 3600 13840
rect 3664 13776 4464 13840
rect 4528 13776 4592 13840
rect 4656 13839 6448 13840
rect 4656 13776 5456 13839
rect 0 13766 1287 13776
rect 0 13702 456 13766
rect 520 13702 536 13766
rect 600 13702 616 13766
rect 680 13702 696 13766
rect 760 13702 776 13766
rect 840 13702 856 13766
rect 920 13702 936 13766
rect 1000 13702 1016 13766
rect 1080 13702 1096 13766
rect 1160 13712 1287 13766
rect 1351 13712 1375 13776
rect 1439 13712 1463 13776
rect 1527 13712 1551 13776
rect 1615 13712 1639 13776
rect 1703 13712 1727 13776
rect 1791 13712 1815 13776
rect 1879 13775 5456 13776
rect 5520 13775 5584 13839
rect 5648 13776 6448 13839
rect 6512 13776 6576 13840
rect 6640 13776 7440 13840
rect 7504 13776 7568 13840
rect 7632 13776 8432 13840
rect 8496 13776 8560 13840
rect 8624 13776 9424 13840
rect 9488 13776 9552 13840
rect 9616 13776 10416 13840
rect 10480 13776 10544 13840
rect 10608 13776 11408 13840
rect 11472 13776 11536 13840
rect 11600 13776 12400 13840
rect 12464 13776 12528 13840
rect 12592 13776 13392 13840
rect 13456 13776 13520 13840
rect 13584 13789 13777 13840
rect 13841 13789 13863 13853
rect 13927 13789 13949 13853
rect 14013 13789 14035 13853
rect 14099 13789 14121 13853
rect 14185 13789 14207 13853
rect 14271 13789 14293 13853
rect 14357 13789 14379 13853
rect 14443 13789 14465 13853
rect 14529 13789 15000 13853
rect 13584 13776 15000 13789
rect 5648 13775 15000 13776
rect 1879 13772 15000 13775
rect 1879 13759 13777 13772
rect 1879 13712 2480 13759
rect 1160 13702 2480 13712
rect 0 13695 2480 13702
rect 2544 13695 2608 13759
rect 2672 13695 3472 13759
rect 3536 13695 3600 13759
rect 3664 13695 4464 13759
rect 4528 13695 4592 13759
rect 4656 13758 6448 13759
rect 4656 13695 5456 13758
rect 0 13685 1287 13695
rect 0 13621 456 13685
rect 520 13621 536 13685
rect 600 13621 616 13685
rect 680 13621 696 13685
rect 760 13621 776 13685
rect 840 13621 856 13685
rect 920 13621 936 13685
rect 1000 13621 1016 13685
rect 1080 13621 1096 13685
rect 1160 13631 1287 13685
rect 1351 13631 1375 13695
rect 1439 13631 1463 13695
rect 1527 13631 1551 13695
rect 1615 13631 1639 13695
rect 1703 13631 1727 13695
rect 1791 13631 1815 13695
rect 1879 13694 5456 13695
rect 5520 13694 5584 13758
rect 5648 13695 6448 13758
rect 6512 13695 6576 13759
rect 6640 13695 7440 13759
rect 7504 13695 7568 13759
rect 7632 13695 8432 13759
rect 8496 13695 8560 13759
rect 8624 13695 9424 13759
rect 9488 13695 9552 13759
rect 9616 13695 10416 13759
rect 10480 13695 10544 13759
rect 10608 13695 11408 13759
rect 11472 13695 11536 13759
rect 11600 13695 12400 13759
rect 12464 13695 12528 13759
rect 12592 13695 13392 13759
rect 13456 13695 13520 13759
rect 13584 13708 13777 13759
rect 13841 13708 13863 13772
rect 13927 13708 13949 13772
rect 14013 13708 14035 13772
rect 14099 13708 14121 13772
rect 14185 13708 14207 13772
rect 14271 13708 14293 13772
rect 14357 13708 14379 13772
rect 14443 13708 14465 13772
rect 14529 13708 15000 13772
rect 13584 13695 15000 13708
rect 5648 13694 15000 13695
rect 1879 13691 15000 13694
rect 1879 13678 13777 13691
rect 1879 13631 2480 13678
rect 1160 13621 2480 13631
rect 0 13614 2480 13621
rect 2544 13614 2608 13678
rect 2672 13614 3472 13678
rect 3536 13614 3600 13678
rect 3664 13614 4464 13678
rect 4528 13614 4592 13678
rect 4656 13677 6448 13678
rect 4656 13614 5456 13677
rect 0 13613 5456 13614
rect 5520 13613 5584 13677
rect 5648 13614 6448 13677
rect 6512 13614 6576 13678
rect 6640 13614 7440 13678
rect 7504 13614 7568 13678
rect 7632 13614 8432 13678
rect 8496 13614 8560 13678
rect 8624 13614 9424 13678
rect 9488 13614 9552 13678
rect 9616 13614 10416 13678
rect 10480 13614 10544 13678
rect 10608 13614 11408 13678
rect 11472 13614 11536 13678
rect 11600 13614 12400 13678
rect 12464 13614 12528 13678
rect 12592 13614 13392 13678
rect 13456 13614 13520 13678
rect 13584 13627 13777 13678
rect 13841 13627 13863 13691
rect 13927 13627 13949 13691
rect 14013 13627 14035 13691
rect 14099 13627 14121 13691
rect 14185 13627 14207 13691
rect 14271 13627 14293 13691
rect 14357 13627 14379 13691
rect 14443 13627 14465 13691
rect 14529 13627 15000 13691
rect 13584 13614 15000 13627
rect 5648 13613 15000 13614
rect 0 13607 15000 13613
rect 0 12417 15000 13307
rect 0 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 9929 15000 10165
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 15000 9213
rect 0 8835 15000 8847
rect 0 8771 204 8835
rect 268 8771 287 8835
rect 351 8771 370 8835
rect 434 8771 453 8835
rect 517 8771 536 8835
rect 600 8771 618 8835
rect 682 8771 700 8835
rect 764 8771 782 8835
rect 846 8771 864 8835
rect 928 8771 946 8835
rect 1010 8771 1028 8835
rect 1092 8771 1110 8835
rect 1174 8771 1192 8835
rect 1256 8829 15000 8835
rect 1256 8771 8224 8829
rect 0 8765 8224 8771
rect 8288 8765 8305 8829
rect 8369 8765 8386 8829
rect 8450 8765 8466 8829
rect 8530 8765 8546 8829
rect 8610 8765 8626 8829
rect 8690 8765 8706 8829
rect 8770 8765 8786 8829
rect 8850 8765 8866 8829
rect 8930 8765 8946 8829
rect 9010 8765 9026 8829
rect 9090 8765 9106 8829
rect 9170 8765 9186 8829
rect 9250 8765 15000 8829
rect 0 8751 15000 8765
rect 0 8687 204 8751
rect 268 8687 287 8751
rect 351 8687 370 8751
rect 434 8687 453 8751
rect 517 8687 536 8751
rect 600 8687 618 8751
rect 682 8687 700 8751
rect 764 8687 782 8751
rect 846 8687 864 8751
rect 928 8687 946 8751
rect 1010 8687 1028 8751
rect 1092 8687 1110 8751
rect 1174 8687 1192 8751
rect 1256 8745 15000 8751
rect 1256 8687 8224 8745
rect 0 8681 8224 8687
rect 8288 8681 8305 8745
rect 8369 8681 8386 8745
rect 8450 8681 8466 8745
rect 8530 8681 8546 8745
rect 8610 8681 8626 8745
rect 8690 8681 8706 8745
rect 8770 8681 8786 8745
rect 8850 8681 8866 8745
rect 8930 8681 8946 8745
rect 9010 8681 9026 8745
rect 9090 8681 9106 8745
rect 9170 8681 9186 8745
rect 9250 8681 15000 8745
rect 0 8667 15000 8681
rect 0 8603 204 8667
rect 268 8603 287 8667
rect 351 8603 370 8667
rect 434 8603 453 8667
rect 517 8603 536 8667
rect 600 8603 618 8667
rect 682 8603 700 8667
rect 764 8603 782 8667
rect 846 8603 864 8667
rect 928 8603 946 8667
rect 1010 8603 1028 8667
rect 1092 8603 1110 8667
rect 1174 8603 1192 8667
rect 1256 8661 15000 8667
rect 1256 8603 8224 8661
rect 0 8597 8224 8603
rect 8288 8597 8305 8661
rect 8369 8597 8386 8661
rect 8450 8597 8466 8661
rect 8530 8597 8546 8661
rect 8610 8597 8626 8661
rect 8690 8597 8706 8661
rect 8770 8597 8786 8661
rect 8850 8597 8866 8661
rect 8930 8597 8946 8661
rect 9010 8597 9026 8661
rect 9090 8597 9106 8661
rect 9170 8597 9186 8661
rect 9250 8597 15000 8661
rect 0 8583 15000 8597
rect 0 8519 204 8583
rect 268 8519 287 8583
rect 351 8519 370 8583
rect 434 8519 453 8583
rect 517 8519 536 8583
rect 600 8519 618 8583
rect 682 8519 700 8583
rect 764 8519 782 8583
rect 846 8519 864 8583
rect 928 8519 946 8583
rect 1010 8519 1028 8583
rect 1092 8519 1110 8583
rect 1174 8519 1192 8583
rect 1256 8577 15000 8583
rect 1256 8519 8224 8577
rect 0 8513 8224 8519
rect 8288 8513 8305 8577
rect 8369 8513 8386 8577
rect 8450 8513 8466 8577
rect 8530 8513 8546 8577
rect 8610 8513 8626 8577
rect 8690 8513 8706 8577
rect 8770 8513 8786 8577
rect 8850 8513 8866 8577
rect 8930 8513 8946 8577
rect 9010 8513 9026 8577
rect 9090 8513 9106 8577
rect 9170 8513 9186 8577
rect 9250 8513 15000 8577
rect 0 8499 15000 8513
rect 0 8435 204 8499
rect 268 8435 287 8499
rect 351 8435 370 8499
rect 434 8435 453 8499
rect 517 8435 536 8499
rect 600 8435 618 8499
rect 682 8435 700 8499
rect 764 8435 782 8499
rect 846 8435 864 8499
rect 928 8435 946 8499
rect 1010 8435 1028 8499
rect 1092 8435 1110 8499
rect 1174 8435 1192 8499
rect 1256 8493 15000 8499
rect 1256 8435 8224 8493
rect 0 8429 8224 8435
rect 8288 8429 8305 8493
rect 8369 8429 8386 8493
rect 8450 8429 8466 8493
rect 8530 8429 8546 8493
rect 8610 8429 8626 8493
rect 8690 8429 8706 8493
rect 8770 8429 8786 8493
rect 8850 8429 8866 8493
rect 8930 8429 8946 8493
rect 9010 8429 9026 8493
rect 9090 8429 9106 8493
rect 9170 8429 9186 8493
rect 9250 8429 15000 8493
rect 0 8415 15000 8429
rect 0 8351 204 8415
rect 268 8351 287 8415
rect 351 8351 370 8415
rect 434 8351 453 8415
rect 517 8351 536 8415
rect 600 8351 618 8415
rect 682 8351 700 8415
rect 764 8351 782 8415
rect 846 8351 864 8415
rect 928 8351 946 8415
rect 1010 8351 1028 8415
rect 1092 8351 1110 8415
rect 1174 8351 1192 8415
rect 1256 8409 15000 8415
rect 1256 8351 8224 8409
rect 0 8345 8224 8351
rect 8288 8345 8305 8409
rect 8369 8345 8386 8409
rect 8450 8345 8466 8409
rect 8530 8345 8546 8409
rect 8610 8345 8626 8409
rect 8690 8345 8706 8409
rect 8770 8345 8786 8409
rect 8850 8345 8866 8409
rect 8930 8345 8946 8409
rect 9010 8345 9026 8409
rect 9090 8345 9106 8409
rect 9170 8345 9186 8409
rect 9250 8345 15000 8409
rect 0 8331 15000 8345
rect 0 8267 204 8331
rect 268 8267 287 8331
rect 351 8267 370 8331
rect 434 8267 453 8331
rect 517 8267 536 8331
rect 600 8267 618 8331
rect 682 8267 700 8331
rect 764 8267 782 8331
rect 846 8267 864 8331
rect 928 8267 946 8331
rect 1010 8267 1028 8331
rect 1092 8267 1110 8331
rect 1174 8267 1192 8331
rect 1256 8325 15000 8331
rect 1256 8267 8224 8325
rect 0 8261 8224 8267
rect 8288 8261 8305 8325
rect 8369 8261 8386 8325
rect 8450 8261 8466 8325
rect 8530 8261 8546 8325
rect 8610 8261 8626 8325
rect 8690 8261 8706 8325
rect 8770 8261 8786 8325
rect 8850 8261 8866 8325
rect 8930 8261 8946 8325
rect 9010 8261 9026 8325
rect 9090 8261 9106 8325
rect 9170 8261 9186 8325
rect 9250 8261 15000 8325
rect 0 8247 15000 8261
rect 0 8183 204 8247
rect 268 8183 287 8247
rect 351 8183 370 8247
rect 434 8183 453 8247
rect 517 8183 536 8247
rect 600 8183 618 8247
rect 682 8183 700 8247
rect 764 8183 782 8247
rect 846 8183 864 8247
rect 928 8183 946 8247
rect 1010 8183 1028 8247
rect 1092 8183 1110 8247
rect 1174 8183 1192 8247
rect 1256 8241 15000 8247
rect 1256 8183 8224 8241
rect 0 8177 8224 8183
rect 8288 8177 8305 8241
rect 8369 8177 8386 8241
rect 8450 8177 8466 8241
rect 8530 8177 8546 8241
rect 8610 8177 8626 8241
rect 8690 8177 8706 8241
rect 8770 8177 8786 8241
rect 8850 8177 8866 8241
rect 8930 8177 8946 8241
rect 9010 8177 9026 8241
rect 9090 8177 9106 8241
rect 9170 8177 9186 8241
rect 9250 8177 15000 8241
rect 0 8163 15000 8177
rect 0 8099 204 8163
rect 268 8099 287 8163
rect 351 8099 370 8163
rect 434 8099 453 8163
rect 517 8099 536 8163
rect 600 8099 618 8163
rect 682 8099 700 8163
rect 764 8099 782 8163
rect 846 8099 864 8163
rect 928 8099 946 8163
rect 1010 8099 1028 8163
rect 1092 8099 1110 8163
rect 1174 8099 1192 8163
rect 1256 8157 15000 8163
rect 1256 8099 8224 8157
rect 0 8093 8224 8099
rect 8288 8093 8305 8157
rect 8369 8093 8386 8157
rect 8450 8093 8466 8157
rect 8530 8093 8546 8157
rect 8610 8093 8626 8157
rect 8690 8093 8706 8157
rect 8770 8093 8786 8157
rect 8850 8093 8866 8157
rect 8930 8093 8946 8157
rect 9010 8093 9026 8157
rect 9090 8093 9106 8157
rect 9170 8093 9186 8157
rect 9250 8093 15000 8157
rect 0 8079 15000 8093
rect 0 8015 204 8079
rect 268 8015 287 8079
rect 351 8015 370 8079
rect 434 8015 453 8079
rect 517 8015 536 8079
rect 600 8015 618 8079
rect 682 8015 700 8079
rect 764 8015 782 8079
rect 846 8015 864 8079
rect 928 8015 946 8079
rect 1010 8015 1028 8079
rect 1092 8015 1110 8079
rect 1174 8015 1192 8079
rect 1256 8073 15000 8079
rect 1256 8015 8224 8073
rect 0 8009 8224 8015
rect 8288 8009 8305 8073
rect 8369 8009 8386 8073
rect 8450 8009 8466 8073
rect 8530 8009 8546 8073
rect 8610 8009 8626 8073
rect 8690 8009 8706 8073
rect 8770 8009 8786 8073
rect 8850 8009 8866 8073
rect 8930 8009 8946 8073
rect 9010 8009 9026 8073
rect 9090 8009 9106 8073
rect 9170 8009 9186 8073
rect 9250 8009 15000 8073
rect 0 7995 15000 8009
rect 0 7931 204 7995
rect 268 7931 287 7995
rect 351 7931 370 7995
rect 434 7931 453 7995
rect 517 7931 536 7995
rect 600 7931 618 7995
rect 682 7931 700 7995
rect 764 7931 782 7995
rect 846 7931 864 7995
rect 928 7931 946 7995
rect 1010 7931 1028 7995
rect 1092 7931 1110 7995
rect 1174 7931 1192 7995
rect 1256 7989 15000 7995
rect 1256 7931 8224 7989
rect 0 7925 8224 7931
rect 8288 7925 8305 7989
rect 8369 7925 8386 7989
rect 8450 7925 8466 7989
rect 8530 7925 8546 7989
rect 8610 7925 8626 7989
rect 8690 7925 8706 7989
rect 8770 7925 8786 7989
rect 8850 7925 8866 7989
rect 8930 7925 8946 7989
rect 9010 7925 9026 7989
rect 9090 7925 9106 7989
rect 9170 7925 9186 7989
rect 9250 7925 15000 7989
rect 0 7917 15000 7925
rect 0 6947 15000 7637
rect 0 5977 15000 6667
rect 0 4767 15000 5697
rect 0 3557 15000 4487
rect 0 2587 15000 3277
rect 0 1377 15000 2307
rect 0 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 6271 26615 8730 30317
rect 0 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_io__com_busses  sky130_fd_io__com_busses_0
timestamp 1701704242
transform 1 0 0 0 1 149
box 0 -142 15000 39451
use sky130_fd_io__top_analog_pad_pddrvr_strong  sky130_fd_io__top_analog_pad_pddrvr_strong_0
timestamp 1701704242
transform 1 0 0 0 -1 36357
box -80 307 15080 9520
use sky130_fd_io__top_analog_pad_pudrvr_strong  sky130_fd_io__top_analog_pad_pudrvr_strong_0
timestamp 1701704242
transform 1 0 -525 0 1 19219
box 493 -790 15554 5464
<< labels >>
flabel metal5 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 vssio
port 1 nsew ground bidirectional
flabel metal5 s 14746 4787 15000 5677 3 FreeSans 520 180 0 0 vssio
port 1 nsew ground bidirectional
flabel metal5 s 0 34757 254 39600 3 FreeSans 520 0 0 0 vssio
port 1 nsew ground bidirectional
flabel metal5 s 0 4787 254 5677 3 FreeSans 520 0 0 0 vssio
port 1 nsew ground bidirectional
flabel metal5 s 14746 1397 15000 2287 3 FreeSans 520 180 0 0 vccd
port 2 nsew power bidirectional
flabel metal5 s 0 1397 254 2287 3 FreeSans 520 0 0 0 vccd
port 2 nsew power bidirectional
flabel metal5 s 14746 12437 15000 13287 3 FreeSans 520 180 0 0 vddio_q
port 3 nsew power bidirectional
flabel metal5 s 0 12437 254 13287 3 FreeSans 520 0 0 0 vddio_q
port 3 nsew power bidirectional
flabel metal5 s 14746 9147 15000 10947 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 14746 6968 15000 7617 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 0 9147 254 10947 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 0 6968 254 7617 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 14746 13607 15000 18597 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 14746 3577 15000 4467 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 0 13607 254 18597 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 0 3577 254 4467 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 14746 27 15000 1077 3 FreeSans 520 180 0 0 vcchib
port 6 nsew power bidirectional
flabel metal5 s 0 27 254 1077 3 FreeSans 520 0 0 0 vcchib
port 6 nsew power bidirectional
flabel metal5 s 14746 5997 15000 6647 3 FreeSans 520 180 0 0 vswitch
port 7 nsew power bidirectional
flabel metal5 s 0 5997 254 6647 3 FreeSans 520 0 0 0 vswitch
port 7 nsew power bidirectional
flabel metal5 s 14746 11267 15000 12117 3 FreeSans 520 180 0 0 vssio_q
port 8 nsew ground bidirectional
flabel metal5 s 0 11267 254 12117 3 FreeSans 520 0 0 0 vssio_q
port 8 nsew ground bidirectional
flabel metal5 s 14807 2607 15000 3257 3 FreeSans 520 180 0 0 vdda
port 9 nsew power bidirectional
flabel metal5 s 0 2607 193 3257 3 FreeSans 520 0 0 0 vdda
port 9 nsew power bidirectional
flabel metal5 s 14746 7937 15000 8827 3 FreeSans 520 180 0 0 vssd
port 10 nsew ground bidirectional
flabel metal5 s 0 7937 254 8827 3 FreeSans 520 0 0 0 vssd
port 10 nsew ground bidirectional
flabel metal5 s 6271 26615 8730 30317 3 FreeSans 520 0 0 0 pad
port 11 nsew signal bidirectional
flabel metal5 s 14873 37921 14873 37921 3 FreeSans 520 180 0 0 vssio
flabel metal5 s 127 37921 127 37921 3 FreeSans 520 0 0 0 vssio
flabel metal5 s 127 37178 127 37178 0 FreeSans 512 0 0 0 vssio
flabel metal5 s 14873 37178 14873 37178 0 FreeSans 512 0 0 0 vssio
flabel metal4 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 vssio
port 1 nsew ground bidirectional
flabel metal4 s 14746 4767 15000 5697 3 FreeSans 520 180 0 0 vssio
port 1 nsew ground bidirectional
flabel metal4 s 0 34757 254 39600 3 FreeSans 520 0 0 0 vssio
port 1 nsew ground bidirectional
flabel metal4 s 0 4767 254 5697 3 FreeSans 520 0 0 0 vssio
port 1 nsew ground bidirectional
flabel metal4 s 14746 9273 15000 9869 3 FreeSans 520 180 0 0 amuxbus_b
port 12 nsew signal bidirectional
flabel metal4 s 0 9273 254 9869 3 FreeSans 520 0 0 0 amuxbus_b
port 12 nsew signal bidirectional
flabel metal4 s 14746 1377 15000 2307 3 FreeSans 520 180 0 0 vccd
port 2 nsew power bidirectional
flabel metal4 s 0 1377 254 2307 3 FreeSans 520 0 0 0 vccd
port 2 nsew power bidirectional
flabel metal4 s 14746 12417 15000 13307 3 FreeSans 520 180 0 0 vddio_q
port 3 nsew power bidirectional
flabel metal4 s 0 12417 254 13307 3 FreeSans 520 0 0 0 vddio_q
port 3 nsew power bidirectional
flabel metal4 s 14746 6947 15000 7637 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 14746 9147 15000 9213 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 14746 10881 15000 10947 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 14746 9929 15000 10165 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 0 9147 254 9213 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 0 9929 254 10165 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 0 10881 254 10947 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 0 6947 254 7637 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 14746 3557 15000 4487 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 14746 13607 15000 18600 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 0 3557 254 4487 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 0 13607 254 18600 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 14746 7 15000 1097 3 FreeSans 520 180 0 0 vcchib
port 6 nsew power bidirectional
flabel metal4 s 0 7 254 1097 3 FreeSans 520 0 0 0 vcchib
port 6 nsew power bidirectional
flabel metal4 s 14746 5977 15000 6667 3 FreeSans 520 180 0 0 vswitch
port 7 nsew power bidirectional
flabel metal4 s 0 5977 254 6667 3 FreeSans 520 0 0 0 vswitch
port 7 nsew power bidirectional
flabel metal4 s 14746 11247 15000 12137 3 FreeSans 520 180 0 0 vssio_q
port 8 nsew ground bidirectional
flabel metal4 s 0 11247 254 12137 3 FreeSans 520 0 0 0 vssio_q
port 8 nsew ground bidirectional
flabel metal4 s 14807 2587 15000 3277 3 FreeSans 520 180 0 0 vdda
port 9 nsew power bidirectional
flabel metal4 s 0 2587 193 3277 3 FreeSans 520 0 0 0 vdda
port 9 nsew power bidirectional
flabel metal4 s 14746 7917 15000 8847 3 FreeSans 520 180 0 0 vssd
port 10 nsew ground bidirectional
flabel metal4 s 0 7917 254 8847 3 FreeSans 520 0 0 0 vssd
port 10 nsew ground bidirectional
flabel metal4 s 14746 10225 15000 10821 3 FreeSans 520 180 0 0 amuxbus_a
port 13 nsew signal bidirectional
flabel metal4 s 0 10225 254 10821 3 FreeSans 520 0 0 0 amuxbus_a
port 13 nsew signal bidirectional
flabel metal4 s 14873 37921 14873 37921 3 FreeSans 520 180 0 0 vssio
flabel metal4 s 0 4767 15000 5697 3 FreeSans 520 0 0 0 vssio
port 15 nsew ground bidirectional
flabel metal4 s 0 34757 15000 39600 0 FreeSans 96 0 0 0 vssio
port 16 nsew ground bidirectional
flabel metal4 s 14873 37178 14873 37178 0 FreeSans 96 0 0 0 vssio
flabel metal3 s 7766 0 9562 977 0 FreeSans 96 0 0 0 pad_core
port 14 nsew signal bidirectional
rlabel metal4 s 0 1377 15000 2307 1 vccd
port 2 nsew power bidirectional
rlabel metal4 s 0 12417 15000 13307 1 vddio_q
port 3 nsew power bidirectional
rlabel metal5 s 0 9147 15000 10947 1 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 6947 15000 7637 1 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 1 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 9929 15000 10165 1 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 1 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 0 13607 15000 18597 1 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 3557 15000 4487 1 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 13607 15000 18600 1 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 7 15000 1097 1 vcchib
port 6 nsew power bidirectional
rlabel metal4 s 0 5977 15000 6667 1 vswitch
port 7 nsew power bidirectional
rlabel metal4 s 0 11247 15000 12137 1 vssio_q
port 8 nsew ground bidirectional
rlabel metal4 s 0 2587 15000 3277 1 vdda
port 9 nsew power bidirectional
rlabel metal4 s 0 7917 15000 8847 1 vssd
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string GDS_END 16732744
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 14492232
string LEFclass BLOCK
string LEFsymmetry R90
string path 64.400 340.325 64.400 464.825 
<< end >>
