magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 0 390 304 396
rect 0 0 304 6
<< via3 >>
rect 0 6 304 390
<< metal4 >>
rect -1 390 305 391
rect -1 6 0 390
rect 304 6 305 390
rect -1 5 305 6
<< properties >>
string GDS_END 94170942
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94169530
<< end >>
