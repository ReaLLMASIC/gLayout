magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal1 >>
rect 816 0 844 754
rect 1280 0 1308 754
rect 1440 0 1468 754
rect 1904 0 1932 754
rect 2064 0 2092 754
rect 2528 0 2556 754
rect 2688 0 2716 754
rect 3152 0 3180 754
rect 3312 0 3340 754
rect 3776 0 3804 754
rect 3936 0 3964 754
rect 4400 0 4428 754
rect 4560 0 4588 754
rect 5024 0 5052 754
rect 5184 0 5212 754
rect 5648 0 5676 754
rect 5808 0 5836 754
rect 6272 0 6300 754
rect 6432 0 6460 754
rect 6896 0 6924 754
rect 7056 0 7084 754
rect 7520 0 7548 754
rect 7680 0 7708 754
rect 8144 0 8172 754
rect 8304 0 8332 754
rect 8768 0 8796 754
rect 8928 0 8956 754
rect 9392 0 9420 754
rect 9552 0 9580 754
rect 10016 0 10044 754
rect 10176 0 10204 754
rect 10640 0 10668 754
rect 10800 0 10828 754
rect 11264 0 11292 754
rect 11424 0 11452 754
rect 11888 0 11916 754
rect 12048 0 12076 754
rect 12512 0 12540 754
rect 12672 0 12700 754
rect 13136 0 13164 754
rect 13296 0 13324 754
rect 13760 0 13788 754
rect 13920 0 13948 754
rect 14384 0 14412 754
rect 14544 0 14572 754
rect 15008 0 15036 754
rect 15168 0 15196 754
rect 15632 0 15660 754
rect 15792 0 15820 754
rect 16256 0 16284 754
rect 16416 0 16444 754
rect 16880 0 16908 754
rect 17040 0 17068 754
rect 17504 0 17532 754
rect 17664 0 17692 754
rect 18128 0 18156 754
rect 18288 0 18316 754
rect 18752 0 18780 754
rect 18912 0 18940 754
rect 19376 0 19404 754
rect 19536 0 19564 754
rect 20000 0 20028 754
rect 20160 0 20188 754
rect 20624 0 20652 754
rect 20784 0 20812 754
rect 21248 0 21276 754
rect 21408 0 21436 754
rect 21872 0 21900 754
rect 22032 0 22060 754
rect 22496 0 22524 754
rect 22656 0 22684 754
rect 23120 0 23148 754
rect 23280 0 23308 754
rect 23744 0 23772 754
rect 23904 0 23932 754
rect 24368 0 24396 754
rect 24528 0 24556 754
rect 24992 0 25020 754
rect 25152 0 25180 754
rect 25616 0 25644 754
rect 25776 0 25804 754
rect 26240 0 26268 754
rect 26400 0 26428 754
rect 26864 0 26892 754
rect 27024 0 27052 754
rect 27488 0 27516 754
rect 27648 0 27676 754
rect 28112 0 28140 754
rect 28272 0 28300 754
rect 28736 0 28764 754
rect 28896 0 28924 754
rect 29360 0 29388 754
rect 29520 0 29548 754
rect 29984 0 30012 754
rect 30144 0 30172 754
rect 30608 0 30636 754
rect 30768 0 30796 754
rect 31232 0 31260 754
rect 31392 0 31420 754
rect 31856 0 31884 754
rect 32016 0 32044 754
rect 32480 0 32508 754
rect 32640 0 32668 754
rect 33104 0 33132 754
rect 33264 0 33292 754
rect 33728 0 33756 754
rect 33888 0 33916 754
rect 34352 0 34380 754
rect 34512 0 34540 754
rect 34976 0 35004 754
rect 35136 0 35164 754
rect 35600 0 35628 754
rect 35760 0 35788 754
rect 36224 0 36252 754
rect 36384 0 36412 754
rect 36848 0 36876 754
rect 37008 0 37036 754
rect 37472 0 37500 754
rect 37632 0 37660 754
rect 38096 0 38124 754
rect 38256 0 38284 754
rect 38720 0 38748 754
rect 38880 0 38908 754
rect 39344 0 39372 754
rect 39504 0 39532 754
rect 39968 0 39996 754
rect 40128 0 40156 754
rect 40592 0 40620 754
rect 40752 0 40780 754
rect 41216 0 41244 754
rect 41376 0 41404 754
rect 41840 0 41868 754
rect 42000 0 42028 754
rect 42464 0 42492 754
rect 42624 0 42652 754
rect 43088 0 43116 754
rect 43248 0 43276 754
rect 43712 0 43740 754
rect 43872 0 43900 754
rect 44336 0 44364 754
rect 44496 0 44524 754
rect 44960 0 44988 754
rect 45120 0 45148 754
rect 45584 0 45612 754
rect 45744 0 45772 754
rect 46208 0 46236 754
rect 46368 0 46396 754
rect 46832 0 46860 754
rect 46992 0 47020 754
rect 47456 0 47484 754
rect 47616 0 47644 754
rect 48080 0 48108 754
rect 48240 0 48268 754
rect 48704 0 48732 754
rect 48864 0 48892 754
rect 49328 0 49356 754
rect 49488 0 49516 754
rect 49952 0 49980 754
rect 50112 0 50140 754
rect 50576 0 50604 754
rect 50736 0 50764 754
rect 51200 0 51228 754
rect 51360 0 51388 754
rect 51824 0 51852 754
rect 51984 0 52012 754
rect 52448 0 52476 754
rect 52608 0 52636 754
rect 53072 0 53100 754
rect 53232 0 53260 754
rect 53696 0 53724 754
rect 53856 0 53884 754
rect 54320 0 54348 754
rect 54480 0 54508 754
rect 54944 0 54972 754
rect 55104 0 55132 754
rect 55568 0 55596 754
rect 55728 0 55756 754
rect 56192 0 56220 754
rect 56352 0 56380 754
rect 56816 0 56844 754
rect 56976 0 57004 754
rect 57440 0 57468 754
rect 57600 0 57628 754
rect 58064 0 58092 754
rect 58224 0 58252 754
rect 58688 0 58716 754
rect 58848 0 58876 754
rect 59312 0 59340 754
rect 59472 0 59500 754
rect 59936 0 59964 754
rect 60096 0 60124 754
rect 60560 0 60588 754
rect 60720 0 60748 754
rect 61184 0 61212 754
rect 61344 0 61372 754
rect 61808 0 61836 754
rect 61968 0 61996 754
rect 62432 0 62460 754
rect 62592 0 62620 754
rect 63056 0 63084 754
rect 63216 0 63244 754
rect 63680 0 63708 754
rect 63840 0 63868 754
rect 64304 0 64332 754
rect 64464 0 64492 754
rect 64928 0 64956 754
rect 65088 0 65116 754
rect 65552 0 65580 754
rect 65712 0 65740 754
rect 66176 0 66204 754
rect 66336 0 66364 754
rect 66800 0 66828 754
rect 66960 0 66988 754
rect 67424 0 67452 754
rect 67584 0 67612 754
rect 68048 0 68076 754
rect 68208 0 68236 754
rect 68672 0 68700 754
rect 68832 0 68860 754
rect 69296 0 69324 754
rect 69456 0 69484 754
rect 69920 0 69948 754
rect 70080 0 70108 754
rect 70544 0 70572 754
rect 70704 0 70732 754
rect 71168 0 71196 754
rect 71328 0 71356 754
rect 71792 0 71820 754
rect 71952 0 71980 754
rect 72416 0 72444 754
rect 72576 0 72604 754
rect 73040 0 73068 754
rect 73200 0 73228 754
rect 73664 0 73692 754
rect 73824 0 73852 754
rect 74288 0 74316 754
rect 74448 0 74476 754
rect 74912 0 74940 754
rect 75072 0 75100 754
rect 75536 0 75564 754
rect 75696 0 75724 754
rect 76160 0 76188 754
rect 76320 0 76348 754
rect 76784 0 76812 754
rect 76944 0 76972 754
rect 77408 0 77436 754
rect 77568 0 77596 754
rect 78032 0 78060 754
rect 78192 0 78220 754
rect 78656 0 78684 754
rect 78816 0 78844 754
rect 79280 0 79308 754
rect 79440 0 79468 754
rect 79904 0 79932 754
rect 80064 0 80092 754
rect 80528 0 80556 754
rect 80688 0 80716 754
rect 81152 0 81180 754
<< metal2 >>
rect 1034 53 1090 62
rect 1034 -12 1090 -3
rect 1658 53 1714 62
rect 1658 -12 1714 -3
rect 2282 53 2338 62
rect 2282 -12 2338 -3
rect 2906 53 2962 62
rect 2906 -12 2962 -3
rect 3530 53 3586 62
rect 3530 -12 3586 -3
rect 4154 53 4210 62
rect 4154 -12 4210 -3
rect 4778 53 4834 62
rect 4778 -12 4834 -3
rect 5402 53 5458 62
rect 5402 -12 5458 -3
rect 6026 53 6082 62
rect 6026 -12 6082 -3
rect 6650 53 6706 62
rect 6650 -12 6706 -3
rect 7274 53 7330 62
rect 7274 -12 7330 -3
rect 7898 53 7954 62
rect 7898 -12 7954 -3
rect 8522 53 8578 62
rect 8522 -12 8578 -3
rect 9146 53 9202 62
rect 9146 -12 9202 -3
rect 9770 53 9826 62
rect 9770 -12 9826 -3
rect 10394 53 10450 62
rect 10394 -12 10450 -3
rect 11018 53 11074 62
rect 11018 -12 11074 -3
rect 11642 53 11698 62
rect 11642 -12 11698 -3
rect 12266 53 12322 62
rect 12266 -12 12322 -3
rect 12890 53 12946 62
rect 12890 -12 12946 -3
rect 13514 53 13570 62
rect 13514 -12 13570 -3
rect 14138 53 14194 62
rect 14138 -12 14194 -3
rect 14762 53 14818 62
rect 14762 -12 14818 -3
rect 15386 53 15442 62
rect 15386 -12 15442 -3
rect 16010 53 16066 62
rect 16010 -12 16066 -3
rect 16634 53 16690 62
rect 16634 -12 16690 -3
rect 17258 53 17314 62
rect 17258 -12 17314 -3
rect 17882 53 17938 62
rect 17882 -12 17938 -3
rect 18506 53 18562 62
rect 18506 -12 18562 -3
rect 19130 53 19186 62
rect 19130 -12 19186 -3
rect 19754 53 19810 62
rect 19754 -12 19810 -3
rect 20378 53 20434 62
rect 20378 -12 20434 -3
rect 21002 53 21058 62
rect 21002 -12 21058 -3
rect 21626 53 21682 62
rect 21626 -12 21682 -3
rect 22250 53 22306 62
rect 22250 -12 22306 -3
rect 22874 53 22930 62
rect 22874 -12 22930 -3
rect 23498 53 23554 62
rect 23498 -12 23554 -3
rect 24122 53 24178 62
rect 24122 -12 24178 -3
rect 24746 53 24802 62
rect 24746 -12 24802 -3
rect 25370 53 25426 62
rect 25370 -12 25426 -3
rect 25994 53 26050 62
rect 25994 -12 26050 -3
rect 26618 53 26674 62
rect 26618 -12 26674 -3
rect 27242 53 27298 62
rect 27242 -12 27298 -3
rect 27866 53 27922 62
rect 27866 -12 27922 -3
rect 28490 53 28546 62
rect 28490 -12 28546 -3
rect 29114 53 29170 62
rect 29114 -12 29170 -3
rect 29738 53 29794 62
rect 29738 -12 29794 -3
rect 30362 53 30418 62
rect 30362 -12 30418 -3
rect 30986 53 31042 62
rect 30986 -12 31042 -3
rect 31610 53 31666 62
rect 31610 -12 31666 -3
rect 32234 53 32290 62
rect 32234 -12 32290 -3
rect 32858 53 32914 62
rect 32858 -12 32914 -3
rect 33482 53 33538 62
rect 33482 -12 33538 -3
rect 34106 53 34162 62
rect 34106 -12 34162 -3
rect 34730 53 34786 62
rect 34730 -12 34786 -3
rect 35354 53 35410 62
rect 35354 -12 35410 -3
rect 35978 53 36034 62
rect 35978 -12 36034 -3
rect 36602 53 36658 62
rect 36602 -12 36658 -3
rect 37226 53 37282 62
rect 37226 -12 37282 -3
rect 37850 53 37906 62
rect 37850 -12 37906 -3
rect 38474 53 38530 62
rect 38474 -12 38530 -3
rect 39098 53 39154 62
rect 39098 -12 39154 -3
rect 39722 53 39778 62
rect 39722 -12 39778 -3
rect 40346 53 40402 62
rect 40346 -12 40402 -3
rect 40970 53 41026 62
rect 40970 -12 41026 -3
rect 41594 53 41650 62
rect 41594 -12 41650 -3
rect 42218 53 42274 62
rect 42218 -12 42274 -3
rect 42842 53 42898 62
rect 42842 -12 42898 -3
rect 43466 53 43522 62
rect 43466 -12 43522 -3
rect 44090 53 44146 62
rect 44090 -12 44146 -3
rect 44714 53 44770 62
rect 44714 -12 44770 -3
rect 45338 53 45394 62
rect 45338 -12 45394 -3
rect 45962 53 46018 62
rect 45962 -12 46018 -3
rect 46586 53 46642 62
rect 46586 -12 46642 -3
rect 47210 53 47266 62
rect 47210 -12 47266 -3
rect 47834 53 47890 62
rect 47834 -12 47890 -3
rect 48458 53 48514 62
rect 48458 -12 48514 -3
rect 49082 53 49138 62
rect 49082 -12 49138 -3
rect 49706 53 49762 62
rect 49706 -12 49762 -3
rect 50330 53 50386 62
rect 50330 -12 50386 -3
rect 50954 53 51010 62
rect 50954 -12 51010 -3
rect 51578 53 51634 62
rect 51578 -12 51634 -3
rect 52202 53 52258 62
rect 52202 -12 52258 -3
rect 52826 53 52882 62
rect 52826 -12 52882 -3
rect 53450 53 53506 62
rect 53450 -12 53506 -3
rect 54074 53 54130 62
rect 54074 -12 54130 -3
rect 54698 53 54754 62
rect 54698 -12 54754 -3
rect 55322 53 55378 62
rect 55322 -12 55378 -3
rect 55946 53 56002 62
rect 55946 -12 56002 -3
rect 56570 53 56626 62
rect 56570 -12 56626 -3
rect 57194 53 57250 62
rect 57194 -12 57250 -3
rect 57818 53 57874 62
rect 57818 -12 57874 -3
rect 58442 53 58498 62
rect 58442 -12 58498 -3
rect 59066 53 59122 62
rect 59066 -12 59122 -3
rect 59690 53 59746 62
rect 59690 -12 59746 -3
rect 60314 53 60370 62
rect 60314 -12 60370 -3
rect 60938 53 60994 62
rect 60938 -12 60994 -3
rect 61562 53 61618 62
rect 61562 -12 61618 -3
rect 62186 53 62242 62
rect 62186 -12 62242 -3
rect 62810 53 62866 62
rect 62810 -12 62866 -3
rect 63434 53 63490 62
rect 63434 -12 63490 -3
rect 64058 53 64114 62
rect 64058 -12 64114 -3
rect 64682 53 64738 62
rect 64682 -12 64738 -3
rect 65306 53 65362 62
rect 65306 -12 65362 -3
rect 65930 53 65986 62
rect 65930 -12 65986 -3
rect 66554 53 66610 62
rect 66554 -12 66610 -3
rect 67178 53 67234 62
rect 67178 -12 67234 -3
rect 67802 53 67858 62
rect 67802 -12 67858 -3
rect 68426 53 68482 62
rect 68426 -12 68482 -3
rect 69050 53 69106 62
rect 69050 -12 69106 -3
rect 69674 53 69730 62
rect 69674 -12 69730 -3
rect 70298 53 70354 62
rect 70298 -12 70354 -3
rect 70922 53 70978 62
rect 70922 -12 70978 -3
rect 71546 53 71602 62
rect 71546 -12 71602 -3
rect 72170 53 72226 62
rect 72170 -12 72226 -3
rect 72794 53 72850 62
rect 72794 -12 72850 -3
rect 73418 53 73474 62
rect 73418 -12 73474 -3
rect 74042 53 74098 62
rect 74042 -12 74098 -3
rect 74666 53 74722 62
rect 74666 -12 74722 -3
rect 75290 53 75346 62
rect 75290 -12 75346 -3
rect 75914 53 75970 62
rect 75914 -12 75970 -3
rect 76538 53 76594 62
rect 76538 -12 76594 -3
rect 77162 53 77218 62
rect 77162 -12 77218 -3
rect 77786 53 77842 62
rect 77786 -12 77842 -3
rect 78410 53 78466 62
rect 78410 -12 78466 -3
rect 79034 53 79090 62
rect 79034 -12 79090 -3
rect 79658 53 79714 62
rect 79658 -12 79714 -3
rect 80282 53 80338 62
rect 80282 -12 80338 -3
rect 80906 53 80962 62
rect 80906 -12 80962 -3
<< via2 >>
rect 1034 -3 1090 53
rect 1658 -3 1714 53
rect 2282 -3 2338 53
rect 2906 -3 2962 53
rect 3530 -3 3586 53
rect 4154 -3 4210 53
rect 4778 -3 4834 53
rect 5402 -3 5458 53
rect 6026 -3 6082 53
rect 6650 -3 6706 53
rect 7274 -3 7330 53
rect 7898 -3 7954 53
rect 8522 -3 8578 53
rect 9146 -3 9202 53
rect 9770 -3 9826 53
rect 10394 -3 10450 53
rect 11018 -3 11074 53
rect 11642 -3 11698 53
rect 12266 -3 12322 53
rect 12890 -3 12946 53
rect 13514 -3 13570 53
rect 14138 -3 14194 53
rect 14762 -3 14818 53
rect 15386 -3 15442 53
rect 16010 -3 16066 53
rect 16634 -3 16690 53
rect 17258 -3 17314 53
rect 17882 -3 17938 53
rect 18506 -3 18562 53
rect 19130 -3 19186 53
rect 19754 -3 19810 53
rect 20378 -3 20434 53
rect 21002 -3 21058 53
rect 21626 -3 21682 53
rect 22250 -3 22306 53
rect 22874 -3 22930 53
rect 23498 -3 23554 53
rect 24122 -3 24178 53
rect 24746 -3 24802 53
rect 25370 -3 25426 53
rect 25994 -3 26050 53
rect 26618 -3 26674 53
rect 27242 -3 27298 53
rect 27866 -3 27922 53
rect 28490 -3 28546 53
rect 29114 -3 29170 53
rect 29738 -3 29794 53
rect 30362 -3 30418 53
rect 30986 -3 31042 53
rect 31610 -3 31666 53
rect 32234 -3 32290 53
rect 32858 -3 32914 53
rect 33482 -3 33538 53
rect 34106 -3 34162 53
rect 34730 -3 34786 53
rect 35354 -3 35410 53
rect 35978 -3 36034 53
rect 36602 -3 36658 53
rect 37226 -3 37282 53
rect 37850 -3 37906 53
rect 38474 -3 38530 53
rect 39098 -3 39154 53
rect 39722 -3 39778 53
rect 40346 -3 40402 53
rect 40970 -3 41026 53
rect 41594 -3 41650 53
rect 42218 -3 42274 53
rect 42842 -3 42898 53
rect 43466 -3 43522 53
rect 44090 -3 44146 53
rect 44714 -3 44770 53
rect 45338 -3 45394 53
rect 45962 -3 46018 53
rect 46586 -3 46642 53
rect 47210 -3 47266 53
rect 47834 -3 47890 53
rect 48458 -3 48514 53
rect 49082 -3 49138 53
rect 49706 -3 49762 53
rect 50330 -3 50386 53
rect 50954 -3 51010 53
rect 51578 -3 51634 53
rect 52202 -3 52258 53
rect 52826 -3 52882 53
rect 53450 -3 53506 53
rect 54074 -3 54130 53
rect 54698 -3 54754 53
rect 55322 -3 55378 53
rect 55946 -3 56002 53
rect 56570 -3 56626 53
rect 57194 -3 57250 53
rect 57818 -3 57874 53
rect 58442 -3 58498 53
rect 59066 -3 59122 53
rect 59690 -3 59746 53
rect 60314 -3 60370 53
rect 60938 -3 60994 53
rect 61562 -3 61618 53
rect 62186 -3 62242 53
rect 62810 -3 62866 53
rect 63434 -3 63490 53
rect 64058 -3 64114 53
rect 64682 -3 64738 53
rect 65306 -3 65362 53
rect 65930 -3 65986 53
rect 66554 -3 66610 53
rect 67178 -3 67234 53
rect 67802 -3 67858 53
rect 68426 -3 68482 53
rect 69050 -3 69106 53
rect 69674 -3 69730 53
rect 70298 -3 70354 53
rect 70922 -3 70978 53
rect 71546 -3 71602 53
rect 72170 -3 72226 53
rect 72794 -3 72850 53
rect 73418 -3 73474 53
rect 74042 -3 74098 53
rect 74666 -3 74722 53
rect 75290 -3 75346 53
rect 75914 -3 75970 53
rect 76538 -3 76594 53
rect 77162 -3 77218 53
rect 77786 -3 77842 53
rect 78410 -3 78466 53
rect 79034 -3 79090 53
rect 79658 -3 79714 53
rect 80282 -3 80338 53
rect 80906 -3 80962 53
<< metal3 >>
rect 1132 595 1230 693
rect 1518 595 1616 693
rect 2380 595 2478 693
rect 2766 595 2864 693
rect 3628 595 3726 693
rect 4014 595 4112 693
rect 4876 595 4974 693
rect 5262 595 5360 693
rect 6124 595 6222 693
rect 6510 595 6608 693
rect 7372 595 7470 693
rect 7758 595 7856 693
rect 8620 595 8718 693
rect 9006 595 9104 693
rect 9868 595 9966 693
rect 10254 595 10352 693
rect 11116 595 11214 693
rect 11502 595 11600 693
rect 12364 595 12462 693
rect 12750 595 12848 693
rect 13612 595 13710 693
rect 13998 595 14096 693
rect 14860 595 14958 693
rect 15246 595 15344 693
rect 16108 595 16206 693
rect 16494 595 16592 693
rect 17356 595 17454 693
rect 17742 595 17840 693
rect 18604 595 18702 693
rect 18990 595 19088 693
rect 19852 595 19950 693
rect 20238 595 20336 693
rect 21100 595 21198 693
rect 21486 595 21584 693
rect 22348 595 22446 693
rect 22734 595 22832 693
rect 23596 595 23694 693
rect 23982 595 24080 693
rect 24844 595 24942 693
rect 25230 595 25328 693
rect 26092 595 26190 693
rect 26478 595 26576 693
rect 27340 595 27438 693
rect 27726 595 27824 693
rect 28588 595 28686 693
rect 28974 595 29072 693
rect 29836 595 29934 693
rect 30222 595 30320 693
rect 31084 595 31182 693
rect 31470 595 31568 693
rect 32332 595 32430 693
rect 32718 595 32816 693
rect 33580 595 33678 693
rect 33966 595 34064 693
rect 34828 595 34926 693
rect 35214 595 35312 693
rect 36076 595 36174 693
rect 36462 595 36560 693
rect 37324 595 37422 693
rect 37710 595 37808 693
rect 38572 595 38670 693
rect 38958 595 39056 693
rect 39820 595 39918 693
rect 40206 595 40304 693
rect 41068 595 41166 693
rect 41454 595 41552 693
rect 42316 595 42414 693
rect 42702 595 42800 693
rect 43564 595 43662 693
rect 43950 595 44048 693
rect 44812 595 44910 693
rect 45198 595 45296 693
rect 46060 595 46158 693
rect 46446 595 46544 693
rect 47308 595 47406 693
rect 47694 595 47792 693
rect 48556 595 48654 693
rect 48942 595 49040 693
rect 49804 595 49902 693
rect 50190 595 50288 693
rect 51052 595 51150 693
rect 51438 595 51536 693
rect 52300 595 52398 693
rect 52686 595 52784 693
rect 53548 595 53646 693
rect 53934 595 54032 693
rect 54796 595 54894 693
rect 55182 595 55280 693
rect 56044 595 56142 693
rect 56430 595 56528 693
rect 57292 595 57390 693
rect 57678 595 57776 693
rect 58540 595 58638 693
rect 58926 595 59024 693
rect 59788 595 59886 693
rect 60174 595 60272 693
rect 61036 595 61134 693
rect 61422 595 61520 693
rect 62284 595 62382 693
rect 62670 595 62768 693
rect 63532 595 63630 693
rect 63918 595 64016 693
rect 64780 595 64878 693
rect 65166 595 65264 693
rect 66028 595 66126 693
rect 66414 595 66512 693
rect 67276 595 67374 693
rect 67662 595 67760 693
rect 68524 595 68622 693
rect 68910 595 69008 693
rect 69772 595 69870 693
rect 70158 595 70256 693
rect 71020 595 71118 693
rect 71406 595 71504 693
rect 72268 595 72366 693
rect 72654 595 72752 693
rect 73516 595 73614 693
rect 73902 595 74000 693
rect 74764 595 74862 693
rect 75150 595 75248 693
rect 76012 595 76110 693
rect 76398 595 76496 693
rect 77260 595 77358 693
rect 77646 595 77744 693
rect 78508 595 78606 693
rect 78894 595 78992 693
rect 79756 595 79854 693
rect 80142 595 80240 693
rect 81004 595 81102 693
rect 1029 55 1095 58
rect 1653 55 1719 58
rect 2277 55 2343 58
rect 2901 55 2967 58
rect 3525 55 3591 58
rect 4149 55 4215 58
rect 4773 55 4839 58
rect 5397 55 5463 58
rect 6021 55 6087 58
rect 6645 55 6711 58
rect 7269 55 7335 58
rect 7893 55 7959 58
rect 8517 55 8583 58
rect 9141 55 9207 58
rect 9765 55 9831 58
rect 10389 55 10455 58
rect 11013 55 11079 58
rect 11637 55 11703 58
rect 12261 55 12327 58
rect 12885 55 12951 58
rect 13509 55 13575 58
rect 14133 55 14199 58
rect 14757 55 14823 58
rect 15381 55 15447 58
rect 16005 55 16071 58
rect 16629 55 16695 58
rect 17253 55 17319 58
rect 17877 55 17943 58
rect 18501 55 18567 58
rect 19125 55 19191 58
rect 19749 55 19815 58
rect 20373 55 20439 58
rect 20997 55 21063 58
rect 21621 55 21687 58
rect 22245 55 22311 58
rect 22869 55 22935 58
rect 23493 55 23559 58
rect 24117 55 24183 58
rect 24741 55 24807 58
rect 25365 55 25431 58
rect 25989 55 26055 58
rect 26613 55 26679 58
rect 27237 55 27303 58
rect 27861 55 27927 58
rect 28485 55 28551 58
rect 29109 55 29175 58
rect 29733 55 29799 58
rect 30357 55 30423 58
rect 30981 55 31047 58
rect 31605 55 31671 58
rect 32229 55 32295 58
rect 32853 55 32919 58
rect 33477 55 33543 58
rect 34101 55 34167 58
rect 34725 55 34791 58
rect 35349 55 35415 58
rect 35973 55 36039 58
rect 36597 55 36663 58
rect 37221 55 37287 58
rect 37845 55 37911 58
rect 38469 55 38535 58
rect 39093 55 39159 58
rect 39717 55 39783 58
rect 40341 55 40407 58
rect 40965 55 41031 58
rect 41589 55 41655 58
rect 42213 55 42279 58
rect 42837 55 42903 58
rect 43461 55 43527 58
rect 44085 55 44151 58
rect 44709 55 44775 58
rect 45333 55 45399 58
rect 45957 55 46023 58
rect 46581 55 46647 58
rect 47205 55 47271 58
rect 47829 55 47895 58
rect 48453 55 48519 58
rect 49077 55 49143 58
rect 49701 55 49767 58
rect 50325 55 50391 58
rect 50949 55 51015 58
rect 51573 55 51639 58
rect 52197 55 52263 58
rect 52821 55 52887 58
rect 53445 55 53511 58
rect 54069 55 54135 58
rect 54693 55 54759 58
rect 55317 55 55383 58
rect 55941 55 56007 58
rect 56565 55 56631 58
rect 57189 55 57255 58
rect 57813 55 57879 58
rect 58437 55 58503 58
rect 59061 55 59127 58
rect 59685 55 59751 58
rect 60309 55 60375 58
rect 60933 55 60999 58
rect 61557 55 61623 58
rect 62181 55 62247 58
rect 62805 55 62871 58
rect 63429 55 63495 58
rect 64053 55 64119 58
rect 64677 55 64743 58
rect 65301 55 65367 58
rect 65925 55 65991 58
rect 66549 55 66615 58
rect 67173 55 67239 58
rect 67797 55 67863 58
rect 68421 55 68487 58
rect 69045 55 69111 58
rect 69669 55 69735 58
rect 70293 55 70359 58
rect 70917 55 70983 58
rect 71541 55 71607 58
rect 72165 55 72231 58
rect 72789 55 72855 58
rect 73413 55 73479 58
rect 74037 55 74103 58
rect 74661 55 74727 58
rect 75285 55 75351 58
rect 75909 55 75975 58
rect 76533 55 76599 58
rect 77157 55 77223 58
rect 77781 55 77847 58
rect 78405 55 78471 58
rect 79029 55 79095 58
rect 79653 55 79719 58
rect 80277 55 80343 58
rect 80901 55 80967 58
rect 0 53 81246 55
rect 0 -3 1034 53
rect 1090 -3 1658 53
rect 1714 -3 2282 53
rect 2338 -3 2906 53
rect 2962 -3 3530 53
rect 3586 -3 4154 53
rect 4210 -3 4778 53
rect 4834 -3 5402 53
rect 5458 -3 6026 53
rect 6082 -3 6650 53
rect 6706 -3 7274 53
rect 7330 -3 7898 53
rect 7954 -3 8522 53
rect 8578 -3 9146 53
rect 9202 -3 9770 53
rect 9826 -3 10394 53
rect 10450 -3 11018 53
rect 11074 -3 11642 53
rect 11698 -3 12266 53
rect 12322 -3 12890 53
rect 12946 -3 13514 53
rect 13570 -3 14138 53
rect 14194 -3 14762 53
rect 14818 -3 15386 53
rect 15442 -3 16010 53
rect 16066 -3 16634 53
rect 16690 -3 17258 53
rect 17314 -3 17882 53
rect 17938 -3 18506 53
rect 18562 -3 19130 53
rect 19186 -3 19754 53
rect 19810 -3 20378 53
rect 20434 -3 21002 53
rect 21058 -3 21626 53
rect 21682 -3 22250 53
rect 22306 -3 22874 53
rect 22930 -3 23498 53
rect 23554 -3 24122 53
rect 24178 -3 24746 53
rect 24802 -3 25370 53
rect 25426 -3 25994 53
rect 26050 -3 26618 53
rect 26674 -3 27242 53
rect 27298 -3 27866 53
rect 27922 -3 28490 53
rect 28546 -3 29114 53
rect 29170 -3 29738 53
rect 29794 -3 30362 53
rect 30418 -3 30986 53
rect 31042 -3 31610 53
rect 31666 -3 32234 53
rect 32290 -3 32858 53
rect 32914 -3 33482 53
rect 33538 -3 34106 53
rect 34162 -3 34730 53
rect 34786 -3 35354 53
rect 35410 -3 35978 53
rect 36034 -3 36602 53
rect 36658 -3 37226 53
rect 37282 -3 37850 53
rect 37906 -3 38474 53
rect 38530 -3 39098 53
rect 39154 -3 39722 53
rect 39778 -3 40346 53
rect 40402 -3 40970 53
rect 41026 -3 41594 53
rect 41650 -3 42218 53
rect 42274 -3 42842 53
rect 42898 -3 43466 53
rect 43522 -3 44090 53
rect 44146 -3 44714 53
rect 44770 -3 45338 53
rect 45394 -3 45962 53
rect 46018 -3 46586 53
rect 46642 -3 47210 53
rect 47266 -3 47834 53
rect 47890 -3 48458 53
rect 48514 -3 49082 53
rect 49138 -3 49706 53
rect 49762 -3 50330 53
rect 50386 -3 50954 53
rect 51010 -3 51578 53
rect 51634 -3 52202 53
rect 52258 -3 52826 53
rect 52882 -3 53450 53
rect 53506 -3 54074 53
rect 54130 -3 54698 53
rect 54754 -3 55322 53
rect 55378 -3 55946 53
rect 56002 -3 56570 53
rect 56626 -3 57194 53
rect 57250 -3 57818 53
rect 57874 -3 58442 53
rect 58498 -3 59066 53
rect 59122 -3 59690 53
rect 59746 -3 60314 53
rect 60370 -3 60938 53
rect 60994 -3 61562 53
rect 61618 -3 62186 53
rect 62242 -3 62810 53
rect 62866 -3 63434 53
rect 63490 -3 64058 53
rect 64114 -3 64682 53
rect 64738 -3 65306 53
rect 65362 -3 65930 53
rect 65986 -3 66554 53
rect 66610 -3 67178 53
rect 67234 -3 67802 53
rect 67858 -3 68426 53
rect 68482 -3 69050 53
rect 69106 -3 69674 53
rect 69730 -3 70298 53
rect 70354 -3 70922 53
rect 70978 -3 71546 53
rect 71602 -3 72170 53
rect 72226 -3 72794 53
rect 72850 -3 73418 53
rect 73474 -3 74042 53
rect 74098 -3 74666 53
rect 74722 -3 75290 53
rect 75346 -3 75914 53
rect 75970 -3 76538 53
rect 76594 -3 77162 53
rect 77218 -3 77786 53
rect 77842 -3 78410 53
rect 78466 -3 79034 53
rect 79090 -3 79658 53
rect 79714 -3 80282 53
rect 80338 -3 80906 53
rect 80962 -3 81246 53
rect 0 -5 81246 -3
rect 1029 -8 1095 -5
rect 1653 -8 1719 -5
rect 2277 -8 2343 -5
rect 2901 -8 2967 -5
rect 3525 -8 3591 -5
rect 4149 -8 4215 -5
rect 4773 -8 4839 -5
rect 5397 -8 5463 -5
rect 6021 -8 6087 -5
rect 6645 -8 6711 -5
rect 7269 -8 7335 -5
rect 7893 -8 7959 -5
rect 8517 -8 8583 -5
rect 9141 -8 9207 -5
rect 9765 -8 9831 -5
rect 10389 -8 10455 -5
rect 11013 -8 11079 -5
rect 11637 -8 11703 -5
rect 12261 -8 12327 -5
rect 12885 -8 12951 -5
rect 13509 -8 13575 -5
rect 14133 -8 14199 -5
rect 14757 -8 14823 -5
rect 15381 -8 15447 -5
rect 16005 -8 16071 -5
rect 16629 -8 16695 -5
rect 17253 -8 17319 -5
rect 17877 -8 17943 -5
rect 18501 -8 18567 -5
rect 19125 -8 19191 -5
rect 19749 -8 19815 -5
rect 20373 -8 20439 -5
rect 20997 -8 21063 -5
rect 21621 -8 21687 -5
rect 22245 -8 22311 -5
rect 22869 -8 22935 -5
rect 23493 -8 23559 -5
rect 24117 -8 24183 -5
rect 24741 -8 24807 -5
rect 25365 -8 25431 -5
rect 25989 -8 26055 -5
rect 26613 -8 26679 -5
rect 27237 -8 27303 -5
rect 27861 -8 27927 -5
rect 28485 -8 28551 -5
rect 29109 -8 29175 -5
rect 29733 -8 29799 -5
rect 30357 -8 30423 -5
rect 30981 -8 31047 -5
rect 31605 -8 31671 -5
rect 32229 -8 32295 -5
rect 32853 -8 32919 -5
rect 33477 -8 33543 -5
rect 34101 -8 34167 -5
rect 34725 -8 34791 -5
rect 35349 -8 35415 -5
rect 35973 -8 36039 -5
rect 36597 -8 36663 -5
rect 37221 -8 37287 -5
rect 37845 -8 37911 -5
rect 38469 -8 38535 -5
rect 39093 -8 39159 -5
rect 39717 -8 39783 -5
rect 40341 -8 40407 -5
rect 40965 -8 41031 -5
rect 41589 -8 41655 -5
rect 42213 -8 42279 -5
rect 42837 -8 42903 -5
rect 43461 -8 43527 -5
rect 44085 -8 44151 -5
rect 44709 -8 44775 -5
rect 45333 -8 45399 -5
rect 45957 -8 46023 -5
rect 46581 -8 46647 -5
rect 47205 -8 47271 -5
rect 47829 -8 47895 -5
rect 48453 -8 48519 -5
rect 49077 -8 49143 -5
rect 49701 -8 49767 -5
rect 50325 -8 50391 -5
rect 50949 -8 51015 -5
rect 51573 -8 51639 -5
rect 52197 -8 52263 -5
rect 52821 -8 52887 -5
rect 53445 -8 53511 -5
rect 54069 -8 54135 -5
rect 54693 -8 54759 -5
rect 55317 -8 55383 -5
rect 55941 -8 56007 -5
rect 56565 -8 56631 -5
rect 57189 -8 57255 -5
rect 57813 -8 57879 -5
rect 58437 -8 58503 -5
rect 59061 -8 59127 -5
rect 59685 -8 59751 -5
rect 60309 -8 60375 -5
rect 60933 -8 60999 -5
rect 61557 -8 61623 -5
rect 62181 -8 62247 -5
rect 62805 -8 62871 -5
rect 63429 -8 63495 -5
rect 64053 -8 64119 -5
rect 64677 -8 64743 -5
rect 65301 -8 65367 -5
rect 65925 -8 65991 -5
rect 66549 -8 66615 -5
rect 67173 -8 67239 -5
rect 67797 -8 67863 -5
rect 68421 -8 68487 -5
rect 69045 -8 69111 -5
rect 69669 -8 69735 -5
rect 70293 -8 70359 -5
rect 70917 -8 70983 -5
rect 71541 -8 71607 -5
rect 72165 -8 72231 -5
rect 72789 -8 72855 -5
rect 73413 -8 73479 -5
rect 74037 -8 74103 -5
rect 74661 -8 74727 -5
rect 75285 -8 75351 -5
rect 75909 -8 75975 -5
rect 76533 -8 76599 -5
rect 77157 -8 77223 -5
rect 77781 -8 77847 -5
rect 78405 -8 78471 -5
rect 79029 -8 79095 -5
rect 79653 -8 79719 -5
rect 80277 -8 80343 -5
rect 80901 -8 80967 -5
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1701704242
transform 1 0 1029 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1701704242
transform 1 0 1653 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1701704242
transform 1 0 20373 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1701704242
transform 1 0 19749 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1701704242
transform 1 0 19125 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1701704242
transform 1 0 18501 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1701704242
transform 1 0 17877 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1701704242
transform 1 0 17253 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1701704242
transform 1 0 16629 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1701704242
transform 1 0 16005 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1701704242
transform 1 0 15381 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1701704242
transform 1 0 14757 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1701704242
transform 1 0 14133 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1701704242
transform 1 0 13509 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1701704242
transform 1 0 12885 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1701704242
transform 1 0 12261 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1701704242
transform 1 0 11637 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1701704242
transform 1 0 11013 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1701704242
transform 1 0 10389 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1701704242
transform 1 0 9765 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1701704242
transform 1 0 9141 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1701704242
transform 1 0 8517 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1701704242
transform 1 0 7893 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1701704242
transform 1 0 7269 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1701704242
transform 1 0 6645 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1701704242
transform 1 0 6021 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1701704242
transform 1 0 5397 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1701704242
transform 1 0 4773 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1701704242
transform 1 0 4149 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1701704242
transform 1 0 3525 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1701704242
transform 1 0 2901 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1701704242
transform 1 0 2277 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1701704242
transform 1 0 20997 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1701704242
transform 1 0 40341 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1701704242
transform 1 0 39717 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1701704242
transform 1 0 39093 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1701704242
transform 1 0 38469 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1701704242
transform 1 0 37845 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1701704242
transform 1 0 37221 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1701704242
transform 1 0 36597 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1701704242
transform 1 0 35973 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1701704242
transform 1 0 35349 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1701704242
transform 1 0 34725 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1701704242
transform 1 0 34101 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1701704242
transform 1 0 33477 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1701704242
transform 1 0 32853 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1701704242
transform 1 0 32229 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1701704242
transform 1 0 31605 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1701704242
transform 1 0 30981 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1701704242
transform 1 0 30357 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1701704242
transform 1 0 29733 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1701704242
transform 1 0 29109 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1701704242
transform 1 0 28485 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1701704242
transform 1 0 27861 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1701704242
transform 1 0 27237 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1701704242
transform 1 0 26613 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1701704242
transform 1 0 25989 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1701704242
transform 1 0 25365 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1701704242
transform 1 0 24741 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1701704242
transform 1 0 24117 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1701704242
transform 1 0 23493 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1701704242
transform 1 0 22869 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1701704242
transform 1 0 22245 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1701704242
transform 1 0 21621 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1701704242
transform 1 0 41589 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1701704242
transform 1 0 60933 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1701704242
transform 1 0 60309 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1701704242
transform 1 0 59685 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1701704242
transform 1 0 59061 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1701704242
transform 1 0 58437 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1701704242
transform 1 0 57813 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1701704242
transform 1 0 57189 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1701704242
transform 1 0 56565 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1701704242
transform 1 0 55941 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1701704242
transform 1 0 55317 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1701704242
transform 1 0 54693 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1701704242
transform 1 0 54069 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1701704242
transform 1 0 53445 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1701704242
transform 1 0 52821 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1701704242
transform 1 0 52197 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1701704242
transform 1 0 51573 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1701704242
transform 1 0 50949 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1701704242
transform 1 0 50325 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1701704242
transform 1 0 49701 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1701704242
transform 1 0 49077 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1701704242
transform 1 0 48453 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1701704242
transform 1 0 47829 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1701704242
transform 1 0 47205 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1701704242
transform 1 0 46581 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1701704242
transform 1 0 45957 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1701704242
transform 1 0 45333 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1701704242
transform 1 0 44709 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1701704242
transform 1 0 44085 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1701704242
transform 1 0 43461 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1701704242
transform 1 0 42837 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1701704242
transform 1 0 42213 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1701704242
transform 1 0 80901 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1701704242
transform 1 0 80277 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1701704242
transform 1 0 79653 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1701704242
transform 1 0 79029 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1701704242
transform 1 0 78405 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1701704242
transform 1 0 77781 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1701704242
transform 1 0 77157 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1701704242
transform 1 0 76533 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1701704242
transform 1 0 75909 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1701704242
transform 1 0 75285 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1701704242
transform 1 0 74661 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1701704242
transform 1 0 74037 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1701704242
transform 1 0 73413 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1701704242
transform 1 0 72789 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1701704242
transform 1 0 72165 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1701704242
transform 1 0 71541 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1701704242
transform 1 0 70917 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1701704242
transform 1 0 70293 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1701704242
transform 1 0 69669 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1701704242
transform 1 0 69045 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1701704242
transform 1 0 68421 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1701704242
transform 1 0 67797 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1701704242
transform 1 0 67173 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1701704242
transform 1 0 66549 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1701704242
transform 1 0 65925 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1701704242
transform 1 0 65301 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1701704242
transform 1 0 64677 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1701704242
transform 1 0 64053 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1701704242
transform 1 0 63429 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1701704242
transform 1 0 62805 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1701704242
transform 1 0 62181 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1701704242
transform 1 0 61557 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_128
timestamp 1701704242
transform 1 0 40965 0 1 -12
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_0
timestamp 1701704242
transform -1 0 1374 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_1
timestamp 1701704242
transform 1 0 1374 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_2
timestamp 1701704242
transform 1 0 20094 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_3
timestamp 1701704242
transform -1 0 20094 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_4
timestamp 1701704242
transform 1 0 18846 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_5
timestamp 1701704242
transform -1 0 18846 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_6
timestamp 1701704242
transform 1 0 17598 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_7
timestamp 1701704242
transform -1 0 17598 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_8
timestamp 1701704242
transform 1 0 16350 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_9
timestamp 1701704242
transform -1 0 16350 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_10
timestamp 1701704242
transform 1 0 15102 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_11
timestamp 1701704242
transform -1 0 15102 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_12
timestamp 1701704242
transform 1 0 13854 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_13
timestamp 1701704242
transform -1 0 13854 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_14
timestamp 1701704242
transform 1 0 12606 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_15
timestamp 1701704242
transform -1 0 12606 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_16
timestamp 1701704242
transform 1 0 11358 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_17
timestamp 1701704242
transform -1 0 11358 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_18
timestamp 1701704242
transform 1 0 10110 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_19
timestamp 1701704242
transform -1 0 10110 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_20
timestamp 1701704242
transform 1 0 8862 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_21
timestamp 1701704242
transform -1 0 8862 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_22
timestamp 1701704242
transform 1 0 7614 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_23
timestamp 1701704242
transform -1 0 7614 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_24
timestamp 1701704242
transform 1 0 6366 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_25
timestamp 1701704242
transform -1 0 6366 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_26
timestamp 1701704242
transform 1 0 5118 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_27
timestamp 1701704242
transform -1 0 5118 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_28
timestamp 1701704242
transform 1 0 3870 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_29
timestamp 1701704242
transform -1 0 3870 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_30
timestamp 1701704242
transform 1 0 2622 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_31
timestamp 1701704242
transform -1 0 2622 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_32
timestamp 1701704242
transform 1 0 40062 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_33
timestamp 1701704242
transform -1 0 40062 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_34
timestamp 1701704242
transform 1 0 38814 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_35
timestamp 1701704242
transform -1 0 38814 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_36
timestamp 1701704242
transform 1 0 37566 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_37
timestamp 1701704242
transform -1 0 37566 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_38
timestamp 1701704242
transform 1 0 36318 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_39
timestamp 1701704242
transform -1 0 36318 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_40
timestamp 1701704242
transform 1 0 35070 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_41
timestamp 1701704242
transform -1 0 35070 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_42
timestamp 1701704242
transform 1 0 33822 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_43
timestamp 1701704242
transform -1 0 33822 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_44
timestamp 1701704242
transform 1 0 32574 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_45
timestamp 1701704242
transform -1 0 32574 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_46
timestamp 1701704242
transform 1 0 31326 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_47
timestamp 1701704242
transform -1 0 31326 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_48
timestamp 1701704242
transform 1 0 30078 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_49
timestamp 1701704242
transform -1 0 30078 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_50
timestamp 1701704242
transform 1 0 28830 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_51
timestamp 1701704242
transform -1 0 28830 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_52
timestamp 1701704242
transform 1 0 27582 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_53
timestamp 1701704242
transform -1 0 27582 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_54
timestamp 1701704242
transform 1 0 26334 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_55
timestamp 1701704242
transform -1 0 26334 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_56
timestamp 1701704242
transform 1 0 25086 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_57
timestamp 1701704242
transform -1 0 25086 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_58
timestamp 1701704242
transform 1 0 23838 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_59
timestamp 1701704242
transform -1 0 23838 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_60
timestamp 1701704242
transform 1 0 22590 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_61
timestamp 1701704242
transform -1 0 22590 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_62
timestamp 1701704242
transform 1 0 21342 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_63
timestamp 1701704242
transform -1 0 21342 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_64
timestamp 1701704242
transform 1 0 41310 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_65
timestamp 1701704242
transform -1 0 43806 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_66
timestamp 1701704242
transform 1 0 42558 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_67
timestamp 1701704242
transform -1 0 42558 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_68
timestamp 1701704242
transform 1 0 60030 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_69
timestamp 1701704242
transform -1 0 60030 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_70
timestamp 1701704242
transform 1 0 58782 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_71
timestamp 1701704242
transform -1 0 58782 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_72
timestamp 1701704242
transform 1 0 57534 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_73
timestamp 1701704242
transform -1 0 57534 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_74
timestamp 1701704242
transform 1 0 56286 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_75
timestamp 1701704242
transform -1 0 56286 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_76
timestamp 1701704242
transform 1 0 55038 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_77
timestamp 1701704242
transform -1 0 55038 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_78
timestamp 1701704242
transform 1 0 53790 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_79
timestamp 1701704242
transform -1 0 53790 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_80
timestamp 1701704242
transform 1 0 52542 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_81
timestamp 1701704242
transform -1 0 52542 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_82
timestamp 1701704242
transform 1 0 51294 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_83
timestamp 1701704242
transform -1 0 51294 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_84
timestamp 1701704242
transform 1 0 50046 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_85
timestamp 1701704242
transform -1 0 50046 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_86
timestamp 1701704242
transform 1 0 48798 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_87
timestamp 1701704242
transform -1 0 48798 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_88
timestamp 1701704242
transform 1 0 47550 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_89
timestamp 1701704242
transform -1 0 47550 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_90
timestamp 1701704242
transform 1 0 46302 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_91
timestamp 1701704242
transform -1 0 46302 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_92
timestamp 1701704242
transform 1 0 45054 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_93
timestamp 1701704242
transform -1 0 45054 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_94
timestamp 1701704242
transform 1 0 43806 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_95
timestamp 1701704242
transform -1 0 81246 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_96
timestamp 1701704242
transform 1 0 79998 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_97
timestamp 1701704242
transform -1 0 79998 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_98
timestamp 1701704242
transform 1 0 78750 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_99
timestamp 1701704242
transform -1 0 78750 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_100
timestamp 1701704242
transform 1 0 77502 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_101
timestamp 1701704242
transform -1 0 77502 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_102
timestamp 1701704242
transform 1 0 76254 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_103
timestamp 1701704242
transform -1 0 76254 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_104
timestamp 1701704242
transform 1 0 75006 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_105
timestamp 1701704242
transform -1 0 75006 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_106
timestamp 1701704242
transform 1 0 73758 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_107
timestamp 1701704242
transform -1 0 73758 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_108
timestamp 1701704242
transform 1 0 72510 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_109
timestamp 1701704242
transform -1 0 72510 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_110
timestamp 1701704242
transform 1 0 71262 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_111
timestamp 1701704242
transform -1 0 71262 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_112
timestamp 1701704242
transform 1 0 70014 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_113
timestamp 1701704242
transform -1 0 70014 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_114
timestamp 1701704242
transform 1 0 68766 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_115
timestamp 1701704242
transform -1 0 68766 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_116
timestamp 1701704242
transform 1 0 67518 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_117
timestamp 1701704242
transform -1 0 67518 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_118
timestamp 1701704242
transform 1 0 66270 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_119
timestamp 1701704242
transform -1 0 66270 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_120
timestamp 1701704242
transform 1 0 65022 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_121
timestamp 1701704242
transform -1 0 65022 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_122
timestamp 1701704242
transform 1 0 63774 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_123
timestamp 1701704242
transform -1 0 63774 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_124
timestamp 1701704242
transform 1 0 62526 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_125
timestamp 1701704242
transform -1 0 62526 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_126
timestamp 1701704242
transform 1 0 61278 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_127
timestamp 1701704242
transform -1 0 61278 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_128
timestamp 1701704242
transform -1 0 41310 0 1 0
box 0 -8 624 768
<< labels >>
rlabel metal3 s 48556 595 48654 693 4 vdd
port 1 nsew
rlabel metal3 s 66028 595 66126 693 4 vdd
port 1 nsew
rlabel metal3 s 81004 595 81102 693 4 vdd
port 1 nsew
rlabel metal3 s 45198 595 45296 693 4 vdd
port 1 nsew
rlabel metal3 s 46060 595 46158 693 4 vdd
port 1 nsew
rlabel metal3 s 71020 595 71118 693 4 vdd
port 1 nsew
rlabel metal3 s 43564 595 43662 693 4 vdd
port 1 nsew
rlabel metal3 s 62670 595 62768 693 4 vdd
port 1 nsew
rlabel metal3 s 66414 595 66512 693 4 vdd
port 1 nsew
rlabel metal3 s 55182 595 55280 693 4 vdd
port 1 nsew
rlabel metal3 s 75150 595 75248 693 4 vdd
port 1 nsew
rlabel metal3 s 48942 595 49040 693 4 vdd
port 1 nsew
rlabel metal3 s 63918 595 64016 693 4 vdd
port 1 nsew
rlabel metal3 s 69772 595 69870 693 4 vdd
port 1 nsew
rlabel metal3 s 78508 595 78606 693 4 vdd
port 1 nsew
rlabel metal3 s 65166 595 65264 693 4 vdd
port 1 nsew
rlabel metal3 s 68910 595 69008 693 4 vdd
port 1 nsew
rlabel metal3 s 46446 595 46544 693 4 vdd
port 1 nsew
rlabel metal3 s 52300 595 52398 693 4 vdd
port 1 nsew
rlabel metal3 s 63532 595 63630 693 4 vdd
port 1 nsew
rlabel metal3 s 49804 595 49902 693 4 vdd
port 1 nsew
rlabel metal3 s 44812 595 44910 693 4 vdd
port 1 nsew
rlabel metal3 s 64780 595 64878 693 4 vdd
port 1 nsew
rlabel metal3 s 77260 595 77358 693 4 vdd
port 1 nsew
rlabel metal3 s 67662 595 67760 693 4 vdd
port 1 nsew
rlabel metal3 s 68524 595 68622 693 4 vdd
port 1 nsew
rlabel metal3 s 42702 595 42800 693 4 vdd
port 1 nsew
rlabel metal3 s 56430 595 56528 693 4 vdd
port 1 nsew
rlabel metal3 s 76398 595 76496 693 4 vdd
port 1 nsew
rlabel metal3 s 71406 595 71504 693 4 vdd
port 1 nsew
rlabel metal3 s 53934 595 54032 693 4 vdd
port 1 nsew
rlabel metal3 s 42316 595 42414 693 4 vdd
port 1 nsew
rlabel metal3 s 77646 595 77744 693 4 vdd
port 1 nsew
rlabel metal3 s 58540 595 58638 693 4 vdd
port 1 nsew
rlabel metal3 s 61422 595 61520 693 4 vdd
port 1 nsew
rlabel metal3 s 54796 595 54894 693 4 vdd
port 1 nsew
rlabel metal3 s 53548 595 53646 693 4 vdd
port 1 nsew
rlabel metal3 s 80142 595 80240 693 4 vdd
port 1 nsew
rlabel metal3 s 41454 595 41552 693 4 vdd
port 1 nsew
rlabel metal3 s 70158 595 70256 693 4 vdd
port 1 nsew
rlabel metal3 s 60174 595 60272 693 4 vdd
port 1 nsew
rlabel metal3 s 57678 595 57776 693 4 vdd
port 1 nsew
rlabel metal3 s 61036 595 61134 693 4 vdd
port 1 nsew
rlabel metal3 s 74764 595 74862 693 4 vdd
port 1 nsew
rlabel metal3 s 73516 595 73614 693 4 vdd
port 1 nsew
rlabel metal3 s 47308 595 47406 693 4 vdd
port 1 nsew
rlabel metal3 s 50190 595 50288 693 4 vdd
port 1 nsew
rlabel metal3 s 51052 595 51150 693 4 vdd
port 1 nsew
rlabel metal3 s 73902 595 74000 693 4 vdd
port 1 nsew
rlabel metal3 s 72654 595 72752 693 4 vdd
port 1 nsew
rlabel metal3 s 43950 595 44048 693 4 vdd
port 1 nsew
rlabel metal3 s 78894 595 78992 693 4 vdd
port 1 nsew
rlabel metal3 s 47694 595 47792 693 4 vdd
port 1 nsew
rlabel metal3 s 57292 595 57390 693 4 vdd
port 1 nsew
rlabel metal3 s 67276 595 67374 693 4 vdd
port 1 nsew
rlabel metal3 s 52686 595 52784 693 4 vdd
port 1 nsew
rlabel metal3 s 58926 595 59024 693 4 vdd
port 1 nsew
rlabel metal3 s 79756 595 79854 693 4 vdd
port 1 nsew
rlabel metal3 s 51438 595 51536 693 4 vdd
port 1 nsew
rlabel metal3 s 62284 595 62382 693 4 vdd
port 1 nsew
rlabel metal3 s 56044 595 56142 693 4 vdd
port 1 nsew
rlabel metal3 s 59788 595 59886 693 4 vdd
port 1 nsew
rlabel metal3 s 72268 595 72366 693 4 vdd
port 1 nsew
rlabel metal3 s 76012 595 76110 693 4 vdd
port 1 nsew
rlabel metal3 s 23596 595 23694 693 4 vdd
port 1 nsew
rlabel metal3 s 23982 595 24080 693 4 vdd
port 1 nsew
rlabel metal3 s 1132 595 1230 693 4 vdd
port 1 nsew
rlabel metal3 s 28974 595 29072 693 4 vdd
port 1 nsew
rlabel metal3 s 31470 595 31568 693 4 vdd
port 1 nsew
rlabel metal3 s 38572 595 38670 693 4 vdd
port 1 nsew
rlabel metal3 s 16494 595 16592 693 4 vdd
port 1 nsew
rlabel metal3 s 2380 595 2478 693 4 vdd
port 1 nsew
rlabel metal3 s 9006 595 9104 693 4 vdd
port 1 nsew
rlabel metal3 s 21486 595 21584 693 4 vdd
port 1 nsew
rlabel metal3 s 38958 595 39056 693 4 vdd
port 1 nsew
rlabel metal3 s 12750 595 12848 693 4 vdd
port 1 nsew
rlabel metal3 s 17742 595 17840 693 4 vdd
port 1 nsew
rlabel metal3 s 26478 595 26576 693 4 vdd
port 1 nsew
rlabel metal3 s 21100 595 21198 693 4 vdd
port 1 nsew
rlabel metal3 s 27726 595 27824 693 4 vdd
port 1 nsew
rlabel metal3 s 19852 595 19950 693 4 vdd
port 1 nsew
rlabel metal3 s 26092 595 26190 693 4 vdd
port 1 nsew
rlabel metal3 s 2766 595 2864 693 4 vdd
port 1 nsew
rlabel metal3 s 33580 595 33678 693 4 vdd
port 1 nsew
rlabel metal3 s 10254 595 10352 693 4 vdd
port 1 nsew
rlabel metal3 s 4014 595 4112 693 4 vdd
port 1 nsew
rlabel metal3 s 6124 595 6222 693 4 vdd
port 1 nsew
rlabel metal3 s 17356 595 17454 693 4 vdd
port 1 nsew
rlabel metal3 s 18604 595 18702 693 4 vdd
port 1 nsew
rlabel metal3 s 12364 595 12462 693 4 vdd
port 1 nsew
rlabel metal3 s 36462 595 36560 693 4 vdd
port 1 nsew
rlabel metal3 s 13612 595 13710 693 4 vdd
port 1 nsew
rlabel metal3 s 15246 595 15344 693 4 vdd
port 1 nsew
rlabel metal3 s 28588 595 28686 693 4 vdd
port 1 nsew
rlabel metal3 s 27340 595 27438 693 4 vdd
port 1 nsew
rlabel metal3 s 35214 595 35312 693 4 vdd
port 1 nsew
rlabel metal3 s 9868 595 9966 693 4 vdd
port 1 nsew
rlabel metal3 s 14860 595 14958 693 4 vdd
port 1 nsew
rlabel metal3 s 39820 595 39918 693 4 vdd
port 1 nsew
rlabel metal3 s 5262 595 5360 693 4 vdd
port 1 nsew
rlabel metal3 s 7372 595 7470 693 4 vdd
port 1 nsew
rlabel metal3 s 11502 595 11600 693 4 vdd
port 1 nsew
rlabel metal3 s 18990 595 19088 693 4 vdd
port 1 nsew
rlabel metal3 s 34828 595 34926 693 4 vdd
port 1 nsew
rlabel metal3 s 8620 595 8718 693 4 vdd
port 1 nsew
rlabel metal3 s 7758 595 7856 693 4 vdd
port 1 nsew
rlabel metal3 s 11116 595 11214 693 4 vdd
port 1 nsew
rlabel metal3 s 22348 595 22446 693 4 vdd
port 1 nsew
rlabel metal3 s 22734 595 22832 693 4 vdd
port 1 nsew
rlabel metal3 s 32718 595 32816 693 4 vdd
port 1 nsew
rlabel metal3 s 25230 595 25328 693 4 vdd
port 1 nsew
rlabel metal3 s 40206 595 40304 693 4 vdd
port 1 nsew
rlabel metal3 s 37324 595 37422 693 4 vdd
port 1 nsew
rlabel metal3 s 41068 595 41166 693 4 vdd
port 1 nsew
rlabel metal3 s 32332 595 32430 693 4 vdd
port 1 nsew
rlabel metal3 s 36076 595 36174 693 4 vdd
port 1 nsew
rlabel metal3 s 4876 595 4974 693 4 vdd
port 1 nsew
rlabel metal3 s 16108 595 16206 693 4 vdd
port 1 nsew
rlabel metal3 s 24844 595 24942 693 4 vdd
port 1 nsew
rlabel metal3 s 37710 595 37808 693 4 vdd
port 1 nsew
rlabel metal3 s 6510 595 6608 693 4 vdd
port 1 nsew
rlabel metal3 s 13998 595 14096 693 4 vdd
port 1 nsew
rlabel metal3 s 1518 595 1616 693 4 vdd
port 1 nsew
rlabel metal3 s 3628 595 3726 693 4 vdd
port 1 nsew
rlabel metal3 s 30222 595 30320 693 4 vdd
port 1 nsew
rlabel metal3 s 29836 595 29934 693 4 vdd
port 1 nsew
rlabel metal3 s 31084 595 31182 693 4 vdd
port 1 nsew
rlabel metal3 s 20238 595 20336 693 4 vdd
port 1 nsew
rlabel metal3 s 33966 595 34064 693 4 vdd
port 1 nsew
rlabel metal3 s 0 -5 81246 55 4 en_bar
port 2 nsew
rlabel metal1 s 1280 0 1308 754 4 bl_0
port 3 nsew
rlabel metal1 s 816 0 844 754 4 br_0
port 4 nsew
rlabel metal1 s 1440 0 1468 754 4 bl_1
port 5 nsew
rlabel metal1 s 1904 0 1932 754 4 br_1
port 6 nsew
rlabel metal1 s 2528 0 2556 754 4 bl_2
port 7 nsew
rlabel metal1 s 2064 0 2092 754 4 br_2
port 8 nsew
rlabel metal1 s 2688 0 2716 754 4 bl_3
port 9 nsew
rlabel metal1 s 3152 0 3180 754 4 br_3
port 10 nsew
rlabel metal1 s 3776 0 3804 754 4 bl_4
port 11 nsew
rlabel metal1 s 3312 0 3340 754 4 br_4
port 12 nsew
rlabel metal1 s 3936 0 3964 754 4 bl_5
port 13 nsew
rlabel metal1 s 4400 0 4428 754 4 br_5
port 14 nsew
rlabel metal1 s 5024 0 5052 754 4 bl_6
port 15 nsew
rlabel metal1 s 4560 0 4588 754 4 br_6
port 16 nsew
rlabel metal1 s 5184 0 5212 754 4 bl_7
port 17 nsew
rlabel metal1 s 5648 0 5676 754 4 br_7
port 18 nsew
rlabel metal1 s 6272 0 6300 754 4 bl_8
port 19 nsew
rlabel metal1 s 5808 0 5836 754 4 br_8
port 20 nsew
rlabel metal1 s 6432 0 6460 754 4 bl_9
port 21 nsew
rlabel metal1 s 6896 0 6924 754 4 br_9
port 22 nsew
rlabel metal1 s 7520 0 7548 754 4 bl_10
port 23 nsew
rlabel metal1 s 7056 0 7084 754 4 br_10
port 24 nsew
rlabel metal1 s 7680 0 7708 754 4 bl_11
port 25 nsew
rlabel metal1 s 8144 0 8172 754 4 br_11
port 26 nsew
rlabel metal1 s 8768 0 8796 754 4 bl_12
port 27 nsew
rlabel metal1 s 8304 0 8332 754 4 br_12
port 28 nsew
rlabel metal1 s 8928 0 8956 754 4 bl_13
port 29 nsew
rlabel metal1 s 9392 0 9420 754 4 br_13
port 30 nsew
rlabel metal1 s 10016 0 10044 754 4 bl_14
port 31 nsew
rlabel metal1 s 9552 0 9580 754 4 br_14
port 32 nsew
rlabel metal1 s 10176 0 10204 754 4 bl_15
port 33 nsew
rlabel metal1 s 10640 0 10668 754 4 br_15
port 34 nsew
rlabel metal1 s 11264 0 11292 754 4 bl_16
port 35 nsew
rlabel metal1 s 10800 0 10828 754 4 br_16
port 36 nsew
rlabel metal1 s 11424 0 11452 754 4 bl_17
port 37 nsew
rlabel metal1 s 11888 0 11916 754 4 br_17
port 38 nsew
rlabel metal1 s 12512 0 12540 754 4 bl_18
port 39 nsew
rlabel metal1 s 12048 0 12076 754 4 br_18
port 40 nsew
rlabel metal1 s 12672 0 12700 754 4 bl_19
port 41 nsew
rlabel metal1 s 13136 0 13164 754 4 br_19
port 42 nsew
rlabel metal1 s 13760 0 13788 754 4 bl_20
port 43 nsew
rlabel metal1 s 13296 0 13324 754 4 br_20
port 44 nsew
rlabel metal1 s 13920 0 13948 754 4 bl_21
port 45 nsew
rlabel metal1 s 14384 0 14412 754 4 br_21
port 46 nsew
rlabel metal1 s 15008 0 15036 754 4 bl_22
port 47 nsew
rlabel metal1 s 14544 0 14572 754 4 br_22
port 48 nsew
rlabel metal1 s 15168 0 15196 754 4 bl_23
port 49 nsew
rlabel metal1 s 15632 0 15660 754 4 br_23
port 50 nsew
rlabel metal1 s 16256 0 16284 754 4 bl_24
port 51 nsew
rlabel metal1 s 15792 0 15820 754 4 br_24
port 52 nsew
rlabel metal1 s 16416 0 16444 754 4 bl_25
port 53 nsew
rlabel metal1 s 16880 0 16908 754 4 br_25
port 54 nsew
rlabel metal1 s 17504 0 17532 754 4 bl_26
port 55 nsew
rlabel metal1 s 17040 0 17068 754 4 br_26
port 56 nsew
rlabel metal1 s 17664 0 17692 754 4 bl_27
port 57 nsew
rlabel metal1 s 18128 0 18156 754 4 br_27
port 58 nsew
rlabel metal1 s 18752 0 18780 754 4 bl_28
port 59 nsew
rlabel metal1 s 18288 0 18316 754 4 br_28
port 60 nsew
rlabel metal1 s 18912 0 18940 754 4 bl_29
port 61 nsew
rlabel metal1 s 19376 0 19404 754 4 br_29
port 62 nsew
rlabel metal1 s 20000 0 20028 754 4 bl_30
port 63 nsew
rlabel metal1 s 19536 0 19564 754 4 br_30
port 64 nsew
rlabel metal1 s 20160 0 20188 754 4 bl_31
port 65 nsew
rlabel metal1 s 20624 0 20652 754 4 br_31
port 66 nsew
rlabel metal1 s 20784 0 20812 754 4 br_32
port 67 nsew
rlabel metal1 s 21248 0 21276 754 4 bl_32
port 68 nsew
rlabel metal1 s 21408 0 21436 754 4 bl_33
port 69 nsew
rlabel metal1 s 21872 0 21900 754 4 br_33
port 70 nsew
rlabel metal1 s 22496 0 22524 754 4 bl_34
port 71 nsew
rlabel metal1 s 22032 0 22060 754 4 br_34
port 72 nsew
rlabel metal1 s 22656 0 22684 754 4 bl_35
port 73 nsew
rlabel metal1 s 23120 0 23148 754 4 br_35
port 74 nsew
rlabel metal1 s 23744 0 23772 754 4 bl_36
port 75 nsew
rlabel metal1 s 23280 0 23308 754 4 br_36
port 76 nsew
rlabel metal1 s 23904 0 23932 754 4 bl_37
port 77 nsew
rlabel metal1 s 24368 0 24396 754 4 br_37
port 78 nsew
rlabel metal1 s 24992 0 25020 754 4 bl_38
port 79 nsew
rlabel metal1 s 24528 0 24556 754 4 br_38
port 80 nsew
rlabel metal1 s 25152 0 25180 754 4 bl_39
port 81 nsew
rlabel metal1 s 25616 0 25644 754 4 br_39
port 82 nsew
rlabel metal1 s 26240 0 26268 754 4 bl_40
port 83 nsew
rlabel metal1 s 25776 0 25804 754 4 br_40
port 84 nsew
rlabel metal1 s 26400 0 26428 754 4 bl_41
port 85 nsew
rlabel metal1 s 26864 0 26892 754 4 br_41
port 86 nsew
rlabel metal1 s 27488 0 27516 754 4 bl_42
port 87 nsew
rlabel metal1 s 27024 0 27052 754 4 br_42
port 88 nsew
rlabel metal1 s 27648 0 27676 754 4 bl_43
port 89 nsew
rlabel metal1 s 28112 0 28140 754 4 br_43
port 90 nsew
rlabel metal1 s 28736 0 28764 754 4 bl_44
port 91 nsew
rlabel metal1 s 28272 0 28300 754 4 br_44
port 92 nsew
rlabel metal1 s 28896 0 28924 754 4 bl_45
port 93 nsew
rlabel metal1 s 29360 0 29388 754 4 br_45
port 94 nsew
rlabel metal1 s 29984 0 30012 754 4 bl_46
port 95 nsew
rlabel metal1 s 29520 0 29548 754 4 br_46
port 96 nsew
rlabel metal1 s 30144 0 30172 754 4 bl_47
port 97 nsew
rlabel metal1 s 30608 0 30636 754 4 br_47
port 98 nsew
rlabel metal1 s 31232 0 31260 754 4 bl_48
port 99 nsew
rlabel metal1 s 30768 0 30796 754 4 br_48
port 100 nsew
rlabel metal1 s 31392 0 31420 754 4 bl_49
port 101 nsew
rlabel metal1 s 31856 0 31884 754 4 br_49
port 102 nsew
rlabel metal1 s 32480 0 32508 754 4 bl_50
port 103 nsew
rlabel metal1 s 32016 0 32044 754 4 br_50
port 104 nsew
rlabel metal1 s 32640 0 32668 754 4 bl_51
port 105 nsew
rlabel metal1 s 33104 0 33132 754 4 br_51
port 106 nsew
rlabel metal1 s 33728 0 33756 754 4 bl_52
port 107 nsew
rlabel metal1 s 33264 0 33292 754 4 br_52
port 108 nsew
rlabel metal1 s 33888 0 33916 754 4 bl_53
port 109 nsew
rlabel metal1 s 34352 0 34380 754 4 br_53
port 110 nsew
rlabel metal1 s 34976 0 35004 754 4 bl_54
port 111 nsew
rlabel metal1 s 34512 0 34540 754 4 br_54
port 112 nsew
rlabel metal1 s 35136 0 35164 754 4 bl_55
port 113 nsew
rlabel metal1 s 35600 0 35628 754 4 br_55
port 114 nsew
rlabel metal1 s 36224 0 36252 754 4 bl_56
port 115 nsew
rlabel metal1 s 35760 0 35788 754 4 br_56
port 116 nsew
rlabel metal1 s 36384 0 36412 754 4 bl_57
port 117 nsew
rlabel metal1 s 36848 0 36876 754 4 br_57
port 118 nsew
rlabel metal1 s 37472 0 37500 754 4 bl_58
port 119 nsew
rlabel metal1 s 37008 0 37036 754 4 br_58
port 120 nsew
rlabel metal1 s 37632 0 37660 754 4 bl_59
port 121 nsew
rlabel metal1 s 38096 0 38124 754 4 br_59
port 122 nsew
rlabel metal1 s 38720 0 38748 754 4 bl_60
port 123 nsew
rlabel metal1 s 38256 0 38284 754 4 br_60
port 124 nsew
rlabel metal1 s 38880 0 38908 754 4 bl_61
port 125 nsew
rlabel metal1 s 39344 0 39372 754 4 br_61
port 126 nsew
rlabel metal1 s 39968 0 39996 754 4 bl_62
port 127 nsew
rlabel metal1 s 39504 0 39532 754 4 br_62
port 128 nsew
rlabel metal1 s 40128 0 40156 754 4 bl_63
port 129 nsew
rlabel metal1 s 40592 0 40620 754 4 br_63
port 130 nsew
rlabel metal1 s 40752 0 40780 754 4 br_64
port 131 nsew
rlabel metal1 s 41216 0 41244 754 4 bl_64
port 132 nsew
rlabel metal1 s 41376 0 41404 754 4 bl_65
port 133 nsew
rlabel metal1 s 41840 0 41868 754 4 br_65
port 134 nsew
rlabel metal1 s 42464 0 42492 754 4 bl_66
port 135 nsew
rlabel metal1 s 42000 0 42028 754 4 br_66
port 136 nsew
rlabel metal1 s 42624 0 42652 754 4 bl_67
port 137 nsew
rlabel metal1 s 43088 0 43116 754 4 br_67
port 138 nsew
rlabel metal1 s 43712 0 43740 754 4 bl_68
port 139 nsew
rlabel metal1 s 43248 0 43276 754 4 br_68
port 140 nsew
rlabel metal1 s 43872 0 43900 754 4 bl_69
port 141 nsew
rlabel metal1 s 44336 0 44364 754 4 br_69
port 142 nsew
rlabel metal1 s 44960 0 44988 754 4 bl_70
port 143 nsew
rlabel metal1 s 44496 0 44524 754 4 br_70
port 144 nsew
rlabel metal1 s 45120 0 45148 754 4 bl_71
port 145 nsew
rlabel metal1 s 45584 0 45612 754 4 br_71
port 146 nsew
rlabel metal1 s 46208 0 46236 754 4 bl_72
port 147 nsew
rlabel metal1 s 45744 0 45772 754 4 br_72
port 148 nsew
rlabel metal1 s 46368 0 46396 754 4 bl_73
port 149 nsew
rlabel metal1 s 46832 0 46860 754 4 br_73
port 150 nsew
rlabel metal1 s 47456 0 47484 754 4 bl_74
port 151 nsew
rlabel metal1 s 46992 0 47020 754 4 br_74
port 152 nsew
rlabel metal1 s 47616 0 47644 754 4 bl_75
port 153 nsew
rlabel metal1 s 48080 0 48108 754 4 br_75
port 154 nsew
rlabel metal1 s 48704 0 48732 754 4 bl_76
port 155 nsew
rlabel metal1 s 48240 0 48268 754 4 br_76
port 156 nsew
rlabel metal1 s 48864 0 48892 754 4 bl_77
port 157 nsew
rlabel metal1 s 49328 0 49356 754 4 br_77
port 158 nsew
rlabel metal1 s 49952 0 49980 754 4 bl_78
port 159 nsew
rlabel metal1 s 49488 0 49516 754 4 br_78
port 160 nsew
rlabel metal1 s 50112 0 50140 754 4 bl_79
port 161 nsew
rlabel metal1 s 50576 0 50604 754 4 br_79
port 162 nsew
rlabel metal1 s 51200 0 51228 754 4 bl_80
port 163 nsew
rlabel metal1 s 50736 0 50764 754 4 br_80
port 164 nsew
rlabel metal1 s 51360 0 51388 754 4 bl_81
port 165 nsew
rlabel metal1 s 51824 0 51852 754 4 br_81
port 166 nsew
rlabel metal1 s 52448 0 52476 754 4 bl_82
port 167 nsew
rlabel metal1 s 51984 0 52012 754 4 br_82
port 168 nsew
rlabel metal1 s 52608 0 52636 754 4 bl_83
port 169 nsew
rlabel metal1 s 53072 0 53100 754 4 br_83
port 170 nsew
rlabel metal1 s 53696 0 53724 754 4 bl_84
port 171 nsew
rlabel metal1 s 53232 0 53260 754 4 br_84
port 172 nsew
rlabel metal1 s 53856 0 53884 754 4 bl_85
port 173 nsew
rlabel metal1 s 54320 0 54348 754 4 br_85
port 174 nsew
rlabel metal1 s 54944 0 54972 754 4 bl_86
port 175 nsew
rlabel metal1 s 54480 0 54508 754 4 br_86
port 176 nsew
rlabel metal1 s 55104 0 55132 754 4 bl_87
port 177 nsew
rlabel metal1 s 55568 0 55596 754 4 br_87
port 178 nsew
rlabel metal1 s 56192 0 56220 754 4 bl_88
port 179 nsew
rlabel metal1 s 55728 0 55756 754 4 br_88
port 180 nsew
rlabel metal1 s 56352 0 56380 754 4 bl_89
port 181 nsew
rlabel metal1 s 56816 0 56844 754 4 br_89
port 182 nsew
rlabel metal1 s 57440 0 57468 754 4 bl_90
port 183 nsew
rlabel metal1 s 56976 0 57004 754 4 br_90
port 184 nsew
rlabel metal1 s 57600 0 57628 754 4 bl_91
port 185 nsew
rlabel metal1 s 58064 0 58092 754 4 br_91
port 186 nsew
rlabel metal1 s 58688 0 58716 754 4 bl_92
port 187 nsew
rlabel metal1 s 58224 0 58252 754 4 br_92
port 188 nsew
rlabel metal1 s 58848 0 58876 754 4 bl_93
port 189 nsew
rlabel metal1 s 59312 0 59340 754 4 br_93
port 190 nsew
rlabel metal1 s 59936 0 59964 754 4 bl_94
port 191 nsew
rlabel metal1 s 59472 0 59500 754 4 br_94
port 192 nsew
rlabel metal1 s 60096 0 60124 754 4 bl_95
port 193 nsew
rlabel metal1 s 60560 0 60588 754 4 br_95
port 194 nsew
rlabel metal1 s 60720 0 60748 754 4 br_96
port 195 nsew
rlabel metal1 s 61184 0 61212 754 4 bl_96
port 196 nsew
rlabel metal1 s 61344 0 61372 754 4 bl_97
port 197 nsew
rlabel metal1 s 61808 0 61836 754 4 br_97
port 198 nsew
rlabel metal1 s 62432 0 62460 754 4 bl_98
port 199 nsew
rlabel metal1 s 61968 0 61996 754 4 br_98
port 200 nsew
rlabel metal1 s 62592 0 62620 754 4 bl_99
port 201 nsew
rlabel metal1 s 63056 0 63084 754 4 br_99
port 202 nsew
rlabel metal1 s 63680 0 63708 754 4 bl_100
port 203 nsew
rlabel metal1 s 63216 0 63244 754 4 br_100
port 204 nsew
rlabel metal1 s 63840 0 63868 754 4 bl_101
port 205 nsew
rlabel metal1 s 64304 0 64332 754 4 br_101
port 206 nsew
rlabel metal1 s 64928 0 64956 754 4 bl_102
port 207 nsew
rlabel metal1 s 64464 0 64492 754 4 br_102
port 208 nsew
rlabel metal1 s 65088 0 65116 754 4 bl_103
port 209 nsew
rlabel metal1 s 65552 0 65580 754 4 br_103
port 210 nsew
rlabel metal1 s 66176 0 66204 754 4 bl_104
port 211 nsew
rlabel metal1 s 65712 0 65740 754 4 br_104
port 212 nsew
rlabel metal1 s 66336 0 66364 754 4 bl_105
port 213 nsew
rlabel metal1 s 66800 0 66828 754 4 br_105
port 214 nsew
rlabel metal1 s 67424 0 67452 754 4 bl_106
port 215 nsew
rlabel metal1 s 66960 0 66988 754 4 br_106
port 216 nsew
rlabel metal1 s 67584 0 67612 754 4 bl_107
port 217 nsew
rlabel metal1 s 68048 0 68076 754 4 br_107
port 218 nsew
rlabel metal1 s 68672 0 68700 754 4 bl_108
port 219 nsew
rlabel metal1 s 68208 0 68236 754 4 br_108
port 220 nsew
rlabel metal1 s 68832 0 68860 754 4 bl_109
port 221 nsew
rlabel metal1 s 69296 0 69324 754 4 br_109
port 222 nsew
rlabel metal1 s 69920 0 69948 754 4 bl_110
port 223 nsew
rlabel metal1 s 69456 0 69484 754 4 br_110
port 224 nsew
rlabel metal1 s 70080 0 70108 754 4 bl_111
port 225 nsew
rlabel metal1 s 70544 0 70572 754 4 br_111
port 226 nsew
rlabel metal1 s 71168 0 71196 754 4 bl_112
port 227 nsew
rlabel metal1 s 70704 0 70732 754 4 br_112
port 228 nsew
rlabel metal1 s 71328 0 71356 754 4 bl_113
port 229 nsew
rlabel metal1 s 71792 0 71820 754 4 br_113
port 230 nsew
rlabel metal1 s 72416 0 72444 754 4 bl_114
port 231 nsew
rlabel metal1 s 71952 0 71980 754 4 br_114
port 232 nsew
rlabel metal1 s 72576 0 72604 754 4 bl_115
port 233 nsew
rlabel metal1 s 73040 0 73068 754 4 br_115
port 234 nsew
rlabel metal1 s 73664 0 73692 754 4 bl_116
port 235 nsew
rlabel metal1 s 73200 0 73228 754 4 br_116
port 236 nsew
rlabel metal1 s 73824 0 73852 754 4 bl_117
port 237 nsew
rlabel metal1 s 74288 0 74316 754 4 br_117
port 238 nsew
rlabel metal1 s 74912 0 74940 754 4 bl_118
port 239 nsew
rlabel metal1 s 74448 0 74476 754 4 br_118
port 240 nsew
rlabel metal1 s 75072 0 75100 754 4 bl_119
port 241 nsew
rlabel metal1 s 75536 0 75564 754 4 br_119
port 242 nsew
rlabel metal1 s 76160 0 76188 754 4 bl_120
port 243 nsew
rlabel metal1 s 75696 0 75724 754 4 br_120
port 244 nsew
rlabel metal1 s 76320 0 76348 754 4 bl_121
port 245 nsew
rlabel metal1 s 76784 0 76812 754 4 br_121
port 246 nsew
rlabel metal1 s 77408 0 77436 754 4 bl_122
port 247 nsew
rlabel metal1 s 76944 0 76972 754 4 br_122
port 248 nsew
rlabel metal1 s 77568 0 77596 754 4 bl_123
port 249 nsew
rlabel metal1 s 78032 0 78060 754 4 br_123
port 250 nsew
rlabel metal1 s 78656 0 78684 754 4 bl_124
port 251 nsew
rlabel metal1 s 78192 0 78220 754 4 br_124
port 252 nsew
rlabel metal1 s 78816 0 78844 754 4 bl_125
port 253 nsew
rlabel metal1 s 79280 0 79308 754 4 br_125
port 254 nsew
rlabel metal1 s 79904 0 79932 754 4 bl_126
port 255 nsew
rlabel metal1 s 79440 0 79468 754 4 br_126
port 256 nsew
rlabel metal1 s 80064 0 80092 754 4 bl_127
port 257 nsew
rlabel metal1 s 80528 0 80556 754 4 br_127
port 258 nsew
rlabel metal1 s 81152 0 81180 754 4 bl_128
port 259 nsew
rlabel metal1 s 80688 0 80716 754 4 br_128
port 260 nsew
<< properties >>
string FIXED_BBOX 80901 -12 80967 0
string GDS_END 1610360
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 1522108
<< end >>
