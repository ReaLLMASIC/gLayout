magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 9 157 284 203
rect 642 157 918 203
rect 9 67 918 157
rect 30 -17 64 67
rect 286 21 918 67
<< scnmos >>
rect 87 93 117 177
rect 176 93 206 177
rect 364 47 394 131
rect 455 47 485 131
rect 539 47 569 131
rect 623 47 653 131
rect 721 47 751 177
rect 805 47 835 177
<< scpmoshvt >>
rect 79 410 109 494
rect 368 413 398 497
rect 176 297 206 381
rect 464 297 494 381
rect 536 297 566 381
rect 623 297 653 381
rect 721 297 751 497
rect 805 297 835 497
<< ndiff >>
rect 35 149 87 177
rect 35 115 43 149
rect 77 115 87 149
rect 35 93 87 115
rect 117 149 176 177
rect 117 115 132 149
rect 166 115 176 149
rect 117 93 176 115
rect 206 149 258 177
rect 206 115 216 149
rect 250 115 258 149
rect 668 131 721 177
rect 206 93 258 115
rect 312 97 364 131
rect 312 63 320 97
rect 354 63 364 97
rect 312 47 364 63
rect 394 111 455 131
rect 394 77 405 111
rect 439 77 455 111
rect 394 47 455 77
rect 485 97 539 131
rect 485 63 495 97
rect 529 63 539 97
rect 485 47 539 63
rect 569 111 623 131
rect 569 77 579 111
rect 613 77 623 111
rect 569 47 623 77
rect 653 97 721 131
rect 653 63 673 97
rect 707 63 721 97
rect 653 47 721 63
rect 751 135 805 177
rect 751 101 761 135
rect 795 101 805 135
rect 751 47 805 101
rect 835 163 892 177
rect 835 129 850 163
rect 884 129 892 163
rect 835 95 892 129
rect 835 61 850 95
rect 884 61 892 95
rect 835 47 892 61
<< pdiff >>
rect 27 475 79 494
rect 27 441 35 475
rect 69 441 79 475
rect 27 410 79 441
rect 109 475 161 494
rect 109 441 119 475
rect 153 441 161 475
rect 109 410 161 441
rect 316 475 368 497
rect 316 441 324 475
rect 358 441 368 475
rect 316 413 368 441
rect 398 413 449 497
rect 668 485 721 497
rect 668 451 676 485
rect 710 451 721 485
rect 124 381 161 410
rect 124 297 176 381
rect 206 339 262 381
rect 206 305 216 339
rect 250 305 262 339
rect 206 297 262 305
rect 413 381 449 413
rect 668 417 721 451
rect 668 383 676 417
rect 710 383 721 417
rect 668 381 721 383
rect 413 297 464 381
rect 494 297 536 381
rect 566 297 623 381
rect 653 297 721 381
rect 751 454 805 497
rect 751 420 761 454
rect 795 420 805 454
rect 751 386 805 420
rect 751 352 761 386
rect 795 352 805 386
rect 751 297 805 352
rect 835 485 892 497
rect 835 451 850 485
rect 884 451 892 485
rect 835 417 892 451
rect 835 383 850 417
rect 884 383 892 417
rect 835 349 892 383
rect 835 315 850 349
rect 884 315 892 349
rect 835 297 892 315
<< ndiffc >>
rect 43 115 77 149
rect 132 115 166 149
rect 216 115 250 149
rect 320 63 354 97
rect 405 77 439 111
rect 495 63 529 97
rect 579 77 613 111
rect 673 63 707 97
rect 761 101 795 135
rect 850 129 884 163
rect 850 61 884 95
<< pdiffc >>
rect 35 441 69 475
rect 119 441 153 475
rect 324 441 358 475
rect 676 451 710 485
rect 216 305 250 339
rect 676 383 710 417
rect 761 420 795 454
rect 761 352 795 386
rect 850 451 884 485
rect 850 383 884 417
rect 850 315 884 349
<< poly >>
rect 79 494 109 520
rect 368 497 398 523
rect 721 497 751 523
rect 805 497 835 523
rect 530 484 596 494
rect 530 450 546 484
rect 580 450 596 484
rect 530 440 596 450
rect 79 265 109 410
rect 176 381 206 407
rect 176 265 206 297
rect 368 265 398 413
rect 464 381 494 407
rect 536 381 566 440
rect 623 381 653 407
rect 464 265 494 297
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 174 249 240 265
rect 174 215 190 249
rect 224 215 240 249
rect 174 199 240 215
rect 307 249 398 265
rect 307 215 317 249
rect 351 215 398 249
rect 307 199 398 215
rect 440 249 494 265
rect 440 215 450 249
rect 484 215 494 249
rect 440 199 494 215
rect 87 177 117 199
rect 176 177 206 199
rect 364 131 394 199
rect 455 131 485 199
rect 536 182 566 297
rect 623 265 653 297
rect 721 265 751 297
rect 805 265 835 297
rect 608 249 662 265
rect 608 215 618 249
rect 652 215 662 249
rect 608 199 662 215
rect 704 249 835 265
rect 704 215 714 249
rect 748 215 835 249
rect 704 199 835 215
rect 536 152 569 182
rect 539 131 569 152
rect 623 131 653 199
rect 721 177 751 199
rect 805 177 835 199
rect 87 67 117 93
rect 176 67 206 93
rect 364 21 394 47
rect 455 21 485 47
rect 539 21 569 47
rect 623 21 653 47
rect 721 21 751 47
rect 805 21 835 47
<< polycont >>
rect 546 450 580 484
rect 86 215 120 249
rect 190 215 224 249
rect 317 215 351 249
rect 450 215 484 249
rect 618 215 652 249
rect 714 215 748 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 475 169 527
rect 501 484 629 491
rect 103 441 119 475
rect 153 441 169 475
rect 307 441 324 475
rect 358 441 456 475
rect 17 407 69 441
rect 17 373 388 407
rect 17 165 52 373
rect 86 249 156 339
rect 199 305 216 339
rect 250 305 320 339
rect 120 215 156 249
rect 86 199 156 215
rect 190 249 248 265
rect 224 215 248 249
rect 190 199 248 215
rect 282 249 320 305
rect 354 317 388 373
rect 422 391 456 441
rect 501 450 546 484
rect 580 450 629 484
rect 501 425 629 450
rect 663 485 719 527
rect 663 451 676 485
rect 710 451 719 485
rect 663 417 719 451
rect 422 357 629 391
rect 663 383 676 417
rect 710 383 719 417
rect 663 367 719 383
rect 761 454 816 493
rect 795 420 816 454
rect 761 386 816 420
rect 595 333 629 357
rect 795 352 816 386
rect 354 283 484 317
rect 595 299 727 333
rect 761 299 816 352
rect 450 249 484 283
rect 693 265 727 299
rect 282 215 317 249
rect 351 215 371 249
rect 282 165 320 215
rect 450 199 484 215
rect 528 249 659 265
rect 528 215 618 249
rect 652 215 659 249
rect 528 199 659 215
rect 693 249 748 265
rect 693 215 714 249
rect 693 199 748 215
rect 693 165 727 199
rect 17 149 81 165
rect 17 115 43 149
rect 77 115 81 149
rect 17 90 81 115
rect 132 149 166 165
rect 132 17 166 115
rect 216 149 320 165
rect 250 131 320 149
rect 405 131 727 165
rect 782 152 816 299
rect 850 485 884 527
rect 850 417 884 451
rect 850 349 884 383
rect 850 288 884 315
rect 761 135 816 152
rect 216 90 250 115
rect 405 111 439 131
rect 299 63 320 97
rect 354 63 370 97
rect 299 17 370 63
rect 579 111 613 131
rect 405 61 439 77
rect 479 63 495 97
rect 529 63 545 97
rect 479 17 545 63
rect 795 101 816 135
rect 579 61 613 77
rect 647 63 673 97
rect 707 63 723 97
rect 761 83 816 101
rect 850 163 884 205
rect 850 95 884 129
rect 647 17 723 63
rect 850 17 884 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 586 221 620 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 770 357 804 391 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 586 425 620 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 or4bb_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1105288
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1097680
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
