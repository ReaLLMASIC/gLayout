magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect -50 -112 0 -96
rect -50 -146 -34 -112
rect -50 -162 0 -146
<< polycont >>
rect -34 16 0 50
rect -34 -146 0 -112
<< npolyres >>
rect 0 0 23637 66
rect 23571 -96 23637 0
rect 0 -162 23637 -96
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect -34 -112 0 -96
rect -34 -162 0 -146
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1701704242
transform 1 0 -50 0 1 -162
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1701704242
transform 1 0 -50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 98009526
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98008790
<< end >>
