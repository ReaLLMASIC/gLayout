magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -66 377 4098 897
<< pwell >>
rect 1330 226 1890 230
rect 1064 217 1890 226
rect 2215 217 4028 283
rect 9 43 4028 217
rect -26 -43 4058 43
<< mvnmos >>
rect 92 107 192 191
rect 248 107 348 191
rect 390 107 490 191
rect 546 107 646 191
rect 688 107 788 191
rect 877 107 977 191
rect 1143 116 1243 200
rect 1413 120 1513 204
rect 1569 120 1669 204
rect 1711 120 1811 204
rect 1977 107 2077 191
rect 2119 107 2219 191
rect 2294 107 2394 257
rect 2436 107 2536 257
rect 2615 173 2715 257
rect 2757 173 2857 257
rect 2899 173 2999 257
rect 3207 173 3307 257
rect 3386 107 3486 257
rect 3666 173 3766 257
rect 3845 107 3945 257
<< mvpmos >>
rect 87 569 187 653
rect 243 569 343 653
rect 385 569 485 653
rect 541 569 641 653
rect 683 569 783 653
rect 872 569 972 719
rect 1184 488 1284 638
rect 1454 556 1554 640
rect 1610 556 1710 640
rect 1752 556 1852 640
rect 1924 556 2024 640
rect 2080 556 2180 640
rect 2259 543 2359 743
rect 2401 543 2501 743
rect 2587 543 2687 627
rect 2729 543 2829 627
rect 2899 543 2999 627
rect 3221 443 3321 527
rect 3396 443 3496 743
rect 3666 479 3766 629
rect 3845 479 3945 679
<< mvndiff >>
rect 35 166 92 191
rect 35 132 47 166
rect 81 132 92 166
rect 35 107 92 132
rect 192 166 248 191
rect 192 132 203 166
rect 237 132 248 166
rect 192 107 248 132
rect 348 107 390 191
rect 490 166 546 191
rect 490 132 501 166
rect 535 132 546 166
rect 490 107 546 132
rect 646 107 688 191
rect 788 166 877 191
rect 788 132 799 166
rect 833 132 877 166
rect 788 107 877 132
rect 977 166 1030 191
rect 977 132 988 166
rect 1022 132 1030 166
rect 977 107 1030 132
rect 1090 175 1143 200
rect 1090 141 1098 175
rect 1132 141 1143 175
rect 1090 116 1143 141
rect 1243 175 1296 200
rect 1243 141 1254 175
rect 1288 141 1296 175
rect 1243 116 1296 141
rect 1356 184 1413 204
rect 1356 150 1368 184
rect 1402 150 1413 184
rect 1356 120 1413 150
rect 1513 179 1569 204
rect 1513 145 1524 179
rect 1558 145 1569 179
rect 1513 120 1569 145
rect 1669 120 1711 204
rect 1811 179 1864 204
rect 2241 191 2294 257
rect 1811 145 1822 179
rect 1856 145 1864 179
rect 1811 120 1864 145
rect 1924 166 1977 191
rect 1924 132 1932 166
rect 1966 132 1977 166
rect 1924 107 1977 132
rect 2077 107 2119 191
rect 2219 179 2294 191
rect 2219 145 2249 179
rect 2283 145 2294 179
rect 2219 107 2294 145
rect 2394 107 2436 257
rect 2536 249 2615 257
rect 2536 215 2547 249
rect 2581 215 2615 249
rect 2536 173 2615 215
rect 2715 173 2757 257
rect 2857 173 2899 257
rect 2999 232 3056 257
rect 2999 198 3010 232
rect 3044 198 3056 232
rect 2999 173 3056 198
rect 3150 232 3207 257
rect 3150 198 3162 232
rect 3196 198 3207 232
rect 3150 173 3207 198
rect 3307 249 3386 257
rect 3307 215 3341 249
rect 3375 215 3386 249
rect 3307 173 3386 215
rect 2536 157 2593 173
rect 2536 123 2547 157
rect 2581 123 2593 157
rect 3329 149 3386 173
rect 2536 107 2593 123
rect 3329 115 3341 149
rect 3375 115 3386 149
rect 3329 107 3386 115
rect 3486 249 3543 257
rect 3486 215 3497 249
rect 3531 215 3543 249
rect 3486 149 3543 215
rect 3609 232 3666 257
rect 3609 198 3621 232
rect 3655 198 3666 232
rect 3609 173 3666 198
rect 3766 249 3845 257
rect 3766 215 3800 249
rect 3834 215 3845 249
rect 3766 173 3845 215
rect 3486 115 3497 149
rect 3531 115 3543 149
rect 3788 149 3845 173
rect 3486 107 3543 115
rect 3788 115 3800 149
rect 3834 115 3845 149
rect 3788 107 3845 115
rect 3945 249 4002 257
rect 3945 215 3956 249
rect 3990 215 4002 249
rect 3945 149 4002 215
rect 3945 115 3956 149
rect 3990 115 4002 149
rect 3945 107 4002 115
<< mvpdiff >>
rect 2202 719 2259 743
rect 815 711 872 719
rect 815 677 827 711
rect 861 677 872 711
rect 815 653 872 677
rect 30 628 87 653
rect 30 594 42 628
rect 76 594 87 628
rect 30 569 87 594
rect 187 628 243 653
rect 187 594 198 628
rect 232 594 243 628
rect 187 569 243 594
rect 343 569 385 653
rect 485 628 541 653
rect 485 594 496 628
rect 530 594 541 628
rect 485 569 541 594
rect 641 569 683 653
rect 783 611 872 653
rect 783 577 827 611
rect 861 577 872 611
rect 783 569 872 577
rect 972 691 1029 719
rect 972 657 983 691
rect 1017 657 1029 691
rect 2202 685 2214 719
rect 2248 685 2259 719
rect 972 611 1029 657
rect 2202 640 2259 685
rect 972 577 983 611
rect 1017 577 1029 611
rect 972 569 1029 577
rect 1127 630 1184 638
rect 1127 596 1139 630
rect 1173 596 1184 630
rect 1127 530 1184 596
rect 1127 496 1139 530
rect 1173 496 1184 530
rect 1127 488 1184 496
rect 1284 626 1337 638
rect 1284 592 1295 626
rect 1329 592 1337 626
rect 1284 534 1337 592
rect 1397 615 1454 640
rect 1397 581 1409 615
rect 1443 581 1454 615
rect 1397 556 1454 581
rect 1554 615 1610 640
rect 1554 581 1565 615
rect 1599 581 1610 615
rect 1554 556 1610 581
rect 1710 556 1752 640
rect 1852 629 1924 640
rect 1852 595 1863 629
rect 1897 595 1924 629
rect 1852 556 1924 595
rect 2024 598 2080 640
rect 2024 564 2035 598
rect 2069 564 2080 598
rect 2024 556 2080 564
rect 2180 556 2259 640
rect 1284 500 1295 534
rect 1329 500 1337 534
rect 1284 488 1337 500
rect 2202 543 2259 556
rect 2359 543 2401 743
rect 2501 735 2565 743
rect 2501 701 2519 735
rect 2553 701 2565 735
rect 2501 660 2565 701
rect 2501 626 2519 660
rect 2553 627 2565 660
rect 3343 731 3396 743
rect 3343 697 3351 731
rect 3385 697 3396 731
rect 3343 651 3396 697
rect 2553 626 2587 627
rect 2501 585 2587 626
rect 2501 551 2519 585
rect 2553 551 2587 585
rect 2501 543 2587 551
rect 2687 543 2729 627
rect 2829 614 2899 627
rect 2829 580 2840 614
rect 2874 580 2899 614
rect 2829 543 2899 580
rect 2999 602 3056 627
rect 2999 568 3010 602
rect 3044 568 3056 602
rect 2999 543 3056 568
rect 3343 617 3351 651
rect 3385 617 3396 651
rect 3343 569 3396 617
rect 3343 535 3351 569
rect 3385 535 3396 569
rect 3343 527 3396 535
rect 3141 502 3221 527
rect 3141 468 3153 502
rect 3187 468 3221 502
rect 3141 443 3221 468
rect 3321 489 3396 527
rect 3321 455 3351 489
rect 3385 455 3396 489
rect 3321 443 3396 455
rect 3496 731 3549 743
rect 3496 697 3507 731
rect 3541 697 3549 731
rect 3496 651 3549 697
rect 3788 671 3845 679
rect 3496 617 3507 651
rect 3541 617 3549 651
rect 3788 637 3800 671
rect 3834 637 3845 671
rect 3788 629 3845 637
rect 3496 569 3549 617
rect 3496 535 3507 569
rect 3541 535 3549 569
rect 3496 489 3549 535
rect 3496 455 3507 489
rect 3541 455 3549 489
rect 3609 621 3666 629
rect 3609 587 3621 621
rect 3655 587 3666 621
rect 3609 521 3666 587
rect 3609 487 3621 521
rect 3655 487 3666 521
rect 3609 479 3666 487
rect 3766 596 3845 629
rect 3766 562 3800 596
rect 3834 562 3845 596
rect 3766 521 3845 562
rect 3766 487 3800 521
rect 3834 487 3845 521
rect 3766 479 3845 487
rect 3945 671 4002 679
rect 3945 637 3956 671
rect 3990 637 4002 671
rect 3945 596 4002 637
rect 3945 562 3956 596
rect 3990 562 4002 596
rect 3945 521 4002 562
rect 3945 487 3956 521
rect 3990 487 4002 521
rect 3945 479 4002 487
rect 3496 443 3549 455
<< mvndiffc >>
rect 47 132 81 166
rect 203 132 237 166
rect 501 132 535 166
rect 799 132 833 166
rect 988 132 1022 166
rect 1098 141 1132 175
rect 1254 141 1288 175
rect 1368 150 1402 184
rect 1524 145 1558 179
rect 1822 145 1856 179
rect 1932 132 1966 166
rect 2249 145 2283 179
rect 2547 215 2581 249
rect 3010 198 3044 232
rect 3162 198 3196 232
rect 3341 215 3375 249
rect 2547 123 2581 157
rect 3341 115 3375 149
rect 3497 215 3531 249
rect 3621 198 3655 232
rect 3800 215 3834 249
rect 3497 115 3531 149
rect 3800 115 3834 149
rect 3956 215 3990 249
rect 3956 115 3990 149
<< mvpdiffc >>
rect 827 677 861 711
rect 42 594 76 628
rect 198 594 232 628
rect 496 594 530 628
rect 827 577 861 611
rect 983 657 1017 691
rect 2214 685 2248 719
rect 983 577 1017 611
rect 1139 596 1173 630
rect 1139 496 1173 530
rect 1295 592 1329 626
rect 1409 581 1443 615
rect 1565 581 1599 615
rect 1863 595 1897 629
rect 2035 564 2069 598
rect 1295 500 1329 534
rect 2519 701 2553 735
rect 2519 626 2553 660
rect 3351 697 3385 731
rect 2519 551 2553 585
rect 2840 580 2874 614
rect 3010 568 3044 602
rect 3351 617 3385 651
rect 3351 535 3385 569
rect 3153 468 3187 502
rect 3351 455 3385 489
rect 3507 697 3541 731
rect 3507 617 3541 651
rect 3800 637 3834 671
rect 3507 535 3541 569
rect 3507 455 3541 489
rect 3621 587 3655 621
rect 3621 487 3655 521
rect 3800 562 3834 596
rect 3800 487 3834 521
rect 3956 637 3990 671
rect 3956 562 3990 596
rect 3956 487 3990 521
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
<< poly >>
rect 872 719 972 745
rect 2259 743 2359 769
rect 2401 743 2501 769
rect 3396 743 3496 769
rect 87 653 187 679
rect 243 653 343 679
rect 385 653 485 679
rect 541 653 641 679
rect 683 653 783 679
rect 1184 638 1284 664
rect 1454 640 1554 666
rect 1610 640 1710 666
rect 1752 640 1852 666
rect 1924 640 2024 666
rect 2080 640 2180 666
rect 87 547 187 569
rect 243 547 343 569
rect 87 464 343 547
rect 385 471 485 569
rect 541 543 641 569
rect 87 417 192 464
rect 385 437 411 471
rect 445 437 485 471
rect 385 422 485 437
rect 87 383 138 417
rect 172 383 192 417
rect 87 349 192 383
rect 87 315 138 349
rect 172 315 192 349
rect 87 217 192 315
rect 92 191 192 217
rect 248 403 485 422
rect 248 369 411 403
rect 445 369 485 403
rect 527 521 641 543
rect 527 487 543 521
rect 577 487 641 521
rect 527 453 641 487
rect 527 419 543 453
rect 577 443 641 453
rect 683 543 783 569
rect 683 443 788 543
rect 577 419 627 443
rect 527 399 627 419
rect 248 338 485 369
rect 248 191 348 338
rect 532 337 646 357
rect 532 303 552 337
rect 586 303 646 337
rect 390 263 490 296
rect 390 229 410 263
rect 444 229 490 263
rect 390 191 490 229
rect 532 269 646 303
rect 532 235 552 269
rect 586 235 646 269
rect 532 215 646 235
rect 546 191 646 215
rect 688 339 788 443
rect 688 305 704 339
rect 738 305 788 339
rect 688 271 788 305
rect 872 434 972 569
rect 1454 534 1554 556
rect 1434 508 1554 534
rect 1610 530 1710 556
rect 872 414 977 434
rect 872 380 892 414
rect 926 380 977 414
rect 872 346 977 380
rect 1184 378 1284 488
rect 1434 474 1454 508
rect 1488 474 1554 508
rect 1434 454 1554 474
rect 1602 508 1710 530
rect 1602 474 1656 508
rect 1690 474 1710 508
rect 1602 412 1710 474
rect 1752 486 1852 556
rect 1752 452 1798 486
rect 1832 452 1852 486
rect 872 312 892 346
rect 926 312 977 346
rect 872 292 977 312
rect 688 237 704 271
rect 738 237 788 271
rect 688 191 788 237
rect 877 191 977 292
rect 1143 358 1284 378
rect 1143 324 1163 358
rect 1197 326 1284 358
rect 1413 342 1702 412
rect 1413 326 1513 342
rect 1197 324 1513 326
rect 1143 290 1513 324
rect 1752 300 1852 452
rect 1143 256 1163 290
rect 1197 256 1513 290
rect 1143 226 1513 256
rect 1143 200 1243 226
rect 1413 204 1513 226
rect 1569 280 1669 300
rect 1569 246 1615 280
rect 1649 246 1669 280
rect 1569 204 1669 246
rect 1711 276 1852 300
rect 1711 242 1798 276
rect 1832 242 1852 276
rect 1711 226 1852 242
rect 1924 416 2024 556
rect 1924 382 1970 416
rect 2004 382 2024 416
rect 1924 289 2024 382
rect 2080 431 2180 556
rect 2587 627 2687 653
rect 2729 627 2829 653
rect 2899 627 2999 653
rect 2259 495 2359 543
rect 2259 461 2279 495
rect 2313 461 2359 495
rect 2080 331 2217 431
rect 2259 427 2359 461
rect 2259 393 2279 427
rect 2313 393 2359 427
rect 2401 517 2501 543
rect 2587 521 2687 543
rect 2401 475 2488 517
rect 2543 475 2687 521
rect 2401 441 2421 475
rect 2455 441 2488 475
rect 2401 421 2488 441
rect 2530 459 2687 475
rect 2729 521 2829 543
rect 2729 469 2857 521
rect 2729 463 2803 469
rect 2259 379 2359 393
rect 2530 379 2582 459
rect 2757 435 2803 463
rect 2837 435 2857 469
rect 2259 373 2394 379
rect 1711 204 1811 226
rect 1924 213 2077 289
rect 1977 191 2077 213
rect 2119 276 2219 331
rect 2119 242 2139 276
rect 2173 242 2219 276
rect 2294 257 2394 373
rect 2436 359 2582 379
rect 2436 325 2456 359
rect 2490 325 2582 359
rect 2624 401 2715 417
rect 2624 367 2640 401
rect 2674 367 2715 401
rect 2624 333 2715 367
rect 2436 257 2536 325
rect 2624 299 2640 333
rect 2674 299 2715 333
rect 2624 283 2715 299
rect 2615 257 2715 283
rect 2757 257 2857 435
rect 2899 329 2999 543
rect 3221 527 3321 553
rect 3845 679 3945 705
rect 3666 629 3766 655
rect 3221 419 3321 443
rect 3396 419 3496 443
rect 3666 419 3766 479
rect 2899 295 2919 329
rect 2953 295 2999 329
rect 2899 257 2999 295
rect 3041 399 3766 419
rect 3041 365 3059 399
rect 3093 365 3766 399
rect 3041 331 3766 365
rect 3041 297 3059 331
rect 3093 319 3766 331
rect 3093 297 3307 319
rect 3041 279 3307 297
rect 3207 257 3307 279
rect 3386 257 3486 319
rect 3666 257 3766 319
rect 3845 419 3945 479
rect 3845 385 3865 419
rect 3899 385 3945 419
rect 3845 351 3945 385
rect 3845 317 3865 351
rect 3899 317 3945 351
rect 3845 257 3945 317
rect 2119 191 2219 242
rect 92 81 192 107
rect 248 81 348 107
rect 390 81 490 107
rect 546 81 646 107
rect 688 81 788 107
rect 877 81 977 107
rect 1143 90 1243 116
rect 1413 94 1513 120
rect 1569 94 1669 120
rect 1711 94 1811 120
rect 2615 147 2715 173
rect 2757 147 2857 173
rect 2899 147 2999 173
rect 3207 147 3307 173
rect 3666 147 3766 173
rect 1977 81 2077 107
rect 2119 81 2219 107
rect 2294 81 2394 107
rect 2436 81 2536 107
rect 3386 81 3486 107
rect 3845 81 3945 107
<< polycont >>
rect 411 437 445 471
rect 138 383 172 417
rect 138 315 172 349
rect 411 369 445 403
rect 543 487 577 521
rect 543 419 577 453
rect 552 303 586 337
rect 410 229 444 263
rect 552 235 586 269
rect 704 305 738 339
rect 892 380 926 414
rect 1454 474 1488 508
rect 1656 474 1690 508
rect 1798 452 1832 486
rect 892 312 926 346
rect 704 237 738 271
rect 1163 324 1197 358
rect 1163 256 1197 290
rect 1615 246 1649 280
rect 1798 242 1832 276
rect 1970 382 2004 416
rect 2279 461 2313 495
rect 2279 393 2313 427
rect 2421 441 2455 475
rect 2803 435 2837 469
rect 2139 242 2173 276
rect 2456 325 2490 359
rect 2640 367 2674 401
rect 2640 299 2674 333
rect 2919 295 2953 329
rect 3059 365 3093 399
rect 3059 297 3093 331
rect 3865 385 3899 419
rect 3865 317 3899 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 128 735 318 741
rect 128 701 134 735
rect 168 701 206 735
rect 240 701 278 735
rect 312 701 318 735
rect 26 628 92 661
rect 26 594 42 628
rect 76 594 92 628
rect 26 541 92 594
rect 128 628 318 701
rect 683 735 861 741
rect 717 701 755 735
rect 789 701 827 735
rect 683 677 827 701
rect 128 594 198 628
rect 232 594 318 628
rect 128 577 318 594
rect 480 628 546 661
rect 480 594 496 628
rect 530 611 546 628
rect 683 611 861 677
rect 530 594 647 611
rect 480 577 647 594
rect 26 521 577 541
rect 26 507 543 521
rect 26 263 60 507
rect 527 487 543 507
rect 613 525 647 577
rect 683 577 827 611
rect 683 561 861 577
rect 897 727 1103 761
rect 897 525 931 727
rect 967 657 983 691
rect 1017 657 1033 691
rect 967 611 1033 657
rect 967 577 983 611
rect 1017 577 1033 611
rect 967 561 1033 577
rect 613 491 931 525
rect 395 437 411 471
rect 445 437 461 471
rect 121 417 359 433
rect 121 383 138 417
rect 172 383 359 417
rect 121 349 359 383
rect 395 403 461 437
rect 527 453 577 487
rect 527 419 543 453
rect 527 403 577 419
rect 395 369 411 403
rect 445 369 461 403
rect 121 315 138 349
rect 172 333 359 349
rect 536 337 591 353
rect 536 333 552 337
rect 172 315 552 333
rect 121 303 552 315
rect 586 303 591 337
rect 121 299 591 303
rect 536 269 591 299
rect 26 229 410 263
rect 444 229 460 263
rect 26 219 460 229
rect 536 235 552 269
rect 586 235 591 269
rect 536 219 591 235
rect 26 166 97 219
rect 627 183 661 491
rect 26 132 47 166
rect 81 132 97 166
rect 26 99 97 132
rect 133 166 323 183
rect 133 132 203 166
rect 237 132 323 166
rect 133 113 323 132
rect 133 79 139 113
rect 173 79 211 113
rect 245 79 283 113
rect 317 79 323 113
rect 485 166 661 183
rect 485 132 501 166
rect 535 149 661 166
rect 697 339 738 430
rect 697 305 704 339
rect 697 271 738 305
rect 697 237 704 271
rect 697 162 738 237
rect 876 414 942 430
rect 876 380 892 414
rect 926 380 942 414
rect 876 346 942 380
rect 876 312 892 346
rect 926 312 942 346
rect 876 236 942 312
rect 988 374 1033 561
rect 1069 444 1103 727
rect 1139 735 1173 741
rect 1723 735 1913 741
rect 1139 630 1173 701
rect 1139 530 1173 596
rect 1139 480 1173 496
rect 1209 678 1459 712
rect 1209 444 1243 678
rect 1069 410 1243 444
rect 1279 626 1329 642
rect 1279 592 1295 626
rect 1279 534 1329 592
rect 1279 500 1295 534
rect 1279 458 1329 500
rect 1368 615 1459 678
rect 1723 701 1729 735
rect 1763 701 1801 735
rect 1835 701 1873 735
rect 1907 701 1913 735
rect 1368 581 1409 615
rect 1443 581 1459 615
rect 1368 548 1459 581
rect 1540 615 1599 648
rect 1540 581 1565 615
rect 1723 629 1913 701
rect 2191 735 2381 751
rect 2191 701 2197 735
rect 2231 719 2269 735
rect 2248 701 2269 719
rect 2303 701 2341 735
rect 2375 701 2381 735
rect 2191 685 2214 701
rect 2248 685 2381 701
rect 2191 670 2381 685
rect 2503 735 2569 751
rect 2503 701 2519 735
rect 2553 701 2569 735
rect 1723 595 1863 629
rect 1897 595 1913 629
rect 1723 592 1913 595
rect 1949 634 2155 668
rect 2503 660 2569 701
rect 988 358 1213 374
rect 988 340 1163 358
rect 774 166 952 199
rect 535 132 551 149
rect 485 99 551 132
rect 774 132 799 166
rect 833 132 952 166
rect 774 113 952 132
rect 133 73 323 79
rect 808 79 846 113
rect 880 79 918 113
rect 988 166 1038 340
rect 1147 324 1163 340
rect 1197 324 1213 358
rect 1147 290 1213 324
rect 1147 256 1163 290
rect 1197 256 1213 290
rect 1147 240 1213 256
rect 1279 204 1313 458
rect 1368 212 1402 548
rect 1022 132 1038 166
rect 988 103 1038 132
rect 1074 175 1192 204
rect 1074 141 1098 175
rect 1132 141 1192 175
rect 1074 113 1192 141
rect 774 73 952 79
rect 1074 79 1080 113
rect 1114 79 1152 113
rect 1186 79 1192 113
rect 1074 73 1192 79
rect 1238 175 1313 204
rect 1238 141 1254 175
rect 1288 141 1313 175
rect 1238 87 1313 141
rect 1352 184 1402 212
rect 1352 150 1368 184
rect 1352 123 1402 150
rect 1438 508 1504 512
rect 1438 474 1454 508
rect 1488 474 1504 508
rect 1438 458 1504 474
rect 1438 87 1472 458
rect 1540 416 1599 581
rect 1949 556 1983 634
rect 2121 600 2467 634
rect 1640 522 1983 556
rect 2019 564 2035 598
rect 2069 564 2085 598
rect 1640 508 1706 522
rect 1640 474 1656 508
rect 1690 474 1706 508
rect 2019 486 2085 564
rect 1640 458 1706 474
rect 1782 452 1798 486
rect 1832 452 2085 486
rect 2263 495 2329 511
rect 2263 461 2279 495
rect 2313 461 2329 495
rect 2263 427 2329 461
rect 2263 416 2279 427
rect 1540 382 1970 416
rect 2004 393 2279 416
rect 2313 393 2329 427
rect 2405 475 2467 600
rect 2503 626 2519 660
rect 2553 626 2569 660
rect 2503 585 2569 626
rect 2503 551 2519 585
rect 2553 551 2569 585
rect 2700 735 2890 741
rect 2700 701 2706 735
rect 2740 701 2778 735
rect 2812 701 2850 735
rect 2884 701 2890 735
rect 2700 614 2890 701
rect 3248 735 3438 747
rect 3248 701 3254 735
rect 3288 701 3326 735
rect 3360 731 3398 735
rect 3385 701 3398 731
rect 3432 701 3438 735
rect 3248 697 3351 701
rect 3385 697 3438 701
rect 3248 651 3438 697
rect 2700 580 2840 614
rect 2874 580 2890 614
rect 2700 575 2890 580
rect 2994 602 3060 635
rect 2503 539 2569 551
rect 2994 568 3010 602
rect 3044 568 3060 602
rect 2994 539 3060 568
rect 2503 505 3060 539
rect 3248 617 3351 651
rect 3385 617 3438 651
rect 3248 569 3438 617
rect 3248 535 3351 569
rect 3385 535 3438 569
rect 2405 441 2421 475
rect 2455 459 2467 475
rect 2455 441 2681 459
rect 2405 425 2681 441
rect 2004 382 2329 393
rect 2633 401 2681 425
rect 1540 212 1574 382
rect 2440 359 2506 375
rect 2440 346 2456 359
rect 1508 179 1574 212
rect 1508 145 1524 179
rect 1558 145 1574 179
rect 1508 128 1574 145
rect 1610 325 2456 346
rect 2490 325 2506 359
rect 1610 312 2506 325
rect 2633 367 2640 401
rect 2674 367 2681 401
rect 2633 333 2681 367
rect 1610 280 1665 312
rect 2633 299 2640 333
rect 2674 299 2681 333
rect 2633 283 2681 299
rect 2717 399 2751 505
rect 3137 502 3212 535
rect 3137 469 3153 502
rect 2787 435 2803 469
rect 2837 468 3153 469
rect 3187 468 3212 502
rect 2837 435 3212 468
rect 3248 489 3438 535
rect 3248 455 3351 489
rect 3385 455 3438 489
rect 3248 439 3438 455
rect 3481 731 3557 747
rect 3481 697 3507 731
rect 3541 697 3557 731
rect 3481 651 3557 697
rect 3481 617 3507 651
rect 3541 617 3557 651
rect 3707 735 3897 741
rect 3707 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 3897 735
rect 3707 671 3897 701
rect 3707 637 3800 671
rect 3834 637 3897 671
rect 3481 569 3557 617
rect 3481 535 3507 569
rect 3541 535 3557 569
rect 3481 489 3557 535
rect 3481 455 3507 489
rect 3541 455 3557 489
rect 2717 365 3059 399
rect 3093 365 3109 399
rect 1610 246 1615 280
rect 1649 246 1665 280
rect 1610 230 1665 246
rect 1782 242 1798 276
rect 1832 242 1982 276
rect 2041 242 2139 276
rect 2173 242 2471 276
rect 1610 87 1644 230
rect 1782 228 1982 242
rect 1238 53 1644 87
rect 1682 179 1872 192
rect 1682 145 1822 179
rect 1856 145 1872 179
rect 1682 113 1872 145
rect 1682 79 1688 113
rect 1722 79 1760 113
rect 1794 79 1832 113
rect 1866 79 1872 113
rect 1916 166 1982 228
rect 1916 132 1932 166
rect 1966 132 1982 166
rect 1916 103 1982 132
rect 2109 179 2299 206
rect 2109 145 2249 179
rect 2283 145 2299 179
rect 2109 113 2299 145
rect 1682 73 1872 79
rect 2109 79 2115 113
rect 2149 79 2187 113
rect 2221 79 2259 113
rect 2293 79 2299 113
rect 2109 73 2299 79
rect 2437 87 2471 242
rect 2531 249 2597 265
rect 2531 215 2547 249
rect 2581 215 2597 249
rect 2531 157 2597 215
rect 2717 157 2751 365
rect 3043 331 3109 365
rect 2531 123 2547 157
rect 2581 123 2751 157
rect 2800 295 2919 329
rect 2953 295 2969 329
rect 2800 285 2969 295
rect 3043 297 3059 331
rect 3093 297 3109 331
rect 3043 285 3109 297
rect 2800 87 2834 285
rect 2437 53 2834 87
rect 2870 232 3060 249
rect 2870 198 3010 232
rect 3044 198 3060 232
rect 2870 113 3060 198
rect 3146 232 3212 435
rect 3146 198 3162 232
rect 3196 198 3212 232
rect 3146 165 3212 198
rect 3248 249 3438 265
rect 3248 215 3341 249
rect 3375 215 3438 249
rect 2870 79 2876 113
rect 2910 79 2948 113
rect 2982 79 3020 113
rect 3054 79 3060 113
rect 2870 73 3060 79
rect 3248 149 3438 215
rect 3248 115 3341 149
rect 3375 115 3438 149
rect 3248 113 3438 115
rect 3248 79 3254 113
rect 3288 79 3326 113
rect 3360 79 3398 113
rect 3432 79 3438 113
rect 3481 249 3557 455
rect 3481 215 3497 249
rect 3531 215 3557 249
rect 3481 149 3557 215
rect 3605 621 3671 637
rect 3605 587 3621 621
rect 3655 587 3671 621
rect 3605 521 3671 587
rect 3605 487 3621 521
rect 3655 487 3671 521
rect 3605 335 3671 487
rect 3707 596 3897 637
rect 3707 562 3800 596
rect 3834 562 3897 596
rect 3707 521 3897 562
rect 3707 487 3800 521
rect 3834 487 3897 521
rect 3707 471 3897 487
rect 3940 671 4007 687
rect 3940 637 3956 671
rect 3990 637 4007 671
rect 3940 596 4007 637
rect 3940 562 3956 596
rect 3990 562 4007 596
rect 3940 521 4007 562
rect 3940 487 3956 521
rect 3990 487 4007 521
rect 3940 471 4007 487
rect 3849 419 3915 435
rect 3849 385 3865 419
rect 3899 385 3915 419
rect 3849 351 3915 385
rect 3849 335 3865 351
rect 3605 317 3865 335
rect 3899 317 3915 351
rect 3605 301 3915 317
rect 3605 232 3671 301
rect 3961 265 4007 471
rect 3605 198 3621 232
rect 3655 198 3671 232
rect 3605 165 3671 198
rect 3707 249 3897 265
rect 3707 215 3800 249
rect 3834 215 3897 249
rect 3481 115 3497 149
rect 3531 115 3557 149
rect 3481 99 3557 115
rect 3707 149 3897 215
rect 3707 115 3800 149
rect 3834 115 3897 149
rect 3707 113 3897 115
rect 3248 73 3438 79
rect 3707 79 3713 113
rect 3747 79 3785 113
rect 3819 79 3857 113
rect 3891 79 3897 113
rect 3940 249 4007 265
rect 3940 215 3956 249
rect 3990 215 4007 249
rect 3940 149 4007 215
rect 3940 115 3956 149
rect 3990 115 4007 149
rect 3940 99 4007 115
rect 3707 73 3897 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 134 701 168 735
rect 206 701 240 735
rect 278 701 312 735
rect 683 701 717 735
rect 755 701 789 735
rect 827 711 861 735
rect 827 701 861 711
rect 139 79 173 113
rect 211 79 245 113
rect 283 79 317 113
rect 1139 701 1173 735
rect 1729 701 1763 735
rect 1801 701 1835 735
rect 1873 701 1907 735
rect 2197 719 2231 735
rect 2197 701 2214 719
rect 2214 701 2231 719
rect 2269 701 2303 735
rect 2341 701 2375 735
rect 774 79 808 113
rect 846 79 880 113
rect 918 79 952 113
rect 1080 79 1114 113
rect 1152 79 1186 113
rect 2706 701 2740 735
rect 2778 701 2812 735
rect 2850 701 2884 735
rect 3254 701 3288 735
rect 3326 731 3360 735
rect 3326 701 3351 731
rect 3351 701 3360 731
rect 3398 701 3432 735
rect 3713 701 3747 735
rect 3785 701 3819 735
rect 3857 701 3891 735
rect 1688 79 1722 113
rect 1760 79 1794 113
rect 1832 79 1866 113
rect 2115 79 2149 113
rect 2187 79 2221 113
rect 2259 79 2293 113
rect 2876 79 2910 113
rect 2948 79 2982 113
rect 3020 79 3054 113
rect 3254 79 3288 113
rect 3326 79 3360 113
rect 3398 79 3432 113
rect 3713 79 3747 113
rect 3785 79 3819 113
rect 3857 79 3891 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
<< metal1 >>
rect 0 831 4032 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 0 791 4032 797
rect 0 735 4032 763
rect 0 701 134 735
rect 168 701 206 735
rect 240 701 278 735
rect 312 701 683 735
rect 717 701 755 735
rect 789 701 827 735
rect 861 701 1139 735
rect 1173 701 1729 735
rect 1763 701 1801 735
rect 1835 701 1873 735
rect 1907 701 2197 735
rect 2231 701 2269 735
rect 2303 701 2341 735
rect 2375 701 2706 735
rect 2740 701 2778 735
rect 2812 701 2850 735
rect 2884 701 3254 735
rect 3288 701 3326 735
rect 3360 701 3398 735
rect 3432 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 4032 735
rect 0 689 4032 701
rect 0 113 4032 125
rect 0 79 139 113
rect 173 79 211 113
rect 245 79 283 113
rect 317 79 774 113
rect 808 79 846 113
rect 880 79 918 113
rect 952 79 1080 113
rect 1114 79 1152 113
rect 1186 79 1688 113
rect 1722 79 1760 113
rect 1794 79 1832 113
rect 1866 79 2115 113
rect 2149 79 2187 113
rect 2221 79 2259 113
rect 2293 79 2876 113
rect 2910 79 2948 113
rect 2982 79 3020 113
rect 3054 79 3254 113
rect 3288 79 3326 113
rect 3360 79 3398 113
rect 3432 79 3713 113
rect 3747 79 3785 113
rect 3819 79 3857 113
rect 3891 79 4032 113
rect 0 51 4032 79
rect 0 17 4032 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
rect 0 -23 4032 -17
<< labels >>
flabel comment s 1799 386 1799 386 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 1363 291 1363 291 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfsbp_1
flabel metal1 s 0 51 4032 125 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 0 4032 23 0 FreeSans 340 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 0 689 4032 763 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 791 4032 814 0 FreeSans 340 0 0 0 VPB
port 8 nsew power bidirectional
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 3967 168 4001 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 242 4001 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 316 4001 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 390 4001 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 464 4001 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 538 4001 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 612 4001 646 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3487 168 3521 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 242 3521 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 316 3521 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 390 3521 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 464 3521 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 538 3521 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 612 3521 646 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2143 242 2177 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
rlabel locali s 2109 73 2299 206 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 2870 73 3060 249 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 3248 73 3438 265 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 3707 73 3897 265 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 774 73 952 199 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 1074 73 1192 204 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 1682 73 1872 192 1 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 51 4032 125 1 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 4032 23 1 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 791 4032 837 1 VPB
port 8 nsew power bidirectional
rlabel locali s 2191 670 2381 751 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 2700 575 2890 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 3248 439 3438 747 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 3707 471 3897 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 683 561 861 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 1139 480 1173 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 1723 592 1913 741 1 VPWR
port 9 nsew power bidirectional
rlabel metal1 s 0 689 4032 763 1 VPWR
port 9 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 4032 814
string GDS_END 570340
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 531624
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
