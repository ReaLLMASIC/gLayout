magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1650 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 950 47 980 177
rect 1034 47 1064 177
rect 1118 47 1148 177
rect 1202 47 1232 177
rect 1286 47 1316 177
rect 1370 47 1400 177
rect 1454 47 1484 177
rect 1538 47 1568 177
<< scpmoshvt >>
rect 79 297 109 497
rect 174 309 204 497
rect 258 309 288 497
rect 342 309 372 497
rect 426 309 456 497
rect 510 309 540 497
rect 594 309 624 497
rect 678 309 708 497
rect 762 309 792 497
rect 950 297 980 497
rect 1034 297 1064 497
rect 1118 297 1148 497
rect 1202 297 1232 497
rect 1286 297 1316 497
rect 1370 297 1400 497
rect 1454 297 1484 497
rect 1538 297 1568 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 93 161 177
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 129 267 177
rect 215 95 223 129
rect 257 95 267 129
rect 215 47 267 95
rect 297 89 351 177
rect 297 55 307 89
rect 341 55 351 89
rect 297 47 351 55
rect 381 129 435 177
rect 381 95 391 129
rect 425 95 435 129
rect 381 47 435 95
rect 465 89 519 177
rect 465 55 475 89
rect 509 55 519 89
rect 465 47 519 55
rect 549 129 603 177
rect 549 95 559 129
rect 593 95 603 129
rect 549 47 603 95
rect 633 89 687 177
rect 633 55 643 89
rect 677 55 687 89
rect 633 47 687 55
rect 717 129 771 177
rect 717 95 727 129
rect 761 95 771 129
rect 717 47 771 95
rect 801 89 855 177
rect 801 55 811 89
rect 845 55 855 89
rect 801 47 855 55
rect 885 129 950 177
rect 885 95 901 129
rect 935 95 950 129
rect 885 47 950 95
rect 980 165 1034 177
rect 980 131 990 165
rect 1024 131 1034 165
rect 980 47 1034 131
rect 1064 90 1118 177
rect 1064 56 1074 90
rect 1108 56 1118 90
rect 1064 47 1118 56
rect 1148 165 1202 177
rect 1148 131 1158 165
rect 1192 131 1202 165
rect 1148 47 1202 131
rect 1232 90 1286 177
rect 1232 56 1242 90
rect 1276 56 1286 90
rect 1232 47 1286 56
rect 1316 165 1370 177
rect 1316 131 1326 165
rect 1360 131 1370 165
rect 1316 47 1370 131
rect 1400 90 1454 177
rect 1400 56 1410 90
rect 1444 56 1454 90
rect 1400 47 1454 56
rect 1484 165 1538 177
rect 1484 131 1494 165
rect 1528 131 1538 165
rect 1484 47 1538 131
rect 1568 90 1624 177
rect 1568 56 1578 90
rect 1612 56 1624 90
rect 1568 47 1624 56
<< pdiff >>
rect 27 448 79 497
rect 27 414 35 448
rect 69 414 79 448
rect 27 380 79 414
rect 27 346 35 380
rect 69 346 79 380
rect 27 297 79 346
rect 109 489 174 497
rect 109 455 119 489
rect 153 455 174 489
rect 109 421 174 455
rect 109 387 119 421
rect 153 387 174 421
rect 109 309 174 387
rect 204 448 258 497
rect 204 414 214 448
rect 248 414 258 448
rect 204 380 258 414
rect 204 346 214 380
rect 248 346 258 380
rect 204 309 258 346
rect 288 489 342 497
rect 288 455 298 489
rect 332 455 342 489
rect 288 421 342 455
rect 288 387 298 421
rect 332 387 342 421
rect 288 309 342 387
rect 372 448 426 497
rect 372 414 382 448
rect 416 414 426 448
rect 372 380 426 414
rect 372 346 382 380
rect 416 346 426 380
rect 372 309 426 346
rect 456 489 510 497
rect 456 455 466 489
rect 500 455 510 489
rect 456 421 510 455
rect 456 387 466 421
rect 500 387 510 421
rect 456 309 510 387
rect 540 448 594 497
rect 540 414 550 448
rect 584 414 594 448
rect 540 380 594 414
rect 540 346 550 380
rect 584 346 594 380
rect 540 309 594 346
rect 624 489 678 497
rect 624 455 634 489
rect 668 455 678 489
rect 624 421 678 455
rect 624 387 634 421
rect 668 387 678 421
rect 624 309 678 387
rect 708 448 762 497
rect 708 414 718 448
rect 752 414 762 448
rect 708 380 762 414
rect 708 346 718 380
rect 752 346 762 380
rect 708 309 762 346
rect 792 485 844 497
rect 792 451 802 485
rect 836 451 844 485
rect 792 417 844 451
rect 792 383 802 417
rect 836 383 844 417
rect 792 309 844 383
rect 898 448 950 497
rect 898 414 906 448
rect 940 414 950 448
rect 898 380 950 414
rect 898 346 906 380
rect 940 346 950 380
rect 109 297 159 309
rect 898 297 950 346
rect 980 425 1034 497
rect 980 391 990 425
rect 1024 391 1034 425
rect 980 357 1034 391
rect 980 323 990 357
rect 1024 323 1034 357
rect 980 297 1034 323
rect 1064 477 1118 497
rect 1064 443 1074 477
rect 1108 443 1118 477
rect 1064 409 1118 443
rect 1064 375 1074 409
rect 1108 375 1118 409
rect 1064 297 1118 375
rect 1148 425 1202 497
rect 1148 391 1158 425
rect 1192 391 1202 425
rect 1148 357 1202 391
rect 1148 323 1158 357
rect 1192 323 1202 357
rect 1148 297 1202 323
rect 1232 477 1286 497
rect 1232 443 1242 477
rect 1276 443 1286 477
rect 1232 409 1286 443
rect 1232 375 1242 409
rect 1276 375 1286 409
rect 1232 297 1286 375
rect 1316 425 1370 497
rect 1316 391 1326 425
rect 1360 391 1370 425
rect 1316 357 1370 391
rect 1316 323 1326 357
rect 1360 323 1370 357
rect 1316 297 1370 323
rect 1400 477 1454 497
rect 1400 443 1410 477
rect 1444 443 1454 477
rect 1400 409 1454 443
rect 1400 375 1410 409
rect 1444 375 1454 409
rect 1400 297 1454 375
rect 1484 425 1538 497
rect 1484 391 1494 425
rect 1528 391 1538 425
rect 1484 357 1538 391
rect 1484 323 1494 357
rect 1528 323 1538 357
rect 1484 297 1538 323
rect 1568 477 1620 497
rect 1568 443 1578 477
rect 1612 443 1620 477
rect 1568 409 1620 443
rect 1568 375 1578 409
rect 1612 375 1620 409
rect 1568 297 1620 375
<< ndiffc >>
rect 35 95 69 129
rect 119 59 153 93
rect 223 95 257 129
rect 307 55 341 89
rect 391 95 425 129
rect 475 55 509 89
rect 559 95 593 129
rect 643 55 677 89
rect 727 95 761 129
rect 811 55 845 89
rect 901 95 935 129
rect 990 131 1024 165
rect 1074 56 1108 90
rect 1158 131 1192 165
rect 1242 56 1276 90
rect 1326 131 1360 165
rect 1410 56 1444 90
rect 1494 131 1528 165
rect 1578 56 1612 90
<< pdiffc >>
rect 35 414 69 448
rect 35 346 69 380
rect 119 455 153 489
rect 119 387 153 421
rect 214 414 248 448
rect 214 346 248 380
rect 298 455 332 489
rect 298 387 332 421
rect 382 414 416 448
rect 382 346 416 380
rect 466 455 500 489
rect 466 387 500 421
rect 550 414 584 448
rect 550 346 584 380
rect 634 455 668 489
rect 634 387 668 421
rect 718 414 752 448
rect 718 346 752 380
rect 802 451 836 485
rect 802 383 836 417
rect 906 414 940 448
rect 906 346 940 380
rect 990 391 1024 425
rect 990 323 1024 357
rect 1074 443 1108 477
rect 1074 375 1108 409
rect 1158 391 1192 425
rect 1158 323 1192 357
rect 1242 443 1276 477
rect 1242 375 1276 409
rect 1326 391 1360 425
rect 1326 323 1360 357
rect 1410 443 1444 477
rect 1410 375 1444 409
rect 1494 391 1528 425
rect 1494 323 1528 357
rect 1578 443 1612 477
rect 1578 375 1612 409
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 258 497 288 523
rect 342 497 372 523
rect 426 497 456 523
rect 510 497 540 523
rect 594 497 624 523
rect 678 497 708 523
rect 762 497 792 523
rect 950 497 980 523
rect 1034 497 1064 523
rect 1118 497 1148 523
rect 1202 497 1232 523
rect 1286 497 1316 523
rect 1370 497 1400 523
rect 1454 497 1484 523
rect 1538 497 1568 523
rect 79 265 109 297
rect 174 294 204 309
rect 258 294 288 309
rect 342 294 372 309
rect 426 294 456 309
rect 510 294 540 309
rect 594 294 624 309
rect 678 294 708 309
rect 762 294 792 309
rect 174 265 792 294
rect 950 265 980 297
rect 1034 265 1064 297
rect 1118 265 1148 297
rect 1202 265 1232 297
rect 1286 265 1316 297
rect 1370 265 1400 297
rect 1454 265 1484 297
rect 1538 265 1568 297
rect 22 264 792 265
rect 22 249 204 264
rect 22 215 32 249
rect 66 235 204 249
rect 834 249 888 265
rect 66 215 109 235
rect 834 222 844 249
rect 22 199 109 215
rect 79 177 109 199
rect 267 215 844 222
rect 878 215 888 249
rect 267 199 888 215
rect 950 249 1568 265
rect 950 215 966 249
rect 1000 215 1034 249
rect 1068 215 1102 249
rect 1136 215 1170 249
rect 1204 215 1238 249
rect 1272 215 1306 249
rect 1340 215 1374 249
rect 1408 215 1442 249
rect 1476 215 1510 249
rect 1544 215 1568 249
rect 950 199 1568 215
rect 267 192 885 199
rect 267 177 297 192
rect 351 177 381 192
rect 435 177 465 192
rect 519 177 549 192
rect 603 177 633 192
rect 687 177 717 192
rect 771 177 801 192
rect 855 177 885 192
rect 950 177 980 199
rect 1034 177 1064 199
rect 1118 177 1148 199
rect 1202 177 1232 199
rect 1286 177 1316 199
rect 1370 177 1400 199
rect 1454 177 1484 199
rect 1538 177 1568 199
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 950 21 980 47
rect 1034 21 1064 47
rect 1118 21 1148 47
rect 1202 21 1232 47
rect 1286 21 1316 47
rect 1370 21 1400 47
rect 1454 21 1484 47
rect 1538 21 1568 47
<< polycont >>
rect 32 215 66 249
rect 844 215 878 249
rect 966 215 1000 249
rect 1034 215 1068 249
rect 1102 215 1136 249
rect 1170 215 1204 249
rect 1238 215 1272 249
rect 1306 215 1340 249
rect 1374 215 1408 249
rect 1442 215 1476 249
rect 1510 215 1544 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 18 448 69 493
rect 18 414 35 448
rect 18 380 69 414
rect 18 346 35 380
rect 103 489 169 527
rect 103 455 119 489
rect 153 455 169 489
rect 103 421 169 455
rect 103 387 119 421
rect 153 387 169 421
rect 103 367 169 387
rect 203 448 248 493
rect 203 414 214 448
rect 203 380 248 414
rect 18 333 69 346
rect 203 346 214 380
rect 282 489 348 527
rect 282 455 298 489
rect 332 455 348 489
rect 282 421 348 455
rect 282 387 298 421
rect 332 387 348 421
rect 282 367 348 387
rect 382 448 416 493
rect 382 380 416 414
rect 203 333 248 346
rect 450 489 516 527
rect 450 455 466 489
rect 500 455 516 489
rect 450 421 516 455
rect 450 387 466 421
rect 500 387 516 421
rect 450 367 516 387
rect 550 448 584 493
rect 550 380 584 414
rect 382 333 416 346
rect 618 489 684 527
rect 618 455 634 489
rect 668 455 684 489
rect 618 421 684 455
rect 618 387 634 421
rect 668 387 684 421
rect 618 367 684 387
rect 718 448 752 493
rect 718 380 752 414
rect 550 333 584 346
rect 786 485 856 527
rect 786 451 802 485
rect 836 451 856 485
rect 786 417 856 451
rect 786 383 802 417
rect 836 383 856 417
rect 786 367 856 383
rect 890 477 1639 493
rect 890 459 1074 477
rect 890 448 940 459
rect 890 414 906 448
rect 1108 459 1242 477
rect 890 380 940 414
rect 718 333 752 346
rect 890 346 906 380
rect 890 333 940 346
rect 18 299 169 333
rect 203 299 940 333
rect 974 391 990 425
rect 1024 391 1040 425
rect 974 357 1040 391
rect 1074 409 1108 443
rect 1276 459 1410 477
rect 1074 359 1108 375
rect 1142 391 1158 425
rect 1192 391 1208 425
rect 974 323 990 357
rect 1024 325 1040 357
rect 1142 357 1208 391
rect 1242 409 1276 443
rect 1444 459 1578 477
rect 1242 359 1276 375
rect 1310 391 1326 425
rect 1360 391 1376 425
rect 1142 325 1158 357
rect 1024 323 1158 325
rect 1192 325 1208 357
rect 1310 357 1376 391
rect 1410 409 1444 443
rect 1612 443 1639 477
rect 1410 359 1444 375
rect 1478 391 1494 425
rect 1528 391 1544 425
rect 1310 325 1326 357
rect 1192 323 1326 325
rect 1360 325 1376 357
rect 1478 357 1544 391
rect 1578 409 1639 443
rect 1612 375 1639 409
rect 1578 359 1639 375
rect 1478 325 1494 357
rect 1360 323 1494 325
rect 1528 325 1544 357
rect 1528 323 1639 325
rect 103 265 169 299
rect 974 291 1639 323
rect 18 249 69 265
rect 18 215 32 249
rect 66 215 69 249
rect 18 199 69 215
rect 103 249 895 265
rect 103 215 844 249
rect 878 215 895 249
rect 103 199 895 215
rect 929 249 1560 257
rect 929 215 966 249
rect 1000 215 1034 249
rect 1068 215 1102 249
rect 1136 215 1170 249
rect 1204 215 1238 249
rect 1272 215 1306 249
rect 1340 215 1374 249
rect 1408 215 1442 249
rect 1476 215 1510 249
rect 1544 215 1560 249
rect 929 199 1560 215
rect 103 165 169 199
rect 1594 165 1639 291
rect 18 131 169 165
rect 203 131 940 165
rect 18 129 69 131
rect 18 95 35 129
rect 203 129 257 131
rect 18 51 69 95
rect 103 93 169 97
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 203 95 223 129
rect 391 129 425 131
rect 203 51 257 95
rect 291 89 357 97
rect 291 55 307 89
rect 341 55 357 89
rect 291 17 357 55
rect 559 129 593 131
rect 391 51 425 95
rect 459 89 525 97
rect 459 55 475 89
rect 509 55 525 89
rect 459 17 525 55
rect 727 129 761 131
rect 559 51 593 95
rect 627 89 693 97
rect 627 55 643 89
rect 677 55 693 89
rect 627 17 693 55
rect 897 129 940 131
rect 727 51 761 95
rect 795 89 863 97
rect 795 55 811 89
rect 845 55 863 89
rect 795 17 863 55
rect 897 95 901 129
rect 935 95 940 129
rect 974 131 990 165
rect 1024 131 1158 165
rect 1192 131 1326 165
rect 1360 131 1494 165
rect 1528 131 1639 165
rect 974 124 1639 131
rect 897 90 940 95
rect 897 56 1074 90
rect 1108 56 1242 90
rect 1276 56 1410 90
rect 1444 56 1578 90
rect 1612 56 1639 90
rect 897 51 1639 56
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 1318 221 1352 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1410 221 1444 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1502 221 1536 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1318 357 1352 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1502 357 1536 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1594 153 1628 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1594 221 1628 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 950 221 984 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1134 221 1168 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1226 221 1260 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 einvn_8
rlabel metal1 s 0 -48 1656 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 3027444
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3015180
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 41.400 0.000 
<< end >>
