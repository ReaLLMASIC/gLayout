magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< obsli1 >>
rect 81 96 8535 39476
<< metal1 >>
rect 7727 0 7877 3360
<< obsm1 >>
rect 75 3416 8573 39482
rect 75 62 7671 3416
rect 7933 62 8573 3416
<< obsm2 >>
rect 1938 430 8573 38730
<< metal3 >>
rect 2724 0 5308 1880
rect 5608 0 8218 925
<< obsm3 >>
rect 2724 1960 8218 38735
rect 5388 1005 8218 1960
rect 5388 925 5528 1005
<< labels >>
rlabel metal1 s 7727 0 7877 3360 6 ogc_lvc
port 1 nsew power bidirectional
rlabel metal3 s 2724 0 5308 1880 6 drn_lvc
port 2 nsew power bidirectional
rlabel metal3 s 5608 0 8218 925 6 src_bdy_lvc
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 9579 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 6061972
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2770452
<< end >>
