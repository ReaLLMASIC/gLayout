magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -116 -66 236 1066
<< mvpmos >>
rect 0 0 120 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 120 0 170 1000
<< poly >>
rect 0 1000 120 1032
rect 0 -32 120 0
<< labels >>
flabel comment s -25 500 -25 500 0 FreeSans 300 0 0 0 S
flabel comment s 145 500 145 500 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 12842656
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 12841888
<< end >>
