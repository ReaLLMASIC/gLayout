magic
tech sky130A
timestamp 1701704242
<< metal1 >>
rect 0 0 3 890
rect 285 0 288 890
<< via1 >>
rect 3 0 285 890
<< metal2 >>
rect 0 0 3 890
rect 285 0 288 890
<< properties >>
string GDS_END 93651438
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93635178
<< end >>
