magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 98 157 717 203
rect 1 67 717 157
rect 1 21 191 67
rect 405 21 717 67
rect 30 -17 64 21
<< locali >>
rect 17 199 71 323
rect 182 215 248 326
rect 395 299 719 493
rect 651 165 719 299
rect 625 51 719 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 401 69 493
rect 103 435 169 527
rect 203 401 254 492
rect 288 435 361 527
rect 17 357 148 401
rect 203 360 361 401
rect 105 165 148 357
rect 282 265 361 360
rect 282 215 507 265
rect 282 177 337 215
rect 541 199 617 265
rect 541 181 591 199
rect 17 123 237 165
rect 271 127 337 177
rect 371 147 591 181
rect 17 56 69 123
rect 203 93 237 123
rect 371 93 405 147
rect 103 17 169 89
rect 203 51 405 93
rect 439 17 591 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 17 199 71 323 6 A
port 1 nsew signal input
rlabel locali s 182 215 248 326 6 TE_B
port 2 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 405 21 717 67 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 191 67 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 67 717 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 98 157 717 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 625 51 719 165 6 Z
port 7 nsew signal output
rlabel locali s 651 165 719 299 6 Z
port 7 nsew signal output
rlabel locali s 395 299 719 493 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2924272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2917454
<< end >>
