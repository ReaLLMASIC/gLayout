magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 23 201 1617 203
rect 23 23 1928 201
rect 23 21 473 23
rect 931 21 1121 23
rect 1532 21 1928 23
rect 29 -17 63 21
<< scnmos >>
rect 101 47 131 177
rect 185 47 215 177
rect 271 47 301 177
rect 355 47 385 177
rect 462 93 492 177
rect 685 49 715 177
rect 773 49 803 177
rect 1015 47 1045 177
rect 1201 49 1231 177
rect 1352 49 1382 133
rect 1511 49 1541 177
rect 1631 47 1661 167
rect 1731 47 1761 175
rect 1815 47 1845 175
<< scpmoshvt >>
rect 101 297 131 497
rect 185 297 215 497
rect 275 297 305 497
rect 359 297 389 497
rect 462 297 492 425
rect 672 325 702 493
rect 769 297 799 465
rect 981 297 1011 497
rect 1201 297 1231 465
rect 1352 297 1382 425
rect 1527 329 1557 457
rect 1630 329 1660 497
rect 1731 297 1761 497
rect 1815 297 1845 497
<< ndiff >>
rect 49 129 101 177
rect 49 95 57 129
rect 91 95 101 129
rect 49 47 101 95
rect 131 129 185 177
rect 131 95 141 129
rect 175 95 185 129
rect 131 47 185 95
rect 215 129 271 177
rect 215 95 225 129
rect 259 95 271 129
rect 215 47 271 95
rect 301 129 355 177
rect 301 95 311 129
rect 345 95 355 129
rect 301 47 355 95
rect 385 93 462 177
rect 492 169 577 177
rect 492 135 531 169
rect 565 135 577 169
rect 492 93 577 135
rect 631 165 685 177
rect 631 131 641 165
rect 675 131 685 165
rect 385 89 447 93
rect 385 55 395 89
rect 429 55 447 89
rect 385 47 447 55
rect 631 49 685 131
rect 715 91 773 177
rect 715 57 727 91
rect 761 57 773 91
rect 715 49 773 57
rect 803 91 873 177
rect 803 57 827 91
rect 861 57 873 91
rect 803 49 873 57
rect 957 157 1015 177
rect 957 123 971 157
rect 1005 123 1015 157
rect 957 89 1015 123
rect 957 55 971 89
rect 1005 55 1015 89
rect 957 47 1015 55
rect 1045 165 1097 177
rect 1045 131 1055 165
rect 1089 131 1097 165
rect 1045 124 1097 131
rect 1045 47 1095 124
rect 1151 104 1201 177
rect 1149 97 1201 104
rect 1149 63 1157 97
rect 1191 63 1201 97
rect 1149 49 1201 63
rect 1231 133 1331 177
rect 1407 169 1511 177
rect 1407 135 1453 169
rect 1487 135 1511 169
rect 1407 133 1511 135
rect 1231 126 1352 133
rect 1231 92 1241 126
rect 1275 92 1352 126
rect 1231 49 1352 92
rect 1382 49 1511 133
rect 1541 167 1591 177
rect 1681 167 1731 175
rect 1541 93 1631 167
rect 1541 59 1553 93
rect 1587 59 1631 93
rect 1541 49 1631 59
rect 1558 47 1631 49
rect 1661 142 1731 167
rect 1661 108 1687 142
rect 1721 108 1731 142
rect 1661 47 1731 108
rect 1761 97 1815 175
rect 1761 63 1771 97
rect 1805 63 1815 97
rect 1761 47 1815 63
rect 1845 101 1902 175
rect 1845 67 1855 101
rect 1889 67 1902 101
rect 1845 47 1902 67
<< pdiff >>
rect 49 485 101 497
rect 49 451 57 485
rect 91 451 101 485
rect 49 417 101 451
rect 49 383 57 417
rect 91 383 101 417
rect 49 349 101 383
rect 49 315 57 349
rect 91 315 101 349
rect 49 297 101 315
rect 131 485 185 497
rect 131 451 141 485
rect 175 451 185 485
rect 131 417 185 451
rect 131 383 141 417
rect 175 383 185 417
rect 131 349 185 383
rect 131 315 141 349
rect 175 315 185 349
rect 131 297 185 315
rect 215 485 275 497
rect 215 451 225 485
rect 259 451 275 485
rect 215 417 275 451
rect 215 383 225 417
rect 259 383 275 417
rect 215 349 275 383
rect 215 315 225 349
rect 259 315 275 349
rect 215 297 275 315
rect 305 477 359 497
rect 305 443 315 477
rect 349 443 359 477
rect 305 409 359 443
rect 305 375 315 409
rect 349 375 359 409
rect 305 341 359 375
rect 305 307 315 341
rect 349 307 359 341
rect 305 297 359 307
rect 389 477 447 497
rect 389 443 400 477
rect 434 443 447 477
rect 389 425 447 443
rect 389 297 462 425
rect 492 341 548 425
rect 492 307 502 341
rect 536 307 548 341
rect 607 413 672 493
rect 607 379 628 413
rect 662 379 672 413
rect 607 325 672 379
rect 702 481 754 493
rect 702 447 712 481
rect 746 465 754 481
rect 929 481 981 497
rect 746 447 769 465
rect 702 325 769 447
rect 492 297 548 307
rect 719 297 769 325
rect 799 423 875 465
rect 929 447 937 481
rect 971 447 981 481
rect 929 435 981 447
rect 799 339 876 423
rect 799 305 830 339
rect 864 305 876 339
rect 799 297 876 305
rect 930 297 981 435
rect 1011 343 1063 497
rect 1011 309 1021 343
rect 1055 309 1063 343
rect 1011 297 1063 309
rect 1117 405 1201 465
rect 1117 371 1125 405
rect 1159 371 1201 405
rect 1117 297 1201 371
rect 1231 425 1330 465
rect 1572 489 1630 497
rect 1572 457 1584 489
rect 1442 425 1527 457
rect 1231 409 1352 425
rect 1231 375 1281 409
rect 1315 375 1352 409
rect 1231 341 1352 375
rect 1231 307 1281 341
rect 1315 307 1352 341
rect 1231 297 1352 307
rect 1382 421 1527 425
rect 1382 387 1483 421
rect 1517 387 1527 421
rect 1382 329 1527 387
rect 1557 455 1584 457
rect 1618 455 1630 489
rect 1557 329 1630 455
rect 1660 341 1731 497
rect 1660 329 1687 341
rect 1382 297 1477 329
rect 1675 307 1687 329
rect 1721 307 1731 341
rect 1675 297 1731 307
rect 1761 489 1815 497
rect 1761 455 1771 489
rect 1805 455 1815 489
rect 1761 297 1815 455
rect 1845 477 1902 497
rect 1845 443 1856 477
rect 1890 443 1902 477
rect 1845 409 1902 443
rect 1845 375 1856 409
rect 1890 375 1902 409
rect 1845 297 1902 375
<< ndiffc >>
rect 57 95 91 129
rect 141 95 175 129
rect 225 95 259 129
rect 311 95 345 129
rect 531 135 565 169
rect 641 131 675 165
rect 395 55 429 89
rect 727 57 761 91
rect 827 57 861 91
rect 971 123 1005 157
rect 971 55 1005 89
rect 1055 131 1089 165
rect 1157 63 1191 97
rect 1453 135 1487 169
rect 1241 92 1275 126
rect 1553 59 1587 93
rect 1687 108 1721 142
rect 1771 63 1805 97
rect 1855 67 1889 101
<< pdiffc >>
rect 57 451 91 485
rect 57 383 91 417
rect 57 315 91 349
rect 141 451 175 485
rect 141 383 175 417
rect 141 315 175 349
rect 225 451 259 485
rect 225 383 259 417
rect 225 315 259 349
rect 315 443 349 477
rect 315 375 349 409
rect 315 307 349 341
rect 400 443 434 477
rect 502 307 536 341
rect 628 379 662 413
rect 712 447 746 481
rect 937 447 971 481
rect 830 305 864 339
rect 1021 309 1055 343
rect 1125 371 1159 405
rect 1281 375 1315 409
rect 1281 307 1315 341
rect 1483 387 1517 421
rect 1584 455 1618 489
rect 1687 307 1721 341
rect 1771 455 1805 489
rect 1856 443 1890 477
rect 1856 375 1890 409
<< poly >>
rect 101 497 131 523
rect 185 497 215 523
rect 275 497 305 523
rect 359 497 389 523
rect 672 493 702 519
rect 462 425 492 483
rect 769 465 799 504
rect 981 497 1011 523
rect 101 265 131 297
rect 185 265 215 297
rect 275 265 305 297
rect 359 265 389 297
rect 462 265 492 297
rect 672 271 702 325
rect 1201 493 1557 523
rect 1630 497 1660 523
rect 1731 497 1761 523
rect 1815 497 1845 523
rect 1201 465 1231 493
rect 1527 457 1557 493
rect 1352 425 1382 451
rect 672 265 715 271
rect 769 265 799 297
rect 101 249 420 265
rect 101 215 376 249
rect 410 215 420 249
rect 101 199 420 215
rect 462 249 715 265
rect 462 215 642 249
rect 676 215 715 249
rect 462 199 715 215
rect 757 249 811 265
rect 757 215 767 249
rect 801 215 811 249
rect 981 247 1011 297
rect 1201 247 1231 297
rect 1352 265 1382 297
rect 1527 265 1557 329
rect 981 217 1231 247
rect 757 199 811 215
rect 101 177 131 199
rect 185 177 215 199
rect 271 177 301 199
rect 355 177 385 199
rect 462 177 492 199
rect 685 177 715 199
rect 773 177 803 199
rect 1015 177 1045 217
rect 1201 177 1231 217
rect 1273 249 1382 265
rect 1273 215 1283 249
rect 1317 215 1382 249
rect 1273 199 1382 215
rect 462 67 492 93
rect 101 21 131 47
rect 185 21 215 47
rect 271 21 301 47
rect 355 21 385 47
rect 685 21 715 49
rect 773 21 803 49
rect 1352 133 1382 199
rect 1511 249 1565 265
rect 1630 256 1660 329
rect 1731 265 1761 297
rect 1815 265 1845 297
rect 1630 255 1661 256
rect 1511 215 1521 249
rect 1555 215 1565 249
rect 1511 199 1565 215
rect 1607 239 1661 255
rect 1607 205 1617 239
rect 1651 205 1661 239
rect 1511 177 1541 199
rect 1607 189 1661 205
rect 1703 249 1761 265
rect 1703 215 1713 249
rect 1747 215 1761 249
rect 1703 199 1761 215
rect 1803 249 1857 265
rect 1803 215 1813 249
rect 1847 215 1857 249
rect 1803 199 1857 215
rect 1631 167 1661 189
rect 1731 175 1761 199
rect 1815 175 1845 199
rect 1015 21 1045 47
rect 1201 21 1231 49
rect 1352 23 1382 49
rect 1511 21 1541 49
rect 1631 21 1661 47
rect 1731 21 1761 47
rect 1815 21 1845 47
<< polycont >>
rect 376 215 410 249
rect 642 215 676 249
rect 767 215 801 249
rect 1283 215 1317 249
rect 1521 215 1555 249
rect 1617 205 1651 239
rect 1713 215 1747 249
rect 1813 215 1847 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 57 485 91 527
rect 225 485 259 527
rect 57 417 91 451
rect 57 349 91 383
rect 57 298 91 315
rect 125 451 141 485
rect 175 451 191 485
rect 125 417 191 451
rect 125 383 141 417
rect 175 383 191 417
rect 125 349 191 383
rect 125 315 141 349
rect 175 315 191 349
rect 125 265 191 315
rect 225 417 259 451
rect 225 349 259 383
rect 225 299 259 315
rect 293 477 349 493
rect 293 443 315 477
rect 383 477 450 527
rect 921 481 987 527
rect 1755 489 1822 527
rect 383 443 400 477
rect 434 443 450 477
rect 486 447 712 481
rect 746 447 780 481
rect 921 447 937 481
rect 971 447 987 481
rect 1054 455 1584 489
rect 1618 455 1673 489
rect 1755 455 1771 489
rect 1805 455 1822 489
rect 1856 477 1915 493
rect 293 409 349 443
rect 486 409 520 447
rect 1054 413 1088 455
rect 293 375 315 409
rect 293 341 349 375
rect 293 307 315 341
rect 293 288 349 307
rect 383 375 520 409
rect 588 379 628 413
rect 662 379 1088 413
rect 1125 405 1159 421
rect 293 265 342 288
rect 383 265 417 375
rect 463 307 502 341
rect 536 307 780 341
rect 125 199 342 265
rect 376 249 417 265
rect 410 215 417 249
rect 376 199 417 215
rect 57 129 91 147
rect 57 17 91 95
rect 125 129 175 199
rect 293 185 342 199
rect 125 95 141 129
rect 125 75 175 95
rect 225 129 259 147
rect 225 17 259 95
rect 293 129 345 185
rect 382 173 417 199
rect 382 139 497 173
rect 293 95 311 129
rect 293 70 345 95
rect 379 89 429 105
rect 379 55 395 89
rect 379 17 429 55
rect 463 85 497 139
rect 531 169 565 307
rect 746 265 780 307
rect 814 305 830 339
rect 864 323 891 339
rect 835 289 857 305
rect 835 275 891 289
rect 599 249 712 265
rect 599 215 642 249
rect 676 215 712 249
rect 746 249 801 265
rect 746 215 767 249
rect 746 199 801 215
rect 531 119 565 135
rect 625 165 701 181
rect 625 131 641 165
rect 675 159 701 165
rect 835 159 869 275
rect 925 241 959 379
rect 1005 309 1021 343
rect 1055 309 1089 343
rect 1005 289 1089 309
rect 675 131 869 159
rect 625 125 869 131
rect 903 207 959 241
rect 903 91 937 207
rect 1041 187 1089 289
rect 690 85 727 91
rect 463 57 727 85
rect 761 57 777 91
rect 811 57 827 91
rect 861 57 937 91
rect 971 157 1005 173
rect 971 89 1005 123
rect 463 51 777 57
rect 1075 165 1089 187
rect 1041 131 1055 153
rect 1041 83 1089 131
rect 1125 119 1159 371
rect 1193 178 1227 455
rect 1890 443 1915 477
rect 1856 421 1915 443
rect 1263 375 1281 409
rect 1315 375 1346 409
rect 1263 341 1346 375
rect 1263 307 1281 341
rect 1315 323 1346 341
rect 1453 387 1483 421
rect 1517 409 1915 421
rect 1517 387 1856 409
rect 1315 307 1317 323
rect 1263 289 1317 307
rect 1351 289 1419 323
rect 1266 249 1351 254
rect 1266 215 1283 249
rect 1317 215 1351 249
rect 1266 199 1351 215
rect 1309 187 1351 199
rect 1193 165 1235 178
rect 1193 144 1275 165
rect 1201 131 1275 144
rect 1241 126 1275 131
rect 1309 153 1317 187
rect 1309 126 1351 153
rect 1125 85 1133 119
rect 971 17 1005 55
rect 1125 63 1157 85
rect 1191 63 1207 97
rect 1241 64 1275 92
rect 1385 85 1419 289
rect 1453 169 1487 387
rect 1818 375 1856 387
rect 1890 375 1915 409
rect 1521 289 1637 323
rect 1671 307 1687 341
rect 1721 307 1835 341
rect 1671 299 1835 307
rect 1521 249 1555 289
rect 1801 265 1835 299
rect 1521 199 1555 215
rect 1589 239 1651 255
rect 1589 205 1617 239
rect 1685 249 1767 265
rect 1685 215 1713 249
rect 1747 215 1767 249
rect 1801 249 1847 265
rect 1801 215 1813 249
rect 1589 189 1651 205
rect 1801 199 1847 215
rect 1589 187 1630 189
rect 1589 153 1593 187
rect 1627 153 1630 187
rect 1801 181 1835 199
rect 1589 146 1630 153
rect 1687 150 1835 181
rect 1679 147 1835 150
rect 1453 119 1487 135
rect 1679 142 1737 147
rect 1679 119 1687 142
rect 1521 85 1553 93
rect 1125 53 1207 63
rect 1385 59 1553 85
rect 1587 59 1614 93
rect 1679 85 1685 119
rect 1721 108 1737 142
rect 1881 117 1915 375
rect 1719 85 1737 108
rect 1679 59 1737 85
rect 1771 97 1805 113
rect 1385 51 1614 59
rect 1771 17 1805 63
rect 1855 101 1915 117
rect 1889 67 1915 101
rect 1855 51 1915 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 857 305 864 323
rect 864 305 891 323
rect 857 289 891 305
rect 1041 165 1075 187
rect 1041 153 1055 165
rect 1055 153 1075 165
rect 1317 289 1351 323
rect 1317 153 1351 187
rect 1133 97 1167 119
rect 1133 85 1157 97
rect 1157 85 1167 97
rect 1593 153 1627 187
rect 1685 108 1687 119
rect 1687 108 1719 119
rect 1685 85 1719 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 845 323 903 329
rect 845 289 857 323
rect 891 320 903 323
rect 1305 323 1363 329
rect 1305 320 1317 323
rect 891 292 1317 320
rect 891 289 903 292
rect 845 283 903 289
rect 1305 289 1317 292
rect 1351 289 1363 323
rect 1305 283 1363 289
rect 1029 187 1087 193
rect 1029 153 1041 187
rect 1075 184 1087 187
rect 1305 187 1363 193
rect 1305 184 1317 187
rect 1075 156 1317 184
rect 1075 153 1087 156
rect 1029 147 1087 153
rect 1305 153 1317 156
rect 1351 184 1363 187
rect 1581 187 1639 193
rect 1581 184 1593 187
rect 1351 156 1593 184
rect 1351 153 1363 156
rect 1305 147 1363 153
rect 1581 153 1593 156
rect 1627 153 1639 187
rect 1581 147 1639 153
rect 1121 119 1179 125
rect 1121 85 1133 119
rect 1167 116 1179 119
rect 1673 119 1731 125
rect 1673 116 1685 119
rect 1167 88 1685 116
rect 1167 85 1179 88
rect 1121 79 1179 85
rect 1673 85 1685 88
rect 1719 85 1731 119
rect 1673 79 1731 85
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 305 357 339 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1593 289 1627 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1685 221 1719 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 hkscl5hdv1_xnor3_1
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
rlabel metal1 s 0 -48 1932 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 580264
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 567078
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.660 0.000 
<< end >>
