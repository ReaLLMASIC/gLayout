magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 495 226
<< mvnnmos >>
rect 0 0 180 200
rect 236 0 416 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 180 182 236 200
rect 180 148 191 182
rect 225 148 236 182
rect 180 114 236 148
rect 180 80 191 114
rect 225 80 236 114
rect 180 46 236 80
rect 180 12 191 46
rect 225 12 236 46
rect 180 0 236 12
rect 416 182 469 200
rect 416 148 427 182
rect 461 148 469 182
rect 416 114 469 148
rect 416 80 427 114
rect 461 80 469 114
rect 416 46 469 80
rect 416 12 427 46
rect 461 12 469 46
rect 416 0 469 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 191 148 225 182
rect 191 80 225 114
rect 191 12 225 46
rect 427 148 461 182
rect 427 80 461 114
rect 427 12 461 46
<< poly >>
rect 0 200 180 226
rect 236 200 416 226
rect 0 -26 180 0
rect 236 -26 416 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 191 182 225 198
rect 191 114 225 148
rect 191 46 225 80
rect 191 -4 225 12
rect 427 182 461 198
rect 427 114 461 148
rect 427 46 461 80
rect 427 -4 461 12
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_1
timestamp 1701704242
transform 1 0 416 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1701704242
transform 1 0 180 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 208 97 208 97 0 FreeSans 300 0 0 0 D
flabel comment s 444 97 444 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 96485764
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96484314
<< end >>
