magic
tech sky130A
timestamp 1701704242
<< metal1 >>
rect 0 0 3 154
rect 93 0 96 154
<< via1 >>
rect 3 0 93 154
<< metal2 >>
rect 0 0 3 154
rect 93 0 96 154
<< properties >>
string GDS_END 85424904
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85423812
<< end >>
