magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< poly >>
rect 277 9434 464 9467
rect 277 9400 294 9434
rect 328 9400 362 9434
rect 396 9400 430 9434
rect 277 9367 464 9400
rect 2504 9434 2691 9467
rect 2538 9400 2572 9434
rect 2606 9400 2640 9434
rect 2674 9400 2691 9434
rect 2504 9367 2691 9400
<< polycont >>
rect 294 9400 328 9434
rect 362 9400 396 9434
rect 430 9400 464 9434
rect 2504 9400 2538 9434
rect 2572 9400 2606 9434
rect 2640 9400 2674 9434
<< npolyres >>
rect 464 9367 2504 9467
<< locali >>
rect 2486 9450 2689 9508
rect 278 9440 480 9450
rect 2486 9440 2690 9450
rect 278 9434 481 9440
rect 278 9400 291 9434
rect 328 9400 362 9434
rect 397 9400 430 9434
rect 469 9400 481 9434
rect 278 9394 481 9400
rect 2487 9434 2690 9440
rect 2487 9400 2499 9434
rect 2538 9400 2571 9434
rect 2606 9400 2640 9434
rect 2677 9400 2690 9434
rect 2487 9394 2690 9400
rect 278 9384 480 9394
rect 2488 9384 2690 9394
rect 688 3623 702 7261
rect 14252 3623 14266 7261
<< viali >>
rect 291 9400 294 9434
rect 294 9400 325 9434
rect 363 9400 396 9434
rect 396 9400 397 9434
rect 435 9400 464 9434
rect 464 9400 469 9434
rect 2499 9400 2504 9434
rect 2504 9400 2533 9434
rect 2571 9400 2572 9434
rect 2572 9400 2605 9434
rect 2643 9400 2674 9434
rect 2674 9400 2677 9434
<< metal1 >>
rect 2487 9476 2690 9492
rect 278 9434 357 9446
rect 278 9400 291 9434
rect 325 9400 357 9434
rect 278 9394 357 9400
rect 409 9394 421 9446
rect 473 9394 481 9446
rect 2427 9434 2690 9476
rect 2427 9424 2499 9434
rect 2487 9400 2499 9424
rect 2533 9400 2571 9434
rect 2605 9400 2643 9434
rect 2677 9400 2690 9434
rect 2487 9362 2690 9400
rect 915 4028 1705 4033
rect 785 4021 1705 4028
rect 785 3969 791 4021
rect 843 3969 857 4021
rect 909 3969 1705 4021
rect 785 3957 1705 3969
rect 785 3905 791 3957
rect 843 3905 857 3957
rect 909 3905 1705 3957
rect 785 3903 1705 3905
rect 2135 3981 2141 4033
rect 2193 3981 2207 4033
rect 2259 3981 2265 4033
rect 2135 3955 2265 3981
rect 2135 3903 2141 3955
rect 2193 3903 2207 3955
rect 2259 3903 2265 3955
rect 2697 4026 2827 4033
rect 2697 3974 2703 4026
rect 2755 3974 2769 4026
rect 2821 3974 2827 4026
rect 2697 3962 2827 3974
rect 2697 3910 2703 3962
rect 2755 3910 2769 3962
rect 2821 3910 2827 3962
rect 2697 3903 2827 3910
rect 3257 3903 3757 4033
rect 3810 4026 4189 4033
rect 3810 3974 3816 4026
rect 3868 3974 3895 4026
rect 3947 3974 3974 4026
rect 4026 3974 4053 4026
rect 4105 3974 4131 4026
rect 4183 3974 4189 4026
rect 3810 3962 4189 3974
rect 3810 3910 3816 3962
rect 3868 3910 3895 3962
rect 3947 3910 3974 3962
rect 4026 3910 4053 3962
rect 4105 3910 4131 3962
rect 4183 3910 4189 3962
rect 3810 3903 4189 3910
rect 4249 3903 4681 4033
rect 4686 3903 5678 4033
rect 6103 4028 7095 4033
rect 6103 3976 6109 4028
rect 6161 3976 6174 4028
rect 6226 3976 6239 4028
rect 6291 3976 6304 4028
rect 6356 3976 6368 4028
rect 6420 3976 6432 4028
rect 6484 3976 6496 4028
rect 6548 3976 6560 4028
rect 6612 3976 6624 4028
rect 6676 3976 6688 4028
rect 6740 3976 6752 4028
rect 6804 3976 7095 4028
rect 6103 3956 7095 3976
rect 6103 3904 6109 3956
rect 6161 3904 6174 3956
rect 6226 3904 6239 3956
rect 6291 3904 6304 3956
rect 6356 3904 6368 3956
rect 6420 3904 6432 3956
rect 6484 3904 6496 3956
rect 6548 3904 6560 3956
rect 6612 3904 6624 3956
rect 6676 3904 6688 3956
rect 6740 3904 6752 3956
rect 6804 3904 7095 3956
rect 6103 3903 7095 3904
rect 7657 3981 7663 4033
rect 7715 3981 7729 4033
rect 7781 3981 7787 4033
rect 7657 3955 7787 3981
rect 7657 3903 7663 3955
rect 7715 3903 7729 3955
rect 7781 3903 7787 3955
rect 8232 3981 8595 4033
rect 8647 3981 8660 4033
rect 8712 3981 8724 4033
rect 8776 3981 8788 4033
rect 8840 3981 9202 4033
rect 8232 3959 9202 3981
rect 8232 3907 8595 3959
rect 8647 3907 8660 3959
rect 8712 3907 8724 3959
rect 8776 3907 8788 3959
rect 8840 3907 9202 3959
rect 8232 3903 9202 3907
rect 9769 3986 10750 4033
rect 9769 3934 10220 3986
rect 10272 3934 10286 3986
rect 10338 3934 10352 3986
rect 10404 3934 10418 3986
rect 10470 3934 10483 3986
rect 10535 3934 10548 3986
rect 10600 3934 10613 3986
rect 10665 3934 10678 3986
rect 10730 3934 10750 3986
rect 9769 3903 10750 3934
rect 11193 3987 12185 4033
rect 11193 3935 11631 3987
rect 11683 3935 11696 3987
rect 11748 3935 11761 3987
rect 11813 3935 11826 3987
rect 11878 3935 11891 3987
rect 11943 3935 11956 3987
rect 12008 3935 12021 3987
rect 12073 3935 12185 3987
rect 11193 3903 12185 3935
rect 12747 3981 13053 4033
rect 13105 3981 13120 4033
rect 13172 3981 13187 4033
rect 13239 3981 13254 4033
rect 13306 3981 13321 4033
rect 13373 3981 13388 4033
rect 13440 3981 13455 4033
rect 13507 3981 14039 4033
rect 12747 3955 14039 3981
rect 12747 3903 13053 3955
rect 13105 3903 13120 3955
rect 13172 3903 13187 3955
rect 13239 3903 13254 3955
rect 13306 3903 13321 3955
rect 13373 3903 13388 3955
rect 13440 3903 13455 3955
rect 13507 3903 14039 3955
rect 785 3898 915 3903
rect 441 2973 641 3074
rect 896 953 904 1005
rect 956 953 968 1005
rect 1020 953 1266 1005
rect 1318 953 1330 1005
rect 1382 953 2796 1005
rect 2848 953 2860 1005
rect 2912 953 5653 1005
rect 5705 953 5742 1005
rect 5794 953 5831 1005
rect 5883 953 5920 1005
rect 5972 953 6809 1005
rect 6861 953 6873 1005
rect 6925 953 8511 1005
rect 8563 953 8575 1005
rect 8627 953 9991 1005
rect 10043 953 10055 1005
rect 10107 953 11334 1005
rect 11386 953 11398 1005
rect 11450 953 12768 1005
rect 12820 953 12832 1005
rect 12884 953 14701 1005
rect 14753 953 14765 1005
rect 14817 953 14823 1005
rect 300 915 352 921
tri 352 873 358 879 sw
rect 655 873 663 925
rect 715 873 727 925
rect 779 873 1570 925
rect 1622 873 1634 925
rect 1686 873 3100 925
rect 3152 873 3164 925
rect 3216 873 3875 925
rect 3927 873 3939 925
rect 3991 873 4003 925
rect 4055 873 4067 925
rect 4119 873 4131 925
rect 4183 873 7239 925
rect 7291 873 7303 925
rect 7355 873 8941 925
rect 8993 873 9005 925
rect 9057 873 10421 925
rect 10473 873 10485 925
rect 10537 873 11764 925
rect 11816 873 11828 925
rect 11880 873 13198 925
rect 13250 873 13262 925
rect 13314 873 14781 925
rect 14833 873 14845 925
rect 14897 873 14903 925
rect 352 863 358 873
rect 300 851 358 863
rect 352 845 358 851
tri 358 845 386 873 sw
rect 352 799 421 845
rect 300 793 421 799
rect 473 793 485 845
rect 537 793 1853 845
rect 1905 793 1917 845
rect 1969 793 3383 845
rect 3435 793 3447 845
rect 3499 793 7669 845
rect 7721 793 7733 845
rect 7785 793 9371 845
rect 9423 793 9435 845
rect 9487 793 10851 845
rect 10903 793 10915 845
rect 10967 793 12194 845
rect 12246 793 12258 845
rect 12310 793 13628 845
rect 13680 793 13692 845
rect 13744 793 14772 845
rect 14824 793 14836 845
rect 14888 793 14894 845
<< via1 >>
rect 357 9434 409 9446
rect 357 9400 363 9434
rect 363 9400 397 9434
rect 397 9400 409 9434
rect 357 9394 409 9400
rect 421 9434 473 9446
rect 421 9400 435 9434
rect 435 9400 469 9434
rect 469 9400 473 9434
rect 421 9394 473 9400
rect 791 3969 843 4021
rect 857 3969 909 4021
rect 791 3905 843 3957
rect 857 3905 909 3957
rect 2141 3981 2193 4033
rect 2207 3981 2259 4033
rect 2141 3903 2193 3955
rect 2207 3903 2259 3955
rect 2703 3974 2755 4026
rect 2769 3974 2821 4026
rect 2703 3910 2755 3962
rect 2769 3910 2821 3962
rect 3816 3974 3868 4026
rect 3895 3974 3947 4026
rect 3974 3974 4026 4026
rect 4053 3974 4105 4026
rect 4131 3974 4183 4026
rect 3816 3910 3868 3962
rect 3895 3910 3947 3962
rect 3974 3910 4026 3962
rect 4053 3910 4105 3962
rect 4131 3910 4183 3962
rect 6109 3976 6161 4028
rect 6174 3976 6226 4028
rect 6239 3976 6291 4028
rect 6304 3976 6356 4028
rect 6368 3976 6420 4028
rect 6432 3976 6484 4028
rect 6496 3976 6548 4028
rect 6560 3976 6612 4028
rect 6624 3976 6676 4028
rect 6688 3976 6740 4028
rect 6752 3976 6804 4028
rect 6109 3904 6161 3956
rect 6174 3904 6226 3956
rect 6239 3904 6291 3956
rect 6304 3904 6356 3956
rect 6368 3904 6420 3956
rect 6432 3904 6484 3956
rect 6496 3904 6548 3956
rect 6560 3904 6612 3956
rect 6624 3904 6676 3956
rect 6688 3904 6740 3956
rect 6752 3904 6804 3956
rect 7663 3981 7715 4033
rect 7729 3981 7781 4033
rect 7663 3903 7715 3955
rect 7729 3903 7781 3955
rect 8595 3981 8647 4033
rect 8660 3981 8712 4033
rect 8724 3981 8776 4033
rect 8788 3981 8840 4033
rect 8595 3907 8647 3959
rect 8660 3907 8712 3959
rect 8724 3907 8776 3959
rect 8788 3907 8840 3959
rect 10220 3934 10272 3986
rect 10286 3934 10338 3986
rect 10352 3934 10404 3986
rect 10418 3934 10470 3986
rect 10483 3934 10535 3986
rect 10548 3934 10600 3986
rect 10613 3934 10665 3986
rect 10678 3934 10730 3986
rect 11631 3935 11683 3987
rect 11696 3935 11748 3987
rect 11761 3935 11813 3987
rect 11826 3935 11878 3987
rect 11891 3935 11943 3987
rect 11956 3935 12008 3987
rect 12021 3935 12073 3987
rect 13053 3981 13105 4033
rect 13120 3981 13172 4033
rect 13187 3981 13239 4033
rect 13254 3981 13306 4033
rect 13321 3981 13373 4033
rect 13388 3981 13440 4033
rect 13455 3981 13507 4033
rect 13053 3903 13105 3955
rect 13120 3903 13172 3955
rect 13187 3903 13239 3955
rect 13254 3903 13306 3955
rect 13321 3903 13373 3955
rect 13388 3903 13440 3955
rect 13455 3903 13507 3955
rect 904 953 956 1005
rect 968 953 1020 1005
rect 1266 953 1318 1005
rect 1330 953 1382 1005
rect 2796 953 2848 1005
rect 2860 953 2912 1005
rect 5653 953 5705 1005
rect 5742 953 5794 1005
rect 5831 953 5883 1005
rect 5920 953 5972 1005
rect 6809 953 6861 1005
rect 6873 953 6925 1005
rect 8511 953 8563 1005
rect 8575 953 8627 1005
rect 9991 953 10043 1005
rect 10055 953 10107 1005
rect 11334 953 11386 1005
rect 11398 953 11450 1005
rect 12768 953 12820 1005
rect 12832 953 12884 1005
rect 14701 953 14753 1005
rect 14765 953 14817 1005
rect 300 863 352 915
rect 663 873 715 925
rect 727 873 779 925
rect 1570 873 1622 925
rect 1634 873 1686 925
rect 3100 873 3152 925
rect 3164 873 3216 925
rect 3875 873 3927 925
rect 3939 873 3991 925
rect 4003 873 4055 925
rect 4067 873 4119 925
rect 4131 873 4183 925
rect 7239 873 7291 925
rect 7303 873 7355 925
rect 8941 873 8993 925
rect 9005 873 9057 925
rect 10421 873 10473 925
rect 10485 873 10537 925
rect 11764 873 11816 925
rect 11828 873 11880 925
rect 13198 873 13250 925
rect 13262 873 13314 925
rect 14781 873 14833 925
rect 14845 873 14897 925
rect 300 799 352 851
rect 421 793 473 845
rect 485 793 537 845
rect 1853 793 1905 845
rect 1917 793 1969 845
rect 3383 793 3435 845
rect 3447 793 3499 845
rect 7669 793 7721 845
rect 7733 793 7785 845
rect 9371 793 9423 845
rect 9435 793 9487 845
rect 10851 793 10903 845
rect 10915 793 10967 845
rect 12194 793 12246 845
rect 12258 793 12310 845
rect 13628 793 13680 845
rect 13692 793 13744 845
rect 14772 793 14824 845
rect 14836 793 14888 845
<< metal2 >>
rect 351 9394 357 9446
rect 409 9394 421 9446
rect 473 9394 481 9446
tri 378 9358 414 9394 ne
rect 414 9159 445 9394
tri 445 9358 481 9394 nw
tri 414 9158 415 9159 ne
rect 415 9158 445 9159
tri 445 9158 466 9179 sw
tri 415 9128 445 9158 ne
rect 445 9128 466 9158
tri 445 9107 466 9128 ne
tri 466 9107 517 9158 sw
tri 466 9087 486 9107 ne
tri 444 7391 486 7433 se
rect 486 7422 517 9107
tri 486 7391 517 7422 nw
tri 402 7349 444 7391 se
tri 444 7349 486 7391 nw
tri 360 7307 402 7349 se
tri 402 7307 444 7349 nw
tri 321 7268 360 7307 se
rect 360 7268 363 7307
tri 363 7268 402 7307 nw
tri 304 925 321 942 se
rect 321 925 352 7268
tri 352 7257 363 7268 nw
tri 1802 4028 1807 4033 se
rect 1807 4028 2141 4033
rect 785 4021 915 4028
rect 785 3969 791 4021
rect 843 3969 857 4021
rect 909 3969 915 4021
tri 1755 3981 1802 4028 se
rect 1802 3981 2141 4028
rect 2193 3981 2207 4033
rect 2259 3981 2265 4033
tri 1748 3974 1755 3981 se
rect 1755 3974 2265 3981
rect 785 3957 915 3969
tri 1736 3962 1748 3974 se
rect 1748 3962 2265 3974
rect 785 3905 791 3957
rect 843 3905 857 3957
rect 909 3905 915 3957
tri 1729 3955 1736 3962 se
rect 1736 3955 2265 3962
tri 715 3387 785 3457 se
rect 785 3387 915 3905
tri 1677 3903 1729 3955 se
rect 1729 3903 2141 3955
rect 2193 3903 2207 3955
rect 2259 3903 2265 3955
rect 2697 4026 2827 4033
rect 2697 3974 2703 4026
rect 2755 3974 2769 4026
rect 2821 3974 2827 4026
rect 2697 3962 2827 3974
rect 2697 3910 2703 3962
rect 2755 3910 2769 3962
rect 2821 3910 2827 3962
tri 1623 3849 1677 3903 se
rect 1677 3849 1807 3903
tri 1807 3849 1861 3903 nw
rect 584 3257 915 3387
tri 1497 3723 1623 3849 se
rect 1623 3723 1681 3849
tri 1681 3723 1807 3849 nw
tri 524 1568 584 1628 se
rect 584 1568 714 3257
tri 714 3187 784 3257 nw
tri 1464 1622 1497 1655 se
rect 1497 1622 1627 3723
tri 1627 3669 1681 3723 nw
rect 2697 3319 2827 3910
rect 3810 4026 4189 4033
rect 3810 3974 3816 4026
rect 3868 3974 3895 4026
rect 3947 3974 3974 4026
rect 4026 3974 4053 4026
rect 4105 3974 4131 4026
rect 4183 3974 4189 4026
rect 3810 3962 4189 3974
rect 3810 3910 3816 3962
rect 3868 3910 3895 3962
rect 3947 3910 3974 3962
rect 4026 3910 4053 3962
rect 4105 3910 4131 3962
rect 4183 3910 4189 3962
tri 2827 3319 2852 3344 sw
rect 2697 3290 2852 3319
tri 2697 3135 2852 3290 ne
tri 2852 3135 3036 3319 sw
tri 2852 2951 3036 3135 ne
tri 3036 2951 3220 3135 sw
tri 3036 2897 3090 2951 ne
tri 714 1568 768 1622 sw
tri 1410 1568 1464 1622 se
rect 1464 1568 1627 1622
tri 1627 1568 1714 1655 sw
tri 3003 1568 3090 1655 se
rect 3090 1568 3220 2951
tri 3220 1568 3307 1655 sw
tri 300 921 304 925 se
rect 304 921 352 925
rect 300 915 352 921
rect 300 851 352 863
rect 300 793 352 799
rect 413 1454 1026 1568
rect 413 1402 543 1454
tri 543 1420 577 1454 nw
tri 621 1420 655 1454 ne
rect 414 1400 542 1401
rect 655 1402 785 1454
tri 785 1420 819 1454 nw
tri 862 1420 896 1454 ne
rect 656 1400 784 1401
rect 896 1402 1026 1454
rect 897 1400 1025 1401
rect 1260 1454 1977 1568
rect 1260 1420 1392 1454
tri 1392 1420 1426 1454 nw
tri 1528 1420 1562 1454 ne
rect 1562 1420 1696 1454
tri 1696 1420 1730 1454 nw
tri 1811 1420 1845 1454 ne
rect 1845 1420 1977 1454
rect 1260 1402 1390 1420
tri 1390 1418 1392 1420 nw
tri 1562 1418 1564 1420 ne
rect 1261 1400 1389 1401
rect 1564 1402 1694 1420
tri 1694 1418 1696 1420 nw
tri 1845 1418 1847 1420 ne
rect 1565 1400 1693 1401
rect 1847 1402 1977 1420
rect 1848 1400 1976 1401
rect 2790 1454 3507 1568
rect 2790 1420 2922 1454
tri 2922 1420 2956 1454 nw
tri 3058 1420 3092 1454 ne
rect 3092 1420 3226 1454
tri 3226 1420 3260 1454 nw
tri 3341 1420 3375 1454 ne
rect 3375 1420 3507 1454
rect 2790 1402 2920 1420
tri 2920 1418 2922 1420 nw
tri 3092 1418 3094 1420 ne
rect 2791 1400 2919 1401
rect 3094 1402 3224 1420
tri 3224 1418 3226 1420 nw
tri 3375 1418 3377 1420 ne
rect 3095 1400 3223 1401
rect 3377 1402 3507 1420
rect 3378 1400 3506 1401
rect 413 1100 543 1400
rect 1260 1100 1390 1400
rect 2790 1100 2920 1400
rect 414 1099 542 1100
rect 413 845 543 1098
rect 656 1099 784 1100
rect 655 925 785 1098
rect 897 1099 1025 1100
rect 896 1005 1026 1098
rect 896 953 904 1005
rect 956 953 968 1005
rect 1020 953 1026 1005
rect 1261 1099 1389 1100
rect 1260 1005 1390 1098
rect 1260 953 1266 1005
rect 1318 953 1330 1005
rect 1382 953 1390 1005
rect 1565 1099 1693 1100
rect 655 873 663 925
rect 715 873 727 925
rect 779 873 785 925
rect 1564 925 1694 1098
rect 1564 873 1570 925
rect 1622 873 1634 925
rect 1686 873 1694 925
rect 1848 1099 1976 1100
rect 413 793 421 845
rect 473 793 485 845
rect 537 793 543 845
rect 1847 845 1977 1098
rect 2791 1099 2919 1100
rect 2790 1005 2920 1098
rect 2790 953 2796 1005
rect 2848 953 2860 1005
rect 2912 953 2920 1005
rect 3095 1099 3223 1100
rect 3094 925 3224 1098
rect 3094 873 3100 925
rect 3152 873 3164 925
rect 3216 873 3224 925
rect 3378 1099 3506 1100
rect 1847 793 1853 845
rect 1905 793 1917 845
rect 1969 793 1977 845
rect 3377 845 3507 1098
rect 3810 925 4189 3910
rect 5647 3976 6109 4028
rect 6161 3976 6174 4028
rect 6226 3976 6239 4028
rect 6291 3976 6304 4028
rect 6356 3976 6368 4028
rect 6420 3976 6432 4028
rect 6484 3976 6496 4028
rect 6548 3976 6560 4028
rect 6612 3976 6624 4028
rect 6676 3976 6688 4028
rect 6740 3976 6752 4028
rect 6804 3976 6810 4028
rect 5647 3956 6810 3976
rect 5647 3904 6109 3956
rect 6161 3904 6174 3956
rect 6226 3904 6239 3956
rect 6291 3904 6304 3956
rect 6356 3904 6368 3956
rect 6420 3904 6432 3956
rect 6484 3904 6496 3956
rect 6548 3904 6560 3956
rect 6612 3904 6624 3956
rect 6676 3904 6688 3956
rect 6740 3904 6752 3956
rect 6804 3904 6810 3956
rect 7657 3981 7663 4033
rect 7715 3981 7729 4033
rect 7781 3981 7787 4033
rect 7657 3955 7787 3981
rect 5647 3903 6112 3904
tri 6112 3903 6113 3904 nw
rect 7657 3903 7663 3955
rect 7715 3903 7729 3955
rect 7781 3903 7787 3955
rect 5647 1005 5978 3903
tri 5978 3769 6112 3903 nw
tri 7463 1686 7657 1880 se
rect 7657 1686 7787 3903
rect 8589 3981 8595 4033
rect 8647 3981 8660 4033
rect 8712 3981 8724 4033
rect 8776 3981 8788 4033
rect 8840 3981 8846 4033
rect 8589 3959 8846 3981
rect 8589 3907 8595 3959
rect 8647 3907 8660 3959
rect 8712 3907 8724 3959
rect 8776 3907 8788 3959
rect 8840 3907 8846 3959
tri 7457 1680 7463 1686 se
rect 7463 1680 7787 1686
tri 7787 1680 7793 1686 sw
tri 7389 1612 7457 1680 se
rect 7457 1612 7793 1680
tri 7345 1568 7389 1612 se
rect 7389 1568 7793 1612
tri 8545 1568 8589 1612 se
rect 8589 1568 8846 3907
rect 10214 3986 10736 4017
rect 10214 3934 10220 3986
rect 10272 3934 10286 3986
rect 10338 3934 10352 3986
rect 10404 3934 10418 3986
rect 10470 3934 10483 3986
rect 10535 3934 10548 3986
rect 10600 3934 10613 3986
rect 10665 3934 10678 3986
rect 10730 3934 10736 3986
tri 10132 1618 10214 1700 se
rect 10214 1618 10736 3934
rect 11625 3987 12079 4018
rect 11625 3935 11631 3987
rect 11683 3935 11696 3987
rect 11748 3935 11761 3987
rect 11813 3935 11826 3987
rect 11878 3935 11891 3987
rect 11943 3935 11956 3987
rect 12008 3935 12021 3987
rect 12073 3935 12079 3987
tri 11557 1700 11625 1768 se
rect 11625 1700 12079 3935
rect 13047 3981 13053 4033
rect 13105 3981 13120 4033
rect 13172 3981 13187 4033
rect 13239 3981 13254 4033
rect 13306 3981 13321 4033
rect 13373 3981 13388 4033
rect 13440 3981 13455 4033
rect 13507 3981 13513 4033
rect 13047 3955 13513 3981
rect 13047 3903 13053 3955
rect 13105 3903 13120 3955
rect 13172 3903 13187 3955
rect 13239 3903 13254 3955
rect 13306 3903 13321 3955
rect 13373 3903 13388 3955
rect 13440 3903 13455 3955
rect 13507 3903 13513 3955
tri 13017 1700 13047 1730 se
rect 13047 1700 13513 3903
tri 10736 1618 10818 1700 sw
tri 11475 1618 11557 1700 se
rect 11557 1618 12079 1700
tri 12079 1618 12161 1700 sw
tri 12991 1674 13017 1700 se
rect 13017 1674 13513 1700
tri 12935 1618 12991 1674 se
rect 12991 1618 13513 1674
tri 13513 1618 13569 1674 sw
tri 8846 1568 8896 1618 sw
tri 10082 1568 10132 1618 se
rect 10132 1568 10818 1618
tri 10818 1568 10868 1618 sw
tri 11425 1568 11475 1618 se
rect 11475 1568 12161 1618
tri 12161 1568 12211 1618 sw
tri 12885 1568 12935 1618 se
rect 12935 1568 13569 1618
tri 13569 1568 13619 1618 sw
rect 6803 1454 7793 1568
rect 6803 1402 6933 1454
tri 6933 1418 6969 1454 nw
tri 7197 1418 7233 1454 ne
rect 6804 1400 6932 1401
rect 7233 1402 7363 1454
tri 7363 1418 7399 1454 nw
tri 7627 1418 7663 1454 ne
rect 7234 1400 7362 1401
rect 7663 1402 7793 1454
rect 7664 1400 7792 1401
tri 8505 1528 8545 1568 se
rect 8545 1528 8896 1568
tri 8896 1528 8936 1568 sw
rect 8505 1454 9495 1528
rect 8505 1402 8635 1454
tri 8635 1418 8671 1454 nw
tri 8899 1418 8935 1454 ne
rect 8506 1400 8634 1401
rect 8935 1402 9065 1454
tri 9065 1418 9101 1454 nw
tri 9329 1418 9365 1454 ne
rect 8936 1400 9064 1401
rect 9365 1402 9495 1454
rect 9366 1400 9494 1401
rect 9985 1454 10975 1568
rect 9985 1402 10115 1454
tri 10115 1418 10151 1454 nw
tri 10379 1418 10415 1454 ne
rect 9986 1400 10114 1401
rect 10415 1402 10545 1454
tri 10545 1418 10581 1454 nw
tri 10809 1418 10845 1454 ne
rect 10416 1400 10544 1401
rect 10845 1402 10975 1454
rect 10846 1400 10974 1401
rect 11328 1454 12318 1568
rect 11328 1402 11458 1454
tri 11458 1418 11494 1454 nw
tri 11722 1418 11758 1454 ne
rect 11329 1400 11457 1401
rect 11758 1402 11888 1454
tri 11888 1418 11924 1454 nw
tri 12152 1418 12188 1454 ne
rect 11759 1400 11887 1401
rect 12188 1402 12318 1454
rect 12189 1400 12317 1401
rect 12762 1454 13752 1568
rect 12762 1402 12892 1454
tri 12892 1418 12928 1454 nw
tri 13156 1418 13192 1454 ne
rect 12763 1400 12891 1401
rect 13192 1402 13322 1454
tri 13322 1418 13358 1454 nw
tri 13586 1418 13622 1454 ne
rect 13193 1400 13321 1401
rect 13622 1402 13752 1454
rect 13623 1400 13751 1401
rect 7233 1100 7363 1400
rect 8935 1100 9065 1400
rect 10415 1100 10545 1400
rect 11758 1100 11888 1400
rect 13622 1100 13752 1400
rect 5647 953 5653 1005
rect 5705 953 5742 1005
rect 5794 953 5831 1005
rect 5883 953 5920 1005
rect 5972 953 5978 1005
rect 6804 1099 6932 1100
rect 6803 1005 6933 1098
rect 6803 953 6809 1005
rect 6861 953 6873 1005
rect 6925 953 6933 1005
rect 7234 1099 7362 1100
rect 3810 873 3875 925
rect 3927 873 3939 925
rect 3991 873 4003 925
rect 4055 873 4067 925
rect 4119 873 4131 925
rect 4183 873 4189 925
rect 7233 925 7363 1098
rect 7233 873 7239 925
rect 7291 873 7303 925
rect 7355 873 7363 925
rect 7664 1099 7792 1100
rect 3377 793 3383 845
rect 3435 793 3447 845
rect 3499 793 3507 845
rect 7663 845 7793 1098
rect 8506 1099 8634 1100
rect 8505 1005 8635 1098
rect 8505 953 8511 1005
rect 8563 953 8575 1005
rect 8627 953 8635 1005
rect 8936 1099 9064 1100
rect 8935 925 9065 1098
rect 8935 873 8941 925
rect 8993 873 9005 925
rect 9057 873 9065 925
rect 9366 1099 9494 1100
rect 7663 793 7669 845
rect 7721 793 7733 845
rect 7785 793 7793 845
rect 9365 845 9495 1098
rect 9986 1099 10114 1100
rect 9985 1005 10115 1098
rect 9985 953 9991 1005
rect 10043 953 10055 1005
rect 10107 953 10115 1005
rect 10416 1099 10544 1100
rect 10415 925 10545 1098
rect 10415 873 10421 925
rect 10473 873 10485 925
rect 10537 873 10545 925
rect 10846 1099 10974 1100
rect 9365 793 9371 845
rect 9423 793 9435 845
rect 9487 793 9495 845
rect 10845 845 10975 1098
rect 11329 1099 11457 1100
rect 11328 1005 11458 1098
rect 11328 953 11334 1005
rect 11386 953 11398 1005
rect 11450 953 11458 1005
rect 11759 1099 11887 1100
rect 11758 925 11888 1098
rect 11758 873 11764 925
rect 11816 873 11828 925
rect 11880 873 11888 925
rect 12189 1099 12317 1100
rect 10845 793 10851 845
rect 10903 793 10915 845
rect 10967 793 10975 845
rect 12188 845 12318 1098
rect 12763 1099 12891 1100
rect 12762 1005 12892 1098
rect 12762 953 12768 1005
rect 12820 953 12832 1005
rect 12884 953 12892 1005
rect 13193 1099 13321 1100
rect 13192 925 13322 1098
rect 13192 873 13198 925
rect 13250 873 13262 925
rect 13314 873 13322 925
rect 13623 1099 13751 1100
rect 12188 793 12194 845
rect 12246 793 12258 845
rect 12310 793 12318 845
rect 13622 845 13752 1098
tri 14755 1005 14783 1033 se
rect 14695 953 14701 1005
rect 14753 953 14765 1005
rect 14817 953 14823 1005
tri 14835 925 14863 953 se
rect 14775 873 14781 925
rect 14833 873 14845 925
rect 14897 873 14903 925
tri 14915 845 14943 873 se
rect 13622 793 13628 845
rect 13680 793 13692 845
rect 13744 793 13752 845
rect 14766 793 14772 845
rect 14824 793 14836 845
rect 14888 793 14983 845
<< rmetal2 >>
rect 413 1401 543 1402
rect 413 1400 414 1401
rect 542 1400 543 1401
rect 655 1401 785 1402
rect 655 1400 656 1401
rect 784 1400 785 1401
rect 896 1401 1026 1402
rect 896 1400 897 1401
rect 1025 1400 1026 1401
rect 1260 1401 1390 1402
rect 1260 1400 1261 1401
rect 1389 1400 1390 1401
rect 1564 1401 1694 1402
rect 1564 1400 1565 1401
rect 1693 1400 1694 1401
rect 1847 1401 1977 1402
rect 1847 1400 1848 1401
rect 1976 1400 1977 1401
rect 2790 1401 2920 1402
rect 2790 1400 2791 1401
rect 2919 1400 2920 1401
rect 3094 1401 3224 1402
rect 3094 1400 3095 1401
rect 3223 1400 3224 1401
rect 3377 1401 3507 1402
rect 3377 1400 3378 1401
rect 3506 1400 3507 1401
rect 413 1099 414 1100
rect 542 1099 543 1100
rect 413 1098 543 1099
rect 655 1099 656 1100
rect 784 1099 785 1100
rect 655 1098 785 1099
rect 896 1099 897 1100
rect 1025 1099 1026 1100
rect 896 1098 1026 1099
rect 1260 1099 1261 1100
rect 1389 1099 1390 1100
rect 1260 1098 1390 1099
rect 1564 1099 1565 1100
rect 1693 1099 1694 1100
rect 1564 1098 1694 1099
rect 1847 1099 1848 1100
rect 1976 1099 1977 1100
rect 1847 1098 1977 1099
rect 2790 1099 2791 1100
rect 2919 1099 2920 1100
rect 2790 1098 2920 1099
rect 3094 1099 3095 1100
rect 3223 1099 3224 1100
rect 3094 1098 3224 1099
rect 3377 1099 3378 1100
rect 3506 1099 3507 1100
rect 3377 1098 3507 1099
rect 6803 1401 6933 1402
rect 6803 1400 6804 1401
rect 6932 1400 6933 1401
rect 7233 1401 7363 1402
rect 7233 1400 7234 1401
rect 7362 1400 7363 1401
rect 7663 1401 7793 1402
rect 7663 1400 7664 1401
rect 7792 1400 7793 1401
rect 8505 1401 8635 1402
rect 8505 1400 8506 1401
rect 8634 1400 8635 1401
rect 8935 1401 9065 1402
rect 8935 1400 8936 1401
rect 9064 1400 9065 1401
rect 9365 1401 9495 1402
rect 9365 1400 9366 1401
rect 9494 1400 9495 1401
rect 9985 1401 10115 1402
rect 9985 1400 9986 1401
rect 10114 1400 10115 1401
rect 10415 1401 10545 1402
rect 10415 1400 10416 1401
rect 10544 1400 10545 1401
rect 10845 1401 10975 1402
rect 10845 1400 10846 1401
rect 10974 1400 10975 1401
rect 11328 1401 11458 1402
rect 11328 1400 11329 1401
rect 11457 1400 11458 1401
rect 11758 1401 11888 1402
rect 11758 1400 11759 1401
rect 11887 1400 11888 1401
rect 12188 1401 12318 1402
rect 12188 1400 12189 1401
rect 12317 1400 12318 1401
rect 12762 1401 12892 1402
rect 12762 1400 12763 1401
rect 12891 1400 12892 1401
rect 13192 1401 13322 1402
rect 13192 1400 13193 1401
rect 13321 1400 13322 1401
rect 13622 1401 13752 1402
rect 13622 1400 13623 1401
rect 13751 1400 13752 1401
rect 6803 1099 6804 1100
rect 6932 1099 6933 1100
rect 6803 1098 6933 1099
rect 7233 1099 7234 1100
rect 7362 1099 7363 1100
rect 7233 1098 7363 1099
rect 7663 1099 7664 1100
rect 7792 1099 7793 1100
rect 7663 1098 7793 1099
rect 8505 1099 8506 1100
rect 8634 1099 8635 1100
rect 8505 1098 8635 1099
rect 8935 1099 8936 1100
rect 9064 1099 9065 1100
rect 8935 1098 9065 1099
rect 9365 1099 9366 1100
rect 9494 1099 9495 1100
rect 9365 1098 9495 1099
rect 9985 1099 9986 1100
rect 10114 1099 10115 1100
rect 9985 1098 10115 1099
rect 10415 1099 10416 1100
rect 10544 1099 10545 1100
rect 10415 1098 10545 1099
rect 10845 1099 10846 1100
rect 10974 1099 10975 1100
rect 10845 1098 10975 1099
rect 11328 1099 11329 1100
rect 11457 1099 11458 1100
rect 11328 1098 11458 1099
rect 11758 1099 11759 1100
rect 11887 1099 11888 1100
rect 11758 1098 11888 1099
rect 12188 1099 12189 1100
rect 12317 1099 12318 1100
rect 12188 1098 12318 1099
rect 12762 1099 12763 1100
rect 12891 1099 12892 1100
rect 12762 1098 12892 1099
rect 13192 1099 13193 1100
rect 13321 1099 13322 1100
rect 13192 1098 13322 1099
rect 13622 1099 13623 1100
rect 13751 1099 13752 1100
rect 13622 1098 13752 1099
use sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2  sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0
timestamp 1701704242
transform -1 0 15088 0 -1 8409
box -36 423 15191 5489
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_0
timestamp 1701704242
transform 0 -1 12892 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_1
timestamp 1701704242
transform 0 -1 11458 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_2
timestamp 1701704242
transform 0 -1 10115 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_3
timestamp 1701704242
transform 0 -1 8635 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_4
timestamp 1701704242
transform 0 -1 6933 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_5
timestamp 1701704242
transform 0 -1 13322 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_6
timestamp 1701704242
transform 0 -1 3224 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_7
timestamp 1701704242
transform 0 -1 10975 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_8
timestamp 1701704242
transform 0 -1 9495 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_9
timestamp 1701704242
transform 0 -1 12318 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_10
timestamp 1701704242
transform 0 -1 7793 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_11
timestamp 1701704242
transform 0 -1 3507 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_12
timestamp 1701704242
transform 0 -1 1977 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_13
timestamp 1701704242
transform 0 -1 1694 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_14
timestamp 1701704242
transform 0 1 655 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_15
timestamp 1701704242
transform 0 1 896 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_0
timestamp 1701704242
transform 0 -1 2920 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_1
timestamp 1701704242
transform 0 -1 11888 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_2
timestamp 1701704242
transform 0 -1 7363 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_3
timestamp 1701704242
transform 0 -1 10545 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_4
timestamp 1701704242
transform 0 -1 9065 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_5
timestamp 1701704242
transform 0 -1 13752 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_6
timestamp 1701704242
transform 0 -1 1390 1 0 1046
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_7
timestamp 1701704242
transform 0 1 413 1 0 1046
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1701704242
transform 1 0 464 0 1 9367
box 15 17 2025 18
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1701704242
transform -1 0 2589 0 -1 9417
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1701704242
transform 1 0 379 0 -1 9417
box 0 0 1 1
<< labels >>
flabel comment s 1276 7511 1276 7511 0 FreeSans 440 180 0 0 CONDIODE
flabel comment s 1589 9429 1589 9429 0 FreeSans 440 0 0 0 LEAKER
flabel comment s 2310 1470 2310 1470 0 FreeSans 440 0 0 0 RES
flabel metal1 s 441 2973 641 3074 0 FreeSans 400 0 0 0 VCC_IO
port 2 nsew
flabel metal1 s 14692 953 14777 1005 0 FreeSans 400 0 0 0 PD_H[2]
port 3 nsew
flabel metal1 s 14701 873 14857 925 0 FreeSans 400 0 0 0 PD_H[3]
port 4 nsew
flabel metal1 s 14767 793 14871 845 0 FreeSans 400 0 0 0 TIE_LO_ESD
port 5 nsew
flabel metal1 s 314 9395 405 9439 0 FreeSans 400 0 0 0 TIE_LO_ESD
port 5 nsew
flabel metal1 s 2427 9424 2499 9476 0 FreeSans 400 180 0 0 VGND_IO
port 6 nsew
<< properties >>
string GDS_END 57115692
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 57090256
<< end >>
