magic
tech sky130A
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_0
timestamp 1701704242
transform 1 0 357 0 1 102
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_1
timestamp 1701704242
transform -1 0 653 0 1 102
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808364  sky130_fd_pr__pfet_01v8__example_55959141808364_0
timestamp 1701704242
transform 1 0 490 0 -1 1466
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808364  sky130_fd_pr__pfet_01v8__example_55959141808364_1
timestamp 1701704242
transform 1 0 178 0 -1 1466
box -1 0 257 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1701704242
transform 1 0 251 0 1 1340
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1701704242
transform -1 0 167 0 1 1142
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1701704242
transform -1 0 515 0 1 1142
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1701704242
transform -1 0 791 0 1 1142
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1701704242
transform 1 0 312 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1701704242
transform 1 0 664 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_2
timestamp 1701704242
transform 1 0 601 0 1 912
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1701704242
transform 0 1 121 1 0 735
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1701704242
transform 0 -1 673 1 0 4
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1701704242
transform 0 -1 473 1 0 4
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1701704242
transform 0 1 537 1 0 735
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_1
timestamp 1701704242
transform 0 1 510 -1 0 1564
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_2
timestamp 1701704242
transform 0 1 217 1 0 1498
box 0 0 1 1
<< properties >>
string GDS_END 20880950
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 20876314
<< end >>
