magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 176 626
<< mvnmos >>
rect 0 0 100 600
<< mvndiff >>
rect -50 0 0 600
rect 100 0 150 600
<< poly >>
rect 0 600 100 632
rect 0 -32 100 0
<< metal1 >>
rect -51 -16 -5 546
rect 105 -16 151 546
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 82 626
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_1
timestamp 1701704242
transform 1 0 100 0 1 0
box -26 -26 82 626
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 128 265 128 265 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6695780
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6694886
<< end >>
