magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -191 -26 9693 1426
<< nmos >>
rect 0 0 36 1400
rect 270 0 306 1400
rect 836 0 872 1400
rect 1106 0 1142 1400
rect 1672 0 1708 1400
rect 1942 0 1978 1400
rect 2508 0 2544 1400
rect 2778 0 2814 1400
rect 3344 0 3380 1400
rect 3614 0 3650 1400
rect 4180 0 4216 1400
rect 4450 0 4486 1400
rect 5016 0 5052 1400
rect 5286 0 5322 1400
rect 5852 0 5888 1400
rect 6122 0 6158 1400
rect 6688 0 6724 1400
rect 6958 0 6994 1400
rect 7524 0 7560 1400
rect 7794 0 7830 1400
rect 8360 0 8396 1400
rect 8630 0 8666 1400
rect 9196 0 9232 1400
rect 9466 0 9502 1400
<< ndiff >>
rect -165 0 0 1400
rect 36 0 270 1400
rect 306 0 471 1400
rect 671 0 836 1400
rect 872 0 1106 1400
rect 1142 0 1307 1400
rect 1507 0 1672 1400
rect 1708 0 1942 1400
rect 1978 0 2143 1400
rect 2343 0 2508 1400
rect 2544 0 2778 1400
rect 2814 0 2979 1400
rect 3179 0 3344 1400
rect 3380 0 3614 1400
rect 3650 0 3815 1400
rect 4015 0 4180 1400
rect 4216 0 4450 1400
rect 4486 0 4651 1400
rect 4851 0 5016 1400
rect 5052 0 5286 1400
rect 5322 0 5487 1400
rect 5687 0 5852 1400
rect 5888 0 6122 1400
rect 6158 0 6323 1400
rect 6523 0 6688 1400
rect 6724 0 6958 1400
rect 6994 0 7159 1400
rect 7359 0 7524 1400
rect 7560 0 7794 1400
rect 7830 0 7995 1400
rect 8195 0 8360 1400
rect 8396 0 8630 1400
rect 8666 0 8831 1400
rect 9031 0 9196 1400
rect 9232 0 9466 1400
rect 9502 0 9667 1400
<< poly >>
rect 0 1400 36 1432
rect 270 1400 306 1432
rect 836 1400 872 1432
rect 1106 1400 1142 1432
rect 1672 1400 1708 1432
rect 1942 1400 1978 1432
rect 2508 1400 2544 1432
rect 2778 1400 2814 1432
rect 3344 1400 3380 1432
rect 3614 1400 3650 1432
rect 4180 1400 4216 1432
rect 4450 1400 4486 1432
rect 5016 1400 5052 1432
rect 5286 1400 5322 1432
rect 5852 1400 5888 1432
rect 6122 1400 6158 1432
rect 6688 1400 6724 1432
rect 6958 1400 6994 1432
rect 7524 1400 7560 1432
rect 7794 1400 7830 1432
rect 8360 1400 8396 1432
rect 8630 1400 8666 1432
rect 9196 1400 9232 1432
rect 9466 1400 9502 1432
rect 0 -32 36 0
rect 270 -32 306 0
rect 836 -32 872 0
rect 1106 -32 1142 0
rect 1672 -32 1708 0
rect 1942 -32 1978 0
rect 2508 -32 2544 0
rect 2778 -32 2814 0
rect 3344 -32 3380 0
rect 3614 -32 3650 0
rect 4180 -32 4216 0
rect 4450 -32 4486 0
rect 5016 -32 5052 0
rect 5286 -32 5322 0
rect 5852 -32 5888 0
rect 6122 -32 6158 0
rect 6688 -32 6724 0
rect 6958 -32 6994 0
rect 7524 -32 7560 0
rect 7794 -32 7830 0
rect 8360 -32 8396 0
rect 8630 -32 8666 0
rect 9196 -32 9232 0
rect 9466 -32 9502 0
<< locali >>
rect -354 -4 -176 1354
rect 482 -4 660 1354
rect 1318 -4 1496 1354
rect 2154 -4 2332 1354
rect 2990 -4 3168 1354
rect 3826 -4 4004 1354
rect 4662 -4 4840 1354
rect 5498 -4 5676 1354
rect 6334 -4 6512 1354
rect 7170 -4 7348 1354
rect 8006 -4 8184 1354
rect 8842 -4 9020 1354
rect 9678 -4 9856 1354
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_0
timestamp 1701704242
transform -1 0 -165 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_1
timestamp 1701704242
transform 1 0 471 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_2
timestamp 1701704242
transform 1 0 1307 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_3
timestamp 1701704242
transform 1 0 2143 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_4
timestamp 1701704242
transform 1 0 2979 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_5
timestamp 1701704242
transform 1 0 3815 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_6
timestamp 1701704242
transform 1 0 4651 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_7
timestamp 1701704242
transform 1 0 5487 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_8
timestamp 1701704242
transform 1 0 6323 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_9
timestamp 1701704242
transform 1 0 7159 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_10
timestamp 1701704242
transform 1 0 7995 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_11
timestamp 1701704242
transform 1 0 8831 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_12
timestamp 1701704242
transform 1 0 9667 0 1 0
box -26 -26 226 1426
<< labels >>
flabel comment s 9767 675 9767 675 0 FreeSans 300 0 0 0 S
flabel comment s 9349 700 9349 700 0 FreeSans 300 0 0 0 D
flabel comment s 8931 675 8931 675 0 FreeSans 300 0 0 0 S
flabel comment s 8513 700 8513 700 0 FreeSans 300 0 0 0 D
flabel comment s 8095 675 8095 675 0 FreeSans 300 0 0 0 S
flabel comment s 7677 700 7677 700 0 FreeSans 300 0 0 0 D
flabel comment s 7259 675 7259 675 0 FreeSans 300 0 0 0 S
flabel comment s 6841 700 6841 700 0 FreeSans 300 0 0 0 D
flabel comment s 6423 675 6423 675 0 FreeSans 300 0 0 0 S
flabel comment s 6005 700 6005 700 0 FreeSans 300 0 0 0 D
flabel comment s 5587 675 5587 675 0 FreeSans 300 0 0 0 S
flabel comment s 5169 700 5169 700 0 FreeSans 300 0 0 0 D
flabel comment s 4751 675 4751 675 0 FreeSans 300 0 0 0 S
flabel comment s 4333 700 4333 700 0 FreeSans 300 0 0 0 D
flabel comment s 3915 675 3915 675 0 FreeSans 300 0 0 0 S
flabel comment s 3497 700 3497 700 0 FreeSans 300 0 0 0 D
flabel comment s 3079 675 3079 675 0 FreeSans 300 0 0 0 S
flabel comment s 2661 700 2661 700 0 FreeSans 300 0 0 0 D
flabel comment s 2243 675 2243 675 0 FreeSans 300 0 0 0 S
flabel comment s 1825 700 1825 700 0 FreeSans 300 0 0 0 D
flabel comment s 1407 675 1407 675 0 FreeSans 300 0 0 0 S
flabel comment s 989 700 989 700 0 FreeSans 300 0 0 0 D
flabel comment s 571 675 571 675 0 FreeSans 300 0 0 0 S
flabel comment s 153 700 153 700 0 FreeSans 300 0 0 0 D
flabel comment s -265 675 -265 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 43050326
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43037902
<< end >>
