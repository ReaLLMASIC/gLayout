magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 0 2051 886 2173
<< nsubdiff >>
rect 36 2129 850 2137
rect 36 2095 60 2129
rect 94 2095 128 2129
rect 162 2095 196 2129
rect 230 2095 264 2129
rect 298 2095 332 2129
rect 366 2095 400 2129
rect 434 2095 468 2129
rect 502 2095 536 2129
rect 570 2095 604 2129
rect 638 2095 672 2129
rect 706 2095 740 2129
rect 774 2095 850 2129
rect 36 2087 850 2095
<< nsubdiffcont >>
rect 60 2095 94 2129
rect 128 2095 162 2129
rect 196 2095 230 2129
rect 264 2095 298 2129
rect 332 2095 366 2129
rect 400 2095 434 2129
rect 468 2095 502 2129
rect 536 2095 570 2129
rect 604 2095 638 2129
rect 672 2095 706 2129
rect 740 2095 774 2129
<< poly >>
rect 119 450 239 1753
rect 119 416 182 450
rect 216 416 239 450
rect 119 382 239 416
rect 119 348 182 382
rect 216 348 239 382
rect 119 277 239 348
rect 295 450 415 1753
rect 295 416 337 450
rect 371 416 415 450
rect 295 382 415 416
rect 295 348 337 382
rect 371 348 415 382
rect 295 277 415 348
rect 471 450 591 1753
rect 471 416 510 450
rect 544 416 591 450
rect 471 382 591 416
rect 471 348 510 382
rect 544 348 591 382
rect 471 277 591 348
rect 647 1721 767 1753
rect 647 1687 690 1721
rect 724 1687 767 1721
rect 647 1653 767 1687
rect 647 1619 690 1653
rect 724 1619 767 1653
rect 647 277 767 1619
<< polycont >>
rect 182 416 216 450
rect 182 348 216 382
rect 337 416 371 450
rect 337 348 371 382
rect 510 416 544 450
rect 510 348 544 382
rect 690 1687 724 1721
rect 690 1619 724 1653
<< locali >>
rect 36 2129 850 2137
rect 36 2095 48 2129
rect 94 2095 124 2129
rect 162 2095 196 2129
rect 234 2095 264 2129
rect 310 2095 332 2129
rect 386 2095 400 2129
rect 462 2095 468 2129
rect 502 2095 504 2129
rect 570 2095 579 2129
rect 638 2095 654 2129
rect 706 2095 729 2129
rect 774 2095 804 2129
rect 838 2095 850 2129
rect 36 2087 850 2095
rect 66 1725 119 1985
rect 239 1983 295 2087
rect 591 1983 647 2087
rect 239 1949 250 1983
rect 284 1949 295 1983
rect 239 1911 295 1949
rect 239 1877 250 1911
rect 284 1877 295 1911
rect 239 1781 295 1877
rect 66 1691 76 1725
rect 110 1691 119 1725
rect 66 1653 119 1691
rect 66 1619 76 1653
rect 110 1619 119 1653
rect 66 41 119 1619
rect 415 1725 471 1983
rect 591 1949 602 1983
rect 636 1949 647 1983
rect 591 1911 647 1949
rect 591 1877 602 1911
rect 636 1877 647 1911
rect 591 1781 647 1877
rect 415 1691 426 1725
rect 460 1691 471 1725
rect 415 1653 471 1691
rect 415 1619 426 1653
rect 460 1619 471 1653
rect 415 1607 471 1619
rect 690 1725 724 1737
rect 690 1653 724 1687
rect 690 1603 724 1619
rect 182 450 216 466
rect 182 382 216 416
rect 182 332 216 348
rect 337 450 371 466
rect 337 382 371 416
rect 337 332 371 348
rect 510 450 544 466
rect 510 382 544 416
rect 510 332 544 348
rect 767 41 820 1985
<< viali >>
rect 48 2095 60 2129
rect 60 2095 82 2129
rect 124 2095 128 2129
rect 128 2095 158 2129
rect 200 2095 230 2129
rect 230 2095 234 2129
rect 276 2095 298 2129
rect 298 2095 310 2129
rect 352 2095 366 2129
rect 366 2095 386 2129
rect 428 2095 434 2129
rect 434 2095 462 2129
rect 504 2095 536 2129
rect 536 2095 538 2129
rect 579 2095 604 2129
rect 604 2095 613 2129
rect 654 2095 672 2129
rect 672 2095 688 2129
rect 729 2095 740 2129
rect 740 2095 763 2129
rect 804 2095 838 2129
rect 250 1949 284 1983
rect 250 1877 284 1911
rect 76 1691 110 1725
rect 76 1619 110 1653
rect 602 1949 636 1983
rect 602 1877 636 1911
rect 426 1691 460 1725
rect 426 1619 460 1653
rect 690 1721 724 1725
rect 690 1691 724 1721
rect 690 1619 724 1653
<< metal1 >>
rect 0 2129 886 2135
rect 0 2095 48 2129
rect 82 2095 124 2129
rect 158 2095 200 2129
rect 234 2095 276 2129
rect 310 2095 352 2129
rect 386 2095 428 2129
rect 462 2095 504 2129
rect 538 2095 579 2129
rect 613 2095 654 2129
rect 688 2095 729 2129
rect 763 2095 804 2129
rect 838 2095 886 2129
rect 0 1983 886 2095
rect 0 1949 250 1983
rect 284 1949 602 1983
rect 636 1949 886 1983
rect 0 1911 886 1949
rect 0 1877 250 1911
rect 284 1877 602 1911
rect 636 1877 886 1911
rect 0 1865 886 1877
rect 70 1725 116 1737
rect 420 1725 466 1737
rect 684 1725 730 1737
rect 70 1691 76 1725
rect 110 1695 116 1725
tri 116 1695 146 1725 sw
tri 390 1695 420 1725 se
rect 420 1695 426 1725
rect 110 1691 426 1695
rect 460 1695 466 1725
tri 466 1695 496 1725 sw
tri 654 1695 684 1725 se
rect 684 1695 690 1725
rect 460 1691 690 1695
rect 724 1691 730 1725
rect 70 1653 730 1691
rect 70 1619 76 1653
rect 110 1649 426 1653
rect 110 1619 116 1649
tri 116 1619 146 1649 nw
tri 390 1619 420 1649 ne
rect 420 1619 426 1649
rect 460 1649 690 1653
rect 460 1619 466 1649
tri 466 1619 496 1649 nw
tri 654 1619 684 1649 ne
rect 684 1619 690 1649
rect 724 1619 730 1653
rect 70 1607 116 1619
rect 420 1607 466 1619
rect 684 1607 730 1619
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_0
timestamp 1701704242
transform -1 0 591 0 1 45
box -79 -32 199 232
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_1
timestamp 1701704242
transform -1 0 239 0 1 45
box -79 -32 199 232
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_2
timestamp 1701704242
transform -1 0 415 0 1 45
box -79 -32 199 232
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_3
timestamp 1701704242
transform 1 0 647 0 1 45
box -79 -32 199 232
use pfet_CDNS_52468879185425  pfet_CDNS_52468879185425_0
timestamp 1701704242
transform -1 0 591 0 1 1785
box -119 -66 239 266
use pfet_CDNS_52468879185425  pfet_CDNS_52468879185425_1
timestamp 1701704242
transform -1 0 239 0 1 1785
box -119 -66 239 266
use pfet_CDNS_52468879185425  pfet_CDNS_52468879185425_2
timestamp 1701704242
transform 1 0 295 0 1 1785
box -119 -66 239 266
use pfet_CDNS_52468879185425  pfet_CDNS_52468879185425_3
timestamp 1701704242
transform 1 0 647 0 1 1785
box -119 -66 239 266
<< properties >>
string GDS_END 80615008
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80609178
string path 0.250 52.800 21.900 52.800 
<< end >>
