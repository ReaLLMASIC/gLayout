magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< locali >>
rect 0 2811 1104 2845
rect 179 2136 213 2152
rect 213 2102 817 2136
rect 915 2102 949 2136
rect 179 2086 213 2102
rect 0 1397 1104 1431
rect 179 686 466 705
rect 547 692 834 726
rect 915 692 949 726
rect 547 688 581 692
rect 64 652 98 686
rect 213 671 466 686
rect 179 636 213 652
rect 0 -17 1104 17
<< viali >>
rect 179 2102 213 2136
rect 179 652 213 686
<< metal1 >>
rect 167 2136 225 2142
rect 167 2102 179 2136
rect 213 2102 225 2136
rect 167 2096 225 2102
rect 182 692 210 2096
rect 167 686 225 692
rect 167 652 179 686
rect 213 652 225 686
rect 167 646 225 652
use contact_7  contact_7_0
timestamp 1701704242
transform 1 0 167 0 1 636
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1701704242
transform 1 0 167 0 1 2086
box 0 0 1 1
use pinv_0  pinv_0_0
timestamp 1701704242
transform 1 0 0 0 1 0
box -36 -17 404 1471
use pinv_1  pinv_1_0
timestamp 1701704242
transform 1 0 368 0 1 0
box -36 -17 404 1471
use pinv_2  pinv_2_0
timestamp 1701704242
transform 1 0 736 0 -1 2828
box -36 -17 404 1471
use pinv_2  pinv_2_1
timestamp 1701704242
transform 1 0 736 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 552 0 552 0 4 gnd
port 5 nsew
rlabel locali s 552 2828 552 2828 4 gnd
port 5 nsew
rlabel locali s 932 2119 932 2119 4 Z
port 3 nsew
rlabel locali s 552 1414 552 1414 4 vdd
port 4 nsew
rlabel locali s 81 669 81 669 4 A
port 1 nsew
rlabel locali s 932 709 932 709 4 Zb
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1104 2828
string GDS_END 4849648
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4847828
<< end >>
