magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -85 1532 809 1568
rect -85 800 55 1532
rect 669 800 809 1532
<< pwell >>
rect 679 76 769 728
<< mvpsubdiff >>
rect 705 665 743 702
rect 705 631 707 665
rect 741 631 743 665
rect 705 597 743 631
rect 705 563 707 597
rect 741 563 743 597
rect 705 529 743 563
rect 705 495 707 529
rect 741 495 743 529
rect 705 461 743 495
rect 705 427 707 461
rect 741 427 743 461
rect 705 393 743 427
rect 705 359 707 393
rect 741 359 743 393
rect 705 325 743 359
rect 705 291 707 325
rect 741 291 743 325
rect 705 257 743 291
rect 705 223 707 257
rect 741 223 743 257
rect 705 189 743 223
rect 705 155 707 189
rect 741 155 743 189
rect 705 102 743 155
<< mvnsubdiff >>
rect -19 1413 19 1462
rect -19 1379 -17 1413
rect 17 1379 19 1413
rect -19 1345 19 1379
rect -19 1311 -17 1345
rect 17 1311 19 1345
rect -19 1277 19 1311
rect -19 1243 -17 1277
rect 17 1243 19 1277
rect -19 1209 19 1243
rect -19 1175 -17 1209
rect 17 1175 19 1209
rect -19 1134 19 1175
rect -19 1100 -17 1134
rect 17 1100 19 1134
rect -19 1066 19 1100
rect -19 1032 -17 1066
rect 17 1032 19 1066
rect -19 998 19 1032
rect -19 964 -17 998
rect 17 964 19 998
rect -19 930 19 964
rect -19 896 -17 930
rect 17 896 19 930
rect -19 866 19 896
rect 705 1413 743 1462
rect 705 1379 707 1413
rect 741 1379 743 1413
rect 705 1345 743 1379
rect 705 1311 707 1345
rect 741 1311 743 1345
rect 705 1277 743 1311
rect 705 1243 707 1277
rect 741 1243 743 1277
rect 705 1209 743 1243
rect 705 1175 707 1209
rect 741 1175 743 1209
rect 705 1134 743 1175
rect 705 1100 707 1134
rect 741 1100 743 1134
rect 705 1066 743 1100
rect 705 1032 707 1066
rect 741 1032 743 1066
rect 705 998 743 1032
rect 705 964 707 998
rect 741 964 743 998
rect 705 930 743 964
rect 705 896 707 930
rect 741 896 743 930
rect 705 866 743 896
<< mvpsubdiffcont >>
rect 707 631 741 665
rect 707 563 741 597
rect 707 495 741 529
rect 707 427 741 461
rect 707 359 741 393
rect 707 291 741 325
rect 707 223 741 257
rect 707 155 741 189
<< mvnsubdiffcont >>
rect -17 1379 17 1413
rect -17 1311 17 1345
rect -17 1243 17 1277
rect -17 1175 17 1209
rect -17 1100 17 1134
rect -17 1032 17 1066
rect -17 964 17 998
rect -17 896 17 930
rect 707 1379 741 1413
rect 707 1311 741 1345
rect 707 1243 741 1277
rect 707 1175 741 1209
rect 707 1100 741 1134
rect 707 1032 741 1066
rect 707 964 741 998
rect 707 896 741 930
<< poly >>
rect 126 1548 422 1568
rect 126 1514 155 1548
rect 189 1514 223 1548
rect 257 1514 291 1548
rect 325 1514 359 1548
rect 393 1514 422 1548
rect 126 1492 422 1514
rect 126 793 388 840
rect 126 759 146 793
rect 180 759 214 793
rect 248 759 282 793
rect 316 759 388 793
rect 126 728 388 759
rect 478 783 634 840
rect 478 749 512 783
rect 546 749 580 783
rect 614 749 634 783
rect 478 728 634 749
rect 246 58 388 76
rect 246 24 266 58
rect 300 24 334 58
rect 368 24 388 58
rect 246 8 388 24
rect 444 58 588 76
rect 444 24 466 58
rect 500 24 534 58
rect 568 24 588 58
rect 444 8 588 24
<< polycont >>
rect 155 1514 189 1548
rect 223 1514 257 1548
rect 291 1514 325 1548
rect 359 1514 393 1548
rect 146 759 180 793
rect 214 759 248 793
rect 282 759 316 793
rect 512 749 546 783
rect 580 749 614 783
rect 266 24 300 58
rect 334 24 368 58
rect 466 24 500 58
rect 534 24 568 58
<< locali >>
rect 139 1514 155 1548
rect 189 1514 223 1548
rect 257 1514 291 1548
rect 325 1514 359 1548
rect 393 1514 409 1548
rect -17 1413 17 1454
rect -17 1345 17 1379
rect 707 1413 741 1454
rect 571 1340 609 1374
rect 707 1345 741 1379
rect -17 1277 17 1311
rect -17 1209 17 1243
rect 707 1277 741 1311
rect 707 1209 741 1243
rect -17 1134 17 1175
rect 149 1144 187 1178
rect 361 1144 399 1178
rect -17 1090 17 1100
rect 707 1134 741 1175
rect 707 1090 741 1100
rect -17 1018 17 1032
rect -17 946 17 964
rect 257 1018 291 1056
rect 257 946 291 984
rect 707 1018 741 1032
rect 707 946 741 964
rect -17 874 17 896
rect 609 880 643 928
rect 399 846 643 880
rect 707 874 741 896
rect 130 759 146 793
rect 180 759 214 793
rect 248 759 282 793
rect 316 759 332 793
rect 399 640 433 846
rect 496 749 512 783
rect 546 749 580 783
rect 614 749 630 783
rect 707 665 741 694
rect 707 597 741 631
rect 223 504 257 542
rect 223 432 257 470
rect 575 504 609 542
rect 575 432 609 470
rect 707 529 741 536
rect 707 461 741 464
rect 707 426 741 427
rect 707 325 741 359
rect 707 257 741 291
rect 707 189 741 223
rect 707 110 741 155
rect 250 24 266 58
rect 300 24 334 58
rect 368 24 384 58
rect 450 24 466 58
rect 500 24 534 58
rect 568 24 584 58
<< viali >>
rect 537 1340 571 1374
rect 609 1340 643 1374
rect 115 1144 149 1178
rect 187 1144 221 1178
rect 327 1144 361 1178
rect 399 1144 433 1178
rect -17 1066 17 1090
rect -17 1056 17 1066
rect -17 998 17 1018
rect -17 984 17 998
rect -17 930 17 946
rect -17 912 17 930
rect 257 1056 291 1090
rect 257 984 291 1018
rect 257 912 291 946
rect 707 1066 741 1090
rect 707 1056 741 1066
rect 707 998 741 1018
rect 707 984 741 998
rect 707 930 741 946
rect 707 912 741 930
rect 223 542 257 576
rect 223 470 257 504
rect 223 398 257 432
rect 575 542 609 576
rect 575 470 609 504
rect 575 398 609 432
rect 707 563 741 570
rect 707 536 741 563
rect 707 495 741 498
rect 707 464 741 495
rect 707 393 741 426
rect 707 392 741 393
<< metal1 >>
rect 525 1374 655 1380
rect 525 1340 537 1374
rect 571 1340 609 1374
rect 643 1340 655 1374
rect 525 1334 655 1340
rect 103 1178 445 1184
rect 103 1144 115 1178
rect 149 1144 187 1178
rect 221 1144 327 1178
rect 361 1144 399 1178
rect 433 1144 445 1178
rect 103 1138 445 1144
rect -29 1090 753 1108
rect -29 1056 -17 1090
rect 17 1056 257 1090
rect 291 1056 707 1090
rect 741 1056 753 1090
rect -29 1018 753 1056
rect -29 984 -17 1018
rect 17 984 257 1018
rect 291 984 707 1018
rect 741 984 753 1018
rect -29 946 753 984
rect -29 912 -17 946
rect 17 912 257 946
rect 291 912 707 946
rect 741 912 753 946
rect -29 906 753 912
rect 0 576 753 582
rect 0 542 223 576
rect 257 542 575 576
rect 609 570 753 576
rect 609 542 707 570
rect 0 536 707 542
rect 741 536 753 570
rect 0 504 753 536
rect 0 470 223 504
rect 257 470 575 504
rect 609 498 753 504
rect 609 470 707 498
rect 0 464 707 470
rect 741 464 753 498
rect 0 432 753 464
rect 0 398 223 432
rect 257 398 575 432
rect 609 426 753 432
rect 609 398 707 426
rect 0 392 707 398
rect 741 392 753 426
rect 0 380 753 392
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 221 0 1 1144
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 433 0 1 1144
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 1 0 537 0 1 1340
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1701704242
transform -1 0 741 0 1 912
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1701704242
transform -1 0 741 0 1 392
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1701704242
transform 1 0 223 0 1 398
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_3
timestamp 1701704242
transform 1 0 575 0 1 398
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_4
timestamp 1701704242
transform 1 0 257 0 1 912
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_5
timestamp 1701704242
transform 1 0 -17 0 1 912
box 0 0 1 1
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1701704242
transform -1 0 564 0 1 102
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_1
timestamp 1701704242
transform 1 0 268 0 1 102
box -79 -26 199 626
use pfet_CDNS_52468879185134  pfet_CDNS_52468879185134_0
timestamp 1701704242
transform 1 0 478 0 -1 1466
box -119 -66 239 666
use pfet_CDNS_52468879185137  pfet_CDNS_52468879185137_0
timestamp 1701704242
transform 1 0 126 0 -1 1466
box -119 -66 415 666
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 496 1 0 733
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 0 -1 584 1 0 8
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1701704242
transform 0 -1 384 1 0 8
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 1 130 1 0 743
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform 0 1 139 1 0 1498
box 0 0 1 1
<< labels >>
flabel comment s 334 1166 334 1166 0 FreeSans 200 0 0 0 int
flabel metal1 s 607 1350 607 1350 7 FreeSans 300 180 0 0 pd_h
flabel metal1 s 711 906 753 1108 6 FreeSans 300 180 0 0 vcc_io
port 2 nsew
flabel metal1 s -29 906 13 1108 6 FreeSans 300 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 711 380 753 582 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 0 380 42 582 7 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel locali s 294 759 331 793 6 FreeSans 300 0 0 0 pden_h_n
port 4 nsew
flabel locali s 496 749 530 783 2 FreeSans 300 0 0 0 drvlo_h_n
port 5 nsew
<< properties >>
string GDS_END 87992098
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87986868
<< end >>
