magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 128 2365 10995 3478
rect 128 1020 2015 2365
<< nwell >>
rect 1990 22188 2156 23119
rect 2610 16366 17105 17046
rect -2822 15314 17094 16262
rect 72 1226 374 3538
rect 1807 1226 2109 3538
rect 72 924 2109 1226
<< pwell >>
rect 638 25473 3274 25620
rect 638 23199 1074 25473
rect 2216 24682 3274 25473
rect 3072 23580 3274 24682
rect 444 1512 666 2238
rect 1524 1512 1746 2238
rect 444 1290 1746 1512
rect 4201 2309 4310 2429
<< psubdiff >>
rect 470 2118 640 2146
rect 470 2115 538 2118
rect 504 2084 538 2115
rect 572 2084 606 2118
rect 1550 2118 1720 2146
rect 1550 2117 1618 2118
rect 504 2081 640 2084
rect 470 2048 640 2081
rect 470 2042 538 2048
rect 504 2014 538 2042
rect 572 2014 606 2048
rect 504 2008 640 2014
rect 470 1978 640 2008
rect 470 1969 538 1978
rect 504 1944 538 1969
rect 572 1944 606 1978
rect 504 1935 640 1944
rect 470 1908 640 1935
rect 470 1896 538 1908
rect 504 1874 538 1896
rect 572 1874 606 1908
rect 1584 2084 1618 2117
rect 1652 2115 1720 2118
rect 1652 2084 1686 2115
rect 1584 2083 1686 2084
rect 1550 2081 1686 2083
rect 1550 2048 1720 2081
rect 1550 2046 1618 2048
rect 1584 2014 1618 2046
rect 1652 2042 1720 2048
rect 1652 2014 1686 2042
rect 1584 2012 1686 2014
rect 1550 2008 1686 2012
rect 1550 1978 1720 2008
rect 1550 1976 1618 1978
rect 1584 1944 1618 1976
rect 1652 1969 1720 1978
rect 1652 1944 1686 1969
rect 1584 1942 1686 1944
rect 1550 1935 1686 1942
rect 1550 1908 1720 1935
rect 1550 1906 1618 1908
rect 504 1862 640 1874
rect 470 1838 640 1862
rect 470 1823 538 1838
rect 504 1804 538 1823
rect 572 1804 606 1838
rect 504 1789 640 1804
rect 470 1768 640 1789
rect 470 1750 538 1768
rect 504 1734 538 1750
rect 572 1734 606 1768
rect 504 1716 640 1734
rect 1584 1874 1618 1906
rect 1652 1896 1720 1908
rect 1652 1874 1686 1896
rect 1584 1872 1686 1874
rect 1550 1862 1686 1872
rect 1550 1838 1720 1862
rect 1550 1836 1618 1838
rect 1584 1804 1618 1836
rect 1652 1823 1720 1838
rect 1652 1804 1686 1823
rect 1584 1802 1686 1804
rect 1550 1789 1686 1802
rect 1550 1768 1720 1789
rect 1550 1766 1618 1768
rect 1584 1734 1618 1766
rect 1652 1750 1720 1768
rect 1652 1734 1686 1750
rect 1584 1732 1686 1734
rect 470 1698 640 1716
rect 470 1677 538 1698
rect 504 1664 538 1677
rect 572 1664 606 1698
rect 504 1643 640 1664
rect 470 1628 640 1643
rect 470 1604 538 1628
rect 504 1594 538 1604
rect 572 1594 606 1628
rect 1550 1716 1686 1732
rect 1550 1698 1720 1716
rect 1550 1696 1618 1698
rect 1584 1664 1618 1696
rect 1652 1677 1720 1698
rect 1652 1664 1686 1677
rect 1584 1662 1686 1664
rect 1550 1643 1686 1662
rect 1550 1628 1720 1643
rect 1550 1626 1618 1628
rect 504 1570 640 1594
rect 470 1558 640 1570
rect 470 1531 538 1558
rect 504 1524 538 1531
rect 572 1557 640 1558
rect 572 1524 606 1557
rect 504 1523 606 1524
rect 504 1497 640 1523
rect 470 1488 640 1497
rect 470 1458 538 1488
rect 504 1454 538 1458
rect 572 1486 640 1488
rect 1584 1594 1618 1626
rect 1652 1604 1720 1628
rect 1652 1594 1686 1604
rect 1584 1592 1686 1594
rect 1550 1570 1686 1592
rect 1550 1558 1720 1570
rect 1550 1556 1618 1558
rect 1584 1524 1618 1556
rect 1652 1532 1720 1558
rect 1652 1524 1686 1532
rect 1584 1522 1686 1524
rect 1550 1498 1686 1522
rect 1550 1488 1720 1498
rect 1550 1486 1618 1488
rect 572 1454 606 1486
rect 504 1452 606 1454
rect 640 1452 678 1486
rect 712 1452 750 1486
rect 784 1452 822 1486
rect 856 1452 894 1486
rect 928 1452 966 1486
rect 1000 1452 1039 1486
rect 1073 1452 1112 1486
rect 1146 1452 1185 1486
rect 1219 1452 1258 1486
rect 1292 1452 1331 1486
rect 1365 1452 1404 1486
rect 1438 1452 1477 1486
rect 1511 1452 1550 1486
rect 1584 1454 1618 1486
rect 1652 1460 1720 1488
rect 1652 1454 1686 1460
rect 1584 1452 1686 1454
rect 504 1426 1686 1452
rect 504 1424 1720 1426
rect 470 1418 1720 1424
rect 470 1384 538 1418
rect 572 1384 610 1418
rect 644 1384 682 1418
rect 716 1384 754 1418
rect 788 1384 826 1418
rect 860 1384 898 1418
rect 932 1384 970 1418
rect 1004 1384 1042 1418
rect 1076 1384 1114 1418
rect 1148 1384 1186 1418
rect 1220 1384 1258 1418
rect 1292 1384 1330 1418
rect 1364 1384 1402 1418
rect 1436 1384 1474 1418
rect 1508 1384 1546 1418
rect 1580 1384 1618 1418
rect 1652 1384 1720 1418
rect 504 1350 1720 1384
rect 470 1316 578 1350
rect 612 1316 649 1350
rect 683 1316 720 1350
rect 754 1316 791 1350
rect 825 1316 862 1350
rect 896 1316 933 1350
rect 967 1316 1004 1350
rect 1038 1316 1076 1350
rect 1110 1316 1148 1350
rect 1182 1316 1220 1350
rect 1254 1316 1292 1350
rect 1326 1316 1364 1350
rect 1398 1316 1436 1350
rect 1470 1316 1508 1350
rect 1542 1316 1580 1350
rect 1614 1316 1652 1350
rect 1686 1316 1720 1350
<< mvpsubdiff >>
rect 664 25543 3248 25594
rect 664 25513 2306 25543
rect 664 25003 728 25513
rect 966 25509 2306 25513
rect 2340 25509 2378 25543
rect 2412 25509 2450 25543
rect 2484 25509 2522 25543
rect 2556 25509 2594 25543
rect 2628 25509 2666 25543
rect 2700 25509 2737 25543
rect 2771 25509 2808 25543
rect 2842 25509 2879 25543
rect 2913 25509 2950 25543
rect 2984 25509 3021 25543
rect 3055 25509 3092 25543
rect 3126 25509 3248 25543
rect 966 25499 3248 25509
rect 966 25003 1048 25499
rect 664 24968 1048 25003
rect 664 24934 728 24968
rect 762 24934 796 24968
rect 830 24934 864 24968
rect 898 24934 932 24968
rect 966 24934 1048 24968
rect 664 24899 1048 24934
rect 664 24865 728 24899
rect 762 24865 796 24899
rect 830 24865 864 24899
rect 898 24865 932 24899
rect 966 24865 1048 24899
rect 664 24830 1048 24865
rect 664 24796 728 24830
rect 762 24796 796 24830
rect 830 24796 864 24830
rect 898 24796 932 24830
rect 966 24796 1048 24830
rect 664 24761 1048 24796
rect 664 24727 728 24761
rect 762 24727 796 24761
rect 830 24727 864 24761
rect 898 24727 932 24761
rect 966 24727 1048 24761
rect 664 24692 1048 24727
rect 2242 25475 3248 25499
rect 2242 25441 2306 25475
rect 2340 25441 2378 25475
rect 2412 25441 2450 25475
rect 2484 25441 2522 25475
rect 2556 25441 2594 25475
rect 2628 25441 2666 25475
rect 2700 25441 2737 25475
rect 2771 25441 2808 25475
rect 2842 25441 2879 25475
rect 2913 25441 2950 25475
rect 2984 25441 3021 25475
rect 3055 25441 3092 25475
rect 3126 25441 3248 25475
rect 2242 25407 3248 25441
rect 2242 25373 2306 25407
rect 2340 25373 2378 25407
rect 2412 25373 2450 25407
rect 2484 25373 2522 25407
rect 2556 25373 2594 25407
rect 2628 25373 2666 25407
rect 2700 25373 2737 25407
rect 2771 25373 2808 25407
rect 2842 25373 2879 25407
rect 2913 25373 2950 25407
rect 2984 25373 3021 25407
rect 3055 25373 3092 25407
rect 3126 25373 3248 25407
rect 2242 25339 3248 25373
rect 2242 25305 2306 25339
rect 2340 25305 2378 25339
rect 2412 25305 2450 25339
rect 2484 25305 2522 25339
rect 2556 25305 2594 25339
rect 2628 25305 2666 25339
rect 2700 25305 2737 25339
rect 2771 25305 2808 25339
rect 2842 25305 2879 25339
rect 2913 25305 2950 25339
rect 2984 25305 3021 25339
rect 3055 25305 3092 25339
rect 3126 25305 3248 25339
rect 2242 25271 3248 25305
rect 2242 25237 2306 25271
rect 2340 25237 2378 25271
rect 2412 25237 2450 25271
rect 2484 25237 2522 25271
rect 2556 25237 2594 25271
rect 2628 25237 2666 25271
rect 2700 25237 2737 25271
rect 2771 25237 2808 25271
rect 2842 25237 2879 25271
rect 2913 25237 2950 25271
rect 2984 25237 3021 25271
rect 3055 25237 3092 25271
rect 3126 25237 3248 25271
rect 2242 25203 3248 25237
rect 2242 25169 2306 25203
rect 2340 25169 2378 25203
rect 2412 25169 2450 25203
rect 2484 25169 2522 25203
rect 2556 25169 2594 25203
rect 2628 25169 2666 25203
rect 2700 25169 2737 25203
rect 2771 25169 2808 25203
rect 2842 25169 2879 25203
rect 2913 25169 2950 25203
rect 2984 25169 3021 25203
rect 3055 25169 3092 25203
rect 3126 25169 3248 25203
rect 2242 25135 3248 25169
rect 2242 25101 2306 25135
rect 2340 25101 2378 25135
rect 2412 25101 2450 25135
rect 2484 25101 2522 25135
rect 2556 25101 2594 25135
rect 2628 25101 2666 25135
rect 2700 25101 2737 25135
rect 2771 25101 2808 25135
rect 2842 25101 2879 25135
rect 2913 25101 2950 25135
rect 2984 25101 3021 25135
rect 3055 25101 3092 25135
rect 3126 25101 3248 25135
rect 2242 25067 3248 25101
rect 2242 25033 2306 25067
rect 2340 25033 2378 25067
rect 2412 25033 2450 25067
rect 2484 25033 2522 25067
rect 2556 25033 2594 25067
rect 2628 25033 2666 25067
rect 2700 25033 2737 25067
rect 2771 25033 2808 25067
rect 2842 25033 2879 25067
rect 2913 25033 2950 25067
rect 2984 25033 3021 25067
rect 3055 25033 3092 25067
rect 3126 25033 3248 25067
rect 2242 24999 3248 25033
rect 2242 24965 2306 24999
rect 2340 24965 2378 24999
rect 2412 24965 2450 24999
rect 2484 24965 2522 24999
rect 2556 24965 2594 24999
rect 2628 24965 2666 24999
rect 2700 24965 2737 24999
rect 2771 24965 2808 24999
rect 2842 24965 2879 24999
rect 2913 24965 2950 24999
rect 2984 24965 3021 24999
rect 3055 24965 3092 24999
rect 3126 24965 3248 24999
rect 2242 24931 3248 24965
rect 2242 24897 2306 24931
rect 2340 24897 2378 24931
rect 2412 24897 2450 24931
rect 2484 24897 2522 24931
rect 2556 24897 2594 24931
rect 2628 24897 2666 24931
rect 2700 24897 2737 24931
rect 2771 24897 2808 24931
rect 2842 24897 2879 24931
rect 2913 24897 2950 24931
rect 2984 24897 3021 24931
rect 3055 24897 3092 24931
rect 3126 24897 3248 24931
rect 2242 24863 3248 24897
rect 2242 24829 2306 24863
rect 2340 24829 2378 24863
rect 2412 24829 2450 24863
rect 2484 24829 2522 24863
rect 2556 24829 2594 24863
rect 2628 24829 2666 24863
rect 2700 24829 2737 24863
rect 2771 24829 2808 24863
rect 2842 24829 2879 24863
rect 2913 24829 2950 24863
rect 2984 24829 3021 24863
rect 3055 24829 3092 24863
rect 3126 24829 3248 24863
rect 2242 24795 3248 24829
rect 2242 24761 2306 24795
rect 2340 24761 2378 24795
rect 2412 24761 2450 24795
rect 2484 24761 2522 24795
rect 2556 24761 2594 24795
rect 2628 24761 2666 24795
rect 2700 24761 2737 24795
rect 2771 24761 2808 24795
rect 2842 24761 2879 24795
rect 2913 24761 2950 24795
rect 2984 24761 3021 24795
rect 3055 24761 3092 24795
rect 3126 24761 3248 24795
rect 2242 24708 3248 24761
rect 664 24658 728 24692
rect 762 24658 796 24692
rect 830 24658 864 24692
rect 898 24658 932 24692
rect 966 24658 1048 24692
rect 664 24623 1048 24658
rect 664 24589 728 24623
rect 762 24589 796 24623
rect 830 24589 864 24623
rect 898 24589 932 24623
rect 966 24589 1048 24623
rect 664 24554 1048 24589
rect 664 24520 728 24554
rect 762 24520 796 24554
rect 830 24520 864 24554
rect 898 24520 932 24554
rect 966 24520 1048 24554
rect 664 24485 1048 24520
rect 664 24451 728 24485
rect 762 24451 796 24485
rect 830 24451 864 24485
rect 898 24451 932 24485
rect 966 24451 1048 24485
rect 664 24416 1048 24451
rect 664 24382 728 24416
rect 762 24382 796 24416
rect 830 24382 864 24416
rect 898 24382 932 24416
rect 966 24382 1048 24416
rect 664 24347 1048 24382
rect 664 24313 728 24347
rect 762 24313 796 24347
rect 830 24313 864 24347
rect 898 24313 932 24347
rect 966 24313 1048 24347
rect 664 24278 1048 24313
rect 664 24244 728 24278
rect 762 24244 796 24278
rect 830 24244 864 24278
rect 898 24244 932 24278
rect 966 24244 1048 24278
rect 664 24209 1048 24244
rect 664 24175 728 24209
rect 762 24175 796 24209
rect 830 24175 864 24209
rect 898 24175 932 24209
rect 966 24175 1048 24209
rect 664 24140 1048 24175
rect 664 24106 728 24140
rect 762 24106 796 24140
rect 830 24106 864 24140
rect 898 24106 932 24140
rect 966 24106 1048 24140
rect 664 24071 1048 24106
rect 664 24037 728 24071
rect 762 24037 796 24071
rect 830 24037 864 24071
rect 898 24037 932 24071
rect 966 24037 1048 24071
rect 664 24002 1048 24037
rect 664 23968 728 24002
rect 762 23968 796 24002
rect 830 23968 864 24002
rect 898 23968 932 24002
rect 966 23968 1048 24002
rect 664 23933 1048 23968
rect 664 23899 728 23933
rect 762 23899 796 23933
rect 830 23899 864 23933
rect 898 23899 932 23933
rect 966 23899 1048 23933
rect 664 23864 1048 23899
rect 664 23830 728 23864
rect 762 23830 796 23864
rect 830 23830 864 23864
rect 898 23830 932 23864
rect 966 23830 1048 23864
rect 664 23795 1048 23830
rect 664 23761 728 23795
rect 762 23761 796 23795
rect 830 23761 864 23795
rect 898 23761 932 23795
rect 966 23761 1048 23795
rect 664 23726 1048 23761
rect 664 23692 728 23726
rect 762 23692 796 23726
rect 830 23692 864 23726
rect 898 23692 932 23726
rect 966 23692 1048 23726
rect 664 23657 1048 23692
rect 664 23623 728 23657
rect 762 23623 796 23657
rect 830 23623 864 23657
rect 898 23623 932 23657
rect 966 23623 1048 23657
rect 664 23588 1048 23623
rect 3098 23606 3248 24708
rect 664 23554 728 23588
rect 762 23554 796 23588
rect 830 23554 864 23588
rect 898 23554 932 23588
rect 966 23554 1048 23588
rect 664 23519 1048 23554
rect 664 23485 728 23519
rect 762 23485 796 23519
rect 830 23485 864 23519
rect 898 23485 932 23519
rect 966 23485 1048 23519
rect 664 23450 1048 23485
rect 664 23416 728 23450
rect 762 23416 796 23450
rect 830 23416 864 23450
rect 898 23416 932 23450
rect 966 23416 1048 23450
rect 664 23381 1048 23416
rect 664 23347 728 23381
rect 762 23347 796 23381
rect 830 23347 864 23381
rect 898 23347 932 23381
rect 966 23347 1048 23381
rect 664 23312 1048 23347
rect 664 23278 728 23312
rect 762 23278 796 23312
rect 830 23278 864 23312
rect 898 23278 932 23312
rect 966 23278 1048 23312
rect 664 23225 1048 23278
rect 470 2188 640 2212
rect 504 2154 538 2188
rect 572 2154 606 2188
rect 470 2146 640 2154
rect 1550 2188 1720 2212
rect 1584 2154 1618 2188
rect 1652 2154 1686 2188
rect 1550 2146 1720 2154
<< mvnsubdiff >>
rect 2056 23029 2090 23053
rect 2056 22958 2090 22995
rect 2056 22887 2090 22924
rect 2056 22816 2090 22853
rect 2056 22744 2090 22782
rect 2056 22672 2090 22710
rect 2056 22600 2090 22638
rect 2056 22528 2090 22566
rect 2056 22456 2090 22494
rect 2056 22384 2090 22422
rect 2056 22312 2090 22350
rect 2056 22254 2090 22278
rect 2676 16961 17039 16980
rect 2676 16927 2710 16961
rect 2744 16927 2779 16961
rect 2813 16927 2848 16961
rect 2882 16927 2917 16961
rect 2951 16927 2986 16961
rect 3020 16927 3055 16961
rect 3089 16927 3124 16961
rect 3158 16927 3193 16961
rect 3227 16927 3262 16961
rect 3296 16927 3331 16961
rect 3365 16927 3400 16961
rect 3434 16927 3469 16961
rect 3503 16927 3538 16961
rect 3572 16927 3607 16961
rect 3641 16927 3676 16961
rect 3710 16927 3745 16961
rect 3779 16927 3814 16961
rect 3848 16927 3883 16961
rect 3917 16927 3952 16961
rect 3986 16927 4021 16961
rect 4055 16927 4090 16961
rect 4124 16927 4159 16961
rect 4193 16927 4228 16961
rect 4262 16927 4297 16961
rect 4331 16927 4366 16961
rect 4400 16927 4435 16961
rect 4469 16927 4504 16961
rect 4538 16927 4573 16961
rect 4607 16927 4642 16961
rect 4676 16927 4711 16961
rect 4745 16927 4780 16961
rect 4814 16927 4849 16961
rect 4883 16927 4918 16961
rect 4952 16927 4987 16961
rect 5021 16927 5056 16961
rect 5090 16927 5125 16961
rect 5159 16927 5194 16961
rect 5228 16927 5263 16961
rect 5297 16927 5332 16961
rect 5366 16927 5401 16961
rect 5435 16927 5470 16961
rect 5504 16927 5539 16961
rect 5573 16927 5608 16961
rect 5642 16927 5677 16961
rect 5711 16927 5746 16961
rect 5780 16927 5815 16961
rect 5849 16927 5884 16961
rect 5918 16927 5953 16961
rect 5987 16927 6022 16961
rect 6056 16927 6091 16961
rect 2676 16893 6091 16927
rect 2676 16859 2710 16893
rect 2744 16859 2779 16893
rect 2813 16859 2848 16893
rect 2882 16859 2917 16893
rect 2951 16859 2986 16893
rect 3020 16859 3055 16893
rect 3089 16859 3124 16893
rect 3158 16859 3193 16893
rect 3227 16859 3262 16893
rect 3296 16859 3331 16893
rect 3365 16859 3400 16893
rect 3434 16859 3469 16893
rect 3503 16859 3538 16893
rect 3572 16859 3607 16893
rect 3641 16859 3676 16893
rect 3710 16859 3745 16893
rect 3779 16859 3814 16893
rect 3848 16859 3883 16893
rect 3917 16859 3952 16893
rect 3986 16859 4021 16893
rect 4055 16859 4090 16893
rect 4124 16859 4159 16893
rect 4193 16859 4228 16893
rect 4262 16859 4297 16893
rect 4331 16859 4366 16893
rect 4400 16859 4435 16893
rect 4469 16859 4504 16893
rect 4538 16859 4573 16893
rect 4607 16859 4642 16893
rect 4676 16859 4711 16893
rect 4745 16859 4780 16893
rect 4814 16859 4849 16893
rect 4883 16859 4918 16893
rect 4952 16859 4987 16893
rect 5021 16859 5056 16893
rect 5090 16859 5125 16893
rect 5159 16859 5194 16893
rect 5228 16859 5263 16893
rect 5297 16859 5332 16893
rect 5366 16859 5401 16893
rect 5435 16859 5470 16893
rect 5504 16859 5539 16893
rect 5573 16859 5608 16893
rect 5642 16859 5677 16893
rect 5711 16859 5746 16893
rect 5780 16859 5815 16893
rect 5849 16859 5884 16893
rect 5918 16859 5953 16893
rect 5987 16859 6022 16893
rect 6056 16859 6091 16893
rect 2676 16825 6091 16859
rect 2676 16791 2710 16825
rect 2744 16791 2779 16825
rect 2813 16791 2848 16825
rect 2882 16791 2917 16825
rect 2951 16791 2986 16825
rect 3020 16791 3055 16825
rect 3089 16791 3124 16825
rect 3158 16791 3193 16825
rect 3227 16791 3262 16825
rect 3296 16791 3331 16825
rect 3365 16791 3400 16825
rect 3434 16791 3469 16825
rect 3503 16791 3538 16825
rect 3572 16791 3607 16825
rect 3641 16791 3676 16825
rect 3710 16791 3745 16825
rect 3779 16791 3814 16825
rect 3848 16791 3883 16825
rect 3917 16791 3952 16825
rect 3986 16791 4021 16825
rect 4055 16791 4090 16825
rect 4124 16791 4159 16825
rect 4193 16791 4228 16825
rect 4262 16791 4297 16825
rect 4331 16791 4366 16825
rect 4400 16791 4435 16825
rect 4469 16791 4504 16825
rect 4538 16791 4573 16825
rect 4607 16791 4642 16825
rect 4676 16791 4711 16825
rect 4745 16791 4780 16825
rect 4814 16791 4849 16825
rect 4883 16791 4918 16825
rect 4952 16791 4987 16825
rect 5021 16791 5056 16825
rect 5090 16791 5125 16825
rect 5159 16791 5194 16825
rect 5228 16791 5263 16825
rect 5297 16791 5332 16825
rect 5366 16791 5401 16825
rect 5435 16791 5470 16825
rect 5504 16791 5539 16825
rect 5573 16791 5608 16825
rect 5642 16791 5677 16825
rect 5711 16791 5746 16825
rect 5780 16791 5815 16825
rect 5849 16791 5884 16825
rect 5918 16791 5953 16825
rect 5987 16791 6022 16825
rect 6056 16791 6091 16825
rect 2676 16757 6091 16791
rect 2676 16723 2710 16757
rect 2744 16723 2779 16757
rect 2813 16723 2848 16757
rect 2882 16723 2917 16757
rect 2951 16723 2986 16757
rect 3020 16723 3055 16757
rect 3089 16723 3124 16757
rect 3158 16723 3193 16757
rect 3227 16723 3262 16757
rect 3296 16723 3331 16757
rect 3365 16723 3400 16757
rect 3434 16723 3469 16757
rect 3503 16723 3538 16757
rect 3572 16723 3607 16757
rect 3641 16723 3676 16757
rect 3710 16723 3745 16757
rect 3779 16723 3814 16757
rect 3848 16723 3883 16757
rect 3917 16723 3952 16757
rect 3986 16723 4021 16757
rect 4055 16723 4090 16757
rect 4124 16723 4159 16757
rect 4193 16723 4228 16757
rect 4262 16723 4297 16757
rect 4331 16723 4366 16757
rect 4400 16723 4435 16757
rect 4469 16723 4504 16757
rect 4538 16723 4573 16757
rect 4607 16723 4642 16757
rect 4676 16723 4711 16757
rect 4745 16723 4780 16757
rect 4814 16723 4849 16757
rect 4883 16723 4918 16757
rect 4952 16723 4987 16757
rect 5021 16723 5056 16757
rect 5090 16723 5125 16757
rect 5159 16723 5194 16757
rect 5228 16723 5263 16757
rect 5297 16723 5332 16757
rect 5366 16723 5401 16757
rect 5435 16723 5470 16757
rect 5504 16723 5539 16757
rect 5573 16723 5608 16757
rect 5642 16723 5677 16757
rect 5711 16723 5746 16757
rect 5780 16723 5815 16757
rect 5849 16723 5884 16757
rect 5918 16723 5953 16757
rect 5987 16723 6022 16757
rect 6056 16723 6091 16757
rect 2676 16689 6091 16723
rect 2676 16655 2710 16689
rect 2744 16655 2779 16689
rect 2813 16655 2848 16689
rect 2882 16655 2917 16689
rect 2951 16655 2986 16689
rect 3020 16655 3055 16689
rect 3089 16655 3124 16689
rect 3158 16655 3193 16689
rect 3227 16655 3262 16689
rect 3296 16655 3331 16689
rect 3365 16655 3400 16689
rect 3434 16655 3469 16689
rect 3503 16655 3538 16689
rect 3572 16655 3607 16689
rect 3641 16655 3676 16689
rect 3710 16655 3745 16689
rect 3779 16655 3814 16689
rect 3848 16655 3883 16689
rect 3917 16655 3952 16689
rect 3986 16655 4021 16689
rect 4055 16655 4090 16689
rect 4124 16655 4159 16689
rect 4193 16655 4228 16689
rect 4262 16655 4297 16689
rect 4331 16655 4366 16689
rect 4400 16655 4435 16689
rect 4469 16655 4504 16689
rect 4538 16655 4573 16689
rect 4607 16655 4642 16689
rect 4676 16655 4711 16689
rect 4745 16655 4780 16689
rect 4814 16655 4849 16689
rect 4883 16655 4918 16689
rect 4952 16655 4987 16689
rect 5021 16655 5056 16689
rect 5090 16655 5125 16689
rect 5159 16655 5194 16689
rect 5228 16655 5263 16689
rect 5297 16655 5332 16689
rect 5366 16655 5401 16689
rect 5435 16655 5470 16689
rect 5504 16655 5539 16689
rect 5573 16655 5608 16689
rect 5642 16655 5677 16689
rect 5711 16655 5746 16689
rect 5780 16655 5815 16689
rect 5849 16655 5884 16689
rect 5918 16655 5953 16689
rect 5987 16655 6022 16689
rect 6056 16655 6091 16689
rect 2676 16621 6091 16655
rect 2676 16587 2710 16621
rect 2744 16587 2779 16621
rect 2813 16587 2848 16621
rect 2882 16587 2917 16621
rect 2951 16587 2986 16621
rect 3020 16587 3055 16621
rect 3089 16587 3124 16621
rect 3158 16587 3193 16621
rect 3227 16587 3262 16621
rect 3296 16587 3331 16621
rect 3365 16587 3400 16621
rect 3434 16587 3469 16621
rect 3503 16587 3538 16621
rect 3572 16587 3607 16621
rect 3641 16587 3676 16621
rect 3710 16587 3745 16621
rect 3779 16587 3814 16621
rect 3848 16587 3883 16621
rect 3917 16587 3952 16621
rect 3986 16587 4021 16621
rect 4055 16587 4090 16621
rect 4124 16587 4159 16621
rect 4193 16587 4228 16621
rect 4262 16587 4297 16621
rect 4331 16587 4366 16621
rect 4400 16587 4435 16621
rect 4469 16587 4504 16621
rect 4538 16587 4573 16621
rect 4607 16587 4642 16621
rect 4676 16587 4711 16621
rect 4745 16587 4780 16621
rect 4814 16587 4849 16621
rect 4883 16587 4918 16621
rect 4952 16587 4987 16621
rect 5021 16587 5056 16621
rect 5090 16587 5125 16621
rect 5159 16587 5194 16621
rect 5228 16587 5263 16621
rect 5297 16587 5332 16621
rect 5366 16587 5401 16621
rect 5435 16587 5470 16621
rect 5504 16587 5539 16621
rect 5573 16587 5608 16621
rect 5642 16587 5677 16621
rect 5711 16587 5746 16621
rect 5780 16587 5815 16621
rect 5849 16587 5884 16621
rect 5918 16587 5953 16621
rect 5987 16587 6022 16621
rect 6056 16587 6091 16621
rect 2676 16553 6091 16587
rect 2676 16519 2710 16553
rect 2744 16519 2779 16553
rect 2813 16519 2848 16553
rect 2882 16519 2917 16553
rect 2951 16519 2986 16553
rect 3020 16519 3055 16553
rect 3089 16519 3124 16553
rect 3158 16519 3193 16553
rect 3227 16519 3262 16553
rect 3296 16519 3331 16553
rect 3365 16519 3400 16553
rect 3434 16519 3469 16553
rect 3503 16519 3538 16553
rect 3572 16519 3607 16553
rect 3641 16519 3676 16553
rect 3710 16519 3745 16553
rect 3779 16519 3814 16553
rect 3848 16519 3883 16553
rect 3917 16519 3952 16553
rect 3986 16519 4021 16553
rect 4055 16519 4090 16553
rect 4124 16519 4159 16553
rect 4193 16519 4228 16553
rect 4262 16519 4297 16553
rect 4331 16519 4366 16553
rect 4400 16519 4435 16553
rect 4469 16519 4504 16553
rect 4538 16519 4573 16553
rect 4607 16519 4642 16553
rect 4676 16519 4711 16553
rect 4745 16519 4780 16553
rect 4814 16519 4849 16553
rect 4883 16519 4918 16553
rect 4952 16519 4987 16553
rect 5021 16519 5056 16553
rect 5090 16519 5125 16553
rect 5159 16519 5194 16553
rect 5228 16519 5263 16553
rect 5297 16519 5332 16553
rect 5366 16519 5401 16553
rect 5435 16519 5470 16553
rect 5504 16519 5539 16553
rect 5573 16519 5608 16553
rect 5642 16519 5677 16553
rect 5711 16519 5746 16553
rect 5780 16519 5815 16553
rect 5849 16519 5884 16553
rect 5918 16519 5953 16553
rect 5987 16519 6022 16553
rect 6056 16519 6091 16553
rect 2676 16485 6091 16519
rect 2676 16451 2710 16485
rect 2744 16451 2779 16485
rect 2813 16451 2848 16485
rect 2882 16451 2917 16485
rect 2951 16451 2986 16485
rect 3020 16451 3055 16485
rect 3089 16451 3124 16485
rect 3158 16451 3193 16485
rect 3227 16451 3262 16485
rect 3296 16451 3331 16485
rect 3365 16451 3400 16485
rect 3434 16451 3469 16485
rect 3503 16451 3538 16485
rect 3572 16451 3607 16485
rect 3641 16451 3676 16485
rect 3710 16451 3745 16485
rect 3779 16451 3814 16485
rect 3848 16451 3883 16485
rect 3917 16451 3952 16485
rect 3986 16451 4021 16485
rect 4055 16451 4090 16485
rect 4124 16451 4159 16485
rect 4193 16451 4228 16485
rect 4262 16451 4297 16485
rect 4331 16451 4366 16485
rect 4400 16451 4435 16485
rect 4469 16451 4504 16485
rect 4538 16451 4573 16485
rect 4607 16451 4642 16485
rect 4676 16451 4711 16485
rect 4745 16451 4780 16485
rect 4814 16451 4849 16485
rect 4883 16451 4918 16485
rect 4952 16451 4987 16485
rect 5021 16451 5056 16485
rect 5090 16451 5125 16485
rect 5159 16451 5194 16485
rect 5228 16451 5263 16485
rect 5297 16451 5332 16485
rect 5366 16451 5401 16485
rect 5435 16451 5470 16485
rect 5504 16451 5539 16485
rect 5573 16451 5608 16485
rect 5642 16451 5677 16485
rect 5711 16451 5746 16485
rect 5780 16451 5815 16485
rect 5849 16451 5884 16485
rect 5918 16451 5953 16485
rect 5987 16451 6022 16485
rect 6056 16451 6091 16485
rect 17005 16451 17039 16961
rect 2676 16398 17039 16451
rect -2817 16179 17039 16228
rect -2817 16145 -2732 16179
rect -2698 16145 -2663 16179
rect -2629 16145 -2594 16179
rect -2560 16145 -2525 16179
rect -2491 16145 -2456 16179
rect -2422 16145 -2387 16179
rect -2353 16145 -2318 16179
rect -2284 16145 -2249 16179
rect -2215 16145 -2180 16179
rect -2146 16145 -2111 16179
rect -2077 16145 -2042 16179
rect -2008 16145 -1973 16179
rect -1939 16145 -1904 16179
rect -1870 16145 -1835 16179
rect -1801 16145 -1766 16179
rect -1732 16145 -1697 16179
rect -1663 16145 -1628 16179
rect -1594 16145 -1559 16179
rect -1525 16145 -1490 16179
rect -1456 16145 -1421 16179
rect -1387 16145 -1352 16179
rect -1318 16145 -1283 16179
rect -1249 16145 -1214 16179
rect -1180 16145 -1145 16179
rect -1111 16145 -1076 16179
rect -1042 16145 -1007 16179
rect -973 16145 -938 16179
rect -904 16145 -869 16179
rect -835 16145 -800 16179
rect -766 16145 -731 16179
rect -697 16145 -662 16179
rect -628 16145 -593 16179
rect -559 16145 -524 16179
rect -490 16145 -455 16179
rect -421 16145 -386 16179
rect -352 16145 -317 16179
rect -283 16145 -248 16179
rect -214 16145 -179 16179
rect -145 16145 -110 16179
rect -76 16145 -41 16179
rect -7 16145 28 16179
rect 62 16145 97 16179
rect 131 16145 166 16179
rect 200 16145 235 16179
rect 269 16145 304 16179
rect 338 16145 373 16179
rect 407 16145 442 16179
rect 476 16145 511 16179
rect 545 16145 580 16179
rect 614 16145 649 16179
rect 683 16145 718 16179
rect -2817 16111 718 16145
rect -2817 16077 -2732 16111
rect -2698 16077 -2663 16111
rect -2629 16077 -2594 16111
rect -2560 16077 -2525 16111
rect -2491 16077 -2456 16111
rect -2422 16077 -2387 16111
rect -2353 16077 -2318 16111
rect -2284 16077 -2249 16111
rect -2215 16077 -2180 16111
rect -2146 16077 -2111 16111
rect -2077 16077 -2042 16111
rect -2008 16077 -1973 16111
rect -1939 16077 -1904 16111
rect -1870 16077 -1835 16111
rect -1801 16077 -1766 16111
rect -1732 16077 -1697 16111
rect -1663 16077 -1628 16111
rect -1594 16077 -1559 16111
rect -1525 16077 -1490 16111
rect -1456 16077 -1421 16111
rect -1387 16077 -1352 16111
rect -1318 16077 -1283 16111
rect -1249 16077 -1214 16111
rect -1180 16077 -1145 16111
rect -1111 16077 -1076 16111
rect -1042 16077 -1007 16111
rect -973 16077 -938 16111
rect -904 16077 -869 16111
rect -835 16077 -800 16111
rect -766 16077 -731 16111
rect -697 16077 -662 16111
rect -628 16077 -593 16111
rect -559 16077 -524 16111
rect -490 16077 -455 16111
rect -421 16077 -386 16111
rect -352 16077 -317 16111
rect -283 16077 -248 16111
rect -214 16077 -179 16111
rect -145 16077 -110 16111
rect -76 16077 -41 16111
rect -7 16077 28 16111
rect 62 16077 97 16111
rect 131 16077 166 16111
rect 200 16077 235 16111
rect 269 16077 304 16111
rect 338 16077 373 16111
rect 407 16077 442 16111
rect 476 16077 511 16111
rect 545 16077 580 16111
rect 614 16077 649 16111
rect 683 16077 718 16111
rect -2817 16043 718 16077
rect -2817 16009 -2732 16043
rect -2698 16009 -2663 16043
rect -2629 16009 -2594 16043
rect -2560 16009 -2525 16043
rect -2491 16009 -2456 16043
rect -2422 16009 -2387 16043
rect -2353 16009 -2318 16043
rect -2284 16009 -2249 16043
rect -2215 16009 -2180 16043
rect -2146 16009 -2111 16043
rect -2077 16009 -2042 16043
rect -2008 16009 -1973 16043
rect -1939 16009 -1904 16043
rect -1870 16009 -1835 16043
rect -1801 16009 -1766 16043
rect -1732 16009 -1697 16043
rect -1663 16009 -1628 16043
rect -1594 16009 -1559 16043
rect -1525 16009 -1490 16043
rect -1456 16009 -1421 16043
rect -1387 16009 -1352 16043
rect -1318 16009 -1283 16043
rect -1249 16009 -1214 16043
rect -1180 16009 -1145 16043
rect -1111 16009 -1076 16043
rect -1042 16009 -1007 16043
rect -973 16009 -938 16043
rect -904 16009 -869 16043
rect -835 16009 -800 16043
rect -766 16009 -731 16043
rect -697 16009 -662 16043
rect -628 16009 -593 16043
rect -559 16009 -524 16043
rect -490 16009 -455 16043
rect -421 16009 -386 16043
rect -352 16009 -317 16043
rect -283 16009 -248 16043
rect -214 16009 -179 16043
rect -145 16009 -110 16043
rect -76 16009 -41 16043
rect -7 16009 28 16043
rect 62 16009 97 16043
rect 131 16009 166 16043
rect 200 16009 235 16043
rect 269 16009 304 16043
rect 338 16009 373 16043
rect 407 16009 442 16043
rect 476 16009 511 16043
rect 545 16009 580 16043
rect 614 16009 649 16043
rect 683 16009 718 16043
rect -2817 15975 718 16009
rect -2817 15941 -2732 15975
rect -2698 15941 -2663 15975
rect -2629 15941 -2594 15975
rect -2560 15941 -2525 15975
rect -2491 15941 -2456 15975
rect -2422 15941 -2387 15975
rect -2353 15941 -2318 15975
rect -2284 15941 -2249 15975
rect -2215 15941 -2180 15975
rect -2146 15941 -2111 15975
rect -2077 15941 -2042 15975
rect -2008 15941 -1973 15975
rect -1939 15941 -1904 15975
rect -1870 15941 -1835 15975
rect -1801 15941 -1766 15975
rect -1732 15941 -1697 15975
rect -1663 15941 -1628 15975
rect -1594 15941 -1559 15975
rect -1525 15941 -1490 15975
rect -1456 15941 -1421 15975
rect -1387 15941 -1352 15975
rect -1318 15941 -1283 15975
rect -1249 15941 -1214 15975
rect -1180 15941 -1145 15975
rect -1111 15941 -1076 15975
rect -1042 15941 -1007 15975
rect -973 15941 -938 15975
rect -904 15941 -869 15975
rect -835 15941 -800 15975
rect -766 15941 -731 15975
rect -697 15941 -662 15975
rect -628 15941 -593 15975
rect -559 15941 -524 15975
rect -490 15941 -455 15975
rect -421 15941 -386 15975
rect -352 15941 -317 15975
rect -283 15941 -248 15975
rect -214 15941 -179 15975
rect -145 15941 -110 15975
rect -76 15941 -41 15975
rect -7 15941 28 15975
rect 62 15941 97 15975
rect 131 15941 166 15975
rect 200 15941 235 15975
rect 269 15941 304 15975
rect 338 15941 373 15975
rect 407 15941 442 15975
rect 476 15941 511 15975
rect 545 15941 580 15975
rect 614 15941 649 15975
rect 683 15941 718 15975
rect -2817 15907 718 15941
rect -2817 15873 -2732 15907
rect -2698 15873 -2663 15907
rect -2629 15873 -2594 15907
rect -2560 15873 -2525 15907
rect -2491 15873 -2456 15907
rect -2422 15873 -2387 15907
rect -2353 15873 -2318 15907
rect -2284 15873 -2249 15907
rect -2215 15873 -2180 15907
rect -2146 15873 -2111 15907
rect -2077 15873 -2042 15907
rect -2008 15873 -1973 15907
rect -1939 15873 -1904 15907
rect -1870 15873 -1835 15907
rect -1801 15873 -1766 15907
rect -1732 15873 -1697 15907
rect -1663 15873 -1628 15907
rect -1594 15873 -1559 15907
rect -1525 15873 -1490 15907
rect -1456 15873 -1421 15907
rect -1387 15873 -1352 15907
rect -1318 15873 -1283 15907
rect -1249 15873 -1214 15907
rect -1180 15873 -1145 15907
rect -1111 15873 -1076 15907
rect -1042 15873 -1007 15907
rect -973 15873 -938 15907
rect -904 15873 -869 15907
rect -835 15873 -800 15907
rect -766 15873 -731 15907
rect -697 15873 -662 15907
rect -628 15873 -593 15907
rect -559 15873 -524 15907
rect -490 15873 -455 15907
rect -421 15873 -386 15907
rect -352 15873 -317 15907
rect -283 15873 -248 15907
rect -214 15873 -179 15907
rect -145 15873 -110 15907
rect -76 15873 -41 15907
rect -7 15873 28 15907
rect 62 15873 97 15907
rect 131 15873 166 15907
rect 200 15873 235 15907
rect 269 15873 304 15907
rect 338 15873 373 15907
rect 407 15873 442 15907
rect 476 15873 511 15907
rect 545 15873 580 15907
rect 614 15873 649 15907
rect 683 15873 718 15907
rect -2817 15839 718 15873
rect -2817 15805 -2732 15839
rect -2698 15805 -2663 15839
rect -2629 15805 -2594 15839
rect -2560 15805 -2525 15839
rect -2491 15805 -2456 15839
rect -2422 15805 -2387 15839
rect -2353 15805 -2318 15839
rect -2284 15805 -2249 15839
rect -2215 15805 -2180 15839
rect -2146 15805 -2111 15839
rect -2077 15805 -2042 15839
rect -2008 15805 -1973 15839
rect -1939 15805 -1904 15839
rect -1870 15805 -1835 15839
rect -1801 15805 -1766 15839
rect -1732 15805 -1697 15839
rect -1663 15805 -1628 15839
rect -1594 15805 -1559 15839
rect -1525 15805 -1490 15839
rect -1456 15805 -1421 15839
rect -1387 15805 -1352 15839
rect -1318 15805 -1283 15839
rect -1249 15805 -1214 15839
rect -1180 15805 -1145 15839
rect -1111 15805 -1076 15839
rect -1042 15805 -1007 15839
rect -973 15805 -938 15839
rect -904 15805 -869 15839
rect -835 15805 -800 15839
rect -766 15805 -731 15839
rect -697 15805 -662 15839
rect -628 15805 -593 15839
rect -559 15805 -524 15839
rect -490 15805 -455 15839
rect -421 15805 -386 15839
rect -352 15805 -317 15839
rect -283 15805 -248 15839
rect -214 15805 -179 15839
rect -145 15805 -110 15839
rect -76 15805 -41 15839
rect -7 15805 28 15839
rect 62 15805 97 15839
rect 131 15805 166 15839
rect 200 15805 235 15839
rect 269 15805 304 15839
rect 338 15805 373 15839
rect 407 15805 442 15839
rect 476 15805 511 15839
rect 545 15805 580 15839
rect 614 15805 649 15839
rect 683 15805 718 15839
rect -2817 15771 718 15805
rect -2817 15737 -2732 15771
rect -2698 15737 -2663 15771
rect -2629 15737 -2594 15771
rect -2560 15737 -2525 15771
rect -2491 15737 -2456 15771
rect -2422 15737 -2387 15771
rect -2353 15737 -2318 15771
rect -2284 15737 -2249 15771
rect -2215 15737 -2180 15771
rect -2146 15737 -2111 15771
rect -2077 15737 -2042 15771
rect -2008 15737 -1973 15771
rect -1939 15737 -1904 15771
rect -1870 15737 -1835 15771
rect -1801 15737 -1766 15771
rect -1732 15737 -1697 15771
rect -1663 15737 -1628 15771
rect -1594 15737 -1559 15771
rect -1525 15737 -1490 15771
rect -1456 15737 -1421 15771
rect -1387 15737 -1352 15771
rect -1318 15737 -1283 15771
rect -1249 15737 -1214 15771
rect -1180 15737 -1145 15771
rect -1111 15737 -1076 15771
rect -1042 15737 -1007 15771
rect -973 15737 -938 15771
rect -904 15737 -869 15771
rect -835 15737 -800 15771
rect -766 15737 -731 15771
rect -697 15737 -662 15771
rect -628 15737 -593 15771
rect -559 15737 -524 15771
rect -490 15737 -455 15771
rect -421 15737 -386 15771
rect -352 15737 -317 15771
rect -283 15737 -248 15771
rect -214 15737 -179 15771
rect -145 15737 -110 15771
rect -76 15737 -41 15771
rect -7 15737 28 15771
rect 62 15737 97 15771
rect 131 15737 166 15771
rect 200 15737 235 15771
rect 269 15737 304 15771
rect 338 15737 373 15771
rect 407 15737 442 15771
rect 476 15737 511 15771
rect 545 15737 580 15771
rect 614 15737 649 15771
rect 683 15737 718 15771
rect -2817 15703 718 15737
rect -2817 15669 -2732 15703
rect -2698 15669 -2663 15703
rect -2629 15669 -2594 15703
rect -2560 15669 -2525 15703
rect -2491 15669 -2456 15703
rect -2422 15669 -2387 15703
rect -2353 15669 -2318 15703
rect -2284 15669 -2249 15703
rect -2215 15669 -2180 15703
rect -2146 15669 -2111 15703
rect -2077 15669 -2042 15703
rect -2008 15669 -1973 15703
rect -1939 15669 -1904 15703
rect -1870 15669 -1835 15703
rect -1801 15669 -1766 15703
rect -1732 15669 -1697 15703
rect -1663 15669 -1628 15703
rect -1594 15669 -1559 15703
rect -1525 15669 -1490 15703
rect -1456 15669 -1421 15703
rect -1387 15669 -1352 15703
rect -1318 15669 -1283 15703
rect -1249 15669 -1214 15703
rect -1180 15669 -1145 15703
rect -1111 15669 -1076 15703
rect -1042 15669 -1007 15703
rect -973 15669 -938 15703
rect -904 15669 -869 15703
rect -835 15669 -800 15703
rect -766 15669 -731 15703
rect -697 15669 -662 15703
rect -628 15669 -593 15703
rect -559 15669 -524 15703
rect -490 15669 -455 15703
rect -421 15669 -386 15703
rect -352 15669 -317 15703
rect -283 15669 -248 15703
rect -214 15669 -179 15703
rect -145 15669 -110 15703
rect -76 15669 -41 15703
rect -7 15669 28 15703
rect 62 15669 97 15703
rect 131 15669 166 15703
rect 200 15669 235 15703
rect 269 15669 304 15703
rect 338 15669 373 15703
rect 407 15669 442 15703
rect 476 15669 511 15703
rect 545 15669 580 15703
rect 614 15669 649 15703
rect 683 15669 718 15703
rect -2817 15635 718 15669
rect -2817 15601 -2732 15635
rect -2698 15601 -2663 15635
rect -2629 15601 -2594 15635
rect -2560 15601 -2525 15635
rect -2491 15601 -2456 15635
rect -2422 15601 -2387 15635
rect -2353 15601 -2318 15635
rect -2284 15601 -2249 15635
rect -2215 15601 -2180 15635
rect -2146 15601 -2111 15635
rect -2077 15601 -2042 15635
rect -2008 15601 -1973 15635
rect -1939 15601 -1904 15635
rect -1870 15601 -1835 15635
rect -1801 15601 -1766 15635
rect -1732 15601 -1697 15635
rect -1663 15601 -1628 15635
rect -1594 15601 -1559 15635
rect -1525 15601 -1490 15635
rect -1456 15601 -1421 15635
rect -1387 15601 -1352 15635
rect -1318 15601 -1283 15635
rect -1249 15601 -1214 15635
rect -1180 15601 -1145 15635
rect -1111 15601 -1076 15635
rect -1042 15601 -1007 15635
rect -973 15601 -938 15635
rect -904 15601 -869 15635
rect -835 15601 -800 15635
rect -766 15601 -731 15635
rect -697 15601 -662 15635
rect -628 15601 -593 15635
rect -559 15601 -524 15635
rect -490 15601 -455 15635
rect -421 15601 -386 15635
rect -352 15601 -317 15635
rect -283 15601 -248 15635
rect -214 15601 -179 15635
rect -145 15601 -110 15635
rect -76 15601 -41 15635
rect -7 15601 28 15635
rect 62 15601 97 15635
rect 131 15601 166 15635
rect 200 15601 235 15635
rect 269 15601 304 15635
rect 338 15601 373 15635
rect 407 15601 442 15635
rect 476 15601 511 15635
rect 545 15601 580 15635
rect 614 15601 649 15635
rect 683 15601 718 15635
rect -2817 15567 718 15601
rect -2817 15533 -2732 15567
rect -2698 15533 -2663 15567
rect -2629 15533 -2594 15567
rect -2560 15533 -2525 15567
rect -2491 15533 -2456 15567
rect -2422 15533 -2387 15567
rect -2353 15533 -2318 15567
rect -2284 15533 -2249 15567
rect -2215 15533 -2180 15567
rect -2146 15533 -2111 15567
rect -2077 15533 -2042 15567
rect -2008 15533 -1973 15567
rect -1939 15533 -1904 15567
rect -1870 15533 -1835 15567
rect -1801 15533 -1766 15567
rect -1732 15533 -1697 15567
rect -1663 15533 -1628 15567
rect -1594 15533 -1559 15567
rect -1525 15533 -1490 15567
rect -1456 15533 -1421 15567
rect -1387 15533 -1352 15567
rect -1318 15533 -1283 15567
rect -1249 15533 -1214 15567
rect -1180 15533 -1145 15567
rect -1111 15533 -1076 15567
rect -1042 15533 -1007 15567
rect -973 15533 -938 15567
rect -904 15533 -869 15567
rect -835 15533 -800 15567
rect -766 15533 -731 15567
rect -697 15533 -662 15567
rect -628 15533 -593 15567
rect -559 15533 -524 15567
rect -490 15533 -455 15567
rect -421 15533 -386 15567
rect -352 15533 -317 15567
rect -283 15533 -248 15567
rect -214 15533 -179 15567
rect -145 15533 -110 15567
rect -76 15533 -41 15567
rect -7 15533 28 15567
rect 62 15533 97 15567
rect 131 15533 166 15567
rect 200 15533 235 15567
rect 269 15533 304 15567
rect 338 15533 373 15567
rect 407 15533 442 15567
rect 476 15533 511 15567
rect 545 15533 580 15567
rect 614 15533 649 15567
rect 683 15533 718 15567
rect -2817 15499 718 15533
rect -2817 15465 -2732 15499
rect -2698 15465 -2663 15499
rect -2629 15465 -2594 15499
rect -2560 15465 -2525 15499
rect -2491 15465 -2456 15499
rect -2422 15465 -2387 15499
rect -2353 15465 -2318 15499
rect -2284 15465 -2249 15499
rect -2215 15465 -2180 15499
rect -2146 15465 -2111 15499
rect -2077 15465 -2042 15499
rect -2008 15465 -1973 15499
rect -1939 15465 -1904 15499
rect -1870 15465 -1835 15499
rect -1801 15465 -1766 15499
rect -1732 15465 -1697 15499
rect -1663 15465 -1628 15499
rect -1594 15465 -1559 15499
rect -1525 15465 -1490 15499
rect -1456 15465 -1421 15499
rect -1387 15465 -1352 15499
rect -1318 15465 -1283 15499
rect -1249 15465 -1214 15499
rect -1180 15465 -1145 15499
rect -1111 15465 -1076 15499
rect -1042 15465 -1007 15499
rect -973 15465 -938 15499
rect -904 15465 -869 15499
rect -835 15465 -800 15499
rect -766 15465 -731 15499
rect -697 15465 -662 15499
rect -628 15465 -593 15499
rect -559 15465 -524 15499
rect -490 15465 -455 15499
rect -421 15465 -386 15499
rect -352 15465 -317 15499
rect -283 15465 -248 15499
rect -214 15465 -179 15499
rect -145 15465 -110 15499
rect -76 15465 -41 15499
rect -7 15465 28 15499
rect 62 15465 97 15499
rect 131 15465 166 15499
rect 200 15465 235 15499
rect 269 15465 304 15499
rect 338 15465 373 15499
rect 407 15465 442 15499
rect 476 15465 511 15499
rect 545 15465 580 15499
rect 614 15465 649 15499
rect 683 15465 718 15499
rect -2817 15431 718 15465
rect -2817 15397 -2732 15431
rect -2698 15397 -2663 15431
rect -2629 15397 -2594 15431
rect -2560 15397 -2525 15431
rect -2491 15397 -2456 15431
rect -2422 15397 -2387 15431
rect -2353 15397 -2318 15431
rect -2284 15397 -2249 15431
rect -2215 15397 -2180 15431
rect -2146 15397 -2111 15431
rect -2077 15397 -2042 15431
rect -2008 15397 -1973 15431
rect -1939 15397 -1904 15431
rect -1870 15397 -1835 15431
rect -1801 15397 -1766 15431
rect -1732 15397 -1697 15431
rect -1663 15397 -1628 15431
rect -1594 15397 -1559 15431
rect -1525 15397 -1490 15431
rect -1456 15397 -1421 15431
rect -1387 15397 -1352 15431
rect -1318 15397 -1283 15431
rect -1249 15397 -1214 15431
rect -1180 15397 -1145 15431
rect -1111 15397 -1076 15431
rect -1042 15397 -1007 15431
rect -973 15397 -938 15431
rect -904 15397 -869 15431
rect -835 15397 -800 15431
rect -766 15397 -731 15431
rect -697 15397 -662 15431
rect -628 15397 -593 15431
rect -559 15397 -524 15431
rect -490 15397 -455 15431
rect -421 15397 -386 15431
rect -352 15397 -317 15431
rect -283 15397 -248 15431
rect -214 15397 -179 15431
rect -145 15397 -110 15431
rect -76 15397 -41 15431
rect -7 15397 28 15431
rect 62 15397 97 15431
rect 131 15397 166 15431
rect 200 15397 235 15431
rect 269 15397 304 15431
rect 338 15397 373 15431
rect 407 15397 442 15431
rect 476 15397 511 15431
rect 545 15397 580 15431
rect 614 15397 649 15431
rect 683 15397 718 15431
rect 17004 15397 17039 16179
rect -2817 15380 17039 15397
rect 138 3448 308 3498
rect 172 3414 206 3448
rect 240 3414 274 3448
rect 138 3378 308 3414
rect 172 3344 206 3378
rect 240 3344 274 3378
rect 138 3308 308 3344
rect 172 3274 206 3308
rect 240 3274 274 3308
rect 138 3238 308 3274
rect 172 3204 206 3238
rect 240 3204 274 3238
rect 138 3168 308 3204
rect 172 3134 206 3168
rect 240 3134 274 3168
rect 138 3098 308 3134
rect 172 3064 206 3098
rect 240 3064 274 3098
rect 138 3028 308 3064
rect 172 2994 206 3028
rect 240 2994 274 3028
rect 138 2958 308 2994
rect 172 2924 206 2958
rect 240 2924 274 2958
rect 138 2888 308 2924
rect 172 2854 206 2888
rect 240 2854 274 2888
rect 138 2818 308 2854
rect 172 2784 206 2818
rect 240 2784 274 2818
rect 138 2749 308 2784
rect 172 2715 206 2749
rect 240 2748 308 2749
rect 240 2715 274 2748
rect 138 2714 274 2715
rect 138 2680 308 2714
rect 172 2646 206 2680
rect 240 2678 308 2680
rect 240 2646 274 2678
rect 138 2644 274 2646
rect 138 2611 308 2644
rect 172 2577 206 2611
rect 240 2609 308 2611
rect 240 2577 274 2609
rect 138 2575 274 2577
rect 138 2542 308 2575
rect 172 2508 206 2542
rect 240 2540 308 2542
rect 240 2508 274 2540
rect 138 2506 274 2508
rect 138 2473 308 2506
rect 172 2439 206 2473
rect 240 2471 308 2473
rect 240 2439 274 2471
rect 138 2437 274 2439
rect 138 2404 308 2437
rect 172 2370 206 2404
rect 240 2402 308 2404
rect 240 2370 274 2402
rect 138 2368 274 2370
rect 138 2335 308 2368
rect 172 2301 206 2335
rect 240 2333 308 2335
rect 240 2301 274 2333
rect 138 2299 274 2301
rect 138 2266 308 2299
rect 172 2232 206 2266
rect 240 2264 308 2266
rect 240 2232 274 2264
rect 138 2230 274 2232
rect 138 2197 308 2230
rect 1873 3448 2043 3498
rect 1907 3414 1941 3448
rect 1975 3414 2009 3448
rect 1873 3379 2043 3414
rect 1907 3345 1941 3379
rect 1975 3345 2009 3379
rect 1873 3310 2043 3345
rect 1907 3276 1941 3310
rect 1975 3276 2009 3310
rect 1873 3241 2043 3276
rect 1907 3207 1941 3241
rect 1975 3207 2009 3241
rect 1873 3172 2043 3207
rect 1907 3138 1941 3172
rect 1975 3138 2009 3172
rect 1873 3103 2043 3138
rect 1907 3069 1941 3103
rect 1975 3069 2009 3103
rect 1873 3034 2043 3069
rect 1907 3000 1941 3034
rect 1975 3000 2009 3034
rect 1873 2965 2043 3000
rect 1907 2931 1941 2965
rect 1975 2931 2009 2965
rect 1873 2896 2043 2931
rect 1907 2862 1941 2896
rect 1975 2862 2009 2896
rect 1873 2827 2043 2862
rect 1907 2793 1941 2827
rect 1975 2793 2009 2827
rect 1873 2758 2043 2793
rect 1907 2724 1941 2758
rect 1975 2724 2009 2758
rect 1873 2689 2043 2724
rect 1907 2655 1941 2689
rect 1975 2655 2009 2689
rect 1873 2620 2043 2655
rect 1907 2586 1941 2620
rect 1975 2586 2009 2620
rect 1873 2551 2043 2586
rect 1907 2517 1941 2551
rect 1975 2517 2009 2551
rect 1873 2482 2043 2517
rect 1907 2448 1941 2482
rect 1975 2448 2009 2482
rect 1873 2413 2043 2448
rect 1907 2379 1941 2413
rect 1975 2379 2009 2413
rect 1873 2344 2043 2379
rect 1907 2310 1941 2344
rect 1975 2310 2009 2344
rect 1873 2275 2043 2310
rect 1907 2241 1941 2275
rect 1975 2241 2009 2275
rect 172 2163 206 2197
rect 240 2195 308 2197
rect 240 2163 274 2195
rect 138 2161 274 2163
rect 138 2128 308 2161
rect 172 2094 206 2128
rect 240 2126 308 2128
rect 240 2094 274 2126
rect 138 2092 274 2094
rect 138 2059 308 2092
rect 172 2025 206 2059
rect 240 2057 308 2059
rect 240 2025 274 2057
rect 138 2023 274 2025
rect 138 1990 308 2023
rect 172 1956 206 1990
rect 240 1988 308 1990
rect 240 1956 274 1988
rect 138 1954 274 1956
rect 138 1921 308 1954
rect 172 1887 206 1921
rect 240 1919 308 1921
rect 240 1887 274 1919
rect 138 1885 274 1887
rect 138 1852 308 1885
rect 172 1818 206 1852
rect 240 1850 308 1852
rect 240 1818 274 1850
rect 138 1816 274 1818
rect 138 1783 308 1816
rect 172 1749 206 1783
rect 240 1781 308 1783
rect 240 1749 274 1781
rect 138 1747 274 1749
rect 138 1714 308 1747
rect 172 1680 206 1714
rect 240 1712 308 1714
rect 240 1680 274 1712
rect 138 1678 274 1680
rect 138 1645 308 1678
rect 172 1611 206 1645
rect 240 1643 308 1645
rect 240 1611 274 1643
rect 138 1609 274 1611
rect 138 1576 308 1609
rect 172 1542 206 1576
rect 240 1574 308 1576
rect 240 1542 274 1574
rect 138 1540 274 1542
rect 138 1507 308 1540
rect 172 1473 206 1507
rect 240 1505 308 1507
rect 240 1473 274 1505
rect 138 1471 274 1473
rect 138 1438 308 1471
rect 172 1404 206 1438
rect 240 1436 308 1438
rect 240 1404 274 1436
rect 138 1402 274 1404
rect 138 1369 308 1402
rect 172 1335 206 1369
rect 240 1367 308 1369
rect 240 1335 274 1367
rect 138 1333 274 1335
rect 138 1300 308 1333
rect 1873 2206 2043 2241
rect 1907 2172 1941 2206
rect 1975 2172 2009 2206
rect 1873 2137 2043 2172
rect 1907 2103 1941 2137
rect 1975 2103 2009 2137
rect 1873 2068 2043 2103
rect 1907 2034 1941 2068
rect 1975 2034 2009 2068
rect 1873 1999 2043 2034
rect 1907 1965 1941 1999
rect 1975 1965 2009 1999
rect 1873 1930 2043 1965
rect 1907 1896 1941 1930
rect 1975 1896 2009 1930
rect 1873 1861 2043 1896
rect 1873 1860 1941 1861
rect 1907 1827 1941 1860
rect 1975 1827 2009 1861
rect 1907 1826 2043 1827
rect 1873 1792 2043 1826
rect 1873 1790 1941 1792
rect 1907 1758 1941 1790
rect 1975 1758 2009 1792
rect 1907 1756 2043 1758
rect 1873 1722 2043 1756
rect 1873 1720 1941 1722
rect 1907 1688 1941 1720
rect 1975 1688 2009 1722
rect 1907 1686 2043 1688
rect 1873 1652 2043 1686
rect 1873 1650 1941 1652
rect 1907 1618 1941 1650
rect 1975 1618 2009 1652
rect 1907 1616 2043 1618
rect 1873 1582 2043 1616
rect 1873 1580 1941 1582
rect 1907 1548 1941 1580
rect 1975 1548 2009 1582
rect 1907 1546 2043 1548
rect 1873 1512 2043 1546
rect 1873 1510 1941 1512
rect 1907 1478 1941 1510
rect 1975 1478 2009 1512
rect 1907 1476 2043 1478
rect 1873 1442 2043 1476
rect 1873 1440 1941 1442
rect 1907 1408 1941 1440
rect 1975 1408 2009 1442
rect 1907 1406 2043 1408
rect 1873 1372 2043 1406
rect 1873 1370 1941 1372
rect 1907 1338 1941 1370
rect 1975 1338 2009 1372
rect 1907 1336 2043 1338
rect 172 1266 206 1300
rect 240 1298 308 1300
rect 240 1266 274 1298
rect 138 1264 274 1266
rect 138 1231 308 1264
rect 172 1197 206 1231
rect 240 1229 308 1231
rect 240 1197 274 1229
rect 138 1195 274 1197
rect 138 1162 308 1195
rect 172 1128 206 1162
rect 240 1160 308 1162
rect 1873 1302 2043 1336
rect 1873 1300 1941 1302
rect 1907 1268 1941 1300
rect 1975 1268 2009 1302
rect 1907 1266 2043 1268
rect 1873 1232 2043 1266
rect 1873 1230 1941 1232
rect 1907 1198 1941 1230
rect 1975 1198 2009 1232
rect 1907 1196 2043 1198
rect 1873 1162 2043 1196
rect 1873 1160 1941 1162
rect 240 1128 274 1160
rect 138 1126 274 1128
rect 308 1126 344 1160
rect 378 1126 414 1160
rect 448 1126 484 1160
rect 518 1126 554 1160
rect 588 1126 624 1160
rect 658 1126 694 1160
rect 728 1126 764 1160
rect 798 1126 834 1160
rect 868 1126 904 1160
rect 938 1126 974 1160
rect 1008 1126 1044 1160
rect 1078 1126 1114 1160
rect 1148 1126 1183 1160
rect 1217 1126 1252 1160
rect 1286 1126 1321 1160
rect 1355 1126 1390 1160
rect 1424 1126 1459 1160
rect 1493 1126 1528 1160
rect 1562 1126 1597 1160
rect 1631 1126 1666 1160
rect 1700 1126 1735 1160
rect 1769 1126 1804 1160
rect 1838 1126 1873 1160
rect 1907 1128 1941 1160
rect 1975 1128 2009 1162
rect 1907 1126 2043 1128
rect 138 1093 2043 1126
rect 172 1092 2043 1093
rect 172 1059 206 1092
rect 138 1058 206 1059
rect 240 1058 276 1092
rect 310 1058 346 1092
rect 380 1058 416 1092
rect 450 1058 486 1092
rect 520 1058 556 1092
rect 590 1058 626 1092
rect 660 1058 696 1092
rect 730 1058 766 1092
rect 800 1058 836 1092
rect 870 1058 905 1092
rect 939 1058 974 1092
rect 1008 1058 1043 1092
rect 1077 1058 1112 1092
rect 1146 1058 1181 1092
rect 1215 1058 1250 1092
rect 1284 1058 1319 1092
rect 1353 1058 1388 1092
rect 1422 1058 1457 1092
rect 1491 1058 1526 1092
rect 1560 1058 1595 1092
rect 1629 1058 1664 1092
rect 1698 1058 1733 1092
rect 1767 1058 1802 1092
rect 1836 1058 1871 1092
rect 1905 1058 1941 1092
rect 1975 1058 2009 1092
rect 138 1024 2043 1058
rect 138 990 206 1024
rect 240 990 276 1024
rect 310 990 346 1024
rect 380 990 416 1024
rect 450 990 486 1024
rect 520 990 556 1024
rect 590 990 626 1024
rect 660 990 696 1024
rect 730 990 766 1024
rect 800 990 836 1024
rect 870 990 905 1024
rect 939 990 974 1024
rect 1008 990 1043 1024
rect 1077 990 1112 1024
rect 1146 990 1181 1024
rect 1215 990 1250 1024
rect 1284 990 1319 1024
rect 1353 990 1388 1024
rect 1422 990 1457 1024
rect 1491 990 1526 1024
rect 1560 990 1595 1024
rect 1629 990 1664 1024
rect 1698 990 1733 1024
rect 1767 990 1802 1024
rect 1836 990 1871 1024
rect 1905 990 1940 1024
rect 1974 990 2043 1024
<< psubdiffcont >>
rect 470 2081 504 2115
rect 538 2084 572 2118
rect 606 2084 640 2118
rect 470 2008 504 2042
rect 538 2014 572 2048
rect 606 2014 640 2048
rect 470 1935 504 1969
rect 538 1944 572 1978
rect 606 1944 640 1978
rect 470 1862 504 1896
rect 538 1874 572 1908
rect 606 1874 640 1908
rect 1550 2083 1584 2117
rect 1618 2084 1652 2118
rect 1686 2081 1720 2115
rect 1550 2012 1584 2046
rect 1618 2014 1652 2048
rect 1686 2008 1720 2042
rect 1550 1942 1584 1976
rect 1618 1944 1652 1978
rect 1686 1935 1720 1969
rect 470 1789 504 1823
rect 538 1804 572 1838
rect 606 1804 640 1838
rect 470 1716 504 1750
rect 538 1734 572 1768
rect 606 1734 640 1768
rect 1550 1872 1584 1906
rect 1618 1874 1652 1908
rect 1686 1862 1720 1896
rect 1550 1802 1584 1836
rect 1618 1804 1652 1838
rect 1686 1789 1720 1823
rect 1550 1732 1584 1766
rect 1618 1734 1652 1768
rect 470 1643 504 1677
rect 538 1664 572 1698
rect 606 1664 640 1698
rect 470 1570 504 1604
rect 538 1594 572 1628
rect 606 1594 640 1628
rect 1686 1716 1720 1750
rect 1550 1662 1584 1696
rect 1618 1664 1652 1698
rect 1686 1643 1720 1677
rect 470 1497 504 1531
rect 538 1524 572 1558
rect 606 1523 640 1557
rect 470 1424 504 1458
rect 538 1454 572 1488
rect 1550 1592 1584 1626
rect 1618 1594 1652 1628
rect 1686 1570 1720 1604
rect 1550 1522 1584 1556
rect 1618 1524 1652 1558
rect 1686 1498 1720 1532
rect 606 1452 640 1486
rect 678 1452 712 1486
rect 750 1452 784 1486
rect 822 1452 856 1486
rect 894 1452 928 1486
rect 966 1452 1000 1486
rect 1039 1452 1073 1486
rect 1112 1452 1146 1486
rect 1185 1452 1219 1486
rect 1258 1452 1292 1486
rect 1331 1452 1365 1486
rect 1404 1452 1438 1486
rect 1477 1452 1511 1486
rect 1550 1452 1584 1486
rect 1618 1454 1652 1488
rect 1686 1426 1720 1460
rect 538 1384 572 1418
rect 610 1384 644 1418
rect 682 1384 716 1418
rect 754 1384 788 1418
rect 826 1384 860 1418
rect 898 1384 932 1418
rect 970 1384 1004 1418
rect 1042 1384 1076 1418
rect 1114 1384 1148 1418
rect 1186 1384 1220 1418
rect 1258 1384 1292 1418
rect 1330 1384 1364 1418
rect 1402 1384 1436 1418
rect 1474 1384 1508 1418
rect 1546 1384 1580 1418
rect 1618 1384 1652 1418
rect 470 1350 504 1384
rect 578 1316 612 1350
rect 649 1316 683 1350
rect 720 1316 754 1350
rect 791 1316 825 1350
rect 862 1316 896 1350
rect 933 1316 967 1350
rect 1004 1316 1038 1350
rect 1076 1316 1110 1350
rect 1148 1316 1182 1350
rect 1220 1316 1254 1350
rect 1292 1316 1326 1350
rect 1364 1316 1398 1350
rect 1436 1316 1470 1350
rect 1508 1316 1542 1350
rect 1580 1316 1614 1350
rect 1652 1316 1686 1350
<< mvpsubdiffcont >>
rect 728 25003 966 25513
rect 2306 25509 2340 25543
rect 2378 25509 2412 25543
rect 2450 25509 2484 25543
rect 2522 25509 2556 25543
rect 2594 25509 2628 25543
rect 2666 25509 2700 25543
rect 2737 25509 2771 25543
rect 2808 25509 2842 25543
rect 2879 25509 2913 25543
rect 2950 25509 2984 25543
rect 3021 25509 3055 25543
rect 3092 25509 3126 25543
rect 728 24934 762 24968
rect 796 24934 830 24968
rect 864 24934 898 24968
rect 932 24934 966 24968
rect 728 24865 762 24899
rect 796 24865 830 24899
rect 864 24865 898 24899
rect 932 24865 966 24899
rect 728 24796 762 24830
rect 796 24796 830 24830
rect 864 24796 898 24830
rect 932 24796 966 24830
rect 728 24727 762 24761
rect 796 24727 830 24761
rect 864 24727 898 24761
rect 932 24727 966 24761
rect 2306 25441 2340 25475
rect 2378 25441 2412 25475
rect 2450 25441 2484 25475
rect 2522 25441 2556 25475
rect 2594 25441 2628 25475
rect 2666 25441 2700 25475
rect 2737 25441 2771 25475
rect 2808 25441 2842 25475
rect 2879 25441 2913 25475
rect 2950 25441 2984 25475
rect 3021 25441 3055 25475
rect 3092 25441 3126 25475
rect 2306 25373 2340 25407
rect 2378 25373 2412 25407
rect 2450 25373 2484 25407
rect 2522 25373 2556 25407
rect 2594 25373 2628 25407
rect 2666 25373 2700 25407
rect 2737 25373 2771 25407
rect 2808 25373 2842 25407
rect 2879 25373 2913 25407
rect 2950 25373 2984 25407
rect 3021 25373 3055 25407
rect 3092 25373 3126 25407
rect 2306 25305 2340 25339
rect 2378 25305 2412 25339
rect 2450 25305 2484 25339
rect 2522 25305 2556 25339
rect 2594 25305 2628 25339
rect 2666 25305 2700 25339
rect 2737 25305 2771 25339
rect 2808 25305 2842 25339
rect 2879 25305 2913 25339
rect 2950 25305 2984 25339
rect 3021 25305 3055 25339
rect 3092 25305 3126 25339
rect 2306 25237 2340 25271
rect 2378 25237 2412 25271
rect 2450 25237 2484 25271
rect 2522 25237 2556 25271
rect 2594 25237 2628 25271
rect 2666 25237 2700 25271
rect 2737 25237 2771 25271
rect 2808 25237 2842 25271
rect 2879 25237 2913 25271
rect 2950 25237 2984 25271
rect 3021 25237 3055 25271
rect 3092 25237 3126 25271
rect 2306 25169 2340 25203
rect 2378 25169 2412 25203
rect 2450 25169 2484 25203
rect 2522 25169 2556 25203
rect 2594 25169 2628 25203
rect 2666 25169 2700 25203
rect 2737 25169 2771 25203
rect 2808 25169 2842 25203
rect 2879 25169 2913 25203
rect 2950 25169 2984 25203
rect 3021 25169 3055 25203
rect 3092 25169 3126 25203
rect 2306 25101 2340 25135
rect 2378 25101 2412 25135
rect 2450 25101 2484 25135
rect 2522 25101 2556 25135
rect 2594 25101 2628 25135
rect 2666 25101 2700 25135
rect 2737 25101 2771 25135
rect 2808 25101 2842 25135
rect 2879 25101 2913 25135
rect 2950 25101 2984 25135
rect 3021 25101 3055 25135
rect 3092 25101 3126 25135
rect 2306 25033 2340 25067
rect 2378 25033 2412 25067
rect 2450 25033 2484 25067
rect 2522 25033 2556 25067
rect 2594 25033 2628 25067
rect 2666 25033 2700 25067
rect 2737 25033 2771 25067
rect 2808 25033 2842 25067
rect 2879 25033 2913 25067
rect 2950 25033 2984 25067
rect 3021 25033 3055 25067
rect 3092 25033 3126 25067
rect 2306 24965 2340 24999
rect 2378 24965 2412 24999
rect 2450 24965 2484 24999
rect 2522 24965 2556 24999
rect 2594 24965 2628 24999
rect 2666 24965 2700 24999
rect 2737 24965 2771 24999
rect 2808 24965 2842 24999
rect 2879 24965 2913 24999
rect 2950 24965 2984 24999
rect 3021 24965 3055 24999
rect 3092 24965 3126 24999
rect 2306 24897 2340 24931
rect 2378 24897 2412 24931
rect 2450 24897 2484 24931
rect 2522 24897 2556 24931
rect 2594 24897 2628 24931
rect 2666 24897 2700 24931
rect 2737 24897 2771 24931
rect 2808 24897 2842 24931
rect 2879 24897 2913 24931
rect 2950 24897 2984 24931
rect 3021 24897 3055 24931
rect 3092 24897 3126 24931
rect 2306 24829 2340 24863
rect 2378 24829 2412 24863
rect 2450 24829 2484 24863
rect 2522 24829 2556 24863
rect 2594 24829 2628 24863
rect 2666 24829 2700 24863
rect 2737 24829 2771 24863
rect 2808 24829 2842 24863
rect 2879 24829 2913 24863
rect 2950 24829 2984 24863
rect 3021 24829 3055 24863
rect 3092 24829 3126 24863
rect 2306 24761 2340 24795
rect 2378 24761 2412 24795
rect 2450 24761 2484 24795
rect 2522 24761 2556 24795
rect 2594 24761 2628 24795
rect 2666 24761 2700 24795
rect 2737 24761 2771 24795
rect 2808 24761 2842 24795
rect 2879 24761 2913 24795
rect 2950 24761 2984 24795
rect 3021 24761 3055 24795
rect 3092 24761 3126 24795
rect 728 24658 762 24692
rect 796 24658 830 24692
rect 864 24658 898 24692
rect 932 24658 966 24692
rect 728 24589 762 24623
rect 796 24589 830 24623
rect 864 24589 898 24623
rect 932 24589 966 24623
rect 728 24520 762 24554
rect 796 24520 830 24554
rect 864 24520 898 24554
rect 932 24520 966 24554
rect 728 24451 762 24485
rect 796 24451 830 24485
rect 864 24451 898 24485
rect 932 24451 966 24485
rect 728 24382 762 24416
rect 796 24382 830 24416
rect 864 24382 898 24416
rect 932 24382 966 24416
rect 728 24313 762 24347
rect 796 24313 830 24347
rect 864 24313 898 24347
rect 932 24313 966 24347
rect 728 24244 762 24278
rect 796 24244 830 24278
rect 864 24244 898 24278
rect 932 24244 966 24278
rect 728 24175 762 24209
rect 796 24175 830 24209
rect 864 24175 898 24209
rect 932 24175 966 24209
rect 728 24106 762 24140
rect 796 24106 830 24140
rect 864 24106 898 24140
rect 932 24106 966 24140
rect 728 24037 762 24071
rect 796 24037 830 24071
rect 864 24037 898 24071
rect 932 24037 966 24071
rect 728 23968 762 24002
rect 796 23968 830 24002
rect 864 23968 898 24002
rect 932 23968 966 24002
rect 728 23899 762 23933
rect 796 23899 830 23933
rect 864 23899 898 23933
rect 932 23899 966 23933
rect 728 23830 762 23864
rect 796 23830 830 23864
rect 864 23830 898 23864
rect 932 23830 966 23864
rect 728 23761 762 23795
rect 796 23761 830 23795
rect 864 23761 898 23795
rect 932 23761 966 23795
rect 728 23692 762 23726
rect 796 23692 830 23726
rect 864 23692 898 23726
rect 932 23692 966 23726
rect 728 23623 762 23657
rect 796 23623 830 23657
rect 864 23623 898 23657
rect 932 23623 966 23657
rect 728 23554 762 23588
rect 796 23554 830 23588
rect 864 23554 898 23588
rect 932 23554 966 23588
rect 728 23485 762 23519
rect 796 23485 830 23519
rect 864 23485 898 23519
rect 932 23485 966 23519
rect 728 23416 762 23450
rect 796 23416 830 23450
rect 864 23416 898 23450
rect 932 23416 966 23450
rect 728 23347 762 23381
rect 796 23347 830 23381
rect 864 23347 898 23381
rect 932 23347 966 23381
rect 728 23278 762 23312
rect 796 23278 830 23312
rect 864 23278 898 23312
rect 932 23278 966 23312
rect 470 2154 504 2188
rect 538 2154 572 2188
rect 606 2154 640 2188
rect 1550 2154 1584 2188
rect 1618 2154 1652 2188
rect 1686 2154 1720 2188
<< mvnsubdiffcont >>
rect 2056 22995 2090 23029
rect 2056 22924 2090 22958
rect 2056 22853 2090 22887
rect 2056 22782 2090 22816
rect 2056 22710 2090 22744
rect 2056 22638 2090 22672
rect 2056 22566 2090 22600
rect 2056 22494 2090 22528
rect 2056 22422 2090 22456
rect 2056 22350 2090 22384
rect 2056 22278 2090 22312
rect 2710 16927 2744 16961
rect 2779 16927 2813 16961
rect 2848 16927 2882 16961
rect 2917 16927 2951 16961
rect 2986 16927 3020 16961
rect 3055 16927 3089 16961
rect 3124 16927 3158 16961
rect 3193 16927 3227 16961
rect 3262 16927 3296 16961
rect 3331 16927 3365 16961
rect 3400 16927 3434 16961
rect 3469 16927 3503 16961
rect 3538 16927 3572 16961
rect 3607 16927 3641 16961
rect 3676 16927 3710 16961
rect 3745 16927 3779 16961
rect 3814 16927 3848 16961
rect 3883 16927 3917 16961
rect 3952 16927 3986 16961
rect 4021 16927 4055 16961
rect 4090 16927 4124 16961
rect 4159 16927 4193 16961
rect 4228 16927 4262 16961
rect 4297 16927 4331 16961
rect 4366 16927 4400 16961
rect 4435 16927 4469 16961
rect 4504 16927 4538 16961
rect 4573 16927 4607 16961
rect 4642 16927 4676 16961
rect 4711 16927 4745 16961
rect 4780 16927 4814 16961
rect 4849 16927 4883 16961
rect 4918 16927 4952 16961
rect 4987 16927 5021 16961
rect 5056 16927 5090 16961
rect 5125 16927 5159 16961
rect 5194 16927 5228 16961
rect 5263 16927 5297 16961
rect 5332 16927 5366 16961
rect 5401 16927 5435 16961
rect 5470 16927 5504 16961
rect 5539 16927 5573 16961
rect 5608 16927 5642 16961
rect 5677 16927 5711 16961
rect 5746 16927 5780 16961
rect 5815 16927 5849 16961
rect 5884 16927 5918 16961
rect 5953 16927 5987 16961
rect 6022 16927 6056 16961
rect 2710 16859 2744 16893
rect 2779 16859 2813 16893
rect 2848 16859 2882 16893
rect 2917 16859 2951 16893
rect 2986 16859 3020 16893
rect 3055 16859 3089 16893
rect 3124 16859 3158 16893
rect 3193 16859 3227 16893
rect 3262 16859 3296 16893
rect 3331 16859 3365 16893
rect 3400 16859 3434 16893
rect 3469 16859 3503 16893
rect 3538 16859 3572 16893
rect 3607 16859 3641 16893
rect 3676 16859 3710 16893
rect 3745 16859 3779 16893
rect 3814 16859 3848 16893
rect 3883 16859 3917 16893
rect 3952 16859 3986 16893
rect 4021 16859 4055 16893
rect 4090 16859 4124 16893
rect 4159 16859 4193 16893
rect 4228 16859 4262 16893
rect 4297 16859 4331 16893
rect 4366 16859 4400 16893
rect 4435 16859 4469 16893
rect 4504 16859 4538 16893
rect 4573 16859 4607 16893
rect 4642 16859 4676 16893
rect 4711 16859 4745 16893
rect 4780 16859 4814 16893
rect 4849 16859 4883 16893
rect 4918 16859 4952 16893
rect 4987 16859 5021 16893
rect 5056 16859 5090 16893
rect 5125 16859 5159 16893
rect 5194 16859 5228 16893
rect 5263 16859 5297 16893
rect 5332 16859 5366 16893
rect 5401 16859 5435 16893
rect 5470 16859 5504 16893
rect 5539 16859 5573 16893
rect 5608 16859 5642 16893
rect 5677 16859 5711 16893
rect 5746 16859 5780 16893
rect 5815 16859 5849 16893
rect 5884 16859 5918 16893
rect 5953 16859 5987 16893
rect 6022 16859 6056 16893
rect 2710 16791 2744 16825
rect 2779 16791 2813 16825
rect 2848 16791 2882 16825
rect 2917 16791 2951 16825
rect 2986 16791 3020 16825
rect 3055 16791 3089 16825
rect 3124 16791 3158 16825
rect 3193 16791 3227 16825
rect 3262 16791 3296 16825
rect 3331 16791 3365 16825
rect 3400 16791 3434 16825
rect 3469 16791 3503 16825
rect 3538 16791 3572 16825
rect 3607 16791 3641 16825
rect 3676 16791 3710 16825
rect 3745 16791 3779 16825
rect 3814 16791 3848 16825
rect 3883 16791 3917 16825
rect 3952 16791 3986 16825
rect 4021 16791 4055 16825
rect 4090 16791 4124 16825
rect 4159 16791 4193 16825
rect 4228 16791 4262 16825
rect 4297 16791 4331 16825
rect 4366 16791 4400 16825
rect 4435 16791 4469 16825
rect 4504 16791 4538 16825
rect 4573 16791 4607 16825
rect 4642 16791 4676 16825
rect 4711 16791 4745 16825
rect 4780 16791 4814 16825
rect 4849 16791 4883 16825
rect 4918 16791 4952 16825
rect 4987 16791 5021 16825
rect 5056 16791 5090 16825
rect 5125 16791 5159 16825
rect 5194 16791 5228 16825
rect 5263 16791 5297 16825
rect 5332 16791 5366 16825
rect 5401 16791 5435 16825
rect 5470 16791 5504 16825
rect 5539 16791 5573 16825
rect 5608 16791 5642 16825
rect 5677 16791 5711 16825
rect 5746 16791 5780 16825
rect 5815 16791 5849 16825
rect 5884 16791 5918 16825
rect 5953 16791 5987 16825
rect 6022 16791 6056 16825
rect 2710 16723 2744 16757
rect 2779 16723 2813 16757
rect 2848 16723 2882 16757
rect 2917 16723 2951 16757
rect 2986 16723 3020 16757
rect 3055 16723 3089 16757
rect 3124 16723 3158 16757
rect 3193 16723 3227 16757
rect 3262 16723 3296 16757
rect 3331 16723 3365 16757
rect 3400 16723 3434 16757
rect 3469 16723 3503 16757
rect 3538 16723 3572 16757
rect 3607 16723 3641 16757
rect 3676 16723 3710 16757
rect 3745 16723 3779 16757
rect 3814 16723 3848 16757
rect 3883 16723 3917 16757
rect 3952 16723 3986 16757
rect 4021 16723 4055 16757
rect 4090 16723 4124 16757
rect 4159 16723 4193 16757
rect 4228 16723 4262 16757
rect 4297 16723 4331 16757
rect 4366 16723 4400 16757
rect 4435 16723 4469 16757
rect 4504 16723 4538 16757
rect 4573 16723 4607 16757
rect 4642 16723 4676 16757
rect 4711 16723 4745 16757
rect 4780 16723 4814 16757
rect 4849 16723 4883 16757
rect 4918 16723 4952 16757
rect 4987 16723 5021 16757
rect 5056 16723 5090 16757
rect 5125 16723 5159 16757
rect 5194 16723 5228 16757
rect 5263 16723 5297 16757
rect 5332 16723 5366 16757
rect 5401 16723 5435 16757
rect 5470 16723 5504 16757
rect 5539 16723 5573 16757
rect 5608 16723 5642 16757
rect 5677 16723 5711 16757
rect 5746 16723 5780 16757
rect 5815 16723 5849 16757
rect 5884 16723 5918 16757
rect 5953 16723 5987 16757
rect 6022 16723 6056 16757
rect 2710 16655 2744 16689
rect 2779 16655 2813 16689
rect 2848 16655 2882 16689
rect 2917 16655 2951 16689
rect 2986 16655 3020 16689
rect 3055 16655 3089 16689
rect 3124 16655 3158 16689
rect 3193 16655 3227 16689
rect 3262 16655 3296 16689
rect 3331 16655 3365 16689
rect 3400 16655 3434 16689
rect 3469 16655 3503 16689
rect 3538 16655 3572 16689
rect 3607 16655 3641 16689
rect 3676 16655 3710 16689
rect 3745 16655 3779 16689
rect 3814 16655 3848 16689
rect 3883 16655 3917 16689
rect 3952 16655 3986 16689
rect 4021 16655 4055 16689
rect 4090 16655 4124 16689
rect 4159 16655 4193 16689
rect 4228 16655 4262 16689
rect 4297 16655 4331 16689
rect 4366 16655 4400 16689
rect 4435 16655 4469 16689
rect 4504 16655 4538 16689
rect 4573 16655 4607 16689
rect 4642 16655 4676 16689
rect 4711 16655 4745 16689
rect 4780 16655 4814 16689
rect 4849 16655 4883 16689
rect 4918 16655 4952 16689
rect 4987 16655 5021 16689
rect 5056 16655 5090 16689
rect 5125 16655 5159 16689
rect 5194 16655 5228 16689
rect 5263 16655 5297 16689
rect 5332 16655 5366 16689
rect 5401 16655 5435 16689
rect 5470 16655 5504 16689
rect 5539 16655 5573 16689
rect 5608 16655 5642 16689
rect 5677 16655 5711 16689
rect 5746 16655 5780 16689
rect 5815 16655 5849 16689
rect 5884 16655 5918 16689
rect 5953 16655 5987 16689
rect 6022 16655 6056 16689
rect 2710 16587 2744 16621
rect 2779 16587 2813 16621
rect 2848 16587 2882 16621
rect 2917 16587 2951 16621
rect 2986 16587 3020 16621
rect 3055 16587 3089 16621
rect 3124 16587 3158 16621
rect 3193 16587 3227 16621
rect 3262 16587 3296 16621
rect 3331 16587 3365 16621
rect 3400 16587 3434 16621
rect 3469 16587 3503 16621
rect 3538 16587 3572 16621
rect 3607 16587 3641 16621
rect 3676 16587 3710 16621
rect 3745 16587 3779 16621
rect 3814 16587 3848 16621
rect 3883 16587 3917 16621
rect 3952 16587 3986 16621
rect 4021 16587 4055 16621
rect 4090 16587 4124 16621
rect 4159 16587 4193 16621
rect 4228 16587 4262 16621
rect 4297 16587 4331 16621
rect 4366 16587 4400 16621
rect 4435 16587 4469 16621
rect 4504 16587 4538 16621
rect 4573 16587 4607 16621
rect 4642 16587 4676 16621
rect 4711 16587 4745 16621
rect 4780 16587 4814 16621
rect 4849 16587 4883 16621
rect 4918 16587 4952 16621
rect 4987 16587 5021 16621
rect 5056 16587 5090 16621
rect 5125 16587 5159 16621
rect 5194 16587 5228 16621
rect 5263 16587 5297 16621
rect 5332 16587 5366 16621
rect 5401 16587 5435 16621
rect 5470 16587 5504 16621
rect 5539 16587 5573 16621
rect 5608 16587 5642 16621
rect 5677 16587 5711 16621
rect 5746 16587 5780 16621
rect 5815 16587 5849 16621
rect 5884 16587 5918 16621
rect 5953 16587 5987 16621
rect 6022 16587 6056 16621
rect 2710 16519 2744 16553
rect 2779 16519 2813 16553
rect 2848 16519 2882 16553
rect 2917 16519 2951 16553
rect 2986 16519 3020 16553
rect 3055 16519 3089 16553
rect 3124 16519 3158 16553
rect 3193 16519 3227 16553
rect 3262 16519 3296 16553
rect 3331 16519 3365 16553
rect 3400 16519 3434 16553
rect 3469 16519 3503 16553
rect 3538 16519 3572 16553
rect 3607 16519 3641 16553
rect 3676 16519 3710 16553
rect 3745 16519 3779 16553
rect 3814 16519 3848 16553
rect 3883 16519 3917 16553
rect 3952 16519 3986 16553
rect 4021 16519 4055 16553
rect 4090 16519 4124 16553
rect 4159 16519 4193 16553
rect 4228 16519 4262 16553
rect 4297 16519 4331 16553
rect 4366 16519 4400 16553
rect 4435 16519 4469 16553
rect 4504 16519 4538 16553
rect 4573 16519 4607 16553
rect 4642 16519 4676 16553
rect 4711 16519 4745 16553
rect 4780 16519 4814 16553
rect 4849 16519 4883 16553
rect 4918 16519 4952 16553
rect 4987 16519 5021 16553
rect 5056 16519 5090 16553
rect 5125 16519 5159 16553
rect 5194 16519 5228 16553
rect 5263 16519 5297 16553
rect 5332 16519 5366 16553
rect 5401 16519 5435 16553
rect 5470 16519 5504 16553
rect 5539 16519 5573 16553
rect 5608 16519 5642 16553
rect 5677 16519 5711 16553
rect 5746 16519 5780 16553
rect 5815 16519 5849 16553
rect 5884 16519 5918 16553
rect 5953 16519 5987 16553
rect 6022 16519 6056 16553
rect 2710 16451 2744 16485
rect 2779 16451 2813 16485
rect 2848 16451 2882 16485
rect 2917 16451 2951 16485
rect 2986 16451 3020 16485
rect 3055 16451 3089 16485
rect 3124 16451 3158 16485
rect 3193 16451 3227 16485
rect 3262 16451 3296 16485
rect 3331 16451 3365 16485
rect 3400 16451 3434 16485
rect 3469 16451 3503 16485
rect 3538 16451 3572 16485
rect 3607 16451 3641 16485
rect 3676 16451 3710 16485
rect 3745 16451 3779 16485
rect 3814 16451 3848 16485
rect 3883 16451 3917 16485
rect 3952 16451 3986 16485
rect 4021 16451 4055 16485
rect 4090 16451 4124 16485
rect 4159 16451 4193 16485
rect 4228 16451 4262 16485
rect 4297 16451 4331 16485
rect 4366 16451 4400 16485
rect 4435 16451 4469 16485
rect 4504 16451 4538 16485
rect 4573 16451 4607 16485
rect 4642 16451 4676 16485
rect 4711 16451 4745 16485
rect 4780 16451 4814 16485
rect 4849 16451 4883 16485
rect 4918 16451 4952 16485
rect 4987 16451 5021 16485
rect 5056 16451 5090 16485
rect 5125 16451 5159 16485
rect 5194 16451 5228 16485
rect 5263 16451 5297 16485
rect 5332 16451 5366 16485
rect 5401 16451 5435 16485
rect 5470 16451 5504 16485
rect 5539 16451 5573 16485
rect 5608 16451 5642 16485
rect 5677 16451 5711 16485
rect 5746 16451 5780 16485
rect 5815 16451 5849 16485
rect 5884 16451 5918 16485
rect 5953 16451 5987 16485
rect 6022 16451 6056 16485
rect 6091 16451 17005 16961
rect -2732 16145 -2698 16179
rect -2663 16145 -2629 16179
rect -2594 16145 -2560 16179
rect -2525 16145 -2491 16179
rect -2456 16145 -2422 16179
rect -2387 16145 -2353 16179
rect -2318 16145 -2284 16179
rect -2249 16145 -2215 16179
rect -2180 16145 -2146 16179
rect -2111 16145 -2077 16179
rect -2042 16145 -2008 16179
rect -1973 16145 -1939 16179
rect -1904 16145 -1870 16179
rect -1835 16145 -1801 16179
rect -1766 16145 -1732 16179
rect -1697 16145 -1663 16179
rect -1628 16145 -1594 16179
rect -1559 16145 -1525 16179
rect -1490 16145 -1456 16179
rect -1421 16145 -1387 16179
rect -1352 16145 -1318 16179
rect -1283 16145 -1249 16179
rect -1214 16145 -1180 16179
rect -1145 16145 -1111 16179
rect -1076 16145 -1042 16179
rect -1007 16145 -973 16179
rect -938 16145 -904 16179
rect -869 16145 -835 16179
rect -800 16145 -766 16179
rect -731 16145 -697 16179
rect -662 16145 -628 16179
rect -593 16145 -559 16179
rect -524 16145 -490 16179
rect -455 16145 -421 16179
rect -386 16145 -352 16179
rect -317 16145 -283 16179
rect -248 16145 -214 16179
rect -179 16145 -145 16179
rect -110 16145 -76 16179
rect -41 16145 -7 16179
rect 28 16145 62 16179
rect 97 16145 131 16179
rect 166 16145 200 16179
rect 235 16145 269 16179
rect 304 16145 338 16179
rect 373 16145 407 16179
rect 442 16145 476 16179
rect 511 16145 545 16179
rect 580 16145 614 16179
rect 649 16145 683 16179
rect -2732 16077 -2698 16111
rect -2663 16077 -2629 16111
rect -2594 16077 -2560 16111
rect -2525 16077 -2491 16111
rect -2456 16077 -2422 16111
rect -2387 16077 -2353 16111
rect -2318 16077 -2284 16111
rect -2249 16077 -2215 16111
rect -2180 16077 -2146 16111
rect -2111 16077 -2077 16111
rect -2042 16077 -2008 16111
rect -1973 16077 -1939 16111
rect -1904 16077 -1870 16111
rect -1835 16077 -1801 16111
rect -1766 16077 -1732 16111
rect -1697 16077 -1663 16111
rect -1628 16077 -1594 16111
rect -1559 16077 -1525 16111
rect -1490 16077 -1456 16111
rect -1421 16077 -1387 16111
rect -1352 16077 -1318 16111
rect -1283 16077 -1249 16111
rect -1214 16077 -1180 16111
rect -1145 16077 -1111 16111
rect -1076 16077 -1042 16111
rect -1007 16077 -973 16111
rect -938 16077 -904 16111
rect -869 16077 -835 16111
rect -800 16077 -766 16111
rect -731 16077 -697 16111
rect -662 16077 -628 16111
rect -593 16077 -559 16111
rect -524 16077 -490 16111
rect -455 16077 -421 16111
rect -386 16077 -352 16111
rect -317 16077 -283 16111
rect -248 16077 -214 16111
rect -179 16077 -145 16111
rect -110 16077 -76 16111
rect -41 16077 -7 16111
rect 28 16077 62 16111
rect 97 16077 131 16111
rect 166 16077 200 16111
rect 235 16077 269 16111
rect 304 16077 338 16111
rect 373 16077 407 16111
rect 442 16077 476 16111
rect 511 16077 545 16111
rect 580 16077 614 16111
rect 649 16077 683 16111
rect -2732 16009 -2698 16043
rect -2663 16009 -2629 16043
rect -2594 16009 -2560 16043
rect -2525 16009 -2491 16043
rect -2456 16009 -2422 16043
rect -2387 16009 -2353 16043
rect -2318 16009 -2284 16043
rect -2249 16009 -2215 16043
rect -2180 16009 -2146 16043
rect -2111 16009 -2077 16043
rect -2042 16009 -2008 16043
rect -1973 16009 -1939 16043
rect -1904 16009 -1870 16043
rect -1835 16009 -1801 16043
rect -1766 16009 -1732 16043
rect -1697 16009 -1663 16043
rect -1628 16009 -1594 16043
rect -1559 16009 -1525 16043
rect -1490 16009 -1456 16043
rect -1421 16009 -1387 16043
rect -1352 16009 -1318 16043
rect -1283 16009 -1249 16043
rect -1214 16009 -1180 16043
rect -1145 16009 -1111 16043
rect -1076 16009 -1042 16043
rect -1007 16009 -973 16043
rect -938 16009 -904 16043
rect -869 16009 -835 16043
rect -800 16009 -766 16043
rect -731 16009 -697 16043
rect -662 16009 -628 16043
rect -593 16009 -559 16043
rect -524 16009 -490 16043
rect -455 16009 -421 16043
rect -386 16009 -352 16043
rect -317 16009 -283 16043
rect -248 16009 -214 16043
rect -179 16009 -145 16043
rect -110 16009 -76 16043
rect -41 16009 -7 16043
rect 28 16009 62 16043
rect 97 16009 131 16043
rect 166 16009 200 16043
rect 235 16009 269 16043
rect 304 16009 338 16043
rect 373 16009 407 16043
rect 442 16009 476 16043
rect 511 16009 545 16043
rect 580 16009 614 16043
rect 649 16009 683 16043
rect -2732 15941 -2698 15975
rect -2663 15941 -2629 15975
rect -2594 15941 -2560 15975
rect -2525 15941 -2491 15975
rect -2456 15941 -2422 15975
rect -2387 15941 -2353 15975
rect -2318 15941 -2284 15975
rect -2249 15941 -2215 15975
rect -2180 15941 -2146 15975
rect -2111 15941 -2077 15975
rect -2042 15941 -2008 15975
rect -1973 15941 -1939 15975
rect -1904 15941 -1870 15975
rect -1835 15941 -1801 15975
rect -1766 15941 -1732 15975
rect -1697 15941 -1663 15975
rect -1628 15941 -1594 15975
rect -1559 15941 -1525 15975
rect -1490 15941 -1456 15975
rect -1421 15941 -1387 15975
rect -1352 15941 -1318 15975
rect -1283 15941 -1249 15975
rect -1214 15941 -1180 15975
rect -1145 15941 -1111 15975
rect -1076 15941 -1042 15975
rect -1007 15941 -973 15975
rect -938 15941 -904 15975
rect -869 15941 -835 15975
rect -800 15941 -766 15975
rect -731 15941 -697 15975
rect -662 15941 -628 15975
rect -593 15941 -559 15975
rect -524 15941 -490 15975
rect -455 15941 -421 15975
rect -386 15941 -352 15975
rect -317 15941 -283 15975
rect -248 15941 -214 15975
rect -179 15941 -145 15975
rect -110 15941 -76 15975
rect -41 15941 -7 15975
rect 28 15941 62 15975
rect 97 15941 131 15975
rect 166 15941 200 15975
rect 235 15941 269 15975
rect 304 15941 338 15975
rect 373 15941 407 15975
rect 442 15941 476 15975
rect 511 15941 545 15975
rect 580 15941 614 15975
rect 649 15941 683 15975
rect -2732 15873 -2698 15907
rect -2663 15873 -2629 15907
rect -2594 15873 -2560 15907
rect -2525 15873 -2491 15907
rect -2456 15873 -2422 15907
rect -2387 15873 -2353 15907
rect -2318 15873 -2284 15907
rect -2249 15873 -2215 15907
rect -2180 15873 -2146 15907
rect -2111 15873 -2077 15907
rect -2042 15873 -2008 15907
rect -1973 15873 -1939 15907
rect -1904 15873 -1870 15907
rect -1835 15873 -1801 15907
rect -1766 15873 -1732 15907
rect -1697 15873 -1663 15907
rect -1628 15873 -1594 15907
rect -1559 15873 -1525 15907
rect -1490 15873 -1456 15907
rect -1421 15873 -1387 15907
rect -1352 15873 -1318 15907
rect -1283 15873 -1249 15907
rect -1214 15873 -1180 15907
rect -1145 15873 -1111 15907
rect -1076 15873 -1042 15907
rect -1007 15873 -973 15907
rect -938 15873 -904 15907
rect -869 15873 -835 15907
rect -800 15873 -766 15907
rect -731 15873 -697 15907
rect -662 15873 -628 15907
rect -593 15873 -559 15907
rect -524 15873 -490 15907
rect -455 15873 -421 15907
rect -386 15873 -352 15907
rect -317 15873 -283 15907
rect -248 15873 -214 15907
rect -179 15873 -145 15907
rect -110 15873 -76 15907
rect -41 15873 -7 15907
rect 28 15873 62 15907
rect 97 15873 131 15907
rect 166 15873 200 15907
rect 235 15873 269 15907
rect 304 15873 338 15907
rect 373 15873 407 15907
rect 442 15873 476 15907
rect 511 15873 545 15907
rect 580 15873 614 15907
rect 649 15873 683 15907
rect -2732 15805 -2698 15839
rect -2663 15805 -2629 15839
rect -2594 15805 -2560 15839
rect -2525 15805 -2491 15839
rect -2456 15805 -2422 15839
rect -2387 15805 -2353 15839
rect -2318 15805 -2284 15839
rect -2249 15805 -2215 15839
rect -2180 15805 -2146 15839
rect -2111 15805 -2077 15839
rect -2042 15805 -2008 15839
rect -1973 15805 -1939 15839
rect -1904 15805 -1870 15839
rect -1835 15805 -1801 15839
rect -1766 15805 -1732 15839
rect -1697 15805 -1663 15839
rect -1628 15805 -1594 15839
rect -1559 15805 -1525 15839
rect -1490 15805 -1456 15839
rect -1421 15805 -1387 15839
rect -1352 15805 -1318 15839
rect -1283 15805 -1249 15839
rect -1214 15805 -1180 15839
rect -1145 15805 -1111 15839
rect -1076 15805 -1042 15839
rect -1007 15805 -973 15839
rect -938 15805 -904 15839
rect -869 15805 -835 15839
rect -800 15805 -766 15839
rect -731 15805 -697 15839
rect -662 15805 -628 15839
rect -593 15805 -559 15839
rect -524 15805 -490 15839
rect -455 15805 -421 15839
rect -386 15805 -352 15839
rect -317 15805 -283 15839
rect -248 15805 -214 15839
rect -179 15805 -145 15839
rect -110 15805 -76 15839
rect -41 15805 -7 15839
rect 28 15805 62 15839
rect 97 15805 131 15839
rect 166 15805 200 15839
rect 235 15805 269 15839
rect 304 15805 338 15839
rect 373 15805 407 15839
rect 442 15805 476 15839
rect 511 15805 545 15839
rect 580 15805 614 15839
rect 649 15805 683 15839
rect -2732 15737 -2698 15771
rect -2663 15737 -2629 15771
rect -2594 15737 -2560 15771
rect -2525 15737 -2491 15771
rect -2456 15737 -2422 15771
rect -2387 15737 -2353 15771
rect -2318 15737 -2284 15771
rect -2249 15737 -2215 15771
rect -2180 15737 -2146 15771
rect -2111 15737 -2077 15771
rect -2042 15737 -2008 15771
rect -1973 15737 -1939 15771
rect -1904 15737 -1870 15771
rect -1835 15737 -1801 15771
rect -1766 15737 -1732 15771
rect -1697 15737 -1663 15771
rect -1628 15737 -1594 15771
rect -1559 15737 -1525 15771
rect -1490 15737 -1456 15771
rect -1421 15737 -1387 15771
rect -1352 15737 -1318 15771
rect -1283 15737 -1249 15771
rect -1214 15737 -1180 15771
rect -1145 15737 -1111 15771
rect -1076 15737 -1042 15771
rect -1007 15737 -973 15771
rect -938 15737 -904 15771
rect -869 15737 -835 15771
rect -800 15737 -766 15771
rect -731 15737 -697 15771
rect -662 15737 -628 15771
rect -593 15737 -559 15771
rect -524 15737 -490 15771
rect -455 15737 -421 15771
rect -386 15737 -352 15771
rect -317 15737 -283 15771
rect -248 15737 -214 15771
rect -179 15737 -145 15771
rect -110 15737 -76 15771
rect -41 15737 -7 15771
rect 28 15737 62 15771
rect 97 15737 131 15771
rect 166 15737 200 15771
rect 235 15737 269 15771
rect 304 15737 338 15771
rect 373 15737 407 15771
rect 442 15737 476 15771
rect 511 15737 545 15771
rect 580 15737 614 15771
rect 649 15737 683 15771
rect -2732 15669 -2698 15703
rect -2663 15669 -2629 15703
rect -2594 15669 -2560 15703
rect -2525 15669 -2491 15703
rect -2456 15669 -2422 15703
rect -2387 15669 -2353 15703
rect -2318 15669 -2284 15703
rect -2249 15669 -2215 15703
rect -2180 15669 -2146 15703
rect -2111 15669 -2077 15703
rect -2042 15669 -2008 15703
rect -1973 15669 -1939 15703
rect -1904 15669 -1870 15703
rect -1835 15669 -1801 15703
rect -1766 15669 -1732 15703
rect -1697 15669 -1663 15703
rect -1628 15669 -1594 15703
rect -1559 15669 -1525 15703
rect -1490 15669 -1456 15703
rect -1421 15669 -1387 15703
rect -1352 15669 -1318 15703
rect -1283 15669 -1249 15703
rect -1214 15669 -1180 15703
rect -1145 15669 -1111 15703
rect -1076 15669 -1042 15703
rect -1007 15669 -973 15703
rect -938 15669 -904 15703
rect -869 15669 -835 15703
rect -800 15669 -766 15703
rect -731 15669 -697 15703
rect -662 15669 -628 15703
rect -593 15669 -559 15703
rect -524 15669 -490 15703
rect -455 15669 -421 15703
rect -386 15669 -352 15703
rect -317 15669 -283 15703
rect -248 15669 -214 15703
rect -179 15669 -145 15703
rect -110 15669 -76 15703
rect -41 15669 -7 15703
rect 28 15669 62 15703
rect 97 15669 131 15703
rect 166 15669 200 15703
rect 235 15669 269 15703
rect 304 15669 338 15703
rect 373 15669 407 15703
rect 442 15669 476 15703
rect 511 15669 545 15703
rect 580 15669 614 15703
rect 649 15669 683 15703
rect -2732 15601 -2698 15635
rect -2663 15601 -2629 15635
rect -2594 15601 -2560 15635
rect -2525 15601 -2491 15635
rect -2456 15601 -2422 15635
rect -2387 15601 -2353 15635
rect -2318 15601 -2284 15635
rect -2249 15601 -2215 15635
rect -2180 15601 -2146 15635
rect -2111 15601 -2077 15635
rect -2042 15601 -2008 15635
rect -1973 15601 -1939 15635
rect -1904 15601 -1870 15635
rect -1835 15601 -1801 15635
rect -1766 15601 -1732 15635
rect -1697 15601 -1663 15635
rect -1628 15601 -1594 15635
rect -1559 15601 -1525 15635
rect -1490 15601 -1456 15635
rect -1421 15601 -1387 15635
rect -1352 15601 -1318 15635
rect -1283 15601 -1249 15635
rect -1214 15601 -1180 15635
rect -1145 15601 -1111 15635
rect -1076 15601 -1042 15635
rect -1007 15601 -973 15635
rect -938 15601 -904 15635
rect -869 15601 -835 15635
rect -800 15601 -766 15635
rect -731 15601 -697 15635
rect -662 15601 -628 15635
rect -593 15601 -559 15635
rect -524 15601 -490 15635
rect -455 15601 -421 15635
rect -386 15601 -352 15635
rect -317 15601 -283 15635
rect -248 15601 -214 15635
rect -179 15601 -145 15635
rect -110 15601 -76 15635
rect -41 15601 -7 15635
rect 28 15601 62 15635
rect 97 15601 131 15635
rect 166 15601 200 15635
rect 235 15601 269 15635
rect 304 15601 338 15635
rect 373 15601 407 15635
rect 442 15601 476 15635
rect 511 15601 545 15635
rect 580 15601 614 15635
rect 649 15601 683 15635
rect -2732 15533 -2698 15567
rect -2663 15533 -2629 15567
rect -2594 15533 -2560 15567
rect -2525 15533 -2491 15567
rect -2456 15533 -2422 15567
rect -2387 15533 -2353 15567
rect -2318 15533 -2284 15567
rect -2249 15533 -2215 15567
rect -2180 15533 -2146 15567
rect -2111 15533 -2077 15567
rect -2042 15533 -2008 15567
rect -1973 15533 -1939 15567
rect -1904 15533 -1870 15567
rect -1835 15533 -1801 15567
rect -1766 15533 -1732 15567
rect -1697 15533 -1663 15567
rect -1628 15533 -1594 15567
rect -1559 15533 -1525 15567
rect -1490 15533 -1456 15567
rect -1421 15533 -1387 15567
rect -1352 15533 -1318 15567
rect -1283 15533 -1249 15567
rect -1214 15533 -1180 15567
rect -1145 15533 -1111 15567
rect -1076 15533 -1042 15567
rect -1007 15533 -973 15567
rect -938 15533 -904 15567
rect -869 15533 -835 15567
rect -800 15533 -766 15567
rect -731 15533 -697 15567
rect -662 15533 -628 15567
rect -593 15533 -559 15567
rect -524 15533 -490 15567
rect -455 15533 -421 15567
rect -386 15533 -352 15567
rect -317 15533 -283 15567
rect -248 15533 -214 15567
rect -179 15533 -145 15567
rect -110 15533 -76 15567
rect -41 15533 -7 15567
rect 28 15533 62 15567
rect 97 15533 131 15567
rect 166 15533 200 15567
rect 235 15533 269 15567
rect 304 15533 338 15567
rect 373 15533 407 15567
rect 442 15533 476 15567
rect 511 15533 545 15567
rect 580 15533 614 15567
rect 649 15533 683 15567
rect -2732 15465 -2698 15499
rect -2663 15465 -2629 15499
rect -2594 15465 -2560 15499
rect -2525 15465 -2491 15499
rect -2456 15465 -2422 15499
rect -2387 15465 -2353 15499
rect -2318 15465 -2284 15499
rect -2249 15465 -2215 15499
rect -2180 15465 -2146 15499
rect -2111 15465 -2077 15499
rect -2042 15465 -2008 15499
rect -1973 15465 -1939 15499
rect -1904 15465 -1870 15499
rect -1835 15465 -1801 15499
rect -1766 15465 -1732 15499
rect -1697 15465 -1663 15499
rect -1628 15465 -1594 15499
rect -1559 15465 -1525 15499
rect -1490 15465 -1456 15499
rect -1421 15465 -1387 15499
rect -1352 15465 -1318 15499
rect -1283 15465 -1249 15499
rect -1214 15465 -1180 15499
rect -1145 15465 -1111 15499
rect -1076 15465 -1042 15499
rect -1007 15465 -973 15499
rect -938 15465 -904 15499
rect -869 15465 -835 15499
rect -800 15465 -766 15499
rect -731 15465 -697 15499
rect -662 15465 -628 15499
rect -593 15465 -559 15499
rect -524 15465 -490 15499
rect -455 15465 -421 15499
rect -386 15465 -352 15499
rect -317 15465 -283 15499
rect -248 15465 -214 15499
rect -179 15465 -145 15499
rect -110 15465 -76 15499
rect -41 15465 -7 15499
rect 28 15465 62 15499
rect 97 15465 131 15499
rect 166 15465 200 15499
rect 235 15465 269 15499
rect 304 15465 338 15499
rect 373 15465 407 15499
rect 442 15465 476 15499
rect 511 15465 545 15499
rect 580 15465 614 15499
rect 649 15465 683 15499
rect -2732 15397 -2698 15431
rect -2663 15397 -2629 15431
rect -2594 15397 -2560 15431
rect -2525 15397 -2491 15431
rect -2456 15397 -2422 15431
rect -2387 15397 -2353 15431
rect -2318 15397 -2284 15431
rect -2249 15397 -2215 15431
rect -2180 15397 -2146 15431
rect -2111 15397 -2077 15431
rect -2042 15397 -2008 15431
rect -1973 15397 -1939 15431
rect -1904 15397 -1870 15431
rect -1835 15397 -1801 15431
rect -1766 15397 -1732 15431
rect -1697 15397 -1663 15431
rect -1628 15397 -1594 15431
rect -1559 15397 -1525 15431
rect -1490 15397 -1456 15431
rect -1421 15397 -1387 15431
rect -1352 15397 -1318 15431
rect -1283 15397 -1249 15431
rect -1214 15397 -1180 15431
rect -1145 15397 -1111 15431
rect -1076 15397 -1042 15431
rect -1007 15397 -973 15431
rect -938 15397 -904 15431
rect -869 15397 -835 15431
rect -800 15397 -766 15431
rect -731 15397 -697 15431
rect -662 15397 -628 15431
rect -593 15397 -559 15431
rect -524 15397 -490 15431
rect -455 15397 -421 15431
rect -386 15397 -352 15431
rect -317 15397 -283 15431
rect -248 15397 -214 15431
rect -179 15397 -145 15431
rect -110 15397 -76 15431
rect -41 15397 -7 15431
rect 28 15397 62 15431
rect 97 15397 131 15431
rect 166 15397 200 15431
rect 235 15397 269 15431
rect 304 15397 338 15431
rect 373 15397 407 15431
rect 442 15397 476 15431
rect 511 15397 545 15431
rect 580 15397 614 15431
rect 649 15397 683 15431
rect 718 15397 17004 16179
rect 138 3414 172 3448
rect 206 3414 240 3448
rect 274 3414 308 3448
rect 138 3344 172 3378
rect 206 3344 240 3378
rect 274 3344 308 3378
rect 138 3274 172 3308
rect 206 3274 240 3308
rect 274 3274 308 3308
rect 138 3204 172 3238
rect 206 3204 240 3238
rect 274 3204 308 3238
rect 138 3134 172 3168
rect 206 3134 240 3168
rect 274 3134 308 3168
rect 138 3064 172 3098
rect 206 3064 240 3098
rect 274 3064 308 3098
rect 138 2994 172 3028
rect 206 2994 240 3028
rect 274 2994 308 3028
rect 138 2924 172 2958
rect 206 2924 240 2958
rect 274 2924 308 2958
rect 138 2854 172 2888
rect 206 2854 240 2888
rect 274 2854 308 2888
rect 138 2784 172 2818
rect 206 2784 240 2818
rect 274 2784 308 2818
rect 138 2715 172 2749
rect 206 2715 240 2749
rect 274 2714 308 2748
rect 138 2646 172 2680
rect 206 2646 240 2680
rect 274 2644 308 2678
rect 138 2577 172 2611
rect 206 2577 240 2611
rect 274 2575 308 2609
rect 138 2508 172 2542
rect 206 2508 240 2542
rect 274 2506 308 2540
rect 138 2439 172 2473
rect 206 2439 240 2473
rect 274 2437 308 2471
rect 138 2370 172 2404
rect 206 2370 240 2404
rect 274 2368 308 2402
rect 138 2301 172 2335
rect 206 2301 240 2335
rect 274 2299 308 2333
rect 138 2232 172 2266
rect 206 2232 240 2266
rect 274 2230 308 2264
rect 1873 3414 1907 3448
rect 1941 3414 1975 3448
rect 2009 3414 2043 3448
rect 1873 3345 1907 3379
rect 1941 3345 1975 3379
rect 2009 3345 2043 3379
rect 1873 3276 1907 3310
rect 1941 3276 1975 3310
rect 2009 3276 2043 3310
rect 1873 3207 1907 3241
rect 1941 3207 1975 3241
rect 2009 3207 2043 3241
rect 1873 3138 1907 3172
rect 1941 3138 1975 3172
rect 2009 3138 2043 3172
rect 1873 3069 1907 3103
rect 1941 3069 1975 3103
rect 2009 3069 2043 3103
rect 1873 3000 1907 3034
rect 1941 3000 1975 3034
rect 2009 3000 2043 3034
rect 1873 2931 1907 2965
rect 1941 2931 1975 2965
rect 2009 2931 2043 2965
rect 1873 2862 1907 2896
rect 1941 2862 1975 2896
rect 2009 2862 2043 2896
rect 1873 2793 1907 2827
rect 1941 2793 1975 2827
rect 2009 2793 2043 2827
rect 1873 2724 1907 2758
rect 1941 2724 1975 2758
rect 2009 2724 2043 2758
rect 1873 2655 1907 2689
rect 1941 2655 1975 2689
rect 2009 2655 2043 2689
rect 1873 2586 1907 2620
rect 1941 2586 1975 2620
rect 2009 2586 2043 2620
rect 1873 2517 1907 2551
rect 1941 2517 1975 2551
rect 2009 2517 2043 2551
rect 1873 2448 1907 2482
rect 1941 2448 1975 2482
rect 2009 2448 2043 2482
rect 1873 2379 1907 2413
rect 1941 2379 1975 2413
rect 2009 2379 2043 2413
rect 1873 2310 1907 2344
rect 1941 2310 1975 2344
rect 2009 2310 2043 2344
rect 1873 2241 1907 2275
rect 1941 2241 1975 2275
rect 2009 2241 2043 2275
rect 138 2163 172 2197
rect 206 2163 240 2197
rect 274 2161 308 2195
rect 138 2094 172 2128
rect 206 2094 240 2128
rect 274 2092 308 2126
rect 138 2025 172 2059
rect 206 2025 240 2059
rect 274 2023 308 2057
rect 138 1956 172 1990
rect 206 1956 240 1990
rect 274 1954 308 1988
rect 138 1887 172 1921
rect 206 1887 240 1921
rect 274 1885 308 1919
rect 138 1818 172 1852
rect 206 1818 240 1852
rect 274 1816 308 1850
rect 138 1749 172 1783
rect 206 1749 240 1783
rect 274 1747 308 1781
rect 138 1680 172 1714
rect 206 1680 240 1714
rect 274 1678 308 1712
rect 138 1611 172 1645
rect 206 1611 240 1645
rect 274 1609 308 1643
rect 138 1542 172 1576
rect 206 1542 240 1576
rect 274 1540 308 1574
rect 138 1473 172 1507
rect 206 1473 240 1507
rect 274 1471 308 1505
rect 138 1404 172 1438
rect 206 1404 240 1438
rect 274 1402 308 1436
rect 138 1335 172 1369
rect 206 1335 240 1369
rect 274 1333 308 1367
rect 1873 2172 1907 2206
rect 1941 2172 1975 2206
rect 2009 2172 2043 2206
rect 1873 2103 1907 2137
rect 1941 2103 1975 2137
rect 2009 2103 2043 2137
rect 1873 2034 1907 2068
rect 1941 2034 1975 2068
rect 2009 2034 2043 2068
rect 1873 1965 1907 1999
rect 1941 1965 1975 1999
rect 2009 1965 2043 1999
rect 1873 1896 1907 1930
rect 1941 1896 1975 1930
rect 2009 1896 2043 1930
rect 1873 1826 1907 1860
rect 1941 1827 1975 1861
rect 2009 1827 2043 1861
rect 1873 1756 1907 1790
rect 1941 1758 1975 1792
rect 2009 1758 2043 1792
rect 1873 1686 1907 1720
rect 1941 1688 1975 1722
rect 2009 1688 2043 1722
rect 1873 1616 1907 1650
rect 1941 1618 1975 1652
rect 2009 1618 2043 1652
rect 1873 1546 1907 1580
rect 1941 1548 1975 1582
rect 2009 1548 2043 1582
rect 1873 1476 1907 1510
rect 1941 1478 1975 1512
rect 2009 1478 2043 1512
rect 1873 1406 1907 1440
rect 1941 1408 1975 1442
rect 2009 1408 2043 1442
rect 1873 1336 1907 1370
rect 1941 1338 1975 1372
rect 2009 1338 2043 1372
rect 138 1266 172 1300
rect 206 1266 240 1300
rect 274 1264 308 1298
rect 138 1197 172 1231
rect 206 1197 240 1231
rect 274 1195 308 1229
rect 138 1128 172 1162
rect 206 1128 240 1162
rect 1873 1266 1907 1300
rect 1941 1268 1975 1302
rect 2009 1268 2043 1302
rect 1873 1196 1907 1230
rect 1941 1198 1975 1232
rect 2009 1198 2043 1232
rect 274 1126 308 1160
rect 344 1126 378 1160
rect 414 1126 448 1160
rect 484 1126 518 1160
rect 554 1126 588 1160
rect 624 1126 658 1160
rect 694 1126 728 1160
rect 764 1126 798 1160
rect 834 1126 868 1160
rect 904 1126 938 1160
rect 974 1126 1008 1160
rect 1044 1126 1078 1160
rect 1114 1126 1148 1160
rect 1183 1126 1217 1160
rect 1252 1126 1286 1160
rect 1321 1126 1355 1160
rect 1390 1126 1424 1160
rect 1459 1126 1493 1160
rect 1528 1126 1562 1160
rect 1597 1126 1631 1160
rect 1666 1126 1700 1160
rect 1735 1126 1769 1160
rect 1804 1126 1838 1160
rect 1873 1126 1907 1160
rect 1941 1128 1975 1162
rect 2009 1128 2043 1162
rect 138 1059 172 1093
rect 206 1058 240 1092
rect 276 1058 310 1092
rect 346 1058 380 1092
rect 416 1058 450 1092
rect 486 1058 520 1092
rect 556 1058 590 1092
rect 626 1058 660 1092
rect 696 1058 730 1092
rect 766 1058 800 1092
rect 836 1058 870 1092
rect 905 1058 939 1092
rect 974 1058 1008 1092
rect 1043 1058 1077 1092
rect 1112 1058 1146 1092
rect 1181 1058 1215 1092
rect 1250 1058 1284 1092
rect 1319 1058 1353 1092
rect 1388 1058 1422 1092
rect 1457 1058 1491 1092
rect 1526 1058 1560 1092
rect 1595 1058 1629 1092
rect 1664 1058 1698 1092
rect 1733 1058 1767 1092
rect 1802 1058 1836 1092
rect 1871 1058 1905 1092
rect 1941 1058 1975 1092
rect 2009 1058 2043 1092
rect 206 990 240 1024
rect 276 990 310 1024
rect 346 990 380 1024
rect 416 990 450 1024
rect 486 990 520 1024
rect 556 990 590 1024
rect 626 990 660 1024
rect 696 990 730 1024
rect 766 990 800 1024
rect 836 990 870 1024
rect 905 990 939 1024
rect 974 990 1008 1024
rect 1043 990 1077 1024
rect 1112 990 1146 1024
rect 1181 990 1215 1024
rect 1250 990 1284 1024
rect 1319 990 1353 1024
rect 1388 990 1422 1024
rect 1457 990 1491 1024
rect 1526 990 1560 1024
rect 1595 990 1629 1024
rect 1664 990 1698 1024
rect 1733 990 1767 1024
rect 1802 990 1836 1024
rect 1871 990 1905 1024
rect 1940 990 1974 1024
<< poly >>
rect 872 22886 944 22903
rect 872 22852 888 22886
rect 922 22852 944 22886
rect 872 22803 944 22852
rect 872 22791 938 22803
rect 872 22757 888 22791
rect 922 22757 938 22791
rect 872 22747 938 22757
rect 872 22697 944 22747
rect 872 22663 888 22697
rect 922 22663 944 22697
rect 872 22647 944 22663
rect 872 22499 938 22515
rect 872 22465 888 22499
rect 922 22481 938 22499
rect 922 22465 944 22481
rect 872 22431 944 22465
rect 872 22397 888 22431
rect 922 22397 944 22431
rect 872 22381 944 22397
rect 234 18728 634 18744
rect 234 18694 281 18728
rect 315 18694 349 18728
rect 383 18694 417 18728
rect 451 18694 485 18728
rect 519 18694 553 18728
rect 587 18694 634 18728
rect 234 18665 634 18694
rect 234 16536 634 16565
rect 234 16502 281 16536
rect 315 16502 349 16536
rect 383 16502 417 16536
rect 451 16502 485 16536
rect 519 16502 553 16536
rect 587 16502 634 16536
rect 234 16486 634 16502
rect 672 2092 738 2108
rect 672 2058 688 2092
rect 722 2058 738 2092
rect 672 2024 738 2058
rect 672 1990 688 2024
rect 722 1990 738 2024
rect 672 1956 738 1990
rect 672 1922 688 1956
rect 722 1922 738 1956
rect 672 1906 738 1922
rect 672 1713 738 1729
rect 672 1679 688 1713
rect 722 1679 738 1713
rect 672 1645 738 1679
rect 672 1611 688 1645
rect 722 1611 738 1645
rect 672 1595 738 1611
<< polycont >>
rect 888 22852 922 22886
rect 888 22757 922 22791
rect 888 22663 922 22697
rect 888 22465 922 22499
rect 888 22397 922 22431
rect 281 18694 315 18728
rect 349 18694 383 18728
rect 417 18694 451 18728
rect 485 18694 519 18728
rect 553 18694 587 18728
rect 281 16502 315 16536
rect 349 16502 383 16536
rect 417 16502 451 16536
rect 485 16502 519 16536
rect 553 16502 587 16536
rect 688 2058 722 2092
rect 688 1990 722 2024
rect 688 1922 722 1956
rect 688 1679 722 1713
rect 688 1611 722 1645
<< locali >>
rect 664 25543 3248 25594
rect 664 25533 2306 25543
rect 2340 25533 2378 25543
rect 2412 25533 2450 25543
rect 664 25513 2297 25533
rect 664 25492 728 25513
rect 966 25499 2297 25513
rect 2340 25509 2373 25533
rect 2412 25509 2449 25533
rect 2484 25509 2522 25543
rect 2556 25533 2594 25543
rect 2628 25533 2666 25543
rect 2700 25533 2737 25543
rect 2771 25533 2808 25543
rect 2842 25533 2879 25543
rect 2913 25533 2950 25543
rect 2984 25533 3021 25543
rect 3055 25533 3092 25543
rect 2559 25509 2594 25533
rect 2635 25509 2666 25533
rect 2711 25509 2737 25533
rect 2787 25509 2808 25533
rect 2863 25509 2879 25533
rect 2938 25509 2950 25533
rect 3013 25509 3021 25533
rect 3088 25509 3092 25533
rect 3126 25533 3248 25543
rect 3126 25509 3129 25533
rect 2331 25499 2373 25509
rect 2407 25499 2449 25509
rect 2483 25499 2525 25509
rect 2559 25499 2601 25509
rect 2635 25499 2677 25509
rect 2711 25499 2753 25509
rect 2787 25499 2829 25509
rect 2863 25499 2904 25509
rect 2938 25499 2979 25509
rect 3013 25499 3054 25509
rect 3088 25499 3129 25509
rect 3163 25499 3248 25533
rect 664 25458 703 25492
rect 664 25419 728 25458
rect 664 25385 703 25419
rect 664 25346 728 25385
rect 664 25312 703 25346
rect 664 25273 728 25312
rect 664 25239 703 25273
rect 664 25200 728 25239
rect 664 25166 703 25200
rect 664 25127 728 25166
rect 664 25093 703 25127
rect 664 25054 728 25093
rect 664 25020 703 25054
rect 664 25003 728 25020
rect 966 25003 1048 25499
rect 2242 25475 3248 25499
rect 2242 25461 2306 25475
rect 2340 25461 2378 25475
rect 2412 25461 2450 25475
rect 2242 25427 2297 25461
rect 2340 25441 2373 25461
rect 2412 25441 2449 25461
rect 2484 25441 2522 25475
rect 2556 25461 2594 25475
rect 2628 25461 2666 25475
rect 2700 25461 2737 25475
rect 2771 25461 2808 25475
rect 2842 25461 2879 25475
rect 2913 25461 2950 25475
rect 2984 25461 3021 25475
rect 3055 25461 3092 25475
rect 2559 25441 2594 25461
rect 2635 25441 2666 25461
rect 2711 25441 2737 25461
rect 2787 25441 2808 25461
rect 2863 25441 2879 25461
rect 2938 25441 2950 25461
rect 3013 25441 3021 25461
rect 3088 25441 3092 25461
rect 3126 25461 3248 25475
rect 3126 25441 3129 25461
rect 2331 25427 2373 25441
rect 2407 25427 2449 25441
rect 2483 25427 2525 25441
rect 2559 25427 2601 25441
rect 2635 25427 2677 25441
rect 2711 25427 2753 25441
rect 2787 25427 2829 25441
rect 2863 25427 2904 25441
rect 2938 25427 2979 25441
rect 3013 25427 3054 25441
rect 3088 25427 3129 25441
rect 3163 25427 3248 25461
rect 2242 25407 3248 25427
rect 2242 25389 2306 25407
rect 2340 25389 2378 25407
rect 2412 25389 2450 25407
rect 2242 25355 2297 25389
rect 2340 25373 2373 25389
rect 2412 25373 2449 25389
rect 2484 25373 2522 25407
rect 2556 25389 2594 25407
rect 2628 25389 2666 25407
rect 2700 25389 2737 25407
rect 2771 25389 2808 25407
rect 2842 25389 2879 25407
rect 2913 25389 2950 25407
rect 2984 25389 3021 25407
rect 3055 25389 3092 25407
rect 2559 25373 2594 25389
rect 2635 25373 2666 25389
rect 2711 25373 2737 25389
rect 2787 25373 2808 25389
rect 2863 25373 2879 25389
rect 2938 25373 2950 25389
rect 3013 25373 3021 25389
rect 3088 25373 3092 25389
rect 3126 25389 3248 25407
rect 3126 25373 3129 25389
rect 2331 25355 2373 25373
rect 2407 25355 2449 25373
rect 2483 25355 2525 25373
rect 2559 25355 2601 25373
rect 2635 25355 2677 25373
rect 2711 25355 2753 25373
rect 2787 25355 2829 25373
rect 2863 25355 2904 25373
rect 2938 25355 2979 25373
rect 3013 25355 3054 25373
rect 3088 25355 3129 25373
rect 3163 25355 3248 25389
rect 664 24981 1048 25003
rect 664 24947 703 24981
rect 737 24968 775 24981
rect 809 24968 847 24981
rect 881 24968 919 24981
rect 953 24968 1048 24981
rect 762 24947 775 24968
rect 830 24947 847 24968
rect 898 24947 919 24968
rect 664 24934 728 24947
rect 762 24934 796 24947
rect 830 24934 864 24947
rect 898 24934 932 24947
rect 966 24934 1048 24968
rect 664 24908 1048 24934
rect 664 24874 703 24908
rect 737 24899 775 24908
rect 809 24899 847 24908
rect 881 24899 919 24908
rect 953 24899 1048 24908
rect 762 24874 775 24899
rect 830 24874 847 24899
rect 898 24874 919 24899
rect 664 24865 728 24874
rect 762 24865 796 24874
rect 830 24865 864 24874
rect 898 24865 932 24874
rect 966 24865 1048 24899
rect 664 24835 1048 24865
rect 664 24801 703 24835
rect 737 24830 775 24835
rect 809 24830 847 24835
rect 881 24830 919 24835
rect 953 24830 1048 24835
rect 762 24801 775 24830
rect 830 24801 847 24830
rect 898 24801 919 24830
rect 664 24796 728 24801
rect 762 24796 796 24801
rect 830 24796 864 24801
rect 898 24796 932 24801
rect 966 24796 1048 24830
rect 664 24762 1048 24796
rect 664 24728 703 24762
rect 737 24761 775 24762
rect 809 24761 847 24762
rect 881 24761 919 24762
rect 953 24761 1048 24762
rect 762 24728 775 24761
rect 830 24728 847 24761
rect 898 24728 919 24761
rect 664 24727 728 24728
rect 762 24727 796 24728
rect 830 24727 864 24728
rect 898 24727 932 24728
rect 966 24727 1048 24761
rect 664 24692 1048 24727
rect 664 24689 728 24692
rect 762 24689 796 24692
rect 830 24689 864 24692
rect 898 24689 932 24692
rect 664 24655 703 24689
rect 762 24658 775 24689
rect 830 24658 847 24689
rect 898 24658 919 24689
rect 966 24658 1048 24692
rect 737 24655 775 24658
rect 809 24655 847 24658
rect 881 24655 919 24658
rect 953 24655 1048 24658
rect 664 24623 1048 24655
rect 664 24616 728 24623
rect 762 24616 796 24623
rect 830 24616 864 24623
rect 898 24616 932 24623
rect 664 24582 703 24616
rect 762 24589 775 24616
rect 830 24589 847 24616
rect 898 24589 919 24616
rect 966 24589 1048 24623
rect 737 24582 775 24589
rect 809 24582 847 24589
rect 881 24582 919 24589
rect 953 24582 1048 24589
rect 664 24554 1048 24582
rect 664 24543 728 24554
rect 762 24543 796 24554
rect 830 24543 864 24554
rect 898 24543 932 24554
rect 664 24509 703 24543
rect 762 24520 775 24543
rect 830 24520 847 24543
rect 898 24520 919 24543
rect 966 24520 1048 24554
rect 737 24509 775 24520
rect 809 24509 847 24520
rect 881 24509 919 24520
rect 953 24509 1048 24520
rect 664 24485 1048 24509
rect 664 24470 728 24485
rect 762 24470 796 24485
rect 830 24470 864 24485
rect 898 24470 932 24485
rect 664 24436 703 24470
rect 762 24451 775 24470
rect 830 24451 847 24470
rect 898 24451 919 24470
rect 966 24451 1048 24485
rect 737 24436 775 24451
rect 809 24436 847 24451
rect 881 24436 919 24451
rect 953 24436 1048 24451
rect 664 24416 1048 24436
rect 664 24397 728 24416
rect 762 24397 796 24416
rect 830 24397 864 24416
rect 898 24397 932 24416
rect 664 24363 703 24397
rect 762 24382 775 24397
rect 830 24382 847 24397
rect 898 24382 919 24397
rect 966 24382 1048 24416
rect 737 24363 775 24382
rect 809 24363 847 24382
rect 881 24363 919 24382
rect 953 24363 1048 24382
rect 664 24347 1048 24363
rect 664 24324 728 24347
rect 762 24324 796 24347
rect 830 24324 864 24347
rect 898 24324 932 24347
rect 664 24290 703 24324
rect 762 24313 775 24324
rect 830 24313 847 24324
rect 898 24313 919 24324
rect 966 24313 1048 24347
rect 737 24290 775 24313
rect 809 24290 847 24313
rect 881 24290 919 24313
rect 953 24290 1048 24313
rect 664 24278 1048 24290
rect 664 24251 728 24278
rect 762 24251 796 24278
rect 830 24251 864 24278
rect 898 24251 932 24278
rect 664 24217 703 24251
rect 762 24244 775 24251
rect 830 24244 847 24251
rect 898 24244 919 24251
rect 966 24244 1048 24278
rect 737 24217 775 24244
rect 809 24217 847 24244
rect 881 24217 919 24244
rect 953 24217 1048 24244
rect 664 24209 1048 24217
rect 664 24178 728 24209
rect 762 24178 796 24209
rect 830 24178 864 24209
rect 898 24178 932 24209
rect 664 24144 703 24178
rect 762 24175 775 24178
rect 830 24175 847 24178
rect 898 24175 919 24178
rect 966 24175 1048 24209
rect 737 24144 775 24175
rect 809 24144 847 24175
rect 881 24144 919 24175
rect 953 24144 1048 24175
rect 664 24140 1048 24144
rect 664 24106 728 24140
rect 762 24106 796 24140
rect 830 24106 864 24140
rect 898 24106 932 24140
rect 966 24106 1048 24140
rect 664 24105 1048 24106
rect 664 24071 703 24105
rect 737 24071 775 24105
rect 809 24071 847 24105
rect 881 24071 919 24105
rect 953 24071 1048 24105
rect 664 24037 728 24071
rect 762 24037 796 24071
rect 830 24037 864 24071
rect 898 24037 932 24071
rect 966 24037 1048 24071
rect 664 24031 1048 24037
rect 664 23997 703 24031
rect 737 24002 775 24031
rect 809 24002 847 24031
rect 881 24002 919 24031
rect 953 24002 1048 24031
rect 762 23997 775 24002
rect 830 23997 847 24002
rect 898 23997 919 24002
rect 664 23968 728 23997
rect 762 23968 796 23997
rect 830 23968 864 23997
rect 898 23968 932 23997
rect 966 23968 1048 24002
rect 664 23957 1048 23968
rect 664 23923 703 23957
rect 737 23933 775 23957
rect 809 23933 847 23957
rect 881 23933 919 23957
rect 953 23933 1048 23957
rect 762 23923 775 23933
rect 830 23923 847 23933
rect 898 23923 919 23933
rect 664 23899 728 23923
rect 762 23899 796 23923
rect 830 23899 864 23923
rect 898 23899 932 23923
rect 966 23899 1048 23933
rect 664 23883 1048 23899
rect 664 23849 703 23883
rect 737 23864 775 23883
rect 809 23864 847 23883
rect 881 23864 919 23883
rect 953 23864 1048 23883
rect 762 23849 775 23864
rect 830 23849 847 23864
rect 898 23849 919 23864
rect 664 23830 728 23849
rect 762 23830 796 23849
rect 830 23830 864 23849
rect 898 23830 932 23849
rect 966 23830 1048 23864
rect 664 23809 1048 23830
rect 664 23775 703 23809
rect 737 23795 775 23809
rect 809 23795 847 23809
rect 881 23795 919 23809
rect 953 23795 1048 23809
rect 762 23775 775 23795
rect 830 23775 847 23795
rect 898 23775 919 23795
rect 664 23761 728 23775
rect 762 23761 796 23775
rect 830 23761 864 23775
rect 898 23761 932 23775
rect 966 23761 1048 23795
rect 664 23735 1048 23761
rect 664 23701 703 23735
rect 737 23726 775 23735
rect 809 23726 847 23735
rect 881 23726 919 23735
rect 953 23726 1048 23735
rect 762 23701 775 23726
rect 830 23701 847 23726
rect 898 23701 919 23726
rect 664 23692 728 23701
rect 762 23692 796 23701
rect 830 23692 864 23701
rect 898 23692 932 23701
rect 966 23692 1048 23726
rect 664 23661 1048 23692
rect 664 23627 703 23661
rect 737 23657 775 23661
rect 809 23657 847 23661
rect 881 23657 919 23661
rect 953 23657 1048 23661
rect 762 23627 775 23657
rect 830 23627 847 23657
rect 898 23627 919 23657
rect 664 23623 728 23627
rect 762 23623 796 23627
rect 830 23623 864 23627
rect 898 23623 932 23627
rect 966 23623 1048 23657
rect 664 23588 1048 23623
rect 664 23587 728 23588
rect 762 23587 796 23588
rect 830 23587 864 23588
rect 898 23587 932 23588
rect 664 23553 703 23587
rect 762 23554 775 23587
rect 830 23554 847 23587
rect 898 23554 919 23587
rect 966 23554 1048 23588
rect 737 23553 775 23554
rect 809 23553 847 23554
rect 881 23553 919 23554
rect 953 23553 1048 23554
rect 664 23519 1048 23553
rect 664 23513 728 23519
rect 762 23513 796 23519
rect 830 23513 864 23519
rect 898 23513 932 23519
rect 664 23479 703 23513
rect 762 23485 775 23513
rect 830 23485 847 23513
rect 898 23485 919 23513
rect 966 23485 1048 23519
rect 737 23479 775 23485
rect 809 23479 847 23485
rect 881 23479 919 23485
rect 953 23479 1048 23485
rect 664 23450 1048 23479
rect 664 23439 728 23450
rect 762 23439 796 23450
rect 830 23439 864 23450
rect 898 23439 932 23450
rect 664 23405 703 23439
rect 762 23416 775 23439
rect 830 23416 847 23439
rect 898 23416 919 23439
rect 966 23416 1048 23450
rect 737 23405 775 23416
rect 809 23405 847 23416
rect 881 23405 919 23416
rect 953 23405 1048 23416
rect 664 23381 1048 23405
rect 664 23365 728 23381
rect 762 23365 796 23381
rect 830 23365 864 23381
rect 898 23365 932 23381
rect 664 23331 703 23365
rect 762 23347 775 23365
rect 830 23347 847 23365
rect 898 23347 919 23365
rect 966 23347 1048 23381
rect 737 23331 775 23347
rect 809 23331 847 23347
rect 881 23331 919 23347
rect 953 23331 1048 23347
rect 664 23312 1048 23331
rect 664 23291 728 23312
rect 762 23291 796 23312
rect 830 23291 864 23312
rect 898 23291 932 23312
rect 664 23257 703 23291
rect 762 23278 775 23291
rect 830 23278 847 23291
rect 898 23278 919 23291
rect 966 23278 1048 23312
rect 737 23257 775 23278
rect 809 23257 847 23278
rect 881 23257 919 23278
rect 953 23257 1048 23278
rect 664 23225 1048 23257
rect 1308 25313 1352 25347
rect 1386 25313 1430 25347
rect 1464 25313 1508 25347
rect 1542 25313 1587 25347
rect 1621 25313 1666 25347
rect 1700 25313 1745 25347
rect 1779 25313 1824 25347
rect 1858 25313 1903 25347
rect 1937 25313 1982 25347
rect 1200 25267 1234 25307
rect 1200 25193 1234 25233
rect 1200 25119 1234 25159
rect 1200 25045 1234 25085
rect 1200 24971 1234 25011
rect 1200 24897 1234 24937
rect 1200 24824 1234 24863
rect 1200 24751 1234 24790
rect 1200 24678 1234 24717
rect 1200 24605 1234 24644
rect 1200 24532 1234 24571
rect 1200 24459 1234 24498
rect 1200 24386 1234 24425
rect 1200 24313 1234 24352
rect 1200 24240 1234 24279
rect 1200 24167 1234 24206
rect 1200 24094 1234 24133
rect 1200 24021 1234 24060
rect 1200 23948 1234 23987
rect 1200 23875 1234 23914
rect 1200 23802 1234 23841
rect 1200 23729 1234 23768
rect 1200 23656 1234 23695
rect 1200 23583 1234 23622
rect 1200 23510 1234 23549
rect 1200 23437 1234 23476
rect 1200 23364 1234 23403
rect 1200 23291 1234 23330
rect 1200 23218 1234 23257
rect 1200 23145 1234 23184
rect 2056 25268 2090 25307
rect 2056 25195 2090 25234
rect 2056 25122 2090 25161
rect 2056 25049 2090 25088
rect 2056 24976 2090 25015
rect 2056 24903 2090 24942
rect 2056 24830 2090 24869
rect 2056 24757 2090 24796
rect 2056 24684 2090 24723
rect 2242 25339 3248 25355
rect 2242 25317 2306 25339
rect 2340 25317 2378 25339
rect 2412 25317 2450 25339
rect 2242 25283 2297 25317
rect 2340 25305 2373 25317
rect 2412 25305 2449 25317
rect 2484 25305 2522 25339
rect 2556 25317 2594 25339
rect 2628 25317 2666 25339
rect 2700 25317 2737 25339
rect 2771 25317 2808 25339
rect 2842 25317 2879 25339
rect 2913 25317 2950 25339
rect 2984 25317 3021 25339
rect 3055 25317 3092 25339
rect 2559 25305 2594 25317
rect 2635 25305 2666 25317
rect 2711 25305 2737 25317
rect 2787 25305 2808 25317
rect 2863 25305 2879 25317
rect 2938 25305 2950 25317
rect 3013 25305 3021 25317
rect 3088 25305 3092 25317
rect 3126 25317 3248 25339
rect 3126 25305 3129 25317
rect 2331 25283 2373 25305
rect 2407 25283 2449 25305
rect 2483 25283 2525 25305
rect 2559 25283 2601 25305
rect 2635 25283 2677 25305
rect 2711 25283 2753 25305
rect 2787 25283 2829 25305
rect 2863 25283 2904 25305
rect 2938 25283 2979 25305
rect 3013 25283 3054 25305
rect 3088 25283 3129 25305
rect 3163 25283 3248 25317
rect 2242 25271 3248 25283
rect 2242 25245 2306 25271
rect 2340 25245 2378 25271
rect 2412 25245 2450 25271
rect 2242 25211 2297 25245
rect 2340 25237 2373 25245
rect 2412 25237 2449 25245
rect 2484 25237 2522 25271
rect 2556 25245 2594 25271
rect 2628 25245 2666 25271
rect 2700 25245 2737 25271
rect 2771 25245 2808 25271
rect 2842 25245 2879 25271
rect 2913 25245 2950 25271
rect 2984 25245 3021 25271
rect 3055 25245 3092 25271
rect 2559 25237 2594 25245
rect 2635 25237 2666 25245
rect 2711 25237 2737 25245
rect 2787 25237 2808 25245
rect 2863 25237 2879 25245
rect 2938 25237 2950 25245
rect 3013 25237 3021 25245
rect 3088 25237 3092 25245
rect 3126 25245 3248 25271
rect 3126 25237 3129 25245
rect 2331 25211 2373 25237
rect 2407 25211 2449 25237
rect 2483 25211 2525 25237
rect 2559 25211 2601 25237
rect 2635 25211 2677 25237
rect 2711 25211 2753 25237
rect 2787 25211 2829 25237
rect 2863 25211 2904 25237
rect 2938 25211 2979 25237
rect 3013 25211 3054 25237
rect 3088 25211 3129 25237
rect 3163 25211 3248 25245
rect 2242 25203 3248 25211
rect 2242 25173 2306 25203
rect 2340 25173 2378 25203
rect 2412 25173 2450 25203
rect 2242 25139 2297 25173
rect 2340 25169 2373 25173
rect 2412 25169 2449 25173
rect 2484 25169 2522 25203
rect 2556 25173 2594 25203
rect 2628 25173 2666 25203
rect 2700 25173 2737 25203
rect 2771 25173 2808 25203
rect 2842 25173 2879 25203
rect 2913 25173 2950 25203
rect 2984 25173 3021 25203
rect 3055 25173 3092 25203
rect 2559 25169 2594 25173
rect 2635 25169 2666 25173
rect 2711 25169 2737 25173
rect 2787 25169 2808 25173
rect 2863 25169 2879 25173
rect 2938 25169 2950 25173
rect 3013 25169 3021 25173
rect 3088 25169 3092 25173
rect 3126 25173 3248 25203
rect 3126 25169 3129 25173
rect 2331 25139 2373 25169
rect 2407 25139 2449 25169
rect 2483 25139 2525 25169
rect 2559 25139 2601 25169
rect 2635 25139 2677 25169
rect 2711 25139 2753 25169
rect 2787 25139 2829 25169
rect 2863 25139 2904 25169
rect 2938 25139 2979 25169
rect 3013 25139 3054 25169
rect 3088 25139 3129 25169
rect 3163 25139 3248 25173
rect 2242 25135 3248 25139
rect 2242 25101 2306 25135
rect 2340 25101 2378 25135
rect 2412 25101 2450 25135
rect 2484 25101 2522 25135
rect 2556 25101 2594 25135
rect 2628 25101 2666 25135
rect 2700 25101 2737 25135
rect 2771 25101 2808 25135
rect 2842 25101 2879 25135
rect 2913 25101 2950 25135
rect 2984 25101 3021 25135
rect 3055 25101 3092 25135
rect 3126 25101 3248 25135
rect 2242 25067 2297 25101
rect 2331 25067 2373 25101
rect 2407 25067 2449 25101
rect 2483 25067 2525 25101
rect 2559 25067 2601 25101
rect 2635 25067 2677 25101
rect 2711 25067 2753 25101
rect 2787 25067 2829 25101
rect 2863 25067 2904 25101
rect 2938 25067 2979 25101
rect 3013 25067 3054 25101
rect 3088 25067 3129 25101
rect 3163 25067 3248 25101
rect 2242 25033 2306 25067
rect 2340 25033 2378 25067
rect 2412 25033 2450 25067
rect 2484 25033 2522 25067
rect 2556 25033 2594 25067
rect 2628 25033 2666 25067
rect 2700 25033 2737 25067
rect 2771 25033 2808 25067
rect 2842 25033 2879 25067
rect 2913 25033 2950 25067
rect 2984 25033 3021 25067
rect 3055 25033 3092 25067
rect 3126 25033 3248 25067
rect 2242 25029 3248 25033
rect 2242 24995 2297 25029
rect 2331 24999 2373 25029
rect 2407 24999 2449 25029
rect 2483 24999 2525 25029
rect 2559 24999 2601 25029
rect 2635 24999 2677 25029
rect 2711 24999 2753 25029
rect 2787 24999 2829 25029
rect 2863 24999 2904 25029
rect 2938 24999 2979 25029
rect 3013 24999 3054 25029
rect 3088 24999 3129 25029
rect 2340 24995 2373 24999
rect 2412 24995 2449 24999
rect 2242 24965 2306 24995
rect 2340 24965 2378 24995
rect 2412 24965 2450 24995
rect 2484 24965 2522 24999
rect 2559 24995 2594 24999
rect 2635 24995 2666 24999
rect 2711 24995 2737 24999
rect 2787 24995 2808 24999
rect 2863 24995 2879 24999
rect 2938 24995 2950 24999
rect 3013 24995 3021 24999
rect 3088 24995 3092 24999
rect 2556 24965 2594 24995
rect 2628 24965 2666 24995
rect 2700 24965 2737 24995
rect 2771 24965 2808 24995
rect 2842 24965 2879 24995
rect 2913 24965 2950 24995
rect 2984 24965 3021 24995
rect 3055 24965 3092 24995
rect 3126 24995 3129 24999
rect 3163 24995 3248 25029
rect 3126 24965 3248 24995
rect 2242 24957 3248 24965
rect 2242 24923 2297 24957
rect 2331 24931 2373 24957
rect 2407 24931 2449 24957
rect 2483 24931 2525 24957
rect 2559 24931 2601 24957
rect 2635 24931 2677 24957
rect 2711 24931 2753 24957
rect 2787 24931 2829 24957
rect 2863 24931 2904 24957
rect 2938 24931 2979 24957
rect 3013 24931 3054 24957
rect 3088 24931 3129 24957
rect 2340 24923 2373 24931
rect 2412 24923 2449 24931
rect 2242 24897 2306 24923
rect 2340 24897 2378 24923
rect 2412 24897 2450 24923
rect 2484 24897 2522 24931
rect 2559 24923 2594 24931
rect 2635 24923 2666 24931
rect 2711 24923 2737 24931
rect 2787 24923 2808 24931
rect 2863 24923 2879 24931
rect 2938 24923 2950 24931
rect 3013 24923 3021 24931
rect 3088 24923 3092 24931
rect 2556 24897 2594 24923
rect 2628 24897 2666 24923
rect 2700 24897 2737 24923
rect 2771 24897 2808 24923
rect 2842 24897 2879 24923
rect 2913 24897 2950 24923
rect 2984 24897 3021 24923
rect 3055 24897 3092 24923
rect 3126 24923 3129 24931
rect 3163 24923 3248 24957
rect 3126 24897 3248 24923
rect 2242 24885 3248 24897
rect 2242 24851 2297 24885
rect 2331 24863 2373 24885
rect 2407 24863 2449 24885
rect 2483 24863 2525 24885
rect 2559 24863 2601 24885
rect 2635 24863 2677 24885
rect 2711 24863 2753 24885
rect 2787 24863 2829 24885
rect 2863 24863 2904 24885
rect 2938 24863 2979 24885
rect 3013 24863 3054 24885
rect 3088 24863 3129 24885
rect 2340 24851 2373 24863
rect 2412 24851 2449 24863
rect 2242 24829 2306 24851
rect 2340 24829 2378 24851
rect 2412 24829 2450 24851
rect 2484 24829 2522 24863
rect 2559 24851 2594 24863
rect 2635 24851 2666 24863
rect 2711 24851 2737 24863
rect 2787 24851 2808 24863
rect 2863 24851 2879 24863
rect 2938 24851 2950 24863
rect 3013 24851 3021 24863
rect 3088 24851 3092 24863
rect 2556 24829 2594 24851
rect 2628 24829 2666 24851
rect 2700 24829 2737 24851
rect 2771 24829 2808 24851
rect 2842 24829 2879 24851
rect 2913 24829 2950 24851
rect 2984 24829 3021 24851
rect 3055 24829 3092 24851
rect 3126 24851 3129 24863
rect 3163 24851 3248 24885
rect 3126 24829 3248 24851
rect 2242 24813 3248 24829
rect 2242 24779 2297 24813
rect 2331 24795 2373 24813
rect 2407 24795 2449 24813
rect 2483 24795 2525 24813
rect 2559 24795 2601 24813
rect 2635 24795 2677 24813
rect 2711 24795 2753 24813
rect 2787 24795 2829 24813
rect 2863 24795 2904 24813
rect 2938 24795 2979 24813
rect 3013 24795 3054 24813
rect 3088 24795 3129 24813
rect 2340 24779 2373 24795
rect 2412 24779 2449 24795
rect 2242 24761 2306 24779
rect 2340 24761 2378 24779
rect 2412 24761 2450 24779
rect 2484 24761 2522 24795
rect 2559 24779 2594 24795
rect 2635 24779 2666 24795
rect 2711 24779 2737 24795
rect 2787 24779 2808 24795
rect 2863 24779 2879 24795
rect 2938 24779 2950 24795
rect 3013 24779 3021 24795
rect 3088 24779 3092 24795
rect 2556 24761 2594 24779
rect 2628 24761 2666 24779
rect 2700 24761 2737 24779
rect 2771 24761 2808 24779
rect 2842 24761 2879 24779
rect 2913 24761 2950 24779
rect 2984 24761 3021 24779
rect 3055 24761 3092 24779
rect 3126 24779 3129 24795
rect 3163 24779 3248 24813
rect 3126 24761 3248 24779
rect 2242 24708 3248 24761
rect 2056 24612 2090 24650
rect 2056 24540 2090 24578
rect 2164 24522 2207 24556
rect 2241 24522 2284 24556
rect 2318 24522 2361 24556
rect 2395 24522 2438 24556
rect 2472 24522 2515 24556
rect 2549 24522 2592 24556
rect 2626 24522 2669 24556
rect 2703 24522 2746 24556
rect 2780 24522 2823 24556
rect 2857 24522 2900 24556
rect 2056 24468 2090 24506
rect 2056 24396 2090 24434
rect 2056 24324 2090 24362
rect 2056 24252 2090 24290
rect 2056 24180 2090 24218
rect 2056 24108 2090 24146
rect 2056 24036 2090 24074
rect 2056 23964 2090 24002
rect 2056 23892 2090 23930
rect 2056 23820 2090 23858
rect 2056 23748 2090 23786
rect 2056 23676 2090 23714
rect 2056 23604 2090 23642
rect 2056 23532 2090 23570
rect 2056 23460 2090 23498
rect 2056 23388 2090 23426
rect 2056 23316 2090 23354
rect 2056 23244 2090 23282
rect 2056 23172 2090 23210
rect 2056 23100 2090 23138
rect 816 23039 822 23047
rect 856 23039 894 23073
rect 928 23039 966 23073
rect 1000 23039 1038 23073
rect 1072 23039 1110 23073
rect 1144 23039 1182 23073
rect 1216 23039 1254 23073
rect 1288 23039 1326 23073
rect 1360 23039 1398 23073
rect 1432 23039 1471 23073
rect 1505 23039 1544 23073
rect 1578 23039 1617 23073
rect 1651 23039 1690 23073
rect 1724 23039 1763 23073
rect 1797 23039 1836 23073
rect 1870 23039 1909 23073
rect 1943 23039 1982 23073
rect 816 23001 850 23039
rect 2056 23029 2090 23066
rect 2056 22958 2090 22994
rect 1034 22914 1077 22948
rect 1111 22914 1154 22948
rect 1188 22914 1231 22948
rect 1265 22914 1308 22948
rect 1342 22914 1384 22948
rect 1418 22914 1460 22948
rect 1494 22914 1536 22948
rect 1570 22914 1612 22948
rect 1646 22914 1688 22948
rect 1722 22914 1764 22948
rect 1798 22914 1840 22948
rect 1874 22914 1916 22948
rect 888 22886 949 22903
rect 922 22852 949 22886
rect 888 22791 949 22852
rect 2056 22887 2090 22924
rect 2056 22816 2090 22853
rect 922 22757 949 22791
rect 1033 22758 1076 22792
rect 1110 22758 1153 22792
rect 1187 22758 1230 22792
rect 1264 22758 1307 22792
rect 1341 22758 1384 22792
rect 1418 22758 1460 22792
rect 1494 22758 1536 22792
rect 1570 22758 1612 22792
rect 1646 22758 1688 22792
rect 1722 22758 1764 22792
rect 1798 22758 1840 22792
rect 1874 22758 1916 22792
rect 2056 22762 2090 22782
rect 888 22698 949 22757
rect 888 22697 909 22698
rect 943 22664 949 22698
rect 922 22663 949 22664
rect 888 22647 949 22663
rect 2056 22687 2090 22710
rect 909 22626 943 22647
rect 1034 22602 1077 22636
rect 1111 22602 1154 22636
rect 1188 22602 1231 22636
rect 1265 22602 1308 22636
rect 1342 22602 1384 22636
rect 1418 22602 1460 22636
rect 1494 22602 1536 22636
rect 1570 22602 1612 22636
rect 1646 22602 1688 22636
rect 1722 22602 1764 22636
rect 1798 22602 1840 22636
rect 1874 22602 1916 22636
rect 2056 22612 2090 22638
rect 2056 22536 2090 22566
rect 816 22476 850 22518
rect 816 22400 850 22442
rect 888 22499 949 22515
rect 922 22498 949 22499
rect 888 22464 912 22465
rect 946 22464 949 22498
rect 1033 22492 1076 22526
rect 1110 22492 1153 22526
rect 1187 22492 1230 22526
rect 1264 22492 1307 22526
rect 1341 22492 1384 22526
rect 1418 22492 1460 22526
rect 1494 22492 1536 22526
rect 1570 22492 1612 22526
rect 1646 22492 1688 22526
rect 1722 22492 1764 22526
rect 1798 22492 1840 22526
rect 1874 22492 1916 22526
rect 888 22431 949 22464
rect 922 22426 949 22431
rect 888 22392 912 22397
rect 946 22392 949 22426
rect 888 22381 949 22392
rect 2056 22460 2090 22494
rect 2056 22384 2090 22422
rect 816 22324 850 22366
rect 1033 22336 1076 22370
rect 1110 22336 1153 22370
rect 1187 22336 1230 22370
rect 1264 22336 1307 22370
rect 1341 22336 1384 22370
rect 1418 22336 1460 22370
rect 1494 22336 1536 22370
rect 1570 22336 1612 22370
rect 1646 22336 1688 22370
rect 1722 22336 1764 22370
rect 1798 22336 1840 22370
rect 1874 22336 1916 22370
rect 816 22248 850 22290
rect 816 22172 850 22214
rect 816 22096 850 22138
rect 816 22020 850 22062
rect 816 21943 850 21986
rect 816 21866 850 21909
rect 816 21789 850 21832
rect 816 21712 850 21755
rect 816 21635 850 21678
rect 816 21558 850 21601
rect 816 21481 850 21524
rect 816 21404 850 21447
rect 2056 22312 2090 22350
rect 2056 22232 2090 22274
rect 2056 22156 2090 22198
rect 2056 22080 2090 22122
rect 2056 22004 2090 22046
rect 2056 21928 2090 21970
rect 2056 21852 2090 21894
rect 2912 24388 2946 24427
rect 2912 24315 2946 24354
rect 2912 24242 2946 24281
rect 2912 24169 2946 24208
rect 2912 24096 2946 24135
rect 2912 24023 2946 24062
rect 2912 23950 2946 23989
rect 2912 23877 2946 23916
rect 2912 23804 2946 23843
rect 2912 23731 2946 23770
rect 2912 23658 2946 23697
rect 2912 23585 2946 23624
rect 3098 23606 3248 24708
rect 2912 23512 2946 23551
rect 2912 23439 2946 23478
rect 2912 23365 2946 23405
rect 2912 23291 2946 23331
rect 2912 23217 2946 23257
rect 2912 23143 2946 23183
rect 2912 23069 2946 23109
rect 2912 22995 2946 23035
rect 2912 22921 2946 22961
rect 2912 22847 2946 22887
rect 2912 22773 2946 22813
rect 2912 22699 2946 22739
rect 2912 22625 2946 22665
rect 2912 22551 2946 22591
rect 2912 22477 2946 22517
rect 2912 22403 2946 22443
rect 2912 22329 2946 22369
rect 2912 22255 2946 22295
rect 2912 22181 2946 22221
rect 2912 22107 2946 22147
rect 2912 22033 2946 22073
rect 2912 21959 2946 21999
rect 2912 21885 2946 21925
rect 2056 21776 2090 21818
rect 2056 21700 2090 21742
rect 2056 21624 2090 21666
rect 2912 21645 2946 21685
rect 2056 21548 2090 21590
rect 2056 21472 2090 21514
rect 924 21364 962 21398
rect 996 21364 1034 21398
rect 1068 21364 1106 21398
rect 1140 21364 1178 21398
rect 1212 21364 1250 21398
rect 1284 21364 1322 21398
rect 1356 21364 1394 21398
rect 1428 21364 1466 21398
rect 1500 21364 1538 21398
rect 1572 21364 1610 21398
rect 1644 21364 1682 21398
rect 1716 21364 1754 21398
rect 1788 21364 1826 21398
rect 1860 21364 1898 21398
rect 1932 21364 1970 21398
rect 2004 21364 2042 21398
rect 2076 21364 2115 21398
rect 2149 21364 2188 21398
rect 2222 21364 2261 21398
rect 265 18694 281 18728
rect 315 18694 349 18728
rect 383 18694 417 18728
rect 451 18694 485 18728
rect 519 18694 553 18728
rect 587 18694 603 18728
rect 265 18144 603 18694
rect 515 18038 603 18144
rect 2676 16961 17039 16980
rect 2676 16927 2710 16961
rect 2744 16927 2779 16961
rect 2813 16927 2848 16961
rect 2882 16927 2917 16961
rect 2951 16927 2986 16961
rect 3020 16927 3055 16961
rect 3089 16927 3124 16961
rect 3158 16927 3193 16961
rect 3227 16927 3262 16961
rect 3296 16927 3331 16961
rect 3365 16927 3400 16961
rect 3434 16927 3469 16961
rect 3503 16927 3538 16961
rect 3572 16927 3607 16961
rect 3641 16927 3676 16961
rect 3710 16927 3745 16961
rect 3779 16927 3814 16961
rect 3848 16927 3883 16961
rect 3917 16927 3952 16961
rect 3986 16927 4021 16961
rect 4055 16927 4090 16961
rect 4124 16927 4159 16961
rect 4193 16927 4228 16961
rect 4262 16927 4297 16961
rect 4331 16927 4366 16961
rect 4400 16927 4435 16961
rect 4469 16927 4504 16961
rect 4538 16927 4573 16961
rect 4607 16927 4642 16961
rect 4676 16927 4711 16961
rect 4745 16927 4780 16961
rect 4814 16927 4849 16961
rect 4883 16927 4918 16961
rect 4952 16927 4987 16961
rect 5021 16927 5056 16961
rect 5090 16927 5125 16961
rect 5159 16927 5194 16961
rect 5228 16927 5263 16961
rect 5297 16927 5332 16961
rect 5366 16927 5401 16961
rect 5435 16927 5470 16961
rect 5504 16927 5539 16961
rect 5573 16927 5608 16961
rect 5642 16927 5677 16961
rect 5711 16927 5746 16961
rect 5780 16927 5815 16961
rect 5849 16927 5884 16961
rect 5918 16927 5953 16961
rect 5987 16927 6022 16961
rect 6056 16927 6091 16961
rect 2676 16893 6091 16927
rect 2676 16859 2710 16893
rect 2744 16859 2779 16893
rect 2813 16859 2848 16893
rect 2882 16859 2917 16893
rect 2951 16859 2986 16893
rect 3020 16859 3055 16893
rect 3089 16859 3124 16893
rect 3158 16859 3193 16893
rect 3227 16859 3262 16893
rect 3296 16859 3331 16893
rect 3365 16859 3400 16893
rect 3434 16859 3469 16893
rect 3503 16859 3538 16893
rect 3572 16859 3607 16893
rect 3641 16859 3676 16893
rect 3710 16859 3745 16893
rect 3779 16859 3814 16893
rect 3848 16859 3883 16893
rect 3917 16859 3952 16893
rect 3986 16859 4021 16893
rect 4055 16859 4090 16893
rect 4124 16859 4159 16893
rect 4193 16859 4228 16893
rect 4262 16859 4297 16893
rect 4331 16859 4366 16893
rect 4400 16859 4435 16893
rect 4469 16859 4504 16893
rect 4538 16859 4573 16893
rect 4607 16859 4642 16893
rect 4676 16859 4711 16893
rect 4745 16859 4780 16893
rect 4814 16859 4849 16893
rect 4883 16859 4918 16893
rect 4952 16859 4987 16893
rect 5021 16859 5056 16893
rect 5090 16859 5125 16893
rect 5159 16859 5194 16893
rect 5228 16859 5263 16893
rect 5297 16859 5332 16893
rect 5366 16859 5401 16893
rect 5435 16859 5470 16893
rect 5504 16859 5539 16893
rect 5573 16859 5608 16893
rect 5642 16859 5677 16893
rect 5711 16859 5746 16893
rect 5780 16859 5815 16893
rect 5849 16859 5884 16893
rect 5918 16859 5953 16893
rect 5987 16859 6022 16893
rect 6056 16859 6091 16893
rect 2676 16825 6091 16859
rect 2676 16791 2710 16825
rect 2744 16791 2779 16825
rect 2813 16791 2848 16825
rect 2882 16791 2917 16825
rect 2951 16791 2986 16825
rect 3020 16791 3055 16825
rect 3089 16791 3124 16825
rect 3158 16791 3193 16825
rect 3227 16791 3262 16825
rect 3296 16791 3331 16825
rect 3365 16791 3400 16825
rect 3434 16791 3469 16825
rect 3503 16791 3538 16825
rect 3572 16791 3607 16825
rect 3641 16791 3676 16825
rect 3710 16791 3745 16825
rect 3779 16791 3814 16825
rect 3848 16791 3883 16825
rect 3917 16791 3952 16825
rect 3986 16791 4021 16825
rect 4055 16791 4090 16825
rect 4124 16791 4159 16825
rect 4193 16791 4228 16825
rect 4262 16791 4297 16825
rect 4331 16791 4366 16825
rect 4400 16791 4435 16825
rect 4469 16791 4504 16825
rect 4538 16791 4573 16825
rect 4607 16791 4642 16825
rect 4676 16791 4711 16825
rect 4745 16791 4780 16825
rect 4814 16791 4849 16825
rect 4883 16791 4918 16825
rect 4952 16791 4987 16825
rect 5021 16791 5056 16825
rect 5090 16791 5125 16825
rect 5159 16791 5194 16825
rect 5228 16791 5263 16825
rect 5297 16791 5332 16825
rect 5366 16791 5401 16825
rect 5435 16791 5470 16825
rect 5504 16791 5539 16825
rect 5573 16791 5608 16825
rect 5642 16791 5677 16825
rect 5711 16791 5746 16825
rect 5780 16791 5815 16825
rect 5849 16791 5884 16825
rect 5918 16791 5953 16825
rect 5987 16791 6022 16825
rect 6056 16791 6091 16825
rect 2676 16757 6091 16791
rect 2676 16723 2710 16757
rect 2744 16723 2779 16757
rect 2813 16723 2848 16757
rect 2882 16723 2917 16757
rect 2951 16723 2986 16757
rect 3020 16723 3055 16757
rect 3089 16723 3124 16757
rect 3158 16723 3193 16757
rect 3227 16723 3262 16757
rect 3296 16723 3331 16757
rect 3365 16723 3400 16757
rect 3434 16723 3469 16757
rect 3503 16723 3538 16757
rect 3572 16723 3607 16757
rect 3641 16723 3676 16757
rect 3710 16723 3745 16757
rect 3779 16723 3814 16757
rect 3848 16723 3883 16757
rect 3917 16723 3952 16757
rect 3986 16723 4021 16757
rect 4055 16723 4090 16757
rect 4124 16723 4159 16757
rect 4193 16723 4228 16757
rect 4262 16723 4297 16757
rect 4331 16723 4366 16757
rect 4400 16723 4435 16757
rect 4469 16723 4504 16757
rect 4538 16723 4573 16757
rect 4607 16723 4642 16757
rect 4676 16723 4711 16757
rect 4745 16723 4780 16757
rect 4814 16723 4849 16757
rect 4883 16723 4918 16757
rect 4952 16723 4987 16757
rect 5021 16723 5056 16757
rect 5090 16723 5125 16757
rect 5159 16723 5194 16757
rect 5228 16723 5263 16757
rect 5297 16723 5332 16757
rect 5366 16723 5401 16757
rect 5435 16723 5470 16757
rect 5504 16723 5539 16757
rect 5573 16723 5608 16757
rect 5642 16723 5677 16757
rect 5711 16723 5746 16757
rect 5780 16723 5815 16757
rect 5849 16723 5884 16757
rect 5918 16723 5953 16757
rect 5987 16723 6022 16757
rect 6056 16723 6091 16757
rect 2676 16689 6091 16723
rect 2676 16655 2710 16689
rect 2744 16655 2779 16689
rect 2813 16655 2848 16689
rect 2882 16655 2917 16689
rect 2951 16655 2986 16689
rect 3020 16655 3055 16689
rect 3089 16655 3124 16689
rect 3158 16655 3193 16689
rect 3227 16655 3262 16689
rect 3296 16655 3331 16689
rect 3365 16655 3400 16689
rect 3434 16655 3469 16689
rect 3503 16655 3538 16689
rect 3572 16655 3607 16689
rect 3641 16655 3676 16689
rect 3710 16655 3745 16689
rect 3779 16655 3814 16689
rect 3848 16655 3883 16689
rect 3917 16655 3952 16689
rect 3986 16655 4021 16689
rect 4055 16655 4090 16689
rect 4124 16655 4159 16689
rect 4193 16655 4228 16689
rect 4262 16655 4297 16689
rect 4331 16655 4366 16689
rect 4400 16655 4435 16689
rect 4469 16655 4504 16689
rect 4538 16655 4573 16689
rect 4607 16655 4642 16689
rect 4676 16655 4711 16689
rect 4745 16655 4780 16689
rect 4814 16655 4849 16689
rect 4883 16655 4918 16689
rect 4952 16655 4987 16689
rect 5021 16655 5056 16689
rect 5090 16655 5125 16689
rect 5159 16655 5194 16689
rect 5228 16655 5263 16689
rect 5297 16655 5332 16689
rect 5366 16655 5401 16689
rect 5435 16655 5470 16689
rect 5504 16655 5539 16689
rect 5573 16655 5608 16689
rect 5642 16655 5677 16689
rect 5711 16655 5746 16689
rect 5780 16655 5815 16689
rect 5849 16655 5884 16689
rect 5918 16655 5953 16689
rect 5987 16655 6022 16689
rect 6056 16655 6091 16689
rect 300 16588 341 16622
rect 375 16588 417 16622
rect 451 16588 493 16622
rect 527 16588 569 16622
rect 266 16550 603 16588
rect 300 16536 341 16550
rect 375 16536 417 16550
rect 451 16536 493 16550
rect 527 16536 569 16550
rect 265 16516 266 16536
rect 315 16516 341 16536
rect 265 16502 281 16516
rect 315 16502 349 16516
rect 383 16502 417 16536
rect 451 16502 485 16536
rect 527 16516 553 16536
rect 519 16502 553 16516
rect 587 16502 603 16516
rect 2676 16621 6091 16655
rect 2676 16587 2710 16621
rect 2744 16587 2779 16621
rect 2813 16587 2848 16621
rect 2882 16587 2917 16621
rect 2951 16587 2986 16621
rect 3020 16587 3055 16621
rect 3089 16587 3124 16621
rect 3158 16587 3193 16621
rect 3227 16587 3262 16621
rect 3296 16587 3331 16621
rect 3365 16587 3400 16621
rect 3434 16587 3469 16621
rect 3503 16587 3538 16621
rect 3572 16587 3607 16621
rect 3641 16587 3676 16621
rect 3710 16587 3745 16621
rect 3779 16587 3814 16621
rect 3848 16587 3883 16621
rect 3917 16587 3952 16621
rect 3986 16587 4021 16621
rect 4055 16587 4090 16621
rect 4124 16587 4159 16621
rect 4193 16587 4228 16621
rect 4262 16587 4297 16621
rect 4331 16587 4366 16621
rect 4400 16587 4435 16621
rect 4469 16587 4504 16621
rect 4538 16587 4573 16621
rect 4607 16587 4642 16621
rect 4676 16587 4711 16621
rect 4745 16587 4780 16621
rect 4814 16587 4849 16621
rect 4883 16587 4918 16621
rect 4952 16587 4987 16621
rect 5021 16587 5056 16621
rect 5090 16587 5125 16621
rect 5159 16587 5194 16621
rect 5228 16587 5263 16621
rect 5297 16587 5332 16621
rect 5366 16587 5401 16621
rect 5435 16587 5470 16621
rect 5504 16587 5539 16621
rect 5573 16587 5608 16621
rect 5642 16587 5677 16621
rect 5711 16587 5746 16621
rect 5780 16587 5815 16621
rect 5849 16587 5884 16621
rect 5918 16587 5953 16621
rect 5987 16587 6022 16621
rect 6056 16587 6091 16621
rect 2676 16553 6091 16587
rect 2676 16519 2710 16553
rect 2744 16519 2779 16553
rect 2813 16519 2848 16553
rect 2882 16519 2917 16553
rect 2951 16519 2986 16553
rect 3020 16519 3055 16553
rect 3089 16519 3124 16553
rect 3158 16519 3193 16553
rect 3227 16519 3262 16553
rect 3296 16519 3331 16553
rect 3365 16519 3400 16553
rect 3434 16519 3469 16553
rect 3503 16519 3538 16553
rect 3572 16519 3607 16553
rect 3641 16519 3676 16553
rect 3710 16519 3745 16553
rect 3779 16519 3814 16553
rect 3848 16519 3883 16553
rect 3917 16519 3952 16553
rect 3986 16519 4021 16553
rect 4055 16519 4090 16553
rect 4124 16519 4159 16553
rect 4193 16519 4228 16553
rect 4262 16519 4297 16553
rect 4331 16519 4366 16553
rect 4400 16519 4435 16553
rect 4469 16519 4504 16553
rect 4538 16519 4573 16553
rect 4607 16519 4642 16553
rect 4676 16519 4711 16553
rect 4745 16519 4780 16553
rect 4814 16519 4849 16553
rect 4883 16519 4918 16553
rect 4952 16519 4987 16553
rect 5021 16519 5056 16553
rect 5090 16519 5125 16553
rect 5159 16519 5194 16553
rect 5228 16519 5263 16553
rect 5297 16519 5332 16553
rect 5366 16519 5401 16553
rect 5435 16519 5470 16553
rect 5504 16519 5539 16553
rect 5573 16519 5608 16553
rect 5642 16519 5677 16553
rect 5711 16519 5746 16553
rect 5780 16519 5815 16553
rect 5849 16519 5884 16553
rect 5918 16519 5953 16553
rect 5987 16519 6022 16553
rect 6056 16519 6091 16553
rect 2676 16485 6091 16519
rect 2676 16451 2710 16485
rect 2744 16451 2779 16485
rect 2813 16451 2848 16485
rect 2882 16451 2917 16485
rect 2951 16451 2986 16485
rect 3020 16451 3055 16485
rect 3089 16451 3124 16485
rect 3158 16451 3193 16485
rect 3227 16451 3262 16485
rect 3296 16451 3331 16485
rect 3365 16451 3400 16485
rect 3434 16451 3469 16485
rect 3503 16451 3538 16485
rect 3572 16451 3607 16485
rect 3641 16451 3676 16485
rect 3710 16451 3745 16485
rect 3779 16451 3814 16485
rect 3848 16451 3883 16485
rect 3917 16451 3952 16485
rect 3986 16451 4021 16485
rect 4055 16451 4090 16485
rect 4124 16451 4159 16485
rect 4193 16451 4228 16485
rect 4262 16451 4297 16485
rect 4331 16451 4366 16485
rect 4400 16451 4435 16485
rect 4469 16451 4504 16485
rect 4538 16451 4573 16485
rect 4607 16451 4642 16485
rect 4676 16451 4711 16485
rect 4745 16451 4780 16485
rect 4814 16451 4849 16485
rect 4883 16451 4918 16485
rect 4952 16451 4987 16485
rect 5021 16451 5056 16485
rect 5090 16451 5125 16485
rect 5159 16451 5194 16485
rect 5228 16451 5263 16485
rect 5297 16451 5332 16485
rect 5366 16451 5401 16485
rect 5435 16451 5470 16485
rect 5504 16451 5539 16485
rect 5573 16451 5608 16485
rect 5642 16451 5677 16485
rect 5711 16451 5746 16485
rect 5780 16451 5815 16485
rect 5849 16451 5884 16485
rect 5918 16451 5953 16485
rect 5987 16451 6022 16485
rect 6056 16451 6091 16485
rect 17005 16451 17039 16961
rect 2676 16398 17039 16451
rect -2814 16179 17039 16228
rect -2814 16145 -2732 16179
rect -2698 16145 -2663 16179
rect -2629 16145 -2594 16179
rect -2560 16145 -2525 16179
rect -2491 16145 -2456 16179
rect -2422 16145 -2387 16179
rect -2353 16145 -2318 16179
rect -2284 16145 -2249 16179
rect -2215 16145 -2180 16179
rect -2146 16145 -2111 16179
rect -2077 16145 -2042 16179
rect -2008 16145 -1973 16179
rect -1939 16145 -1904 16179
rect -1870 16145 -1835 16179
rect -1801 16145 -1766 16179
rect -1732 16145 -1697 16179
rect -1663 16145 -1628 16179
rect -1594 16145 -1559 16179
rect -1525 16145 -1490 16179
rect -1456 16145 -1421 16179
rect -1387 16145 -1352 16179
rect -1318 16145 -1283 16179
rect -1249 16145 -1214 16179
rect -1180 16145 -1145 16179
rect -1111 16145 -1076 16179
rect -1042 16145 -1007 16179
rect -973 16145 -938 16179
rect -904 16145 -869 16179
rect -835 16145 -800 16179
rect -766 16145 -731 16179
rect -697 16145 -662 16179
rect -628 16145 -593 16179
rect -559 16145 -524 16179
rect -490 16145 -455 16179
rect -421 16145 -386 16179
rect -352 16145 -317 16179
rect -283 16145 -248 16179
rect -214 16145 -179 16179
rect -145 16145 -110 16179
rect -76 16145 -41 16179
rect -7 16145 28 16179
rect 62 16145 97 16179
rect 131 16145 166 16179
rect 200 16145 235 16179
rect 269 16145 304 16179
rect 338 16145 373 16179
rect 407 16145 442 16179
rect 476 16145 511 16179
rect 545 16145 580 16179
rect 614 16145 649 16179
rect 683 16145 718 16179
rect 17004 16171 17039 16179
rect -2814 16111 718 16145
rect -2814 16077 -2732 16111
rect -2698 16077 -2663 16111
rect -2629 16077 -2594 16111
rect -2560 16077 -2525 16111
rect -2491 16077 -2456 16111
rect -2422 16077 -2387 16111
rect -2353 16077 -2318 16111
rect -2284 16077 -2249 16111
rect -2215 16077 -2180 16111
rect -2146 16077 -2111 16111
rect -2077 16077 -2042 16111
rect -2008 16077 -1973 16111
rect -1939 16077 -1904 16111
rect -1870 16077 -1835 16111
rect -1801 16077 -1766 16111
rect -1732 16077 -1697 16111
rect -1663 16077 -1628 16111
rect -1594 16077 -1559 16111
rect -1525 16077 -1490 16111
rect -1456 16077 -1421 16111
rect -1387 16077 -1352 16111
rect -1318 16077 -1283 16111
rect -1249 16077 -1214 16111
rect -1180 16077 -1145 16111
rect -1111 16077 -1076 16111
rect -1042 16077 -1007 16111
rect -973 16077 -938 16111
rect -904 16077 -869 16111
rect -835 16077 -800 16111
rect -766 16077 -731 16111
rect -697 16077 -662 16111
rect -628 16077 -593 16111
rect -559 16077 -524 16111
rect -490 16077 -455 16111
rect -421 16077 -386 16111
rect -352 16077 -317 16111
rect -283 16077 -248 16111
rect -214 16077 -179 16111
rect -145 16077 -110 16111
rect -76 16077 -41 16111
rect -7 16077 28 16111
rect 62 16077 97 16111
rect 131 16077 166 16111
rect 200 16077 235 16111
rect 269 16077 304 16111
rect 338 16077 373 16111
rect 407 16077 442 16111
rect 476 16077 511 16111
rect 545 16077 580 16111
rect 614 16077 649 16111
rect 683 16077 718 16111
rect -2814 16043 718 16077
rect -2814 16009 -2732 16043
rect -2698 16009 -2663 16043
rect -2629 16009 -2594 16043
rect -2560 16009 -2525 16043
rect -2491 16009 -2456 16043
rect -2422 16009 -2387 16043
rect -2353 16009 -2318 16043
rect -2284 16009 -2249 16043
rect -2215 16009 -2180 16043
rect -2146 16009 -2111 16043
rect -2077 16009 -2042 16043
rect -2008 16009 -1973 16043
rect -1939 16009 -1904 16043
rect -1870 16009 -1835 16043
rect -1801 16009 -1766 16043
rect -1732 16009 -1697 16043
rect -1663 16009 -1628 16043
rect -1594 16009 -1559 16043
rect -1525 16009 -1490 16043
rect -1456 16009 -1421 16043
rect -1387 16009 -1352 16043
rect -1318 16009 -1283 16043
rect -1249 16009 -1214 16043
rect -1180 16009 -1145 16043
rect -1111 16009 -1076 16043
rect -1042 16009 -1007 16043
rect -973 16009 -938 16043
rect -904 16009 -869 16043
rect -835 16009 -800 16043
rect -766 16009 -731 16043
rect -697 16009 -662 16043
rect -628 16009 -593 16043
rect -559 16009 -524 16043
rect -490 16009 -455 16043
rect -421 16009 -386 16043
rect -352 16009 -317 16043
rect -283 16009 -248 16043
rect -214 16009 -179 16043
rect -145 16009 -110 16043
rect -76 16009 -41 16043
rect -7 16009 28 16043
rect 62 16009 97 16043
rect 131 16009 166 16043
rect 200 16009 235 16043
rect 269 16009 304 16043
rect 338 16009 373 16043
rect 407 16009 442 16043
rect 476 16009 511 16043
rect 545 16009 580 16043
rect 614 16009 649 16043
rect 683 16009 718 16043
rect -2814 15975 718 16009
rect -2814 15941 -2732 15975
rect -2698 15941 -2663 15975
rect -2629 15941 -2594 15975
rect -2560 15941 -2525 15975
rect -2491 15941 -2456 15975
rect -2422 15941 -2387 15975
rect -2353 15941 -2318 15975
rect -2284 15941 -2249 15975
rect -2215 15941 -2180 15975
rect -2146 15941 -2111 15975
rect -2077 15941 -2042 15975
rect -2008 15941 -1973 15975
rect -1939 15941 -1904 15975
rect -1870 15941 -1835 15975
rect -1801 15941 -1766 15975
rect -1732 15941 -1697 15975
rect -1663 15941 -1628 15975
rect -1594 15941 -1559 15975
rect -1525 15941 -1490 15975
rect -1456 15941 -1421 15975
rect -1387 15941 -1352 15975
rect -1318 15941 -1283 15975
rect -1249 15941 -1214 15975
rect -1180 15941 -1145 15975
rect -1111 15941 -1076 15975
rect -1042 15941 -1007 15975
rect -973 15941 -938 15975
rect -904 15941 -869 15975
rect -835 15941 -800 15975
rect -766 15941 -731 15975
rect -697 15941 -662 15975
rect -628 15941 -593 15975
rect -559 15941 -524 15975
rect -490 15941 -455 15975
rect -421 15941 -386 15975
rect -352 15941 -317 15975
rect -283 15941 -248 15975
rect -214 15941 -179 15975
rect -145 15941 -110 15975
rect -76 15941 -41 15975
rect -7 15941 28 15975
rect 62 15941 97 15975
rect 131 15941 166 15975
rect 200 15941 235 15975
rect 269 15941 304 15975
rect 338 15941 373 15975
rect 407 15941 442 15975
rect 476 15941 511 15975
rect 545 15941 580 15975
rect 614 15941 649 15975
rect 683 15941 718 15975
rect -2814 15907 718 15941
rect 17018 15921 17039 16171
rect -2814 15873 -2732 15907
rect -2698 15873 -2663 15907
rect -2629 15873 -2594 15907
rect -2560 15873 -2525 15907
rect -2491 15873 -2456 15907
rect -2422 15873 -2387 15907
rect -2353 15873 -2318 15907
rect -2284 15873 -2249 15907
rect -2215 15873 -2180 15907
rect -2146 15873 -2111 15907
rect -2077 15873 -2042 15907
rect -2008 15873 -1973 15907
rect -1939 15873 -1904 15907
rect -1870 15873 -1835 15907
rect -1801 15873 -1766 15907
rect -1732 15873 -1697 15907
rect -1663 15873 -1628 15907
rect -1594 15873 -1559 15907
rect -1525 15873 -1490 15907
rect -1456 15873 -1421 15907
rect -1387 15873 -1352 15907
rect -1318 15873 -1283 15907
rect -1249 15873 -1214 15907
rect -1180 15873 -1145 15907
rect -1111 15873 -1076 15907
rect -1042 15873 -1007 15907
rect -973 15873 -938 15907
rect -904 15873 -869 15907
rect -835 15873 -800 15907
rect -766 15873 -731 15907
rect -697 15873 -662 15907
rect -628 15873 -593 15907
rect -559 15873 -524 15907
rect -490 15873 -455 15907
rect -421 15873 -386 15907
rect -352 15873 -317 15907
rect -283 15873 -248 15907
rect -214 15873 -179 15907
rect -145 15873 -110 15907
rect -76 15873 -41 15907
rect -7 15873 28 15907
rect 62 15873 97 15907
rect 131 15873 166 15907
rect 200 15873 235 15907
rect 269 15873 304 15907
rect 338 15873 373 15907
rect 407 15873 442 15907
rect 476 15873 511 15907
rect 545 15873 580 15907
rect 614 15873 649 15907
rect 683 15873 718 15907
rect -2814 15839 718 15873
rect -2814 15805 -2732 15839
rect -2698 15805 -2663 15839
rect -2629 15805 -2594 15839
rect -2560 15805 -2525 15839
rect -2491 15805 -2456 15839
rect -2422 15805 -2387 15839
rect -2353 15805 -2318 15839
rect -2284 15805 -2249 15839
rect -2215 15805 -2180 15839
rect -2146 15805 -2111 15839
rect -2077 15805 -2042 15839
rect -2008 15805 -1973 15839
rect -1939 15805 -1904 15839
rect -1870 15805 -1835 15839
rect -1801 15805 -1766 15839
rect -1732 15805 -1697 15839
rect -1663 15805 -1628 15839
rect -1594 15805 -1559 15839
rect -1525 15805 -1490 15839
rect -1456 15805 -1421 15839
rect -1387 15805 -1352 15839
rect -1318 15805 -1283 15839
rect -1249 15805 -1214 15839
rect -1180 15805 -1145 15839
rect -1111 15805 -1076 15839
rect -1042 15805 -1007 15839
rect -973 15805 -938 15839
rect -904 15805 -869 15839
rect -835 15805 -800 15839
rect -766 15805 -731 15839
rect -697 15805 -662 15839
rect -628 15805 -593 15839
rect -559 15805 -524 15839
rect -490 15805 -455 15839
rect -421 15805 -386 15839
rect -352 15805 -317 15839
rect -283 15805 -248 15839
rect -214 15805 -179 15839
rect -145 15805 -110 15839
rect -76 15805 -41 15839
rect -7 15805 28 15839
rect 62 15805 97 15839
rect 131 15805 166 15839
rect 200 15805 235 15839
rect 269 15805 304 15839
rect 338 15805 373 15839
rect 407 15805 442 15839
rect 476 15805 511 15839
rect 545 15805 580 15839
rect 614 15805 649 15839
rect 683 15805 718 15839
rect -2814 15771 718 15805
rect -2814 15737 -2732 15771
rect -2698 15737 -2663 15771
rect -2629 15737 -2594 15771
rect -2560 15737 -2525 15771
rect -2491 15737 -2456 15771
rect -2422 15737 -2387 15771
rect -2353 15737 -2318 15771
rect -2284 15737 -2249 15771
rect -2215 15737 -2180 15771
rect -2146 15737 -2111 15771
rect -2077 15737 -2042 15771
rect -2008 15737 -1973 15771
rect -1939 15737 -1904 15771
rect -1870 15737 -1835 15771
rect -1801 15737 -1766 15771
rect -1732 15737 -1697 15771
rect -1663 15737 -1628 15771
rect -1594 15737 -1559 15771
rect -1525 15737 -1490 15771
rect -1456 15737 -1421 15771
rect -1387 15737 -1352 15771
rect -1318 15737 -1283 15771
rect -1249 15737 -1214 15771
rect -1180 15737 -1145 15771
rect -1111 15737 -1076 15771
rect -1042 15737 -1007 15771
rect -973 15737 -938 15771
rect -904 15737 -869 15771
rect -835 15737 -800 15771
rect -766 15737 -731 15771
rect -697 15737 -662 15771
rect -628 15737 -593 15771
rect -559 15737 -524 15771
rect -490 15737 -455 15771
rect -421 15737 -386 15771
rect -352 15737 -317 15771
rect -283 15737 -248 15771
rect -214 15737 -179 15771
rect -145 15737 -110 15771
rect -76 15737 -41 15771
rect -7 15737 28 15771
rect 62 15737 97 15771
rect 131 15737 166 15771
rect 200 15737 235 15771
rect 269 15737 304 15771
rect 338 15737 373 15771
rect 407 15737 442 15771
rect 476 15737 511 15771
rect 545 15737 580 15771
rect 614 15737 649 15771
rect 683 15737 718 15771
rect -2814 15703 718 15737
rect -2814 15669 -2732 15703
rect -2698 15669 -2663 15703
rect -2629 15669 -2594 15703
rect -2560 15669 -2525 15703
rect -2491 15669 -2456 15703
rect -2422 15669 -2387 15703
rect -2353 15669 -2318 15703
rect -2284 15669 -2249 15703
rect -2215 15669 -2180 15703
rect -2146 15669 -2111 15703
rect -2077 15669 -2042 15703
rect -2008 15669 -1973 15703
rect -1939 15669 -1904 15703
rect -1870 15669 -1835 15703
rect -1801 15669 -1766 15703
rect -1732 15669 -1697 15703
rect -1663 15669 -1628 15703
rect -1594 15669 -1559 15703
rect -1525 15669 -1490 15703
rect -1456 15669 -1421 15703
rect -1387 15669 -1352 15703
rect -1318 15669 -1283 15703
rect -1249 15669 -1214 15703
rect -1180 15669 -1145 15703
rect -1111 15669 -1076 15703
rect -1042 15669 -1007 15703
rect -973 15669 -938 15703
rect -904 15669 -869 15703
rect -835 15669 -800 15703
rect -766 15669 -731 15703
rect -697 15669 -662 15703
rect -628 15669 -593 15703
rect -559 15669 -524 15703
rect -490 15669 -455 15703
rect -421 15669 -386 15703
rect -352 15669 -317 15703
rect -283 15669 -248 15703
rect -214 15669 -179 15703
rect -145 15669 -110 15703
rect -76 15669 -41 15703
rect -7 15669 28 15703
rect 62 15669 97 15703
rect 131 15669 166 15703
rect 200 15669 235 15703
rect 269 15669 304 15703
rect 338 15669 373 15703
rect 407 15669 442 15703
rect 476 15669 511 15703
rect 545 15669 580 15703
rect 614 15669 649 15703
rect 683 15669 718 15703
rect -2814 15635 718 15669
rect -2814 15601 -2732 15635
rect -2698 15601 -2663 15635
rect -2629 15601 -2594 15635
rect -2560 15601 -2525 15635
rect -2491 15601 -2456 15635
rect -2422 15601 -2387 15635
rect -2353 15601 -2318 15635
rect -2284 15601 -2249 15635
rect -2215 15601 -2180 15635
rect -2146 15601 -2111 15635
rect -2077 15601 -2042 15635
rect -2008 15601 -1973 15635
rect -1939 15601 -1904 15635
rect -1870 15601 -1835 15635
rect -1801 15601 -1766 15635
rect -1732 15601 -1697 15635
rect -1663 15601 -1628 15635
rect -1594 15601 -1559 15635
rect -1525 15601 -1490 15635
rect -1456 15601 -1421 15635
rect -1387 15601 -1352 15635
rect -1318 15601 -1283 15635
rect -1249 15601 -1214 15635
rect -1180 15601 -1145 15635
rect -1111 15601 -1076 15635
rect -1042 15601 -1007 15635
rect -973 15601 -938 15635
rect -904 15601 -869 15635
rect -835 15601 -800 15635
rect -766 15601 -731 15635
rect -697 15601 -662 15635
rect -628 15601 -593 15635
rect -559 15601 -524 15635
rect -490 15601 -455 15635
rect -421 15601 -386 15635
rect -352 15601 -317 15635
rect -283 15601 -248 15635
rect -214 15601 -179 15635
rect -145 15601 -110 15635
rect -76 15601 -41 15635
rect -7 15601 28 15635
rect 62 15601 97 15635
rect 131 15601 166 15635
rect 200 15601 235 15635
rect 269 15601 304 15635
rect 338 15601 373 15635
rect 407 15601 442 15635
rect 476 15601 511 15635
rect 545 15601 580 15635
rect 614 15601 649 15635
rect 683 15601 718 15635
rect -2814 15567 718 15601
rect -2814 15533 -2732 15567
rect -2698 15533 -2663 15567
rect -2629 15533 -2594 15567
rect -2560 15533 -2525 15567
rect -2491 15533 -2456 15567
rect -2422 15533 -2387 15567
rect -2353 15533 -2318 15567
rect -2284 15533 -2249 15567
rect -2215 15533 -2180 15567
rect -2146 15533 -2111 15567
rect -2077 15533 -2042 15567
rect -2008 15533 -1973 15567
rect -1939 15533 -1904 15567
rect -1870 15533 -1835 15567
rect -1801 15533 -1766 15567
rect -1732 15533 -1697 15567
rect -1663 15533 -1628 15567
rect -1594 15533 -1559 15567
rect -1525 15533 -1490 15567
rect -1456 15533 -1421 15567
rect -1387 15533 -1352 15567
rect -1318 15533 -1283 15567
rect -1249 15533 -1214 15567
rect -1180 15533 -1145 15567
rect -1111 15533 -1076 15567
rect -1042 15533 -1007 15567
rect -973 15533 -938 15567
rect -904 15533 -869 15567
rect -835 15533 -800 15567
rect -766 15533 -731 15567
rect -697 15533 -662 15567
rect -628 15533 -593 15567
rect -559 15533 -524 15567
rect -490 15533 -455 15567
rect -421 15533 -386 15567
rect -352 15533 -317 15567
rect -283 15533 -248 15567
rect -214 15533 -179 15567
rect -145 15533 -110 15567
rect -76 15533 -41 15567
rect -7 15533 28 15567
rect 62 15533 97 15567
rect 131 15533 166 15567
rect 200 15533 235 15567
rect 269 15533 304 15567
rect 338 15533 373 15567
rect 407 15533 442 15567
rect 476 15533 511 15567
rect 545 15533 580 15567
rect 614 15533 649 15567
rect 683 15533 718 15567
rect -2814 15499 718 15533
rect -2814 15465 -2732 15499
rect -2698 15465 -2663 15499
rect -2629 15465 -2594 15499
rect -2560 15465 -2525 15499
rect -2491 15465 -2456 15499
rect -2422 15465 -2387 15499
rect -2353 15465 -2318 15499
rect -2284 15465 -2249 15499
rect -2215 15465 -2180 15499
rect -2146 15465 -2111 15499
rect -2077 15465 -2042 15499
rect -2008 15465 -1973 15499
rect -1939 15465 -1904 15499
rect -1870 15465 -1835 15499
rect -1801 15465 -1766 15499
rect -1732 15465 -1697 15499
rect -1663 15465 -1628 15499
rect -1594 15465 -1559 15499
rect -1525 15465 -1490 15499
rect -1456 15465 -1421 15499
rect -1387 15465 -1352 15499
rect -1318 15465 -1283 15499
rect -1249 15465 -1214 15499
rect -1180 15465 -1145 15499
rect -1111 15465 -1076 15499
rect -1042 15465 -1007 15499
rect -973 15465 -938 15499
rect -904 15465 -869 15499
rect -835 15465 -800 15499
rect -766 15465 -731 15499
rect -697 15465 -662 15499
rect -628 15465 -593 15499
rect -559 15465 -524 15499
rect -490 15465 -455 15499
rect -421 15465 -386 15499
rect -352 15465 -317 15499
rect -283 15465 -248 15499
rect -214 15465 -179 15499
rect -145 15465 -110 15499
rect -76 15465 -41 15499
rect -7 15465 28 15499
rect 62 15465 97 15499
rect 131 15465 166 15499
rect 200 15465 235 15499
rect 269 15465 304 15499
rect 338 15465 373 15499
rect 407 15465 442 15499
rect 476 15465 511 15499
rect 545 15465 580 15499
rect 614 15465 649 15499
rect 683 15465 718 15499
rect -2814 15431 718 15465
rect -2814 15397 -2732 15431
rect -2698 15397 -2663 15431
rect -2629 15397 -2594 15431
rect -2560 15397 -2525 15431
rect -2491 15397 -2456 15431
rect -2422 15397 -2387 15431
rect -2353 15397 -2318 15431
rect -2284 15397 -2249 15431
rect -2215 15397 -2180 15431
rect -2146 15397 -2111 15431
rect -2077 15397 -2042 15431
rect -2008 15397 -1973 15431
rect -1939 15397 -1904 15431
rect -1870 15397 -1835 15431
rect -1801 15397 -1766 15431
rect -1732 15397 -1697 15431
rect -1663 15397 -1628 15431
rect -1594 15397 -1559 15431
rect -1525 15397 -1490 15431
rect -1456 15397 -1421 15431
rect -1387 15397 -1352 15431
rect -1318 15397 -1283 15431
rect -1249 15397 -1214 15431
rect -1180 15397 -1145 15431
rect -1111 15397 -1076 15431
rect -1042 15397 -1007 15431
rect -973 15397 -938 15431
rect -904 15397 -869 15431
rect -835 15397 -800 15431
rect -766 15397 -731 15431
rect -697 15397 -662 15431
rect -628 15397 -593 15431
rect -559 15397 -524 15431
rect -490 15397 -455 15431
rect -421 15397 -386 15431
rect -352 15397 -317 15431
rect -283 15397 -248 15431
rect -214 15397 -179 15431
rect -145 15397 -110 15431
rect -76 15397 -41 15431
rect -7 15397 28 15431
rect 62 15397 97 15431
rect 131 15397 166 15431
rect 200 15397 235 15431
rect 269 15397 304 15431
rect 338 15397 373 15431
rect 407 15397 442 15431
rect 476 15397 511 15431
rect 545 15397 580 15431
rect 614 15397 649 15431
rect 683 15397 718 15431
rect 17004 15397 17039 15921
rect -2814 15380 17039 15397
rect 10855 3498 11477 3500
rect 138 3448 308 3498
rect 1873 3489 11477 3498
rect 172 3414 206 3448
rect 240 3414 274 3448
rect 138 3378 308 3414
rect 172 3344 206 3378
rect 240 3344 274 3378
rect 138 3308 308 3344
rect 172 3274 206 3308
rect 240 3274 274 3308
rect 138 3238 308 3274
rect 172 3204 206 3238
rect 240 3204 274 3238
rect 138 3168 308 3204
rect 172 3134 206 3168
rect 240 3134 274 3168
rect 138 3098 308 3134
rect 172 3064 206 3098
rect 240 3064 274 3098
rect 138 3028 308 3064
rect 172 2994 206 3028
rect 240 2994 274 3028
rect 138 2958 308 2994
rect 1873 3448 2043 3472
rect 1907 3414 1941 3448
rect 1975 3414 2009 3448
rect 1873 3379 2043 3414
rect 1907 3345 1941 3379
rect 1975 3345 2009 3379
rect 1873 3310 2043 3345
rect 1907 3276 1941 3310
rect 1975 3276 2009 3310
rect 1873 3241 2043 3276
rect 1907 3207 1941 3241
rect 1975 3207 2009 3241
rect 1873 3172 2043 3207
rect 1907 3138 1941 3172
rect 1975 3138 2009 3172
rect 1873 3103 2043 3138
rect 1907 3069 1941 3103
rect 1975 3069 2009 3103
rect 1873 3034 2043 3069
rect 1907 3000 1941 3034
rect 1975 3000 2009 3034
rect 172 2924 206 2958
rect 240 2924 274 2958
rect 138 2888 308 2924
rect 172 2854 206 2888
rect 240 2854 274 2888
rect 138 2818 308 2854
rect 172 2784 206 2818
rect 240 2784 274 2818
rect 138 2749 308 2784
rect 172 2715 206 2749
rect 240 2748 308 2749
rect 240 2715 274 2748
rect 138 2714 274 2715
rect 138 2680 308 2714
rect 172 2646 206 2680
rect 240 2678 308 2680
rect 240 2646 274 2678
rect 138 2644 274 2646
rect 138 2611 308 2644
rect 172 2577 206 2611
rect 240 2609 308 2611
rect 240 2577 274 2609
rect 138 2575 274 2577
rect 138 2542 308 2575
rect 172 2508 206 2542
rect 240 2540 308 2542
rect 240 2508 274 2540
rect 138 2506 274 2508
rect 138 2473 308 2506
rect 172 2439 206 2473
rect 240 2471 308 2473
rect 240 2439 274 2471
rect 138 2437 274 2439
rect 138 2404 308 2437
rect 172 2370 206 2404
rect 240 2402 308 2404
rect 240 2370 274 2402
rect 138 2368 274 2370
rect 138 2335 308 2368
rect 172 2301 206 2335
rect 240 2333 308 2335
rect 240 2301 274 2333
rect 138 2299 274 2301
rect 138 2266 308 2299
rect 172 2232 206 2266
rect 240 2264 308 2266
rect 240 2232 274 2264
rect 138 2230 274 2232
rect 138 2197 308 2230
rect 172 2163 206 2197
rect 240 2195 308 2197
rect 240 2163 274 2195
rect 138 2161 274 2163
rect 138 2128 308 2161
rect 172 2094 206 2128
rect 240 2126 308 2128
rect 240 2094 274 2126
rect 138 2092 274 2094
rect 138 2059 308 2092
rect 172 2025 206 2059
rect 240 2057 308 2059
rect 240 2025 274 2057
rect 138 2023 274 2025
rect 138 1990 308 2023
rect 172 1956 206 1990
rect 240 1988 308 1990
rect 240 1956 274 1988
rect 138 1954 274 1956
rect 138 1921 308 1954
rect 172 1887 206 1921
rect 240 1919 308 1921
rect 240 1887 274 1919
rect 138 1885 274 1887
rect 138 1852 308 1885
rect 172 1818 206 1852
rect 240 1850 308 1852
rect 240 1818 274 1850
rect 138 1816 274 1818
rect 138 1783 308 1816
rect 172 1749 206 1783
rect 240 1781 308 1783
rect 240 1749 274 1781
rect 138 1747 274 1749
rect 138 1714 308 1747
rect 172 1680 206 1714
rect 240 1712 308 1714
rect 240 1680 274 1712
rect 138 1678 274 1680
rect 138 1645 308 1678
rect 172 1611 206 1645
rect 240 1643 308 1645
rect 240 1611 274 1643
rect 138 1609 274 1611
rect 138 1576 308 1609
rect 172 1542 206 1576
rect 240 1574 308 1576
rect 240 1542 274 1574
rect 138 1540 274 1542
rect 138 1507 308 1540
rect 172 1473 206 1507
rect 240 1505 308 1507
rect 240 1473 274 1505
rect 138 1471 274 1473
rect 138 1438 308 1471
rect 172 1404 206 1438
rect 240 1436 308 1438
rect 240 1404 274 1436
rect 138 1402 274 1404
rect 138 1369 308 1402
rect 172 1335 206 1369
rect 240 1367 308 1369
rect 240 1335 274 1367
rect 138 1333 274 1335
rect 138 1300 308 1333
rect 470 2188 640 2212
rect 504 2154 538 2188
rect 572 2154 606 2188
rect 470 2118 640 2154
rect 470 2115 538 2118
rect 504 2084 538 2115
rect 572 2084 606 2118
rect 504 2081 640 2084
rect 470 2048 640 2081
rect 470 2042 538 2048
rect 504 2014 538 2042
rect 572 2014 606 2048
rect 504 2008 640 2014
rect 470 1978 640 2008
rect 470 1969 538 1978
rect 504 1944 538 1969
rect 572 1944 606 1978
rect 504 1935 640 1944
rect 470 1908 640 1935
rect 470 1896 538 1908
rect 504 1874 538 1896
rect 572 1874 606 1908
rect 504 1862 640 1874
rect 470 1838 640 1862
rect 470 1823 538 1838
rect 504 1804 538 1823
rect 572 1804 606 1838
rect 504 1789 640 1804
rect 470 1768 640 1789
rect 470 1750 538 1768
rect 504 1734 538 1750
rect 572 1734 606 1768
rect 504 1716 640 1734
rect 470 1698 640 1716
rect 470 1677 538 1698
rect 504 1664 538 1677
rect 572 1664 606 1698
rect 504 1643 640 1664
rect 470 1628 640 1643
rect 470 1604 538 1628
rect 504 1594 538 1604
rect 572 1594 606 1628
rect 676 2176 737 2979
rect 1873 2965 2043 3000
rect 1907 2931 1941 2965
rect 1975 2931 2009 2965
rect 1873 2896 2043 2931
rect 1616 2854 1654 2888
rect 1582 2815 1688 2854
rect 1582 2813 1654 2815
rect 1616 2781 1654 2813
rect 1616 2779 1688 2781
rect 1582 2742 1688 2779
rect 1582 2738 1654 2742
rect 1616 2708 1654 2738
rect 1616 2704 1688 2708
rect 1582 2669 1688 2704
rect 1582 2663 1654 2669
rect 1616 2635 1654 2663
rect 1616 2629 1688 2635
rect 1582 2596 1688 2629
rect 1582 2588 1654 2596
rect 1616 2562 1654 2588
rect 1616 2554 1688 2562
rect 1582 2523 1688 2554
rect 1582 2513 1654 2523
rect 1616 2489 1654 2513
rect 1616 2479 1688 2489
rect 1582 2450 1688 2479
rect 1582 2438 1654 2450
rect 1616 2416 1654 2438
rect 1616 2404 1688 2416
rect 1582 2377 1688 2404
rect 1582 2363 1654 2377
rect 1616 2343 1654 2363
rect 1616 2329 1688 2343
rect 1582 2304 1688 2329
rect 1582 2288 1654 2304
rect 1616 2270 1654 2288
rect 1616 2254 1688 2270
rect 1582 2231 1688 2254
rect 1582 2213 1654 2231
rect 1550 2188 1582 2212
rect 1616 2197 1654 2213
rect 1907 2862 1941 2896
rect 1975 2862 2009 2896
rect 1873 2827 2043 2862
rect 1907 2793 1941 2827
rect 1975 2793 2009 2827
rect 1873 2758 2043 2793
rect 1907 2724 1941 2758
rect 1975 2724 2009 2758
rect 1873 2689 2043 2724
rect 1907 2655 1941 2689
rect 1975 2655 2009 2689
rect 1873 2620 2043 2655
rect 1907 2586 1941 2620
rect 1975 2586 2009 2620
rect 1873 2551 2043 2586
rect 1907 2517 1941 2551
rect 1975 2517 2009 2551
rect 1873 2482 2043 2517
rect 1907 2448 1941 2482
rect 1975 2448 2009 2482
rect 1873 2413 2043 2448
rect 1907 2379 1941 2413
rect 1975 2379 2009 2413
rect 1873 2344 2043 2379
rect 1907 2310 1941 2344
rect 1975 2310 2009 2344
rect 4227 3461 11477 3489
rect 4227 2335 4284 3461
rect 10855 2498 11477 3461
rect 1873 2275 2043 2310
rect 1907 2241 1941 2275
rect 1975 2241 2009 2275
rect 1688 2197 1720 2212
rect 1616 2188 1720 2197
rect 676 2142 686 2176
rect 720 2142 737 2176
rect 820 2146 861 2180
rect 895 2146 936 2180
rect 970 2146 1010 2180
rect 1044 2146 1084 2180
rect 1118 2146 1158 2180
rect 1192 2146 1232 2180
rect 1266 2146 1306 2180
rect 1616 2179 1618 2188
rect 1584 2154 1618 2179
rect 1652 2158 1686 2188
rect 1652 2154 1654 2158
rect 676 2104 737 2142
rect 676 2070 686 2104
rect 720 2092 737 2104
rect 676 2058 688 2070
rect 722 2058 737 2092
rect 676 2024 737 2058
rect 1550 2138 1654 2154
rect 1550 2117 1582 2138
rect 1616 2124 1654 2138
rect 1688 2124 1720 2154
rect 1616 2118 1720 2124
rect 1616 2104 1618 2118
rect 1584 2084 1618 2104
rect 1652 2115 1720 2118
rect 1652 2085 1686 2115
rect 1652 2084 1654 2085
rect 1584 2083 1654 2084
rect 1550 2062 1654 2083
rect 1550 2046 1582 2062
rect 1616 2051 1654 2062
rect 1688 2051 1720 2081
rect 1616 2048 1720 2051
rect 1616 2028 1618 2048
rect 676 1990 688 2024
rect 722 1990 737 2024
rect 813 1990 855 2024
rect 889 1990 931 2024
rect 965 1990 1007 2024
rect 1041 1990 1083 2024
rect 1117 1990 1159 2024
rect 1193 1990 1234 2024
rect 1584 2014 1618 2028
rect 1652 2042 1720 2048
rect 1652 2014 1686 2042
rect 1584 2012 1686 2014
rect 676 1956 737 1990
rect 676 1922 688 1956
rect 722 1922 737 1956
rect 676 1713 737 1922
rect 1550 1986 1654 2012
rect 1550 1976 1582 1986
rect 1616 1978 1654 1986
rect 1688 1978 1720 2008
rect 1616 1952 1618 1978
rect 1584 1944 1618 1952
rect 1652 1969 1720 1978
rect 1652 1944 1686 1969
rect 1584 1942 1686 1944
rect 1550 1938 1686 1942
rect 1550 1910 1654 1938
rect 1550 1906 1582 1910
rect 1616 1908 1654 1910
rect 1616 1876 1618 1908
rect 1584 1874 1618 1876
rect 1652 1904 1654 1908
rect 1688 1904 1720 1935
rect 1652 1896 1720 1904
rect 1652 1874 1686 1896
rect 1584 1872 1686 1874
rect 814 1834 856 1868
rect 890 1834 931 1868
rect 965 1834 1006 1868
rect 1040 1834 1081 1868
rect 1115 1834 1156 1868
rect 1190 1834 1231 1868
rect 1265 1834 1306 1868
rect 1550 1864 1686 1872
rect 1550 1838 1654 1864
rect 1550 1836 1618 1838
rect 1584 1834 1618 1836
rect 1616 1804 1618 1834
rect 1652 1830 1654 1838
rect 1688 1830 1720 1862
rect 1652 1823 1720 1830
rect 1652 1804 1686 1823
rect 1550 1800 1582 1802
rect 1616 1800 1686 1804
rect 1550 1790 1686 1800
rect 1550 1768 1654 1790
rect 1550 1766 1618 1768
rect 1584 1758 1618 1766
rect 820 1724 861 1758
rect 895 1724 936 1758
rect 970 1724 1010 1758
rect 1044 1724 1084 1758
rect 1118 1724 1158 1758
rect 1192 1724 1232 1758
rect 1266 1724 1306 1758
rect 1616 1734 1618 1758
rect 1652 1756 1654 1768
rect 1688 1756 1720 1789
rect 1652 1750 1720 1756
rect 1652 1734 1686 1750
rect 1550 1724 1582 1732
rect 1616 1724 1686 1734
rect 676 1679 688 1713
rect 722 1679 737 1713
rect 676 1645 737 1679
rect 676 1611 688 1645
rect 722 1611 737 1645
rect 676 1594 737 1611
rect 1550 1716 1686 1724
rect 1550 1698 1654 1716
rect 1550 1696 1618 1698
rect 1584 1682 1618 1696
rect 1616 1664 1618 1682
rect 1652 1682 1654 1698
rect 1688 1682 1720 1716
rect 1652 1677 1720 1682
rect 1652 1664 1686 1677
rect 1550 1648 1582 1662
rect 1616 1648 1686 1664
rect 1550 1643 1686 1648
rect 1550 1642 1720 1643
rect 1550 1628 1654 1642
rect 1550 1626 1618 1628
rect 1584 1606 1618 1626
rect 504 1570 640 1594
rect 470 1558 640 1570
rect 820 1568 861 1602
rect 895 1568 936 1602
rect 970 1568 1010 1602
rect 1044 1568 1084 1602
rect 1118 1568 1158 1602
rect 1192 1568 1232 1602
rect 1266 1568 1306 1602
rect 1616 1594 1618 1606
rect 1652 1608 1654 1628
rect 1688 1608 1720 1642
rect 1652 1604 1720 1608
rect 1652 1594 1686 1604
rect 1550 1572 1582 1592
rect 1616 1572 1686 1594
rect 1550 1570 1686 1572
rect 1550 1568 1720 1570
rect 470 1531 538 1558
rect 504 1524 538 1531
rect 572 1557 640 1558
rect 572 1524 606 1557
rect 504 1523 606 1524
rect 504 1511 640 1523
rect 470 1477 502 1497
rect 536 1488 640 1511
rect 536 1477 538 1488
rect 470 1458 538 1477
rect 504 1454 538 1458
rect 572 1486 640 1488
rect 1550 1558 1654 1568
rect 1550 1556 1618 1558
rect 1584 1530 1618 1556
rect 1616 1524 1618 1530
rect 1652 1534 1654 1558
rect 1688 1534 1720 1568
rect 1652 1532 1720 1534
rect 1652 1524 1686 1532
rect 1550 1496 1582 1522
rect 1616 1498 1686 1524
rect 1616 1496 1720 1498
rect 1550 1494 1720 1496
rect 1550 1488 1654 1494
rect 1550 1486 1618 1488
rect 572 1454 606 1486
rect 640 1454 678 1486
rect 712 1454 750 1486
rect 784 1454 822 1486
rect 856 1454 894 1486
rect 928 1454 966 1486
rect 1000 1454 1039 1486
rect 1073 1454 1112 1486
rect 504 1424 574 1454
rect 640 1452 646 1454
rect 712 1452 718 1454
rect 784 1452 790 1454
rect 856 1452 862 1454
rect 928 1452 934 1454
rect 1000 1452 1006 1454
rect 1073 1452 1078 1454
rect 470 1420 574 1424
rect 608 1420 646 1452
rect 680 1420 718 1452
rect 752 1420 790 1452
rect 824 1420 862 1452
rect 896 1420 934 1452
rect 968 1420 1006 1452
rect 1040 1420 1078 1452
rect 1146 1454 1185 1486
rect 1146 1452 1150 1454
rect 1112 1420 1150 1452
rect 1184 1452 1185 1454
rect 1219 1454 1258 1486
rect 1219 1452 1222 1454
rect 1184 1420 1222 1452
rect 1256 1452 1258 1454
rect 1292 1454 1331 1486
rect 1292 1452 1294 1454
rect 1256 1420 1294 1452
rect 1328 1452 1331 1454
rect 1365 1454 1404 1486
rect 1365 1452 1366 1454
rect 1328 1420 1366 1452
rect 1400 1452 1404 1454
rect 1438 1454 1477 1486
rect 1511 1454 1550 1486
rect 1584 1454 1618 1486
rect 1652 1460 1654 1488
rect 1688 1460 1720 1494
rect 1652 1454 1686 1460
rect 1400 1420 1438 1452
rect 1472 1452 1477 1454
rect 1544 1452 1550 1454
rect 1472 1420 1510 1452
rect 1544 1420 1582 1452
rect 1616 1426 1686 1454
rect 1616 1420 1720 1426
rect 470 1418 1654 1420
rect 470 1384 538 1418
rect 572 1384 610 1418
rect 644 1384 682 1418
rect 716 1384 754 1418
rect 788 1384 826 1418
rect 860 1384 898 1418
rect 932 1384 970 1418
rect 1004 1384 1042 1418
rect 1076 1384 1114 1418
rect 1148 1384 1186 1418
rect 1220 1384 1258 1418
rect 1292 1384 1330 1418
rect 1364 1384 1402 1418
rect 1436 1384 1474 1418
rect 1508 1384 1546 1418
rect 1580 1384 1618 1418
rect 1652 1386 1654 1418
rect 1688 1386 1720 1420
rect 1652 1384 1720 1386
rect 504 1382 1720 1384
rect 504 1350 540 1382
rect 470 1348 540 1350
rect 574 1350 617 1382
rect 651 1350 694 1382
rect 728 1350 771 1382
rect 805 1350 848 1382
rect 882 1350 925 1382
rect 959 1350 1002 1382
rect 1036 1350 1079 1382
rect 1113 1350 1156 1382
rect 1190 1350 1232 1382
rect 1266 1350 1308 1382
rect 1342 1350 1384 1382
rect 1418 1350 1460 1382
rect 1494 1350 1536 1382
rect 1570 1350 1720 1382
rect 574 1348 578 1350
rect 470 1316 578 1348
rect 612 1348 617 1350
rect 683 1348 694 1350
rect 754 1348 771 1350
rect 825 1348 848 1350
rect 896 1348 925 1350
rect 967 1348 1002 1350
rect 612 1316 649 1348
rect 683 1316 720 1348
rect 754 1316 791 1348
rect 825 1316 862 1348
rect 896 1316 933 1348
rect 967 1316 1004 1348
rect 1038 1316 1076 1350
rect 1113 1348 1148 1350
rect 1190 1348 1220 1350
rect 1266 1348 1292 1350
rect 1342 1348 1364 1350
rect 1418 1348 1436 1350
rect 1494 1348 1508 1350
rect 1570 1348 1580 1350
rect 1110 1316 1148 1348
rect 1182 1316 1220 1348
rect 1254 1316 1292 1348
rect 1326 1316 1364 1348
rect 1398 1316 1436 1348
rect 1470 1316 1508 1348
rect 1542 1316 1580 1348
rect 1614 1316 1652 1350
rect 1686 1316 1720 1350
rect 1873 2206 2043 2241
rect 1907 2172 1941 2206
rect 1975 2172 2009 2206
rect 1873 2137 2043 2172
rect 1907 2103 1941 2137
rect 1975 2103 2009 2137
rect 1873 2068 2043 2103
rect 1907 2034 1941 2068
rect 1975 2034 2009 2068
rect 1873 1999 2043 2034
rect 1907 1965 1941 1999
rect 1975 1965 2009 1999
rect 1873 1930 2043 1965
rect 1907 1896 1941 1930
rect 1975 1896 2009 1930
rect 1873 1861 2043 1896
rect 1873 1860 1941 1861
rect 1907 1827 1941 1860
rect 1975 1827 2009 1861
rect 1907 1826 2043 1827
rect 1873 1792 2043 1826
rect 1873 1790 1941 1792
rect 1907 1758 1941 1790
rect 1975 1758 2009 1792
rect 1907 1756 2043 1758
rect 1873 1722 2043 1756
rect 1873 1720 1941 1722
rect 1907 1688 1941 1720
rect 1975 1688 2009 1722
rect 1907 1686 2043 1688
rect 1873 1652 2043 1686
rect 1873 1650 1941 1652
rect 1907 1618 1941 1650
rect 1975 1618 2009 1652
rect 1907 1616 2043 1618
rect 1873 1582 2043 1616
rect 1873 1580 1941 1582
rect 1907 1548 1941 1580
rect 1975 1548 2009 1582
rect 1907 1546 2043 1548
rect 1873 1512 2043 1546
rect 1873 1510 1941 1512
rect 1907 1478 1941 1510
rect 1975 1478 2009 1512
rect 1907 1476 2043 1478
rect 1873 1442 2043 1476
rect 1873 1440 1941 1442
rect 1907 1408 1941 1440
rect 1975 1408 2009 1442
rect 1907 1406 2043 1408
rect 1873 1372 2043 1406
rect 1873 1370 1941 1372
rect 1907 1338 1941 1370
rect 1975 1338 2009 1372
rect 1907 1336 2043 1338
rect 172 1266 206 1300
rect 240 1298 308 1300
rect 240 1266 274 1298
rect 138 1264 274 1266
rect 138 1231 308 1264
rect 172 1197 206 1231
rect 240 1229 308 1231
rect 240 1197 274 1229
rect 138 1195 274 1197
rect 138 1162 308 1195
rect 172 1128 206 1162
rect 240 1160 308 1162
rect 1873 1302 2043 1336
rect 1873 1300 1941 1302
rect 1907 1268 1941 1300
rect 1975 1268 2009 1302
rect 1907 1266 2043 1268
rect 1873 1232 2043 1266
rect 1873 1230 1941 1232
rect 1907 1198 1941 1230
rect 1975 1198 2009 1232
rect 1907 1196 2043 1198
rect 1873 1162 2043 1196
rect 1873 1160 1941 1162
rect 240 1128 274 1160
rect 138 1126 274 1128
rect 308 1126 344 1160
rect 378 1126 414 1160
rect 448 1126 484 1160
rect 518 1126 554 1160
rect 588 1126 624 1160
rect 658 1126 694 1160
rect 728 1126 764 1160
rect 798 1126 834 1160
rect 868 1126 904 1160
rect 938 1126 974 1160
rect 1008 1126 1044 1160
rect 1078 1126 1114 1160
rect 1148 1126 1183 1160
rect 1217 1126 1252 1160
rect 1286 1126 1321 1160
rect 1355 1126 1390 1160
rect 1424 1126 1459 1160
rect 1493 1126 1528 1160
rect 1562 1126 1597 1160
rect 1631 1126 1666 1160
rect 1700 1126 1735 1160
rect 1769 1126 1804 1160
rect 1838 1126 1873 1160
rect 1907 1128 1941 1160
rect 1975 1128 2009 1162
rect 1907 1126 2043 1128
rect 138 1093 2043 1126
rect 172 1092 2043 1093
rect 172 1059 206 1092
rect 138 1058 206 1059
rect 240 1058 276 1092
rect 310 1058 346 1092
rect 380 1058 416 1092
rect 450 1058 486 1092
rect 520 1058 556 1092
rect 590 1058 626 1092
rect 660 1058 696 1092
rect 730 1058 766 1092
rect 800 1058 836 1092
rect 870 1058 905 1092
rect 939 1058 974 1092
rect 1008 1058 1043 1092
rect 1077 1058 1112 1092
rect 1146 1058 1181 1092
rect 1215 1058 1250 1092
rect 1284 1058 1319 1092
rect 1353 1058 1388 1092
rect 1422 1058 1457 1092
rect 1491 1058 1526 1092
rect 1560 1058 1595 1092
rect 1629 1058 1664 1092
rect 1698 1058 1733 1092
rect 1767 1058 1802 1092
rect 1836 1058 1871 1092
rect 1905 1058 1941 1092
rect 1975 1058 2009 1092
rect 138 1024 2043 1058
rect 138 990 206 1024
rect 240 990 276 1024
rect 310 990 346 1024
rect 380 990 416 1024
rect 450 990 486 1024
rect 520 990 556 1024
rect 590 990 626 1024
rect 660 990 696 1024
rect 730 990 766 1024
rect 800 990 836 1024
rect 870 990 905 1024
rect 939 990 974 1024
rect 1008 990 1043 1024
rect 1077 990 1112 1024
rect 1146 990 1181 1024
rect 1215 990 1250 1024
rect 1284 990 1319 1024
rect 1353 990 1388 1024
rect 1422 990 1457 1024
rect 1491 990 1526 1024
rect 1560 990 1595 1024
rect 1629 990 1664 1024
rect 1698 990 1733 1024
rect 1767 990 1802 1024
rect 1836 990 1871 1024
rect 1905 990 1940 1024
rect 1974 990 2043 1024
<< viali >>
rect 2297 25509 2306 25533
rect 2306 25509 2331 25533
rect 2373 25509 2378 25533
rect 2378 25509 2407 25533
rect 2449 25509 2450 25533
rect 2450 25509 2483 25533
rect 2525 25509 2556 25533
rect 2556 25509 2559 25533
rect 2601 25509 2628 25533
rect 2628 25509 2635 25533
rect 2677 25509 2700 25533
rect 2700 25509 2711 25533
rect 2753 25509 2771 25533
rect 2771 25509 2787 25533
rect 2829 25509 2842 25533
rect 2842 25509 2863 25533
rect 2904 25509 2913 25533
rect 2913 25509 2938 25533
rect 2979 25509 2984 25533
rect 2984 25509 3013 25533
rect 3054 25509 3055 25533
rect 3055 25509 3088 25533
rect 2297 25499 2331 25509
rect 2373 25499 2407 25509
rect 2449 25499 2483 25509
rect 2525 25499 2559 25509
rect 2601 25499 2635 25509
rect 2677 25499 2711 25509
rect 2753 25499 2787 25509
rect 2829 25499 2863 25509
rect 2904 25499 2938 25509
rect 2979 25499 3013 25509
rect 3054 25499 3088 25509
rect 3129 25499 3163 25533
rect 703 25458 728 25492
rect 728 25458 737 25492
rect 775 25458 809 25492
rect 847 25458 881 25492
rect 919 25458 953 25492
rect 703 25385 728 25419
rect 728 25385 737 25419
rect 775 25385 809 25419
rect 847 25385 881 25419
rect 919 25385 953 25419
rect 703 25312 728 25346
rect 728 25312 737 25346
rect 775 25312 809 25346
rect 847 25312 881 25346
rect 919 25312 953 25346
rect 703 25239 728 25273
rect 728 25239 737 25273
rect 775 25239 809 25273
rect 847 25239 881 25273
rect 919 25239 953 25273
rect 703 25166 728 25200
rect 728 25166 737 25200
rect 775 25166 809 25200
rect 847 25166 881 25200
rect 919 25166 953 25200
rect 703 25093 728 25127
rect 728 25093 737 25127
rect 775 25093 809 25127
rect 847 25093 881 25127
rect 919 25093 953 25127
rect 703 25020 728 25054
rect 728 25020 737 25054
rect 775 25020 809 25054
rect 847 25020 881 25054
rect 919 25020 953 25054
rect 2297 25441 2306 25461
rect 2306 25441 2331 25461
rect 2373 25441 2378 25461
rect 2378 25441 2407 25461
rect 2449 25441 2450 25461
rect 2450 25441 2483 25461
rect 2525 25441 2556 25461
rect 2556 25441 2559 25461
rect 2601 25441 2628 25461
rect 2628 25441 2635 25461
rect 2677 25441 2700 25461
rect 2700 25441 2711 25461
rect 2753 25441 2771 25461
rect 2771 25441 2787 25461
rect 2829 25441 2842 25461
rect 2842 25441 2863 25461
rect 2904 25441 2913 25461
rect 2913 25441 2938 25461
rect 2979 25441 2984 25461
rect 2984 25441 3013 25461
rect 3054 25441 3055 25461
rect 3055 25441 3088 25461
rect 2297 25427 2331 25441
rect 2373 25427 2407 25441
rect 2449 25427 2483 25441
rect 2525 25427 2559 25441
rect 2601 25427 2635 25441
rect 2677 25427 2711 25441
rect 2753 25427 2787 25441
rect 2829 25427 2863 25441
rect 2904 25427 2938 25441
rect 2979 25427 3013 25441
rect 3054 25427 3088 25441
rect 3129 25427 3163 25461
rect 2297 25373 2306 25389
rect 2306 25373 2331 25389
rect 2373 25373 2378 25389
rect 2378 25373 2407 25389
rect 2449 25373 2450 25389
rect 2450 25373 2483 25389
rect 2525 25373 2556 25389
rect 2556 25373 2559 25389
rect 2601 25373 2628 25389
rect 2628 25373 2635 25389
rect 2677 25373 2700 25389
rect 2700 25373 2711 25389
rect 2753 25373 2771 25389
rect 2771 25373 2787 25389
rect 2829 25373 2842 25389
rect 2842 25373 2863 25389
rect 2904 25373 2913 25389
rect 2913 25373 2938 25389
rect 2979 25373 2984 25389
rect 2984 25373 3013 25389
rect 3054 25373 3055 25389
rect 3055 25373 3088 25389
rect 2297 25355 2331 25373
rect 2373 25355 2407 25373
rect 2449 25355 2483 25373
rect 2525 25355 2559 25373
rect 2601 25355 2635 25373
rect 2677 25355 2711 25373
rect 2753 25355 2787 25373
rect 2829 25355 2863 25373
rect 2904 25355 2938 25373
rect 2979 25355 3013 25373
rect 3054 25355 3088 25373
rect 3129 25355 3163 25389
rect 703 24968 737 24981
rect 775 24968 809 24981
rect 847 24968 881 24981
rect 919 24968 953 24981
rect 703 24947 728 24968
rect 728 24947 737 24968
rect 775 24947 796 24968
rect 796 24947 809 24968
rect 847 24947 864 24968
rect 864 24947 881 24968
rect 919 24947 932 24968
rect 932 24947 953 24968
rect 703 24899 737 24908
rect 775 24899 809 24908
rect 847 24899 881 24908
rect 919 24899 953 24908
rect 703 24874 728 24899
rect 728 24874 737 24899
rect 775 24874 796 24899
rect 796 24874 809 24899
rect 847 24874 864 24899
rect 864 24874 881 24899
rect 919 24874 932 24899
rect 932 24874 953 24899
rect 703 24830 737 24835
rect 775 24830 809 24835
rect 847 24830 881 24835
rect 919 24830 953 24835
rect 703 24801 728 24830
rect 728 24801 737 24830
rect 775 24801 796 24830
rect 796 24801 809 24830
rect 847 24801 864 24830
rect 864 24801 881 24830
rect 919 24801 932 24830
rect 932 24801 953 24830
rect 703 24761 737 24762
rect 775 24761 809 24762
rect 847 24761 881 24762
rect 919 24761 953 24762
rect 703 24728 728 24761
rect 728 24728 737 24761
rect 775 24728 796 24761
rect 796 24728 809 24761
rect 847 24728 864 24761
rect 864 24728 881 24761
rect 919 24728 932 24761
rect 932 24728 953 24761
rect 703 24658 728 24689
rect 728 24658 737 24689
rect 775 24658 796 24689
rect 796 24658 809 24689
rect 847 24658 864 24689
rect 864 24658 881 24689
rect 919 24658 932 24689
rect 932 24658 953 24689
rect 703 24655 737 24658
rect 775 24655 809 24658
rect 847 24655 881 24658
rect 919 24655 953 24658
rect 703 24589 728 24616
rect 728 24589 737 24616
rect 775 24589 796 24616
rect 796 24589 809 24616
rect 847 24589 864 24616
rect 864 24589 881 24616
rect 919 24589 932 24616
rect 932 24589 953 24616
rect 703 24582 737 24589
rect 775 24582 809 24589
rect 847 24582 881 24589
rect 919 24582 953 24589
rect 703 24520 728 24543
rect 728 24520 737 24543
rect 775 24520 796 24543
rect 796 24520 809 24543
rect 847 24520 864 24543
rect 864 24520 881 24543
rect 919 24520 932 24543
rect 932 24520 953 24543
rect 703 24509 737 24520
rect 775 24509 809 24520
rect 847 24509 881 24520
rect 919 24509 953 24520
rect 703 24451 728 24470
rect 728 24451 737 24470
rect 775 24451 796 24470
rect 796 24451 809 24470
rect 847 24451 864 24470
rect 864 24451 881 24470
rect 919 24451 932 24470
rect 932 24451 953 24470
rect 703 24436 737 24451
rect 775 24436 809 24451
rect 847 24436 881 24451
rect 919 24436 953 24451
rect 703 24382 728 24397
rect 728 24382 737 24397
rect 775 24382 796 24397
rect 796 24382 809 24397
rect 847 24382 864 24397
rect 864 24382 881 24397
rect 919 24382 932 24397
rect 932 24382 953 24397
rect 703 24363 737 24382
rect 775 24363 809 24382
rect 847 24363 881 24382
rect 919 24363 953 24382
rect 703 24313 728 24324
rect 728 24313 737 24324
rect 775 24313 796 24324
rect 796 24313 809 24324
rect 847 24313 864 24324
rect 864 24313 881 24324
rect 919 24313 932 24324
rect 932 24313 953 24324
rect 703 24290 737 24313
rect 775 24290 809 24313
rect 847 24290 881 24313
rect 919 24290 953 24313
rect 703 24244 728 24251
rect 728 24244 737 24251
rect 775 24244 796 24251
rect 796 24244 809 24251
rect 847 24244 864 24251
rect 864 24244 881 24251
rect 919 24244 932 24251
rect 932 24244 953 24251
rect 703 24217 737 24244
rect 775 24217 809 24244
rect 847 24217 881 24244
rect 919 24217 953 24244
rect 703 24175 728 24178
rect 728 24175 737 24178
rect 775 24175 796 24178
rect 796 24175 809 24178
rect 847 24175 864 24178
rect 864 24175 881 24178
rect 919 24175 932 24178
rect 932 24175 953 24178
rect 703 24144 737 24175
rect 775 24144 809 24175
rect 847 24144 881 24175
rect 919 24144 953 24175
rect 703 24071 737 24105
rect 775 24071 809 24105
rect 847 24071 881 24105
rect 919 24071 953 24105
rect 703 24002 737 24031
rect 775 24002 809 24031
rect 847 24002 881 24031
rect 919 24002 953 24031
rect 703 23997 728 24002
rect 728 23997 737 24002
rect 775 23997 796 24002
rect 796 23997 809 24002
rect 847 23997 864 24002
rect 864 23997 881 24002
rect 919 23997 932 24002
rect 932 23997 953 24002
rect 703 23933 737 23957
rect 775 23933 809 23957
rect 847 23933 881 23957
rect 919 23933 953 23957
rect 703 23923 728 23933
rect 728 23923 737 23933
rect 775 23923 796 23933
rect 796 23923 809 23933
rect 847 23923 864 23933
rect 864 23923 881 23933
rect 919 23923 932 23933
rect 932 23923 953 23933
rect 703 23864 737 23883
rect 775 23864 809 23883
rect 847 23864 881 23883
rect 919 23864 953 23883
rect 703 23849 728 23864
rect 728 23849 737 23864
rect 775 23849 796 23864
rect 796 23849 809 23864
rect 847 23849 864 23864
rect 864 23849 881 23864
rect 919 23849 932 23864
rect 932 23849 953 23864
rect 703 23795 737 23809
rect 775 23795 809 23809
rect 847 23795 881 23809
rect 919 23795 953 23809
rect 703 23775 728 23795
rect 728 23775 737 23795
rect 775 23775 796 23795
rect 796 23775 809 23795
rect 847 23775 864 23795
rect 864 23775 881 23795
rect 919 23775 932 23795
rect 932 23775 953 23795
rect 703 23726 737 23735
rect 775 23726 809 23735
rect 847 23726 881 23735
rect 919 23726 953 23735
rect 703 23701 728 23726
rect 728 23701 737 23726
rect 775 23701 796 23726
rect 796 23701 809 23726
rect 847 23701 864 23726
rect 864 23701 881 23726
rect 919 23701 932 23726
rect 932 23701 953 23726
rect 703 23657 737 23661
rect 775 23657 809 23661
rect 847 23657 881 23661
rect 919 23657 953 23661
rect 703 23627 728 23657
rect 728 23627 737 23657
rect 775 23627 796 23657
rect 796 23627 809 23657
rect 847 23627 864 23657
rect 864 23627 881 23657
rect 919 23627 932 23657
rect 932 23627 953 23657
rect 703 23554 728 23587
rect 728 23554 737 23587
rect 775 23554 796 23587
rect 796 23554 809 23587
rect 847 23554 864 23587
rect 864 23554 881 23587
rect 919 23554 932 23587
rect 932 23554 953 23587
rect 703 23553 737 23554
rect 775 23553 809 23554
rect 847 23553 881 23554
rect 919 23553 953 23554
rect 703 23485 728 23513
rect 728 23485 737 23513
rect 775 23485 796 23513
rect 796 23485 809 23513
rect 847 23485 864 23513
rect 864 23485 881 23513
rect 919 23485 932 23513
rect 932 23485 953 23513
rect 703 23479 737 23485
rect 775 23479 809 23485
rect 847 23479 881 23485
rect 919 23479 953 23485
rect 703 23416 728 23439
rect 728 23416 737 23439
rect 775 23416 796 23439
rect 796 23416 809 23439
rect 847 23416 864 23439
rect 864 23416 881 23439
rect 919 23416 932 23439
rect 932 23416 953 23439
rect 703 23405 737 23416
rect 775 23405 809 23416
rect 847 23405 881 23416
rect 919 23405 953 23416
rect 703 23347 728 23365
rect 728 23347 737 23365
rect 775 23347 796 23365
rect 796 23347 809 23365
rect 847 23347 864 23365
rect 864 23347 881 23365
rect 919 23347 932 23365
rect 932 23347 953 23365
rect 703 23331 737 23347
rect 775 23331 809 23347
rect 847 23331 881 23347
rect 919 23331 953 23347
rect 703 23278 728 23291
rect 728 23278 737 23291
rect 775 23278 796 23291
rect 796 23278 809 23291
rect 847 23278 864 23291
rect 864 23278 881 23291
rect 919 23278 932 23291
rect 932 23278 953 23291
rect 703 23257 737 23278
rect 775 23257 809 23278
rect 847 23257 881 23278
rect 919 23257 953 23278
rect 1200 25307 1234 25341
rect 1274 25313 1308 25347
rect 1352 25313 1386 25347
rect 1430 25313 1464 25347
rect 1508 25313 1542 25347
rect 1587 25313 1621 25347
rect 1666 25313 1700 25347
rect 1745 25313 1779 25347
rect 1824 25313 1858 25347
rect 1903 25313 1937 25347
rect 1982 25313 2016 25347
rect 1200 25233 1234 25267
rect 1200 25159 1234 25193
rect 1200 25085 1234 25119
rect 1200 25011 1234 25045
rect 1200 24937 1234 24971
rect 1200 24863 1234 24897
rect 1200 24790 1234 24824
rect 1200 24717 1234 24751
rect 1200 24644 1234 24678
rect 1200 24571 1234 24605
rect 1200 24498 1234 24532
rect 1200 24425 1234 24459
rect 1200 24352 1234 24386
rect 1200 24279 1234 24313
rect 1200 24206 1234 24240
rect 1200 24133 1234 24167
rect 1200 24060 1234 24094
rect 1200 23987 1234 24021
rect 1200 23914 1234 23948
rect 1200 23841 1234 23875
rect 1200 23768 1234 23802
rect 1200 23695 1234 23729
rect 1200 23622 1234 23656
rect 1200 23549 1234 23583
rect 1200 23476 1234 23510
rect 1200 23403 1234 23437
rect 1200 23330 1234 23364
rect 1200 23257 1234 23291
rect 1200 23184 1234 23218
rect 1200 23111 1234 23145
rect 2056 25307 2090 25341
rect 2056 25234 2090 25268
rect 2056 25161 2090 25195
rect 2056 25088 2090 25122
rect 2056 25015 2090 25049
rect 2056 24942 2090 24976
rect 2056 24869 2090 24903
rect 2056 24796 2090 24830
rect 2056 24723 2090 24757
rect 2297 25305 2306 25317
rect 2306 25305 2331 25317
rect 2373 25305 2378 25317
rect 2378 25305 2407 25317
rect 2449 25305 2450 25317
rect 2450 25305 2483 25317
rect 2525 25305 2556 25317
rect 2556 25305 2559 25317
rect 2601 25305 2628 25317
rect 2628 25305 2635 25317
rect 2677 25305 2700 25317
rect 2700 25305 2711 25317
rect 2753 25305 2771 25317
rect 2771 25305 2787 25317
rect 2829 25305 2842 25317
rect 2842 25305 2863 25317
rect 2904 25305 2913 25317
rect 2913 25305 2938 25317
rect 2979 25305 2984 25317
rect 2984 25305 3013 25317
rect 3054 25305 3055 25317
rect 3055 25305 3088 25317
rect 2297 25283 2331 25305
rect 2373 25283 2407 25305
rect 2449 25283 2483 25305
rect 2525 25283 2559 25305
rect 2601 25283 2635 25305
rect 2677 25283 2711 25305
rect 2753 25283 2787 25305
rect 2829 25283 2863 25305
rect 2904 25283 2938 25305
rect 2979 25283 3013 25305
rect 3054 25283 3088 25305
rect 3129 25283 3163 25317
rect 2297 25237 2306 25245
rect 2306 25237 2331 25245
rect 2373 25237 2378 25245
rect 2378 25237 2407 25245
rect 2449 25237 2450 25245
rect 2450 25237 2483 25245
rect 2525 25237 2556 25245
rect 2556 25237 2559 25245
rect 2601 25237 2628 25245
rect 2628 25237 2635 25245
rect 2677 25237 2700 25245
rect 2700 25237 2711 25245
rect 2753 25237 2771 25245
rect 2771 25237 2787 25245
rect 2829 25237 2842 25245
rect 2842 25237 2863 25245
rect 2904 25237 2913 25245
rect 2913 25237 2938 25245
rect 2979 25237 2984 25245
rect 2984 25237 3013 25245
rect 3054 25237 3055 25245
rect 3055 25237 3088 25245
rect 2297 25211 2331 25237
rect 2373 25211 2407 25237
rect 2449 25211 2483 25237
rect 2525 25211 2559 25237
rect 2601 25211 2635 25237
rect 2677 25211 2711 25237
rect 2753 25211 2787 25237
rect 2829 25211 2863 25237
rect 2904 25211 2938 25237
rect 2979 25211 3013 25237
rect 3054 25211 3088 25237
rect 3129 25211 3163 25245
rect 2297 25169 2306 25173
rect 2306 25169 2331 25173
rect 2373 25169 2378 25173
rect 2378 25169 2407 25173
rect 2449 25169 2450 25173
rect 2450 25169 2483 25173
rect 2525 25169 2556 25173
rect 2556 25169 2559 25173
rect 2601 25169 2628 25173
rect 2628 25169 2635 25173
rect 2677 25169 2700 25173
rect 2700 25169 2711 25173
rect 2753 25169 2771 25173
rect 2771 25169 2787 25173
rect 2829 25169 2842 25173
rect 2842 25169 2863 25173
rect 2904 25169 2913 25173
rect 2913 25169 2938 25173
rect 2979 25169 2984 25173
rect 2984 25169 3013 25173
rect 3054 25169 3055 25173
rect 3055 25169 3088 25173
rect 2297 25139 2331 25169
rect 2373 25139 2407 25169
rect 2449 25139 2483 25169
rect 2525 25139 2559 25169
rect 2601 25139 2635 25169
rect 2677 25139 2711 25169
rect 2753 25139 2787 25169
rect 2829 25139 2863 25169
rect 2904 25139 2938 25169
rect 2979 25139 3013 25169
rect 3054 25139 3088 25169
rect 3129 25139 3163 25173
rect 2297 25067 2331 25101
rect 2373 25067 2407 25101
rect 2449 25067 2483 25101
rect 2525 25067 2559 25101
rect 2601 25067 2635 25101
rect 2677 25067 2711 25101
rect 2753 25067 2787 25101
rect 2829 25067 2863 25101
rect 2904 25067 2938 25101
rect 2979 25067 3013 25101
rect 3054 25067 3088 25101
rect 3129 25067 3163 25101
rect 2297 24999 2331 25029
rect 2373 24999 2407 25029
rect 2449 24999 2483 25029
rect 2525 24999 2559 25029
rect 2601 24999 2635 25029
rect 2677 24999 2711 25029
rect 2753 24999 2787 25029
rect 2829 24999 2863 25029
rect 2904 24999 2938 25029
rect 2979 24999 3013 25029
rect 3054 24999 3088 25029
rect 2297 24995 2306 24999
rect 2306 24995 2331 24999
rect 2373 24995 2378 24999
rect 2378 24995 2407 24999
rect 2449 24995 2450 24999
rect 2450 24995 2483 24999
rect 2525 24995 2556 24999
rect 2556 24995 2559 24999
rect 2601 24995 2628 24999
rect 2628 24995 2635 24999
rect 2677 24995 2700 24999
rect 2700 24995 2711 24999
rect 2753 24995 2771 24999
rect 2771 24995 2787 24999
rect 2829 24995 2842 24999
rect 2842 24995 2863 24999
rect 2904 24995 2913 24999
rect 2913 24995 2938 24999
rect 2979 24995 2984 24999
rect 2984 24995 3013 24999
rect 3054 24995 3055 24999
rect 3055 24995 3088 24999
rect 3129 24995 3163 25029
rect 2297 24931 2331 24957
rect 2373 24931 2407 24957
rect 2449 24931 2483 24957
rect 2525 24931 2559 24957
rect 2601 24931 2635 24957
rect 2677 24931 2711 24957
rect 2753 24931 2787 24957
rect 2829 24931 2863 24957
rect 2904 24931 2938 24957
rect 2979 24931 3013 24957
rect 3054 24931 3088 24957
rect 2297 24923 2306 24931
rect 2306 24923 2331 24931
rect 2373 24923 2378 24931
rect 2378 24923 2407 24931
rect 2449 24923 2450 24931
rect 2450 24923 2483 24931
rect 2525 24923 2556 24931
rect 2556 24923 2559 24931
rect 2601 24923 2628 24931
rect 2628 24923 2635 24931
rect 2677 24923 2700 24931
rect 2700 24923 2711 24931
rect 2753 24923 2771 24931
rect 2771 24923 2787 24931
rect 2829 24923 2842 24931
rect 2842 24923 2863 24931
rect 2904 24923 2913 24931
rect 2913 24923 2938 24931
rect 2979 24923 2984 24931
rect 2984 24923 3013 24931
rect 3054 24923 3055 24931
rect 3055 24923 3088 24931
rect 3129 24923 3163 24957
rect 2297 24863 2331 24885
rect 2373 24863 2407 24885
rect 2449 24863 2483 24885
rect 2525 24863 2559 24885
rect 2601 24863 2635 24885
rect 2677 24863 2711 24885
rect 2753 24863 2787 24885
rect 2829 24863 2863 24885
rect 2904 24863 2938 24885
rect 2979 24863 3013 24885
rect 3054 24863 3088 24885
rect 2297 24851 2306 24863
rect 2306 24851 2331 24863
rect 2373 24851 2378 24863
rect 2378 24851 2407 24863
rect 2449 24851 2450 24863
rect 2450 24851 2483 24863
rect 2525 24851 2556 24863
rect 2556 24851 2559 24863
rect 2601 24851 2628 24863
rect 2628 24851 2635 24863
rect 2677 24851 2700 24863
rect 2700 24851 2711 24863
rect 2753 24851 2771 24863
rect 2771 24851 2787 24863
rect 2829 24851 2842 24863
rect 2842 24851 2863 24863
rect 2904 24851 2913 24863
rect 2913 24851 2938 24863
rect 2979 24851 2984 24863
rect 2984 24851 3013 24863
rect 3054 24851 3055 24863
rect 3055 24851 3088 24863
rect 3129 24851 3163 24885
rect 2297 24795 2331 24813
rect 2373 24795 2407 24813
rect 2449 24795 2483 24813
rect 2525 24795 2559 24813
rect 2601 24795 2635 24813
rect 2677 24795 2711 24813
rect 2753 24795 2787 24813
rect 2829 24795 2863 24813
rect 2904 24795 2938 24813
rect 2979 24795 3013 24813
rect 3054 24795 3088 24813
rect 2297 24779 2306 24795
rect 2306 24779 2331 24795
rect 2373 24779 2378 24795
rect 2378 24779 2407 24795
rect 2449 24779 2450 24795
rect 2450 24779 2483 24795
rect 2525 24779 2556 24795
rect 2556 24779 2559 24795
rect 2601 24779 2628 24795
rect 2628 24779 2635 24795
rect 2677 24779 2700 24795
rect 2700 24779 2711 24795
rect 2753 24779 2771 24795
rect 2771 24779 2787 24795
rect 2829 24779 2842 24795
rect 2842 24779 2863 24795
rect 2904 24779 2913 24795
rect 2913 24779 2938 24795
rect 2979 24779 2984 24795
rect 2984 24779 3013 24795
rect 3054 24779 3055 24795
rect 3055 24779 3088 24795
rect 3129 24779 3163 24813
rect 2056 24650 2090 24684
rect 2056 24578 2090 24612
rect 2056 24506 2090 24540
rect 2130 24522 2164 24556
rect 2207 24522 2241 24556
rect 2284 24522 2318 24556
rect 2361 24522 2395 24556
rect 2438 24522 2472 24556
rect 2515 24522 2549 24556
rect 2592 24522 2626 24556
rect 2669 24522 2703 24556
rect 2746 24522 2780 24556
rect 2823 24522 2857 24556
rect 2900 24522 2934 24556
rect 2056 24434 2090 24468
rect 2056 24362 2090 24396
rect 2056 24290 2090 24324
rect 2056 24218 2090 24252
rect 2056 24146 2090 24180
rect 2056 24074 2090 24108
rect 2056 24002 2090 24036
rect 2056 23930 2090 23964
rect 2056 23858 2090 23892
rect 2056 23786 2090 23820
rect 2056 23714 2090 23748
rect 2056 23642 2090 23676
rect 2056 23570 2090 23604
rect 2056 23498 2090 23532
rect 2056 23426 2090 23460
rect 2056 23354 2090 23388
rect 2056 23282 2090 23316
rect 2056 23210 2090 23244
rect 2056 23138 2090 23172
rect 822 23039 856 23073
rect 894 23039 928 23073
rect 966 23039 1000 23073
rect 1038 23039 1072 23073
rect 1110 23039 1144 23073
rect 1182 23039 1216 23073
rect 1254 23039 1288 23073
rect 1326 23039 1360 23073
rect 1398 23039 1432 23073
rect 1471 23039 1505 23073
rect 1544 23039 1578 23073
rect 1617 23039 1651 23073
rect 1690 23039 1724 23073
rect 1763 23039 1797 23073
rect 1836 23039 1870 23073
rect 1909 23039 1943 23073
rect 1982 23039 2016 23073
rect 2056 23066 2090 23100
rect 816 22967 850 23001
rect 2056 22995 2090 23028
rect 2056 22994 2090 22995
rect 1000 22914 1034 22948
rect 1077 22914 1111 22948
rect 1154 22914 1188 22948
rect 1231 22914 1265 22948
rect 1308 22914 1342 22948
rect 1384 22914 1418 22948
rect 1460 22914 1494 22948
rect 1536 22914 1570 22948
rect 1612 22914 1646 22948
rect 1688 22914 1722 22948
rect 1764 22914 1798 22948
rect 1840 22914 1874 22948
rect 1916 22914 1950 22948
rect 999 22758 1033 22792
rect 1076 22758 1110 22792
rect 1153 22758 1187 22792
rect 1230 22758 1264 22792
rect 1307 22758 1341 22792
rect 1384 22758 1418 22792
rect 1460 22758 1494 22792
rect 1536 22758 1570 22792
rect 1612 22758 1646 22792
rect 1688 22758 1722 22792
rect 1764 22758 1798 22792
rect 1840 22758 1874 22792
rect 1916 22758 1950 22792
rect 909 22697 943 22698
rect 909 22664 922 22697
rect 922 22664 943 22697
rect 2056 22744 2090 22762
rect 2056 22728 2090 22744
rect 2056 22672 2090 22687
rect 2056 22653 2090 22672
rect 909 22592 943 22626
rect 1000 22602 1034 22636
rect 1077 22602 1111 22636
rect 1154 22602 1188 22636
rect 1231 22602 1265 22636
rect 1308 22602 1342 22636
rect 1384 22602 1418 22636
rect 1460 22602 1494 22636
rect 1536 22602 1570 22636
rect 1612 22602 1646 22636
rect 1688 22602 1722 22636
rect 1764 22602 1798 22636
rect 1840 22602 1874 22636
rect 1916 22602 1950 22636
rect 2056 22600 2090 22612
rect 2056 22578 2090 22600
rect 816 22518 850 22552
rect 2056 22528 2090 22536
rect 816 22442 850 22476
rect 816 22366 850 22400
rect 912 22465 922 22498
rect 922 22465 946 22498
rect 912 22464 946 22465
rect 999 22492 1033 22526
rect 1076 22492 1110 22526
rect 1153 22492 1187 22526
rect 1230 22492 1264 22526
rect 1307 22492 1341 22526
rect 1384 22492 1418 22526
rect 1460 22492 1494 22526
rect 1536 22492 1570 22526
rect 1612 22492 1646 22526
rect 1688 22492 1722 22526
rect 1764 22492 1798 22526
rect 1840 22492 1874 22526
rect 1916 22492 1950 22526
rect 2056 22502 2090 22528
rect 912 22397 922 22426
rect 922 22397 946 22426
rect 912 22392 946 22397
rect 2056 22456 2090 22460
rect 2056 22426 2090 22456
rect 999 22336 1033 22370
rect 1076 22336 1110 22370
rect 1153 22336 1187 22370
rect 1230 22336 1264 22370
rect 1307 22336 1341 22370
rect 1384 22336 1418 22370
rect 1460 22336 1494 22370
rect 1536 22336 1570 22370
rect 1612 22336 1646 22370
rect 1688 22336 1722 22370
rect 1764 22336 1798 22370
rect 1840 22336 1874 22370
rect 1916 22336 1950 22370
rect 2056 22350 2090 22384
rect 816 22290 850 22324
rect 816 22214 850 22248
rect 816 22138 850 22172
rect 816 22062 850 22096
rect 816 21986 850 22020
rect 816 21909 850 21943
rect 816 21832 850 21866
rect 816 21755 850 21789
rect 816 21678 850 21712
rect 816 21601 850 21635
rect 816 21524 850 21558
rect 816 21447 850 21481
rect 2056 22278 2090 22308
rect 2056 22274 2090 22278
rect 2056 22198 2090 22232
rect 2056 22122 2090 22156
rect 2056 22046 2090 22080
rect 2056 21970 2090 22004
rect 2056 21894 2090 21928
rect 2056 21818 2090 21852
rect 2912 24427 2946 24461
rect 2912 24354 2946 24388
rect 2912 24281 2946 24315
rect 2912 24208 2946 24242
rect 2912 24135 2946 24169
rect 2912 24062 2946 24096
rect 2912 23989 2946 24023
rect 2912 23916 2946 23950
rect 2912 23843 2946 23877
rect 2912 23770 2946 23804
rect 2912 23697 2946 23731
rect 2912 23624 2946 23658
rect 2912 23551 2946 23585
rect 2912 23478 2946 23512
rect 2912 23405 2946 23439
rect 2912 23331 2946 23365
rect 2912 23257 2946 23291
rect 2912 23183 2946 23217
rect 2912 23109 2946 23143
rect 2912 23035 2946 23069
rect 2912 22961 2946 22995
rect 2912 22887 2946 22921
rect 2912 22813 2946 22847
rect 2912 22739 2946 22773
rect 2912 22665 2946 22699
rect 2912 22591 2946 22625
rect 2912 22517 2946 22551
rect 2912 22443 2946 22477
rect 2912 22369 2946 22403
rect 2912 22295 2946 22329
rect 2912 22221 2946 22255
rect 2912 22147 2946 22181
rect 2912 22073 2946 22107
rect 2912 21999 2946 22033
rect 2912 21925 2946 21959
rect 2912 21851 2946 21885
rect 2056 21742 2090 21776
rect 2056 21666 2090 21700
rect 2056 21590 2090 21624
rect 2912 21685 2946 21719
rect 2912 21611 2946 21645
rect 2056 21514 2090 21548
rect 2056 21438 2090 21472
rect 816 21370 850 21404
rect 890 21364 924 21398
rect 962 21364 996 21398
rect 1034 21364 1068 21398
rect 1106 21364 1140 21398
rect 1178 21364 1212 21398
rect 1250 21364 1284 21398
rect 1322 21364 1356 21398
rect 1394 21364 1428 21398
rect 1466 21364 1500 21398
rect 1538 21364 1572 21398
rect 1610 21364 1644 21398
rect 1682 21364 1716 21398
rect 1754 21364 1788 21398
rect 1826 21364 1860 21398
rect 1898 21364 1932 21398
rect 1970 21364 2004 21398
rect 2042 21364 2076 21398
rect 2115 21364 2149 21398
rect 2188 21364 2222 21398
rect 2261 21364 2295 21398
rect 265 18038 515 18144
rect 266 16588 300 16622
rect 341 16588 375 16622
rect 417 16588 451 16622
rect 493 16588 527 16622
rect 569 16588 603 16622
rect 266 16536 300 16550
rect 341 16536 375 16550
rect 417 16536 451 16550
rect 493 16536 527 16550
rect 569 16536 603 16550
rect 266 16516 281 16536
rect 281 16516 300 16536
rect 341 16516 349 16536
rect 349 16516 375 16536
rect 417 16516 451 16536
rect 493 16516 519 16536
rect 519 16516 527 16536
rect 569 16516 587 16536
rect 587 16516 603 16536
rect 2231 16137 2265 16171
rect 2304 16137 2338 16171
rect 2377 16137 2411 16171
rect 2450 16137 2484 16171
rect 2523 16137 2557 16171
rect 2596 16137 2630 16171
rect 2669 16137 2703 16171
rect 2742 16137 2776 16171
rect 2815 16137 2849 16171
rect 2888 16137 2922 16171
rect 2961 16137 2995 16171
rect 3034 16137 3068 16171
rect 3107 16137 3141 16171
rect 3180 16137 3214 16171
rect 3253 16137 3287 16171
rect 3326 16137 3360 16171
rect 3399 16137 3433 16171
rect 3472 16137 3506 16171
rect 3545 16137 3579 16171
rect 3618 16137 3652 16171
rect 3691 16137 3725 16171
rect 3764 16137 3798 16171
rect 3837 16137 3871 16171
rect 3910 16137 3944 16171
rect 3983 16137 4017 16171
rect 4056 16137 4090 16171
rect 4129 16137 4163 16171
rect 4202 16137 4236 16171
rect 4275 16137 4309 16171
rect 4348 16137 4382 16171
rect 4421 16137 4455 16171
rect 4494 16137 4528 16171
rect 4567 16137 4601 16171
rect 4640 16137 4674 16171
rect 4713 16137 4747 16171
rect 4786 16137 4820 16171
rect 4859 16137 4893 16171
rect 4932 16137 4966 16171
rect 5005 16137 5039 16171
rect 5078 16137 5112 16171
rect 5151 16137 5185 16171
rect 5224 16137 5258 16171
rect 5297 16137 5331 16171
rect 5370 16137 5404 16171
rect 5443 16137 5477 16171
rect 5516 16137 5550 16171
rect 5589 16137 5623 16171
rect 5662 16137 5696 16171
rect 5735 16137 5769 16171
rect 5808 16137 5842 16171
rect 5881 16137 5915 16171
rect 5954 16137 5988 16171
rect 6027 16137 6061 16171
rect 6100 16137 6134 16171
rect 6173 16137 6207 16171
rect 6246 16137 6280 16171
rect 6319 16137 6353 16171
rect 6392 16137 6426 16171
rect 6465 16137 6499 16171
rect 6538 16137 6572 16171
rect 6611 16137 6645 16171
rect 6684 16137 6718 16171
rect 6757 16137 6791 16171
rect 6830 16137 6864 16171
rect 6903 16137 6937 16171
rect 2231 16065 2265 16099
rect 2304 16065 2338 16099
rect 2377 16065 2411 16099
rect 2450 16065 2484 16099
rect 2523 16065 2557 16099
rect 2596 16065 2630 16099
rect 2669 16065 2703 16099
rect 2742 16065 2776 16099
rect 2815 16065 2849 16099
rect 2888 16065 2922 16099
rect 2961 16065 2995 16099
rect 3034 16065 3068 16099
rect 3107 16065 3141 16099
rect 3180 16065 3214 16099
rect 3253 16065 3287 16099
rect 3326 16065 3360 16099
rect 3399 16065 3433 16099
rect 3472 16065 3506 16099
rect 3545 16065 3579 16099
rect 3618 16065 3652 16099
rect 3691 16065 3725 16099
rect 3764 16065 3798 16099
rect 3837 16065 3871 16099
rect 3910 16065 3944 16099
rect 3983 16065 4017 16099
rect 4056 16065 4090 16099
rect 4129 16065 4163 16099
rect 4202 16065 4236 16099
rect 4275 16065 4309 16099
rect 4348 16065 4382 16099
rect 4421 16065 4455 16099
rect 4494 16065 4528 16099
rect 4567 16065 4601 16099
rect 4640 16065 4674 16099
rect 4713 16065 4747 16099
rect 4786 16065 4820 16099
rect 4859 16065 4893 16099
rect 4932 16065 4966 16099
rect 5005 16065 5039 16099
rect 5078 16065 5112 16099
rect 5151 16065 5185 16099
rect 5224 16065 5258 16099
rect 5297 16065 5331 16099
rect 5370 16065 5404 16099
rect 5443 16065 5477 16099
rect 5516 16065 5550 16099
rect 5589 16065 5623 16099
rect 5662 16065 5696 16099
rect 5735 16065 5769 16099
rect 5808 16065 5842 16099
rect 5881 16065 5915 16099
rect 5954 16065 5988 16099
rect 6027 16065 6061 16099
rect 6100 16065 6134 16099
rect 6173 16065 6207 16099
rect 6246 16065 6280 16099
rect 6319 16065 6353 16099
rect 6392 16065 6426 16099
rect 6465 16065 6499 16099
rect 6538 16065 6572 16099
rect 6611 16065 6645 16099
rect 6684 16065 6718 16099
rect 6757 16065 6791 16099
rect 6830 16065 6864 16099
rect 6903 16065 6937 16099
rect 2231 15993 2265 16027
rect 2304 15993 2338 16027
rect 2377 15993 2411 16027
rect 2450 15993 2484 16027
rect 2523 15993 2557 16027
rect 2596 15993 2630 16027
rect 2669 15993 2703 16027
rect 2742 15993 2776 16027
rect 2815 15993 2849 16027
rect 2888 15993 2922 16027
rect 2961 15993 2995 16027
rect 3034 15993 3068 16027
rect 3107 15993 3141 16027
rect 3180 15993 3214 16027
rect 3253 15993 3287 16027
rect 3326 15993 3360 16027
rect 3399 15993 3433 16027
rect 3472 15993 3506 16027
rect 3545 15993 3579 16027
rect 3618 15993 3652 16027
rect 3691 15993 3725 16027
rect 3764 15993 3798 16027
rect 3837 15993 3871 16027
rect 3910 15993 3944 16027
rect 3983 15993 4017 16027
rect 4056 15993 4090 16027
rect 4129 15993 4163 16027
rect 4202 15993 4236 16027
rect 4275 15993 4309 16027
rect 4348 15993 4382 16027
rect 4421 15993 4455 16027
rect 4494 15993 4528 16027
rect 4567 15993 4601 16027
rect 4640 15993 4674 16027
rect 4713 15993 4747 16027
rect 4786 15993 4820 16027
rect 4859 15993 4893 16027
rect 4932 15993 4966 16027
rect 5005 15993 5039 16027
rect 5078 15993 5112 16027
rect 5151 15993 5185 16027
rect 5224 15993 5258 16027
rect 5297 15993 5331 16027
rect 5370 15993 5404 16027
rect 5443 15993 5477 16027
rect 5516 15993 5550 16027
rect 5589 15993 5623 16027
rect 5662 15993 5696 16027
rect 5735 15993 5769 16027
rect 5808 15993 5842 16027
rect 5881 15993 5915 16027
rect 5954 15993 5988 16027
rect 6027 15993 6061 16027
rect 6100 15993 6134 16027
rect 6173 15993 6207 16027
rect 6246 15993 6280 16027
rect 6319 15993 6353 16027
rect 6392 15993 6426 16027
rect 6465 15993 6499 16027
rect 6538 15993 6572 16027
rect 6611 15993 6645 16027
rect 6684 15993 6718 16027
rect 6757 15993 6791 16027
rect 6830 15993 6864 16027
rect 6903 15993 6937 16027
rect 2231 15921 2265 15955
rect 2304 15921 2338 15955
rect 2377 15921 2411 15955
rect 2450 15921 2484 15955
rect 2523 15921 2557 15955
rect 2596 15921 2630 15955
rect 2669 15921 2703 15955
rect 2742 15921 2776 15955
rect 2815 15921 2849 15955
rect 2888 15921 2922 15955
rect 2961 15921 2995 15955
rect 3034 15921 3068 15955
rect 3107 15921 3141 15955
rect 3180 15921 3214 15955
rect 3253 15921 3287 15955
rect 3326 15921 3360 15955
rect 3399 15921 3433 15955
rect 3472 15921 3506 15955
rect 3545 15921 3579 15955
rect 3618 15921 3652 15955
rect 3691 15921 3725 15955
rect 3764 15921 3798 15955
rect 3837 15921 3871 15955
rect 3910 15921 3944 15955
rect 3983 15921 4017 15955
rect 4056 15921 4090 15955
rect 4129 15921 4163 15955
rect 4202 15921 4236 15955
rect 4275 15921 4309 15955
rect 4348 15921 4382 15955
rect 4421 15921 4455 15955
rect 4494 15921 4528 15955
rect 4567 15921 4601 15955
rect 4640 15921 4674 15955
rect 4713 15921 4747 15955
rect 4786 15921 4820 15955
rect 4859 15921 4893 15955
rect 4932 15921 4966 15955
rect 5005 15921 5039 15955
rect 5078 15921 5112 15955
rect 5151 15921 5185 15955
rect 5224 15921 5258 15955
rect 5297 15921 5331 15955
rect 5370 15921 5404 15955
rect 5443 15921 5477 15955
rect 5516 15921 5550 15955
rect 5589 15921 5623 15955
rect 5662 15921 5696 15955
rect 5735 15921 5769 15955
rect 5808 15921 5842 15955
rect 5881 15921 5915 15955
rect 5954 15921 5988 15955
rect 6027 15921 6061 15955
rect 6100 15921 6134 15955
rect 6173 15921 6207 15955
rect 6246 15921 6280 15955
rect 6319 15921 6353 15955
rect 6392 15921 6426 15955
rect 6465 15921 6499 15955
rect 6538 15921 6572 15955
rect 6611 15921 6645 15955
rect 6684 15921 6718 15955
rect 6757 15921 6791 15955
rect 6830 15921 6864 15955
rect 6903 15921 6937 15955
rect 6976 15921 17004 16171
rect 17004 15921 17018 16171
rect 1582 2854 1616 2888
rect 1654 2854 1688 2888
rect 1582 2779 1616 2813
rect 1654 2781 1688 2815
rect 1582 2704 1616 2738
rect 1654 2708 1688 2742
rect 1582 2629 1616 2663
rect 1654 2635 1688 2669
rect 1582 2554 1616 2588
rect 1654 2562 1688 2596
rect 1582 2479 1616 2513
rect 1654 2489 1688 2523
rect 1582 2404 1616 2438
rect 1654 2416 1688 2450
rect 1582 2329 1616 2363
rect 1654 2343 1688 2377
rect 1582 2254 1616 2288
rect 1654 2270 1688 2304
rect 1582 2188 1616 2213
rect 1654 2197 1688 2231
rect 686 2142 720 2176
rect 786 2146 820 2180
rect 861 2146 895 2180
rect 936 2146 970 2180
rect 1010 2146 1044 2180
rect 1084 2146 1118 2180
rect 1158 2146 1192 2180
rect 1232 2146 1266 2180
rect 1306 2146 1340 2180
rect 1582 2179 1584 2188
rect 1584 2179 1616 2188
rect 1654 2154 1686 2158
rect 1686 2154 1688 2158
rect 686 2092 720 2104
rect 686 2070 688 2092
rect 688 2070 720 2092
rect 1582 2117 1616 2138
rect 1654 2124 1688 2154
rect 1582 2104 1584 2117
rect 1584 2104 1616 2117
rect 1654 2081 1686 2085
rect 1686 2081 1688 2085
rect 1582 2046 1616 2062
rect 1654 2051 1688 2081
rect 1582 2028 1584 2046
rect 1584 2028 1616 2046
rect 779 1990 813 2024
rect 855 1990 889 2024
rect 931 1990 965 2024
rect 1007 1990 1041 2024
rect 1083 1990 1117 2024
rect 1159 1990 1193 2024
rect 1234 1990 1268 2024
rect 1654 2008 1686 2012
rect 1686 2008 1688 2012
rect 1582 1976 1616 1986
rect 1654 1978 1688 2008
rect 1582 1952 1584 1976
rect 1584 1952 1616 1976
rect 1654 1935 1686 1938
rect 1686 1935 1688 1938
rect 1582 1906 1616 1910
rect 1582 1876 1584 1906
rect 1584 1876 1616 1906
rect 1654 1904 1688 1935
rect 780 1834 814 1868
rect 856 1834 890 1868
rect 931 1834 965 1868
rect 1006 1834 1040 1868
rect 1081 1834 1115 1868
rect 1156 1834 1190 1868
rect 1231 1834 1265 1868
rect 1306 1834 1340 1868
rect 1654 1862 1686 1864
rect 1686 1862 1688 1864
rect 1582 1802 1584 1834
rect 1584 1802 1616 1834
rect 1654 1830 1688 1862
rect 1582 1800 1616 1802
rect 1654 1789 1686 1790
rect 1686 1789 1688 1790
rect 786 1724 820 1758
rect 861 1724 895 1758
rect 936 1724 970 1758
rect 1010 1724 1044 1758
rect 1084 1724 1118 1758
rect 1158 1724 1192 1758
rect 1232 1724 1266 1758
rect 1306 1724 1340 1758
rect 1582 1732 1584 1758
rect 1584 1732 1616 1758
rect 1654 1756 1688 1789
rect 1582 1724 1616 1732
rect 1582 1662 1584 1682
rect 1584 1662 1616 1682
rect 1654 1682 1688 1716
rect 1582 1648 1616 1662
rect 786 1568 820 1602
rect 861 1568 895 1602
rect 936 1568 970 1602
rect 1010 1568 1044 1602
rect 1084 1568 1118 1602
rect 1158 1568 1192 1602
rect 1232 1568 1266 1602
rect 1306 1568 1340 1602
rect 1582 1592 1584 1606
rect 1584 1592 1616 1606
rect 1654 1608 1688 1642
rect 1582 1572 1616 1592
rect 502 1497 504 1511
rect 504 1497 536 1511
rect 502 1477 536 1497
rect 1582 1522 1584 1530
rect 1584 1522 1616 1530
rect 1654 1534 1688 1568
rect 1582 1496 1616 1522
rect 574 1452 606 1454
rect 606 1452 608 1454
rect 646 1452 678 1454
rect 678 1452 680 1454
rect 718 1452 750 1454
rect 750 1452 752 1454
rect 790 1452 822 1454
rect 822 1452 824 1454
rect 862 1452 894 1454
rect 894 1452 896 1454
rect 934 1452 966 1454
rect 966 1452 968 1454
rect 1006 1452 1039 1454
rect 1039 1452 1040 1454
rect 574 1420 608 1452
rect 646 1420 680 1452
rect 718 1420 752 1452
rect 790 1420 824 1452
rect 862 1420 896 1452
rect 934 1420 968 1452
rect 1006 1420 1040 1452
rect 1078 1420 1112 1454
rect 1150 1420 1184 1454
rect 1222 1420 1256 1454
rect 1294 1420 1328 1454
rect 1366 1420 1400 1454
rect 1654 1460 1688 1494
rect 1438 1420 1472 1454
rect 1510 1452 1511 1454
rect 1511 1452 1544 1454
rect 1582 1452 1584 1454
rect 1584 1452 1616 1454
rect 1510 1420 1544 1452
rect 1582 1420 1616 1452
rect 1654 1386 1688 1420
rect 540 1348 574 1382
rect 617 1350 651 1382
rect 694 1350 728 1382
rect 771 1350 805 1382
rect 848 1350 882 1382
rect 925 1350 959 1382
rect 1002 1350 1036 1382
rect 1079 1350 1113 1382
rect 1156 1350 1190 1382
rect 1232 1350 1266 1382
rect 1308 1350 1342 1382
rect 1384 1350 1418 1382
rect 1460 1350 1494 1382
rect 1536 1350 1570 1382
rect 617 1348 649 1350
rect 649 1348 651 1350
rect 694 1348 720 1350
rect 720 1348 728 1350
rect 771 1348 791 1350
rect 791 1348 805 1350
rect 848 1348 862 1350
rect 862 1348 882 1350
rect 925 1348 933 1350
rect 933 1348 959 1350
rect 1002 1348 1004 1350
rect 1004 1348 1036 1350
rect 1079 1348 1110 1350
rect 1110 1348 1113 1350
rect 1156 1348 1182 1350
rect 1182 1348 1190 1350
rect 1232 1348 1254 1350
rect 1254 1348 1266 1350
rect 1308 1348 1326 1350
rect 1326 1348 1342 1350
rect 1384 1348 1398 1350
rect 1398 1348 1418 1350
rect 1460 1348 1470 1350
rect 1470 1348 1494 1350
rect 1536 1348 1542 1350
rect 1542 1348 1570 1350
<< metal1 >>
rect 520 25492 984 25686
rect 520 25458 703 25492
rect 737 25458 775 25492
rect 809 25458 847 25492
rect 881 25458 919 25492
rect 953 25458 984 25492
rect 520 25419 984 25458
rect 520 25385 703 25419
rect 737 25385 775 25419
rect 809 25385 847 25419
rect 881 25385 919 25419
rect 953 25385 984 25419
rect 520 25346 984 25385
rect 520 25312 703 25346
rect 737 25312 775 25346
rect 809 25312 847 25346
rect 881 25312 919 25346
rect 953 25312 984 25346
rect 520 25273 984 25312
rect 520 25239 703 25273
rect 737 25239 775 25273
rect 809 25239 847 25273
rect 881 25239 919 25273
rect 953 25239 984 25273
rect 520 25200 984 25239
rect 520 25166 703 25200
rect 737 25166 775 25200
rect 809 25166 847 25200
rect 881 25166 919 25200
rect 953 25166 984 25200
rect 520 25127 984 25166
rect 520 25093 703 25127
rect 737 25093 775 25127
rect 809 25093 847 25127
rect 881 25093 919 25127
rect 953 25093 984 25127
rect 520 25054 984 25093
rect 520 25020 703 25054
rect 737 25020 775 25054
rect 809 25020 847 25054
rect 881 25020 919 25054
rect 953 25020 984 25054
rect 520 24981 984 25020
rect 520 24947 703 24981
rect 737 24947 775 24981
rect 809 24947 847 24981
rect 881 24947 919 24981
rect 953 24947 984 24981
rect 520 24908 984 24947
rect 520 24874 703 24908
rect 737 24874 775 24908
rect 809 24874 847 24908
rect 881 24874 919 24908
rect 953 24874 984 24908
rect 520 24835 984 24874
rect 520 24801 703 24835
rect 737 24801 775 24835
rect 809 24801 847 24835
rect 881 24801 919 24835
rect 953 24801 984 24835
rect 520 24762 984 24801
rect 520 24728 703 24762
rect 737 24728 775 24762
rect 809 24728 847 24762
rect 881 24728 919 24762
rect 953 24728 984 24762
rect 520 24689 984 24728
rect 520 24655 703 24689
rect 737 24655 775 24689
rect 809 24655 847 24689
rect 881 24655 919 24689
rect 953 24655 984 24689
rect 520 24616 984 24655
rect 520 24582 703 24616
rect 737 24582 775 24616
rect 809 24582 847 24616
rect 881 24582 919 24616
rect 953 24582 984 24616
rect 520 24543 984 24582
rect 520 24509 703 24543
rect 737 24509 775 24543
rect 809 24509 847 24543
rect 881 24509 919 24543
rect 953 24509 984 24543
rect 520 24470 984 24509
rect 520 24436 703 24470
rect 737 24436 775 24470
rect 809 24436 847 24470
rect 881 24436 919 24470
rect 953 24436 984 24470
rect 520 24397 984 24436
rect 520 24363 703 24397
rect 737 24363 775 24397
rect 809 24363 847 24397
rect 881 24363 919 24397
rect 953 24363 984 24397
rect 520 24324 984 24363
rect 520 24290 703 24324
rect 737 24290 775 24324
rect 809 24290 847 24324
rect 881 24290 919 24324
rect 953 24290 984 24324
rect 520 24251 984 24290
rect 520 24217 703 24251
rect 737 24217 775 24251
rect 809 24217 847 24251
rect 881 24217 919 24251
rect 953 24217 984 24251
rect 520 24178 984 24217
rect 520 24144 703 24178
rect 737 24144 775 24178
rect 809 24144 847 24178
rect 881 24144 919 24178
rect 953 24144 984 24178
rect 520 24105 984 24144
rect 520 24071 703 24105
rect 737 24071 775 24105
rect 809 24071 847 24105
rect 881 24071 919 24105
rect 953 24071 984 24105
rect 520 24031 984 24071
rect 520 23997 703 24031
rect 737 23997 775 24031
rect 809 23997 847 24031
rect 881 23997 919 24031
rect 953 23997 984 24031
rect 520 23957 984 23997
rect 520 23923 703 23957
rect 737 23923 775 23957
rect 809 23923 847 23957
rect 881 23923 919 23957
rect 953 23923 984 23957
rect 520 23883 984 23923
rect 520 23849 703 23883
rect 737 23849 775 23883
rect 809 23849 847 23883
rect 881 23849 919 23883
rect 953 23849 984 23883
rect 520 23809 984 23849
rect 520 23775 703 23809
rect 737 23775 775 23809
rect 809 23775 847 23809
rect 881 23775 919 23809
rect 953 23775 984 23809
rect 520 23735 984 23775
rect 520 23701 703 23735
rect 737 23701 775 23735
rect 809 23701 847 23735
rect 881 23701 919 23735
rect 953 23701 984 23735
rect 520 23661 984 23701
rect 520 23627 703 23661
rect 737 23627 775 23661
rect 809 23627 847 23661
rect 881 23627 919 23661
rect 953 23627 984 23661
rect 520 23587 984 23627
rect 520 23553 703 23587
rect 737 23553 775 23587
rect 809 23553 847 23587
rect 881 23553 919 23587
rect 953 23553 984 23587
rect 520 23513 984 23553
rect 520 23479 703 23513
rect 737 23479 775 23513
rect 809 23479 847 23513
rect 881 23479 919 23513
rect 953 23479 984 23513
rect 520 23439 984 23479
rect 520 23405 703 23439
rect 737 23405 775 23439
rect 809 23405 847 23439
rect 881 23405 919 23439
rect 953 23405 984 23439
rect 520 23365 984 23405
rect 520 23331 703 23365
rect 737 23331 775 23365
rect 809 23331 847 23365
rect 881 23331 919 23365
rect 953 23331 984 23365
rect 520 23291 984 23331
rect 520 23257 703 23291
rect 737 23257 775 23291
rect 809 23257 847 23291
rect 881 23257 919 23291
rect 953 23257 984 23291
rect 520 23245 984 23257
rect 520 23244 683 23245
tri 683 23244 684 23245 nw
rect 520 23218 657 23244
tri 657 23218 683 23244 nw
rect 520 23194 633 23218
tri 633 23194 657 23218 nw
tri 1031 23194 1034 23197 se
rect 1034 23194 1086 25744
tri 1021 23184 1031 23194 se
rect 1031 23184 1086 23194
tri 1020 23183 1021 23184 se
rect 1021 23183 1086 23184
tri 1009 23172 1020 23183 se
rect 1020 23172 1086 23183
rect 1034 23120 1086 23172
rect 1114 23242 1166 25744
rect 1194 25533 3320 25686
rect 1194 25520 2297 25533
tri 2068 25499 2089 25520 ne
rect 2089 25499 2297 25520
rect 2331 25499 2373 25533
rect 2407 25499 2449 25533
rect 2483 25499 2525 25533
rect 2559 25499 2601 25533
rect 2635 25499 2677 25533
rect 2711 25499 2753 25533
rect 2787 25499 2829 25533
rect 2863 25499 2904 25533
rect 2938 25499 2979 25533
rect 3013 25499 3054 25533
rect 3088 25499 3129 25533
rect 3163 25499 3320 25533
tri 2089 25461 2127 25499 ne
rect 2127 25461 3320 25499
tri 2127 25427 2161 25461 ne
rect 2161 25427 2297 25461
rect 2331 25427 2373 25461
rect 2407 25427 2449 25461
rect 2483 25427 2525 25461
rect 2559 25427 2601 25461
rect 2635 25427 2677 25461
rect 2711 25427 2753 25461
rect 2787 25427 2829 25461
rect 2863 25427 2904 25461
rect 2938 25427 2979 25461
rect 3013 25427 3054 25461
rect 3088 25427 3129 25461
rect 3163 25427 3320 25461
tri 2161 25389 2199 25427 ne
rect 2199 25389 3320 25427
tri 2199 25355 2233 25389 ne
rect 2233 25355 2297 25389
rect 2331 25355 2373 25389
rect 2407 25355 2449 25389
rect 2483 25355 2525 25389
rect 2559 25355 2601 25389
rect 2635 25355 2677 25389
rect 2711 25355 2753 25389
rect 2787 25355 2829 25389
rect 2863 25355 2904 25389
rect 2938 25355 2979 25389
rect 3013 25355 3054 25389
rect 3088 25355 3129 25389
rect 3163 25355 3320 25389
tri 2233 25353 2235 25355 ne
rect 2235 25353 3320 25355
rect 1114 23178 1166 23190
rect 1114 23120 1166 23126
rect 1194 25347 2099 25353
rect 1194 25341 1274 25347
rect 1194 25307 1200 25341
rect 1234 25313 1274 25341
rect 1308 25313 1352 25347
rect 1386 25313 1430 25347
rect 1464 25313 1508 25347
rect 1542 25313 1587 25347
rect 1621 25313 1666 25347
rect 1700 25313 1745 25347
rect 1779 25313 1824 25347
rect 1858 25313 1903 25347
rect 1937 25313 1982 25347
rect 2016 25341 2099 25347
rect 2016 25313 2056 25341
rect 1234 25307 2056 25313
rect 2090 25307 2099 25341
tri 2235 25337 2251 25353 ne
rect 1194 25283 1241 25307
tri 1241 25283 1265 25307 nw
tri 2022 25283 2046 25307 ne
rect 2046 25283 2099 25307
rect 1194 25267 1240 25283
tri 1240 25282 1241 25283 nw
tri 2046 25282 2047 25283 ne
rect 1194 25233 1200 25267
rect 1234 25233 1240 25267
rect 1194 25193 1240 25233
rect 1194 25159 1200 25193
rect 1234 25159 1240 25193
rect 2047 25268 2099 25283
rect 2047 25234 2056 25268
rect 2090 25234 2099 25268
rect 2047 25195 2099 25234
rect 1194 25119 1240 25159
rect 1194 25085 1200 25119
rect 1234 25085 1240 25119
rect 1194 25045 1240 25085
rect 1194 25011 1200 25045
rect 1234 25011 1240 25045
rect 1194 24971 1240 25011
rect 1194 24937 1200 24971
rect 1234 24937 1240 24971
rect 1194 24897 1240 24937
rect 1194 24863 1200 24897
rect 1234 24863 1240 24897
rect 1194 24824 1240 24863
rect 1194 24790 1200 24824
rect 1234 24790 1240 24824
rect 1194 24751 1240 24790
rect 1194 24717 1200 24751
rect 1234 24717 1240 24751
rect 1194 24678 1240 24717
rect 1194 24644 1200 24678
rect 1234 24644 1240 24678
rect 1194 24605 1240 24644
rect 1194 24571 1200 24605
rect 1234 24571 1240 24605
rect 1194 24532 1240 24571
rect 1194 24498 1200 24532
rect 1234 24498 1240 24532
rect 1194 24459 1240 24498
rect 1194 24425 1200 24459
rect 1234 24425 1240 24459
rect 1194 24386 1240 24425
rect 1194 24352 1200 24386
rect 1234 24352 1240 24386
rect 1194 24313 1240 24352
rect 1194 24279 1200 24313
rect 1234 24279 1240 24313
rect 1194 24240 1240 24279
rect 1194 24206 1200 24240
rect 1234 24206 1240 24240
rect 1194 24167 1240 24206
rect 1194 24133 1200 24167
rect 1234 24133 1240 24167
rect 1194 24094 1240 24133
rect 1194 24060 1200 24094
rect 1234 24060 1240 24094
rect 1194 24021 1240 24060
rect 1194 23987 1200 24021
rect 1234 23987 1240 24021
rect 1307 23998 1359 25170
rect 1619 23999 1671 25170
rect 1931 24934 1983 25170
tri 1906 24923 1917 24934 ne
rect 1917 24923 1983 24934
tri 1917 24909 1931 24923 ne
rect 1194 23948 1240 23987
rect 1194 23914 1200 23948
rect 1234 23914 1240 23948
rect 1194 23875 1240 23914
rect 1194 23841 1200 23875
rect 1234 23841 1240 23875
rect 1194 23802 1240 23841
rect 1194 23768 1200 23802
rect 1234 23768 1240 23802
rect 1194 23729 1240 23768
rect 1194 23695 1200 23729
rect 1234 23695 1240 23729
rect 1194 23656 1240 23695
rect 1194 23622 1200 23656
rect 1234 23622 1240 23656
rect 1194 23583 1240 23622
rect 1194 23549 1200 23583
rect 1234 23549 1240 23583
rect 1931 23984 1983 24923
rect 2047 25161 2056 25195
rect 2090 25161 2099 25195
rect 2047 25122 2099 25161
rect 2047 25088 2056 25122
rect 2090 25088 2099 25122
rect 2047 25049 2099 25088
rect 2047 25015 2056 25049
rect 2090 25015 2099 25049
rect 2047 24976 2099 25015
rect 2047 24942 2056 24976
rect 2090 24942 2099 24976
rect 2047 24903 2099 24942
rect 2047 24869 2056 24903
rect 2090 24869 2099 24903
rect 2047 24830 2099 24869
rect 2047 24796 2056 24830
rect 2090 24796 2099 24830
rect 2047 24757 2099 24796
rect 2047 24723 2056 24757
rect 2090 24723 2099 24757
rect 2251 25317 3320 25353
rect 2251 25283 2297 25317
rect 2331 25283 2373 25317
rect 2407 25283 2449 25317
rect 2483 25283 2525 25317
rect 2559 25283 2601 25317
rect 2635 25283 2677 25317
rect 2711 25283 2753 25317
rect 2787 25283 2829 25317
rect 2863 25283 2904 25317
rect 2938 25283 2979 25317
rect 3013 25283 3054 25317
rect 3088 25283 3129 25317
rect 3163 25283 3320 25317
rect 2251 25245 3320 25283
rect 2251 25211 2297 25245
rect 2331 25211 2373 25245
rect 2407 25211 2449 25245
rect 2483 25211 2525 25245
rect 2559 25211 2601 25245
rect 2635 25211 2677 25245
rect 2711 25211 2753 25245
rect 2787 25211 2829 25245
rect 2863 25211 2904 25245
rect 2938 25211 2979 25245
rect 3013 25211 3054 25245
rect 3088 25211 3129 25245
rect 3163 25211 3320 25245
rect 2251 25173 3320 25211
rect 2251 25139 2297 25173
rect 2331 25139 2373 25173
rect 2407 25139 2449 25173
rect 2483 25139 2525 25173
rect 2559 25139 2601 25173
rect 2635 25139 2677 25173
rect 2711 25139 2753 25173
rect 2787 25139 2829 25173
rect 2863 25139 2904 25173
rect 2938 25139 2979 25173
rect 3013 25139 3054 25173
rect 3088 25139 3129 25173
rect 3163 25139 3320 25173
rect 2251 25101 3320 25139
rect 2251 25067 2297 25101
rect 2331 25067 2373 25101
rect 2407 25067 2449 25101
rect 2483 25067 2525 25101
rect 2559 25067 2601 25101
rect 2635 25067 2677 25101
rect 2711 25067 2753 25101
rect 2787 25067 2829 25101
rect 2863 25067 2904 25101
rect 2938 25067 2979 25101
rect 3013 25067 3054 25101
rect 3088 25067 3129 25101
rect 3163 25067 3320 25101
rect 2251 25029 3320 25067
rect 2251 24995 2297 25029
rect 2331 24995 2373 25029
rect 2407 24995 2449 25029
rect 2483 24995 2525 25029
rect 2559 24995 2601 25029
rect 2635 24995 2677 25029
rect 2711 24995 2753 25029
rect 2787 24995 2829 25029
rect 2863 24995 2904 25029
rect 2938 24995 2979 25029
rect 3013 24995 3054 25029
rect 3088 24995 3129 25029
rect 3163 24995 3320 25029
rect 2251 24957 3320 24995
rect 2251 24923 2297 24957
rect 2331 24923 2373 24957
rect 2407 24923 2449 24957
rect 2483 24923 2525 24957
rect 2559 24923 2601 24957
rect 2635 24923 2677 24957
rect 2711 24923 2753 24957
rect 2787 24923 2829 24957
rect 2863 24923 2904 24957
rect 2938 24923 2979 24957
rect 3013 24923 3054 24957
rect 3088 24923 3129 24957
rect 3163 24923 3320 24957
rect 2251 24885 3320 24923
rect 2251 24851 2297 24885
rect 2331 24851 2373 24885
rect 2407 24851 2449 24885
rect 2483 24851 2525 24885
rect 2559 24851 2601 24885
rect 2635 24851 2677 24885
rect 2711 24851 2753 24885
rect 2787 24851 2829 24885
rect 2863 24851 2904 24885
rect 2938 24851 2979 24885
rect 3013 24851 3054 24885
rect 3088 24851 3129 24885
rect 3163 24851 3320 24885
rect 2251 24813 3320 24851
rect 2251 24779 2297 24813
rect 2331 24779 2373 24813
rect 2407 24779 2449 24813
rect 2483 24779 2525 24813
rect 2559 24779 2601 24813
rect 2635 24779 2677 24813
rect 2711 24779 2753 24813
rect 2787 24779 2829 24813
rect 2863 24779 2904 24813
rect 2938 24779 2979 24813
rect 3013 24779 3054 24813
rect 3088 24779 3129 24813
rect 3163 24779 3320 24813
rect 2251 24736 3320 24779
rect 2047 24684 2099 24723
rect 2047 24650 2056 24684
rect 2090 24650 2099 24684
rect 2047 24612 2099 24650
rect 2047 24578 2056 24612
rect 2090 24578 2099 24612
tri 3139 24587 3288 24736 ne
rect 3288 24587 3320 24736
rect 2047 24562 2099 24578
tri 2099 24562 2124 24587 sw
tri 3288 24583 3292 24587 ne
rect 3292 24583 3320 24587
rect 2047 24556 2955 24562
rect 2047 24540 2130 24556
rect 2047 24506 2056 24540
rect 2090 24522 2130 24540
rect 2164 24522 2207 24556
rect 2241 24522 2284 24556
rect 2318 24522 2361 24556
rect 2395 24522 2438 24556
rect 2472 24522 2515 24556
rect 2549 24522 2592 24556
rect 2626 24522 2669 24556
rect 2703 24522 2746 24556
rect 2780 24522 2823 24556
rect 2857 24522 2900 24556
rect 2934 24522 2955 24556
rect 2090 24516 2955 24522
rect 2090 24506 2099 24516
rect 2047 24468 2099 24506
tri 2099 24491 2124 24516 nw
tri 2878 24491 2903 24516 ne
rect 2047 24434 2056 24468
rect 2090 24434 2099 24468
rect 2047 24427 2099 24434
rect 2903 24461 2955 24516
rect 2903 24427 2912 24461
rect 2946 24427 2955 24461
rect 2047 24363 2056 24375
rect 2090 24363 2099 24375
rect 2047 24299 2056 24311
rect 2090 24299 2099 24311
rect 2047 24235 2056 24247
rect 2090 24235 2099 24247
rect 2047 24180 2099 24183
rect 2047 24171 2056 24180
rect 2090 24171 2099 24180
rect 2047 24108 2099 24119
rect 2047 24074 2056 24108
rect 2090 24074 2099 24108
rect 2047 24036 2099 24074
rect 2047 24002 2056 24036
rect 2090 24002 2099 24036
rect 1619 23935 1671 23947
rect 1619 23871 1671 23883
rect 1619 23807 1671 23819
rect 1619 23743 1671 23755
rect 1619 23679 1671 23691
rect 1619 23615 1671 23627
rect 1619 23557 1671 23563
rect 2047 23964 2099 24002
rect 2047 23930 2056 23964
rect 2090 23930 2099 23964
rect 2047 23892 2099 23930
rect 2047 23858 2056 23892
rect 2090 23858 2099 23892
rect 2047 23820 2099 23858
rect 2047 23786 2056 23820
rect 2090 23786 2099 23820
rect 2047 23748 2099 23786
rect 2047 23714 2056 23748
rect 2090 23714 2099 23748
rect 2047 23676 2099 23714
rect 2047 23642 2056 23676
rect 2090 23642 2099 23676
rect 2047 23604 2099 23642
rect 2047 23570 2056 23604
rect 2090 23570 2099 23604
rect 1194 23510 1240 23549
rect 1194 23476 1200 23510
rect 1234 23476 1240 23510
rect 1194 23437 1240 23476
rect 1194 23403 1200 23437
rect 1234 23403 1240 23437
rect 1194 23364 1240 23403
rect 1194 23330 1200 23364
rect 1234 23330 1240 23364
rect 2047 23532 2099 23570
rect 2047 23498 2056 23532
rect 2090 23498 2099 23532
rect 2047 23460 2099 23498
rect 2047 23426 2056 23460
rect 2090 23426 2099 23460
rect 2047 23388 2099 23426
rect 1194 23291 1240 23330
rect 1194 23257 1200 23291
rect 1234 23257 1240 23291
rect 1194 23218 1240 23257
rect 1194 23184 1200 23218
rect 1234 23184 1240 23218
rect 1307 23216 1359 23358
rect 2047 23354 2056 23388
rect 2090 23354 2099 23388
rect 2047 23316 2099 23354
rect 2047 23282 2056 23316
rect 2090 23282 2099 23316
rect 1466 23216 1472 23268
rect 1524 23216 1536 23268
rect 1588 23216 1600 23268
rect 1652 23216 1664 23268
rect 1716 23216 1728 23268
rect 1780 23216 1786 23268
rect 2047 23244 2099 23282
rect 1194 23145 1240 23184
rect 2047 23210 2056 23244
rect 2090 23210 2099 23244
rect 2047 23172 2099 23210
rect 1194 23111 1200 23145
rect 1234 23111 1240 23145
tri 1190 23100 1194 23104 se
rect 1194 23100 1240 23111
rect 1406 23107 1412 23159
rect 1464 23107 1476 23159
rect 1528 23107 1534 23159
rect 2047 23138 2056 23172
rect 2090 23138 2099 23172
tri 1240 23100 1244 23104 sw
tri 2043 23100 2047 23104 se
rect 2047 23100 2099 23138
tri 1169 23079 1190 23100 se
rect 1190 23079 1244 23100
tri 1244 23079 1265 23100 sw
tri 2022 23079 2043 23100 se
rect 2043 23079 2056 23100
rect 810 23073 2056 23079
rect 810 23039 822 23073
rect 856 23039 894 23073
rect 928 23039 966 23073
rect 1000 23039 1038 23073
rect 1072 23039 1110 23073
rect 1144 23039 1182 23073
rect 1216 23039 1254 23073
rect 1288 23039 1326 23073
rect 1360 23039 1398 23073
rect 1432 23039 1471 23073
rect 1505 23039 1544 23073
rect 1578 23039 1617 23073
rect 1651 23039 1690 23073
rect 1724 23039 1763 23073
rect 1797 23039 1836 23073
rect 1870 23039 1909 23073
rect 1943 23039 1982 23073
rect 2016 23066 2056 23073
rect 2090 23066 2099 23100
rect 2016 23039 2099 23066
rect 2163 24257 2215 24426
rect 2475 24257 2527 24426
rect 2787 24257 2839 24426
rect 2163 24242 2225 24257
tri 2225 24242 2240 24257 nw
tri 2450 24242 2465 24257 ne
rect 2465 24242 2537 24257
tri 2537 24242 2552 24257 nw
tri 2762 24242 2777 24257 ne
rect 2777 24242 2839 24257
rect 2163 23051 2215 24242
tri 2215 24232 2225 24242 nw
tri 2465 24232 2475 24242 ne
rect 2475 23221 2527 24242
tri 2527 24232 2537 24242 nw
tri 2777 24232 2787 24242 ne
rect 2787 23221 2839 24242
rect 2903 24363 2912 24375
rect 2946 24363 2955 24375
rect 2903 24299 2912 24311
rect 2946 24299 2955 24311
rect 2903 24242 2955 24247
rect 2903 24235 2912 24242
rect 2946 24235 2955 24242
rect 2903 24171 2955 24183
rect 2903 24096 2955 24119
rect 2903 24062 2912 24096
rect 2946 24062 2955 24096
rect 2903 24023 2955 24062
rect 2903 23989 2912 24023
rect 2946 23989 2955 24023
rect 2903 23950 2955 23989
rect 2903 23916 2912 23950
rect 2946 23916 2955 23950
rect 2903 23877 2955 23916
rect 2903 23843 2912 23877
rect 2946 23843 2955 23877
rect 2903 23804 2955 23843
rect 2903 23770 2912 23804
rect 2946 23770 2955 23804
rect 2903 23731 2955 23770
rect 2903 23697 2912 23731
rect 2946 23697 2955 23731
rect 2903 23658 2955 23697
rect 2903 23624 2912 23658
rect 2946 23624 2955 23658
rect 2903 23585 2955 23624
rect 2903 23551 2912 23585
rect 2946 23551 2955 23585
rect 2903 23512 2955 23551
rect 2903 23478 2912 23512
rect 2946 23478 2955 23512
rect 2903 23439 2955 23478
rect 2903 23405 2912 23439
rect 2946 23405 2955 23439
rect 2903 23365 2955 23405
rect 2903 23331 2912 23365
rect 2946 23331 2955 23365
rect 2903 23291 2955 23331
rect 2903 23257 2912 23291
rect 2946 23257 2955 23291
rect 2903 23217 2955 23257
rect 2903 23183 2912 23217
rect 2946 23183 2955 23217
rect 2903 23143 2955 23183
rect 2903 23109 2912 23143
rect 2946 23109 2955 23143
rect 2903 23069 2955 23109
rect 810 23033 2099 23039
rect 810 23028 876 23033
tri 876 23028 881 23033 nw
tri 2022 23028 2027 23033 ne
rect 2027 23028 2099 23033
rect 810 23001 856 23028
tri 856 23008 876 23028 nw
tri 2027 23008 2047 23028 ne
tri 808 22967 810 22969 se
rect 810 22967 816 23001
rect 850 22967 856 23001
rect 2047 22994 2056 23028
rect 2090 22994 2099 23028
rect 2047 22982 2099 22994
rect 2903 23035 2912 23069
rect 2946 23035 2955 23069
rect 2903 22995 2955 23035
tri 802 22961 808 22967 se
rect 808 22961 856 22967
tri 795 22954 802 22961 se
rect 802 22954 856 22961
rect 2903 22961 2912 22995
rect 2946 22961 2955 22995
tri 790 22949 795 22954 se
rect 795 22949 856 22954
tri 789 22948 790 22949 se
rect 790 22948 855 22949
tri 855 22948 856 22949 nw
rect 988 22948 2225 22954
tri 755 22914 789 22948 se
rect 789 22914 821 22948
tri 821 22914 855 22948 nw
rect 1040 22914 1077 22948
rect 1111 22914 1154 22948
rect 1188 22914 1231 22948
rect 1265 22914 1308 22948
rect 1342 22914 1384 22948
rect 1418 22914 1460 22948
rect 1494 22914 1536 22948
rect 1570 22914 1612 22948
rect 1646 22914 1688 22948
rect 1722 22914 1764 22948
rect 1798 22914 1840 22948
rect 1874 22914 1916 22948
rect 1950 22914 2225 22948
tri 753 22912 755 22914 se
rect 755 22912 799 22914
rect 753 22728 799 22912
tri 799 22892 821 22914 nw
rect 1040 22908 2225 22914
rect 2903 22921 2955 22961
rect 1040 22896 1044 22908
rect 988 22887 1044 22896
tri 1044 22887 1065 22908 nw
rect 2903 22887 2912 22921
rect 2946 22887 2955 22921
rect 988 22884 1040 22887
rect 827 22874 879 22880
tri 1040 22883 1044 22887 nw
rect 988 22826 1040 22832
rect 1077 22828 1083 22880
rect 1135 22828 1147 22880
rect 1199 22828 2322 22880
rect 1077 22826 2322 22828
tri 2120 22823 2123 22826 ne
rect 2123 22823 2322 22826
rect 827 22813 879 22822
tri 879 22813 889 22823 sw
tri 2123 22813 2133 22823 ne
rect 2133 22813 2322 22823
rect 827 22810 889 22813
rect 879 22798 889 22810
tri 889 22798 904 22813 sw
tri 2133 22798 2148 22813 ne
rect 2148 22798 2322 22813
rect 879 22792 1962 22798
rect 879 22758 999 22792
rect 1033 22758 1076 22792
rect 1110 22758 1153 22792
rect 1187 22758 1230 22792
rect 1264 22758 1307 22792
rect 1341 22758 1384 22792
rect 1418 22758 1460 22792
rect 1494 22758 1536 22792
rect 1570 22758 1612 22792
rect 1646 22758 1688 22792
rect 1722 22758 1764 22792
rect 1798 22758 1840 22792
rect 1874 22758 1916 22792
rect 1950 22758 1962 22792
tri 2148 22774 2172 22798 ne
rect 2172 22774 2322 22798
rect 827 22752 1962 22758
rect 2047 22762 2099 22774
tri 2172 22773 2173 22774 ne
rect 2173 22773 2322 22774
tri 799 22728 811 22740 sw
rect 2047 22728 2056 22762
rect 2090 22728 2099 22762
tri 2173 22739 2207 22773 ne
rect 2207 22739 2322 22773
rect 753 22724 811 22728
tri 811 22724 815 22728 sw
rect 753 22720 815 22724
tri 753 22699 774 22720 ne
rect 774 22710 815 22720
tri 815 22710 829 22724 sw
rect 988 22718 1040 22724
rect 774 22699 829 22710
tri 829 22699 840 22710 sw
tri 774 22698 775 22699 ne
rect 775 22698 840 22699
tri 840 22698 841 22699 sw
rect 901 22698 959 22710
tri 775 22683 790 22698 ne
rect 790 22683 841 22698
tri 841 22683 856 22698 sw
tri 790 22674 799 22683 ne
rect 799 22674 856 22683
tri 799 22664 809 22674 ne
rect 809 22664 856 22674
tri 809 22663 810 22664 ne
rect 810 22552 856 22664
rect 810 22518 816 22552
rect 850 22518 856 22552
rect 810 22476 856 22518
rect 810 22442 816 22476
rect 850 22442 856 22476
rect 810 22400 856 22442
rect 810 22366 816 22400
rect 850 22366 856 22400
rect 810 22324 856 22366
rect 810 22290 816 22324
rect 850 22290 856 22324
rect 810 22248 856 22290
rect 810 22214 816 22248
rect 850 22214 856 22248
rect 810 22172 856 22214
rect 810 22138 816 22172
rect 850 22138 856 22172
rect 810 22096 856 22138
rect 810 22062 816 22096
rect 850 22062 856 22096
rect 810 22020 856 22062
rect 810 21986 816 22020
rect 850 21986 856 22020
rect 810 21943 856 21986
rect 810 21909 816 21943
rect 850 21909 856 21943
rect 810 21866 856 21909
rect 810 21832 816 21866
rect 850 21832 856 21866
rect 810 21789 856 21832
rect 810 21755 816 21789
rect 850 21755 856 21789
rect 810 21712 856 21755
rect 810 21678 816 21712
rect 850 21678 856 21712
rect 810 21635 856 21678
rect 810 21601 816 21635
rect 850 21601 856 21635
rect 810 21558 856 21601
rect 810 21524 816 21558
rect 850 21524 856 21558
rect 901 22664 909 22698
rect 943 22664 959 22698
rect 901 22626 959 22664
rect 901 22592 909 22626
rect 943 22592 959 22626
rect 2047 22687 2099 22728
tri 2207 22699 2247 22739 ne
rect 2247 22699 2322 22739
rect 988 22654 1040 22666
tri 1040 22653 1054 22667 sw
rect 2047 22653 2056 22687
rect 2090 22653 2099 22687
tri 2247 22685 2261 22699 ne
rect 2261 22685 2322 22699
rect 2903 22847 2955 22887
rect 2903 22813 2912 22847
rect 2946 22813 2955 22847
rect 2903 22773 2955 22813
rect 2903 22739 2912 22773
rect 2946 22739 2955 22773
rect 2903 22699 2955 22739
rect 1040 22642 1054 22653
tri 1054 22642 1065 22653 sw
rect 1040 22636 1962 22642
rect 1040 22602 1077 22636
rect 1111 22602 1154 22636
rect 1188 22602 1231 22636
rect 1265 22602 1308 22636
rect 1342 22602 1384 22636
rect 1418 22602 1460 22636
rect 1494 22602 1536 22636
rect 1570 22602 1612 22636
rect 1646 22602 1688 22636
rect 1722 22602 1764 22636
rect 1798 22602 1840 22636
rect 1874 22602 1916 22636
rect 1950 22602 1962 22636
rect 988 22596 1962 22602
rect 2047 22612 2099 22653
rect 901 22498 959 22592
rect 2047 22578 2056 22612
rect 2090 22578 2099 22612
tri 1222 22551 1228 22557 se
rect 1228 22551 1280 22557
tri 1280 22551 1286 22557 sw
tri 1212 22541 1222 22551 se
rect 1222 22541 1286 22551
tri 1286 22541 1296 22551 sw
tri 1207 22536 1212 22541 se
rect 1212 22536 1296 22541
tri 1296 22536 1301 22541 sw
rect 2047 22536 2099 22578
tri 1203 22532 1207 22536 se
rect 1207 22535 1301 22536
rect 1207 22532 1228 22535
rect 901 22464 912 22498
rect 946 22464 959 22498
rect 987 22526 1228 22532
rect 1280 22532 1301 22535
tri 1301 22532 1305 22536 sw
rect 1280 22526 1962 22532
rect 987 22492 999 22526
rect 1033 22492 1076 22526
rect 1110 22492 1153 22526
rect 1187 22492 1228 22526
rect 1280 22492 1307 22526
rect 1341 22492 1384 22526
rect 1418 22492 1460 22526
rect 1494 22492 1536 22526
rect 1570 22492 1612 22526
rect 1646 22492 1688 22526
rect 1722 22492 1764 22526
rect 1798 22492 1840 22526
rect 1874 22492 1916 22526
rect 1950 22492 1962 22526
rect 987 22486 1228 22492
tri 1203 22477 1212 22486 ne
rect 1212 22483 1228 22486
rect 1280 22486 1962 22492
rect 2047 22502 2056 22536
rect 2090 22502 2099 22536
rect 1280 22483 1297 22486
rect 1212 22478 1297 22483
tri 1297 22478 1305 22486 nw
rect 1212 22477 1296 22478
tri 1296 22477 1297 22478 nw
rect 901 22426 959 22464
tri 1212 22461 1228 22477 ne
rect 1228 22471 1280 22477
rect 901 22392 912 22426
rect 946 22392 959 22426
tri 1280 22461 1296 22477 nw
rect 2047 22460 2099 22502
rect 1228 22413 1280 22419
rect 1308 22443 1360 22449
rect 901 21732 959 22392
tri 1291 22384 1308 22401 se
rect 2047 22426 2056 22460
rect 2090 22426 2099 22460
rect 1308 22384 1360 22391
tri 1360 22384 1377 22401 sw
rect 2047 22384 2099 22426
tri 1283 22376 1291 22384 se
rect 1291 22379 1377 22384
rect 1291 22376 1308 22379
rect 987 22370 1308 22376
rect 1360 22376 1377 22379
tri 1377 22376 1385 22384 sw
rect 1360 22370 1962 22376
rect 987 22336 999 22370
rect 1033 22336 1076 22370
rect 1110 22336 1153 22370
rect 1187 22336 1230 22370
rect 1264 22336 1307 22370
rect 1360 22336 1384 22370
rect 1418 22336 1460 22370
rect 1494 22336 1536 22370
rect 1570 22336 1612 22370
rect 1646 22336 1688 22370
rect 1722 22336 1764 22370
rect 1798 22336 1840 22370
rect 1874 22336 1916 22370
rect 1950 22336 1962 22370
rect 987 22330 1308 22336
tri 1283 22329 1284 22330 ne
rect 1284 22329 1308 22330
tri 1284 22321 1292 22329 ne
rect 1292 22327 1308 22329
rect 1360 22330 1962 22336
rect 2047 22350 2056 22384
rect 2090 22350 2099 22384
rect 2047 22330 2099 22350
rect 1360 22329 1384 22330
tri 1384 22329 1385 22330 nw
rect 1360 22327 1376 22329
rect 1292 22321 1376 22327
tri 1376 22321 1384 22329 nw
tri 1292 22308 1305 22321 ne
rect 1305 22308 1363 22321
tri 1363 22308 1376 22321 nw
tri 1305 22305 1308 22308 ne
rect 1308 22305 1360 22308
tri 1360 22305 1363 22308 nw
rect 2047 22274 2056 22278
rect 2090 22274 2099 22278
rect 2047 22266 2099 22274
tri 1363 22198 1385 22220 ne
rect 1385 22198 1388 22220
tri 1385 22195 1388 22198 ne
rect 1440 22198 1443 22220
tri 1443 22198 1465 22220 nw
rect 2047 22202 2056 22214
rect 2090 22202 2099 22214
tri 1440 22195 1443 22198 nw
rect 2047 22138 2056 22150
rect 2090 22138 2099 22150
tri 1455 22122 1468 22135 se
tri 1443 22110 1455 22122 se
rect 1455 22110 1468 22122
tri 1520 22122 1533 22135 sw
rect 1520 22110 1533 22122
tri 1533 22110 1545 22122 sw
rect 2047 22080 2099 22086
rect 2047 22074 2056 22080
rect 2090 22074 2099 22080
tri 1443 22046 1461 22064 ne
rect 1461 22046 1468 22064
tri 1461 22039 1468 22046 ne
rect 1520 22046 1527 22064
tri 1527 22046 1545 22064 nw
tri 1520 22039 1527 22046 nw
rect 2047 22010 2099 22022
tri 1379 21970 1388 21979 se
tri 1368 21959 1379 21970 se
rect 1379 21959 1388 21970
tri 1363 21954 1368 21959 se
rect 1368 21954 1388 21959
tri 1440 21970 1449 21979 sw
rect 1440 21959 1449 21970
tri 1449 21959 1460 21970 sw
rect 1440 21954 1460 21959
tri 1460 21954 1465 21959 sw
rect 2047 21928 2099 21958
rect 2047 21894 2056 21928
rect 2090 21894 2099 21928
rect 2047 21852 2099 21894
rect 2047 21818 2056 21852
rect 2090 21818 2099 21852
tri 1523 21776 1545 21798 ne
rect 1545 21776 1548 21798
tri 1545 21773 1548 21776 ne
rect 1600 21776 1603 21798
tri 1603 21776 1625 21798 nw
rect 2047 21776 2099 21818
tri 1600 21773 1603 21776 nw
rect 901 21680 907 21732
rect 2047 21742 2056 21776
rect 2090 21742 2099 21776
tri 1615 21700 1628 21713 se
tri 1603 21688 1615 21700 se
rect 1615 21688 1628 21700
tri 1680 21700 1693 21713 sw
rect 2047 21700 2099 21742
rect 1680 21688 1693 21700
tri 1693 21688 1705 21700 sw
rect 901 21668 959 21680
rect 901 21616 907 21668
rect 2047 21666 2056 21700
rect 2090 21666 2099 21700
tri 1603 21624 1621 21642 ne
rect 1621 21624 1628 21642
tri 1621 21617 1628 21624 ne
rect 1680 21624 1687 21642
tri 1687 21624 1705 21642 nw
rect 2047 21624 2099 21666
tri 1680 21617 1687 21624 nw
rect 901 21604 959 21616
rect 901 21552 907 21604
rect 2047 21590 2056 21624
rect 2090 21590 2099 21624
rect 901 21546 959 21552
tri 1539 21548 1548 21557 se
tri 1537 21546 1539 21548 se
rect 1539 21546 1548 21548
tri 1523 21532 1537 21546 se
rect 1537 21532 1548 21546
tri 1600 21548 1609 21557 sw
rect 2047 21548 2099 21590
rect 1600 21532 1609 21548
tri 1609 21532 1625 21548 sw
rect 810 21481 856 21524
rect 810 21447 816 21481
rect 850 21447 856 21481
rect 810 21404 856 21447
rect 2047 21514 2056 21548
rect 2090 21514 2099 21548
rect 2163 22664 2215 22685
tri 2261 22670 2276 22685 ne
rect 2276 22670 2322 22685
tri 2276 22665 2281 22670 ne
rect 2281 22665 2322 22670
tri 2281 22625 2321 22665 ne
rect 2321 22625 2322 22665
tri 2321 22624 2322 22625 ne
rect 2475 22664 2527 22685
rect 2163 22600 2215 22612
rect 2163 22536 2215 22548
rect 2163 21731 2215 22484
rect 2475 22600 2527 22612
rect 2475 22536 2527 22548
tri 2215 21731 2219 21735 sw
tri 2471 21731 2475 21735 se
rect 2475 21731 2527 22484
rect 2787 22664 2839 22685
rect 2787 22600 2839 22612
rect 2787 22536 2839 22548
tri 2527 21731 2531 21735 sw
tri 2783 21731 2787 21735 se
rect 2787 21731 2839 22484
rect 2903 22665 2912 22699
rect 2946 22665 2955 22699
rect 2903 22625 2955 22665
rect 2903 22591 2912 22625
rect 2946 22591 2955 22625
rect 2903 22551 2955 22591
rect 2903 22517 2912 22551
rect 2946 22517 2955 22551
rect 2903 22477 2955 22517
rect 2903 22443 2912 22477
rect 2946 22443 2955 22477
rect 2903 22403 2955 22443
rect 2903 22369 2912 22403
rect 2946 22369 2955 22403
rect 2903 22330 2955 22369
rect 2903 22266 2955 22278
rect 2903 22202 2955 22214
rect 2903 22147 2912 22150
rect 2946 22147 2955 22150
rect 2903 22138 2955 22147
rect 2903 22074 2912 22086
rect 2946 22074 2955 22086
rect 2903 22010 2912 22022
rect 2946 22010 2955 22022
rect 2903 21925 2912 21958
rect 2946 21925 2955 21958
rect 2903 21885 2955 21925
rect 2903 21851 2912 21885
rect 2946 21851 2955 21885
rect 2903 21839 2955 21851
tri 17229 21737 17254 21762 ne
tri 17382 21737 17407 21762 nw
rect 2163 21719 2219 21731
tri 2219 21719 2231 21731 sw
tri 2459 21719 2471 21731 se
rect 2471 21719 2531 21731
tri 2531 21719 2543 21731 sw
tri 2771 21719 2783 21731 se
rect 2783 21719 2839 21731
rect 2163 21710 2231 21719
tri 2231 21710 2240 21719 sw
tri 2450 21710 2459 21719 se
rect 2459 21710 2543 21719
tri 2543 21710 2552 21719 sw
tri 2762 21710 2771 21719 se
rect 2771 21710 2839 21719
rect 2163 21541 2215 21710
rect 2475 21541 2527 21710
rect 2787 21541 2839 21710
rect 2906 21719 2952 21731
rect 2906 21685 2912 21719
rect 2946 21685 2952 21719
rect 2906 21645 2952 21685
rect 2906 21611 2912 21645
rect 2946 21611 2952 21645
rect 2906 21599 2952 21611
rect 2047 21472 2099 21514
rect 2047 21438 2056 21472
rect 2090 21438 2099 21472
tri 856 21404 881 21429 sw
tri 2044 21426 2047 21429 se
rect 2047 21426 2099 21438
tri 2099 21426 2102 21429 sw
tri 2022 21404 2044 21426 se
rect 2044 21404 2102 21426
tri 2102 21404 2124 21426 sw
rect 810 21370 816 21404
rect 850 21398 2307 21404
rect 850 21370 890 21398
rect 810 21364 890 21370
rect 924 21364 962 21398
rect 996 21364 1034 21398
rect 1068 21364 1106 21398
rect 1140 21364 1178 21398
rect 1212 21364 1250 21398
rect 1284 21364 1322 21398
rect 1356 21364 1394 21398
rect 1428 21364 1466 21398
rect 1500 21364 1538 21398
rect 1572 21364 1610 21398
rect 1644 21364 1682 21398
rect 1716 21364 1754 21398
rect 1788 21364 1826 21398
rect 1860 21364 1898 21398
rect 1932 21364 1970 21398
rect 2004 21364 2042 21398
rect 2076 21364 2115 21398
rect 2149 21364 2188 21398
rect 2222 21364 2261 21398
rect 2295 21364 2307 21398
rect 810 21358 2307 21364
rect 2850 21089 2958 21143
tri 857 20295 882 20320 nw
rect 1334 20273 2002 20279
rect 1386 20227 2002 20273
rect 2054 20227 2066 20279
rect 2118 20227 2124 20279
rect 1334 20209 1386 20221
tri 1386 20202 1411 20227 nw
rect 1334 20151 1386 20157
rect 1174 19965 1226 19971
rect 1174 19911 1226 19913
tri 1226 19911 1235 19920 sw
rect 1174 19901 1235 19911
rect 1226 19895 1235 19901
tri 1235 19895 1251 19911 sw
tri 1980 19895 1996 19911 se
rect 1996 19895 2002 19911
rect 1226 19859 2002 19895
rect 2054 19859 2066 19911
rect 2118 19859 2124 19911
rect 1226 19849 2124 19859
rect 1174 19843 2124 19849
tri 956 19562 981 19587 se
rect 1014 19434 2232 19440
rect 1066 19388 2232 19434
rect 1014 19370 1066 19382
tri 1066 19363 1091 19388 nw
tri 2079 19363 2104 19388 ne
rect 1014 19312 1066 19318
rect 534 19230 586 19236
rect 534 19166 586 19178
rect 534 19108 586 19114
tri 586 19108 591 19113 sw
rect 534 19088 591 19108
tri 591 19088 611 19108 sw
rect 534 19036 1410 19088
tri 1280 18922 1394 19036 ne
rect 1394 19029 1410 19036
tri 1410 19029 1469 19088 sw
rect 2104 19029 2232 19388
rect 1394 18977 1469 19029
tri 1469 18977 1521 19029 sw
rect 2104 18977 2110 19029
rect 2162 18977 2174 19029
rect 2226 18977 2232 19029
rect 1394 18922 1521 18977
tri 1521 18922 1576 18977 sw
tri 1394 18906 1410 18922 ne
rect 1410 18906 1576 18922
tri 1410 18853 1463 18906 ne
rect 1463 18853 1576 18906
tri 1576 18853 1645 18922 sw
rect 593 18847 1131 18853
rect 645 18795 1131 18847
rect 593 18783 1131 18795
rect 645 18775 1131 18783
tri 645 18750 670 18775 nw
tri 704 18750 729 18775 ne
rect 729 18750 1131 18775
tri 1463 18750 1566 18853 ne
rect 1566 18750 1645 18853
tri 1645 18750 1748 18853 sw
tri 1566 18740 1576 18750 ne
rect 1576 18740 1748 18750
tri 1748 18740 1758 18750 sw
rect 593 18719 645 18731
rect 593 18655 645 18667
rect 593 18591 645 18603
tri 1576 18558 1758 18740 ne
tri 1758 18558 1940 18740 sw
rect 593 18533 645 18539
tri 1758 18533 1783 18558 ne
rect 1783 18533 1940 18558
tri 1940 18533 1965 18558 sw
tri 1783 18376 1940 18533 ne
rect 1940 18376 1965 18533
tri 1965 18376 2122 18533 sw
tri 1940 18354 1962 18376 ne
rect 1962 18354 2122 18376
tri 1137 18308 1183 18354 se
rect 1183 18308 1416 18354
tri 1416 18308 1462 18354 sw
tri 1962 18322 1994 18354 ne
tri 1109 18280 1137 18308 se
rect 1137 18302 1462 18308
rect 1137 18280 1183 18302
tri 1183 18280 1205 18302 nw
tri 1385 18280 1407 18302 ne
rect 1407 18280 1462 18302
tri 1108 18279 1109 18280 se
rect 1109 18279 1182 18280
tri 1182 18279 1183 18280 nw
tri 1407 18279 1408 18280 ne
rect 1408 18279 1462 18280
rect 253 18218 906 18224
rect 253 18166 854 18218
rect 253 18154 906 18166
rect 253 18144 854 18154
rect 253 18038 265 18144
rect 515 18102 854 18144
rect 515 18090 906 18102
rect 515 18038 854 18090
rect 253 18032 906 18038
tri 1107 18032 1108 18033 se
rect 1108 18032 1160 18279
tri 1160 18257 1182 18279 nw
tri 1408 18277 1410 18279 ne
rect 253 17763 527 18032
tri 527 18007 552 18032 nw
tri 1082 18007 1107 18032 se
rect 1107 18011 1160 18032
rect 1107 18007 1108 18011
tri 1034 17959 1082 18007 se
rect 1082 17959 1108 18007
tri 1108 17959 1160 18011 nw
tri 1020 17945 1034 17959 se
rect 1034 17945 1094 17959
tri 1094 17945 1108 17959 nw
rect 614 17939 1042 17945
rect 666 17893 1042 17939
tri 1042 17893 1094 17945 nw
rect 614 17875 666 17887
tri 666 17868 691 17893 nw
rect 614 17817 666 17823
rect 254 17761 526 17762
rect 254 17460 526 17461
rect 253 16628 527 17459
rect 1410 17214 1462 18279
rect 1994 18103 2122 18354
rect 1994 18051 2000 18103
rect 2052 18051 2064 18103
rect 2116 18051 2122 18103
tri 1462 17214 1695 17447 sw
rect 1410 17098 2000 17214
rect 2116 17098 2122 17214
tri 527 16628 615 16716 sw
rect 253 16622 615 16628
rect 253 16588 266 16622
rect 300 16588 341 16622
rect 375 16588 417 16622
rect 451 16588 493 16622
rect 527 16588 569 16622
rect 603 16588 615 16622
rect 253 16554 615 16588
tri 1218 16555 1241 16578 se
rect 1241 16555 1373 16683
tri 615 16554 616 16555 sw
tri 728 16554 729 16555 se
tri 1217 16554 1218 16555 se
rect 1218 16554 1373 16555
rect 253 16550 616 16554
rect 253 16516 266 16550
rect 300 16516 341 16550
rect 375 16516 417 16550
rect 451 16516 493 16550
rect 527 16516 569 16550
rect 603 16530 616 16550
tri 616 16530 640 16554 sw
tri 704 16530 728 16554 se
rect 728 16530 729 16554
rect 603 16516 729 16530
rect 253 16480 729 16516
tri 1131 16529 1156 16554 sw
tri 1192 16529 1217 16554 se
rect 1217 16529 1373 16554
rect 1131 16480 1373 16529
rect 253 16406 1373 16480
rect 174 16254 2124 16378
rect 5161 16365 5473 16371
rect 5161 16313 5163 16365
rect 5215 16313 5227 16365
rect 5279 16313 5291 16365
rect 5343 16313 5355 16365
rect 5407 16313 5419 16365
rect 5471 16313 5473 16365
rect 5161 16295 5473 16313
rect 292 16210 437 16254
tri 437 16210 481 16254 nw
tri 1913 16210 1957 16254 ne
rect 1957 16210 2000 16254
rect 5161 16243 5163 16295
rect 5215 16243 5227 16295
rect 5279 16243 5291 16295
rect 5343 16243 5355 16295
rect 5407 16243 5419 16295
rect 5471 16243 5473 16295
rect 5161 16225 5473 16243
rect 5161 16210 5163 16225
rect 292 16171 398 16210
tri 398 16171 437 16210 nw
tri 1957 16171 1996 16210 ne
rect 1996 16171 2000 16210
rect 292 16137 364 16171
tri 364 16137 398 16171 nw
tri 1996 16167 2000 16171 ne
rect 2219 16173 5163 16210
rect 5215 16173 5227 16225
rect 5279 16173 5291 16225
rect 5343 16173 5355 16225
rect 5407 16173 5419 16225
rect 5471 16210 5473 16225
rect 7741 16365 8053 16371
rect 7741 16313 7743 16365
rect 7795 16313 7807 16365
rect 7859 16313 7871 16365
rect 7923 16313 7935 16365
rect 7987 16313 7999 16365
rect 8051 16313 8053 16365
rect 7741 16295 8053 16313
rect 7741 16243 7743 16295
rect 7795 16243 7807 16295
rect 7859 16243 7871 16295
rect 7923 16243 7935 16295
rect 7987 16243 7999 16295
rect 8051 16243 8053 16295
rect 7741 16225 8053 16243
rect 7741 16210 7743 16225
rect 5471 16173 7743 16210
rect 7795 16173 7807 16225
rect 7859 16173 7871 16225
rect 7923 16173 7935 16225
rect 7987 16173 7999 16225
rect 8051 16210 8053 16225
rect 8514 16365 8826 16371
rect 8514 16313 8516 16365
rect 8568 16313 8580 16365
rect 8632 16313 8644 16365
rect 8696 16313 8708 16365
rect 8760 16313 8772 16365
rect 8824 16313 8826 16365
rect 8514 16295 8826 16313
rect 8514 16243 8516 16295
rect 8568 16243 8580 16295
rect 8632 16243 8644 16295
rect 8696 16243 8708 16295
rect 8760 16243 8772 16295
rect 8824 16243 8826 16295
rect 8514 16225 8826 16243
rect 8514 16210 8516 16225
rect 8051 16173 8516 16210
rect 8568 16173 8580 16225
rect 8632 16173 8644 16225
rect 8696 16173 8708 16225
rect 8760 16173 8772 16225
rect 8824 16210 8826 16225
rect 9338 16365 9650 16371
rect 9338 16313 9340 16365
rect 9392 16313 9404 16365
rect 9456 16313 9468 16365
rect 9520 16313 9532 16365
rect 9584 16313 9596 16365
rect 9648 16313 9650 16365
rect 9338 16295 9650 16313
rect 9338 16243 9340 16295
rect 9392 16243 9404 16295
rect 9456 16243 9468 16295
rect 9520 16243 9532 16295
rect 9584 16243 9596 16295
rect 9648 16243 9650 16295
rect 9338 16225 9650 16243
rect 9338 16210 9340 16225
rect 8824 16173 9340 16210
rect 9392 16173 9404 16225
rect 9456 16173 9468 16225
rect 9520 16173 9532 16225
rect 9584 16173 9596 16225
rect 9648 16210 9650 16225
rect 10321 16365 10633 16371
rect 10321 16313 10323 16365
rect 10375 16313 10387 16365
rect 10439 16313 10451 16365
rect 10503 16313 10515 16365
rect 10567 16313 10579 16365
rect 10631 16313 10633 16365
rect 10321 16295 10633 16313
rect 10321 16243 10323 16295
rect 10375 16243 10387 16295
rect 10439 16243 10451 16295
rect 10503 16243 10515 16295
rect 10567 16243 10579 16295
rect 10631 16243 10633 16295
rect 10321 16225 10633 16243
rect 10321 16210 10323 16225
rect 9648 16173 10323 16210
rect 10375 16173 10387 16225
rect 10439 16173 10451 16225
rect 10503 16173 10515 16225
rect 10567 16173 10579 16225
rect 10631 16210 10633 16225
rect 11811 16365 12123 16371
rect 11811 16313 11813 16365
rect 11865 16313 11877 16365
rect 11929 16313 11941 16365
rect 11993 16313 12005 16365
rect 12057 16313 12069 16365
rect 12121 16313 12123 16365
rect 11811 16295 12123 16313
rect 11811 16243 11813 16295
rect 11865 16243 11877 16295
rect 11929 16243 11941 16295
rect 11993 16243 12005 16295
rect 12057 16243 12069 16295
rect 12121 16243 12123 16295
rect 11811 16225 12123 16243
rect 11811 16210 11813 16225
rect 10631 16173 11813 16210
rect 11865 16173 11877 16225
rect 11929 16173 11941 16225
rect 11993 16173 12005 16225
rect 12057 16173 12069 16225
rect 12121 16210 12123 16225
rect 12633 16365 12945 16371
rect 12633 16313 12635 16365
rect 12687 16313 12699 16365
rect 12751 16313 12763 16365
rect 12815 16313 12827 16365
rect 12879 16313 12891 16365
rect 12943 16313 12945 16365
rect 12633 16295 12945 16313
rect 12633 16243 12635 16295
rect 12687 16243 12699 16295
rect 12751 16243 12763 16295
rect 12815 16243 12827 16295
rect 12879 16243 12891 16295
rect 12943 16243 12945 16295
rect 12633 16225 12945 16243
rect 12633 16210 12635 16225
rect 12121 16173 12635 16210
rect 12687 16173 12699 16225
rect 12751 16173 12763 16225
rect 12815 16173 12827 16225
rect 12879 16173 12891 16225
rect 12943 16210 12945 16225
rect 13456 16365 13768 16371
rect 13456 16313 13458 16365
rect 13510 16313 13522 16365
rect 13574 16313 13586 16365
rect 13638 16313 13650 16365
rect 13702 16313 13714 16365
rect 13766 16313 13768 16365
rect 13456 16295 13768 16313
rect 13456 16243 13458 16295
rect 13510 16243 13522 16295
rect 13574 16243 13586 16295
rect 13638 16243 13650 16295
rect 13702 16243 13714 16295
rect 13766 16243 13768 16295
rect 13456 16225 13768 16243
rect 13456 16210 13458 16225
rect 12943 16173 13458 16210
rect 13510 16173 13522 16225
rect 13574 16173 13586 16225
rect 13638 16173 13650 16225
rect 13702 16173 13714 16225
rect 13766 16210 13768 16225
rect 14285 16365 14597 16371
rect 14285 16313 14287 16365
rect 14339 16313 14351 16365
rect 14403 16313 14415 16365
rect 14467 16313 14479 16365
rect 14531 16313 14543 16365
rect 14595 16313 14597 16365
rect 14285 16295 14597 16313
rect 14285 16243 14287 16295
rect 14339 16243 14351 16295
rect 14403 16243 14415 16295
rect 14467 16243 14479 16295
rect 14531 16243 14543 16295
rect 14595 16243 14597 16295
rect 14285 16225 14597 16243
rect 14285 16210 14287 16225
rect 13766 16173 14287 16210
rect 14339 16173 14351 16225
rect 14403 16173 14415 16225
rect 14467 16173 14479 16225
rect 14531 16173 14543 16225
rect 14595 16210 14597 16225
rect 15109 16365 15421 16371
rect 15109 16313 15111 16365
rect 15163 16313 15175 16365
rect 15227 16313 15239 16365
rect 15291 16313 15303 16365
rect 15355 16313 15367 16365
rect 15419 16313 15421 16365
rect 15109 16295 15421 16313
rect 15109 16243 15111 16295
rect 15163 16243 15175 16295
rect 15227 16243 15239 16295
rect 15291 16243 15303 16295
rect 15355 16243 15367 16295
rect 15419 16243 15421 16295
rect 15109 16225 15421 16243
rect 15109 16210 15111 16225
rect 14595 16173 15111 16210
rect 15163 16173 15175 16225
rect 15227 16173 15239 16225
rect 15291 16173 15303 16225
rect 15355 16173 15367 16225
rect 15419 16210 15421 16225
rect 15932 16365 16244 16371
rect 15932 16313 15934 16365
rect 15986 16313 15998 16365
rect 16050 16313 16062 16365
rect 16114 16313 16126 16365
rect 16178 16313 16190 16365
rect 16242 16313 16244 16365
rect 15932 16295 16244 16313
rect 15932 16243 15934 16295
rect 15986 16243 15998 16295
rect 16050 16243 16062 16295
rect 16114 16243 16126 16295
rect 16178 16243 16190 16295
rect 16242 16243 16244 16295
rect 15932 16225 16244 16243
rect 15932 16210 15934 16225
rect 15419 16173 15934 16210
rect 15986 16173 15998 16225
rect 16050 16173 16062 16225
rect 16114 16173 16126 16225
rect 16178 16173 16190 16225
rect 16242 16210 16244 16225
rect 16747 16212 17025 16218
rect 16747 16210 16764 16212
rect 16242 16173 16764 16210
rect 2219 16171 16764 16173
rect 16816 16171 16828 16212
rect 16880 16171 16892 16212
rect 16944 16171 16956 16212
rect 17008 16210 17025 16212
rect 17008 16171 17030 16210
rect 2219 16137 2231 16171
rect 2265 16137 2304 16171
rect 2338 16137 2377 16171
rect 2411 16137 2450 16171
rect 2484 16137 2523 16171
rect 2557 16137 2596 16171
rect 2630 16137 2669 16171
rect 2703 16137 2742 16171
rect 2776 16137 2815 16171
rect 2849 16137 2888 16171
rect 2922 16137 2961 16171
rect 2995 16137 3034 16171
rect 3068 16137 3107 16171
rect 3141 16137 3180 16171
rect 3214 16137 3253 16171
rect 3287 16137 3326 16171
rect 3360 16137 3399 16171
rect 3433 16137 3472 16171
rect 3506 16137 3545 16171
rect 3579 16137 3618 16171
rect 3652 16137 3691 16171
rect 3725 16137 3764 16171
rect 3798 16137 3837 16171
rect 3871 16137 3910 16171
rect 3944 16137 3983 16171
rect 4017 16137 4056 16171
rect 4090 16137 4129 16171
rect 4163 16137 4202 16171
rect 4236 16137 4275 16171
rect 4309 16137 4348 16171
rect 4382 16137 4421 16171
rect 4455 16137 4494 16171
rect 4528 16137 4567 16171
rect 4601 16137 4640 16171
rect 4674 16137 4713 16171
rect 4747 16137 4786 16171
rect 4820 16137 4859 16171
rect 4893 16137 4932 16171
rect 4966 16137 5005 16171
rect 5039 16137 5078 16171
rect 5112 16137 5151 16171
rect 5185 16155 5224 16171
rect 5258 16155 5297 16171
rect 5331 16155 5370 16171
rect 5404 16155 5443 16171
rect 5215 16137 5224 16155
rect 292 16099 326 16137
tri 326 16099 364 16137 nw
rect 2219 16103 5163 16137
rect 5215 16103 5227 16137
rect 5279 16103 5291 16155
rect 5343 16103 5355 16155
rect 5407 16103 5419 16155
rect 5477 16137 5516 16171
rect 5550 16137 5589 16171
rect 5623 16137 5662 16171
rect 5696 16137 5735 16171
rect 5769 16137 5808 16171
rect 5842 16137 5881 16171
rect 5915 16137 5954 16171
rect 5988 16137 6027 16171
rect 6061 16137 6100 16171
rect 6134 16137 6173 16171
rect 6207 16137 6246 16171
rect 6280 16137 6319 16171
rect 6353 16137 6392 16171
rect 6426 16137 6465 16171
rect 6499 16137 6538 16171
rect 6572 16137 6611 16171
rect 6645 16137 6684 16171
rect 6718 16137 6757 16171
rect 6791 16137 6830 16171
rect 6864 16137 6903 16171
rect 6937 16137 6976 16171
rect 5471 16103 6976 16137
rect 2219 16099 6976 16103
tri 292 16065 326 16099 nw
rect 2219 16065 2231 16099
rect 2265 16065 2304 16099
rect 2338 16065 2377 16099
rect 2411 16065 2450 16099
rect 2484 16065 2523 16099
rect 2557 16065 2596 16099
rect 2630 16065 2669 16099
rect 2703 16065 2742 16099
rect 2776 16065 2815 16099
rect 2849 16065 2888 16099
rect 2922 16065 2961 16099
rect 2995 16065 3034 16099
rect 3068 16065 3107 16099
rect 3141 16065 3180 16099
rect 3214 16065 3253 16099
rect 3287 16065 3326 16099
rect 3360 16065 3399 16099
rect 3433 16065 3472 16099
rect 3506 16065 3545 16099
rect 3579 16065 3618 16099
rect 3652 16065 3691 16099
rect 3725 16065 3764 16099
rect 3798 16065 3837 16099
rect 3871 16065 3910 16099
rect 3944 16065 3983 16099
rect 4017 16065 4056 16099
rect 4090 16065 4129 16099
rect 4163 16065 4202 16099
rect 4236 16065 4275 16099
rect 4309 16065 4348 16099
rect 4382 16065 4421 16099
rect 4455 16065 4494 16099
rect 4528 16065 4567 16099
rect 4601 16065 4640 16099
rect 4674 16065 4713 16099
rect 4747 16065 4786 16099
rect 4820 16065 4859 16099
rect 4893 16065 4932 16099
rect 4966 16065 5005 16099
rect 5039 16065 5078 16099
rect 5112 16065 5151 16099
rect 5185 16085 5224 16099
rect 5258 16085 5297 16099
rect 5331 16085 5370 16099
rect 5404 16085 5443 16099
rect 5215 16065 5224 16085
rect 2219 16033 5163 16065
rect 5215 16033 5227 16065
rect 5279 16033 5291 16085
rect 5343 16033 5355 16085
rect 5407 16033 5419 16085
rect 5477 16065 5516 16099
rect 5550 16065 5589 16099
rect 5623 16065 5662 16099
rect 5696 16065 5735 16099
rect 5769 16065 5808 16099
rect 5842 16065 5881 16099
rect 5915 16065 5954 16099
rect 5988 16065 6027 16099
rect 6061 16065 6100 16099
rect 6134 16065 6173 16099
rect 6207 16065 6246 16099
rect 6280 16065 6319 16099
rect 6353 16065 6392 16099
rect 6426 16065 6465 16099
rect 6499 16065 6538 16099
rect 6572 16065 6611 16099
rect 6645 16065 6684 16099
rect 6718 16065 6757 16099
rect 6791 16065 6830 16099
rect 6864 16065 6903 16099
rect 6937 16065 6976 16099
rect 5471 16033 6976 16065
rect 2219 16027 6976 16033
rect 2219 15993 2231 16027
rect 2265 15993 2304 16027
rect 2338 15993 2377 16027
rect 2411 15993 2450 16027
rect 2484 15993 2523 16027
rect 2557 15993 2596 16027
rect 2630 15993 2669 16027
rect 2703 15993 2742 16027
rect 2776 15993 2815 16027
rect 2849 15993 2888 16027
rect 2922 15993 2961 16027
rect 2995 15993 3034 16027
rect 3068 15993 3107 16027
rect 3141 15993 3180 16027
rect 3214 15993 3253 16027
rect 3287 15993 3326 16027
rect 3360 15993 3399 16027
rect 3433 15993 3472 16027
rect 3506 15993 3545 16027
rect 3579 15993 3618 16027
rect 3652 15993 3691 16027
rect 3725 15993 3764 16027
rect 3798 15993 3837 16027
rect 3871 15993 3910 16027
rect 3944 15993 3983 16027
rect 4017 15993 4056 16027
rect 4090 15993 4129 16027
rect 4163 15993 4202 16027
rect 4236 15993 4275 16027
rect 4309 15993 4348 16027
rect 4382 15993 4421 16027
rect 4455 15993 4494 16027
rect 4528 15993 4567 16027
rect 4601 15993 4640 16027
rect 4674 15993 4713 16027
rect 4747 15993 4786 16027
rect 4820 15993 4859 16027
rect 4893 15993 4932 16027
rect 4966 15993 5005 16027
rect 5039 15993 5078 16027
rect 5112 15993 5151 16027
rect 5185 16015 5224 16027
rect 5258 16015 5297 16027
rect 5331 16015 5370 16027
rect 5404 16015 5443 16027
rect 5215 15993 5224 16015
rect 2219 15963 5163 15993
rect 5215 15963 5227 15993
rect 5279 15963 5291 16015
rect 5343 15963 5355 16015
rect 5407 15963 5419 16015
rect 5477 15993 5516 16027
rect 5550 15993 5589 16027
rect 5623 15993 5662 16027
rect 5696 15993 5735 16027
rect 5769 15993 5808 16027
rect 5842 15993 5881 16027
rect 5915 15993 5954 16027
rect 5988 15993 6027 16027
rect 6061 15993 6100 16027
rect 6134 15993 6173 16027
rect 6207 15993 6246 16027
rect 6280 15993 6319 16027
rect 6353 15993 6392 16027
rect 6426 15993 6465 16027
rect 6499 15993 6538 16027
rect 6572 15993 6611 16027
rect 6645 15993 6684 16027
rect 6718 15993 6757 16027
rect 6791 15993 6830 16027
rect 6864 15993 6903 16027
rect 6937 15993 6976 16027
rect 5471 15963 6976 15993
rect 2219 15955 6976 15963
rect 2219 15921 2231 15955
rect 2265 15921 2304 15955
rect 2338 15921 2377 15955
rect 2411 15921 2450 15955
rect 2484 15921 2523 15955
rect 2557 15921 2596 15955
rect 2630 15921 2669 15955
rect 2703 15921 2742 15955
rect 2776 15921 2815 15955
rect 2849 15921 2888 15955
rect 2922 15921 2961 15955
rect 2995 15921 3034 15955
rect 3068 15921 3107 15955
rect 3141 15921 3180 15955
rect 3214 15921 3253 15955
rect 3287 15921 3326 15955
rect 3360 15921 3399 15955
rect 3433 15921 3472 15955
rect 3506 15921 3545 15955
rect 3579 15921 3618 15955
rect 3652 15921 3691 15955
rect 3725 15921 3764 15955
rect 3798 15921 3837 15955
rect 3871 15921 3910 15955
rect 3944 15921 3983 15955
rect 4017 15921 4056 15955
rect 4090 15921 4129 15955
rect 4163 15921 4202 15955
rect 4236 15921 4275 15955
rect 4309 15921 4348 15955
rect 4382 15921 4421 15955
rect 4455 15921 4494 15955
rect 4528 15921 4567 15955
rect 4601 15921 4640 15955
rect 4674 15921 4713 15955
rect 4747 15921 4786 15955
rect 4820 15921 4859 15955
rect 4893 15921 4932 15955
rect 4966 15921 5005 15955
rect 5039 15921 5078 15955
rect 5112 15921 5151 15955
rect 5185 15945 5224 15955
rect 5258 15945 5297 15955
rect 5331 15945 5370 15955
rect 5404 15945 5443 15955
rect 5215 15921 5224 15945
rect 2219 15893 5163 15921
rect 5215 15893 5227 15921
rect 5279 15893 5291 15945
rect 5343 15893 5355 15945
rect 5407 15893 5419 15945
rect 5477 15921 5516 15955
rect 5550 15921 5589 15955
rect 5623 15921 5662 15955
rect 5696 15921 5735 15955
rect 5769 15921 5808 15955
rect 5842 15921 5881 15955
rect 5915 15921 5954 15955
rect 5988 15921 6027 15955
rect 6061 15921 6100 15955
rect 6134 15921 6173 15955
rect 6207 15921 6246 15955
rect 6280 15921 6319 15955
rect 6353 15921 6392 15955
rect 6426 15921 6465 15955
rect 6499 15921 6538 15955
rect 6572 15921 6611 15955
rect 6645 15921 6684 15955
rect 6718 15921 6757 15955
rect 6791 15921 6830 15955
rect 6864 15921 6903 15955
rect 6937 15921 6976 15955
rect 17018 15921 17030 16171
rect 5471 15893 7743 15921
rect 7795 15893 7807 15921
rect 7859 15893 7871 15921
rect 7923 15893 7935 15921
rect 7987 15893 7999 15921
rect 8051 15893 8516 15921
rect 8568 15893 8580 15921
rect 8632 15893 8644 15921
rect 8696 15893 8708 15921
rect 8760 15893 8772 15921
rect 8824 15893 9340 15921
rect 9392 15893 9404 15921
rect 9456 15893 9468 15921
rect 9520 15893 9532 15921
rect 9584 15893 9596 15921
rect 9648 15893 10323 15921
rect 10375 15893 10387 15921
rect 10439 15893 10451 15921
rect 10503 15893 10515 15921
rect 10567 15893 10579 15921
rect 10631 15893 11813 15921
rect 11865 15893 11877 15921
rect 11929 15893 11941 15921
rect 11993 15893 12005 15921
rect 12057 15893 12069 15921
rect 12121 15893 12635 15921
rect 12687 15893 12699 15921
rect 12751 15893 12763 15921
rect 12815 15893 12827 15921
rect 12879 15893 12891 15921
rect 12943 15893 13458 15921
rect 13510 15893 13522 15921
rect 13574 15893 13586 15921
rect 13638 15893 13650 15921
rect 13702 15893 13714 15921
rect 13766 15893 14287 15921
rect 14339 15893 14351 15921
rect 14403 15893 14415 15921
rect 14467 15893 14479 15921
rect 14531 15893 14543 15921
rect 14595 15893 15111 15921
rect 15163 15893 15175 15921
rect 15227 15893 15239 15921
rect 15291 15893 15303 15921
rect 15355 15893 15367 15921
rect 15419 15893 15934 15921
rect 15986 15893 15998 15921
rect 16050 15893 16062 15921
rect 16114 15893 16126 15921
rect 16178 15893 16190 15921
rect 16242 15893 16764 15921
rect 16816 15893 16828 15921
rect 16880 15893 16892 15921
rect 16944 15893 16956 15921
rect 17008 15893 17030 15921
rect 2219 15882 17030 15893
rect 17059 13801 17254 13943
tri 17254 13801 17396 13943 sw
rect 17059 10736 17564 13801
tri 17564 10736 17713 10885 sw
rect 17059 10492 17713 10736
rect 17059 10263 17254 10492
tri 17254 10263 17483 10492 nw
rect 15650 4379 15656 4431
rect 15708 4379 15720 4431
rect 15772 4379 15778 4431
rect 16040 4345 16418 4397
rect 16470 4345 16482 4397
rect 16534 4345 16540 4397
rect 15897 4271 16540 4274
rect 15718 4253 15770 4259
rect 15897 4219 16333 4271
rect 16385 4219 16397 4271
rect 16449 4219 16540 4271
rect 15897 4216 16540 4219
rect 15718 4189 15770 4201
rect 15598 4137 15718 4188
rect 15598 4131 15770 4137
rect 16415 4173 16467 4179
rect 16415 4109 16467 4121
rect 15656 4057 16415 4103
rect 15656 4046 16467 4057
rect 15718 3828 15770 3834
tri 16616 3791 16654 3829 se
rect 16654 3828 16706 3834
rect 15718 3764 15770 3776
tri 15770 3761 15800 3791 sw
tri 16586 3761 16616 3791 se
rect 16616 3776 16654 3791
rect 16616 3764 16706 3776
rect 16616 3761 16654 3764
rect 15770 3712 16654 3761
rect 15718 3706 16706 3712
rect 3900 3681 4892 3685
rect 3900 3629 3906 3681
rect 3958 3629 3973 3681
rect 4025 3629 4040 3681
rect 4092 3629 4107 3681
rect 4159 3629 4174 3681
rect 4226 3629 4240 3681
rect 4292 3629 4306 3681
rect 4358 3629 4372 3681
rect 4424 3629 4438 3681
rect 4490 3629 4504 3681
rect 4556 3629 4570 3681
rect 4622 3629 4636 3681
rect 4688 3629 4702 3681
rect 4754 3629 4768 3681
rect 4820 3629 4834 3681
rect 4886 3629 4892 3681
rect 3900 3617 4892 3629
rect 3900 3565 3906 3617
rect 3958 3565 3973 3617
rect 4025 3565 4040 3617
rect 4092 3565 4107 3617
rect 4159 3565 4174 3617
rect 4226 3565 4240 3617
rect 4292 3565 4306 3617
rect 4358 3565 4372 3617
rect 4424 3565 4438 3617
rect 4490 3565 4504 3617
rect 4556 3565 4570 3617
rect 4622 3565 4636 3617
rect 4688 3565 4702 3617
rect 4754 3565 4768 3617
rect 4820 3565 4834 3617
rect 4886 3565 4892 3617
rect 3900 3561 4892 3565
rect 5775 3682 6697 3686
rect 5775 3630 5781 3682
rect 5833 3630 5847 3682
rect 5899 3630 5913 3682
rect 5965 3630 5979 3682
rect 6031 3630 6045 3682
rect 6097 3630 6111 3682
rect 6163 3630 6177 3682
rect 6229 3630 6243 3682
rect 6295 3630 6309 3682
rect 6361 3630 6375 3682
rect 6427 3630 6441 3682
rect 6493 3630 6507 3682
rect 6559 3630 6573 3682
rect 6625 3630 6639 3682
rect 6691 3630 6697 3682
rect 5775 3618 6697 3630
rect 5775 3566 5781 3618
rect 5833 3566 5847 3618
rect 5899 3566 5913 3618
rect 5965 3566 5979 3618
rect 6031 3566 6045 3618
rect 6097 3566 6111 3618
rect 6163 3566 6177 3618
rect 6229 3566 6243 3618
rect 6295 3566 6309 3618
rect 6361 3566 6375 3618
rect 6427 3566 6441 3618
rect 6493 3566 6507 3618
rect 6559 3566 6573 3618
rect 6625 3566 6639 3618
rect 6691 3566 6697 3618
rect 5775 3562 6697 3566
rect 7504 3682 8502 3686
rect 7504 3630 7510 3682
rect 7562 3630 7577 3682
rect 7629 3630 7644 3682
rect 7696 3630 7711 3682
rect 7763 3630 7778 3682
rect 7830 3630 7845 3682
rect 7897 3630 7912 3682
rect 7964 3630 7979 3682
rect 8031 3630 8046 3682
rect 8098 3630 8113 3682
rect 8165 3630 8180 3682
rect 8232 3630 8246 3682
rect 8298 3630 8312 3682
rect 8364 3630 8378 3682
rect 8430 3630 8444 3682
rect 8496 3630 8502 3682
rect 7504 3618 8502 3630
rect 7504 3566 7510 3618
rect 7562 3566 7577 3618
rect 7629 3566 7644 3618
rect 7696 3566 7711 3618
rect 7763 3566 7778 3618
rect 7830 3566 7845 3618
rect 7897 3566 7912 3618
rect 7964 3566 7979 3618
rect 8031 3566 8046 3618
rect 8098 3566 8113 3618
rect 8165 3566 8180 3618
rect 8232 3566 8246 3618
rect 8298 3566 8312 3618
rect 8364 3566 8378 3618
rect 8430 3566 8444 3618
rect 8496 3566 8502 3618
rect 7504 3562 8502 3566
rect 9316 3681 10308 3685
rect 9316 3629 9322 3681
rect 9374 3629 9389 3681
rect 9441 3629 9456 3681
rect 9508 3629 9523 3681
rect 9575 3629 9590 3681
rect 9642 3629 9656 3681
rect 9708 3629 9722 3681
rect 9774 3629 9788 3681
rect 9840 3629 9854 3681
rect 9906 3629 9920 3681
rect 9972 3629 9986 3681
rect 10038 3629 10052 3681
rect 10104 3629 10118 3681
rect 10170 3629 10184 3681
rect 10236 3629 10250 3681
rect 10302 3629 10308 3681
rect 9316 3617 10308 3629
rect 9316 3565 9322 3617
rect 9374 3565 9389 3617
rect 9441 3565 9456 3617
rect 9508 3565 9523 3617
rect 9575 3565 9590 3617
rect 9642 3565 9656 3617
rect 9708 3565 9722 3617
rect 9774 3565 9788 3617
rect 9840 3565 9854 3617
rect 9906 3565 9920 3617
rect 9972 3565 9986 3617
rect 10038 3565 10052 3617
rect 10104 3565 10118 3617
rect 10170 3565 10184 3617
rect 10236 3565 10250 3617
rect 10302 3565 10308 3617
rect 9316 3561 10308 3565
rect 11118 3681 12110 3685
rect 11118 3629 11124 3681
rect 11176 3629 11191 3681
rect 11243 3629 11258 3681
rect 11310 3629 11325 3681
rect 11377 3629 11392 3681
rect 11444 3629 11458 3681
rect 11510 3629 11524 3681
rect 11576 3629 11590 3681
rect 11642 3629 11656 3681
rect 11708 3629 11722 3681
rect 11774 3629 11788 3681
rect 11840 3629 11854 3681
rect 11906 3629 11920 3681
rect 11972 3629 11986 3681
rect 12038 3629 12052 3681
rect 12104 3629 12110 3681
rect 11118 3617 12110 3629
rect 11118 3565 11124 3617
rect 11176 3565 11191 3617
rect 11243 3565 11258 3617
rect 11310 3565 11325 3617
rect 11377 3565 11392 3617
rect 11444 3565 11458 3617
rect 11510 3565 11524 3617
rect 11576 3565 11590 3617
rect 11642 3565 11656 3617
rect 11708 3565 11722 3617
rect 11774 3565 11788 3617
rect 11840 3565 11854 3617
rect 11906 3565 11920 3617
rect 11972 3565 11986 3617
rect 12038 3565 12052 3617
rect 12104 3565 12110 3617
rect 11118 3561 12110 3565
rect 12922 3681 13914 3685
rect 12922 3629 12928 3681
rect 12980 3629 12995 3681
rect 13047 3629 13062 3681
rect 13114 3629 13129 3681
rect 13181 3629 13196 3681
rect 13248 3629 13262 3681
rect 13314 3629 13328 3681
rect 13380 3629 13394 3681
rect 13446 3629 13460 3681
rect 13512 3629 13526 3681
rect 13578 3629 13592 3681
rect 13644 3629 13658 3681
rect 13710 3629 13724 3681
rect 13776 3629 13790 3681
rect 13842 3629 13856 3681
rect 13908 3629 13914 3681
rect 12922 3617 13914 3629
rect 12922 3565 12928 3617
rect 12980 3565 12995 3617
rect 13047 3565 13062 3617
rect 13114 3565 13129 3617
rect 13181 3565 13196 3617
rect 13248 3565 13262 3617
rect 13314 3565 13328 3617
rect 13380 3565 13394 3617
rect 13446 3565 13460 3617
rect 13512 3565 13526 3617
rect 13578 3565 13592 3617
rect 13644 3565 13658 3617
rect 13710 3565 13724 3617
rect 13776 3565 13790 3617
rect 13842 3565 13856 3617
rect 13908 3565 13914 3617
rect 12922 3561 13914 3565
rect 14720 3681 15568 3685
rect 14720 3629 14726 3681
rect 14778 3629 14792 3681
rect 14844 3629 14858 3681
rect 14910 3629 14924 3681
rect 14976 3629 14990 3681
rect 15042 3629 15055 3681
rect 15107 3629 15120 3681
rect 15172 3629 15185 3681
rect 15237 3629 15250 3681
rect 15302 3629 15315 3681
rect 15367 3629 15380 3681
rect 15432 3629 15445 3681
rect 15497 3629 15510 3681
rect 15562 3629 15568 3681
rect 14720 3617 15568 3629
rect 14720 3565 14726 3617
rect 14778 3565 14792 3617
rect 14844 3565 14858 3617
rect 14910 3565 14924 3617
rect 14976 3565 14990 3617
rect 15042 3565 15055 3617
rect 15107 3565 15120 3617
rect 15172 3565 15185 3617
rect 15237 3565 15250 3617
rect 15302 3565 15315 3617
rect 15367 3565 15380 3617
rect 15432 3565 15445 3617
rect 15497 3565 15510 3617
rect 15562 3565 15568 3617
rect 14720 3561 15568 3565
rect 17100 3559 17254 3667
tri 16817 3453 16923 3559 ne
rect 16923 3453 17254 3559
tri -2738 3403 -2688 3453 sw
tri 16923 3403 16973 3453 ne
rect 16973 3403 17254 3453
tri 16973 3281 17095 3403 ne
rect 17095 3281 17254 3403
rect -3110 3244 -3058 3250
rect 5168 3229 5174 3281
rect 5226 3229 5240 3281
rect 5292 3229 5306 3281
rect 5358 3229 5372 3281
rect 5424 3229 5438 3281
rect 5490 3229 5503 3281
rect 5555 3229 5568 3281
rect 5620 3229 5633 3281
rect 5685 3229 5691 3281
rect -3110 3180 -3058 3192
tri -3058 3158 -3008 3208 sw
rect 5168 3185 5691 3229
rect -3058 3128 2738 3158
rect -3110 3122 2738 3128
tri 2738 3122 2774 3158 sw
rect 5168 3133 5174 3185
rect 5226 3133 5240 3185
rect 5292 3133 5306 3185
rect 5358 3133 5372 3185
rect 5424 3133 5438 3185
rect 5490 3133 5503 3185
rect 5555 3133 5568 3185
rect 5620 3133 5633 3185
rect 5685 3133 5691 3185
tri 2724 3114 2732 3122 ne
rect 2732 3114 2774 3122
tri 2774 3114 2782 3122 sw
tri 2732 3108 2738 3114 ne
rect 2738 3108 2782 3114
tri 2738 3094 2752 3108 ne
rect 2752 3094 2782 3108
tri 2782 3094 2802 3114 sw
tri -2154 3074 -2134 3094 se
rect -2134 3074 2696 3094
rect -3190 3017 -3138 3023
rect -3106 3022 -3100 3074
rect -3048 3022 -3036 3074
rect -2984 3064 2696 3074
tri 2696 3064 2726 3094 sw
tri 2752 3064 2782 3094 ne
rect 2782 3064 2802 3094
tri 2802 3064 2832 3094 sw
rect -2984 3058 2726 3064
rect -2984 3050 -2102 3058
tri -2102 3050 -2094 3058 nw
tri 2682 3050 2690 3058 ne
rect 2690 3050 2726 3058
tri 2726 3050 2740 3064 sw
tri 2782 3050 2796 3064 ne
rect 2796 3050 2832 3064
tri 2832 3050 2846 3064 sw
rect -2984 3044 -2108 3050
tri -2108 3044 -2102 3050 nw
tri 2690 3044 2696 3050 ne
rect 2696 3044 2740 3050
rect -2984 3038 -2114 3044
tri -2114 3038 -2108 3044 nw
tri 2696 3038 2702 3044 ne
rect 2702 3038 2740 3044
rect -2984 3023 -2977 3038
tri -2977 3023 -2962 3038 nw
tri 2702 3023 2717 3038 ne
rect 2717 3023 2740 3038
tri 2740 3023 2767 3050 sw
tri 2796 3023 2823 3050 ne
rect 2823 3023 2846 3050
tri 2846 3023 2873 3050 sw
rect -2984 3022 -2978 3023
tri -2978 3022 -2977 3023 nw
tri 2717 3022 2718 3023 ne
rect 2718 3022 2767 3023
tri -3196 2977 -3190 2983 se
tri 2718 3005 2735 3022 ne
rect 2735 3014 2767 3022
tri 2767 3014 2776 3023 sw
tri 2823 3014 2832 3023 ne
rect 2832 3014 2873 3023
tri 2873 3014 2882 3023 sw
rect 6097 3022 6149 3056
rect 2735 3005 2776 3014
tri -3138 3000 -3133 3005 sw
tri 2735 3000 2740 3005 ne
rect 2740 3000 2776 3005
tri 2776 3000 2790 3014 sw
tri 2832 3000 2846 3014 ne
rect 2846 3000 2882 3014
tri 2882 3000 2896 3014 sw
rect -3138 2977 -3133 3000
tri -3133 2977 -3110 3000 sw
tri 2740 2977 2763 3000 ne
rect 2763 2977 2790 3000
rect -3190 2953 -3138 2965
tri -3196 2919 -3190 2925 ne
tri 2763 2950 2790 2977 ne
tri 2790 2964 2826 3000 sw
tri 2846 2964 2882 3000 ne
rect 2882 2964 2896 3000
tri 2896 2964 2932 3000 sw
rect 2790 2950 2826 2964
tri 2826 2950 2840 2964 sw
tri 2882 2950 2896 2964 ne
rect 2896 2950 2932 2964
tri 2932 2950 2946 2964 sw
tri 2790 2925 2815 2950 ne
rect 2815 2925 2840 2950
rect -3138 2901 -3135 2925
rect -3190 2900 -3135 2901
tri -3135 2900 -3110 2925 nw
tri 2815 2900 2840 2925 ne
tri 2840 2914 2876 2950 sw
tri 2896 2914 2932 2950 ne
rect 2932 2914 2946 2950
tri 2946 2914 2982 2950 sw
rect 5005 2937 5011 2989
rect 5063 2937 5075 2989
rect 5127 2937 5133 2989
rect 2840 2900 2876 2914
tri 2876 2900 2890 2914 sw
tri 2932 2900 2946 2914 ne
rect 2946 2900 2982 2914
tri 2982 2900 2996 2914 sw
rect -3190 2895 -3138 2900
tri -3138 2897 -3135 2900 nw
rect 1576 2888 1694 2900
tri -2422 2874 -2419 2877 sw
rect 1576 2854 1582 2888
rect 1616 2854 1654 2888
rect 1688 2854 1694 2888
tri -2422 2825 -2419 2828 nw
rect 1576 2815 1694 2854
tri 2840 2850 2890 2900 ne
tri 2890 2864 2926 2900 sw
tri 2946 2864 2982 2900 ne
rect 2982 2864 2996 2900
tri 2996 2864 3032 2900 sw
rect 2890 2850 2926 2864
tri 2926 2850 2940 2864 sw
tri 2982 2850 2996 2864 ne
rect 2996 2850 3032 2864
tri 3032 2850 3046 2864 sw
rect 1576 2813 1654 2815
rect 1576 2779 1582 2813
rect 1616 2781 1654 2813
rect 1688 2781 1694 2815
tri 2890 2800 2940 2850 ne
tri 2940 2814 2976 2850 sw
tri 2996 2814 3032 2850 ne
rect 3032 2814 3046 2850
tri 3046 2814 3082 2850 sw
rect 2940 2800 2976 2814
tri 2976 2800 2990 2814 sw
tri 3032 2800 3046 2814 ne
rect 3046 2800 3082 2814
tri 3082 2800 3096 2814 sw
rect 1616 2779 1694 2781
tri 1252 2742 1254 2744 se
tri 1248 2738 1252 2742 se
rect 1252 2738 1254 2742
tri 1228 2718 1248 2738 se
rect 1248 2718 1254 2738
rect 1576 2742 1694 2779
tri 2940 2750 2990 2800 ne
tri 2990 2764 3026 2800 sw
tri 3046 2764 3082 2800 ne
rect 3082 2764 3096 2800
tri 3096 2764 3132 2800 sw
rect 2990 2750 3026 2764
tri 3026 2750 3040 2764 sw
tri 3082 2750 3096 2764 ne
rect 3096 2750 3132 2764
tri 3132 2750 3146 2764 sw
rect 1576 2738 1654 2742
rect 1576 2704 1582 2738
rect 1616 2708 1654 2738
rect 1688 2708 1694 2742
rect 1616 2704 1694 2708
rect -2502 2669 -2499 2672
tri -2499 2669 -2496 2672 nw
rect 1576 2669 1694 2704
tri 2990 2700 3040 2750 ne
tri 3040 2714 3076 2750 sw
tri 3096 2714 3132 2750 ne
rect 3132 2714 3146 2750
tri 3146 2714 3182 2750 sw
rect 5214 2745 5220 2797
rect 5272 2745 5286 2797
rect 5338 2745 5351 2797
rect 5403 2745 5416 2797
rect 5468 2745 5481 2797
rect 5533 2745 5546 2797
rect 5598 2745 5611 2797
rect 5663 2745 5676 2797
rect 5728 2745 5741 2797
rect 5793 2745 5806 2797
rect 5858 2745 5871 2797
rect 5923 2745 5936 2797
rect 5988 2745 5994 2797
rect 3040 2700 3076 2714
tri 3076 2700 3090 2714 sw
tri 3132 2700 3146 2714 ne
rect 3146 2700 3182 2714
tri 3182 2700 3196 2714 sw
rect 5214 2703 5994 2745
tri -2502 2666 -2499 2669 nw
rect 1576 2663 1654 2669
tri -2738 2629 -2731 2636 sw
rect 1576 2629 1582 2663
rect 1616 2635 1654 2663
rect 1688 2635 1694 2669
tri 3040 2650 3090 2700 ne
tri 3090 2664 3126 2700 sw
tri 3146 2664 3182 2700 ne
rect 3182 2664 3196 2700
tri 3196 2664 3232 2700 sw
rect 3090 2650 3126 2664
tri 3126 2650 3140 2664 sw
tri 3182 2650 3196 2664 ne
rect 3196 2651 3232 2664
tri 3232 2651 3245 2664 sw
rect 5214 2651 5220 2703
rect 5272 2651 5286 2703
rect 5338 2651 5351 2703
rect 5403 2651 5416 2703
rect 5468 2651 5481 2703
rect 5533 2651 5546 2703
rect 5598 2651 5611 2703
rect 5663 2651 5676 2703
rect 5728 2651 5741 2703
rect 5793 2651 5806 2703
rect 5858 2651 5871 2703
rect 5923 2651 5936 2703
rect 5988 2651 5994 2703
rect 6864 2651 7192 3281
rect 8522 3229 8528 3281
rect 8580 3229 8594 3281
rect 8646 3229 8660 3281
rect 8712 3229 8726 3281
rect 8778 3229 8792 3281
rect 8844 3229 8857 3281
rect 8909 3229 8922 3281
rect 8974 3229 8980 3281
rect 8522 3215 8980 3229
rect 8522 3163 8528 3215
rect 8580 3163 8594 3215
rect 8646 3163 8660 3215
rect 8712 3163 8726 3215
rect 8778 3163 8792 3215
rect 8844 3163 8857 3215
rect 8909 3163 8922 3215
rect 8974 3163 8980 3215
tri 17095 3163 17213 3281 ne
rect 17213 3163 17254 3281
tri 17213 3159 17217 3163 ne
rect 17217 3159 17254 3163
rect 8181 3017 8187 3069
rect 8239 3017 8251 3069
rect 8303 3017 8309 3069
rect 7714 2937 7720 2989
rect 7772 2937 7784 2989
rect 7836 2937 7842 2989
rect 8411 2745 8417 2797
rect 8469 2745 8482 2797
rect 8534 2745 8547 2797
rect 8599 2745 8612 2797
rect 8664 2745 8677 2797
rect 8729 2745 8741 2797
rect 8793 2745 8805 2797
rect 8857 2745 8863 2797
rect 8411 2703 8863 2745
rect 8411 2651 8417 2703
rect 8469 2651 8482 2703
rect 8534 2651 8547 2703
rect 8599 2651 8612 2703
rect 8664 2651 8677 2703
rect 8729 2651 8741 2703
rect 8793 2651 8805 2703
rect 8857 2651 8863 2703
rect 3196 2650 3245 2651
tri 3245 2650 3246 2651 sw
rect 1616 2629 1694 2635
rect -2738 2608 -2731 2629
tri -2731 2608 -2710 2629 sw
rect 1576 2596 1694 2629
tri 3090 2600 3140 2650 ne
tri 3140 2614 3176 2650 sw
tri 3196 2614 3232 2650 ne
rect 3232 2614 3246 2650
tri 3246 2614 3282 2650 sw
rect 3140 2600 3176 2614
tri 3176 2600 3190 2614 sw
tri 3232 2600 3246 2614 ne
rect 3246 2600 3282 2614
tri 3282 2600 3296 2614 sw
rect 1576 2588 1654 2596
rect -2738 2554 -2726 2562
tri -2726 2554 -2718 2562 nw
rect 1576 2554 1582 2588
rect 1616 2562 1654 2588
rect 1688 2562 1694 2596
rect 1616 2554 1694 2562
tri -2738 2542 -2726 2554 nw
rect 1576 2523 1694 2554
tri 3140 2550 3190 2600 ne
tri 3190 2564 3226 2600 sw
tri 3246 2564 3282 2600 ne
rect 3282 2564 3296 2600
tri 3296 2564 3332 2600 sw
rect 3190 2550 3226 2564
tri 3226 2550 3240 2564 sw
tri 3282 2550 3296 2564 ne
rect 3296 2550 3332 2564
tri 3332 2550 3346 2564 sw
rect 1576 2513 1654 2523
rect 1576 2479 1582 2513
rect 1616 2489 1654 2513
rect 1688 2489 1694 2523
tri 3190 2500 3240 2550 ne
tri 3240 2514 3276 2550 sw
tri 3296 2514 3332 2550 ne
rect 3332 2514 3346 2550
tri 3346 2514 3382 2550 sw
rect 3240 2500 3276 2514
tri 3276 2500 3290 2514 sw
tri 3332 2500 3346 2514 ne
rect 3346 2500 3382 2514
tri 3382 2500 3396 2514 sw
rect 1616 2479 1694 2489
tri 1226 2456 1248 2478 sw
tri -2582 2453 -2579 2456 sw
rect 1226 2453 1248 2456
tri 1248 2453 1251 2456 sw
tri 779 2452 780 2453 sw
rect 1226 2452 1251 2453
tri 1251 2452 1252 2453 sw
rect 1576 2450 1694 2479
tri 3240 2450 3290 2500 ne
tri 3290 2464 3326 2500 sw
tri 3346 2464 3382 2500 ne
rect 3382 2464 3396 2500
tri 3396 2464 3432 2500 sw
rect 3290 2450 3326 2464
tri 3326 2450 3340 2464 sw
tri 3382 2450 3396 2464 ne
rect 3396 2450 3432 2464
tri 3432 2450 3446 2464 sw
rect 1576 2438 1654 2450
tri -2582 2404 -2579 2407 nw
tri 778 2406 779 2407 ne
rect 1226 2404 1250 2406
tri 1250 2404 1252 2406 nw
rect 1576 2404 1582 2438
rect 1616 2416 1654 2438
rect 1688 2416 1694 2450
rect 1616 2404 1694 2416
tri 1226 2380 1250 2404 nw
rect 1576 2377 1694 2404
tri 3290 2400 3340 2450 ne
tri 3340 2414 3376 2450 sw
tri 3396 2414 3432 2450 ne
rect 3432 2414 3446 2450
tri 3446 2414 3482 2450 sw
rect 3340 2400 3376 2414
tri 3376 2400 3390 2414 sw
tri 3432 2400 3446 2414 ne
rect 3446 2400 3482 2414
tri 3482 2400 3496 2414 sw
rect 1576 2363 1654 2377
rect 1576 2329 1582 2363
rect 1616 2343 1654 2363
rect 1688 2343 1694 2377
tri 3340 2350 3390 2400 ne
tri 3390 2364 3426 2400 sw
tri 3446 2364 3482 2400 ne
rect 3482 2364 3496 2400
tri 3496 2364 3532 2400 sw
rect 3390 2350 3426 2364
tri 3426 2350 3440 2364 sw
tri 3482 2350 3496 2364 ne
rect 3496 2350 3532 2364
tri 3532 2350 3546 2364 sw
rect 1616 2329 1694 2343
rect 1576 2304 1694 2329
rect 1576 2288 1654 2304
rect -3190 2264 -3138 2270
rect 1576 2254 1582 2288
rect 1616 2270 1654 2288
rect 1688 2270 1694 2304
tri 3390 2300 3440 2350 ne
tri 3440 2314 3476 2350 sw
tri 3496 2314 3532 2350 ne
rect 3532 2314 3546 2350
tri 3546 2314 3582 2350 sw
rect 3440 2300 3476 2314
tri 3476 2300 3490 2314 sw
tri 3532 2300 3546 2314 ne
rect 3546 2300 3582 2314
tri 3582 2300 3596 2314 sw
rect 1616 2254 1694 2270
rect 1576 2231 1694 2254
tri 3440 2250 3490 2300 ne
tri 3490 2264 3526 2300 sw
tri 3546 2264 3582 2300 ne
rect 3582 2280 3596 2300
tri 3596 2280 3616 2300 sw
rect 3582 2264 3616 2280
tri 3616 2264 3632 2280 sw
tri 7698 2264 7714 2280 se
rect 7714 2264 7720 2280
rect 3490 2250 3526 2264
tri 3526 2250 3540 2264 sw
tri 3582 2250 3596 2264 ne
rect 3596 2250 7720 2264
tri -3138 2213 -3135 2216 sw
rect 1576 2213 1654 2231
rect -3138 2212 -3135 2213
rect -3190 2200 -3135 2212
rect -3138 2188 -3135 2200
tri -3135 2188 -3110 2213 sw
rect -3138 2176 746 2188
rect -3138 2148 686 2176
rect -3190 2142 686 2148
rect 720 2142 746 2176
tri 654 2138 658 2142 ne
rect 658 2138 746 2142
rect 774 2180 1352 2186
rect 774 2146 786 2180
rect 820 2146 861 2180
rect 895 2146 936 2180
rect 970 2146 1010 2180
rect 1044 2146 1084 2180
rect 1118 2146 1158 2180
rect 1192 2146 1232 2180
rect 1266 2146 1306 2180
rect 1340 2158 1352 2180
rect 1576 2179 1582 2213
rect 1616 2197 1654 2213
rect 1688 2197 1694 2231
tri 3490 2200 3540 2250 ne
tri 3540 2228 3562 2250 sw
tri 3596 2228 3618 2250 ne
rect 3618 2228 7720 2250
rect 7772 2228 7784 2280
rect 7836 2264 7842 2280
tri 7842 2264 7858 2280 sw
rect 7836 2228 7858 2264
rect 3540 2200 3562 2228
tri 3562 2200 3590 2228 sw
rect 1616 2179 1694 2197
tri 1352 2158 1358 2164 sw
rect 1576 2158 1694 2179
tri 3540 2164 3576 2200 ne
rect 3576 2164 5011 2200
rect 1340 2146 1358 2158
rect 774 2140 1358 2146
tri 1358 2140 1376 2158 sw
tri 1310 2138 1312 2140 ne
rect 1312 2138 1376 2140
tri 1376 2138 1378 2140 sw
rect 1576 2138 1654 2158
tri 658 2116 680 2138 ne
rect -3350 2106 -3298 2112
rect 680 2104 746 2138
tri 1312 2130 1320 2138 ne
rect 1320 2130 1378 2138
tri 1378 2130 1386 2138 sw
tri 1320 2120 1330 2130 ne
rect 1330 2120 1386 2130
tri 1330 2110 1340 2120 ne
rect 680 2070 686 2104
rect 720 2070 746 2104
rect 680 2058 746 2070
rect -3350 2042 -3298 2054
tri -3298 2030 -3272 2056 sw
rect -3298 2024 1280 2030
rect -3298 1990 779 2024
rect 813 1990 855 2024
rect 889 1990 931 2024
rect 965 1990 1007 2024
rect 1041 1990 1083 2024
rect 1117 1990 1159 2024
rect 1193 1990 1234 2024
rect 1268 1990 1280 2024
rect -3350 1984 1280 1990
rect -3430 1950 -3378 1956
rect -3430 1886 -3378 1898
tri -3378 1876 -3349 1905 sw
tri 1312 1876 1340 1904 se
rect 1340 1884 1386 2120
rect 1340 1876 1378 1884
tri 1378 1876 1386 1884 nw
rect 1576 2104 1582 2138
rect 1616 2124 1654 2138
rect 1688 2124 1694 2158
tri 4947 2148 4963 2164 ne
rect 4963 2148 5011 2164
rect 5063 2148 5075 2200
rect 5127 2148 5133 2200
rect 1616 2104 1694 2124
rect 1576 2085 1694 2104
rect 1576 2062 1654 2085
rect 1576 2028 1582 2062
rect 1616 2051 1654 2062
rect 1688 2051 1694 2085
rect 1616 2028 1694 2051
rect 1576 2012 1694 2028
rect 1576 1986 1654 2012
rect 1576 1952 1582 1986
rect 1616 1978 1654 1986
rect 1688 1978 1694 2012
rect 1616 1952 1694 1978
rect 1576 1938 1694 1952
rect 1576 1910 1654 1938
rect 1576 1876 1582 1910
rect 1616 1904 1654 1910
rect 1688 1904 1694 1938
rect 1616 1876 1694 1904
rect -3378 1874 -3349 1876
tri -3349 1874 -3347 1876 sw
tri 1310 1874 1312 1876 se
rect 1312 1874 1376 1876
tri 1376 1874 1378 1876 nw
rect -3378 1868 1366 1874
rect -3378 1834 780 1868
rect 814 1834 856 1868
rect 890 1834 931 1868
rect 965 1834 1006 1868
rect 1040 1834 1081 1868
rect 1115 1834 1156 1868
rect 1190 1834 1231 1868
rect 1265 1834 1306 1868
rect 1340 1864 1366 1868
tri 1366 1864 1376 1874 nw
rect 1576 1864 1694 1876
rect 1340 1834 1352 1864
tri 1352 1850 1366 1864 nw
rect -3430 1828 1352 1834
rect 1576 1834 1654 1864
rect 1576 1800 1582 1834
rect 1616 1830 1654 1834
rect 1688 1850 1694 1864
tri 1694 1850 1720 1876 sw
rect 1688 1849 3618 1850
tri 3618 1849 3619 1850 sw
rect 1688 1830 3623 1849
rect 1616 1818 3623 1830
rect 1616 1800 3212 1818
rect 1576 1790 3212 1800
tri 919 1774 934 1789 se
rect 934 1774 986 1789
tri 986 1774 1001 1789 sw
rect -2950 1773 -2898 1774
tri -2898 1773 -2897 1774 sw
tri 918 1773 919 1774 se
rect 919 1773 1001 1774
tri 1001 1773 1002 1774 sw
rect -2950 1768 -2897 1773
rect -2898 1764 -2897 1768
tri -2897 1764 -2888 1773 sw
tri 909 1764 918 1773 se
rect 918 1767 1002 1773
rect 918 1764 934 1767
rect -2898 1758 934 1764
rect 986 1764 1002 1767
tri 1002 1764 1011 1773 sw
rect 986 1758 1352 1764
rect -2898 1724 786 1758
rect 820 1724 861 1758
rect 895 1724 934 1758
rect 986 1724 1010 1758
rect 1044 1724 1084 1758
rect 1118 1724 1158 1758
rect 1192 1724 1232 1758
rect 1266 1724 1306 1758
rect 1340 1724 1352 1758
rect -2898 1718 934 1724
rect -2898 1716 -2874 1718
tri -2874 1716 -2872 1718 nw
tri 909 1716 911 1718 ne
rect 911 1716 934 1718
rect -2950 1704 -2897 1716
rect -2898 1693 -2897 1704
tri -2897 1693 -2874 1716 nw
tri 911 1693 934 1716 ne
rect 986 1718 1352 1724
rect 1576 1758 1654 1790
rect 1576 1724 1582 1758
rect 1616 1756 1654 1758
rect 1688 1766 3212 1790
rect 3264 1766 3283 1818
rect 3335 1766 3354 1818
rect 3406 1766 3425 1818
rect 3477 1766 3495 1818
rect 3547 1766 3565 1818
rect 3617 1766 3623 1818
rect 1688 1756 3623 1766
rect 1616 1735 3623 1756
rect 1616 1724 1694 1735
rect 986 1716 1009 1718
tri 1009 1716 1011 1718 nw
rect 1576 1716 1694 1724
rect 934 1703 986 1715
tri -2898 1692 -2897 1693 nw
rect -2950 1646 -2898 1652
tri 986 1693 1009 1716 nw
rect 1576 1682 1654 1716
rect 1688 1682 1694 1716
tri 1694 1709 1720 1735 nw
rect 934 1645 986 1651
rect 1014 1675 1066 1681
tri 989 1608 1014 1633 se
rect 1576 1648 1582 1682
rect 1616 1648 1694 1682
rect 1576 1642 1694 1648
rect 1014 1611 1066 1623
rect -2870 1556 -2864 1608
rect -2812 1556 -2800 1608
rect -2748 1602 1014 1608
tri 1066 1608 1091 1633 sw
rect 1576 1608 1654 1642
rect 1688 1608 1694 1642
rect 1066 1602 1352 1608
rect -2748 1568 786 1602
rect 820 1568 861 1602
rect 895 1568 936 1602
rect 970 1568 1010 1602
rect 1066 1568 1084 1602
rect 1118 1568 1158 1602
rect 1192 1568 1232 1602
rect 1266 1568 1306 1602
rect 1340 1568 1352 1602
rect -2748 1562 1014 1568
rect -2748 1556 -2742 1562
tri -2742 1556 -2736 1562 nw
tri 989 1556 995 1562 ne
rect 995 1559 1014 1562
rect 1066 1562 1352 1568
rect 1576 1606 1694 1608
rect 1576 1572 1582 1606
rect 1616 1572 1694 1606
rect 1576 1568 1694 1572
rect 1066 1559 1082 1562
rect 995 1556 1082 1559
tri 995 1553 998 1556 ne
rect 998 1553 1082 1556
tri 1082 1553 1091 1562 nw
tri 998 1537 1014 1553 ne
rect 1014 1537 1066 1553
tri 1066 1537 1082 1553 nw
rect 1576 1534 1654 1568
rect 1688 1534 1694 1568
rect 1576 1530 1694 1534
rect 496 1511 614 1523
rect 496 1477 502 1511
rect 536 1477 614 1511
rect 1576 1496 1582 1530
rect 1616 1496 1694 1530
rect 1576 1494 1694 1496
tri 1575 1485 1576 1486 se
rect 1576 1485 1654 1494
rect 496 1460 614 1477
tri 614 1460 639 1485 sw
tri 1550 1460 1575 1485 se
rect 1575 1460 1654 1485
rect 1688 1460 1694 1494
rect 496 1454 1694 1460
rect 496 1420 574 1454
rect 608 1420 646 1454
rect 680 1420 718 1454
rect 752 1420 790 1454
rect 824 1420 862 1454
rect 896 1420 934 1454
rect 968 1420 1006 1454
rect 1040 1420 1078 1454
rect 1112 1420 1150 1454
rect 1184 1420 1222 1454
rect 1256 1420 1294 1454
rect 1328 1420 1366 1454
rect 1400 1420 1438 1454
rect 1472 1420 1510 1454
rect 1544 1420 1582 1454
rect 1616 1420 1694 1454
rect 496 1386 1654 1420
rect 1688 1386 1694 1420
rect 496 1382 1694 1386
rect 496 1348 540 1382
rect 574 1348 617 1382
rect 651 1348 694 1382
rect 728 1348 771 1382
rect 805 1348 848 1382
rect 882 1348 925 1382
rect 959 1348 1002 1382
rect 1036 1348 1079 1382
rect 1113 1348 1156 1382
rect 1190 1348 1232 1382
rect 1266 1348 1308 1382
rect 1342 1348 1384 1382
rect 1418 1348 1460 1382
rect 1494 1348 1536 1382
rect 1570 1348 1694 1382
rect 496 1342 1694 1348
<< rmetal1 >>
rect 253 17762 527 17763
rect 253 17761 254 17762
rect 526 17761 527 17762
rect 253 17460 254 17461
rect 526 17460 527 17461
rect 253 17459 527 17460
<< via1 >>
rect 1114 23190 1166 23242
rect 1114 23126 1166 23178
rect 1619 23947 1671 23999
rect 2047 24396 2099 24427
rect 2047 24375 2056 24396
rect 2056 24375 2090 24396
rect 2090 24375 2099 24396
rect 2047 24362 2056 24363
rect 2056 24362 2090 24363
rect 2090 24362 2099 24363
rect 2047 24324 2099 24362
rect 2047 24311 2056 24324
rect 2056 24311 2090 24324
rect 2090 24311 2099 24324
rect 2047 24290 2056 24299
rect 2056 24290 2090 24299
rect 2090 24290 2099 24299
rect 2047 24252 2099 24290
rect 2047 24247 2056 24252
rect 2056 24247 2090 24252
rect 2090 24247 2099 24252
rect 2047 24218 2056 24235
rect 2056 24218 2090 24235
rect 2090 24218 2099 24235
rect 2047 24183 2099 24218
rect 2047 24146 2056 24171
rect 2056 24146 2090 24171
rect 2090 24146 2099 24171
rect 2047 24119 2099 24146
rect 1619 23883 1671 23935
rect 1619 23819 1671 23871
rect 1619 23755 1671 23807
rect 1619 23691 1671 23743
rect 1619 23627 1671 23679
rect 1619 23563 1671 23615
rect 1472 23216 1524 23268
rect 1536 23216 1588 23268
rect 1600 23216 1652 23268
rect 1664 23216 1716 23268
rect 1728 23216 1780 23268
rect 1412 23107 1464 23159
rect 1476 23107 1528 23159
rect 2903 24388 2955 24427
rect 2903 24375 2912 24388
rect 2912 24375 2946 24388
rect 2946 24375 2955 24388
rect 2903 24354 2912 24363
rect 2912 24354 2946 24363
rect 2946 24354 2955 24363
rect 2903 24315 2955 24354
rect 2903 24311 2912 24315
rect 2912 24311 2946 24315
rect 2946 24311 2955 24315
rect 2903 24281 2912 24299
rect 2912 24281 2946 24299
rect 2946 24281 2955 24299
rect 2903 24247 2955 24281
rect 2903 24208 2912 24235
rect 2912 24208 2946 24235
rect 2946 24208 2955 24235
rect 2903 24183 2955 24208
rect 2903 24169 2955 24171
rect 2903 24135 2912 24169
rect 2912 24135 2946 24169
rect 2946 24135 2955 24169
rect 2903 24119 2955 24135
rect 988 22914 1000 22948
rect 1000 22914 1034 22948
rect 1034 22914 1040 22948
rect 988 22896 1040 22914
rect 827 22822 879 22874
rect 988 22832 1040 22884
rect 1083 22828 1135 22880
rect 1147 22828 1199 22880
rect 827 22758 879 22810
rect 988 22666 1040 22718
rect 988 22636 1040 22654
rect 988 22602 1000 22636
rect 1000 22602 1034 22636
rect 1034 22602 1040 22636
rect 1228 22526 1280 22535
rect 1228 22492 1230 22526
rect 1230 22492 1264 22526
rect 1264 22492 1280 22526
rect 1228 22483 1280 22492
rect 1228 22419 1280 22471
rect 1308 22391 1360 22443
rect 1308 22370 1360 22379
rect 1308 22336 1341 22370
rect 1341 22336 1360 22370
rect 1308 22327 1360 22336
rect 2047 22308 2099 22330
rect 2047 22278 2056 22308
rect 2056 22278 2090 22308
rect 2090 22278 2099 22308
rect 2047 22232 2099 22266
rect 2047 22214 2056 22232
rect 2056 22214 2090 22232
rect 2090 22214 2099 22232
rect 2047 22198 2056 22202
rect 2056 22198 2090 22202
rect 2090 22198 2099 22202
rect 2047 22156 2099 22198
rect 2047 22150 2056 22156
rect 2056 22150 2090 22156
rect 2090 22150 2099 22156
rect 2047 22122 2056 22138
rect 2056 22122 2090 22138
rect 2090 22122 2099 22138
rect 2047 22086 2099 22122
rect 2047 22046 2056 22074
rect 2056 22046 2090 22074
rect 2090 22046 2099 22074
rect 2047 22022 2099 22046
rect 2047 22004 2099 22010
rect 2047 21970 2056 22004
rect 2056 21970 2090 22004
rect 2090 21970 2099 22004
rect 2047 21958 2099 21970
rect 907 21680 959 21732
rect 907 21616 959 21668
rect 907 21552 959 21604
rect 2163 22612 2215 22664
rect 2163 22548 2215 22600
rect 2163 22484 2215 22536
rect 2475 22612 2527 22664
rect 2475 22548 2527 22600
rect 2475 22484 2527 22536
rect 2787 22612 2839 22664
rect 2787 22548 2839 22600
rect 2787 22484 2839 22536
rect 2903 22329 2955 22330
rect 2903 22295 2912 22329
rect 2912 22295 2946 22329
rect 2946 22295 2955 22329
rect 2903 22278 2955 22295
rect 2903 22255 2955 22266
rect 2903 22221 2912 22255
rect 2912 22221 2946 22255
rect 2946 22221 2955 22255
rect 2903 22214 2955 22221
rect 2903 22181 2955 22202
rect 2903 22150 2912 22181
rect 2912 22150 2946 22181
rect 2946 22150 2955 22181
rect 2903 22107 2955 22138
rect 2903 22086 2912 22107
rect 2912 22086 2946 22107
rect 2946 22086 2955 22107
rect 2903 22073 2912 22074
rect 2912 22073 2946 22074
rect 2946 22073 2955 22074
rect 2903 22033 2955 22073
rect 2903 22022 2912 22033
rect 2912 22022 2946 22033
rect 2946 22022 2955 22033
rect 2903 21999 2912 22010
rect 2912 21999 2946 22010
rect 2946 21999 2955 22010
rect 2903 21959 2955 21999
rect 2903 21958 2912 21959
rect 2912 21958 2946 21959
rect 2946 21958 2955 21959
rect 1334 20221 1386 20273
rect 2002 20227 2054 20279
rect 2066 20227 2118 20279
rect 1334 20157 1386 20209
rect 1174 19913 1226 19965
rect 1174 19849 1226 19901
rect 2002 19859 2054 19911
rect 2066 19859 2118 19911
rect 1014 19382 1066 19434
rect 1014 19318 1066 19370
rect 534 19178 586 19230
rect 534 19114 586 19166
rect 2110 18977 2162 19029
rect 2174 18977 2226 19029
rect 593 18795 645 18847
rect 593 18731 645 18783
rect 593 18667 645 18719
rect 593 18603 645 18655
rect 593 18539 645 18591
rect 854 18166 906 18218
rect 854 18102 906 18154
rect 854 18038 906 18090
rect 614 17887 666 17939
rect 614 17823 666 17875
rect 2000 18051 2052 18103
rect 2064 18051 2116 18103
rect 2000 17098 2116 17214
rect 5163 16313 5215 16365
rect 5227 16313 5279 16365
rect 5291 16313 5343 16365
rect 5355 16313 5407 16365
rect 5419 16313 5471 16365
rect 5163 16243 5215 16295
rect 5227 16243 5279 16295
rect 5291 16243 5343 16295
rect 5355 16243 5407 16295
rect 5419 16243 5471 16295
rect 5163 16173 5215 16225
rect 5227 16173 5279 16225
rect 5291 16173 5343 16225
rect 5355 16173 5407 16225
rect 5419 16173 5471 16225
rect 7743 16313 7795 16365
rect 7807 16313 7859 16365
rect 7871 16313 7923 16365
rect 7935 16313 7987 16365
rect 7999 16313 8051 16365
rect 7743 16243 7795 16295
rect 7807 16243 7859 16295
rect 7871 16243 7923 16295
rect 7935 16243 7987 16295
rect 7999 16243 8051 16295
rect 7743 16173 7795 16225
rect 7807 16173 7859 16225
rect 7871 16173 7923 16225
rect 7935 16173 7987 16225
rect 7999 16173 8051 16225
rect 8516 16313 8568 16365
rect 8580 16313 8632 16365
rect 8644 16313 8696 16365
rect 8708 16313 8760 16365
rect 8772 16313 8824 16365
rect 8516 16243 8568 16295
rect 8580 16243 8632 16295
rect 8644 16243 8696 16295
rect 8708 16243 8760 16295
rect 8772 16243 8824 16295
rect 8516 16173 8568 16225
rect 8580 16173 8632 16225
rect 8644 16173 8696 16225
rect 8708 16173 8760 16225
rect 8772 16173 8824 16225
rect 9340 16313 9392 16365
rect 9404 16313 9456 16365
rect 9468 16313 9520 16365
rect 9532 16313 9584 16365
rect 9596 16313 9648 16365
rect 9340 16243 9392 16295
rect 9404 16243 9456 16295
rect 9468 16243 9520 16295
rect 9532 16243 9584 16295
rect 9596 16243 9648 16295
rect 9340 16173 9392 16225
rect 9404 16173 9456 16225
rect 9468 16173 9520 16225
rect 9532 16173 9584 16225
rect 9596 16173 9648 16225
rect 10323 16313 10375 16365
rect 10387 16313 10439 16365
rect 10451 16313 10503 16365
rect 10515 16313 10567 16365
rect 10579 16313 10631 16365
rect 10323 16243 10375 16295
rect 10387 16243 10439 16295
rect 10451 16243 10503 16295
rect 10515 16243 10567 16295
rect 10579 16243 10631 16295
rect 10323 16173 10375 16225
rect 10387 16173 10439 16225
rect 10451 16173 10503 16225
rect 10515 16173 10567 16225
rect 10579 16173 10631 16225
rect 11813 16313 11865 16365
rect 11877 16313 11929 16365
rect 11941 16313 11993 16365
rect 12005 16313 12057 16365
rect 12069 16313 12121 16365
rect 11813 16243 11865 16295
rect 11877 16243 11929 16295
rect 11941 16243 11993 16295
rect 12005 16243 12057 16295
rect 12069 16243 12121 16295
rect 11813 16173 11865 16225
rect 11877 16173 11929 16225
rect 11941 16173 11993 16225
rect 12005 16173 12057 16225
rect 12069 16173 12121 16225
rect 12635 16313 12687 16365
rect 12699 16313 12751 16365
rect 12763 16313 12815 16365
rect 12827 16313 12879 16365
rect 12891 16313 12943 16365
rect 12635 16243 12687 16295
rect 12699 16243 12751 16295
rect 12763 16243 12815 16295
rect 12827 16243 12879 16295
rect 12891 16243 12943 16295
rect 12635 16173 12687 16225
rect 12699 16173 12751 16225
rect 12763 16173 12815 16225
rect 12827 16173 12879 16225
rect 12891 16173 12943 16225
rect 13458 16313 13510 16365
rect 13522 16313 13574 16365
rect 13586 16313 13638 16365
rect 13650 16313 13702 16365
rect 13714 16313 13766 16365
rect 13458 16243 13510 16295
rect 13522 16243 13574 16295
rect 13586 16243 13638 16295
rect 13650 16243 13702 16295
rect 13714 16243 13766 16295
rect 13458 16173 13510 16225
rect 13522 16173 13574 16225
rect 13586 16173 13638 16225
rect 13650 16173 13702 16225
rect 13714 16173 13766 16225
rect 14287 16313 14339 16365
rect 14351 16313 14403 16365
rect 14415 16313 14467 16365
rect 14479 16313 14531 16365
rect 14543 16313 14595 16365
rect 14287 16243 14339 16295
rect 14351 16243 14403 16295
rect 14415 16243 14467 16295
rect 14479 16243 14531 16295
rect 14543 16243 14595 16295
rect 14287 16173 14339 16225
rect 14351 16173 14403 16225
rect 14415 16173 14467 16225
rect 14479 16173 14531 16225
rect 14543 16173 14595 16225
rect 15111 16313 15163 16365
rect 15175 16313 15227 16365
rect 15239 16313 15291 16365
rect 15303 16313 15355 16365
rect 15367 16313 15419 16365
rect 15111 16243 15163 16295
rect 15175 16243 15227 16295
rect 15239 16243 15291 16295
rect 15303 16243 15355 16295
rect 15367 16243 15419 16295
rect 15111 16173 15163 16225
rect 15175 16173 15227 16225
rect 15239 16173 15291 16225
rect 15303 16173 15355 16225
rect 15367 16173 15419 16225
rect 15934 16313 15986 16365
rect 15998 16313 16050 16365
rect 16062 16313 16114 16365
rect 16126 16313 16178 16365
rect 16190 16313 16242 16365
rect 15934 16243 15986 16295
rect 15998 16243 16050 16295
rect 16062 16243 16114 16295
rect 16126 16243 16178 16295
rect 16190 16243 16242 16295
rect 15934 16173 15986 16225
rect 15998 16173 16050 16225
rect 16062 16173 16114 16225
rect 16126 16173 16178 16225
rect 16190 16173 16242 16225
rect 16764 16171 16816 16212
rect 16828 16171 16880 16212
rect 16892 16171 16944 16212
rect 16956 16171 17008 16212
rect 5163 16137 5185 16155
rect 5185 16137 5215 16155
rect 5227 16137 5258 16155
rect 5258 16137 5279 16155
rect 5163 16103 5215 16137
rect 5227 16103 5279 16137
rect 5291 16137 5297 16155
rect 5297 16137 5331 16155
rect 5331 16137 5343 16155
rect 5291 16103 5343 16137
rect 5355 16137 5370 16155
rect 5370 16137 5404 16155
rect 5404 16137 5407 16155
rect 5355 16103 5407 16137
rect 5419 16137 5443 16155
rect 5443 16137 5471 16155
rect 16764 16160 16816 16171
rect 16828 16160 16880 16171
rect 16892 16160 16944 16171
rect 16956 16160 17008 16171
rect 5419 16103 5471 16137
rect 7743 16103 7795 16155
rect 7807 16103 7859 16155
rect 7871 16103 7923 16155
rect 7935 16103 7987 16155
rect 7999 16103 8051 16155
rect 8516 16103 8568 16155
rect 8580 16103 8632 16155
rect 8644 16103 8696 16155
rect 8708 16103 8760 16155
rect 8772 16103 8824 16155
rect 9340 16103 9392 16155
rect 9404 16103 9456 16155
rect 9468 16103 9520 16155
rect 9532 16103 9584 16155
rect 9596 16103 9648 16155
rect 10323 16103 10375 16155
rect 10387 16103 10439 16155
rect 10451 16103 10503 16155
rect 10515 16103 10567 16155
rect 10579 16103 10631 16155
rect 11813 16103 11865 16155
rect 11877 16103 11929 16155
rect 11941 16103 11993 16155
rect 12005 16103 12057 16155
rect 12069 16103 12121 16155
rect 12635 16103 12687 16155
rect 12699 16103 12751 16155
rect 12763 16103 12815 16155
rect 12827 16103 12879 16155
rect 12891 16103 12943 16155
rect 13458 16103 13510 16155
rect 13522 16103 13574 16155
rect 13586 16103 13638 16155
rect 13650 16103 13702 16155
rect 13714 16103 13766 16155
rect 14287 16103 14339 16155
rect 14351 16103 14403 16155
rect 14415 16103 14467 16155
rect 14479 16103 14531 16155
rect 14543 16103 14595 16155
rect 15111 16103 15163 16155
rect 15175 16103 15227 16155
rect 15239 16103 15291 16155
rect 15303 16103 15355 16155
rect 15367 16103 15419 16155
rect 15934 16103 15986 16155
rect 15998 16103 16050 16155
rect 16062 16103 16114 16155
rect 16126 16103 16178 16155
rect 16190 16103 16242 16155
rect 5163 16065 5185 16085
rect 5185 16065 5215 16085
rect 5227 16065 5258 16085
rect 5258 16065 5279 16085
rect 5163 16033 5215 16065
rect 5227 16033 5279 16065
rect 5291 16065 5297 16085
rect 5297 16065 5331 16085
rect 5331 16065 5343 16085
rect 5291 16033 5343 16065
rect 5355 16065 5370 16085
rect 5370 16065 5404 16085
rect 5404 16065 5407 16085
rect 5355 16033 5407 16065
rect 5419 16065 5443 16085
rect 5443 16065 5471 16085
rect 16764 16094 16816 16146
rect 16828 16094 16880 16146
rect 16892 16094 16944 16146
rect 16956 16094 17008 16146
rect 5419 16033 5471 16065
rect 7743 16033 7795 16085
rect 7807 16033 7859 16085
rect 7871 16033 7923 16085
rect 7935 16033 7987 16085
rect 7999 16033 8051 16085
rect 8516 16033 8568 16085
rect 8580 16033 8632 16085
rect 8644 16033 8696 16085
rect 8708 16033 8760 16085
rect 8772 16033 8824 16085
rect 9340 16033 9392 16085
rect 9404 16033 9456 16085
rect 9468 16033 9520 16085
rect 9532 16033 9584 16085
rect 9596 16033 9648 16085
rect 10323 16033 10375 16085
rect 10387 16033 10439 16085
rect 10451 16033 10503 16085
rect 10515 16033 10567 16085
rect 10579 16033 10631 16085
rect 11813 16033 11865 16085
rect 11877 16033 11929 16085
rect 11941 16033 11993 16085
rect 12005 16033 12057 16085
rect 12069 16033 12121 16085
rect 12635 16033 12687 16085
rect 12699 16033 12751 16085
rect 12763 16033 12815 16085
rect 12827 16033 12879 16085
rect 12891 16033 12943 16085
rect 13458 16033 13510 16085
rect 13522 16033 13574 16085
rect 13586 16033 13638 16085
rect 13650 16033 13702 16085
rect 13714 16033 13766 16085
rect 14287 16033 14339 16085
rect 14351 16033 14403 16085
rect 14415 16033 14467 16085
rect 14479 16033 14531 16085
rect 14543 16033 14595 16085
rect 15111 16033 15163 16085
rect 15175 16033 15227 16085
rect 15239 16033 15291 16085
rect 15303 16033 15355 16085
rect 15367 16033 15419 16085
rect 15934 16033 15986 16085
rect 15998 16033 16050 16085
rect 16062 16033 16114 16085
rect 16126 16033 16178 16085
rect 16190 16033 16242 16085
rect 16764 16027 16816 16079
rect 16828 16027 16880 16079
rect 16892 16027 16944 16079
rect 16956 16027 17008 16079
rect 5163 15993 5185 16015
rect 5185 15993 5215 16015
rect 5227 15993 5258 16015
rect 5258 15993 5279 16015
rect 5163 15963 5215 15993
rect 5227 15963 5279 15993
rect 5291 15993 5297 16015
rect 5297 15993 5331 16015
rect 5331 15993 5343 16015
rect 5291 15963 5343 15993
rect 5355 15993 5370 16015
rect 5370 15993 5404 16015
rect 5404 15993 5407 16015
rect 5355 15963 5407 15993
rect 5419 15993 5443 16015
rect 5443 15993 5471 16015
rect 5419 15963 5471 15993
rect 7743 15963 7795 16015
rect 7807 15963 7859 16015
rect 7871 15963 7923 16015
rect 7935 15963 7987 16015
rect 7999 15963 8051 16015
rect 8516 15963 8568 16015
rect 8580 15963 8632 16015
rect 8644 15963 8696 16015
rect 8708 15963 8760 16015
rect 8772 15963 8824 16015
rect 9340 15963 9392 16015
rect 9404 15963 9456 16015
rect 9468 15963 9520 16015
rect 9532 15963 9584 16015
rect 9596 15963 9648 16015
rect 10323 15963 10375 16015
rect 10387 15963 10439 16015
rect 10451 15963 10503 16015
rect 10515 15963 10567 16015
rect 10579 15963 10631 16015
rect 11813 15963 11865 16015
rect 11877 15963 11929 16015
rect 11941 15963 11993 16015
rect 12005 15963 12057 16015
rect 12069 15963 12121 16015
rect 12635 15963 12687 16015
rect 12699 15963 12751 16015
rect 12763 15963 12815 16015
rect 12827 15963 12879 16015
rect 12891 15963 12943 16015
rect 13458 15963 13510 16015
rect 13522 15963 13574 16015
rect 13586 15963 13638 16015
rect 13650 15963 13702 16015
rect 13714 15963 13766 16015
rect 14287 15963 14339 16015
rect 14351 15963 14403 16015
rect 14415 15963 14467 16015
rect 14479 15963 14531 16015
rect 14543 15963 14595 16015
rect 15111 15963 15163 16015
rect 15175 15963 15227 16015
rect 15239 15963 15291 16015
rect 15303 15963 15355 16015
rect 15367 15963 15419 16015
rect 15934 15963 15986 16015
rect 15998 15963 16050 16015
rect 16062 15963 16114 16015
rect 16126 15963 16178 16015
rect 16190 15963 16242 16015
rect 16764 15960 16816 16012
rect 16828 15960 16880 16012
rect 16892 15960 16944 16012
rect 16956 15960 17008 16012
rect 5163 15921 5185 15945
rect 5185 15921 5215 15945
rect 5227 15921 5258 15945
rect 5258 15921 5279 15945
rect 5163 15893 5215 15921
rect 5227 15893 5279 15921
rect 5291 15921 5297 15945
rect 5297 15921 5331 15945
rect 5331 15921 5343 15945
rect 5291 15893 5343 15921
rect 5355 15921 5370 15945
rect 5370 15921 5404 15945
rect 5404 15921 5407 15945
rect 5355 15893 5407 15921
rect 5419 15921 5443 15945
rect 5443 15921 5471 15945
rect 7743 15921 7795 15945
rect 7807 15921 7859 15945
rect 7871 15921 7923 15945
rect 7935 15921 7987 15945
rect 7999 15921 8051 15945
rect 8516 15921 8568 15945
rect 8580 15921 8632 15945
rect 8644 15921 8696 15945
rect 8708 15921 8760 15945
rect 8772 15921 8824 15945
rect 9340 15921 9392 15945
rect 9404 15921 9456 15945
rect 9468 15921 9520 15945
rect 9532 15921 9584 15945
rect 9596 15921 9648 15945
rect 10323 15921 10375 15945
rect 10387 15921 10439 15945
rect 10451 15921 10503 15945
rect 10515 15921 10567 15945
rect 10579 15921 10631 15945
rect 11813 15921 11865 15945
rect 11877 15921 11929 15945
rect 11941 15921 11993 15945
rect 12005 15921 12057 15945
rect 12069 15921 12121 15945
rect 12635 15921 12687 15945
rect 12699 15921 12751 15945
rect 12763 15921 12815 15945
rect 12827 15921 12879 15945
rect 12891 15921 12943 15945
rect 13458 15921 13510 15945
rect 13522 15921 13574 15945
rect 13586 15921 13638 15945
rect 13650 15921 13702 15945
rect 13714 15921 13766 15945
rect 14287 15921 14339 15945
rect 14351 15921 14403 15945
rect 14415 15921 14467 15945
rect 14479 15921 14531 15945
rect 14543 15921 14595 15945
rect 15111 15921 15163 15945
rect 15175 15921 15227 15945
rect 15239 15921 15291 15945
rect 15303 15921 15355 15945
rect 15367 15921 15419 15945
rect 15934 15921 15986 15945
rect 15998 15921 16050 15945
rect 16062 15921 16114 15945
rect 16126 15921 16178 15945
rect 16190 15921 16242 15945
rect 16764 15921 16816 15945
rect 16828 15921 16880 15945
rect 16892 15921 16944 15945
rect 16956 15921 17008 15945
rect 5419 15893 5471 15921
rect 7743 15893 7795 15921
rect 7807 15893 7859 15921
rect 7871 15893 7923 15921
rect 7935 15893 7987 15921
rect 7999 15893 8051 15921
rect 8516 15893 8568 15921
rect 8580 15893 8632 15921
rect 8644 15893 8696 15921
rect 8708 15893 8760 15921
rect 8772 15893 8824 15921
rect 9340 15893 9392 15921
rect 9404 15893 9456 15921
rect 9468 15893 9520 15921
rect 9532 15893 9584 15921
rect 9596 15893 9648 15921
rect 10323 15893 10375 15921
rect 10387 15893 10439 15921
rect 10451 15893 10503 15921
rect 10515 15893 10567 15921
rect 10579 15893 10631 15921
rect 11813 15893 11865 15921
rect 11877 15893 11929 15921
rect 11941 15893 11993 15921
rect 12005 15893 12057 15921
rect 12069 15893 12121 15921
rect 12635 15893 12687 15921
rect 12699 15893 12751 15921
rect 12763 15893 12815 15921
rect 12827 15893 12879 15921
rect 12891 15893 12943 15921
rect 13458 15893 13510 15921
rect 13522 15893 13574 15921
rect 13586 15893 13638 15921
rect 13650 15893 13702 15921
rect 13714 15893 13766 15921
rect 14287 15893 14339 15921
rect 14351 15893 14403 15921
rect 14415 15893 14467 15921
rect 14479 15893 14531 15921
rect 14543 15893 14595 15921
rect 15111 15893 15163 15921
rect 15175 15893 15227 15921
rect 15239 15893 15291 15921
rect 15303 15893 15355 15921
rect 15367 15893 15419 15921
rect 15934 15893 15986 15921
rect 15998 15893 16050 15921
rect 16062 15893 16114 15921
rect 16126 15893 16178 15921
rect 16190 15893 16242 15921
rect 16764 15893 16816 15921
rect 16828 15893 16880 15921
rect 16892 15893 16944 15921
rect 16956 15893 17008 15921
rect 15656 4379 15708 4431
rect 15720 4379 15772 4431
rect 16418 4345 16470 4397
rect 16482 4345 16534 4397
rect 15718 4201 15770 4253
rect 16333 4219 16385 4271
rect 16397 4219 16449 4271
rect 15718 4137 15770 4189
rect 16415 4121 16467 4173
rect 16415 4057 16467 4109
rect 15718 3776 15770 3828
rect 15718 3712 15770 3764
rect 16654 3776 16706 3828
rect 16654 3712 16706 3764
rect 3906 3629 3958 3681
rect 3973 3629 4025 3681
rect 4040 3629 4092 3681
rect 4107 3629 4159 3681
rect 4174 3629 4226 3681
rect 4240 3629 4292 3681
rect 4306 3629 4358 3681
rect 4372 3629 4424 3681
rect 4438 3629 4490 3681
rect 4504 3629 4556 3681
rect 4570 3629 4622 3681
rect 4636 3629 4688 3681
rect 4702 3629 4754 3681
rect 4768 3629 4820 3681
rect 4834 3629 4886 3681
rect 3906 3565 3958 3617
rect 3973 3565 4025 3617
rect 4040 3565 4092 3617
rect 4107 3565 4159 3617
rect 4174 3565 4226 3617
rect 4240 3565 4292 3617
rect 4306 3565 4358 3617
rect 4372 3565 4424 3617
rect 4438 3565 4490 3617
rect 4504 3565 4556 3617
rect 4570 3565 4622 3617
rect 4636 3565 4688 3617
rect 4702 3565 4754 3617
rect 4768 3565 4820 3617
rect 4834 3565 4886 3617
rect 5781 3630 5833 3682
rect 5847 3630 5899 3682
rect 5913 3630 5965 3682
rect 5979 3630 6031 3682
rect 6045 3630 6097 3682
rect 6111 3630 6163 3682
rect 6177 3630 6229 3682
rect 6243 3630 6295 3682
rect 6309 3630 6361 3682
rect 6375 3630 6427 3682
rect 6441 3630 6493 3682
rect 6507 3630 6559 3682
rect 6573 3630 6625 3682
rect 6639 3630 6691 3682
rect 5781 3566 5833 3618
rect 5847 3566 5899 3618
rect 5913 3566 5965 3618
rect 5979 3566 6031 3618
rect 6045 3566 6097 3618
rect 6111 3566 6163 3618
rect 6177 3566 6229 3618
rect 6243 3566 6295 3618
rect 6309 3566 6361 3618
rect 6375 3566 6427 3618
rect 6441 3566 6493 3618
rect 6507 3566 6559 3618
rect 6573 3566 6625 3618
rect 6639 3566 6691 3618
rect 7510 3630 7562 3682
rect 7577 3630 7629 3682
rect 7644 3630 7696 3682
rect 7711 3630 7763 3682
rect 7778 3630 7830 3682
rect 7845 3630 7897 3682
rect 7912 3630 7964 3682
rect 7979 3630 8031 3682
rect 8046 3630 8098 3682
rect 8113 3630 8165 3682
rect 8180 3630 8232 3682
rect 8246 3630 8298 3682
rect 8312 3630 8364 3682
rect 8378 3630 8430 3682
rect 8444 3630 8496 3682
rect 7510 3566 7562 3618
rect 7577 3566 7629 3618
rect 7644 3566 7696 3618
rect 7711 3566 7763 3618
rect 7778 3566 7830 3618
rect 7845 3566 7897 3618
rect 7912 3566 7964 3618
rect 7979 3566 8031 3618
rect 8046 3566 8098 3618
rect 8113 3566 8165 3618
rect 8180 3566 8232 3618
rect 8246 3566 8298 3618
rect 8312 3566 8364 3618
rect 8378 3566 8430 3618
rect 8444 3566 8496 3618
rect 9322 3629 9374 3681
rect 9389 3629 9441 3681
rect 9456 3629 9508 3681
rect 9523 3629 9575 3681
rect 9590 3629 9642 3681
rect 9656 3629 9708 3681
rect 9722 3629 9774 3681
rect 9788 3629 9840 3681
rect 9854 3629 9906 3681
rect 9920 3629 9972 3681
rect 9986 3629 10038 3681
rect 10052 3629 10104 3681
rect 10118 3629 10170 3681
rect 10184 3629 10236 3681
rect 10250 3629 10302 3681
rect 9322 3565 9374 3617
rect 9389 3565 9441 3617
rect 9456 3565 9508 3617
rect 9523 3565 9575 3617
rect 9590 3565 9642 3617
rect 9656 3565 9708 3617
rect 9722 3565 9774 3617
rect 9788 3565 9840 3617
rect 9854 3565 9906 3617
rect 9920 3565 9972 3617
rect 9986 3565 10038 3617
rect 10052 3565 10104 3617
rect 10118 3565 10170 3617
rect 10184 3565 10236 3617
rect 10250 3565 10302 3617
rect 11124 3629 11176 3681
rect 11191 3629 11243 3681
rect 11258 3629 11310 3681
rect 11325 3629 11377 3681
rect 11392 3629 11444 3681
rect 11458 3629 11510 3681
rect 11524 3629 11576 3681
rect 11590 3629 11642 3681
rect 11656 3629 11708 3681
rect 11722 3629 11774 3681
rect 11788 3629 11840 3681
rect 11854 3629 11906 3681
rect 11920 3629 11972 3681
rect 11986 3629 12038 3681
rect 12052 3629 12104 3681
rect 11124 3565 11176 3617
rect 11191 3565 11243 3617
rect 11258 3565 11310 3617
rect 11325 3565 11377 3617
rect 11392 3565 11444 3617
rect 11458 3565 11510 3617
rect 11524 3565 11576 3617
rect 11590 3565 11642 3617
rect 11656 3565 11708 3617
rect 11722 3565 11774 3617
rect 11788 3565 11840 3617
rect 11854 3565 11906 3617
rect 11920 3565 11972 3617
rect 11986 3565 12038 3617
rect 12052 3565 12104 3617
rect 12928 3629 12980 3681
rect 12995 3629 13047 3681
rect 13062 3629 13114 3681
rect 13129 3629 13181 3681
rect 13196 3629 13248 3681
rect 13262 3629 13314 3681
rect 13328 3629 13380 3681
rect 13394 3629 13446 3681
rect 13460 3629 13512 3681
rect 13526 3629 13578 3681
rect 13592 3629 13644 3681
rect 13658 3629 13710 3681
rect 13724 3629 13776 3681
rect 13790 3629 13842 3681
rect 13856 3629 13908 3681
rect 12928 3565 12980 3617
rect 12995 3565 13047 3617
rect 13062 3565 13114 3617
rect 13129 3565 13181 3617
rect 13196 3565 13248 3617
rect 13262 3565 13314 3617
rect 13328 3565 13380 3617
rect 13394 3565 13446 3617
rect 13460 3565 13512 3617
rect 13526 3565 13578 3617
rect 13592 3565 13644 3617
rect 13658 3565 13710 3617
rect 13724 3565 13776 3617
rect 13790 3565 13842 3617
rect 13856 3565 13908 3617
rect 14726 3629 14778 3681
rect 14792 3629 14844 3681
rect 14858 3629 14910 3681
rect 14924 3629 14976 3681
rect 14990 3629 15042 3681
rect 15055 3629 15107 3681
rect 15120 3629 15172 3681
rect 15185 3629 15237 3681
rect 15250 3629 15302 3681
rect 15315 3629 15367 3681
rect 15380 3629 15432 3681
rect 15445 3629 15497 3681
rect 15510 3629 15562 3681
rect 14726 3565 14778 3617
rect 14792 3565 14844 3617
rect 14858 3565 14910 3617
rect 14924 3565 14976 3617
rect 14990 3565 15042 3617
rect 15055 3565 15107 3617
rect 15120 3565 15172 3617
rect 15185 3565 15237 3617
rect 15250 3565 15302 3617
rect 15315 3565 15367 3617
rect 15380 3565 15432 3617
rect 15445 3565 15497 3617
rect 15510 3565 15562 3617
rect -3110 3192 -3058 3244
rect 5174 3229 5226 3281
rect 5240 3229 5292 3281
rect 5306 3229 5358 3281
rect 5372 3229 5424 3281
rect 5438 3229 5490 3281
rect 5503 3229 5555 3281
rect 5568 3229 5620 3281
rect 5633 3229 5685 3281
rect -3110 3128 -3058 3180
rect 5174 3133 5226 3185
rect 5240 3133 5292 3185
rect 5306 3133 5358 3185
rect 5372 3133 5424 3185
rect 5438 3133 5490 3185
rect 5503 3133 5555 3185
rect 5568 3133 5620 3185
rect 5633 3133 5685 3185
rect -3100 3022 -3048 3074
rect -3036 3022 -2984 3074
rect -3190 2965 -3138 3017
rect -3190 2901 -3138 2953
rect 5011 2937 5063 2989
rect 5075 2937 5127 2989
rect 5220 2745 5272 2797
rect 5286 2745 5338 2797
rect 5351 2745 5403 2797
rect 5416 2745 5468 2797
rect 5481 2745 5533 2797
rect 5546 2745 5598 2797
rect 5611 2745 5663 2797
rect 5676 2745 5728 2797
rect 5741 2745 5793 2797
rect 5806 2745 5858 2797
rect 5871 2745 5923 2797
rect 5936 2745 5988 2797
rect 5220 2651 5272 2703
rect 5286 2651 5338 2703
rect 5351 2651 5403 2703
rect 5416 2651 5468 2703
rect 5481 2651 5533 2703
rect 5546 2651 5598 2703
rect 5611 2651 5663 2703
rect 5676 2651 5728 2703
rect 5741 2651 5793 2703
rect 5806 2651 5858 2703
rect 5871 2651 5923 2703
rect 5936 2651 5988 2703
rect 8528 3229 8580 3281
rect 8594 3229 8646 3281
rect 8660 3229 8712 3281
rect 8726 3229 8778 3281
rect 8792 3229 8844 3281
rect 8857 3229 8909 3281
rect 8922 3229 8974 3281
rect 8528 3163 8580 3215
rect 8594 3163 8646 3215
rect 8660 3163 8712 3215
rect 8726 3163 8778 3215
rect 8792 3163 8844 3215
rect 8857 3163 8909 3215
rect 8922 3163 8974 3215
rect 8187 3017 8239 3069
rect 8251 3017 8303 3069
rect 7720 2937 7772 2989
rect 7784 2937 7836 2989
rect 8417 2745 8469 2797
rect 8482 2745 8534 2797
rect 8547 2745 8599 2797
rect 8612 2745 8664 2797
rect 8677 2745 8729 2797
rect 8741 2745 8793 2797
rect 8805 2745 8857 2797
rect 8417 2651 8469 2703
rect 8482 2651 8534 2703
rect 8547 2651 8599 2703
rect 8612 2651 8664 2703
rect 8677 2651 8729 2703
rect 8741 2651 8793 2703
rect 8805 2651 8857 2703
rect -3190 2212 -3138 2264
rect -3190 2148 -3138 2200
rect 7720 2228 7772 2280
rect 7784 2228 7836 2280
rect -3350 2054 -3298 2106
rect -3350 1990 -3298 2042
rect -3430 1898 -3378 1950
rect -3430 1834 -3378 1886
rect 5011 2148 5063 2200
rect 5075 2148 5127 2200
rect -2950 1716 -2898 1768
rect 934 1758 986 1767
rect 934 1724 936 1758
rect 936 1724 970 1758
rect 970 1724 986 1758
rect -2950 1652 -2898 1704
rect 934 1715 986 1724
rect 3212 1766 3264 1818
rect 3283 1766 3335 1818
rect 3354 1766 3406 1818
rect 3425 1766 3477 1818
rect 3495 1766 3547 1818
rect 3565 1766 3617 1818
rect 934 1651 986 1703
rect 1014 1623 1066 1675
rect -2864 1556 -2812 1608
rect -2800 1556 -2748 1608
rect 1014 1602 1066 1611
rect 1014 1568 1044 1602
rect 1044 1568 1066 1602
rect 1014 1559 1066 1568
<< metal2 >>
rect 2045 24427 3611 24453
rect 2045 24375 2047 24427
rect 2099 24375 2903 24427
rect 2955 24375 3611 24427
rect 2045 24363 3611 24375
rect 2045 24311 2047 24363
rect 2099 24311 2903 24363
rect 2955 24311 3611 24363
rect 2045 24299 3611 24311
rect 2045 24247 2047 24299
rect 2099 24247 2903 24299
rect 2955 24247 3611 24299
rect 2045 24235 3611 24247
rect 2045 24183 2047 24235
rect 2099 24183 2903 24235
rect 2955 24183 3611 24235
rect 2045 24171 3611 24183
rect 2045 24119 2047 24171
rect 2099 24119 2903 24171
rect 2955 24119 3611 24171
rect 2045 24113 3611 24119
rect 1302 23999 4458 24005
rect 1302 23947 1619 23999
rect 1671 23947 4458 23999
rect 1302 23935 4458 23947
rect 1302 23883 1619 23935
rect 1671 23883 4458 23935
rect 1302 23871 4458 23883
rect 1302 23819 1619 23871
rect 1671 23819 4458 23871
rect 1302 23807 4458 23819
rect 1302 23755 1619 23807
rect 1671 23755 4458 23807
rect 1302 23743 4458 23755
rect 1302 23691 1619 23743
rect 1671 23691 4458 23743
rect 1302 23679 4458 23691
rect 1302 23627 1619 23679
rect 1671 23627 4458 23679
rect 1302 23615 4458 23627
rect 1302 23563 1619 23615
rect 1671 23563 4458 23615
rect 1302 23358 4458 23563
tri 1378 23326 1410 23358 ne
tri 1776 23326 1808 23358 ne
rect 1808 23326 4458 23358
tri 1808 23268 1866 23326 ne
rect 1866 23268 4458 23326
tri 1316 23248 1336 23268 se
rect 1336 23248 1472 23268
rect 1114 23242 1166 23248
rect 1114 23178 1166 23190
tri 1086 23042 1114 23070 se
rect 1114 23056 1166 23126
rect 1114 23042 1152 23056
tri 1152 23042 1166 23056 nw
tri 1295 23227 1316 23248 se
rect 1316 23227 1472 23248
rect 1295 23216 1472 23227
rect 1524 23216 1536 23268
rect 1588 23216 1600 23268
rect 1652 23216 1664 23268
rect 1716 23216 1728 23268
rect 1780 23216 1786 23268
tri 1866 23216 1918 23268 ne
rect 1918 23216 4458 23268
tri 907 22995 954 23042 se
rect 954 22995 1105 23042
tri 1105 22995 1152 23042 nw
rect 907 22990 1100 22995
tri 1100 22990 1105 22995 nw
rect 827 22874 879 22880
rect 827 22810 879 22822
rect 827 22324 879 22758
rect 907 22324 959 22990
tri 959 22965 984 22990 nw
rect 988 22948 1040 22954
rect 988 22884 1040 22896
rect 988 22718 1040 22832
rect 988 22654 1040 22666
rect 988 22324 1040 22602
rect 1068 22828 1083 22880
rect 1135 22828 1147 22880
rect 1199 22828 1205 22880
rect 1068 22324 1120 22828
tri 1120 22803 1145 22828 nw
tri 1286 22803 1295 22812 se
rect 1295 22803 1347 23216
tri 1347 23191 1372 23216 nw
tri 1918 23191 1943 23216 ne
rect 1943 23191 4458 23216
tri 1943 23172 1962 23191 ne
tri 1221 22738 1286 22803 se
rect 1286 22790 1347 22803
rect 1286 22738 1295 22790
tri 1295 22738 1347 22790 nw
rect 1406 23107 1412 23159
rect 1464 23107 1476 23159
rect 1528 23107 1534 23159
tri 1190 22707 1221 22738 se
rect 1221 22707 1264 22738
tri 1264 22707 1295 22738 nw
tri 1153 22670 1190 22707 se
rect 1190 22670 1227 22707
tri 1227 22670 1264 22707 nw
tri 1369 22670 1406 22707 se
rect 1406 22685 1458 23107
tri 1458 23082 1483 23107 nw
rect 1406 22670 1443 22685
tri 1443 22670 1458 22685 nw
tri 1148 22665 1153 22670 se
rect 1153 22665 1222 22670
tri 1222 22665 1227 22670 nw
tri 1364 22665 1369 22670 se
rect 1369 22665 1437 22670
rect 1148 22664 1221 22665
tri 1221 22664 1222 22665 nw
tri 1363 22664 1364 22665 se
rect 1364 22664 1437 22665
tri 1437 22664 1443 22670 nw
rect 1962 22664 4458 23191
rect 1148 22324 1200 22664
tri 1200 22643 1221 22664 nw
tri 1342 22643 1363 22664 se
rect 1363 22643 1406 22664
tri 1332 22633 1342 22643 se
rect 1342 22633 1406 22643
tri 1406 22633 1437 22664 nw
tri 1311 22612 1332 22633 se
rect 1332 22612 1385 22633
tri 1385 22612 1406 22633 nw
rect 1962 22612 2163 22664
rect 2215 22612 2475 22664
rect 2527 22612 2787 22664
rect 2839 22612 4458 22664
tri 1308 22609 1311 22612 se
rect 1311 22609 1382 22612
tri 1382 22609 1385 22612 nw
rect 1308 22600 1373 22609
tri 1373 22600 1382 22609 nw
rect 1962 22600 4458 22612
rect 1228 22535 1280 22541
rect 1228 22471 1280 22483
rect 1228 22324 1280 22419
rect 1308 22443 1360 22600
tri 1360 22587 1373 22600 nw
rect 1962 22548 2163 22600
rect 2215 22548 2475 22600
rect 2527 22548 2787 22600
rect 2839 22548 4458 22600
rect 1962 22536 4458 22548
rect 1962 22484 2163 22536
rect 2215 22484 2475 22536
rect 2527 22484 2787 22536
rect 2839 22484 4458 22536
rect 1962 22458 4458 22484
tri 3198 22429 3227 22458 ne
tri 3781 22429 3810 22458 nw
tri 5002 22429 5031 22458 ne
tri 5585 22429 5614 22458 nw
tri 6800 22429 6829 22458 ne
tri 7383 22429 7412 22458 nw
tri 10156 22429 10184 22457 ne
rect 10184 22429 10191 22457
tri 10184 22422 10191 22429 ne
tri 10451 22422 10486 22457 nw
tri 10983 22422 11018 22457 ne
tri 11266 22422 11301 22457 nw
rect 1308 22379 1360 22391
rect 1308 22321 1360 22327
rect 2037 22330 4407 22350
rect 2037 22278 2047 22330
rect 2099 22278 2903 22330
rect 2955 22278 4407 22330
rect 2037 22266 4407 22278
rect 2037 22214 2047 22266
rect 2099 22214 2903 22266
rect 2955 22214 4407 22266
rect 2037 22202 4407 22214
rect 2037 22150 2047 22202
rect 2099 22150 2903 22202
rect 2955 22150 4407 22202
rect 2037 22138 4407 22150
rect 2037 22086 2047 22138
rect 2099 22086 2903 22138
rect 2955 22086 4407 22138
rect 2037 22074 4407 22086
rect 2037 22022 2047 22074
rect 2099 22022 2903 22074
rect 2955 22022 4407 22074
rect 2037 22010 4407 22022
rect 2037 21958 2047 22010
rect 2099 21958 2903 22010
rect 2955 21958 4407 22010
rect 2037 21952 4407 21958
rect 907 21732 959 21738
rect 907 21668 959 21680
rect 907 21604 959 21616
tri 1680 21574 1705 21599 nw
rect 907 21546 959 21552
rect 17254 20895 17382 20935
rect 1334 20273 1386 20279
rect 1996 20227 2002 20279
rect 2054 20227 2066 20279
rect 2118 20227 2124 20279
rect 1334 20209 1386 20221
rect 1334 20151 1386 20157
rect 1174 19965 1226 19971
rect 1174 19901 1226 19913
rect 1996 19859 2002 19911
rect 2054 19859 2066 19911
rect 2118 19859 2124 19911
rect 1174 19843 1226 19849
rect 1014 19434 1066 19440
rect 1014 19370 1066 19382
rect 1014 19312 1066 19318
rect 534 19230 586 19236
rect 534 19166 586 19178
rect 534 19108 586 19114
rect 2104 18977 2110 19029
rect 2162 18977 2174 19029
rect 2226 18977 2232 19029
rect 593 18847 746 18902
rect 645 18795 746 18847
rect 593 18783 746 18795
rect 645 18731 746 18783
rect 593 18719 746 18731
rect 645 18667 746 18719
rect 593 18655 746 18667
rect 645 18603 746 18655
rect 593 18591 746 18603
rect 645 18539 746 18591
rect 593 18508 746 18539
rect 854 18218 906 18224
rect 854 18154 906 18166
rect 854 18090 906 18102
rect 1994 18051 2000 18103
rect 2052 18051 2064 18103
rect 2116 18051 2122 18103
rect 854 18032 906 18038
rect 614 17939 666 17945
rect 614 17875 666 17887
rect 614 17817 666 17823
tri 432 16706 454 16728 se
rect 454 16706 506 17432
tri 377 16651 432 16706 se
rect 432 16694 494 16706
tri 494 16694 506 16706 nw
rect 432 16685 485 16694
tri 485 16685 494 16694 nw
tri 525 16685 534 16694 se
rect 534 16685 586 17432
rect 432 16651 451 16685
tri 451 16651 485 16685 nw
tri 512 16672 525 16685 se
rect 525 16672 586 16685
tri 491 16651 512 16672 se
rect 512 16651 565 16672
tri 565 16651 586 16672 nw
tri 605 16651 614 16660 se
rect 614 16651 666 17432
tri 355 16629 377 16651 se
rect 377 16645 445 16651
tri 445 16645 451 16651 nw
tri 485 16645 491 16651 se
rect 491 16645 559 16651
tri 559 16645 565 16651 nw
tri 599 16645 605 16651 se
rect 605 16645 666 16651
rect 377 16629 429 16645
tri 429 16629 445 16645 nw
tri 469 16629 485 16645 se
rect 485 16638 552 16645
tri 552 16638 559 16645 nw
tri 592 16638 599 16645 se
rect 599 16638 666 16645
rect 485 16629 543 16638
tri 543 16629 552 16638 nw
tri 583 16629 592 16638 se
rect 592 16629 657 16638
tri 657 16629 666 16638 nw
tri -2869 16555 -2795 16629 se
rect -2795 16611 411 16629
tri 411 16611 429 16629 nw
tri 451 16611 469 16629 se
rect 469 16611 519 16629
rect -2795 16577 377 16611
tri 377 16577 411 16611 nw
tri 417 16577 451 16611 se
rect 451 16605 519 16611
tri 519 16605 543 16629 nw
tri 559 16605 583 16629 se
rect 583 16626 654 16629
tri 654 16626 657 16629 nw
rect 583 16605 627 16626
rect 451 16577 491 16605
tri 491 16577 519 16605 nw
tri 531 16577 559 16605 se
rect 559 16599 627 16605
tri 627 16599 654 16626 nw
tri 672 16604 694 16626 se
rect 694 16604 746 17432
tri 667 16599 672 16604 se
rect 672 16599 734 16604
rect 559 16577 605 16599
tri 605 16577 627 16599 nw
tri 645 16577 667 16599 se
rect 667 16592 734 16599
tri 734 16592 746 16604 nw
rect 667 16577 719 16592
tri 719 16577 734 16592 nw
tri 759 16577 774 16592 se
rect 774 16577 826 17432
tri -2795 16555 -2773 16577 nw
tri 411 16571 417 16577 se
rect 417 16571 485 16577
tri 485 16571 491 16577 nw
tri 525 16571 531 16577 se
rect 531 16571 599 16577
tri 599 16571 605 16577 nw
tri 639 16571 645 16577 se
rect 645 16571 713 16577
tri 713 16571 719 16577 nw
tri 753 16571 759 16577 se
rect 759 16571 826 16577
tri 395 16555 411 16571 se
rect 411 16565 479 16571
tri 479 16565 485 16571 nw
tri 519 16565 525 16571 se
rect 525 16565 593 16571
tri 593 16565 599 16571 nw
tri 633 16565 639 16571 se
rect 639 16565 707 16571
tri 707 16565 713 16571 nw
tri 752 16570 753 16571 se
rect 753 16570 826 16571
tri 747 16565 752 16570 se
rect 752 16565 821 16570
tri 821 16565 826 16570 nw
rect 411 16555 469 16565
tri 469 16555 479 16565 nw
tri 509 16555 519 16565 se
rect 519 16559 587 16565
tri 587 16559 593 16565 nw
tri 627 16559 633 16565 se
rect 633 16559 701 16565
tri 701 16559 707 16565 nw
tri 741 16559 747 16565 se
rect 747 16559 815 16565
tri 815 16559 821 16565 nw
rect 519 16555 583 16559
tri 583 16555 587 16559 nw
tri 623 16555 627 16559 se
rect 627 16555 697 16559
tri 697 16555 701 16559 nw
tri 737 16555 741 16559 se
rect 741 16555 811 16559
tri 811 16555 815 16559 nw
tri 851 16555 854 16558 se
rect 854 16555 906 17432
tri -2943 16481 -2869 16555 se
rect -2869 16549 -2801 16555
tri -2801 16549 -2795 16555 nw
tri 389 16549 395 16555 se
rect 395 16549 463 16555
tri 463 16549 469 16555 nw
tri 503 16549 509 16555 se
rect 509 16549 577 16555
tri 577 16549 583 16555 nw
tri 617 16549 623 16555 se
rect 623 16553 695 16555
tri 695 16553 697 16555 nw
tri 735 16553 737 16555 se
rect 737 16553 809 16555
tri 809 16553 811 16555 nw
tri 849 16553 851 16555 se
rect 851 16553 906 16555
rect 623 16549 691 16553
tri 691 16549 695 16553 nw
tri 731 16549 735 16553 se
rect 735 16549 805 16553
tri 805 16549 809 16553 nw
tri 845 16549 849 16553 se
rect 849 16549 906 16553
rect -2869 16515 -2835 16549
tri -2835 16515 -2801 16549 nw
tri -2795 16515 -2761 16549 se
rect -2761 16531 445 16549
tri 445 16531 463 16549 nw
tri 485 16531 503 16549 se
rect 503 16531 553 16549
rect -2761 16515 411 16531
tri -2869 16481 -2835 16515 nw
tri -2829 16481 -2795 16515 se
rect -2795 16497 411 16515
tri 411 16497 445 16531 nw
tri 451 16497 485 16531 se
rect 485 16525 553 16531
tri 553 16525 577 16549 nw
tri 593 16525 617 16549 se
rect 617 16525 661 16549
rect 485 16497 525 16525
tri 525 16497 553 16525 nw
tri 565 16497 593 16525 se
rect 593 16519 661 16525
tri 661 16519 691 16549 nw
tri 701 16519 731 16549 se
rect 731 16536 792 16549
tri 792 16536 805 16549 nw
tri 832 16536 845 16549 se
rect 845 16536 906 16549
rect 731 16519 769 16536
rect 593 16497 639 16519
tri 639 16497 661 16519 nw
tri 679 16497 701 16519 se
rect 701 16513 769 16519
tri 769 16513 792 16536 nw
tri 809 16513 832 16536 se
rect 832 16524 894 16536
tri 894 16524 906 16536 nw
rect 832 16513 877 16524
rect 701 16497 753 16513
tri 753 16497 769 16513 nw
tri 793 16497 809 16513 se
rect 809 16507 877 16513
tri 877 16507 894 16524 nw
tri 917 16507 934 16524 se
rect 934 16507 986 17432
rect 809 16497 867 16507
tri 867 16497 877 16507 nw
tri 912 16502 917 16507 se
rect 917 16502 986 16507
tri 907 16497 912 16502 se
rect 912 16497 981 16502
tri 981 16497 986 16502 nw
rect -2795 16481 -2761 16497
tri -3017 16407 -2943 16481 se
rect -2943 16475 -2875 16481
tri -2875 16475 -2869 16481 nw
tri -2835 16475 -2829 16481 se
rect -2829 16475 -2761 16481
tri -2761 16475 -2739 16497 nw
tri 445 16491 451 16497 se
rect 451 16491 519 16497
tri 519 16491 525 16497 nw
tri 559 16491 565 16497 se
rect 565 16491 633 16497
tri 633 16491 639 16497 nw
tri 673 16491 679 16497 se
rect 679 16491 747 16497
tri 747 16491 753 16497 nw
tri 787 16491 793 16497 se
rect 793 16491 861 16497
tri 861 16491 867 16497 nw
tri 901 16491 907 16497 se
rect 907 16491 975 16497
tri 975 16491 981 16497 nw
tri 429 16475 445 16491 se
rect 445 16485 513 16491
tri 513 16485 519 16491 nw
tri 553 16485 559 16491 se
rect 559 16485 627 16491
tri 627 16485 633 16491 nw
tri 667 16485 673 16491 se
rect 673 16485 741 16491
tri 741 16485 747 16491 nw
tri 781 16485 787 16491 se
rect 787 16485 855 16491
tri 855 16485 861 16491 nw
tri 895 16485 901 16491 se
rect 901 16485 969 16491
tri 969 16485 975 16491 nw
tri 1009 16485 1014 16490 se
rect 1014 16485 1066 17432
rect 445 16475 503 16485
tri 503 16475 513 16485 nw
tri 543 16475 553 16485 se
rect 553 16479 621 16485
tri 621 16479 627 16485 nw
tri 661 16479 667 16485 se
rect 667 16479 735 16485
tri 735 16479 741 16485 nw
tri 775 16479 781 16485 se
rect 781 16479 849 16485
tri 849 16479 855 16485 nw
tri 889 16479 895 16485 se
rect 895 16479 963 16485
tri 963 16479 969 16485 nw
tri 1003 16479 1009 16485 se
rect 1009 16479 1066 16485
rect 553 16475 617 16479
tri 617 16475 621 16479 nw
tri 657 16475 661 16479 se
rect 661 16475 731 16479
tri 731 16475 735 16479 nw
tri 771 16475 775 16479 se
rect 775 16475 845 16479
tri 845 16475 849 16479 nw
tri 885 16475 889 16479 se
rect 889 16475 959 16479
tri 959 16475 963 16479 nw
tri 999 16475 1003 16479 se
rect 1003 16475 1066 16479
rect -2943 16441 -2909 16475
tri -2909 16441 -2875 16475 nw
tri -2869 16441 -2835 16475 se
rect -2835 16469 -2767 16475
tri -2767 16469 -2761 16475 nw
tri 423 16469 429 16475 se
rect 429 16469 497 16475
tri 497 16469 503 16475 nw
tri 537 16469 543 16475 se
rect 543 16469 611 16475
tri 611 16469 617 16475 nw
tri 651 16469 657 16475 se
rect 657 16473 729 16475
tri 729 16473 731 16475 nw
tri 769 16473 771 16475 se
rect 771 16473 843 16475
tri 843 16473 845 16475 nw
tri 883 16473 885 16475 se
rect 885 16473 957 16475
tri 957 16473 959 16475 nw
tri 997 16473 999 16475 se
rect 999 16473 1066 16475
rect 657 16469 725 16473
tri 725 16469 729 16473 nw
tri 765 16469 769 16473 se
rect 769 16469 839 16473
tri 839 16469 843 16473 nw
tri 879 16469 883 16473 se
rect 883 16469 953 16473
tri 953 16469 957 16473 nw
tri 993 16469 997 16473 se
rect 997 16469 1066 16473
rect -2835 16441 -2801 16469
tri -2943 16407 -2909 16441 nw
tri -2903 16407 -2869 16441 se
rect -2869 16435 -2801 16441
tri -2801 16435 -2767 16469 nw
tri -2761 16435 -2727 16469 se
rect -2727 16451 479 16469
tri 479 16451 497 16469 nw
tri 519 16451 537 16469 se
rect 537 16451 587 16469
rect -2727 16435 445 16451
rect -2869 16407 -2835 16435
tri -3053 16371 -3017 16407 se
rect -3017 16401 -2949 16407
tri -2949 16401 -2943 16407 nw
tri -2909 16401 -2903 16407 se
rect -2903 16401 -2835 16407
tri -2835 16401 -2801 16435 nw
tri -2795 16401 -2761 16435 se
rect -2761 16417 445 16435
tri 445 16417 479 16451 nw
tri 485 16417 519 16451 se
rect 519 16445 587 16451
tri 587 16445 611 16469 nw
tri 627 16445 651 16469 se
rect 651 16445 695 16469
rect 519 16417 559 16445
tri 559 16417 587 16445 nw
tri 599 16417 627 16445 se
rect 627 16439 695 16445
tri 695 16439 725 16469 nw
tri 735 16439 765 16469 se
rect 765 16467 837 16469
tri 837 16467 839 16469 nw
tri 877 16467 879 16469 se
rect 879 16467 951 16469
tri 951 16467 953 16469 nw
tri 992 16468 993 16469 se
rect 993 16468 1066 16469
tri 991 16467 992 16468 se
rect 992 16467 1065 16468
tri 1065 16467 1066 16468 nw
rect 765 16439 803 16467
rect 627 16417 673 16439
tri 673 16417 695 16439 nw
tri 713 16417 735 16439 se
rect 735 16433 803 16439
tri 803 16433 837 16467 nw
tri 843 16433 877 16467 se
rect 877 16461 945 16467
tri 945 16461 951 16467 nw
tri 985 16461 991 16467 se
rect 991 16461 1059 16467
tri 1059 16461 1065 16467 nw
rect 877 16433 911 16461
rect 735 16417 787 16433
tri 787 16417 803 16433 nw
tri 827 16417 843 16433 se
rect 843 16427 911 16433
tri 911 16427 945 16461 nw
tri 951 16427 985 16461 se
rect 985 16434 1032 16461
tri 1032 16434 1059 16461 nw
tri 1072 16434 1094 16456 se
rect 1094 16434 1146 17432
rect 985 16427 1019 16434
rect 843 16417 901 16427
tri 901 16417 911 16427 nw
tri 941 16417 951 16427 se
rect 951 16421 1019 16427
tri 1019 16421 1032 16434 nw
tri 1059 16421 1072 16434 se
rect 1072 16422 1134 16434
tri 1134 16422 1146 16434 nw
rect 1072 16421 1129 16422
rect 951 16417 1015 16421
tri 1015 16417 1019 16421 nw
tri 1055 16417 1059 16421 se
rect 1059 16417 1129 16421
tri 1129 16417 1134 16422 nw
tri 1169 16417 1174 16422 se
rect 1174 16417 1226 17432
rect -2761 16401 -2727 16417
rect -3017 16371 -2979 16401
tri -2979 16371 -2949 16401 nw
tri -2939 16371 -2909 16401 se
rect -2909 16395 -2841 16401
tri -2841 16395 -2835 16401 nw
tri -2801 16395 -2795 16401 se
rect -2795 16395 -2727 16401
tri -2727 16395 -2705 16417 nw
tri 479 16411 485 16417 se
rect 485 16411 553 16417
tri 553 16411 559 16417 nw
tri 593 16411 599 16417 se
rect 599 16411 667 16417
tri 667 16411 673 16417 nw
tri 707 16411 713 16417 se
rect 713 16411 781 16417
tri 781 16411 787 16417 nw
tri 821 16411 827 16417 se
rect 827 16411 895 16417
tri 895 16411 901 16417 nw
tri 935 16411 941 16417 se
rect 941 16411 1009 16417
tri 1009 16411 1015 16417 nw
tri 1049 16411 1055 16417 se
rect 1055 16415 1127 16417
tri 1127 16415 1129 16417 nw
tri 1167 16415 1169 16417 se
rect 1169 16415 1226 16417
rect 1055 16411 1123 16415
tri 1123 16411 1127 16415 nw
tri 1163 16411 1167 16415 se
rect 1167 16411 1226 16415
tri 463 16395 479 16411 se
rect 479 16405 547 16411
tri 547 16405 553 16411 nw
tri 587 16405 593 16411 se
rect 593 16405 661 16411
tri 661 16405 667 16411 nw
tri 701 16405 707 16411 se
rect 707 16405 775 16411
tri 775 16405 781 16411 nw
tri 815 16405 821 16411 se
rect 821 16405 889 16411
tri 889 16405 895 16411 nw
tri 929 16405 935 16411 se
rect 935 16405 1003 16411
tri 1003 16405 1009 16411 nw
tri 1043 16405 1049 16411 se
rect 1049 16405 1117 16411
tri 1117 16405 1123 16411 nw
tri 1157 16405 1163 16411 se
rect 1163 16405 1226 16411
rect 479 16395 537 16405
tri 537 16395 547 16405 nw
tri 577 16395 587 16405 se
rect 587 16399 655 16405
tri 655 16399 661 16405 nw
tri 695 16399 701 16405 se
rect 701 16399 769 16405
tri 769 16399 775 16405 nw
tri 809 16399 815 16405 se
rect 815 16399 883 16405
tri 883 16399 889 16405 nw
tri 923 16399 929 16405 se
rect 929 16399 997 16405
tri 997 16399 1003 16405 nw
tri 1037 16399 1043 16405 se
rect 1043 16399 1111 16405
tri 1111 16399 1117 16405 nw
tri 1152 16400 1157 16405 se
rect 1157 16400 1226 16405
tri 1151 16399 1152 16400 se
rect 1152 16399 1225 16400
tri 1225 16399 1226 16400 nw
rect 587 16395 651 16399
tri 651 16395 655 16399 nw
tri 691 16395 695 16399 se
rect 695 16395 765 16399
tri 765 16395 769 16399 nw
tri 805 16395 809 16399 se
rect 809 16395 879 16399
tri 879 16395 883 16399 nw
tri 919 16395 923 16399 se
rect 923 16395 993 16399
tri 993 16395 997 16399 nw
tri 1033 16395 1037 16399 se
rect 1037 16395 1107 16399
tri 1107 16395 1111 16399 nw
tri 1147 16395 1151 16399 se
rect 1151 16395 1221 16399
tri 1221 16395 1225 16399 nw
rect -2909 16371 -2865 16395
tri -2865 16371 -2841 16395 nw
tri -2825 16371 -2801 16395 se
rect -2801 16389 -2733 16395
tri -2733 16389 -2727 16395 nw
tri 457 16389 463 16395 se
rect 463 16389 531 16395
tri 531 16389 537 16395 nw
tri 571 16389 577 16395 se
rect 577 16389 645 16395
tri 645 16389 651 16395 nw
tri 685 16389 691 16395 se
rect 691 16393 763 16395
tri 763 16393 765 16395 nw
tri 803 16393 805 16395 se
rect 805 16393 877 16395
tri 877 16393 879 16395 nw
tri 917 16393 919 16395 se
rect 919 16393 991 16395
tri 991 16393 993 16395 nw
tri 1031 16393 1033 16395 se
rect 1033 16393 1105 16395
tri 1105 16393 1107 16395 nw
tri 1145 16393 1147 16395 se
rect 1147 16393 1219 16395
tri 1219 16393 1221 16395 nw
rect 691 16389 759 16393
tri 759 16389 763 16393 nw
tri 799 16389 803 16393 se
rect 803 16389 873 16393
tri 873 16389 877 16393 nw
tri 913 16389 917 16393 se
rect 917 16389 987 16393
tri 987 16389 991 16393 nw
tri 1027 16389 1031 16393 se
rect 1031 16389 1101 16393
tri 1101 16389 1105 16393 nw
tri 1141 16389 1145 16393 se
rect 1145 16389 1215 16393
tri 1215 16389 1219 16393 nw
rect -2801 16371 -2751 16389
tri -2751 16371 -2733 16389 nw
tri -2711 16371 -2693 16389 se
rect -2693 16371 513 16389
tri 513 16371 531 16389 nw
tri 553 16371 571 16389 se
rect 571 16371 627 16389
tri 627 16371 645 16389 nw
tri 667 16371 685 16389 se
rect 685 16371 741 16389
tri 741 16371 759 16389 nw
tri 781 16371 799 16389 se
rect 799 16387 871 16389
tri 871 16387 873 16389 nw
tri 911 16387 913 16389 se
rect 913 16387 985 16389
tri 985 16387 987 16389 nw
tri 1025 16387 1027 16389 se
rect 1027 16387 1099 16389
tri 1099 16387 1101 16389 nw
tri 1139 16387 1141 16389 se
rect 1141 16387 1213 16389
tri 1213 16387 1215 16389 nw
tri 1253 16387 1254 16388 se
rect 1254 16387 1306 17432
rect 799 16371 855 16387
tri 855 16371 871 16387 nw
tri 895 16371 911 16387 se
rect 911 16381 979 16387
tri 979 16381 985 16387 nw
tri 1019 16381 1025 16387 se
rect 1025 16381 1093 16387
tri 1093 16381 1099 16387 nw
tri 1133 16381 1139 16387 se
rect 1139 16381 1207 16387
tri 1207 16381 1213 16387 nw
tri 1247 16381 1253 16387 se
rect 1253 16381 1306 16387
rect 911 16371 969 16381
tri 969 16371 979 16381 nw
tri 1009 16371 1019 16381 se
rect 1019 16375 1087 16381
tri 1087 16375 1093 16381 nw
tri 1127 16375 1133 16381 se
rect 1133 16375 1201 16381
tri 1201 16375 1207 16381 nw
tri 1241 16375 1247 16381 se
rect 1247 16375 1306 16381
rect 1019 16371 1083 16375
tri 1083 16371 1087 16375 nw
tri 1123 16371 1127 16375 se
rect 1127 16371 1197 16375
tri 1197 16371 1201 16375 nw
tri 1237 16371 1241 16375 se
rect 1241 16371 1306 16375
tri -3059 16365 -3053 16371 se
rect -3053 16367 -2983 16371
tri -2983 16367 -2979 16371 nw
tri -2943 16367 -2939 16371 se
rect -2939 16367 -2871 16371
rect -3053 16365 -2985 16367
tri -2985 16365 -2983 16367 nw
tri -2945 16365 -2943 16367 se
rect -2943 16365 -2871 16367
tri -2871 16365 -2865 16371 nw
tri -2831 16365 -2825 16371 se
rect -2825 16365 -2757 16371
tri -2757 16365 -2751 16371 nw
tri -2717 16365 -2711 16371 se
rect -2711 16365 507 16371
tri 507 16365 513 16371 nw
tri 547 16365 553 16371 se
rect 553 16365 621 16371
tri 621 16365 627 16371 nw
tri 661 16365 667 16371 se
rect 667 16365 735 16371
tri 735 16365 741 16371 nw
tri 775 16365 781 16371 se
rect 781 16365 849 16371
tri 849 16365 855 16371 nw
tri 889 16365 895 16371 se
rect 895 16365 963 16371
tri 963 16365 969 16371 nw
tri 1003 16365 1009 16371 se
rect 1009 16365 1077 16371
tri 1077 16365 1083 16371 nw
tri 1117 16365 1123 16371 se
rect 1123 16366 1192 16371
tri 1192 16366 1197 16371 nw
tri 1232 16366 1237 16371 se
rect 1237 16366 1306 16371
rect 1123 16365 1191 16366
tri 1191 16365 1192 16366 nw
tri 1231 16365 1232 16366 se
rect 1232 16365 1305 16366
tri 1305 16365 1306 16366 nw
tri -3091 16333 -3059 16365 se
rect -3059 16333 -3017 16365
tri -3017 16333 -2985 16365 nw
tri -2977 16333 -2945 16365 se
rect -2945 16361 -2875 16365
tri -2875 16361 -2871 16365 nw
tri -2835 16361 -2831 16365 se
rect -2831 16361 -2767 16365
rect -2945 16333 -2909 16361
tri -3111 16313 -3091 16333 se
rect -3091 16327 -3023 16333
tri -3023 16327 -3017 16333 nw
tri -2983 16327 -2977 16333 se
rect -2977 16327 -2909 16333
tri -2909 16327 -2875 16361 nw
tri -2869 16327 -2835 16361 se
rect -2835 16355 -2767 16361
tri -2767 16355 -2757 16365 nw
tri -2727 16355 -2717 16365 se
rect -2717 16355 479 16365
rect -2835 16327 -2801 16355
rect -3091 16313 -3037 16327
tri -3037 16313 -3023 16327 nw
tri -2997 16313 -2983 16327 se
rect -2983 16321 -2915 16327
tri -2915 16321 -2909 16327 nw
tri -2875 16321 -2869 16327 se
rect -2869 16321 -2801 16327
tri -2801 16321 -2767 16355 nw
tri -2761 16321 -2727 16355 se
rect -2727 16337 479 16355
tri 479 16337 507 16365 nw
tri 519 16337 547 16365 se
rect 547 16337 593 16365
tri 593 16337 621 16365 nw
tri 633 16337 661 16365 se
rect 661 16359 729 16365
tri 729 16359 735 16365 nw
tri 769 16359 775 16365 se
rect 775 16359 837 16365
rect 661 16337 707 16359
tri 707 16337 729 16359 nw
tri 747 16337 769 16359 se
rect 769 16353 837 16359
tri 837 16353 849 16365 nw
tri 877 16353 889 16365 se
rect 889 16353 945 16365
rect 769 16337 821 16353
tri 821 16337 837 16353 nw
tri 861 16337 877 16353 se
rect 877 16347 945 16353
tri 945 16347 963 16365 nw
tri 985 16347 1003 16365 se
rect 1003 16347 1053 16365
rect 877 16337 935 16347
tri 935 16337 945 16347 nw
tri 975 16337 985 16347 se
rect 985 16341 1053 16347
tri 1053 16341 1077 16365 nw
tri 1093 16341 1117 16365 se
rect 1117 16341 1163 16365
rect 985 16337 1049 16341
tri 1049 16337 1053 16341 nw
tri 1089 16337 1093 16341 se
rect 1093 16337 1163 16341
tri 1163 16337 1191 16365 nw
tri 1203 16337 1231 16365 se
rect 1231 16354 1294 16365
tri 1294 16354 1305 16365 nw
rect 1231 16337 1277 16354
tri 1277 16337 1294 16354 nw
tri 1317 16337 1334 16354 se
rect 1334 16337 1386 17432
rect 1994 17098 2000 17214
rect 2116 17098 2122 17214
tri 8364 16498 8506 16640 se
rect 8506 16498 8834 20546
tri 8834 16498 8976 16640 sw
tri 9188 16498 9330 16640 se
rect 9330 16498 9658 20546
tri 9658 16498 9800 16640 sw
tri 11660 16498 11802 16640 se
rect 11802 16498 12130 20546
tri 12130 16498 12272 16640 sw
tri 12484 16498 12626 16640 se
rect 12626 16498 12954 20546
tri 12954 16498 13096 16640 sw
tri 13308 16498 13450 16640 se
rect 13450 16498 13778 20546
tri 13778 16498 13920 16640 sw
tri 14132 16498 14274 16640 se
rect 14274 16498 14602 20546
tri 14602 16498 14744 16640 sw
tri 14956 16498 15098 16640 se
rect 15098 16498 15426 20546
rect 15922 19548 16250 20546
rect 16746 20011 17074 20546
tri 17560 20154 17561 20155 se
rect 17561 20154 17871 20586
rect 17927 20546 18667 20586
tri 17074 20011 17217 20154 sw
tri 17417 20011 17560 20154 se
rect 17560 20035 17871 20154
rect 17560 20011 17847 20035
tri 17847 20011 17871 20035 nw
tri 15922 19516 15954 19548 ne
rect 15954 19516 16250 19548
tri 16250 19516 16417 19683 sw
tri 15954 19381 16089 19516 ne
tri 15922 17541 16089 17708 se
rect 16089 17572 16417 19516
rect 16089 17541 16386 17572
tri 16386 17541 16417 17572 nw
tri 15426 16498 15568 16640 sw
tri 15780 16498 15922 16640 se
rect 15922 16498 16250 17541
tri 16250 17405 16386 17541 nw
tri 16250 16498 16392 16640 sw
tri 16604 16498 16746 16640 se
rect 16746 16498 17254 20011
tri 17254 19418 17847 20011 nw
tri 3737 16458 3777 16498 se
rect 3777 16458 17254 16498
rect -2727 16321 -2693 16337
rect -2983 16313 -2923 16321
tri -2923 16313 -2915 16321 nw
tri -2883 16313 -2875 16321 se
rect -2875 16315 -2807 16321
tri -2807 16315 -2801 16321 nw
tri -2767 16315 -2761 16321 se
rect -2761 16315 -2693 16321
tri -2693 16315 -2671 16337 nw
tri 513 16331 519 16337 se
rect 519 16331 587 16337
tri 587 16331 593 16337 nw
tri 627 16331 633 16337 se
rect 633 16331 701 16337
tri 701 16331 707 16337 nw
tri 741 16331 747 16337 se
rect 747 16331 815 16337
tri 815 16331 821 16337 nw
tri 855 16331 861 16337 se
rect 861 16331 929 16337
tri 929 16331 935 16337 nw
tri 969 16331 975 16337 se
rect 975 16331 1043 16337
tri 1043 16331 1049 16337 nw
tri 1083 16331 1089 16337 se
rect 1089 16335 1161 16337
tri 1161 16335 1163 16337 nw
tri 1201 16335 1203 16337 se
rect 1203 16335 1271 16337
rect 1089 16331 1157 16335
tri 1157 16331 1161 16335 nw
tri 1197 16331 1201 16335 se
rect 1201 16331 1271 16335
tri 1271 16331 1277 16337 nw
tri 1312 16332 1317 16337 se
rect 1317 16332 1386 16337
tri 1311 16331 1312 16332 se
rect 1312 16331 1385 16332
tri 1385 16331 1386 16332 nw
rect 2002 16411 2042 16458
tri 2042 16411 2089 16458 sw
tri 3690 16411 3737 16458 se
rect 3737 16411 17079 16458
rect 2002 16378 2594 16411
tri 2594 16378 2627 16411 sw
tri 3657 16378 3690 16411 se
rect 3690 16378 17079 16411
rect 2002 16365 17079 16378
tri 497 16315 513 16331 se
rect 513 16325 581 16331
tri 581 16325 587 16331 nw
tri 621 16325 627 16331 se
rect 627 16325 695 16331
tri 695 16325 701 16331 nw
tri 735 16325 741 16331 se
rect 741 16325 809 16331
tri 809 16325 815 16331 nw
tri 849 16325 855 16331 se
rect 855 16325 923 16331
tri 923 16325 929 16331 nw
tri 963 16325 969 16331 se
rect 969 16325 1037 16331
tri 1037 16325 1043 16331 nw
tri 1077 16325 1083 16331 se
rect 1083 16325 1151 16331
tri 1151 16325 1157 16331 nw
tri 1191 16325 1197 16331 se
rect 1197 16329 1269 16331
tri 1269 16329 1271 16331 nw
tri 1309 16329 1311 16331 se
rect 1311 16329 1379 16331
rect 1197 16325 1265 16329
tri 1265 16325 1269 16329 nw
tri 1305 16325 1309 16329 se
rect 1309 16325 1379 16329
tri 1379 16325 1385 16331 nw
rect 513 16315 571 16325
tri 571 16315 581 16325 nw
tri 611 16315 621 16325 se
rect 621 16319 689 16325
tri 689 16319 695 16325 nw
tri 729 16319 735 16325 se
rect 735 16319 803 16325
tri 803 16319 809 16325 nw
tri 843 16319 849 16325 se
rect 849 16319 917 16325
tri 917 16319 923 16325 nw
tri 957 16319 963 16325 se
rect 963 16319 1031 16325
tri 1031 16319 1037 16325 nw
tri 1071 16319 1077 16325 se
rect 1077 16319 1145 16325
tri 1145 16319 1151 16325 nw
tri 1185 16319 1191 16325 se
rect 1191 16319 1259 16325
tri 1259 16319 1265 16325 nw
tri 1299 16319 1305 16325 se
rect 1305 16319 1373 16325
tri 1373 16319 1379 16325 nw
rect 621 16315 685 16319
tri 685 16315 689 16319 nw
tri 725 16315 729 16319 se
rect 729 16315 799 16319
tri 799 16315 803 16319 nw
tri 839 16315 843 16319 se
rect 843 16315 913 16319
tri 913 16315 917 16319 nw
tri 953 16315 957 16319 se
rect 957 16315 1027 16319
tri 1027 16315 1031 16319 nw
tri 1067 16315 1071 16319 se
rect 1071 16315 1141 16319
tri 1141 16315 1145 16319 nw
tri 1181 16315 1185 16319 se
rect 1185 16315 1255 16319
tri 1255 16315 1259 16319 nw
tri 1295 16315 1299 16319 se
rect 1299 16315 1369 16319
tri 1369 16315 1373 16319 nw
rect -2875 16313 -2809 16315
tri -2809 16313 -2807 16315 nw
tri -2769 16313 -2767 16315 se
rect -2767 16313 -2695 16315
tri -2695 16313 -2693 16315 nw
tri 495 16313 497 16315 se
rect 497 16313 569 16315
tri 569 16313 571 16315 nw
tri 609 16313 611 16315 se
rect 611 16313 683 16315
tri 683 16313 685 16315 nw
tri 723 16313 725 16315 se
rect 725 16313 797 16315
tri 797 16313 799 16315 nw
tri 837 16313 839 16315 se
rect 839 16313 911 16315
tri 911 16313 913 16315 nw
tri 951 16313 953 16315 se
rect 953 16313 1025 16315
tri 1025 16313 1027 16315 nw
tri 1065 16313 1067 16315 se
rect 1067 16313 1139 16315
tri 1139 16313 1141 16315 nw
tri 1179 16313 1181 16315 se
rect 1181 16313 1253 16315
tri 1253 16313 1255 16315 nw
tri 1293 16313 1295 16315 se
rect 1295 16313 1367 16315
tri 1367 16313 1369 16315 nw
rect 2002 16313 5163 16365
rect 5215 16313 5227 16365
rect 5279 16313 5291 16365
rect 5343 16313 5355 16365
rect 5407 16313 5419 16365
rect 5471 16313 7743 16365
rect 7795 16313 7807 16365
rect 7859 16313 7871 16365
rect 7923 16313 7935 16365
rect 7987 16313 7999 16365
rect 8051 16313 8516 16365
rect 8568 16313 8580 16365
rect 8632 16313 8644 16365
rect 8696 16313 8708 16365
rect 8760 16313 8772 16365
rect 8824 16313 9340 16365
rect 9392 16313 9404 16365
rect 9456 16313 9468 16365
rect 9520 16313 9532 16365
rect 9584 16313 9596 16365
rect 9648 16313 10323 16365
rect 10375 16313 10387 16365
rect 10439 16313 10451 16365
rect 10503 16313 10515 16365
rect 10567 16313 10579 16365
rect 10631 16313 11813 16365
rect 11865 16313 11877 16365
rect 11929 16313 11941 16365
rect 11993 16313 12005 16365
rect 12057 16313 12069 16365
rect 12121 16313 12635 16365
rect 12687 16313 12699 16365
rect 12751 16313 12763 16365
rect 12815 16313 12827 16365
rect 12879 16313 12891 16365
rect 12943 16313 13458 16365
rect 13510 16313 13522 16365
rect 13574 16313 13586 16365
rect 13638 16313 13650 16365
rect 13702 16313 13714 16365
rect 13766 16313 14287 16365
rect 14339 16313 14351 16365
rect 14403 16313 14415 16365
rect 14467 16313 14479 16365
rect 14531 16313 14543 16365
rect 14595 16313 15111 16365
rect 15163 16313 15175 16365
rect 15227 16313 15239 16365
rect 15291 16313 15303 16365
rect 15355 16313 15367 16365
rect 15419 16313 15934 16365
rect 15986 16313 15998 16365
rect 16050 16313 16062 16365
rect 16114 16313 16126 16365
rect 16178 16313 16190 16365
rect 16242 16313 17079 16365
tri -3115 16309 -3111 16313 se
rect -3111 16309 -3041 16313
tri -3041 16309 -3037 16313 nw
tri -3001 16309 -2997 16313 se
rect -2997 16309 -2927 16313
tri -2927 16309 -2923 16313 nw
tri -2887 16309 -2883 16313 se
rect -2883 16309 -2813 16313
tri -2813 16309 -2809 16313 nw
tri -2773 16309 -2769 16313 se
rect -2769 16309 -2699 16313
tri -2699 16309 -2695 16313 nw
tri 491 16309 495 16313 se
rect 495 16309 565 16313
tri 565 16309 569 16313 nw
tri 605 16309 609 16313 se
rect 609 16309 679 16313
tri 679 16309 683 16313 nw
tri 719 16309 723 16313 se
rect 723 16309 793 16313
tri 793 16309 797 16313 nw
tri 833 16309 837 16313 se
rect 837 16309 907 16313
tri 907 16309 911 16313 nw
tri 947 16309 951 16313 se
rect 951 16309 1021 16313
tri 1021 16309 1025 16313 nw
tri 1061 16309 1065 16313 se
rect 1065 16309 1135 16313
tri 1135 16309 1139 16313 nw
tri 1175 16309 1179 16313 se
rect 1179 16309 1249 16313
tri 1249 16309 1253 16313 nw
tri 1289 16309 1293 16313 se
rect 1293 16309 1363 16313
tri 1363 16309 1367 16313 nw
tri -3129 16295 -3115 16309 se
rect -3115 16295 -3055 16309
tri -3055 16295 -3041 16309 nw
tri -3015 16295 -3001 16309 se
rect -3001 16295 -2941 16309
tri -2941 16295 -2927 16309 nw
tri -2901 16295 -2887 16309 se
rect -2887 16295 -2827 16309
tri -2827 16295 -2813 16309 nw
tri -2787 16295 -2773 16309 se
rect -2773 16295 -2713 16309
tri -2713 16295 -2699 16309 nw
tri -2673 16295 -2659 16309 se
rect -2659 16295 551 16309
tri 551 16295 565 16309 nw
tri 591 16295 605 16309 se
rect 605 16295 665 16309
tri 665 16295 679 16309 nw
tri 705 16295 719 16309 se
rect 719 16295 779 16309
tri 779 16295 793 16309 nw
tri 819 16295 833 16309 se
rect 833 16307 905 16309
tri 905 16307 907 16309 nw
tri 945 16307 947 16309 se
rect 947 16307 1019 16309
tri 1019 16307 1021 16309 nw
tri 1059 16307 1061 16309 se
rect 1061 16307 1133 16309
tri 1133 16307 1135 16309 nw
tri 1173 16307 1175 16309 se
rect 1175 16307 1247 16309
tri 1247 16307 1249 16309 nw
tri 1287 16307 1289 16309 se
rect 1289 16307 1361 16309
tri 1361 16307 1363 16309 nw
rect 833 16295 893 16307
tri 893 16295 905 16307 nw
tri 933 16295 945 16307 se
rect 945 16301 1013 16307
tri 1013 16301 1019 16307 nw
tri 1053 16301 1059 16307 se
rect 1059 16301 1127 16307
tri 1127 16301 1133 16307 nw
tri 1167 16301 1173 16307 se
rect 1173 16301 1241 16307
tri 1241 16301 1247 16307 nw
tri 1281 16301 1287 16307 se
rect 1287 16301 1355 16307
tri 1355 16301 1361 16307 nw
rect 945 16295 1007 16301
tri 1007 16295 1013 16301 nw
tri 1047 16295 1053 16301 se
rect 1053 16295 1121 16301
tri 1121 16295 1127 16301 nw
tri 1161 16295 1167 16301 se
rect 1167 16295 1235 16301
tri 1235 16295 1241 16301 nw
tri 1275 16295 1281 16301 se
rect 1281 16295 1349 16301
tri 1349 16295 1355 16301 nw
rect 2002 16295 17079 16313
tri -3165 16259 -3129 16295 se
rect -3129 16293 -3057 16295
tri -3057 16293 -3055 16295 nw
tri -3017 16293 -3015 16295 se
rect -3015 16293 -2949 16295
rect -3129 16259 -3091 16293
tri -3091 16259 -3057 16293 nw
tri -3051 16259 -3017 16293 se
rect -3017 16287 -2949 16293
tri -2949 16287 -2941 16295 nw
tri -2909 16287 -2901 16295 se
rect -2901 16287 -2841 16295
rect -3017 16259 -2983 16287
tri -3181 16243 -3165 16259 se
rect -3165 16253 -3097 16259
tri -3097 16253 -3091 16259 nw
tri -3057 16253 -3051 16259 se
rect -3051 16253 -2983 16259
tri -2983 16253 -2949 16287 nw
tri -2943 16253 -2909 16287 se
rect -2909 16281 -2841 16287
tri -2841 16281 -2827 16295 nw
tri -2801 16281 -2787 16295 se
rect -2787 16281 -2733 16295
rect -2909 16253 -2875 16281
rect -3165 16243 -3107 16253
tri -3107 16243 -3097 16253 nw
tri -3067 16243 -3057 16253 se
rect -3057 16247 -2989 16253
tri -2989 16247 -2983 16253 nw
tri -2949 16247 -2943 16253 se
rect -2943 16247 -2875 16253
tri -2875 16247 -2841 16281 nw
tri -2835 16247 -2801 16281 se
rect -2801 16275 -2733 16281
tri -2733 16275 -2713 16295 nw
tri -2693 16275 -2673 16295 se
rect -2673 16291 547 16295
tri 547 16291 551 16295 nw
tri 587 16291 591 16295 se
rect 591 16291 655 16295
rect -2673 16275 513 16291
rect -2801 16247 -2765 16275
rect -3057 16243 -2993 16247
tri -2993 16243 -2989 16247 nw
tri -2953 16243 -2949 16247 se
rect -2949 16243 -2879 16247
tri -2879 16243 -2875 16247 nw
tri -2839 16243 -2835 16247 se
rect -2835 16243 -2765 16247
tri -2765 16243 -2733 16275 nw
tri -2725 16243 -2693 16275 se
rect -2693 16257 513 16275
tri 513 16257 547 16291 nw
tri 553 16257 587 16291 se
rect 587 16285 655 16291
tri 655 16285 665 16295 nw
tri 695 16285 705 16295 se
rect 705 16285 763 16295
rect 587 16257 627 16285
tri 627 16257 655 16285 nw
tri 667 16257 695 16285 se
rect 695 16279 763 16285
tri 763 16279 779 16295 nw
tri 803 16279 819 16295 se
rect 819 16279 871 16295
rect 695 16257 741 16279
tri 741 16257 763 16279 nw
tri 781 16257 803 16279 se
rect 803 16273 871 16279
tri 871 16273 893 16295 nw
tri 911 16273 933 16295 se
rect 933 16273 979 16295
rect 803 16257 855 16273
tri 855 16257 871 16273 nw
tri 895 16257 911 16273 se
rect 911 16267 979 16273
tri 979 16267 1007 16295 nw
tri 1019 16267 1047 16295 se
rect 1047 16267 1087 16295
rect 911 16257 969 16267
tri 969 16257 979 16267 nw
tri 1009 16257 1019 16267 se
rect 1019 16261 1087 16267
tri 1087 16261 1121 16295 nw
tri 1127 16261 1161 16295 se
rect 1161 16289 1229 16295
tri 1229 16289 1235 16295 nw
tri 1269 16289 1275 16295 se
rect 1275 16289 1343 16295
tri 1343 16289 1349 16295 nw
rect 1161 16261 1197 16289
rect 1019 16257 1083 16261
tri 1083 16257 1087 16261 nw
tri 1123 16257 1127 16261 se
rect 1127 16257 1197 16261
tri 1197 16257 1229 16289 nw
tri 1237 16257 1269 16289 se
rect 1269 16257 1311 16289
tri 1311 16257 1343 16289 nw
rect -2693 16243 -2651 16257
tri -2651 16243 -2637 16257 nw
tri 547 16251 553 16257 se
rect 553 16251 621 16257
tri 621 16251 627 16257 nw
tri 661 16251 667 16257 se
rect 667 16251 735 16257
tri 735 16251 741 16257 nw
tri 775 16251 781 16257 se
rect 781 16251 849 16257
tri 849 16251 855 16257 nw
tri 889 16251 895 16257 se
rect 895 16251 963 16257
tri 963 16251 969 16257 nw
tri 1003 16251 1009 16257 se
rect 1009 16251 1077 16257
tri 1077 16251 1083 16257 nw
tri 1117 16251 1123 16257 se
rect 1123 16255 1195 16257
tri 1195 16255 1197 16257 nw
tri 1235 16255 1237 16257 se
rect 1237 16255 1305 16257
rect 1123 16251 1191 16255
tri 1191 16251 1195 16255 nw
tri 1231 16251 1235 16255 se
rect 1235 16251 1305 16255
tri 1305 16251 1311 16257 nw
tri 539 16243 547 16251 se
rect 547 16245 615 16251
tri 615 16245 621 16251 nw
tri 655 16245 661 16251 se
rect 661 16245 729 16251
tri 729 16245 735 16251 nw
tri 769 16245 775 16251 se
rect 775 16245 843 16251
tri 843 16245 849 16251 nw
tri 883 16245 889 16251 se
rect 889 16245 957 16251
tri 957 16245 963 16251 nw
tri 997 16245 1003 16251 se
rect 1003 16245 1071 16251
tri 1071 16245 1077 16251 nw
tri 1111 16245 1117 16251 se
rect 1117 16245 1185 16251
tri 1185 16245 1191 16251 nw
tri 1225 16245 1231 16251 se
rect 1231 16245 1299 16251
tri 1299 16245 1305 16251 nw
rect 547 16243 613 16245
tri 613 16243 615 16245 nw
tri 653 16243 655 16245 se
rect 655 16243 727 16245
tri 727 16243 729 16245 nw
tri 767 16243 769 16245 se
rect 769 16243 841 16245
tri 841 16243 843 16245 nw
tri 881 16243 883 16245 se
rect 883 16243 955 16245
tri 955 16243 957 16245 nw
tri 995 16243 997 16245 se
rect 997 16243 1069 16245
tri 1069 16243 1071 16245 nw
tri 1109 16243 1111 16245 se
rect 1111 16243 1183 16245
tri 1183 16243 1185 16245 nw
tri 1223 16243 1225 16245 se
rect 1225 16243 1297 16245
tri 1297 16243 1299 16245 nw
rect 2002 16243 5163 16295
rect 5215 16243 5227 16295
rect 5279 16243 5291 16295
rect 5343 16243 5355 16295
rect 5407 16243 5419 16295
rect 5471 16243 7743 16295
rect 7795 16243 7807 16295
rect 7859 16243 7871 16295
rect 7923 16243 7935 16295
rect 7987 16243 7999 16295
rect 8051 16243 8516 16295
rect 8568 16243 8580 16295
rect 8632 16243 8644 16295
rect 8696 16243 8708 16295
rect 8760 16243 8772 16295
rect 8824 16243 9340 16295
rect 9392 16243 9404 16295
rect 9456 16243 9468 16295
rect 9520 16243 9532 16295
rect 9584 16243 9596 16295
rect 9648 16243 10323 16295
rect 10375 16243 10387 16295
rect 10439 16243 10451 16295
rect 10503 16243 10515 16295
rect 10567 16243 10579 16295
rect 10631 16243 11813 16295
rect 11865 16243 11877 16295
rect 11929 16243 11941 16295
rect 11993 16243 12005 16295
rect 12057 16243 12069 16295
rect 12121 16243 12635 16295
rect 12687 16243 12699 16295
rect 12751 16243 12763 16295
rect 12815 16243 12827 16295
rect 12879 16243 12891 16295
rect 12943 16243 13458 16295
rect 13510 16243 13522 16295
rect 13574 16243 13586 16295
rect 13638 16243 13650 16295
rect 13702 16243 13714 16295
rect 13766 16243 14287 16295
rect 14339 16243 14351 16295
rect 14403 16243 14415 16295
rect 14467 16243 14479 16295
rect 14531 16243 14543 16295
rect 14595 16243 15111 16295
rect 15163 16243 15175 16295
rect 15227 16243 15239 16295
rect 15291 16243 15303 16295
rect 15355 16243 15367 16295
rect 15419 16243 15934 16295
rect 15986 16243 15998 16295
rect 16050 16243 16062 16295
rect 16114 16243 16126 16295
rect 16178 16243 16190 16295
rect 16242 16243 17079 16295
tri -3189 16235 -3181 16243 se
rect -3181 16235 -3115 16243
tri -3115 16235 -3107 16243 nw
tri -3075 16235 -3067 16243 se
rect -3067 16235 -3001 16243
tri -3001 16235 -2993 16243 nw
tri -2961 16235 -2953 16243 se
rect -2953 16241 -2881 16243
tri -2881 16241 -2879 16243 nw
tri -2841 16241 -2839 16243 se
rect -2839 16241 -2767 16243
tri -2767 16241 -2765 16243 nw
tri -2727 16241 -2725 16243 se
rect -2725 16241 -2659 16243
rect -2953 16235 -2887 16241
tri -2887 16235 -2881 16241 nw
tri -2847 16235 -2841 16241 se
rect -2841 16235 -2773 16241
tri -2773 16235 -2767 16241 nw
tri -2733 16235 -2727 16241 se
rect -2727 16235 -2659 16241
tri -2659 16235 -2651 16243 nw
tri 531 16235 539 16243 se
rect 539 16235 605 16243
tri 605 16235 613 16243 nw
tri 645 16235 653 16243 se
rect 653 16239 723 16243
tri 723 16239 727 16243 nw
tri 763 16239 767 16243 se
rect 767 16239 837 16243
tri 837 16239 841 16243 nw
tri 877 16239 881 16243 se
rect 881 16239 951 16243
tri 951 16239 955 16243 nw
tri 991 16239 995 16243 se
rect 995 16239 1065 16243
tri 1065 16239 1069 16243 nw
tri 1105 16239 1109 16243 se
rect 1109 16239 1179 16243
tri 1179 16239 1183 16243 nw
tri 1219 16239 1223 16243 se
rect 1223 16239 1293 16243
tri 1293 16239 1297 16243 nw
rect 653 16235 719 16239
tri 719 16235 723 16239 nw
tri 759 16235 763 16239 se
rect 763 16235 833 16239
tri 833 16235 837 16239 nw
tri 873 16235 877 16239 se
rect 877 16235 947 16239
tri 947 16235 951 16239 nw
tri 987 16235 991 16239 se
rect 991 16235 1061 16239
tri 1061 16235 1065 16239 nw
tri 1101 16235 1105 16239 se
rect 1105 16235 1175 16239
tri 1175 16235 1179 16239 nw
tri 1215 16235 1219 16239 se
rect 1219 16235 1289 16239
tri 1289 16235 1293 16239 nw
tri -3199 16225 -3189 16235 se
rect -3189 16225 -3125 16235
tri -3125 16225 -3115 16235 nw
tri -3085 16225 -3075 16235 se
rect -3075 16225 -3011 16235
tri -3011 16225 -3001 16235 nw
tri -2971 16225 -2961 16235 se
rect -2961 16225 -2897 16235
tri -2897 16225 -2887 16235 nw
tri -2857 16225 -2847 16235 se
rect -2847 16225 -2783 16235
tri -2783 16225 -2773 16235 nw
tri -2743 16225 -2733 16235 se
rect -2733 16229 -2665 16235
tri -2665 16229 -2659 16235 nw
tri 525 16229 531 16235 se
rect 531 16229 599 16235
tri 599 16229 605 16235 nw
tri 639 16229 645 16235 se
rect 645 16229 713 16235
tri 713 16229 719 16235 nw
tri 753 16229 759 16235 se
rect 759 16233 831 16235
tri 831 16233 833 16235 nw
tri 871 16233 873 16235 se
rect 873 16233 945 16235
tri 945 16233 947 16235 nw
tri 985 16233 987 16235 se
rect 987 16233 1059 16235
tri 1059 16233 1061 16235 nw
tri 1099 16233 1101 16235 se
rect 1101 16233 1173 16235
tri 1173 16233 1175 16235 nw
tri 1213 16233 1215 16235 se
rect 1215 16233 1287 16235
tri 1287 16233 1289 16235 nw
rect 759 16229 827 16233
tri 827 16229 831 16233 nw
tri 867 16229 871 16233 se
rect 871 16229 941 16233
tri 941 16229 945 16233 nw
tri 981 16229 985 16233 se
rect 985 16229 1055 16233
tri 1055 16229 1059 16233 nw
tri 1095 16229 1099 16233 se
rect 1099 16229 1169 16233
tri 1169 16229 1173 16233 nw
tri 1209 16229 1213 16233 se
rect 1213 16229 1283 16233
tri 1283 16229 1287 16233 nw
rect -2733 16225 -2669 16229
tri -2669 16225 -2665 16229 nw
tri -2629 16225 -2625 16229 se
rect -2625 16225 595 16229
tri 595 16225 599 16229 nw
tri 635 16225 639 16229 se
rect 639 16225 709 16229
tri 709 16225 713 16229 nw
tri 749 16225 753 16229 se
rect 753 16225 823 16229
tri 823 16225 827 16229 nw
tri 863 16225 867 16229 se
rect 867 16227 939 16229
tri 939 16227 941 16229 nw
tri 979 16227 981 16229 se
rect 981 16227 1053 16229
tri 1053 16227 1055 16229 nw
tri 1093 16227 1095 16229 se
rect 1095 16227 1167 16229
tri 1167 16227 1169 16229 nw
tri 1207 16227 1209 16229 se
rect 1209 16227 1281 16229
tri 1281 16227 1283 16229 nw
rect 867 16225 937 16227
tri 937 16225 939 16227 nw
tri 977 16225 979 16227 se
rect 979 16225 1051 16227
tri 1051 16225 1053 16227 nw
tri 1091 16225 1093 16227 se
rect 1093 16225 1165 16227
tri 1165 16225 1167 16227 nw
tri 1205 16225 1207 16227 se
rect 1207 16225 1279 16227
tri 1279 16225 1281 16227 nw
rect 2002 16225 17079 16243
tri -3239 16185 -3199 16225 se
rect -3199 16219 -3131 16225
tri -3131 16219 -3125 16225 nw
tri -3091 16219 -3085 16225 se
rect -3085 16219 -3023 16225
rect -3199 16185 -3165 16219
tri -3165 16185 -3131 16219 nw
tri -3125 16185 -3091 16219 se
rect -3091 16213 -3023 16219
tri -3023 16213 -3011 16225 nw
tri -2983 16213 -2971 16225 se
rect -2971 16213 -2915 16225
rect -3091 16185 -3057 16213
tri -3251 16173 -3239 16185 se
rect -3239 16179 -3171 16185
tri -3171 16179 -3165 16185 nw
tri -3131 16179 -3125 16185 se
rect -3125 16179 -3057 16185
tri -3057 16179 -3023 16213 nw
tri -3017 16179 -2983 16213 se
rect -2983 16207 -2915 16213
tri -2915 16207 -2897 16225 nw
tri -2875 16207 -2857 16225 se
rect -2857 16207 -2807 16225
rect -2983 16179 -2949 16207
rect -3239 16173 -3177 16179
tri -3177 16173 -3171 16179 nw
tri -3137 16173 -3131 16179 se
rect -3131 16173 -3063 16179
tri -3063 16173 -3057 16179 nw
tri -3023 16173 -3017 16179 se
rect -3017 16173 -2949 16179
tri -2949 16173 -2915 16207 nw
tri -2909 16173 -2875 16207 se
rect -2875 16201 -2807 16207
tri -2807 16201 -2783 16225 nw
tri -2767 16201 -2743 16225 se
rect -2743 16201 -2699 16225
rect -2875 16173 -2835 16201
tri -2835 16173 -2807 16201 nw
tri -2795 16173 -2767 16201 se
rect -2767 16195 -2699 16201
tri -2699 16195 -2669 16225 nw
tri -2659 16195 -2629 16225 se
rect -2629 16211 581 16225
tri 581 16211 595 16225 nw
tri 621 16211 635 16225 se
rect 635 16211 689 16225
rect -2629 16195 547 16211
rect -2767 16173 -2721 16195
tri -2721 16173 -2699 16195 nw
tri -2681 16173 -2659 16195 se
rect -2659 16177 547 16195
tri 547 16177 581 16211 nw
tri 587 16177 621 16211 se
rect 621 16205 689 16211
tri 689 16205 709 16225 nw
tri 729 16205 749 16225 se
rect 749 16205 797 16225
rect 621 16177 661 16205
tri 661 16177 689 16205 nw
tri 701 16177 729 16205 se
rect 729 16199 797 16205
tri 797 16199 823 16225 nw
tri 837 16199 863 16225 se
rect 863 16199 905 16225
rect 729 16177 775 16199
tri 775 16177 797 16199 nw
tri 815 16177 837 16199 se
rect 837 16193 905 16199
tri 905 16193 937 16225 nw
tri 945 16193 977 16225 se
rect 977 16221 1047 16225
tri 1047 16221 1051 16225 nw
tri 1087 16221 1091 16225 se
rect 1091 16221 1161 16225
tri 1161 16221 1165 16225 nw
tri 1201 16221 1205 16225 se
rect 1205 16221 1275 16225
tri 1275 16221 1279 16225 nw
rect 977 16193 1013 16221
rect 837 16177 889 16193
tri 889 16177 905 16193 nw
tri 929 16177 945 16193 se
rect 945 16187 1013 16193
tri 1013 16187 1047 16221 nw
tri 1053 16187 1087 16221 se
rect 1087 16215 1155 16221
tri 1155 16215 1161 16221 nw
tri 1195 16215 1201 16221 se
rect 1201 16215 1269 16221
tri 1269 16215 1275 16221 nw
rect 1087 16187 1121 16215
rect 945 16177 1003 16187
tri 1003 16177 1013 16187 nw
tri 1043 16177 1053 16187 se
rect 1053 16181 1121 16187
tri 1121 16181 1155 16215 nw
tri 1161 16181 1195 16215 se
rect 1195 16181 1231 16215
rect 1053 16177 1117 16181
tri 1117 16177 1121 16181 nw
tri 1157 16177 1161 16181 se
rect 1161 16177 1231 16181
tri 1231 16177 1269 16215 nw
rect -2659 16173 -2607 16177
tri -2607 16173 -2603 16177 nw
tri 583 16173 587 16177 se
rect 587 16173 657 16177
tri 657 16173 661 16177 nw
tri 697 16173 701 16177 se
rect 701 16173 771 16177
tri 771 16173 775 16177 nw
tri 811 16173 815 16177 se
rect 815 16173 885 16177
tri 885 16173 889 16177 nw
tri 925 16173 929 16177 se
rect 929 16173 999 16177
tri 999 16173 1003 16177 nw
tri 1039 16173 1043 16177 se
rect 1043 16173 1113 16177
tri 1113 16173 1117 16177 nw
tri 1153 16173 1157 16177 se
rect 1157 16173 1227 16177
tri 1227 16173 1231 16177 nw
rect 2002 16173 5163 16225
rect 5215 16173 5227 16225
rect 5279 16173 5291 16225
rect 5343 16173 5355 16225
rect 5407 16173 5419 16225
rect 5471 16173 7743 16225
rect 7795 16173 7807 16225
rect 7859 16173 7871 16225
rect 7923 16173 7935 16225
rect 7987 16173 7999 16225
rect 8051 16173 8516 16225
rect 8568 16173 8580 16225
rect 8632 16173 8644 16225
rect 8696 16173 8708 16225
rect 8760 16173 8772 16225
rect 8824 16173 9340 16225
rect 9392 16173 9404 16225
rect 9456 16173 9468 16225
rect 9520 16173 9532 16225
rect 9584 16173 9596 16225
rect 9648 16173 10323 16225
rect 10375 16173 10387 16225
rect 10439 16173 10451 16225
rect 10503 16173 10515 16225
rect 10567 16173 10579 16225
rect 10631 16173 11813 16225
rect 11865 16173 11877 16225
rect 11929 16173 11941 16225
rect 11993 16173 12005 16225
rect 12057 16173 12069 16225
rect 12121 16173 12635 16225
rect 12687 16173 12699 16225
rect 12751 16173 12763 16225
rect 12815 16173 12827 16225
rect 12879 16173 12891 16225
rect 12943 16173 13458 16225
rect 13510 16173 13522 16225
rect 13574 16173 13586 16225
rect 13638 16173 13650 16225
rect 13702 16173 13714 16225
rect 13766 16173 14287 16225
rect 14339 16173 14351 16225
rect 14403 16173 14415 16225
rect 14467 16173 14479 16225
rect 14531 16173 14543 16225
rect 14595 16173 15111 16225
rect 15163 16173 15175 16225
rect 15227 16173 15239 16225
rect 15291 16173 15303 16225
rect 15355 16173 15367 16225
rect 15419 16173 15934 16225
rect 15986 16173 15998 16225
rect 16050 16173 16062 16225
rect 16114 16173 16126 16225
rect 16178 16173 16190 16225
rect 16242 16212 17079 16225
rect 16242 16173 16764 16212
tri -3263 16161 -3251 16173 se
rect -3251 16161 -3189 16173
tri -3189 16161 -3177 16173 nw
tri -3149 16161 -3137 16173 se
rect -3137 16161 -3075 16173
tri -3075 16161 -3063 16173 nw
tri -3035 16161 -3023 16173 se
rect -3023 16167 -2955 16173
tri -2955 16167 -2949 16173 nw
tri -2915 16167 -2909 16173 se
rect -2909 16167 -2841 16173
tri -2841 16167 -2835 16173 nw
tri -2801 16167 -2795 16173 se
rect -2795 16167 -2733 16173
rect -3023 16161 -2961 16167
tri -2961 16161 -2955 16167 nw
tri -2921 16161 -2915 16167 se
rect -2915 16161 -2847 16167
tri -2847 16161 -2841 16167 nw
tri -2807 16161 -2801 16167 se
rect -2801 16161 -2733 16167
tri -2733 16161 -2721 16173 nw
tri -2693 16161 -2681 16173 se
rect -2681 16161 -2620 16173
tri -3264 16160 -3263 16161 se
rect -3263 16160 -3190 16161
tri -3190 16160 -3189 16161 nw
tri -3150 16160 -3149 16161 se
rect -3149 16160 -3076 16161
tri -3076 16160 -3075 16161 nw
tri -3036 16160 -3035 16161 se
rect -3035 16160 -2962 16161
tri -2962 16160 -2961 16161 nw
tri -2922 16160 -2921 16161 se
rect -2921 16160 -2848 16161
tri -2848 16160 -2847 16161 nw
tri -2808 16160 -2807 16161 se
rect -2807 16160 -2734 16161
tri -2734 16160 -2733 16161 nw
tri -2694 16160 -2693 16161 se
rect -2693 16160 -2620 16161
tri -2620 16160 -2607 16173 nw
tri 581 16171 583 16173 se
rect 583 16171 655 16173
tri 655 16171 657 16173 nw
tri 695 16171 697 16173 se
rect 697 16171 769 16173
tri 769 16171 771 16173 nw
tri 809 16171 811 16173 se
rect 811 16171 883 16173
tri 883 16171 885 16173 nw
tri 923 16171 925 16173 se
rect 925 16171 997 16173
tri 997 16171 999 16173 nw
tri 1037 16171 1039 16173 se
rect 1039 16171 1111 16173
tri 1111 16171 1113 16173 nw
tri 1151 16171 1153 16173 se
rect 1153 16171 1225 16173
tri 1225 16171 1227 16173 nw
tri 570 16160 581 16171 se
rect 581 16165 649 16171
tri 649 16165 655 16171 nw
tri 689 16165 695 16171 se
rect 695 16165 763 16171
tri 763 16165 769 16171 nw
tri 803 16165 809 16171 se
rect 809 16165 877 16171
tri 877 16165 883 16171 nw
tri 917 16165 923 16171 se
rect 923 16165 991 16171
tri 991 16165 997 16171 nw
tri 1031 16165 1037 16171 se
rect 1037 16165 1105 16171
tri 1105 16165 1111 16171 nw
tri 1145 16165 1151 16171 se
rect 1151 16165 1219 16171
tri 1219 16165 1225 16171 nw
rect 581 16160 644 16165
tri 644 16160 649 16165 nw
tri 684 16160 689 16165 se
rect 689 16160 758 16165
tri 758 16160 763 16165 nw
tri 798 16160 803 16165 se
rect 803 16160 872 16165
tri 872 16160 877 16165 nw
tri 912 16160 917 16165 se
rect 917 16160 986 16165
tri 986 16160 991 16165 nw
tri 1026 16160 1031 16165 se
rect 1031 16160 1100 16165
tri 1100 16160 1105 16165 nw
tri 1140 16160 1145 16165 se
rect 1145 16160 1214 16165
tri 1214 16160 1219 16165 nw
rect 2002 16160 16764 16173
rect 16816 16160 16828 16212
rect 16880 16160 16892 16212
rect 16944 16160 16956 16212
rect 17008 16160 17079 16212
tri -3269 16155 -3264 16160 se
rect -3264 16155 -3195 16160
tri -3195 16155 -3190 16160 nw
tri -3155 16155 -3150 16160 se
rect -3150 16155 -3081 16160
tri -3081 16155 -3076 16160 nw
tri -3041 16155 -3036 16160 se
rect -3036 16155 -2967 16160
tri -2967 16155 -2962 16160 nw
tri -2927 16155 -2922 16160 se
rect -2922 16155 -2853 16160
tri -2853 16155 -2848 16160 nw
tri -2813 16155 -2808 16160 se
rect -2808 16155 -2739 16160
tri -2739 16155 -2734 16160 nw
tri -2699 16155 -2694 16160 se
rect -2694 16155 -2625 16160
tri -2625 16155 -2620 16160 nw
tri 565 16155 570 16160 se
rect 570 16155 639 16160
tri 639 16155 644 16160 nw
tri 679 16155 684 16160 se
rect 684 16159 757 16160
tri 757 16159 758 16160 nw
tri 797 16159 798 16160 se
rect 798 16159 871 16160
tri 871 16159 872 16160 nw
tri 911 16159 912 16160 se
rect 912 16159 985 16160
tri 985 16159 986 16160 nw
tri 1025 16159 1026 16160 se
rect 1026 16159 1099 16160
tri 1099 16159 1100 16160 nw
tri 1139 16159 1140 16160 se
rect 1140 16159 1213 16160
tri 1213 16159 1214 16160 nw
rect 684 16155 753 16159
tri 753 16155 757 16159 nw
tri 793 16155 797 16159 se
rect 797 16155 867 16159
tri 867 16155 871 16159 nw
tri 907 16155 911 16159 se
rect 911 16155 981 16159
tri 981 16155 985 16159 nw
tri 1021 16155 1025 16159 se
rect 1025 16155 1095 16159
tri 1095 16155 1099 16159 nw
tri 1135 16155 1139 16159 se
rect 1139 16155 1209 16159
tri 1209 16155 1213 16159 nw
rect 2002 16155 17079 16160
tri -3313 16111 -3269 16155 se
rect -3269 16145 -3205 16155
tri -3205 16145 -3195 16155 nw
tri -3165 16145 -3155 16155 se
rect -3155 16145 -3097 16155
rect -3269 16111 -3239 16145
tri -3239 16111 -3205 16145 nw
tri -3199 16111 -3165 16145 se
rect -3165 16139 -3097 16145
tri -3097 16139 -3081 16155 nw
tri -3057 16139 -3041 16155 se
rect -3041 16139 -2989 16155
rect -3165 16111 -3131 16139
tri -3321 16103 -3313 16111 se
rect -3313 16105 -3245 16111
tri -3245 16105 -3239 16111 nw
tri -3205 16105 -3199 16111 se
rect -3199 16105 -3131 16111
tri -3131 16105 -3097 16139 nw
tri -3091 16105 -3057 16139 se
rect -3057 16133 -2989 16139
tri -2989 16133 -2967 16155 nw
tri -2949 16133 -2927 16155 se
rect -2927 16133 -2881 16155
rect -3057 16105 -3019 16133
rect -3313 16103 -3247 16105
tri -3247 16103 -3245 16105 nw
tri -3207 16103 -3205 16105 se
rect -3205 16103 -3133 16105
tri -3133 16103 -3131 16105 nw
tri -3093 16103 -3091 16105 se
rect -3091 16103 -3019 16105
tri -3019 16103 -2989 16133 nw
tri -2979 16103 -2949 16133 se
rect -2949 16127 -2881 16133
tri -2881 16127 -2853 16155 nw
tri -2841 16127 -2813 16155 se
rect -2813 16127 -2773 16155
rect -2949 16103 -2905 16127
tri -2905 16103 -2881 16127 nw
tri -2865 16103 -2841 16127 se
rect -2841 16121 -2773 16127
tri -2773 16121 -2739 16155 nw
tri -2733 16121 -2699 16155 se
rect -2699 16149 -2631 16155
tri -2631 16149 -2625 16155 nw
tri 559 16149 565 16155 se
rect 565 16149 633 16155
tri 633 16149 639 16155 nw
tri 673 16149 679 16155 se
rect 679 16149 747 16155
tri 747 16149 753 16155 nw
tri 787 16149 793 16155 se
rect 793 16153 865 16155
tri 865 16153 867 16155 nw
tri 905 16153 907 16155 se
rect 907 16153 979 16155
tri 979 16153 981 16155 nw
tri 1019 16153 1021 16155 se
rect 1021 16153 1093 16155
tri 1093 16153 1095 16155 nw
tri 1133 16153 1135 16155 se
rect 1135 16153 1207 16155
tri 1207 16153 1209 16155 nw
rect 793 16149 861 16153
tri 861 16149 865 16153 nw
tri 901 16149 905 16153 se
rect 905 16149 975 16153
tri 975 16149 979 16153 nw
tri 1015 16149 1019 16153 se
rect 1019 16149 1089 16153
tri 1089 16149 1093 16153 nw
tri 1129 16149 1133 16153 se
rect 1133 16149 1203 16153
tri 1203 16149 1207 16153 nw
rect -2699 16121 -2665 16149
rect -2841 16103 -2791 16121
tri -2791 16103 -2773 16121 nw
tri -2751 16103 -2733 16121 se
rect -2733 16115 -2665 16121
tri -2665 16115 -2631 16149 nw
tri -2625 16115 -2591 16149 se
rect -2591 16131 615 16149
tri 615 16131 633 16149 nw
tri 655 16131 673 16149 se
rect 673 16131 723 16149
rect -2591 16115 587 16131
rect -2733 16103 -2677 16115
tri -2677 16103 -2665 16115 nw
tri -2637 16103 -2625 16115 se
rect -2625 16103 587 16115
tri 587 16103 615 16131 nw
tri 627 16103 655 16131 se
rect 655 16125 723 16131
tri 723 16125 747 16149 nw
tri 763 16125 787 16149 se
rect 787 16125 831 16149
rect 655 16103 701 16125
tri 701 16103 723 16125 nw
tri 741 16103 763 16125 se
rect 763 16119 831 16125
tri 831 16119 861 16149 nw
tri 871 16119 901 16149 se
rect 901 16147 973 16149
tri 973 16147 975 16149 nw
tri 1013 16147 1015 16149 se
rect 1015 16147 1087 16149
tri 1087 16147 1089 16149 nw
tri 1127 16147 1129 16149 se
rect 1129 16147 1201 16149
tri 1201 16147 1203 16149 nw
rect 901 16119 939 16147
rect 763 16103 815 16119
tri 815 16103 831 16119 nw
tri 855 16103 871 16119 se
rect 871 16113 939 16119
tri 939 16113 973 16147 nw
tri 979 16113 1013 16147 se
rect 1013 16141 1081 16147
tri 1081 16141 1087 16147 nw
tri 1121 16141 1127 16147 se
rect 1127 16141 1195 16147
tri 1195 16141 1201 16147 nw
rect 1013 16113 1047 16141
rect 871 16103 929 16113
tri 929 16103 939 16113 nw
tri 969 16103 979 16113 se
rect 979 16107 1047 16113
tri 1047 16107 1081 16141 nw
tri 1087 16107 1121 16141 se
rect 1121 16107 1157 16141
rect 979 16103 1043 16107
tri 1043 16103 1047 16107 nw
tri 1083 16103 1087 16107 se
rect 1087 16103 1157 16107
tri 1157 16103 1195 16141 nw
rect 2002 16103 5163 16155
rect 5215 16103 5227 16155
rect 5279 16103 5291 16155
rect 5343 16103 5355 16155
rect 5407 16103 5419 16155
rect 5471 16103 7743 16155
rect 7795 16103 7807 16155
rect 7859 16103 7871 16155
rect 7923 16103 7935 16155
rect 7987 16103 7999 16155
rect 8051 16103 8516 16155
rect 8568 16103 8580 16155
rect 8632 16103 8644 16155
rect 8696 16103 8708 16155
rect 8760 16103 8772 16155
rect 8824 16103 9340 16155
rect 9392 16103 9404 16155
rect 9456 16103 9468 16155
rect 9520 16103 9532 16155
rect 9584 16103 9596 16155
rect 9648 16103 10323 16155
rect 10375 16103 10387 16155
rect 10439 16103 10451 16155
rect 10503 16103 10515 16155
rect 10567 16103 10579 16155
rect 10631 16103 11813 16155
rect 11865 16103 11877 16155
rect 11929 16103 11941 16155
rect 11993 16103 12005 16155
rect 12057 16103 12069 16155
rect 12121 16103 12635 16155
rect 12687 16103 12699 16155
rect 12751 16103 12763 16155
rect 12815 16103 12827 16155
rect 12879 16103 12891 16155
rect 12943 16103 13458 16155
rect 13510 16103 13522 16155
rect 13574 16103 13586 16155
rect 13638 16103 13650 16155
rect 13702 16103 13714 16155
rect 13766 16103 14287 16155
rect 14339 16103 14351 16155
rect 14403 16103 14415 16155
rect 14467 16103 14479 16155
rect 14531 16103 14543 16155
rect 14595 16103 15111 16155
rect 15163 16103 15175 16155
rect 15227 16103 15239 16155
rect 15291 16103 15303 16155
rect 15355 16103 15367 16155
rect 15419 16103 15934 16155
rect 15986 16103 15998 16155
rect 16050 16103 16062 16155
rect 16114 16103 16126 16155
rect 16178 16103 16190 16155
rect 16242 16146 17079 16155
rect 16242 16103 16764 16146
tri -3330 16094 -3321 16103 se
rect -3321 16094 -3256 16103
tri -3256 16094 -3247 16103 nw
tri -3216 16094 -3207 16103 se
rect -3207 16099 -3137 16103
tri -3137 16099 -3133 16103 nw
tri -3097 16099 -3093 16103 se
rect -3093 16099 -3023 16103
tri -3023 16099 -3019 16103 nw
tri -2983 16099 -2979 16103 se
rect -2979 16099 -2914 16103
rect -3207 16094 -3142 16099
tri -3142 16094 -3137 16099 nw
tri -3102 16094 -3097 16099 se
rect -3097 16094 -3028 16099
tri -3028 16094 -3023 16099 nw
tri -2988 16094 -2983 16099 se
rect -2983 16094 -2914 16099
tri -2914 16094 -2905 16103 nw
tri -2874 16094 -2865 16103 se
rect -2865 16094 -2800 16103
tri -2800 16094 -2791 16103 nw
tri -2760 16094 -2751 16103 se
rect -2751 16094 -2686 16103
tri -2686 16094 -2677 16103 nw
tri -2646 16094 -2637 16103 se
rect -2637 16097 581 16103
tri 581 16097 587 16103 nw
tri 621 16097 627 16103 se
rect 627 16097 695 16103
tri 695 16097 701 16103 nw
tri 735 16097 741 16103 se
rect 741 16097 809 16103
tri 809 16097 815 16103 nw
tri 849 16097 855 16103 se
rect 855 16097 923 16103
tri 923 16097 929 16103 nw
tri 963 16097 969 16103 se
rect 969 16097 1037 16103
tri 1037 16097 1043 16103 nw
tri 1077 16097 1083 16103 se
rect 1083 16097 1151 16103
tri 1151 16097 1157 16103 nw
rect -2637 16094 -2572 16097
tri -2572 16094 -2569 16097 nw
tri 618 16094 621 16097 se
rect 621 16094 692 16097
tri 692 16094 695 16097 nw
tri 732 16094 735 16097 se
rect 735 16094 806 16097
tri 806 16094 809 16097 nw
tri 846 16094 849 16097 se
rect 849 16094 920 16097
tri 920 16094 923 16097 nw
tri 960 16094 963 16097 se
rect 963 16094 1034 16097
tri 1034 16094 1037 16097 nw
tri 1074 16094 1077 16097 se
rect 1077 16094 1148 16097
tri 1148 16094 1151 16097 nw
rect 2002 16094 16764 16103
rect 16816 16094 16828 16146
rect 16880 16094 16892 16146
rect 16944 16094 16956 16146
rect 17008 16094 17079 16146
tri -3337 16087 -3330 16094 se
rect -3330 16087 -3263 16094
tri -3263 16087 -3256 16094 nw
tri -3223 16087 -3216 16094 se
rect -3216 16087 -3149 16094
tri -3149 16087 -3142 16094 nw
tri -3109 16087 -3102 16094 se
rect -3102 16093 -3029 16094
tri -3029 16093 -3028 16094 nw
tri -2989 16093 -2988 16094 se
rect -2988 16093 -2915 16094
tri -2915 16093 -2914 16094 nw
tri -2875 16093 -2874 16094 se
rect -2874 16093 -2807 16094
rect -3102 16087 -3035 16093
tri -3035 16087 -3029 16093 nw
tri -2995 16087 -2989 16093 se
rect -2989 16087 -2921 16093
tri -2921 16087 -2915 16093 nw
tri -2881 16087 -2875 16093 se
rect -2875 16087 -2807 16093
tri -2807 16087 -2800 16094 nw
tri -2767 16087 -2760 16094 se
rect -2760 16087 -2695 16094
tri -3339 16085 -3337 16087 se
rect -3337 16085 -3265 16087
tri -3265 16085 -3263 16087 nw
tri -3225 16085 -3223 16087 se
rect -3223 16085 -3151 16087
tri -3151 16085 -3149 16087 nw
tri -3111 16085 -3109 16087 se
rect -3109 16085 -3037 16087
tri -3037 16085 -3035 16087 nw
tri -2997 16085 -2995 16087 se
rect -2995 16085 -2923 16087
tri -2923 16085 -2921 16087 nw
tri -2883 16085 -2881 16087 se
rect -2881 16085 -2809 16087
tri -2809 16085 -2807 16087 nw
tri -2769 16085 -2767 16087 se
rect -2767 16085 -2695 16087
tri -2695 16085 -2686 16094 nw
tri -2655 16085 -2646 16094 se
rect -2646 16085 -2581 16094
tri -2581 16085 -2572 16094 nw
tri 615 16091 618 16094 se
rect 618 16091 689 16094
tri 689 16091 692 16094 nw
tri 729 16091 732 16094 se
rect 732 16091 803 16094
tri 803 16091 806 16094 nw
tri 843 16091 846 16094 se
rect 846 16091 917 16094
tri 917 16091 920 16094 nw
tri 957 16091 960 16094 se
rect 960 16091 1031 16094
tri 1031 16091 1034 16094 nw
tri 1071 16091 1074 16094 se
rect 1074 16091 1145 16094
tri 1145 16091 1148 16094 nw
tri 609 16085 615 16091 se
rect 615 16085 683 16091
tri 683 16085 689 16091 nw
tri 723 16085 729 16091 se
rect 729 16085 797 16091
tri 797 16085 803 16091 nw
tri 837 16085 843 16091 se
rect 843 16085 911 16091
tri 911 16085 917 16091 nw
tri 951 16085 957 16091 se
rect 957 16085 1025 16091
tri 1025 16085 1031 16091 nw
tri 1065 16085 1071 16091 se
rect 1071 16085 1139 16091
tri 1139 16085 1145 16091 nw
rect 2002 16085 17079 16094
tri -3387 16037 -3339 16085 se
rect -3339 16071 -3279 16085
tri -3279 16071 -3265 16085 nw
tri -3239 16071 -3225 16085 se
rect -3225 16071 -3171 16085
rect -3339 16037 -3313 16071
tri -3313 16037 -3279 16071 nw
tri -3273 16037 -3239 16071 se
rect -3239 16065 -3171 16071
tri -3171 16065 -3151 16085 nw
tri -3131 16065 -3111 16085 se
rect -3111 16065 -3063 16085
rect -3239 16037 -3203 16065
tri -3391 16033 -3387 16037 se
rect -3387 16033 -3317 16037
tri -3317 16033 -3313 16037 nw
tri -3277 16033 -3273 16037 se
rect -3273 16033 -3203 16037
tri -3203 16033 -3171 16065 nw
tri -3163 16033 -3131 16065 se
rect -3131 16059 -3063 16065
tri -3063 16059 -3037 16085 nw
tri -3023 16059 -2997 16085 se
rect -2997 16059 -2955 16085
rect -3131 16033 -3089 16059
tri -3089 16033 -3063 16059 nw
tri -3049 16033 -3023 16059 se
rect -3023 16053 -2955 16059
tri -2955 16053 -2923 16085 nw
tri -2915 16053 -2883 16085 se
rect -2883 16081 -2813 16085
tri -2813 16081 -2809 16085 nw
tri -2773 16081 -2769 16085 se
rect -2769 16081 -2699 16085
tri -2699 16081 -2695 16085 nw
tri -2659 16081 -2655 16085 se
rect -2655 16081 -2591 16085
rect -2883 16053 -2847 16081
rect -3023 16033 -2975 16053
tri -2975 16033 -2955 16053 nw
tri -2935 16033 -2915 16053 se
rect -2915 16047 -2847 16053
tri -2847 16047 -2813 16081 nw
tri -2807 16047 -2773 16081 se
rect -2773 16075 -2705 16081
tri -2705 16075 -2699 16081 nw
tri -2665 16075 -2659 16081 se
rect -2659 16075 -2591 16081
tri -2591 16075 -2581 16085 nw
tri 599 16075 609 16085 se
rect 609 16075 673 16085
tri 673 16075 683 16085 nw
tri 713 16075 723 16085 se
rect 723 16079 791 16085
tri 791 16079 797 16085 nw
tri 831 16079 837 16085 se
rect 837 16079 905 16085
tri 905 16079 911 16085 nw
tri 945 16079 951 16085 se
rect 951 16079 1019 16085
tri 1019 16079 1025 16085 nw
tri 1059 16079 1065 16085 se
rect 1065 16079 1133 16085
tri 1133 16079 1139 16085 nw
rect 723 16075 787 16079
tri 787 16075 791 16079 nw
tri 827 16075 831 16079 se
rect 831 16075 901 16079
tri 901 16075 905 16079 nw
tri 941 16075 945 16079 se
rect 945 16075 1015 16079
tri 1015 16075 1019 16079 nw
tri 1055 16075 1059 16079 se
rect 1059 16075 1129 16079
tri 1129 16075 1133 16079 nw
rect -2773 16047 -2739 16075
rect -2915 16033 -2861 16047
tri -2861 16033 -2847 16047 nw
tri -2821 16033 -2807 16047 se
rect -2807 16041 -2739 16047
tri -2739 16041 -2705 16075 nw
tri -2699 16041 -2665 16075 se
rect -2665 16069 -2597 16075
tri -2597 16069 -2591 16075 nw
tri 593 16069 599 16075 se
rect 599 16069 667 16075
tri 667 16069 673 16075 nw
tri 707 16069 713 16075 se
rect 713 16069 781 16075
tri 781 16069 787 16075 nw
tri 821 16069 827 16075 se
rect 827 16073 899 16075
tri 899 16073 901 16075 nw
tri 939 16073 941 16075 se
rect 941 16073 1013 16075
tri 1013 16073 1015 16075 nw
tri 1053 16073 1055 16075 se
rect 1055 16073 1127 16075
tri 1127 16073 1129 16075 nw
rect 827 16069 895 16073
tri 895 16069 899 16073 nw
tri 935 16069 939 16073 se
rect 939 16069 1009 16073
tri 1009 16069 1013 16073 nw
tri 1049 16069 1053 16073 se
rect 1053 16069 1123 16073
tri 1123 16069 1127 16073 nw
rect -2665 16041 -2631 16069
rect -2807 16033 -2747 16041
tri -2747 16033 -2739 16041 nw
tri -2707 16033 -2699 16041 se
rect -2699 16035 -2631 16041
tri -2631 16035 -2597 16069 nw
tri -2591 16035 -2557 16069 se
rect -2557 16051 649 16069
tri 649 16051 667 16069 nw
tri 689 16051 707 16069 se
rect 707 16051 757 16069
rect -2557 16035 631 16051
rect -2699 16033 -2633 16035
tri -2633 16033 -2631 16035 nw
tri -2593 16033 -2591 16035 se
rect -2591 16033 631 16035
tri 631 16033 649 16051 nw
tri 671 16033 689 16051 se
rect 689 16045 757 16051
tri 757 16045 781 16069 nw
tri 797 16045 821 16069 se
rect 821 16045 865 16069
rect 689 16033 745 16045
tri 745 16033 757 16045 nw
tri 785 16033 797 16045 se
rect 797 16039 865 16045
tri 865 16039 895 16069 nw
tri 905 16039 935 16069 se
rect 935 16067 1007 16069
tri 1007 16067 1009 16069 nw
tri 1047 16067 1049 16069 se
rect 1049 16067 1121 16069
tri 1121 16067 1123 16069 nw
rect 935 16039 973 16067
rect 797 16033 859 16039
tri 859 16033 865 16039 nw
tri 899 16033 905 16039 se
rect 905 16033 973 16039
tri 973 16033 1007 16067 nw
tri 1013 16033 1047 16067 se
rect 1047 16033 1087 16067
tri 1087 16033 1121 16067 nw
rect 2002 16033 5163 16085
rect 5215 16033 5227 16085
rect 5279 16033 5291 16085
rect 5343 16033 5355 16085
rect 5407 16033 5419 16085
rect 5471 16033 7743 16085
rect 7795 16033 7807 16085
rect 7859 16033 7871 16085
rect 7923 16033 7935 16085
rect 7987 16033 7999 16085
rect 8051 16033 8516 16085
rect 8568 16033 8580 16085
rect 8632 16033 8644 16085
rect 8696 16033 8708 16085
rect 8760 16033 8772 16085
rect 8824 16033 9340 16085
rect 9392 16033 9404 16085
rect 9456 16033 9468 16085
rect 9520 16033 9532 16085
rect 9584 16033 9596 16085
rect 9648 16033 10323 16085
rect 10375 16033 10387 16085
rect 10439 16033 10451 16085
rect 10503 16033 10515 16085
rect 10567 16033 10579 16085
rect 10631 16033 11813 16085
rect 11865 16033 11877 16085
rect 11929 16033 11941 16085
rect 11993 16033 12005 16085
rect 12057 16033 12069 16085
rect 12121 16033 12635 16085
rect 12687 16033 12699 16085
rect 12751 16033 12763 16085
rect 12815 16033 12827 16085
rect 12879 16033 12891 16085
rect 12943 16033 13458 16085
rect 13510 16033 13522 16085
rect 13574 16033 13586 16085
rect 13638 16033 13650 16085
rect 13702 16033 13714 16085
rect 13766 16033 14287 16085
rect 14339 16033 14351 16085
rect 14403 16033 14415 16085
rect 14467 16033 14479 16085
rect 14531 16033 14543 16085
rect 14595 16033 15111 16085
rect 15163 16033 15175 16085
rect 15227 16033 15239 16085
rect 15291 16033 15303 16085
rect 15355 16033 15367 16085
rect 15419 16033 15934 16085
rect 15986 16033 15998 16085
rect 16050 16033 16062 16085
rect 16114 16033 16126 16085
rect 16178 16033 16190 16085
rect 16242 16079 17079 16085
rect 16242 16033 16764 16079
tri -3397 16027 -3391 16033 se
rect -3391 16031 -3319 16033
tri -3319 16031 -3317 16033 nw
tri -3279 16031 -3277 16033 se
rect -3277 16031 -3205 16033
tri -3205 16031 -3203 16033 nw
tri -3165 16031 -3163 16033 se
rect -3163 16031 -3095 16033
rect -3391 16027 -3323 16031
tri -3323 16027 -3319 16031 nw
tri -3283 16027 -3279 16031 se
rect -3279 16027 -3209 16031
tri -3209 16027 -3205 16031 nw
tri -3169 16027 -3165 16031 se
rect -3165 16027 -3095 16031
tri -3095 16027 -3089 16033 nw
tri -3055 16027 -3049 16033 se
rect -3049 16027 -2981 16033
tri -2981 16027 -2975 16033 nw
tri -2941 16027 -2935 16033 se
rect -2935 16027 -2867 16033
tri -2867 16027 -2861 16033 nw
tri -2827 16027 -2821 16033 se
rect -2821 16027 -2753 16033
tri -2753 16027 -2747 16033 nw
tri -2713 16027 -2707 16033 se
rect -2707 16027 -2639 16033
tri -2639 16027 -2633 16033 nw
tri -2599 16027 -2593 16033 se
rect -2593 16027 625 16033
tri 625 16027 631 16033 nw
tri 665 16027 671 16033 se
rect 671 16027 739 16033
tri 739 16027 745 16033 nw
tri 779 16027 785 16033 se
rect 785 16027 853 16033
tri 853 16027 859 16033 nw
tri 893 16027 899 16033 se
rect 899 16027 967 16033
tri 967 16027 973 16033 nw
tri 1007 16027 1013 16033 se
rect 1013 16027 1081 16033
tri 1081 16027 1087 16033 nw
rect 2002 16027 16764 16033
rect 16816 16027 16828 16079
rect 16880 16027 16892 16079
rect 16944 16027 16956 16079
rect 17008 16027 17079 16079
tri -3409 16015 -3397 16027 se
rect -3397 16015 -3335 16027
tri -3335 16015 -3323 16027 nw
tri -3295 16015 -3283 16027 se
rect -3283 16025 -3211 16027
tri -3211 16025 -3209 16027 nw
tri -3171 16025 -3169 16027 se
rect -3169 16025 -3097 16027
tri -3097 16025 -3095 16027 nw
tri -3057 16025 -3055 16027 se
rect -3055 16025 -2989 16027
rect -3283 16015 -3221 16025
tri -3221 16015 -3211 16025 nw
tri -3181 16015 -3171 16025 se
rect -3171 16019 -3103 16025
tri -3103 16019 -3097 16025 nw
tri -3063 16019 -3057 16025 se
rect -3057 16019 -2989 16025
tri -2989 16019 -2981 16027 nw
tri -2949 16019 -2941 16027 se
rect -2941 16019 -2879 16027
rect -3171 16015 -3107 16019
tri -3107 16015 -3103 16019 nw
tri -3067 16015 -3063 16019 se
rect -3063 16015 -2993 16019
tri -2993 16015 -2989 16019 nw
tri -2953 16015 -2949 16019 se
rect -2949 16015 -2879 16019
tri -2879 16015 -2867 16027 nw
tri -2839 16015 -2827 16027 se
rect -2827 16015 -2765 16027
tri -2765 16015 -2753 16027 nw
tri -2725 16015 -2713 16027 se
rect -2713 16015 -2651 16027
tri -2651 16015 -2639 16027 nw
tri -2611 16015 -2599 16027 se
rect -2599 16017 615 16027
tri 615 16017 625 16027 nw
tri 655 16017 665 16027 se
rect 665 16017 729 16027
tri 729 16017 739 16027 nw
tri 769 16017 779 16027 se
rect 779 16017 843 16027
tri 843 16017 853 16027 nw
tri 883 16017 893 16027 se
rect 893 16017 957 16027
tri 957 16017 967 16027 nw
tri 997 16017 1007 16027 se
rect 1007 16017 1071 16027
tri 1071 16017 1081 16027 nw
rect -2599 16015 -2537 16017
tri -2537 16015 -2535 16017 nw
tri 653 16015 655 16017 se
rect 655 16015 727 16017
tri 727 16015 729 16017 nw
tri 767 16015 769 16017 se
rect 769 16015 841 16017
tri 841 16015 843 16017 nw
tri 881 16015 883 16017 se
rect 883 16015 955 16017
tri 955 16015 957 16017 nw
tri 995 16015 997 16017 se
rect 997 16015 1069 16017
tri 1069 16015 1071 16017 nw
rect 2002 16015 17079 16027
tri -3411 16013 -3409 16015 se
rect -3409 16013 -3337 16015
tri -3337 16013 -3335 16015 nw
tri -3297 16013 -3295 16015 se
rect -3295 16013 -3223 16015
tri -3223 16013 -3221 16015 nw
tri -3183 16013 -3181 16015 se
rect -3181 16013 -3109 16015
tri -3109 16013 -3107 16015 nw
tri -3069 16013 -3067 16015 se
rect -3067 16013 -2995 16015
tri -2995 16013 -2993 16015 nw
tri -2955 16013 -2953 16015 se
rect -2953 16013 -2881 16015
tri -2881 16013 -2879 16015 nw
tri -2841 16013 -2839 16015 se
rect -2839 16013 -2773 16015
tri -3430 15994 -3411 16013 se
rect -3411 16000 -3350 16013
tri -3350 16000 -3337 16013 nw
tri -3310 16000 -3297 16013 se
rect -3297 16000 -3245 16013
rect -3411 15994 -3356 16000
tri -3356 15994 -3350 16000 nw
tri -3316 15994 -3310 16000 se
rect -3310 15994 -3245 16000
rect -3430 15989 -3361 15994
tri -3361 15989 -3356 15994 nw
tri -3321 15989 -3316 15994 se
rect -3316 15991 -3245 15994
tri -3245 15991 -3223 16013 nw
tri -3205 15991 -3183 16013 se
rect -3183 15991 -3133 16013
rect -3316 15989 -3247 15991
tri -3247 15989 -3245 15991 nw
tri -3207 15989 -3205 15991 se
rect -3205 15989 -3133 15991
tri -3133 15989 -3109 16013 nw
tri -3093 15989 -3069 16013 se
rect -3069 15989 -3019 16013
tri -3019 15989 -2995 16013 nw
tri -2979 15989 -2955 16013 se
rect -2955 16007 -2887 16013
tri -2887 16007 -2881 16013 nw
tri -2847 16007 -2841 16013 se
rect -2841 16007 -2773 16013
tri -2773 16007 -2765 16015 nw
tri -2733 16007 -2725 16015 se
rect -2725 16007 -2665 16015
rect -2955 15989 -2905 16007
tri -2905 15989 -2887 16007 nw
tri -2865 15989 -2847 16007 se
rect -2847 16001 -2779 16007
tri -2779 16001 -2773 16007 nw
tri -2739 16001 -2733 16007 se
rect -2733 16001 -2665 16007
tri -2665 16001 -2651 16015 nw
tri -2625 16001 -2611 16015 se
rect -2611 16001 -2557 16015
rect -2847 15989 -2791 16001
tri -2791 15989 -2779 16001 nw
tri -2751 15989 -2739 16001 se
rect -2739 15995 -2671 16001
tri -2671 15995 -2665 16001 nw
tri -2631 15995 -2625 16001 se
rect -2625 15995 -2557 16001
tri -2557 15995 -2537 16015 nw
tri 649 16011 653 16015 se
rect 653 16011 723 16015
tri 723 16011 727 16015 nw
tri 763 16011 767 16015 se
rect 767 16011 837 16015
tri 837 16011 841 16015 nw
tri 877 16011 881 16015 se
rect 881 16011 951 16015
tri 951 16011 955 16015 nw
tri 991 16011 995 16015 se
rect 995 16011 1065 16015
tri 1065 16011 1069 16015 nw
tri 633 15995 649 16011 se
rect 649 16005 717 16011
tri 717 16005 723 16011 nw
tri 757 16005 763 16011 se
rect 763 16005 831 16011
tri 831 16005 837 16011 nw
tri 871 16005 877 16011 se
rect 877 16005 945 16011
tri 945 16005 951 16011 nw
tri 985 16005 991 16011 se
rect 991 16005 1059 16011
tri 1059 16005 1065 16011 nw
rect 649 15995 707 16005
tri 707 15995 717 16005 nw
tri 747 15995 757 16005 se
rect 757 15999 825 16005
tri 825 15999 831 16005 nw
tri 865 15999 871 16005 se
rect 871 15999 939 16005
tri 939 15999 945 16005 nw
tri 979 15999 985 16005 se
rect 985 15999 1053 16005
tri 1053 15999 1059 16005 nw
rect 757 15995 821 15999
tri 821 15995 825 15999 nw
tri 861 15995 865 15999 se
rect 865 15995 935 15999
tri 935 15995 939 15999 nw
tri 975 15995 979 15999 se
rect 979 15995 1049 15999
tri 1049 15995 1053 15999 nw
rect -2739 15989 -2677 15995
tri -2677 15989 -2671 15995 nw
tri -2637 15989 -2631 15995 se
rect -2631 15989 -2563 15995
tri -2563 15989 -2557 15995 nw
tri 627 15989 633 15995 se
rect 633 15989 701 15995
tri 701 15989 707 15995 nw
tri 741 15989 747 15995 se
rect 747 15989 815 15995
tri 815 15989 821 15995 nw
tri 855 15989 861 15995 se
rect 861 15993 933 15995
tri 933 15993 935 15995 nw
tri 973 15993 975 15995 se
rect 975 15993 1047 15995
tri 1047 15993 1049 15995 nw
rect 861 15989 929 15993
tri 929 15989 933 15993 nw
tri 969 15989 973 15993 se
rect 973 15989 1043 15993
tri 1043 15989 1047 15993 nw
rect -3430 1950 -3378 15989
tri -3378 15972 -3361 15989 nw
tri -3338 15972 -3321 15989 se
rect -3321 15972 -3273 15989
tri -3347 15963 -3338 15972 se
rect -3338 15963 -3273 15972
tri -3273 15963 -3247 15989 nw
tri -3233 15963 -3207 15989 se
rect -3207 15985 -3137 15989
tri -3137 15985 -3133 15989 nw
tri -3097 15985 -3093 15989 se
rect -3093 15985 -3029 15989
rect -3207 15963 -3159 15985
tri -3159 15963 -3137 15985 nw
tri -3119 15963 -3097 15985 se
rect -3097 15979 -3029 15985
tri -3029 15979 -3019 15989 nw
tri -2989 15979 -2979 15989 se
rect -2979 15979 -2921 15989
rect -3097 15963 -3045 15979
tri -3045 15963 -3029 15979 nw
tri -3005 15963 -2989 15979 se
rect -2989 15973 -2921 15979
tri -2921 15973 -2905 15989 nw
tri -2881 15973 -2865 15989 se
rect -2865 15973 -2813 15989
rect -2989 15963 -2931 15973
tri -2931 15963 -2921 15973 nw
tri -2891 15963 -2881 15973 se
rect -2881 15967 -2813 15973
tri -2813 15967 -2791 15989 nw
tri -2773 15967 -2751 15989 se
rect -2751 15967 -2703 15989
rect -2881 15963 -2817 15967
tri -2817 15963 -2813 15967 nw
tri -2777 15963 -2773 15967 se
rect -2773 15963 -2703 15967
tri -2703 15963 -2677 15989 nw
tri -2663 15963 -2637 15989 se
rect -2637 15963 -2589 15989
tri -2589 15963 -2563 15989 nw
tri -2549 15963 -2523 15989 se
rect -2523 15971 683 15989
tri 683 15971 701 15989 nw
tri 723 15971 741 15989 se
rect 741 15971 791 15989
rect -2523 15963 675 15971
tri 675 15963 683 15971 nw
tri 715 15963 723 15971 se
rect 723 15965 791 15971
tri 791 15965 815 15989 nw
tri 831 15965 855 15989 se
rect 855 15965 903 15989
rect 723 15963 789 15965
tri 789 15963 791 15965 nw
tri 829 15963 831 15965 se
rect 831 15963 903 15965
tri 903 15963 929 15989 nw
tri 943 15963 969 15989 se
rect 969 15963 1017 15989
tri 1017 15963 1043 15989 nw
rect 2002 15963 5163 16015
rect 5215 15963 5227 16015
rect 5279 15963 5291 16015
rect 5343 15963 5355 16015
rect 5407 15963 5419 16015
rect 5471 15963 7743 16015
rect 7795 15963 7807 16015
rect 7859 15963 7871 16015
rect 7923 15963 7935 16015
rect 7987 15963 7999 16015
rect 8051 15963 8516 16015
rect 8568 15963 8580 16015
rect 8632 15963 8644 16015
rect 8696 15963 8708 16015
rect 8760 15963 8772 16015
rect 8824 15963 9340 16015
rect 9392 15963 9404 16015
rect 9456 15963 9468 16015
rect 9520 15963 9532 16015
rect 9584 15963 9596 16015
rect 9648 15963 10323 16015
rect 10375 15963 10387 16015
rect 10439 15963 10451 16015
rect 10503 15963 10515 16015
rect 10567 15963 10579 16015
rect 10631 15963 11813 16015
rect 11865 15963 11877 16015
rect 11929 15963 11941 16015
rect 11993 15963 12005 16015
rect 12057 15963 12069 16015
rect 12121 15963 12635 16015
rect 12687 15963 12699 16015
rect 12751 15963 12763 16015
rect 12815 15963 12827 16015
rect 12879 15963 12891 16015
rect 12943 15963 13458 16015
rect 13510 15963 13522 16015
rect 13574 15963 13586 16015
rect 13638 15963 13650 16015
rect 13702 15963 13714 16015
rect 13766 15963 14287 16015
rect 14339 15963 14351 16015
rect 14403 15963 14415 16015
rect 14467 15963 14479 16015
rect 14531 15963 14543 16015
rect 14595 15963 15111 16015
rect 15163 15963 15175 16015
rect 15227 15963 15239 16015
rect 15291 15963 15303 16015
rect 15355 15963 15367 16015
rect 15419 15963 15934 16015
rect 15986 15963 15998 16015
rect 16050 15963 16062 16015
rect 16114 15963 16126 16015
rect 16178 15963 16190 16015
rect 16242 16012 17079 16015
rect 16242 15963 16764 16012
rect -3430 1886 -3378 1898
rect -3430 1828 -3378 1834
tri -3350 15960 -3347 15963 se
rect -3347 15960 -3276 15963
tri -3276 15960 -3273 15963 nw
tri -3236 15960 -3233 15963 se
rect -3233 15960 -3162 15963
tri -3162 15960 -3159 15963 nw
tri -3122 15960 -3119 15963 se
rect -3119 15960 -3048 15963
tri -3048 15960 -3045 15963 nw
tri -3008 15960 -3005 15963 se
rect -3005 15960 -2934 15963
tri -2934 15960 -2931 15963 nw
tri -2894 15960 -2891 15963 se
rect -2891 15960 -2820 15963
tri -2820 15960 -2817 15963 nw
tri -2780 15960 -2777 15963 se
rect -2777 15961 -2705 15963
tri -2705 15961 -2703 15963 nw
tri -2665 15961 -2663 15963 se
rect -2663 15961 -2592 15963
rect -2777 15960 -2706 15961
tri -2706 15960 -2705 15961 nw
tri -2666 15960 -2665 15961 se
rect -2665 15960 -2592 15961
tri -2592 15960 -2589 15963 nw
tri -2552 15960 -2549 15963 se
rect -2549 15960 672 15963
tri 672 15960 675 15963 nw
tri 712 15960 715 15963 se
rect 715 15960 786 15963
tri 786 15960 789 15963 nw
tri 826 15960 829 15963 se
rect 829 15960 900 15963
tri 900 15960 903 15963 nw
tri 940 15960 943 15963 se
rect 943 15960 1014 15963
tri 1014 15960 1017 15963 nw
rect 2002 15960 16764 15963
rect 16816 15960 16828 16012
rect 16880 15960 16892 16012
rect 16944 15960 16956 16012
rect 17008 15960 17079 16012
rect -3350 15945 -3291 15960
tri -3291 15945 -3276 15960 nw
tri -3245 15951 -3236 15960 se
rect -3236 15951 -3171 15960
tri -3171 15951 -3162 15960 nw
tri -3131 15951 -3122 15960 se
rect -3122 15951 -3063 15960
tri -3251 15945 -3245 15951 se
rect -3245 15945 -3177 15951
tri -3177 15945 -3171 15951 nw
tri -3137 15945 -3131 15951 se
rect -3131 15945 -3063 15951
tri -3063 15945 -3048 15960 nw
tri -3023 15945 -3008 15960 se
rect -3008 15945 -2949 15960
tri -2949 15945 -2934 15960 nw
tri -2909 15945 -2894 15960 se
rect -2894 15945 -2835 15960
tri -2835 15945 -2820 15960 nw
tri -2795 15945 -2780 15960 se
rect -2780 15945 -2721 15960
tri -2721 15945 -2706 15960 nw
tri -2681 15945 -2666 15960 se
rect -2666 15955 -2597 15960
tri -2597 15955 -2592 15960 nw
tri -2557 15955 -2552 15960 se
rect -2552 15955 657 15960
rect -2666 15945 -2607 15955
tri -2607 15945 -2597 15955 nw
tri -2567 15945 -2557 15955 se
rect -2557 15945 657 15955
tri 657 15945 672 15960 nw
tri 697 15945 712 15960 se
rect 712 15945 771 15960
tri 771 15945 786 15960 nw
tri 811 15945 826 15960 se
rect 826 15959 899 15960
tri 899 15959 900 15960 nw
tri 939 15959 940 15960 se
rect 940 15959 999 15960
rect 826 15945 885 15959
tri 885 15945 899 15959 nw
tri 925 15945 939 15959 se
rect 939 15945 999 15959
tri 999 15945 1014 15960 nw
rect 2002 15945 17079 15960
rect -3350 15939 -3297 15945
tri -3297 15939 -3291 15945 nw
tri -3257 15939 -3251 15945 se
rect -3251 15939 -3183 15945
tri -3183 15939 -3177 15945 nw
tri -3143 15939 -3137 15945 se
rect -3137 15939 -3069 15945
tri -3069 15939 -3063 15945 nw
tri -3029 15939 -3023 15945 se
rect -3023 15939 -2955 15945
tri -2955 15939 -2949 15945 nw
tri -2915 15939 -2909 15945 se
rect -2909 15939 -2847 15945
rect -3350 2106 -3298 15939
tri -3298 15938 -3297 15939 nw
tri -3258 15938 -3257 15939 se
rect -3257 15938 -3190 15939
tri -3270 15926 -3258 15938 se
rect -3258 15932 -3190 15938
tri -3190 15932 -3183 15939 nw
tri -3150 15932 -3143 15939 se
rect -3143 15932 -3093 15939
rect -3258 15926 -3196 15932
tri -3196 15926 -3190 15932 nw
tri -3156 15926 -3150 15932 se
rect -3150 15926 -3093 15932
rect -3270 15915 -3207 15926
tri -3207 15915 -3196 15926 nw
tri -3167 15915 -3156 15926 se
rect -3156 15915 -3093 15926
tri -3093 15915 -3069 15939 nw
tri -3053 15915 -3029 15939 se
rect -3029 15933 -2961 15939
tri -2961 15933 -2955 15939 nw
tri -2921 15933 -2915 15939 se
rect -2915 15933 -2847 15939
tri -2847 15933 -2835 15945 nw
tri -2807 15933 -2795 15945 se
rect -2795 15933 -2739 15945
rect -3029 15915 -2979 15933
tri -2979 15915 -2961 15933 nw
tri -2939 15915 -2921 15933 se
rect -2921 15927 -2853 15933
tri -2853 15927 -2847 15933 nw
tri -2813 15927 -2807 15933 se
rect -2807 15927 -2739 15933
tri -2739 15927 -2721 15945 nw
tri -2699 15927 -2681 15945 se
rect -2681 15927 -2631 15945
rect -2921 15915 -2865 15927
tri -2865 15915 -2853 15927 nw
tri -2825 15915 -2813 15927 se
rect -2813 15921 -2745 15927
tri -2745 15921 -2739 15927 nw
tri -2705 15921 -2699 15927 se
rect -2699 15921 -2631 15927
tri -2631 15921 -2607 15945 nw
tri -2591 15921 -2567 15945 se
rect -2567 15937 649 15945
tri 649 15937 657 15945 nw
tri 689 15937 697 15945 se
rect 697 15937 763 15945
tri 763 15937 771 15945 nw
tri 803 15937 811 15945 se
rect 811 15937 877 15945
tri 877 15937 885 15945 nw
tri 917 15937 925 15945 se
rect 925 15937 991 15945
tri 991 15937 999 15945 nw
rect -2567 15921 -2523 15937
rect -2813 15915 -2751 15921
tri -2751 15915 -2745 15921 nw
tri -2711 15915 -2705 15921 se
rect -2705 15915 -2637 15921
tri -2637 15915 -2631 15921 nw
tri -2597 15915 -2591 15921 se
rect -2591 15915 -2523 15921
tri -2523 15915 -2501 15937 nw
tri 683 15931 689 15937 se
rect 689 15931 757 15937
tri 757 15931 763 15937 nw
tri 797 15931 803 15937 se
rect 803 15931 871 15937
tri 871 15931 877 15937 nw
tri 911 15931 917 15937 se
rect 917 15931 985 15937
tri 985 15931 991 15937 nw
tri 667 15915 683 15931 se
rect 683 15925 751 15931
tri 751 15925 757 15931 nw
tri 791 15925 797 15931 se
rect 797 15925 865 15931
tri 865 15925 871 15931 nw
tri 905 15925 911 15931 se
rect 911 15925 979 15931
tri 979 15925 985 15931 nw
rect 683 15915 741 15925
tri 741 15915 751 15925 nw
tri 781 15915 791 15925 se
rect 791 15919 859 15925
tri 859 15919 865 15925 nw
tri 899 15919 905 15925 se
rect 905 15919 973 15925
tri 973 15919 979 15925 nw
rect 791 15915 855 15919
tri 855 15915 859 15919 nw
tri 895 15915 899 15919 se
rect 899 15915 969 15919
tri 969 15915 973 15919 nw
rect -3270 2230 -3218 15915
tri -3218 15904 -3207 15915 nw
tri -3178 15904 -3167 15915 se
rect -3167 15905 -3103 15915
tri -3103 15905 -3093 15915 nw
tri -3063 15905 -3053 15915 se
rect -3053 15905 -2995 15915
rect -3167 15904 -3115 15905
tri -3189 15893 -3178 15904 se
rect -3178 15893 -3115 15904
tri -3115 15893 -3103 15905 nw
tri -3075 15893 -3063 15905 se
rect -3063 15899 -2995 15905
tri -2995 15899 -2979 15915 nw
tri -2955 15899 -2939 15915 se
rect -2939 15899 -2887 15915
rect -3063 15893 -3001 15899
tri -3001 15893 -2995 15899 nw
tri -2961 15893 -2955 15899 se
rect -2955 15893 -2887 15899
tri -2887 15893 -2865 15915 nw
tri -2847 15893 -2825 15915 se
rect -2825 15893 -2773 15915
tri -2773 15893 -2751 15915 nw
tri -2733 15893 -2711 15915 se
rect -2711 15893 -2659 15915
tri -2659 15893 -2637 15915 nw
tri -2619 15893 -2597 15915 se
rect -2597 15909 -2529 15915
tri -2529 15909 -2523 15915 nw
tri 661 15909 667 15915 se
rect 667 15909 735 15915
tri 735 15909 741 15915 nw
tri 775 15909 781 15915 se
rect 781 15909 849 15915
tri 849 15909 855 15915 nw
tri 889 15909 895 15915 se
rect 895 15909 963 15915
tri 963 15909 969 15915 nw
rect -2597 15893 -2545 15909
tri -2545 15893 -2529 15909 nw
tri -2505 15893 -2489 15909 se
rect -2489 15893 719 15909
tri 719 15893 735 15909 nw
tri 759 15893 775 15909 se
rect 775 15893 833 15909
tri 833 15893 849 15909 nw
tri 873 15893 889 15909 se
rect 889 15893 947 15909
tri 947 15893 963 15909 nw
rect 2002 15893 5163 15945
rect 5215 15893 5227 15945
rect 5279 15893 5291 15945
rect 5343 15893 5355 15945
rect 5407 15893 5419 15945
rect 5471 15893 7743 15945
rect 7795 15893 7807 15945
rect 7859 15893 7871 15945
rect 7923 15893 7935 15945
rect 7987 15893 7999 15945
rect 8051 15893 8516 15945
rect 8568 15893 8580 15945
rect 8632 15893 8644 15945
rect 8696 15893 8708 15945
rect 8760 15893 8772 15945
rect 8824 15893 9340 15945
rect 9392 15893 9404 15945
rect 9456 15893 9468 15945
rect 9520 15893 9532 15945
rect 9584 15893 9596 15945
rect 9648 15893 10323 15945
rect 10375 15893 10387 15945
rect 10439 15893 10451 15945
rect 10503 15893 10515 15945
rect 10567 15893 10579 15945
rect 10631 15893 11813 15945
rect 11865 15893 11877 15945
rect 11929 15893 11941 15945
rect 11993 15893 12005 15945
rect 12057 15893 12069 15945
rect 12121 15893 12635 15945
rect 12687 15893 12699 15945
rect 12751 15893 12763 15945
rect 12815 15893 12827 15945
rect 12879 15893 12891 15945
rect 12943 15893 13458 15945
rect 13510 15893 13522 15945
rect 13574 15893 13586 15945
rect 13638 15893 13650 15945
rect 13702 15893 13714 15945
rect 13766 15893 14287 15945
rect 14339 15893 14351 15945
rect 14403 15893 14415 15945
rect 14467 15893 14479 15945
rect 14531 15893 14543 15945
rect 14595 15893 15111 15945
rect 15163 15893 15175 15945
rect 15227 15893 15239 15945
rect 15291 15893 15303 15945
rect 15355 15893 15367 15945
rect 15419 15893 15934 15945
rect 15986 15893 15998 15945
rect 16050 15893 16062 15945
rect 16114 15893 16126 15945
rect 16178 15893 16190 15945
rect 16242 15893 16764 15945
rect 16816 15893 16828 15945
rect 16880 15893 16892 15945
rect 16944 15893 16956 15945
rect 17008 15893 17079 15945
tri -3190 15892 -3189 15893 se
rect -3189 15892 -3116 15893
tri -3116 15892 -3115 15893 nw
tri -3076 15892 -3075 15893 se
rect -3075 15892 -3007 15893
rect -3190 15887 -3121 15892
tri -3121 15887 -3116 15892 nw
tri -3081 15887 -3076 15892 se
rect -3076 15887 -3007 15892
tri -3007 15887 -3001 15893 nw
tri -2967 15887 -2961 15893 se
rect -2961 15887 -2893 15893
tri -2893 15887 -2887 15893 nw
tri -2853 15887 -2847 15893 se
rect -2847 15887 -2779 15893
tri -2779 15887 -2773 15893 nw
tri -2739 15887 -2733 15893 se
rect -2733 15887 -2665 15893
tri -2665 15887 -2659 15893 nw
tri -2625 15887 -2619 15893 se
rect -2619 15887 -2551 15893
tri -2551 15887 -2545 15893 nw
tri -2511 15887 -2505 15893 se
rect -2505 15891 717 15893
tri 717 15891 719 15893 nw
tri 757 15891 759 15893 se
rect 759 15891 827 15893
rect -2505 15887 713 15891
tri 713 15887 717 15891 nw
tri 753 15887 757 15891 se
rect 757 15887 827 15891
tri 827 15887 833 15893 nw
tri 867 15887 873 15893 se
rect 873 15887 941 15893
tri 941 15887 947 15893 nw
rect -3190 15881 -3127 15887
tri -3127 15881 -3121 15887 nw
tri -3087 15881 -3081 15887 se
rect -3081 15881 -3013 15887
tri -3013 15881 -3007 15887 nw
tri -2973 15881 -2967 15887 se
rect -2967 15881 -2899 15887
tri -2899 15881 -2893 15887 nw
tri -2859 15881 -2853 15887 se
rect -2853 15881 -2785 15887
tri -2785 15881 -2779 15887 nw
tri -2745 15881 -2739 15887 se
rect -2739 15881 -2671 15887
tri -2671 15881 -2665 15887 nw
tri -2631 15881 -2625 15887 se
rect -2625 15881 -2557 15887
tri -2557 15881 -2551 15887 nw
tri -2517 15881 -2511 15887 se
rect -2511 15881 683 15887
rect -3190 3017 -3138 15881
tri -3138 15870 -3127 15881 nw
tri -3098 15870 -3087 15881 se
rect -3087 15870 -3029 15881
tri -3103 15865 -3098 15870 se
rect -3098 15865 -3029 15870
tri -3029 15865 -3013 15881 nw
tri -2989 15865 -2973 15881 se
rect -2973 15865 -2921 15881
tri -3110 15858 -3103 15865 se
rect -3103 15859 -3035 15865
tri -3035 15859 -3029 15865 nw
tri -2995 15859 -2989 15865 se
rect -2989 15859 -2921 15865
tri -2921 15859 -2899 15881 nw
tri -2881 15859 -2859 15881 se
rect -2859 15859 -2813 15881
rect -3103 15858 -3036 15859
tri -3036 15858 -3035 15859 nw
tri -2996 15858 -2995 15859 se
rect -2995 15858 -2927 15859
rect -3110 15841 -3053 15858
tri -3053 15841 -3036 15858 nw
tri -3013 15841 -2996 15858 se
rect -2996 15853 -2927 15858
tri -2927 15853 -2921 15859 nw
tri -2887 15853 -2881 15859 se
rect -2881 15853 -2813 15859
tri -2813 15853 -2785 15881 nw
tri -2773 15853 -2745 15881 se
rect -2745 15853 -2705 15881
rect -2996 15841 -2939 15853
tri -2939 15841 -2927 15853 nw
tri -2899 15841 -2887 15853 se
rect -2887 15847 -2819 15853
tri -2819 15847 -2813 15853 nw
tri -2779 15847 -2773 15853 se
rect -2773 15847 -2705 15853
tri -2705 15847 -2671 15881 nw
tri -2665 15847 -2631 15881 se
rect -2631 15875 -2563 15881
tri -2563 15875 -2557 15881 nw
tri -2523 15875 -2517 15881 se
rect -2517 15875 683 15881
rect -2631 15847 -2597 15875
rect -2887 15841 -2825 15847
tri -2825 15841 -2819 15847 nw
tri -2785 15841 -2779 15847 se
rect -2779 15841 -2711 15847
tri -2711 15841 -2705 15847 nw
tri -2671 15841 -2665 15847 se
rect -2665 15841 -2597 15847
tri -2597 15841 -2563 15875 nw
tri -2557 15841 -2523 15875 se
rect -2523 15857 683 15875
tri 683 15857 713 15887 nw
tri 723 15857 753 15887 se
rect 753 15885 825 15887
tri 825 15885 827 15887 nw
tri 865 15885 867 15887 se
rect 867 15885 911 15887
rect 753 15857 797 15885
tri 797 15857 825 15885 nw
tri 837 15857 865 15885 se
rect 865 15857 911 15885
tri 911 15857 941 15887 nw
rect 2002 15881 17079 15893
rect 2002 15878 15026 15881
tri 15026 15878 15029 15881 nw
tri 15440 15878 15443 15881 ne
rect 15443 15878 17079 15881
rect 2002 15857 2123 15878
tri 2123 15857 2144 15878 nw
tri 4993 15857 5014 15878 ne
rect 5014 15857 5027 15878
rect -2523 15841 -2489 15857
rect -3110 3244 -3058 15841
tri -3058 15836 -3053 15841 nw
tri -3018 15836 -3013 15841 se
rect -3013 15836 -2950 15841
tri -3025 15829 -3018 15836 se
rect -3018 15830 -2950 15836
tri -2950 15830 -2939 15841 nw
tri -2910 15830 -2899 15841 se
rect -2899 15830 -2837 15841
rect -3018 15829 -2951 15830
tri -2951 15829 -2950 15830 nw
tri -2911 15829 -2910 15830 se
rect -2910 15829 -2837 15830
tri -2837 15829 -2825 15841 nw
tri -2797 15829 -2785 15841 se
rect -2785 15829 -2723 15841
tri -2723 15829 -2711 15841 nw
tri -2683 15829 -2671 15841 se
rect -2671 15835 -2603 15841
tri -2603 15835 -2597 15841 nw
tri -2563 15835 -2557 15841 se
rect -2557 15835 -2489 15841
tri -2489 15835 -2467 15857 nw
tri 717 15851 723 15857 se
rect 723 15851 791 15857
tri 791 15851 797 15857 nw
tri 831 15851 837 15857 se
rect 837 15851 905 15857
tri 905 15851 911 15857 nw
rect 2002 15851 2117 15857
tri 2117 15851 2123 15857 nw
tri 5014 15851 5020 15857 ne
rect 5020 15851 5027 15857
tri 701 15835 717 15851 se
rect 717 15845 785 15851
tri 785 15845 791 15851 nw
tri 825 15845 831 15851 se
rect 831 15845 899 15851
tri 899 15845 905 15851 nw
rect 2002 15845 2111 15851
tri 2111 15845 2117 15851 nw
tri 5020 15845 5026 15851 ne
rect 5026 15845 5027 15851
rect 717 15835 775 15845
tri 775 15835 785 15845 nw
tri 815 15835 825 15845 se
rect 825 15835 889 15845
tri 889 15835 899 15845 nw
rect 2002 15844 2110 15845
tri 2110 15844 2111 15845 nw
tri 5026 15844 5027 15845 ne
rect 5593 15857 5606 15878
tri 5606 15857 5627 15878 nw
tri 10282 15857 10303 15878 ne
rect 10303 15871 11159 15878
tri 11159 15871 11166 15878 nw
rect 12626 15871 12954 15878
tri 12954 15871 12961 15878 nw
tri 13639 15871 13646 15878 ne
rect 13646 15871 13983 15878
rect 10303 15857 11023 15871
rect 5593 15851 5600 15857
tri 5600 15851 5606 15857 nw
tri 10303 15851 10309 15857 ne
rect 10309 15851 11023 15857
rect 5593 15845 5594 15851
tri 5594 15845 5600 15851 nw
tri 10309 15845 10315 15851 ne
rect 10315 15845 11023 15851
tri 5593 15844 5594 15845 nw
tri 10315 15844 10316 15845 ne
rect 10316 15844 11023 15845
rect 2002 15835 2101 15844
tri 2101 15835 2110 15844 nw
tri 10316 15835 10325 15844 ne
rect 10325 15835 11023 15844
rect -2671 15829 -2609 15835
tri -2609 15829 -2603 15835 nw
tri -2569 15829 -2563 15835 se
rect -2563 15829 -2495 15835
tri -2495 15829 -2489 15835 nw
tri 695 15829 701 15835 se
rect 701 15829 769 15835
tri 769 15829 775 15835 nw
tri 809 15829 815 15835 se
rect 815 15829 883 15835
tri 883 15829 889 15835 nw
rect 2002 15829 2095 15835
tri 2095 15829 2101 15835 nw
tri 10325 15829 10331 15835 ne
rect 10331 15829 11023 15835
rect -3110 3180 -3058 3192
rect -3110 3122 -3058 3128
tri -3030 15824 -3025 15829 se
rect -3025 15824 -2956 15829
tri -2956 15824 -2951 15829 nw
tri -2916 15824 -2911 15829 se
rect -2911 15824 -2853 15829
rect -3030 3074 -2978 15824
tri -2978 15802 -2956 15824 nw
tri -2938 15802 -2916 15824 se
rect -2916 15813 -2853 15824
tri -2853 15813 -2837 15829 nw
tri -2813 15813 -2797 15829 se
rect -2797 15813 -2745 15829
rect -2916 15802 -2876 15813
rect -3106 3022 -3100 3074
rect -3048 3022 -3036 3074
rect -2984 3022 -2978 3074
tri -2950 15790 -2938 15802 se
rect -2938 15790 -2876 15802
tri -2876 15790 -2853 15813 nw
tri -2836 15790 -2813 15813 se
rect -2813 15807 -2745 15813
tri -2745 15807 -2723 15829 nw
tri -2705 15807 -2683 15829 se
rect -2683 15807 -2637 15829
rect -2813 15790 -2779 15807
rect -3190 2953 -3138 2965
rect -3190 2264 -3138 2901
rect -3190 2200 -3138 2212
rect -3190 2142 -3138 2148
rect -3350 2042 -3298 2054
rect -3350 1832 -3298 1990
rect -2950 1768 -2898 15790
tri -2898 15768 -2876 15790 nw
tri -2853 15773 -2836 15790 se
rect -2836 15773 -2779 15790
tri -2779 15773 -2745 15807 nw
tri -2739 15773 -2705 15807 se
rect -2705 15801 -2637 15807
tri -2637 15801 -2609 15829 nw
tri -2597 15801 -2569 15829 se
rect -2569 15801 -2529 15829
rect -2705 15773 -2671 15801
tri -2858 15768 -2853 15773 se
rect -2853 15768 -2785 15773
tri -2859 15767 -2858 15768 se
rect -2858 15767 -2785 15768
tri -2785 15767 -2779 15773 nw
tri -2745 15767 -2739 15773 se
rect -2739 15767 -2671 15773
tri -2671 15767 -2637 15801 nw
tri -2631 15767 -2597 15801 se
rect -2597 15795 -2529 15801
tri -2529 15795 -2495 15829 nw
tri -2489 15795 -2455 15829 se
rect -2455 15811 751 15829
tri 751 15811 769 15829 nw
tri 791 15811 809 15829 se
rect 809 15811 831 15829
rect -2455 15795 717 15811
rect -2597 15767 -2563 15795
rect -2950 1704 -2898 1716
rect -2950 1645 -2898 1652
tri -2870 15756 -2859 15767 se
rect -2859 15756 -2796 15767
tri -2796 15756 -2785 15767 nw
tri -2756 15756 -2745 15767 se
rect -2745 15761 -2677 15767
tri -2677 15761 -2671 15767 nw
tri -2637 15761 -2631 15767 se
rect -2631 15761 -2563 15767
tri -2563 15761 -2529 15795 nw
tri -2523 15761 -2489 15795 se
rect -2489 15777 717 15795
tri 717 15777 751 15811 nw
tri 757 15777 791 15811 se
rect 791 15777 831 15811
tri 831 15777 883 15829 nw
rect 2002 15777 2043 15829
tri 2043 15777 2095 15829 nw
tri 10331 15777 10383 15829 ne
rect 10383 15777 11023 15829
rect -2489 15761 -2455 15777
rect -2745 15756 -2683 15761
rect -2870 15755 -2797 15756
tri -2797 15755 -2796 15756 nw
tri -2757 15755 -2756 15756 se
rect -2756 15755 -2683 15756
tri -2683 15755 -2677 15761 nw
tri -2643 15755 -2637 15761 se
rect -2637 15755 -2569 15761
tri -2569 15755 -2563 15761 nw
tri -2529 15755 -2523 15761 se
rect -2523 15755 -2455 15761
tri -2455 15755 -2433 15777 nw
tri 751 15771 757 15777 se
rect 757 15771 825 15777
tri 825 15771 831 15777 nw
rect 2002 15771 2037 15777
tri 2037 15771 2043 15777 nw
tri 10383 15771 10389 15777 ne
rect 10389 15771 11023 15777
tri 735 15755 751 15771 se
rect 751 15755 809 15771
tri 809 15755 825 15771 nw
rect 2002 15755 2021 15771
tri 2021 15755 2037 15771 nw
tri 10389 15755 10405 15771 ne
rect 10405 15755 11023 15771
rect -2870 1623 -2818 15755
tri -2818 15734 -2797 15755 nw
tri -2778 15734 -2757 15755 se
rect -2757 15734 -2710 15755
tri -2790 15722 -2778 15734 se
rect -2778 15728 -2710 15734
tri -2710 15728 -2683 15755 nw
tri -2670 15728 -2643 15755 se
rect -2643 15728 -2603 15755
rect -2778 15722 -2716 15728
tri -2716 15722 -2710 15728 nw
tri -2676 15722 -2670 15728 se
rect -2670 15722 -2603 15728
rect -2790 2241 -2738 15722
tri -2738 15700 -2716 15722 nw
tri -2698 15700 -2676 15722 se
rect -2676 15721 -2603 15722
tri -2603 15721 -2569 15755 nw
tri -2563 15721 -2529 15755 se
rect -2529 15749 -2461 15755
tri -2461 15749 -2455 15755 nw
tri 729 15749 735 15755 se
rect 735 15749 803 15755
tri 803 15749 809 15755 nw
rect 2002 15749 2015 15755
tri 2015 15749 2021 15755 nw
tri 10405 15749 10411 15755 ne
rect 10411 15749 11023 15755
rect -2529 15721 -2495 15749
rect -2676 15700 -2636 15721
tri -2710 15688 -2698 15700 se
rect -2698 15688 -2636 15700
tri -2636 15688 -2603 15721 nw
tri -2596 15688 -2563 15721 se
rect -2563 15715 -2495 15721
tri -2495 15715 -2461 15749 nw
tri -2455 15715 -2421 15749 se
rect -2421 15715 751 15749
rect -2563 15688 -2529 15715
rect -2710 15681 -2643 15688
tri -2643 15681 -2636 15688 nw
tri -2603 15681 -2596 15688 se
rect -2596 15681 -2529 15688
tri -2529 15681 -2495 15715 nw
tri -2489 15681 -2455 15715 se
rect -2455 15697 751 15715
tri 751 15697 803 15749 nw
tri 2002 15736 2015 15749 nw
tri 10411 15736 10424 15749 ne
rect -2455 15681 -2421 15697
rect -2710 2404 -2658 15681
tri -2658 15666 -2643 15681 nw
tri -2618 15666 -2603 15681 se
rect -2603 15675 -2535 15681
tri -2535 15675 -2529 15681 nw
tri -2495 15675 -2489 15681 se
rect -2489 15675 -2421 15681
tri -2421 15675 -2399 15697 nw
rect -2603 15666 -2550 15675
tri -2630 15654 -2618 15666 se
rect -2618 15660 -2550 15666
tri -2550 15660 -2535 15675 nw
tri -2510 15660 -2495 15675 se
rect -2495 15660 -2476 15675
rect -2618 15654 -2556 15660
tri -2556 15654 -2550 15660 nw
tri -2516 15654 -2510 15660 se
rect -2510 15654 -2476 15660
rect -2630 2666 -2578 15654
tri -2578 15632 -2556 15654 nw
tri -2538 15632 -2516 15654 se
rect -2516 15632 -2476 15654
tri -2550 15620 -2538 15632 se
rect -2538 15620 -2476 15632
tri -2476 15620 -2421 15675 nw
rect -2550 14329 -2498 15620
tri -2498 15598 -2476 15620 nw
tri -2187 8512 -2162 8537 ne
tri 10222 8277 10424 8479 se
rect 10424 8385 11023 15749
tri 11023 15735 11159 15871 nw
tri 13646 15736 13781 15871 ne
rect 13781 15736 13983 15871
tri 13983 15736 14125 15878 nw
tri 14539 15736 14681 15878 ne
rect 14681 15736 14882 15878
tri 14681 15735 14682 15736 ne
rect 14682 15735 14882 15736
tri 14682 15734 14683 15735 ne
rect 14683 15734 14882 15735
tri 14882 15734 15026 15878 nw
tri 15443 15736 15585 15878 ne
rect 15585 15736 15787 15878
tri 15787 15736 15929 15878 nw
tri 16315 15736 16457 15878 ne
rect 16457 15736 17079 15878
tri 16457 15734 16459 15736 ne
rect 16459 15734 17079 15736
tri 16459 15669 16524 15734 ne
rect 16524 15669 17079 15734
tri 11023 8385 11133 8495 sw
rect 10424 8277 11133 8385
tri 11133 8277 11241 8385 sw
tri 16635 8277 16743 8385 se
rect 16743 8277 17079 15669
rect 1940 7561 16555 8277
tri 16595 8237 16635 8277 se
rect 16635 8237 17079 8277
rect 1940 7418 2207 7561
tri 2207 7418 2350 7561 nw
tri 2858 7418 3001 7561 ne
rect 3001 7418 4015 7561
tri 4015 7418 4158 7561 nw
tri 4666 7418 4809 7561 ne
rect 4809 7418 5815 7561
tri 5815 7418 5958 7561 nw
tri 6466 7418 6609 7561 ne
rect 6609 7418 7622 7561
tri 7622 7418 7765 7561 nw
tri 8273 7418 8416 7561 ne
rect 8416 7418 9423 7561
tri 9423 7418 9566 7561 nw
tri 10074 7418 10217 7561 ne
rect 10217 7418 11233 7561
tri 11233 7418 11376 7561 nw
tri 11884 7418 12027 7561 ne
rect 12027 7418 13034 7561
tri 13034 7418 13177 7561 nw
tri 13685 7418 13828 7561 ne
rect 13828 7418 14833 7561
tri 14833 7418 14976 7561 nw
tri 15484 7418 15627 7561 ne
rect 15627 7418 16555 7561
rect 1940 7394 2183 7418
tri 2183 7394 2207 7418 nw
tri 3001 7394 3025 7418 ne
rect 1940 6975 2156 7394
tri 2156 7367 2183 7394 nw
tri 2156 6975 2173 6992 sw
tri 3008 6975 3025 6992 se
rect 3025 6975 4015 7418
tri 4809 7394 4833 7418 ne
tri 4808 6975 4833 7000 se
rect 4833 6975 5815 7418
tri 6609 7394 6633 7418 ne
tri 6608 6975 6633 7000 se
rect 6633 6975 7622 7418
tri 8416 7394 8440 7418 ne
tri 8415 6975 8440 7000 se
rect 8440 6975 9423 7418
tri 10217 7394 10241 7418 ne
tri 10216 6975 10241 7000 se
rect 10241 6975 11233 7418
tri 12027 7394 12051 7418 ne
tri 12026 6975 12051 7000 se
rect 12051 6975 13034 7418
tri 13828 7394 13852 7418 ne
tri 13827 6975 13852 7000 se
rect 13852 6975 14833 7418
tri 15627 7394 15651 7418 ne
tri 15626 6975 15651 7000 se
rect 15651 6975 16555 7418
rect 1940 6833 2173 6975
tri 2173 6833 2315 6975 sw
tri 2866 6833 3008 6975 se
rect 3008 6833 4015 6975
tri 4015 6833 4157 6975 sw
tri 4666 6833 4808 6975 se
rect 4808 6833 5815 6975
tri 5815 6833 5957 6975 sw
tri 6466 6833 6608 6975 se
rect 6608 6833 7622 6975
tri 7622 6833 7764 6975 sw
tri 8273 6833 8415 6975 se
rect 8415 6833 9423 6975
tri 9423 6833 9565 6975 sw
tri 10074 6833 10216 6975 se
rect 10216 6833 11233 6975
tri 11233 6833 11375 6975 sw
tri 11884 6833 12026 6975 se
rect 12026 6833 13034 6975
tri 13034 6833 13176 6975 sw
tri 13685 6833 13827 6975 se
rect 13827 6833 14833 6975
tri 14833 6833 14975 6975 sw
tri 15484 6833 15626 6975 se
rect 15626 6833 16555 6975
rect 1940 6670 16555 6833
rect 1940 6630 14073 6670
tri 14073 6630 14113 6670 nw
tri 14528 6630 14568 6670 ne
rect 14568 6630 15719 6670
tri 1910 6478 2062 6630 ne
rect 2062 6478 3097 6630
tri 3097 6480 3247 6630 nw
tri 3748 6480 3898 6630 ne
rect 3898 6480 4899 6630
tri 3898 6478 3900 6480 ne
tri 2062 6442 2098 6478 ne
rect 1414 6025 1630 6370
rect 1658 3438 1938 6112
rect -2550 3398 -2498 3432
rect 2098 3398 3097 6478
rect 3206 3438 3750 6370
rect 3900 3681 4899 6480
tri 4899 6478 5051 6630 nw
tri 5565 6478 5717 6630 ne
rect 5717 6478 6697 6630
tri 6697 6478 6849 6630 nw
tri 7352 6625 7357 6630 ne
rect 7357 6625 8654 6630
tri 7357 6620 7362 6625 ne
rect 7362 6624 8654 6625
tri 8654 6624 8660 6630 nw
tri 9162 6624 9168 6630 ne
rect 9168 6624 10313 6630
rect 7362 6620 8648 6624
tri 7362 6615 7367 6620 ne
rect 7367 6618 8648 6620
tri 8648 6618 8654 6624 nw
tri 9168 6618 9174 6624 ne
rect 9174 6618 10313 6624
rect 7367 6615 8642 6618
tri 7367 6610 7372 6615 ne
rect 7372 6612 8642 6615
tri 8642 6612 8648 6618 nw
tri 9174 6612 9180 6618 ne
rect 9180 6612 10313 6618
rect 7372 6610 8636 6612
tri 7372 6605 7377 6610 ne
rect 7377 6606 8636 6610
tri 8636 6606 8642 6612 nw
tri 9180 6606 9186 6612 ne
rect 9186 6606 10313 6612
rect 7377 6605 8630 6606
tri 7377 6600 7382 6605 ne
rect 7382 6600 8630 6605
tri 8630 6600 8636 6606 nw
tri 9186 6600 9192 6606 ne
rect 9192 6600 10313 6606
tri 7382 6595 7387 6600 ne
rect 7387 6595 8624 6600
tri 7387 6590 7392 6595 ne
rect 7392 6594 8624 6595
tri 8624 6594 8630 6600 nw
tri 9192 6594 9198 6600 ne
rect 9198 6594 10313 6600
rect 7392 6590 8618 6594
tri 7392 6585 7397 6590 ne
rect 7397 6588 8618 6590
tri 8618 6588 8624 6594 nw
tri 9198 6588 9204 6594 ne
rect 9204 6588 10313 6594
rect 7397 6585 8612 6588
tri 7397 6580 7402 6585 ne
rect 7402 6582 8612 6585
tri 8612 6582 8618 6588 nw
tri 9204 6582 9210 6588 ne
rect 9210 6582 10313 6588
rect 7402 6580 8606 6582
tri 7402 6575 7407 6580 ne
rect 7407 6576 8606 6580
tri 8606 6576 8612 6582 nw
tri 9210 6576 9216 6582 ne
rect 9216 6576 10313 6582
rect 7407 6575 8600 6576
tri 7407 6570 7412 6575 ne
rect 7412 6570 8600 6575
tri 8600 6570 8606 6576 nw
tri 9216 6570 9222 6576 ne
rect 9222 6570 10313 6576
tri 7412 6565 7417 6570 ne
rect 7417 6565 8594 6570
tri 7417 6560 7422 6565 ne
rect 7422 6564 8594 6565
tri 8594 6564 8600 6570 nw
tri 9222 6564 9228 6570 ne
rect 9228 6564 10313 6570
rect 7422 6560 8588 6564
tri 7422 6555 7427 6560 ne
rect 7427 6558 8588 6560
tri 8588 6558 8594 6564 nw
tri 9228 6558 9234 6564 ne
rect 9234 6558 10313 6564
rect 7427 6556 8586 6558
tri 8586 6556 8588 6558 nw
tri 9234 6556 9236 6558 ne
rect 9236 6556 10313 6558
rect 7427 6555 8580 6556
tri 7427 6553 7429 6555 ne
rect 7429 6553 8580 6555
tri 7429 6548 7434 6553 ne
rect 7434 6550 8580 6553
tri 8580 6550 8586 6556 nw
tri 9236 6550 9242 6556 ne
rect 9242 6550 10313 6556
rect 7434 6548 8574 6550
tri 7434 6543 7439 6548 ne
rect 7439 6544 8574 6548
tri 8574 6544 8580 6550 nw
tri 9242 6544 9248 6550 ne
rect 9248 6544 10313 6550
rect 7439 6543 8568 6544
tri 7439 6538 7444 6543 ne
rect 7444 6538 8568 6543
tri 8568 6538 8574 6544 nw
tri 9248 6538 9254 6544 ne
rect 9254 6538 10313 6544
tri 7444 6533 7449 6538 ne
rect 7449 6533 8562 6538
tri 7449 6528 7454 6533 ne
rect 7454 6532 8562 6533
tri 8562 6532 8568 6538 nw
tri 9254 6532 9260 6538 ne
rect 9260 6532 10313 6538
rect 7454 6528 8556 6532
tri 7454 6523 7459 6528 ne
rect 7459 6526 8556 6528
tri 8556 6526 8562 6532 nw
tri 9260 6526 9266 6532 ne
rect 9266 6526 10313 6532
rect 7459 6523 8550 6526
tri 7459 6518 7464 6523 ne
rect 7464 6520 8550 6523
tri 8550 6520 8556 6526 nw
tri 9266 6520 9272 6526 ne
rect 9272 6520 10313 6526
rect 7464 6518 8544 6520
tri 7464 6513 7469 6518 ne
rect 7469 6514 8544 6518
tri 8544 6514 8550 6520 nw
tri 9272 6514 9278 6520 ne
rect 9278 6514 10313 6520
rect 7469 6513 8538 6514
tri 7469 6508 7474 6513 ne
rect 7474 6508 8538 6513
tri 8538 6508 8544 6514 nw
tri 9278 6508 9284 6514 ne
rect 9284 6508 10313 6514
tri 7474 6503 7479 6508 ne
rect 7479 6503 8532 6508
tri 7479 6498 7484 6503 ne
rect 7484 6502 8532 6503
tri 8532 6502 8538 6508 nw
tri 9284 6502 9290 6508 ne
rect 9290 6502 10313 6508
rect 7484 6498 8526 6502
tri 7484 6493 7489 6498 ne
rect 7489 6496 8526 6498
tri 8526 6496 8532 6502 nw
tri 9290 6496 9296 6502 ne
rect 9296 6496 10313 6502
rect 7489 6493 8520 6496
tri 7489 6488 7494 6493 ne
rect 7494 6490 8520 6493
tri 8520 6490 8526 6496 nw
tri 9296 6490 9302 6496 ne
rect 9302 6490 10313 6496
rect 7494 6488 8514 6490
tri 7494 6483 7499 6488 ne
rect 7499 6484 8514 6488
tri 8514 6484 8520 6490 nw
tri 9302 6484 9308 6490 ne
rect 9308 6484 10313 6490
rect 7499 6483 8508 6484
tri 7499 6478 7504 6483 ne
tri 5717 6420 5775 6478 ne
rect 3900 3629 3906 3681
rect 3958 3629 3973 3681
rect 4025 3629 4040 3681
rect 4092 3629 4107 3681
rect 4159 3629 4174 3681
rect 4226 3629 4240 3681
rect 4292 3629 4306 3681
rect 4358 3629 4372 3681
rect 4424 3629 4438 3681
rect 4490 3629 4504 3681
rect 4556 3629 4570 3681
rect 4622 3629 4636 3681
rect 4688 3629 4702 3681
rect 4754 3629 4768 3681
rect 4820 3629 4834 3681
rect 4886 3629 4899 3681
rect 3900 3617 4899 3629
rect 3900 3565 3906 3617
rect 3958 3565 3973 3617
rect 4025 3565 4040 3617
rect 4092 3565 4107 3617
rect 4159 3565 4174 3617
rect 4226 3565 4240 3617
rect 4292 3565 4306 3617
rect 4358 3565 4372 3617
rect 4424 3565 4438 3617
rect 4490 3565 4504 3617
rect 4556 3565 4570 3617
rect 4622 3565 4636 3617
rect 4688 3565 4702 3617
rect 4754 3565 4768 3617
rect 4820 3565 4834 3617
rect 4886 3565 4899 3617
rect 3900 3398 4899 3565
rect 5010 3398 5610 6370
rect 5775 3682 6697 6478
rect 5775 3630 5781 3682
rect 5833 3630 5847 3682
rect 5899 3630 5913 3682
rect 5965 3630 5979 3682
rect 6031 3630 6045 3682
rect 6097 3630 6111 3682
rect 6163 3630 6177 3682
rect 6229 3630 6243 3682
rect 6295 3630 6309 3682
rect 6361 3630 6375 3682
rect 6427 3630 6441 3682
rect 6493 3630 6507 3682
rect 6559 3630 6573 3682
rect 6625 3630 6639 3682
rect 6691 3630 6697 3682
rect 5775 3618 6697 3630
rect 5775 3566 5781 3618
rect 5833 3566 5847 3618
rect 5899 3566 5913 3618
rect 5965 3566 5979 3618
rect 6031 3566 6045 3618
rect 6097 3566 6111 3618
rect 6163 3566 6177 3618
rect 6229 3566 6243 3618
rect 6295 3566 6309 3618
rect 6361 3566 6375 3618
rect 6427 3566 6441 3618
rect 6493 3566 6507 3618
rect 6559 3566 6573 3618
rect 6625 3566 6639 3618
rect 6691 3566 6697 3618
rect 5775 3398 6697 3566
rect 7504 3682 8508 6483
tri 8508 6478 8514 6484 nw
tri 9308 6478 9314 6484 ne
rect 7504 3630 7510 3682
rect 7562 3630 7577 3682
rect 7629 3630 7644 3682
rect 7696 3630 7711 3682
rect 7763 3630 7778 3682
rect 7830 3630 7845 3682
rect 7897 3630 7912 3682
rect 7964 3630 7979 3682
rect 8031 3630 8046 3682
rect 8098 3630 8113 3682
rect 8165 3630 8180 3682
rect 8232 3630 8246 3682
rect 8298 3630 8312 3682
rect 8364 3630 8378 3682
rect 8430 3630 8444 3682
rect 8496 3630 8508 3682
rect 7504 3618 8508 3630
rect 7504 3566 7510 3618
rect 7562 3566 7577 3618
rect 7629 3566 7644 3618
rect 7696 3566 7711 3618
rect 7763 3566 7778 3618
rect 7830 3566 7845 3618
rect 7897 3566 7912 3618
rect 7964 3566 7979 3618
rect 8031 3566 8046 3618
rect 8098 3566 8113 3618
rect 8165 3566 8180 3618
rect 8232 3566 8246 3618
rect 8298 3566 8312 3618
rect 8364 3566 8378 3618
rect 8430 3566 8444 3618
rect 8496 3566 8508 3618
rect 7504 3560 8508 3566
rect 7504 3558 8502 3560
rect 8618 3398 9218 6370
rect 9314 3681 10313 6484
tri 10313 6478 10465 6630 nw
tri 10965 6478 11117 6630 ne
rect 9314 3629 9322 3681
rect 9374 3629 9389 3681
rect 9441 3629 9456 3681
rect 9508 3629 9523 3681
rect 9575 3629 9590 3681
rect 9642 3629 9656 3681
rect 9708 3629 9722 3681
rect 9774 3629 9788 3681
rect 9840 3629 9854 3681
rect 9906 3629 9920 3681
rect 9972 3629 9986 3681
rect 10038 3629 10052 3681
rect 10104 3629 10118 3681
rect 10170 3629 10184 3681
rect 10236 3629 10250 3681
rect 10302 3629 10313 3681
rect 9314 3617 10313 3629
rect 9314 3565 9322 3617
rect 9374 3565 9389 3617
rect 9441 3565 9456 3617
rect 9508 3565 9523 3617
rect 9575 3565 9590 3617
rect 9642 3565 9656 3617
rect 9708 3565 9722 3617
rect 9774 3565 9788 3617
rect 9840 3565 9854 3617
rect 9906 3565 9920 3617
rect 9972 3565 9986 3617
rect 10038 3565 10052 3617
rect 10104 3565 10118 3617
rect 10170 3565 10184 3617
rect 10236 3565 10250 3617
rect 10302 3565 10313 3617
rect 9314 3398 10313 3565
tri 10421 6194 10597 6370 se
rect 10597 6194 11022 6370
rect 10421 3398 11022 6194
rect 11117 4665 12117 6630
tri 12117 6478 12269 6630 nw
tri 12770 6478 12922 6630 ne
tri 11117 4492 11290 4665 ne
tri 11117 3846 11290 4019 se
rect 11290 3846 12117 4665
rect 12922 4627 13921 6630
tri 13921 6478 14073 6630 nw
tri 14568 6478 14720 6630 ne
rect 12922 4617 13911 4627
tri 13911 4617 13921 4627 nw
tri 12922 4477 13062 4617 ne
rect 11117 3681 12117 3846
rect 11117 3629 11124 3681
rect 11176 3629 11191 3681
rect 11243 3629 11258 3681
rect 11310 3629 11325 3681
rect 11377 3629 11392 3681
rect 11444 3629 11458 3681
rect 11510 3629 11524 3681
rect 11576 3629 11590 3681
rect 11642 3629 11656 3681
rect 11708 3629 11722 3681
rect 11774 3629 11788 3681
rect 11840 3629 11854 3681
rect 11906 3629 11920 3681
rect 11972 3629 11986 3681
rect 12038 3629 12052 3681
rect 12104 3629 12117 3681
rect 11117 3617 12117 3629
rect 11117 3565 11124 3617
rect 11176 3565 11191 3617
rect 11243 3565 11258 3617
rect 11310 3565 11325 3617
rect 11377 3565 11392 3617
rect 11444 3565 11458 3617
rect 11510 3565 11524 3617
rect 11576 3565 11590 3617
rect 11642 3565 11656 3617
rect 11708 3565 11722 3617
rect 11774 3565 11788 3617
rect 11840 3565 11854 3617
rect 11906 3565 11920 3617
rect 11972 3565 11986 3617
rect 12038 3565 12052 3617
rect 12104 3565 12117 3617
rect 11117 3398 12117 3565
tri 12922 3896 13062 4036 se
rect 13062 3896 13776 4617
tri 13776 4482 13911 4617 nw
tri 13776 3896 13905 4025 sw
rect 12922 3880 13905 3896
tri 13905 3880 13921 3896 sw
rect 12922 3681 13921 3880
rect 12922 3629 12928 3681
rect 12980 3629 12995 3681
rect 13047 3629 13062 3681
rect 13114 3629 13129 3681
rect 13181 3629 13196 3681
rect 13248 3629 13262 3681
rect 13314 3629 13328 3681
rect 13380 3629 13394 3681
rect 13446 3629 13460 3681
rect 13512 3629 13526 3681
rect 13578 3629 13592 3681
rect 13644 3629 13658 3681
rect 13710 3629 13724 3681
rect 13776 3629 13790 3681
rect 13842 3629 13856 3681
rect 13908 3629 13921 3681
rect 12922 3617 13921 3629
rect 12922 3565 12928 3617
rect 12980 3565 12995 3617
rect 13047 3565 13062 3617
rect 13114 3565 13129 3617
rect 13181 3565 13196 3617
rect 13248 3565 13262 3617
rect 13314 3565 13328 3617
rect 13380 3565 13394 3617
rect 13446 3565 13460 3617
rect 13512 3565 13526 3617
rect 13578 3565 13592 3617
rect 13644 3565 13658 3617
rect 13710 3565 13724 3617
rect 13776 3565 13790 3617
rect 13842 3565 13856 3617
rect 13908 3565 13921 3617
rect 12411 3438 12633 3512
rect 12922 3398 13921 3565
rect 14029 3398 14629 6370
rect 14720 4620 15719 6630
tri 15719 6478 15911 6670 nw
rect 14720 3681 15573 4620
tri 15573 4474 15719 4620 nw
rect 14720 3629 14726 3681
rect 14778 3629 14792 3681
rect 14844 3629 14858 3681
rect 14910 3629 14924 3681
rect 14976 3629 14990 3681
rect 15042 3629 15055 3681
rect 15107 3629 15120 3681
rect 15172 3629 15185 3681
rect 15237 3629 15250 3681
rect 15302 3629 15315 3681
rect 15367 3629 15380 3681
rect 15432 3629 15445 3681
rect 15497 3629 15510 3681
rect 15562 3629 15573 3681
rect 14720 3617 15573 3629
rect 14720 3565 14726 3617
rect 14778 3565 14792 3617
rect 14844 3565 14858 3617
rect 14910 3565 14924 3617
rect 14976 3565 14990 3617
rect 15042 3565 15055 3617
rect 15107 3565 15120 3617
rect 15172 3565 15185 3617
rect 15237 3565 15250 3617
rect 15302 3565 15315 3617
rect 15367 3565 15380 3617
rect 15432 3565 15445 3617
rect 15497 3565 15510 3617
rect 15562 3565 15573 3617
rect 14720 3398 15573 3565
rect 15632 4379 15656 4431
rect 15708 4379 15720 4431
rect 15772 4379 15778 4431
rect 15632 4345 15693 4379
tri 15693 4345 15727 4379 nw
rect 16412 4345 16418 4397
rect 16470 4345 16482 4397
rect 16534 4345 16654 4397
tri 16654 4345 16706 4397 sw
rect 15632 3398 15690 4345
tri 15690 4342 15693 4345 nw
tri 16602 4342 16605 4345 ne
rect 16605 4342 16706 4345
tri 16706 4342 16709 4345 sw
tri 16605 4296 16651 4342 ne
rect 15718 4253 15770 4259
rect 15718 4189 15770 4201
rect 15718 3828 15770 4137
rect 15718 3764 15770 3776
rect 15718 3706 15770 3712
rect 16327 4219 16333 4271
rect 16385 4219 16397 4271
rect 16449 4219 16455 4271
rect 16019 3438 16241 3512
rect 16327 3455 16385 4219
tri 16385 4189 16415 4219 nw
rect 16415 4173 16467 4179
rect 16415 4109 16467 4121
tri 16467 4103 16495 4131 sw
rect 16467 4071 16591 4103
tri 16591 4071 16623 4103 sw
rect 16467 4057 16623 4071
rect 16415 4051 16623 4057
tri 16540 4026 16565 4051 ne
tri 16385 3455 16470 3540 sw
rect 16327 3422 16470 3455
tri 16327 3398 16351 3422 ne
rect 16351 3398 16470 3422
rect 16565 3398 16623 4051
rect 16651 3969 16709 4342
rect 16651 3828 16709 3834
rect 16651 3776 16654 3828
rect 16706 3776 16709 3828
rect 16651 3764 16709 3776
rect 16651 3712 16654 3764
rect 16706 3712 16709 3764
rect 16651 3398 16709 3712
rect 16791 3398 17111 7366
rect 3206 1818 3623 3398
tri 16351 3337 16412 3398 ne
rect 16412 3337 16470 3398
rect 5168 3229 5174 3281
rect 5226 3229 5240 3281
rect 5292 3229 5306 3281
rect 5358 3229 5372 3281
rect 5424 3229 5438 3281
rect 5490 3229 5503 3281
rect 5555 3229 5568 3281
rect 5620 3229 5633 3281
rect 5685 3229 5691 3281
rect 5168 3185 5691 3229
rect 5168 3133 5174 3185
rect 5226 3133 5240 3185
rect 5292 3133 5306 3185
rect 5358 3133 5372 3185
rect 5424 3133 5438 3185
rect 5490 3133 5503 3185
rect 5555 3133 5568 3185
rect 5620 3133 5633 3185
rect 5685 3133 5691 3185
rect 8522 3229 8528 3281
rect 8580 3229 8594 3281
rect 8646 3229 8660 3281
rect 8712 3229 8726 3281
rect 8778 3229 8792 3281
rect 8844 3229 8857 3281
rect 8909 3229 8922 3281
rect 8974 3229 8980 3281
rect 8522 3215 8980 3229
rect 8522 3163 8528 3215
rect 8580 3163 8594 3215
rect 8646 3163 8660 3215
rect 8712 3163 8726 3215
rect 8778 3163 8792 3215
rect 8844 3163 8857 3215
rect 8909 3163 8922 3215
rect 8974 3163 8980 3215
rect 8181 3017 8187 3069
rect 8239 3017 8251 3069
rect 8303 3017 8309 3069
rect 5005 2937 5011 2989
rect 5063 2937 5075 2989
rect 5127 2937 5133 2989
rect 5005 2200 5133 2937
rect 7714 2937 7720 2989
rect 7772 2937 7784 2989
rect 7836 2937 7842 2989
rect 5214 2745 5220 2797
rect 5272 2745 5286 2797
rect 5338 2745 5351 2797
rect 5403 2745 5416 2797
rect 5468 2745 5481 2797
rect 5533 2745 5546 2797
rect 5598 2745 5611 2797
rect 5663 2745 5676 2797
rect 5728 2745 5741 2797
rect 5793 2745 5806 2797
rect 5858 2745 5871 2797
rect 5923 2745 5936 2797
rect 5988 2745 5994 2797
rect 5214 2703 5994 2745
rect 5214 2651 5220 2703
rect 5272 2651 5286 2703
rect 5338 2651 5351 2703
rect 5403 2651 5416 2703
rect 5468 2651 5481 2703
rect 5533 2651 5546 2703
rect 5598 2651 5611 2703
rect 5663 2651 5676 2703
rect 5728 2651 5741 2703
rect 5793 2651 5806 2703
rect 5858 2651 5871 2703
rect 5923 2651 5936 2703
rect 5988 2651 5994 2703
rect 7714 2280 7842 2937
rect 8411 2745 8417 2797
rect 8469 2745 8482 2797
rect 8534 2745 8547 2797
rect 8599 2745 8612 2797
rect 8664 2745 8677 2797
rect 8729 2745 8741 2797
rect 8793 2745 8805 2797
rect 8857 2745 8863 2797
rect 8411 2703 8863 2745
rect 8411 2651 8417 2703
rect 8469 2651 8482 2703
rect 8534 2651 8547 2703
rect 8599 2651 8612 2703
rect 8664 2651 8677 2703
rect 8729 2651 8741 2703
rect 8793 2651 8805 2703
rect 8857 2651 8863 2703
rect 7714 2228 7720 2280
rect 7772 2228 7784 2280
rect 7836 2228 7842 2280
rect 5005 2148 5011 2200
rect 5063 2148 5075 2200
rect 5127 2148 5133 2200
rect 934 1767 986 1773
rect 3206 1766 3212 1818
rect 3264 1766 3283 1818
rect 3335 1766 3354 1818
rect 3406 1766 3425 1818
rect 3477 1766 3495 1818
rect 3547 1766 3565 1818
rect 3617 1766 3623 1818
rect 3206 1735 3623 1766
rect 934 1703 986 1715
rect 934 1645 986 1651
rect 1014 1675 1066 1681
tri -2818 1623 -2807 1634 sw
rect -2870 1611 -2807 1623
tri -2807 1611 -2795 1623 sw
rect 1014 1611 1066 1623
rect -2870 1608 -2795 1611
tri -2795 1608 -2792 1611 sw
rect -2870 1556 -2864 1608
rect -2812 1556 -2800 1608
rect -2748 1556 -2742 1608
rect 1014 1553 1066 1559
<< metal3 >>
tri 4137 21945 4350 22158 se
rect 4350 21945 5052 22158
rect 4137 21924 5052 21945
rect 4137 21632 4903 21924
tri 4903 21775 5052 21924 nw
rect 5594 21911 6804 22158
rect 5594 21879 6772 21911
tri 6772 21879 6804 21911 nw
rect 7242 21885 8452 22158
tri 7395 21879 7401 21885 ne
rect 7401 21879 8452 21885
tri 5594 21775 5698 21879 ne
rect 5698 21775 6495 21879
rect 4137 21426 4697 21632
tri 4697 21426 4903 21632 nw
tri 5698 21538 5935 21775 ne
rect 5935 21516 6495 21775
tri 6495 21602 6772 21879 nw
tri 7401 21602 7678 21879 ne
rect 7678 21752 8452 21879
rect 8890 21753 10103 22163
rect 7678 21602 8302 21752
tri 8302 21602 8452 21752 nw
tri 9221 21602 9372 21753 ne
rect 9372 21602 10103 21753
tri 7678 21538 7742 21602 ne
rect 7742 21516 8302 21602
tri 9372 21516 9458 21602 ne
rect 9458 21516 10103 21602
tri 9458 21426 9548 21516 ne
rect 9548 21426 10103 21516
tri 9548 21302 9672 21426 ne
rect 9672 21302 10103 21426
rect 11353 21911 12574 22163
rect 11353 21302 11913 21911
tri 11913 21563 12261 21911 nw
rect 13010 21890 14220 22163
rect 14658 21927 17131 22163
rect 14658 21911 15900 21927
tri 15900 21911 15916 21927 nw
tri 14658 21890 14679 21911 ne
rect 14679 21890 15605 21911
rect 13010 21757 13714 21890
tri 13010 21629 13138 21757 ne
rect 13138 21629 13714 21757
tri 13714 21629 13975 21890 nw
tri 14679 21629 14940 21890 ne
rect 14940 21629 15605 21890
tri 13138 21613 13154 21629 ne
rect 13154 21521 13714 21629
tri 14940 21616 14953 21629 ne
rect 14953 21616 15605 21629
tri 15605 21616 15900 21911 nw
rect 14953 21516 15513 21616
tri 15513 21524 15605 21616 nw
tri 530 18875 861 19206 se
rect 861 18875 1322 19206
rect 530 18543 1322 18875
tri 530 18212 861 18543 ne
rect 861 18212 1322 18543
rect 17111 6972 17113 7368
rect -147 278 16368 2138
rect -2317 -3054 16526 -220
<< metal4 >>
rect 8571 22045 8790 22259
rect 8137 6971 8540 7328
rect 15060 6929 17133 7395
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 1 912 -1 0 22498
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 1 686 1 0 2070
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 1 909 1 0 22592
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 879 -1 0 22880
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 1386 -1 0 20279
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 666 -1 0 17945
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 -1 586 -1 0 19236
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 -1 1066 -1 0 19440
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 -1 1226 -1 0 19971
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 -1 -3138 1 0 2142
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 -1 1360 1 0 22321
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 -1 1280 1 0 22413
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 0 -1 1040 1 0 22596
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 0 -1 1040 1 0 22826
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 0 -1 -3138 1 0 2895
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 0 -1 986 1 0 1645
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 0 -1 1066 1 0 1553
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 0 -1 1166 1 0 23120
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform 0 -1 16467 1 0 4051
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform 1 0 1077 0 -1 22880
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1701704242
transform 1 0 1996 0 -1 20279
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1701704242
transform 1 0 1996 0 -1 19911
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1701704242
transform 1 0 1406 0 1 23107
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1701704242
transform 1 0 15650 0 1 4379
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1701704242
transform 1 0 16327 0 1 4219
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1701704242
transform 1 0 16412 0 1 4345
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1701704242
transform 1 0 1994 0 1 18051
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1701704242
transform 1 0 2104 0 1 18977
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1701704242
transform 1 0 1754 0 1 21064
box 0 0 256 116
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform 1 0 1994 0 1 17098
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1701704242
transform 0 1 593 1 0 18533
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1701704242
transform 0 -1 2099 1 0 24113
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1701704242
transform 0 -1 2955 1 0 24113
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_3
timestamp 1701704242
transform 1 0 1466 0 1 23216
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1701704242
transform 0 -1 959 1 0 21546
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1701704242
transform 0 -1 2839 1 0 22478
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1701704242
transform 0 -1 2527 1 0 22478
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1701704242
transform 0 -1 2215 1 0 22478
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_4
timestamp 1701704242
transform 0 -1 906 1 0 18032
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_0
timestamp 1701704242
transform 0 -1 2955 1 0 21952
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_1
timestamp 1701704242
transform 0 -1 2099 1 0 21952
box 0 0 1 1
use M1M2_CDNS_52468879185963  M1M2_CDNS_52468879185963_0
timestamp 1701704242
transform -1 0 3077 0 -1 3681
box 0 0 960 116
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_0
timestamp 1701704242
transform 0 -1 959 1 0 22194
box 0 0 512 52
use M1M2_CDNS_524688791851113  M1M2_CDNS_524688791851113_0
timestamp 1701704242
transform 0 -1 1671 -1 0 24005
box 0 0 1 1
use M1M2_CDNS_524688791851496  M1M2_CDNS_524688791851496_0
timestamp 1701704242
transform 1 0 3625 0 1 21967
box 0 0 768 372
use M1M2_CDNS_524688791851497  M1M2_CDNS_524688791851497_0
timestamp 1701704242
transform 0 -1 1359 -1 0 23998
box 0 0 640 52
use M1M2_CDNS_524688791851498  M1M2_CDNS_524688791851498_0
timestamp 1701704242
transform 0 -1 2527 1 0 23221
box 0 0 768 52
use M1M2_CDNS_524688791851498  M1M2_CDNS_524688791851498_1
timestamp 1701704242
transform 0 -1 2839 1 0 23221
box 0 0 768 52
use M1M2_CDNS_524688791851498  M1M2_CDNS_524688791851498_2
timestamp 1701704242
transform 0 -1 1983 1 0 23216
box 0 0 768 52
use M1M2_CDNS_524688791851499  M1M2_CDNS_524688791851499_0
timestamp 1701704242
transform 0 -1 2215 1 0 23051
box 0 0 896 52
use M1M2_CDNS_524688791851500  M1M2_CDNS_524688791851500_0
timestamp 1701704242
transform 0 1 17066 1 0 16416
box 0 0 768 116
use M2M3_CDNS_524688791851501  M2M3_CDNS_524688791851501_0
timestamp 1701704242
transform 1 0 610 0 1 18508
box -5 0 141 394
use M2M3_CDNS_524688791851502  M2M3_CDNS_524688791851502_0
timestamp 1701704242
transform 1 0 16812 0 1 6972
box -5 0 301 394
use M3M4_CDNS_524688791851495  M3M4_CDNS_524688791851495_0
timestamp 1701704242
transform 1 0 16807 0 1 6972
box -1 0 305 396
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_0
timestamp 1701704242
transform 0 -1 1360 -1 0 1713
box -79 -26 179 626
use nfet_CDNS_52468879185391  nfet_CDNS_52468879185391_0
timestamp 1701704242
transform 0 -1 1360 1 0 1879
box -79 -26 335 626
use pfet_CDNS_52468879185352  pfet_CDNS_52468879185352_0
timestamp 1701704242
transform 0 -1 1970 1 0 22381
box -119 -66 219 1066
use pfet_CDNS_52468879185397  pfet_CDNS_52468879185397_0
timestamp 1701704242
transform 0 -1 1970 1 0 22647
box -119 -66 375 1066
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 1 0 672 0 1 1595
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 1 0 672 0 1 1906
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1701704242
transform 0 1 265 -1 0 18744
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_1
timestamp 1701704242
transform 0 1 265 1 0 16486
box 0 0 1 1
use PYres_CDNS_524688791851556  PYres_CDNS_524688791851556_0
timestamp 1701704242
transform 0 1 234 1 0 16615
box -50 0 2050 400
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1701704242
transform 0 -1 1132 1 0 16480
box 0 0 2270 404
use sky130_fd_io__sio_pddrvr_strong  sky130_fd_io__sio_pddrvr_strong_0
timestamp 1701704242
transform 1 0 2124 0 1 3398
box -5205 -800 15185 20567
use sky130_fd_io__sio_pddrvr_strong_slow  sky130_fd_io__sio_pddrvr_strong_slow_0
timestamp 1701704242
transform 0 1 4217 -1 0 3529
box 0 0 1126 2895
use sky130_fd_io__sio_pddrvr_weak  sky130_fd_io__sio_pddrvr_weak_0
timestamp 1701704242
transform 0 -1 10956 -1 0 3529
box 0 0 1126 4012
use sky130_fd_io__sio_pudrvr_strong  sky130_fd_io__sio_pudrvr_strong_0
timestamp 1701704242
transform 1 0 298 0 1 -1977
box -3494 4163 18774 27929
use sky130_fd_io__sio_pudrvr_strong_slow  sky130_fd_io__sio_pudrvr_strong_slow_0
timestamp 1701704242
transform 1 0 1134 0 -1 25413
box 0 0 1022 2440
use sky130_fd_io__sio_pudrvr_weak  sky130_fd_io__sio_pudrvr_weak_0
timestamp 1701704242
transform -1 0 3012 0 1 21298
box 0 0 1022 3324
use sky130_fd_io__sio_res_weak  sky130_fd_io__sio_res_weak_0
timestamp 1701704242
transform 1 0 456 0 1 16482
box 0 4 1954 4112
use sky130_fd_io__tk_em1o_CDNS_524688791851503  sky130_fd_io__tk_em1o_CDNS_524688791851503_0
timestamp 1701704242
transform 0 1 253 -1 0 17815
box 0 0 1 1
<< labels >>
flabel comment s 2739 3836 2739 3836 0 FreeSans 1000 0 0 0 condiode
flabel comment s 2739 15266 2739 15266 0 FreeSans 1000 0 0 0 condiode
flabel comment s 794 1278 794 1278 0 FreeSans 440 0 0 0 condiode
flabel comment s 7766 3311 7766 3311 0 FreeSans 440 0 0 0 condiode
flabel comment s 4891 3314 4891 3314 0 FreeSans 440 0 0 0 condiode
flabel comment s 1807 3427 1807 3427 0 FreeSans 300 0 0 0 vnb
flabel comment s 797 7187 797 7187 0 FreeSans 200 90 0 0 pd_h<1>
flabel comment s 936 16563 936 16563 0 FreeSans 400 180 0 0 pad_r250
flabel comment s 878 7191 878 7191 0 FreeSans 200 90 0 0 pd_h<0>
flabel comment s 16959 3438 16959 3438 0 FreeSans 300 0 0 0 pad
flabel metal1 s 6097 3022 6149 3056 0 FreeSans 400 0 0 0 pd_h<1>
port 3 nsew
flabel metal1 s 8611 2726 8611 2726 0 FreeSans 440 0 0 0 vgnd_io
flabel metal1 s 697 16478 697 16478 3 FreeSans 200 90 0 0 pad_r250
flabel metal1 s 15598 4131 15656 4188 3 FreeSans 200 180 0 0 pd_h<4>
port 2 nsew
flabel metal1 s 2850 21089 2958 21143 0 FreeSans 200 0 0 0 vgnd
port 4 nsew
flabel metal4 s 8571 22045 8790 22259 0 FreeSans 200 0 0 0 pad
port 5 nsew
flabel metal4 s 8137 6971 8540 7328 0 FreeSans 200 0 0 0 pad
port 5 nsew
flabel metal3 s 914 18586 1133 18800 0 FreeSans 200 0 0 0 pad
port 5 nsew
flabel metal2 s 8193 3026 8245 3060 0 FreeSans 400 0 0 0 pd_h<0>
port 6 nsew
flabel metal2 s -3270 3398 -3218 3432 0 FreeSans 200 90 0 0 pghs_h
port 7 nsew
flabel metal2 s 17561 20546 17871 20586 0 FreeSans 200 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 2188 3398 2370 3472 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 4363 3398 4545 3472 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 6109 3398 6291 3472 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 9706 3398 9888 3472 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 11516 3398 11698 3472 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 15085 3398 15267 3472 0 FreeSans 400 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 16019 3438 16241 3512 0 FreeSans 400 0 0 0 vgnd_io
port 9 nsew
flabel metal2 s 12411 3438 12633 3512 0 FreeSans 400 0 0 0 vgnd_io
port 9 nsew
flabel metal2 s 10607 3438 10829 3512 0 FreeSans 400 0 0 0 vgnd_io
port 9 nsew
flabel metal2 s 8803 3438 9025 3512 0 FreeSans 400 0 0 0 vgnd_io
port 9 nsew
flabel metal2 s 5195 3438 5417 3512 0 FreeSans 400 0 0 0 vgnd_io
port 9 nsew
flabel metal2 s 3391 3438 3613 3512 0 FreeSans 400 0 0 0 vgnd_io
port 9 nsew
flabel metal2 s -2550 3398 -2498 3432 3 FreeSans 200 90 0 0 pug<3>
port 10 nsew
flabel metal2 s -2524 3416 -2524 3416 3 FreeSans 200 90 0 0 pug<3>
flabel metal2 s 16791 3398 17111 3463 0 FreeSans 200 0 0 0 pad
port 5 nsew
flabel metal2 s -2950 3398 -2898 3432 3 FreeSans 200 90 0 0 pu_h_n<1>
port 11 nsew
flabel metal2 s 15632 3398 15690 3455 3 FreeSans 200 90 0 0 pd_h<2>
port 12 nsew
flabel metal2 s 16412 3398 16470 3455 3 FreeSans 200 90 0 0 pd_h<3>
port 13 nsew
flabel metal2 s 17927 20546 18667 20586 0 FreeSans 200 0 0 0 vpb_drvr
port 14 nsew
flabel metal2 s 16565 3398 16623 3456 3 FreeSans 200 90 0 0 tie_lo_esd
port 15 nsew
flabel metal2 s -2710 3398 -2658 3432 3 FreeSans 200 90 0 0 pug<2>
port 16 nsew
flabel metal2 s -2790 3398 -2738 3432 3 FreeSans 200 90 0 0 pu_h_n<2>
port 17 nsew
flabel metal2 s -3190 3398 -3138 3432 3 FreeSans 200 90 0 0 nghs_h
port 18 nsew
flabel metal2 s -2870 3398 -2818 3432 3 FreeSans 200 90 0 0 pug<1>
port 19 nsew
flabel metal2 s -3350 3397 -3298 3431 3 FreeSans 200 90 0 0 pug<0>
port 20 nsew
<< properties >>
string GDS_END 94738568
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94182702
string path 393.600 103.275 393.600 106.475 
<< end >>
