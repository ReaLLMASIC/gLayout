magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -68 -26 1361 126
<< ndiff >>
rect -42 67 0 100
rect -42 33 -34 67
rect -42 0 0 33
rect 1293 67 1335 100
rect 1327 33 1335 67
rect 1293 0 1335 33
<< ndiffc >>
rect -34 33 0 67
rect 1293 33 1327 67
<< ndiffres >>
rect 0 0 1293 100
<< locali >>
rect -34 67 0 83
rect -34 17 0 33
rect 1293 67 1327 83
rect 1293 17 1327 33
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform -1 0 8 0 1 21
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 1 0 1285 0 1 21
box 0 0 1 1
<< properties >>
string GDS_END 79453528
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79453026
<< end >>
