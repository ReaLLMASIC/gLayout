magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 59 1532 865 1568
<< poly >>
rect 178 1548 434 1568
rect 178 1514 233 1548
rect 267 1514 301 1548
rect 335 1514 369 1548
rect 403 1514 434 1548
rect 178 1492 434 1514
rect 490 1548 746 1568
rect 490 1514 526 1548
rect 560 1514 594 1548
rect 628 1514 662 1548
rect 696 1514 746 1548
rect 490 1492 746 1514
rect 117 785 434 840
rect 117 751 137 785
rect 171 751 205 785
rect 239 751 434 785
rect 117 728 434 751
rect 533 785 746 840
rect 533 751 553 785
rect 587 751 621 785
rect 655 751 689 785
rect 723 751 746 785
rect 533 728 746 751
rect 335 54 477 76
rect 335 20 355 54
rect 389 20 423 54
rect 457 20 477 54
rect 335 0 477 20
rect 533 54 677 76
rect 533 20 555 54
rect 589 20 623 54
rect 657 20 677 54
rect 533 0 677 20
<< polycont >>
rect 233 1514 267 1548
rect 301 1514 335 1548
rect 369 1514 403 1548
rect 526 1514 560 1548
rect 594 1514 628 1548
rect 662 1514 696 1548
rect 137 751 171 785
rect 205 751 239 785
rect 553 751 587 785
rect 621 751 655 785
rect 689 751 723 785
rect 355 20 389 54
rect 423 20 457 54
rect 555 20 589 54
rect 623 20 657 54
<< locali >>
rect 217 1514 233 1548
rect 267 1514 301 1548
rect 335 1514 369 1548
rect 403 1514 419 1548
rect 510 1514 526 1548
rect 560 1514 594 1548
rect 628 1514 662 1548
rect 696 1514 712 1548
rect 285 1340 323 1374
rect 183 1142 221 1176
rect 443 1142 481 1176
rect 703 1142 741 1176
rect 601 1018 635 1056
rect 601 946 635 984
rect 121 751 137 785
rect 171 751 205 785
rect 239 751 255 785
rect 289 708 323 928
rect 537 751 553 785
rect 587 751 621 785
rect 655 751 689 785
rect 723 751 739 785
rect 289 674 522 708
rect 488 640 522 674
rect 312 504 346 542
rect 312 432 346 470
rect 664 504 698 542
rect 664 432 698 470
rect 339 20 355 54
rect 389 20 423 54
rect 457 20 473 54
rect 539 20 555 54
rect 589 20 623 54
rect 657 20 673 54
<< viali >>
rect 251 1340 285 1374
rect 323 1340 357 1374
rect 149 1142 183 1176
rect 221 1142 255 1176
rect 409 1142 443 1176
rect 481 1142 515 1176
rect 669 1142 703 1176
rect 741 1142 775 1176
rect 601 1056 635 1090
rect 601 984 635 1018
rect 601 912 635 946
rect 312 542 346 576
rect 312 470 346 504
rect 312 398 346 432
rect 664 542 698 576
rect 664 470 698 504
rect 664 398 698 432
<< metal1 >>
rect 239 1374 369 1380
rect 239 1340 251 1374
rect 285 1340 323 1374
rect 357 1340 369 1374
rect 239 1334 369 1340
rect 137 1176 787 1182
rect 137 1142 149 1176
rect 183 1142 221 1176
rect 255 1142 409 1176
rect 443 1142 481 1176
rect 515 1142 669 1176
rect 703 1142 741 1176
rect 775 1142 787 1176
rect 137 1136 787 1142
rect 0 1090 872 1108
rect 0 1056 601 1090
rect 635 1056 872 1090
rect 0 1018 872 1056
rect 0 984 601 1018
rect 635 984 872 1018
rect 0 946 872 984
rect 0 912 601 946
rect 635 912 872 946
rect 0 906 872 912
rect 0 576 872 582
rect 0 542 312 576
rect 346 542 664 576
rect 698 542 872 576
rect 0 504 872 542
rect 0 470 312 504
rect 346 470 664 504
rect 698 470 872 504
rect 0 432 872 470
rect 0 398 312 432
rect 346 398 664 432
rect 698 398 872 432
rect 0 380 872 398
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 775 0 1 1142
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 515 0 1 1142
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 255 0 1 1142
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 1 0 251 0 1 1340
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1701704242
transform 1 0 601 0 1 912
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1701704242
transform 1 0 664 0 1 398
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1701704242
transform 1 0 312 0 1 398
box 0 0 1 1
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1701704242
transform -1 0 653 0 1 102
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_1
timestamp 1701704242
transform 1 0 357 0 1 102
box -79 -26 199 626
use pfet_CDNS_52468879185368  pfet_CDNS_52468879185368_0
timestamp 1701704242
transform 1 0 178 0 -1 1466
box -119 -66 375 666
use pfet_CDNS_52468879185368  pfet_CDNS_52468879185368_1
timestamp 1701704242
transform 1 0 490 0 -1 1466
box -119 -66 375 666
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 121 1 0 735
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 0 -1 473 1 0 4
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1701704242
transform 0 -1 673 1 0 4
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 1 510 -1 0 1564
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1701704242
transform 0 1 217 1 0 1498
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1701704242
transform 0 1 537 1 0 735
box 0 0 1 1
<< labels >>
flabel comment s 544 1164 544 1164 0 FreeSans 200 0 0 0 int
flabel metal1 s 239 1334 285 1380 7 FreeSans 300 0 0 0 pd_h
port 1 nsew
flabel metal1 s 830 380 872 582 7 FreeSans 300 180 0 0 vgnd_io
port 2 nsew
flabel metal1 s 830 906 872 1108 7 FreeSans 300 180 0 0 vcc_io
port 3 nsew
flabel metal1 s 0 380 42 582 7 FreeSans 300 0 0 0 vgnd_io
port 2 nsew
flabel metal1 s 0 906 42 1108 6 FreeSans 300 0 0 0 vcc_io
port 3 nsew
flabel locali s 705 751 739 785 3 FreeSans 300 180 0 0 pden_h_n
port 5 nsew
flabel locali s 133 751 167 785 3 FreeSans 300 0 0 0 drvlo_h_n
port 6 nsew
<< properties >>
string GDS_END 87996930
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87993748
<< end >>
