magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 319 150
<< mvpmos >>
rect 0 0 200 84
<< mvpdiff >>
rect -53 46 0 84
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 200 46 253 84
rect 200 12 211 46
rect 245 12 253 46
rect 200 0 253 12
<< mvpdiffc >>
rect -45 12 -11 46
rect 211 12 245 46
<< poly >>
rect 0 84 200 116
rect 0 -32 200 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 211 46 245 62
rect 211 -4 245 12
use DFL1sd_CDNS_52468879185322  DFL1sd_CDNS_52468879185322_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185322  DFL1sd_CDNS_52468879185322_1
timestamp 1701704242
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 228 29 228 29 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 7542256
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7541242
<< end >>
