magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -116 -66 13132 1066
<< mvpmos >>
rect 0 0 120 1000
rect 430 0 550 1000
rect 992 0 1112 1000
rect 1422 0 1542 1000
rect 1984 0 2104 1000
rect 2414 0 2534 1000
rect 2976 0 3096 1000
rect 3406 0 3526 1000
rect 3968 0 4088 1000
rect 4398 0 4518 1000
rect 4960 0 5080 1000
rect 5390 0 5510 1000
rect 5952 0 6072 1000
rect 6382 0 6502 1000
rect 6944 0 7064 1000
rect 7374 0 7494 1000
rect 7936 0 8056 1000
rect 8366 0 8486 1000
rect 8928 0 9048 1000
rect 9358 0 9478 1000
rect 9920 0 10040 1000
rect 10350 0 10470 1000
rect 10912 0 11032 1000
rect 11342 0 11462 1000
rect 11904 0 12024 1000
rect 12334 0 12454 1000
rect 12896 0 13016 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 120 0 430 1000
rect 550 0 641 1000
rect 901 0 992 1000
rect 1112 0 1422 1000
rect 1542 0 1633 1000
rect 1893 0 1984 1000
rect 2104 0 2414 1000
rect 2534 0 2625 1000
rect 2885 0 2976 1000
rect 3096 0 3406 1000
rect 3526 0 3617 1000
rect 3877 0 3968 1000
rect 4088 0 4398 1000
rect 4518 0 4609 1000
rect 4869 0 4960 1000
rect 5080 0 5390 1000
rect 5510 0 5601 1000
rect 5861 0 5952 1000
rect 6072 0 6382 1000
rect 6502 0 6593 1000
rect 6853 0 6944 1000
rect 7064 0 7374 1000
rect 7494 0 7585 1000
rect 7845 0 7936 1000
rect 8056 0 8366 1000
rect 8486 0 8577 1000
rect 8837 0 8928 1000
rect 9048 0 9358 1000
rect 9478 0 9569 1000
rect 9829 0 9920 1000
rect 10040 0 10350 1000
rect 10470 0 10561 1000
rect 10821 0 10912 1000
rect 11032 0 11342 1000
rect 11462 0 11553 1000
rect 11813 0 11904 1000
rect 12024 0 12334 1000
rect 12454 0 12545 1000
rect 12805 0 12896 1000
rect 13016 0 13066 1000
<< poly >>
rect 0 1000 120 1032
rect 430 1000 550 1032
rect 992 1000 1112 1032
rect 1422 1000 1542 1032
rect 1984 1000 2104 1032
rect 2414 1000 2534 1032
rect 2976 1000 3096 1032
rect 3406 1000 3526 1032
rect 3968 1000 4088 1032
rect 4398 1000 4518 1032
rect 4960 1000 5080 1032
rect 5390 1000 5510 1032
rect 5952 1000 6072 1032
rect 6382 1000 6502 1032
rect 6944 1000 7064 1032
rect 7374 1000 7494 1032
rect 7936 1000 8056 1032
rect 8366 1000 8486 1032
rect 8928 1000 9048 1032
rect 9358 1000 9478 1032
rect 9920 1000 10040 1032
rect 10350 1000 10470 1032
rect 10912 1000 11032 1032
rect 11342 1000 11462 1032
rect 11904 1000 12024 1032
rect 12334 1000 12454 1032
rect 12896 1000 13016 1032
rect 0 -32 120 0
rect 430 -32 550 0
rect 992 -32 1112 0
rect 1422 -32 1542 0
rect 1984 -32 2104 0
rect 2414 -32 2534 0
rect 2976 -32 3096 0
rect 3406 -32 3526 0
rect 3968 -32 4088 0
rect 4398 -32 4518 0
rect 4960 -32 5080 0
rect 5390 -32 5510 0
rect 5952 -32 6072 0
rect 6382 -32 6502 0
rect 6944 -32 7064 0
rect 7374 -32 7494 0
rect 7936 -32 8056 0
rect 8366 -32 8486 0
rect 8928 -32 9048 0
rect 9358 -32 9478 0
rect 9920 -32 10040 0
rect 10350 -32 10470 0
rect 10912 -32 11032 0
rect 11342 -32 11462 0
rect 11904 -32 12024 0
rect 12334 -32 12454 0
rect 12896 -32 13016 0
<< metal1 >>
rect 748 -16 794 978
rect 1740 -16 1786 978
rect 2732 -16 2778 978
rect 3724 -16 3770 978
rect 4716 -16 4762 978
rect 5708 -16 5754 978
rect 6700 -16 6746 978
rect 7692 -16 7738 978
rect 8684 -16 8730 978
rect 9676 -16 9722 978
rect 10668 -16 10714 978
rect 11660 -16 11706 978
rect 12652 -16 12698 978
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_0
timestamp 1701704242
transform 1 0 12545 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_1
timestamp 1701704242
transform 1 0 11553 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_2
timestamp 1701704242
transform 1 0 10561 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_3
timestamp 1701704242
transform 1 0 9569 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_4
timestamp 1701704242
transform 1 0 8577 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_5
timestamp 1701704242
transform 1 0 7585 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_6
timestamp 1701704242
transform 1 0 6593 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_7
timestamp 1701704242
transform 1 0 5601 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_8
timestamp 1701704242
transform 1 0 4609 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_9
timestamp 1701704242
transform 1 0 3617 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_10
timestamp 1701704242
transform 1 0 2625 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_11
timestamp 1701704242
transform 1 0 1633 0 1 0
box -26 -26 286 1026
use hvDFTPM1s2_CDNS_524688791853  hvDFTPM1s2_CDNS_524688791853_12
timestamp 1701704242
transform 1 0 641 0 1 0
box -26 -26 286 1026
<< labels >>
flabel comment s -25 500 -25 500 0 FreeSans 300 0 0 0 S
flabel comment s 275 500 275 500 0 FreeSans 300 0 0 0 D
flabel comment s 771 481 771 481 0 FreeSans 300 0 0 0 S
flabel comment s 1267 500 1267 500 0 FreeSans 300 0 0 0 D
flabel comment s 1763 481 1763 481 0 FreeSans 300 0 0 0 S
flabel comment s 2259 500 2259 500 0 FreeSans 300 0 0 0 D
flabel comment s 2755 481 2755 481 0 FreeSans 300 0 0 0 S
flabel comment s 3251 500 3251 500 0 FreeSans 300 0 0 0 D
flabel comment s 3747 481 3747 481 0 FreeSans 300 0 0 0 S
flabel comment s 4243 500 4243 500 0 FreeSans 300 0 0 0 D
flabel comment s 4739 481 4739 481 0 FreeSans 300 0 0 0 S
flabel comment s 5235 500 5235 500 0 FreeSans 300 0 0 0 D
flabel comment s 5731 481 5731 481 0 FreeSans 300 0 0 0 S
flabel comment s 6227 500 6227 500 0 FreeSans 300 0 0 0 D
flabel comment s 6723 481 6723 481 0 FreeSans 300 0 0 0 S
flabel comment s 7219 500 7219 500 0 FreeSans 300 0 0 0 D
flabel comment s 7715 481 7715 481 0 FreeSans 300 0 0 0 S
flabel comment s 8211 500 8211 500 0 FreeSans 300 0 0 0 D
flabel comment s 8707 481 8707 481 0 FreeSans 300 0 0 0 S
flabel comment s 9203 500 9203 500 0 FreeSans 300 0 0 0 D
flabel comment s 9699 481 9699 481 0 FreeSans 300 0 0 0 S
flabel comment s 10195 500 10195 500 0 FreeSans 300 0 0 0 D
flabel comment s 10691 481 10691 481 0 FreeSans 300 0 0 0 S
flabel comment s 11187 500 11187 500 0 FreeSans 300 0 0 0 D
flabel comment s 11683 481 11683 481 0 FreeSans 300 0 0 0 S
flabel comment s 12179 500 12179 500 0 FreeSans 300 0 0 0 D
flabel comment s 12675 481 12675 481 0 FreeSans 300 0 0 0 S
flabel comment s 13041 500 13041 500 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 12841834
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 12827962
<< end >>
