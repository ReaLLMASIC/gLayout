magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 1047 326
<< mvnmos >>
rect 0 0 200 300
rect 256 0 456 300
rect 512 0 712 300
rect 768 0 968 300
<< mvndiff >>
rect -53 250 0 300
rect -53 216 -45 250
rect -11 216 0 250
rect -53 182 0 216
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 200 250 256 300
rect 200 216 211 250
rect 245 216 256 250
rect 200 182 256 216
rect 200 148 211 182
rect 245 148 256 182
rect 200 114 256 148
rect 200 80 211 114
rect 245 80 256 114
rect 200 46 256 80
rect 200 12 211 46
rect 245 12 256 46
rect 200 0 256 12
rect 456 250 512 300
rect 456 216 467 250
rect 501 216 512 250
rect 456 182 512 216
rect 456 148 467 182
rect 501 148 512 182
rect 456 114 512 148
rect 456 80 467 114
rect 501 80 512 114
rect 456 46 512 80
rect 456 12 467 46
rect 501 12 512 46
rect 456 0 512 12
rect 712 250 768 300
rect 712 216 723 250
rect 757 216 768 250
rect 712 182 768 216
rect 712 148 723 182
rect 757 148 768 182
rect 712 114 768 148
rect 712 80 723 114
rect 757 80 768 114
rect 712 46 768 80
rect 712 12 723 46
rect 757 12 768 46
rect 712 0 768 12
rect 968 250 1021 300
rect 968 216 979 250
rect 1013 216 1021 250
rect 968 182 1021 216
rect 968 148 979 182
rect 1013 148 1021 182
rect 968 114 1021 148
rect 968 80 979 114
rect 1013 80 1021 114
rect 968 46 1021 80
rect 968 12 979 46
rect 1013 12 1021 46
rect 968 0 1021 12
<< mvndiffc >>
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 211 216 245 250
rect 211 148 245 182
rect 211 80 245 114
rect 211 12 245 46
rect 467 216 501 250
rect 467 148 501 182
rect 467 80 501 114
rect 467 12 501 46
rect 723 216 757 250
rect 723 148 757 182
rect 723 80 757 114
rect 723 12 757 46
rect 979 216 1013 250
rect 979 148 1013 182
rect 979 80 1013 114
rect 979 12 1013 46
<< poly >>
rect 0 300 200 326
rect 256 300 456 326
rect 512 300 712 326
rect 768 300 968 326
rect 0 -26 200 0
rect 256 -26 456 0
rect 512 -26 712 0
rect 768 -26 968 0
<< locali >>
rect -45 250 -11 266
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 211 250 245 266
rect 211 182 245 216
rect 211 114 245 148
rect 211 46 245 80
rect 211 -4 245 12
rect 467 250 501 266
rect 467 182 501 216
rect 467 114 501 148
rect 467 46 501 80
rect 467 -4 501 12
rect 723 250 757 266
rect 723 182 757 216
rect 723 114 757 148
rect 723 46 757 80
rect 723 -4 757 12
rect 979 250 1013 266
rect 979 182 1013 216
rect 979 114 1013 148
rect 979 46 1013 80
rect 979 -4 1013 12
use hvDFL1sd2_CDNS_52468879185238  hvDFL1sd2_CDNS_52468879185238_0
timestamp 1701704242
transform 1 0 712 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185238  hvDFL1sd2_CDNS_52468879185238_1
timestamp 1701704242
transform 1 0 456 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185238  hvDFL1sd2_CDNS_52468879185238_2
timestamp 1701704242
transform 1 0 200 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185376  hvDFL1sd_CDNS_52468879185376_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185376  hvDFL1sd_CDNS_52468879185376_1
timestamp 1701704242
transform 1 0 968 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
flabel comment s 228 131 228 131 0 FreeSans 300 0 0 0 D
flabel comment s 484 131 484 131 0 FreeSans 300 0 0 0 S
flabel comment s 740 131 740 131 0 FreeSans 300 0 0 0 D
flabel comment s 996 131 996 131 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 97993312
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97990922
<< end >>
