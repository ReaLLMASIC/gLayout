magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -91 3928 83 4014
rect 2203 3928 2377 4014
rect -91 3631 2377 3928
rect 117 3109 2169 3631
rect 117 2023 2425 3109
rect 117 819 2169 2023
rect 117 59 2425 819
rect 2203 -27 2425 59
<< mvnnmos >>
tri 143 3557 163 3577 sw
tri 2123 3557 2143 3577 se
rect 143 3157 2143 3557
tri 143 3137 163 3157 nw
tri 2123 3137 2143 3157 ne
tri 143 1975 163 1995 sw
tri 2123 1975 2143 1995 se
rect 143 1575 2143 1975
tri 143 1555 163 1575 nw
tri 2123 1555 2143 1575 ne
tri 143 1267 163 1287 sw
tri 2123 1267 2143 1287 se
rect 143 1195 2143 1267
<< nmoslvt >>
rect 143 867 2143 1195
tri 143 847 163 867 nw
tri 2123 847 2143 867 ne
<< ndiff >>
rect 143 3762 2143 3902
rect 143 3660 242 3762
rect 1976 3660 2143 3762
rect 143 3654 2143 3660
tri 143 847 163 867 se
rect 163 847 2123 867
tri 2123 847 2143 867 sw
rect 143 327 2143 847
rect 143 225 242 327
rect 1976 225 2143 327
rect 143 85 2143 225
<< mvndiff >>
rect 143 3577 2143 3654
tri 143 3557 163 3577 ne
rect 163 3557 2123 3577
tri 2123 3557 2143 3577 nw
tri 143 3137 163 3157 se
rect 163 3137 2123 3157
tri 2123 3137 2143 3157 sw
rect 143 2617 2143 3137
rect 143 2515 242 2617
rect 1976 2515 2143 2617
rect 143 1995 2143 2515
tri 143 1975 163 1995 ne
rect 163 1975 2123 1995
tri 2123 1975 2143 1995 nw
tri 143 1555 163 1575 se
rect 163 1555 2123 1575
tri 2123 1555 2143 1575 sw
rect 143 1472 2143 1555
rect 143 1370 242 1472
rect 1976 1370 2143 1472
rect 143 1287 2143 1370
tri 143 1267 163 1287 ne
rect 163 1267 2123 1287
tri 2123 1267 2143 1287 nw
<< ndiffc >>
rect 242 3660 1976 3762
rect 242 225 1976 327
<< mvndiffc >>
rect 242 2515 1976 2617
rect 242 1370 1976 1472
<< psubdiff >>
rect -65 3936 57 3988
rect -65 3902 -45 3936
rect -11 3902 23 3936
rect 2229 3936 2351 3988
rect 2263 3902 2297 3936
rect 2331 3902 2351 3936
rect -65 3862 57 3902
rect -65 3828 -45 3862
rect -11 3828 23 3862
rect -65 3788 57 3828
rect -65 3754 -45 3788
rect -11 3754 23 3788
rect -65 3715 57 3754
rect -65 3681 -45 3715
rect -11 3681 23 3715
rect -65 3657 57 3681
rect 2229 3862 2351 3902
rect 2263 3828 2297 3862
rect 2331 3828 2351 3862
rect 2229 3788 2351 3828
rect 2263 3754 2297 3788
rect 2331 3754 2351 3788
rect 2229 3715 2351 3754
rect 2263 3681 2297 3715
rect 2331 3681 2351 3715
rect 2229 3657 2351 3681
rect 2229 3059 2399 3083
rect 2229 2049 2399 2073
rect 2229 769 2399 793
rect 2263 735 2297 769
rect 2331 735 2365 769
rect 2229 699 2399 735
rect 2263 665 2297 699
rect 2331 665 2365 699
rect 2229 629 2399 665
rect 2263 595 2297 629
rect 2331 595 2365 629
rect 2229 559 2399 595
rect 2263 525 2297 559
rect 2331 525 2365 559
rect 2229 489 2399 525
rect 2263 455 2297 489
rect 2331 455 2365 489
rect 2229 419 2399 455
rect 2263 385 2297 419
rect 2331 385 2365 419
rect 2229 349 2399 385
rect 2263 315 2297 349
rect 2331 315 2365 349
rect 2229 279 2399 315
rect 2263 245 2297 279
rect 2331 245 2365 279
rect 2229 209 2399 245
rect 2263 175 2297 209
rect 2331 175 2365 209
rect 2229 138 2399 175
rect 2263 104 2297 138
rect 2331 104 2365 138
rect 2229 67 2399 104
rect 2263 33 2297 67
rect 2331 33 2365 67
rect 2229 -1 2399 33
<< psubdiffcont >>
rect -45 3902 -11 3936
rect 23 3902 57 3936
rect 2229 3902 2263 3936
rect 2297 3902 2331 3936
rect -45 3828 -11 3862
rect 23 3828 57 3862
rect -45 3754 -11 3788
rect 23 3754 57 3788
rect -45 3681 -11 3715
rect 23 3681 57 3715
rect 2229 3828 2263 3862
rect 2297 3828 2331 3862
rect 2229 3754 2263 3788
rect 2297 3754 2331 3788
rect 2229 3681 2263 3715
rect 2297 3681 2331 3715
rect 2229 2073 2399 3059
rect 2229 735 2263 769
rect 2297 735 2331 769
rect 2365 735 2399 769
rect 2229 665 2263 699
rect 2297 665 2331 699
rect 2365 665 2399 699
rect 2229 595 2263 629
rect 2297 595 2331 629
rect 2365 595 2399 629
rect 2229 525 2263 559
rect 2297 525 2331 559
rect 2365 525 2399 559
rect 2229 455 2263 489
rect 2297 455 2331 489
rect 2365 455 2399 489
rect 2229 385 2263 419
rect 2297 385 2331 419
rect 2365 385 2399 419
rect 2229 315 2263 349
rect 2297 315 2331 349
rect 2365 315 2399 349
rect 2229 245 2263 279
rect 2297 245 2331 279
rect 2365 245 2399 279
rect 2229 175 2263 209
rect 2297 175 2331 209
rect 2365 175 2399 209
rect 2229 104 2263 138
rect 2297 104 2331 138
rect 2365 104 2399 138
rect 2229 33 2263 67
rect 2297 33 2331 67
rect 2365 33 2399 67
<< poly >>
rect -61 3581 123 3597
rect -61 3547 -45 3581
rect -11 3577 123 3581
tri 123 3577 143 3597 sw
tri 2143 3577 2163 3597 se
rect 2163 3581 2347 3597
rect 2163 3577 2297 3581
rect -11 3547 143 3577
rect -61 3512 143 3547
rect -61 3478 -45 3512
rect -11 3478 143 3512
rect -61 3443 143 3478
rect -61 3409 -45 3443
rect -11 3409 143 3443
rect -61 3374 143 3409
rect -61 3340 -45 3374
rect -11 3340 143 3374
rect -61 3305 143 3340
rect -61 3271 -45 3305
rect -11 3271 143 3305
rect -61 3236 143 3271
rect -61 3202 -45 3236
rect -11 3202 143 3236
rect -61 3167 143 3202
rect -61 3133 -45 3167
rect -11 3137 143 3167
rect 2143 3547 2297 3577
rect 2331 3547 2347 3581
rect 2143 3512 2347 3547
rect 2143 3478 2297 3512
rect 2331 3478 2347 3512
rect 2143 3443 2347 3478
rect 2143 3409 2297 3443
rect 2331 3409 2347 3443
rect 2143 3374 2347 3409
rect 2143 3340 2297 3374
rect 2331 3340 2347 3374
rect 2143 3305 2347 3340
rect 2143 3271 2297 3305
rect 2331 3271 2347 3305
rect 2143 3236 2347 3271
rect 2143 3202 2297 3236
rect 2331 3202 2347 3236
rect 2143 3167 2347 3202
rect 2143 3137 2297 3167
rect -11 3133 123 3137
rect -61 3117 123 3133
tri 123 3117 143 3137 nw
tri 2143 3117 2163 3137 ne
rect 2163 3133 2297 3137
rect 2331 3133 2347 3167
rect 2163 3117 2347 3133
rect -61 1999 123 2015
rect -61 1965 -45 1999
rect -11 1995 123 1999
tri 123 1995 143 2015 sw
tri 2143 1995 2163 2015 se
rect 2163 1999 2347 2015
rect 2163 1995 2297 1999
rect -11 1965 143 1995
rect -61 1930 143 1965
rect -61 1896 -45 1930
rect -11 1896 143 1930
rect -61 1861 143 1896
rect -61 1827 -45 1861
rect -11 1827 143 1861
rect -61 1792 143 1827
rect -61 1758 -45 1792
rect -11 1758 143 1792
rect -61 1723 143 1758
rect -61 1689 -45 1723
rect -11 1689 143 1723
rect -61 1654 143 1689
rect -61 1620 -45 1654
rect -11 1620 143 1654
rect -61 1585 143 1620
rect -61 1551 -45 1585
rect -11 1555 143 1585
rect 2143 1965 2297 1995
rect 2331 1965 2347 1999
rect 2143 1930 2347 1965
rect 2143 1896 2297 1930
rect 2331 1896 2347 1930
rect 2143 1861 2347 1896
rect 2143 1827 2297 1861
rect 2331 1827 2347 1861
rect 2143 1792 2347 1827
rect 2143 1758 2297 1792
rect 2331 1758 2347 1792
rect 2143 1723 2347 1758
rect 2143 1689 2297 1723
rect 2331 1689 2347 1723
rect 2143 1654 2347 1689
rect 2143 1620 2297 1654
rect 2331 1620 2347 1654
rect 2143 1585 2347 1620
rect 2143 1555 2297 1585
rect -11 1551 123 1555
rect -61 1535 123 1551
tri 123 1535 143 1555 nw
tri 2143 1535 2163 1555 ne
rect 2163 1551 2297 1555
rect 2331 1551 2347 1585
rect 2163 1535 2347 1551
rect -61 1291 123 1307
rect -61 1257 -45 1291
rect -11 1287 123 1291
tri 123 1287 143 1307 sw
tri 2143 1287 2163 1307 se
rect 2163 1291 2347 1307
rect 2163 1287 2297 1291
rect -11 1257 143 1287
rect -61 1222 143 1257
rect -61 1188 -45 1222
rect -11 1188 143 1222
rect 2143 1257 2297 1287
rect 2331 1257 2347 1291
rect 2143 1222 2347 1257
rect -61 1153 143 1188
rect -61 1119 -45 1153
rect -11 1119 143 1153
rect -61 1084 143 1119
rect -61 1050 -45 1084
rect -11 1050 143 1084
rect -61 1015 143 1050
rect -61 981 -45 1015
rect -11 981 143 1015
rect -61 946 143 981
rect -61 912 -45 946
rect -11 912 143 946
rect -61 877 143 912
rect -61 843 -45 877
rect -11 847 143 877
rect 2143 1188 2297 1222
rect 2331 1188 2347 1222
rect 2143 1153 2347 1188
rect 2143 1119 2297 1153
rect 2331 1119 2347 1153
rect 2143 1084 2347 1119
rect 2143 1050 2297 1084
rect 2331 1050 2347 1084
rect 2143 1015 2347 1050
rect 2143 981 2297 1015
rect 2331 981 2347 1015
rect 2143 946 2347 981
rect 2143 912 2297 946
rect 2331 912 2347 946
rect 2143 877 2347 912
rect 2143 847 2297 877
rect -11 843 123 847
rect -61 827 123 843
tri 123 827 143 847 nw
tri 2143 827 2163 847 ne
rect 2163 843 2297 847
rect 2331 843 2347 877
rect 2163 827 2347 843
<< polycont >>
rect -45 3547 -11 3581
rect -45 3478 -11 3512
rect -45 3409 -11 3443
rect -45 3340 -11 3374
rect -45 3271 -11 3305
rect -45 3202 -11 3236
rect -45 3133 -11 3167
rect 2297 3547 2331 3581
rect 2297 3478 2331 3512
rect 2297 3409 2331 3443
rect 2297 3340 2331 3374
rect 2297 3271 2331 3305
rect 2297 3202 2331 3236
rect 2297 3133 2331 3167
rect -45 1965 -11 1999
rect -45 1896 -11 1930
rect -45 1827 -11 1861
rect -45 1758 -11 1792
rect -45 1689 -11 1723
rect -45 1620 -11 1654
rect -45 1551 -11 1585
rect 2297 1965 2331 1999
rect 2297 1896 2331 1930
rect 2297 1827 2331 1861
rect 2297 1758 2331 1792
rect 2297 1689 2331 1723
rect 2297 1620 2331 1654
rect 2297 1551 2331 1585
rect -45 1257 -11 1291
rect -45 1188 -11 1222
rect 2297 1257 2331 1291
rect -45 1119 -11 1153
rect -45 1050 -11 1084
rect -45 981 -11 1015
rect -45 912 -11 946
rect -45 843 -11 877
rect 2297 1188 2331 1222
rect 2297 1119 2331 1153
rect 2297 1050 2331 1084
rect 2297 981 2331 1015
rect 2297 912 2331 946
rect 2297 843 2331 877
<< locali >>
rect -65 3936 57 3988
rect -65 3902 -45 3936
rect -11 3902 23 3936
rect 2229 3936 2351 3988
rect 2263 3902 2297 3936
rect 2331 3902 2351 3936
rect -65 3862 57 3902
rect -65 3828 -45 3862
rect -11 3828 23 3862
rect -65 3788 57 3828
rect -65 3754 -45 3788
rect -11 3754 23 3788
rect -65 3715 57 3754
rect -65 3681 -45 3715
rect -11 3681 23 3715
rect -65 3657 57 3681
rect 143 3764 2143 3902
rect 143 3658 242 3764
rect 276 3762 315 3764
rect 349 3762 388 3764
rect 422 3762 461 3764
rect 495 3762 534 3764
rect 568 3762 607 3764
rect 641 3762 680 3764
rect 714 3762 753 3764
rect 787 3762 826 3764
rect 860 3762 900 3764
rect 934 3762 974 3764
rect 1008 3762 1048 3764
rect 1082 3762 1122 3764
rect 1156 3762 1196 3764
rect 1230 3762 1270 3764
rect 1304 3762 1344 3764
rect 1378 3762 1418 3764
rect 1452 3762 1492 3764
rect 1526 3762 1566 3764
rect 1600 3762 1640 3764
rect 1674 3762 1714 3764
rect 1748 3762 1788 3764
rect 1822 3762 1862 3764
rect 1896 3762 1936 3764
rect 1970 3762 2010 3764
rect 1976 3730 2010 3762
rect 2044 3730 2143 3764
rect 1976 3692 2143 3730
rect 1976 3660 2010 3692
rect 276 3658 315 3660
rect 349 3658 388 3660
rect 422 3658 461 3660
rect 495 3658 534 3660
rect 568 3658 607 3660
rect 641 3658 680 3660
rect 714 3658 753 3660
rect 787 3658 826 3660
rect 860 3658 900 3660
rect 934 3658 974 3660
rect 1008 3658 1048 3660
rect 1082 3658 1122 3660
rect 1156 3658 1196 3660
rect 1230 3658 1270 3660
rect 1304 3658 1344 3660
rect 1378 3658 1418 3660
rect 1452 3658 1492 3660
rect 1526 3658 1566 3660
rect 1600 3658 1640 3660
rect 1674 3658 1714 3660
rect 1748 3658 1788 3660
rect 1822 3658 1862 3660
rect 1896 3658 1936 3660
rect 1970 3658 2010 3660
rect 2044 3658 2143 3692
rect -45 3581 -11 3597
rect -45 3512 -11 3547
rect -45 3443 -11 3478
rect 143 3435 2143 3658
rect 2229 3862 2351 3902
rect 2263 3828 2297 3862
rect 2331 3828 2351 3862
rect 2229 3788 2351 3828
rect 2263 3754 2297 3788
rect 2331 3754 2351 3788
rect 2229 3715 2351 3754
rect 2263 3681 2297 3715
rect 2331 3681 2351 3715
rect 2229 3657 2351 3681
rect 2297 3581 2331 3597
rect 2297 3512 2331 3547
rect 2297 3443 2331 3478
rect -45 3401 -11 3409
rect 2297 3401 2331 3409
rect -45 3374 2331 3401
rect -11 3340 2297 3374
rect -45 3305 2331 3340
rect -11 3271 2297 3305
rect -45 3236 2331 3271
rect -11 3202 2297 3236
rect -45 3167 2331 3202
rect -11 3133 2297 3167
rect -45 3117 2331 3133
rect -45 3059 2399 3083
rect -45 2876 2229 3059
rect 143 2619 2143 2842
rect 143 2513 242 2619
rect 276 2617 315 2619
rect 349 2617 388 2619
rect 422 2617 461 2619
rect 495 2617 534 2619
rect 568 2617 607 2619
rect 641 2617 680 2619
rect 714 2617 753 2619
rect 787 2617 826 2619
rect 860 2617 900 2619
rect 934 2617 974 2619
rect 1008 2617 1048 2619
rect 1082 2617 1122 2619
rect 1156 2617 1196 2619
rect 1230 2617 1270 2619
rect 1304 2617 1344 2619
rect 1378 2617 1418 2619
rect 1452 2617 1492 2619
rect 1526 2617 1566 2619
rect 1600 2617 1640 2619
rect 1674 2617 1714 2619
rect 1748 2617 1788 2619
rect 1822 2617 1862 2619
rect 1896 2617 1936 2619
rect 1970 2617 2010 2619
rect 1976 2585 2010 2617
rect 2044 2585 2143 2619
rect 1976 2547 2143 2585
rect 1976 2515 2010 2547
rect 276 2513 315 2515
rect 349 2513 388 2515
rect 422 2513 461 2515
rect 495 2513 534 2515
rect 568 2513 607 2515
rect 641 2513 680 2515
rect 714 2513 753 2515
rect 787 2513 826 2515
rect 860 2513 900 2515
rect 934 2513 974 2515
rect 1008 2513 1048 2515
rect 1082 2513 1122 2515
rect 1156 2513 1196 2515
rect 1230 2513 1270 2515
rect 1304 2513 1344 2515
rect 1378 2513 1418 2515
rect 1452 2513 1492 2515
rect 1526 2513 1566 2515
rect 1600 2513 1640 2515
rect 1674 2513 1714 2515
rect 1748 2513 1788 2515
rect 1822 2513 1862 2515
rect 1896 2513 1936 2515
rect 1970 2513 2010 2515
rect 2044 2513 2143 2547
rect 143 2290 2143 2513
rect -45 2073 2229 2256
rect -45 2049 2399 2073
rect -45 1999 2331 2015
rect -11 1965 2297 1999
rect -45 1930 2331 1965
rect -11 1896 2297 1930
rect -45 1861 2331 1896
rect -11 1827 2297 1861
rect -45 1792 2331 1827
rect -11 1758 2297 1792
rect -45 1731 2331 1758
rect -45 1723 -11 1731
rect 2297 1723 2331 1731
rect -45 1654 -11 1689
rect -45 1585 -11 1620
rect -45 1535 -11 1551
rect 143 1474 2143 1697
rect 2297 1654 2331 1689
rect 2297 1585 2331 1620
rect 2297 1535 2331 1551
rect 143 1368 242 1474
rect 276 1472 315 1474
rect 349 1472 388 1474
rect 422 1472 461 1474
rect 495 1472 534 1474
rect 568 1472 607 1474
rect 641 1472 680 1474
rect 714 1472 753 1474
rect 787 1472 826 1474
rect 860 1472 900 1474
rect 934 1472 974 1474
rect 1008 1472 1048 1474
rect 1082 1472 1122 1474
rect 1156 1472 1196 1474
rect 1230 1472 1270 1474
rect 1304 1472 1344 1474
rect 1378 1472 1418 1474
rect 1452 1472 1492 1474
rect 1526 1472 1566 1474
rect 1600 1472 1640 1474
rect 1674 1472 1714 1474
rect 1748 1472 1788 1474
rect 1822 1472 1862 1474
rect 1896 1472 1936 1474
rect 1970 1472 2010 1474
rect 1976 1440 2010 1472
rect 2044 1440 2143 1474
rect 1976 1402 2143 1440
rect 1976 1370 2010 1402
rect 276 1368 315 1370
rect 349 1368 388 1370
rect 422 1368 461 1370
rect 495 1368 534 1370
rect 568 1368 607 1370
rect 641 1368 680 1370
rect 714 1368 753 1370
rect 787 1368 826 1370
rect 860 1368 900 1370
rect 934 1368 974 1370
rect 1008 1368 1048 1370
rect 1082 1368 1122 1370
rect 1156 1368 1196 1370
rect 1230 1368 1270 1370
rect 1304 1368 1344 1370
rect 1378 1368 1418 1370
rect 1452 1368 1492 1370
rect 1526 1368 1566 1370
rect 1600 1368 1640 1370
rect 1674 1368 1714 1370
rect 1748 1368 1788 1370
rect 1822 1368 1862 1370
rect 1896 1368 1936 1370
rect 1970 1368 2010 1370
rect 2044 1368 2143 1402
rect -45 1291 -11 1307
rect -45 1222 -11 1257
rect -45 1153 -11 1188
rect 143 1145 2143 1368
rect 2297 1291 2331 1307
rect 2297 1222 2331 1257
rect 2297 1153 2331 1188
rect -45 1111 -11 1119
rect 2297 1111 2331 1119
rect -45 1084 2331 1111
rect -11 1050 2297 1084
rect -45 1015 2331 1050
rect -11 981 2297 1015
rect -45 946 2331 981
rect -11 912 2297 946
rect -45 877 2331 912
rect -11 843 2297 877
rect -45 827 2331 843
rect -45 769 2399 793
rect -45 735 2229 769
rect 2263 735 2297 769
rect 2331 735 2365 769
rect -45 699 2399 735
rect -45 665 2229 699
rect 2263 665 2297 699
rect 2331 665 2365 699
rect -45 629 2399 665
rect -45 595 2229 629
rect 2263 595 2297 629
rect 2331 595 2365 629
rect -45 586 2399 595
rect 2229 559 2399 586
rect 143 329 2143 552
rect 143 223 242 329
rect 276 327 315 329
rect 349 327 388 329
rect 422 327 461 329
rect 495 327 534 329
rect 568 327 607 329
rect 641 327 680 329
rect 714 327 753 329
rect 787 327 826 329
rect 860 327 900 329
rect 934 327 974 329
rect 1008 327 1048 329
rect 1082 327 1122 329
rect 1156 327 1196 329
rect 1230 327 1270 329
rect 1304 327 1344 329
rect 1378 327 1418 329
rect 1452 327 1492 329
rect 1526 327 1566 329
rect 1600 327 1640 329
rect 1674 327 1714 329
rect 1748 327 1788 329
rect 1822 327 1862 329
rect 1896 327 1936 329
rect 1970 327 2010 329
rect 1976 295 2010 327
rect 2044 295 2143 329
rect 1976 257 2143 295
rect 1976 225 2010 257
rect 276 223 315 225
rect 349 223 388 225
rect 422 223 461 225
rect 495 223 534 225
rect 568 223 607 225
rect 641 223 680 225
rect 714 223 753 225
rect 787 223 826 225
rect 860 223 900 225
rect 934 223 974 225
rect 1008 223 1048 225
rect 1082 223 1122 225
rect 1156 223 1196 225
rect 1230 223 1270 225
rect 1304 223 1344 225
rect 1378 223 1418 225
rect 1452 223 1492 225
rect 1526 223 1566 225
rect 1600 223 1640 225
rect 1674 223 1714 225
rect 1748 223 1788 225
rect 1822 223 1862 225
rect 1896 223 1936 225
rect 1970 223 2010 225
rect 2044 223 2143 257
rect 143 85 2143 223
rect 2263 525 2297 559
rect 2331 525 2365 559
rect 2229 489 2399 525
rect 2263 455 2297 489
rect 2331 455 2365 489
rect 2229 419 2399 455
rect 2263 385 2297 419
rect 2331 385 2365 419
rect 2229 349 2399 385
rect 2263 315 2297 349
rect 2331 315 2365 349
rect 2229 279 2399 315
rect 2263 245 2297 279
rect 2331 245 2365 279
rect 2229 209 2399 245
rect 2263 175 2297 209
rect 2331 175 2365 209
rect 2229 138 2399 175
rect 2263 104 2297 138
rect 2331 104 2365 138
rect 2229 67 2399 104
rect 2263 33 2297 67
rect 2331 33 2365 67
rect 2229 -1 2399 33
<< viali >>
rect 242 3762 276 3764
rect 315 3762 349 3764
rect 388 3762 422 3764
rect 461 3762 495 3764
rect 534 3762 568 3764
rect 607 3762 641 3764
rect 680 3762 714 3764
rect 753 3762 787 3764
rect 826 3762 860 3764
rect 900 3762 934 3764
rect 974 3762 1008 3764
rect 1048 3762 1082 3764
rect 1122 3762 1156 3764
rect 1196 3762 1230 3764
rect 1270 3762 1304 3764
rect 1344 3762 1378 3764
rect 1418 3762 1452 3764
rect 1492 3762 1526 3764
rect 1566 3762 1600 3764
rect 1640 3762 1674 3764
rect 1714 3762 1748 3764
rect 1788 3762 1822 3764
rect 1862 3762 1896 3764
rect 1936 3762 1970 3764
rect 242 3730 276 3762
rect 315 3730 349 3762
rect 388 3730 422 3762
rect 461 3730 495 3762
rect 534 3730 568 3762
rect 607 3730 641 3762
rect 680 3730 714 3762
rect 753 3730 787 3762
rect 826 3730 860 3762
rect 900 3730 934 3762
rect 974 3730 1008 3762
rect 1048 3730 1082 3762
rect 1122 3730 1156 3762
rect 1196 3730 1230 3762
rect 1270 3730 1304 3762
rect 1344 3730 1378 3762
rect 1418 3730 1452 3762
rect 1492 3730 1526 3762
rect 1566 3730 1600 3762
rect 1640 3730 1674 3762
rect 1714 3730 1748 3762
rect 1788 3730 1822 3762
rect 1862 3730 1896 3762
rect 1936 3730 1970 3762
rect 2010 3730 2044 3764
rect 242 3660 276 3692
rect 315 3660 349 3692
rect 388 3660 422 3692
rect 461 3660 495 3692
rect 534 3660 568 3692
rect 607 3660 641 3692
rect 680 3660 714 3692
rect 753 3660 787 3692
rect 826 3660 860 3692
rect 900 3660 934 3692
rect 974 3660 1008 3692
rect 1048 3660 1082 3692
rect 1122 3660 1156 3692
rect 1196 3660 1230 3692
rect 1270 3660 1304 3692
rect 1344 3660 1378 3692
rect 1418 3660 1452 3692
rect 1492 3660 1526 3692
rect 1566 3660 1600 3692
rect 1640 3660 1674 3692
rect 1714 3660 1748 3692
rect 1788 3660 1822 3692
rect 1862 3660 1896 3692
rect 1936 3660 1970 3692
rect 242 3658 276 3660
rect 315 3658 349 3660
rect 388 3658 422 3660
rect 461 3658 495 3660
rect 534 3658 568 3660
rect 607 3658 641 3660
rect 680 3658 714 3660
rect 753 3658 787 3660
rect 826 3658 860 3660
rect 900 3658 934 3660
rect 974 3658 1008 3660
rect 1048 3658 1082 3660
rect 1122 3658 1156 3660
rect 1196 3658 1230 3660
rect 1270 3658 1304 3660
rect 1344 3658 1378 3660
rect 1418 3658 1452 3660
rect 1492 3658 1526 3660
rect 1566 3658 1600 3660
rect 1640 3658 1674 3660
rect 1714 3658 1748 3660
rect 1788 3658 1822 3660
rect 1862 3658 1896 3660
rect 1936 3658 1970 3660
rect 2010 3658 2044 3692
rect 242 2617 276 2619
rect 315 2617 349 2619
rect 388 2617 422 2619
rect 461 2617 495 2619
rect 534 2617 568 2619
rect 607 2617 641 2619
rect 680 2617 714 2619
rect 753 2617 787 2619
rect 826 2617 860 2619
rect 900 2617 934 2619
rect 974 2617 1008 2619
rect 1048 2617 1082 2619
rect 1122 2617 1156 2619
rect 1196 2617 1230 2619
rect 1270 2617 1304 2619
rect 1344 2617 1378 2619
rect 1418 2617 1452 2619
rect 1492 2617 1526 2619
rect 1566 2617 1600 2619
rect 1640 2617 1674 2619
rect 1714 2617 1748 2619
rect 1788 2617 1822 2619
rect 1862 2617 1896 2619
rect 1936 2617 1970 2619
rect 242 2585 276 2617
rect 315 2585 349 2617
rect 388 2585 422 2617
rect 461 2585 495 2617
rect 534 2585 568 2617
rect 607 2585 641 2617
rect 680 2585 714 2617
rect 753 2585 787 2617
rect 826 2585 860 2617
rect 900 2585 934 2617
rect 974 2585 1008 2617
rect 1048 2585 1082 2617
rect 1122 2585 1156 2617
rect 1196 2585 1230 2617
rect 1270 2585 1304 2617
rect 1344 2585 1378 2617
rect 1418 2585 1452 2617
rect 1492 2585 1526 2617
rect 1566 2585 1600 2617
rect 1640 2585 1674 2617
rect 1714 2585 1748 2617
rect 1788 2585 1822 2617
rect 1862 2585 1896 2617
rect 1936 2585 1970 2617
rect 2010 2585 2044 2619
rect 242 2515 276 2547
rect 315 2515 349 2547
rect 388 2515 422 2547
rect 461 2515 495 2547
rect 534 2515 568 2547
rect 607 2515 641 2547
rect 680 2515 714 2547
rect 753 2515 787 2547
rect 826 2515 860 2547
rect 900 2515 934 2547
rect 974 2515 1008 2547
rect 1048 2515 1082 2547
rect 1122 2515 1156 2547
rect 1196 2515 1230 2547
rect 1270 2515 1304 2547
rect 1344 2515 1378 2547
rect 1418 2515 1452 2547
rect 1492 2515 1526 2547
rect 1566 2515 1600 2547
rect 1640 2515 1674 2547
rect 1714 2515 1748 2547
rect 1788 2515 1822 2547
rect 1862 2515 1896 2547
rect 1936 2515 1970 2547
rect 242 2513 276 2515
rect 315 2513 349 2515
rect 388 2513 422 2515
rect 461 2513 495 2515
rect 534 2513 568 2515
rect 607 2513 641 2515
rect 680 2513 714 2515
rect 753 2513 787 2515
rect 826 2513 860 2515
rect 900 2513 934 2515
rect 974 2513 1008 2515
rect 1048 2513 1082 2515
rect 1122 2513 1156 2515
rect 1196 2513 1230 2515
rect 1270 2513 1304 2515
rect 1344 2513 1378 2515
rect 1418 2513 1452 2515
rect 1492 2513 1526 2515
rect 1566 2513 1600 2515
rect 1640 2513 1674 2515
rect 1714 2513 1748 2515
rect 1788 2513 1822 2515
rect 1862 2513 1896 2515
rect 1936 2513 1970 2515
rect 2010 2513 2044 2547
rect 242 1472 276 1474
rect 315 1472 349 1474
rect 388 1472 422 1474
rect 461 1472 495 1474
rect 534 1472 568 1474
rect 607 1472 641 1474
rect 680 1472 714 1474
rect 753 1472 787 1474
rect 826 1472 860 1474
rect 900 1472 934 1474
rect 974 1472 1008 1474
rect 1048 1472 1082 1474
rect 1122 1472 1156 1474
rect 1196 1472 1230 1474
rect 1270 1472 1304 1474
rect 1344 1472 1378 1474
rect 1418 1472 1452 1474
rect 1492 1472 1526 1474
rect 1566 1472 1600 1474
rect 1640 1472 1674 1474
rect 1714 1472 1748 1474
rect 1788 1472 1822 1474
rect 1862 1472 1896 1474
rect 1936 1472 1970 1474
rect 242 1440 276 1472
rect 315 1440 349 1472
rect 388 1440 422 1472
rect 461 1440 495 1472
rect 534 1440 568 1472
rect 607 1440 641 1472
rect 680 1440 714 1472
rect 753 1440 787 1472
rect 826 1440 860 1472
rect 900 1440 934 1472
rect 974 1440 1008 1472
rect 1048 1440 1082 1472
rect 1122 1440 1156 1472
rect 1196 1440 1230 1472
rect 1270 1440 1304 1472
rect 1344 1440 1378 1472
rect 1418 1440 1452 1472
rect 1492 1440 1526 1472
rect 1566 1440 1600 1472
rect 1640 1440 1674 1472
rect 1714 1440 1748 1472
rect 1788 1440 1822 1472
rect 1862 1440 1896 1472
rect 1936 1440 1970 1472
rect 2010 1440 2044 1474
rect 242 1370 276 1402
rect 315 1370 349 1402
rect 388 1370 422 1402
rect 461 1370 495 1402
rect 534 1370 568 1402
rect 607 1370 641 1402
rect 680 1370 714 1402
rect 753 1370 787 1402
rect 826 1370 860 1402
rect 900 1370 934 1402
rect 974 1370 1008 1402
rect 1048 1370 1082 1402
rect 1122 1370 1156 1402
rect 1196 1370 1230 1402
rect 1270 1370 1304 1402
rect 1344 1370 1378 1402
rect 1418 1370 1452 1402
rect 1492 1370 1526 1402
rect 1566 1370 1600 1402
rect 1640 1370 1674 1402
rect 1714 1370 1748 1402
rect 1788 1370 1822 1402
rect 1862 1370 1896 1402
rect 1936 1370 1970 1402
rect 242 1368 276 1370
rect 315 1368 349 1370
rect 388 1368 422 1370
rect 461 1368 495 1370
rect 534 1368 568 1370
rect 607 1368 641 1370
rect 680 1368 714 1370
rect 753 1368 787 1370
rect 826 1368 860 1370
rect 900 1368 934 1370
rect 974 1368 1008 1370
rect 1048 1368 1082 1370
rect 1122 1368 1156 1370
rect 1196 1368 1230 1370
rect 1270 1368 1304 1370
rect 1344 1368 1378 1370
rect 1418 1368 1452 1370
rect 1492 1368 1526 1370
rect 1566 1368 1600 1370
rect 1640 1368 1674 1370
rect 1714 1368 1748 1370
rect 1788 1368 1822 1370
rect 1862 1368 1896 1370
rect 1936 1368 1970 1370
rect 2010 1368 2044 1402
rect 242 327 276 329
rect 315 327 349 329
rect 388 327 422 329
rect 461 327 495 329
rect 534 327 568 329
rect 607 327 641 329
rect 680 327 714 329
rect 753 327 787 329
rect 826 327 860 329
rect 900 327 934 329
rect 974 327 1008 329
rect 1048 327 1082 329
rect 1122 327 1156 329
rect 1196 327 1230 329
rect 1270 327 1304 329
rect 1344 327 1378 329
rect 1418 327 1452 329
rect 1492 327 1526 329
rect 1566 327 1600 329
rect 1640 327 1674 329
rect 1714 327 1748 329
rect 1788 327 1822 329
rect 1862 327 1896 329
rect 1936 327 1970 329
rect 242 295 276 327
rect 315 295 349 327
rect 388 295 422 327
rect 461 295 495 327
rect 534 295 568 327
rect 607 295 641 327
rect 680 295 714 327
rect 753 295 787 327
rect 826 295 860 327
rect 900 295 934 327
rect 974 295 1008 327
rect 1048 295 1082 327
rect 1122 295 1156 327
rect 1196 295 1230 327
rect 1270 295 1304 327
rect 1344 295 1378 327
rect 1418 295 1452 327
rect 1492 295 1526 327
rect 1566 295 1600 327
rect 1640 295 1674 327
rect 1714 295 1748 327
rect 1788 295 1822 327
rect 1862 295 1896 327
rect 1936 295 1970 327
rect 2010 295 2044 329
rect 242 225 276 257
rect 315 225 349 257
rect 388 225 422 257
rect 461 225 495 257
rect 534 225 568 257
rect 607 225 641 257
rect 680 225 714 257
rect 753 225 787 257
rect 826 225 860 257
rect 900 225 934 257
rect 974 225 1008 257
rect 1048 225 1082 257
rect 1122 225 1156 257
rect 1196 225 1230 257
rect 1270 225 1304 257
rect 1344 225 1378 257
rect 1418 225 1452 257
rect 1492 225 1526 257
rect 1566 225 1600 257
rect 1640 225 1674 257
rect 1714 225 1748 257
rect 1788 225 1822 257
rect 1862 225 1896 257
rect 1936 225 1970 257
rect 242 223 276 225
rect 315 223 349 225
rect 388 223 422 225
rect 461 223 495 225
rect 534 223 568 225
rect 607 223 641 225
rect 680 223 714 225
rect 753 223 787 225
rect 826 223 860 225
rect 900 223 934 225
rect 974 223 1008 225
rect 1048 223 1082 225
rect 1122 223 1156 225
rect 1196 223 1230 225
rect 1270 223 1304 225
rect 1344 223 1378 225
rect 1418 223 1452 225
rect 1492 223 1526 225
rect 1566 223 1600 225
rect 1640 223 1674 225
rect 1714 223 1748 225
rect 1788 223 1822 225
rect 1862 223 1896 225
rect 1936 223 1970 225
rect 2010 223 2044 257
<< metal1 >>
tri 230 3940 277 3987 se
rect 277 3940 2009 3987
tri 2009 3940 2056 3987 sw
rect 230 3764 2056 3940
rect 230 3730 242 3764
rect 276 3730 315 3764
rect 349 3730 388 3764
rect 422 3730 461 3764
rect 495 3730 534 3764
rect 568 3730 607 3764
rect 641 3730 680 3764
rect 714 3730 753 3764
rect 787 3730 826 3764
rect 860 3730 900 3764
rect 934 3730 974 3764
rect 1008 3730 1048 3764
rect 1082 3730 1122 3764
rect 1156 3730 1196 3764
rect 1230 3730 1270 3764
rect 1304 3730 1344 3764
rect 1378 3730 1418 3764
rect 1452 3730 1492 3764
rect 1526 3730 1566 3764
rect 1600 3730 1640 3764
rect 1674 3730 1714 3764
rect 1748 3730 1788 3764
rect 1822 3730 1862 3764
rect 1896 3730 1936 3764
rect 1970 3730 2010 3764
rect 2044 3730 2056 3764
rect 230 3692 2056 3730
rect 230 3658 242 3692
rect 276 3658 315 3692
rect 349 3658 388 3692
rect 422 3658 461 3692
rect 495 3658 534 3692
rect 568 3658 607 3692
rect 641 3658 680 3692
rect 714 3658 753 3692
rect 787 3658 826 3692
rect 860 3658 900 3692
rect 934 3658 974 3692
rect 1008 3658 1048 3692
rect 1082 3658 1122 3692
rect 1156 3658 1196 3692
rect 1230 3658 1270 3692
rect 1304 3658 1344 3692
rect 1378 3658 1418 3692
rect 1452 3658 1492 3692
rect 1526 3658 1566 3692
rect 1600 3658 1640 3692
rect 1674 3658 1714 3692
rect 1748 3658 1788 3692
rect 1822 3658 1862 3692
rect 1896 3658 1936 3692
rect 1970 3658 2010 3692
rect 2044 3658 2056 3692
rect 230 3482 2056 3658
tri 230 3435 277 3482 ne
rect 277 3435 2009 3482
tri 2009 3435 2056 3482 nw
tri 230 2795 277 2842 se
rect 277 2795 2009 2842
tri 2009 2795 2056 2842 sw
rect 230 2619 2056 2795
rect 230 2585 242 2619
rect 276 2585 315 2619
rect 349 2585 388 2619
rect 422 2585 461 2619
rect 495 2585 534 2619
rect 568 2585 607 2619
rect 641 2585 680 2619
rect 714 2585 753 2619
rect 787 2585 826 2619
rect 860 2585 900 2619
rect 934 2585 974 2619
rect 1008 2585 1048 2619
rect 1082 2585 1122 2619
rect 1156 2585 1196 2619
rect 1230 2585 1270 2619
rect 1304 2585 1344 2619
rect 1378 2585 1418 2619
rect 1452 2585 1492 2619
rect 1526 2585 1566 2619
rect 1600 2585 1640 2619
rect 1674 2585 1714 2619
rect 1748 2585 1788 2619
rect 1822 2585 1862 2619
rect 1896 2585 1936 2619
rect 1970 2585 2010 2619
rect 2044 2585 2056 2619
rect 230 2547 2056 2585
rect 230 2513 242 2547
rect 276 2513 315 2547
rect 349 2513 388 2547
rect 422 2513 461 2547
rect 495 2513 534 2547
rect 568 2513 607 2547
rect 641 2513 680 2547
rect 714 2513 753 2547
rect 787 2513 826 2547
rect 860 2513 900 2547
rect 934 2513 974 2547
rect 1008 2513 1048 2547
rect 1082 2513 1122 2547
rect 1156 2513 1196 2547
rect 1230 2513 1270 2547
rect 1304 2513 1344 2547
rect 1378 2513 1418 2547
rect 1452 2513 1492 2547
rect 1526 2513 1566 2547
rect 1600 2513 1640 2547
rect 1674 2513 1714 2547
rect 1748 2513 1788 2547
rect 1822 2513 1862 2547
rect 1896 2513 1936 2547
rect 1970 2513 2010 2547
rect 2044 2513 2056 2547
rect 230 2290 2056 2513
rect 231 2288 2055 2289
rect 230 2232 2056 2288
rect 231 2231 2055 2232
rect 230 2178 2056 2230
tri 230 1576 351 1697 se
rect 351 1576 1935 1697
tri 1935 1576 2056 1697 sw
rect 230 1474 2056 1576
rect 230 1440 242 1474
rect 276 1440 315 1474
rect 349 1440 388 1474
rect 422 1440 461 1474
rect 495 1440 534 1474
rect 568 1440 607 1474
rect 641 1440 680 1474
rect 714 1440 753 1474
rect 787 1440 826 1474
rect 860 1440 900 1474
rect 934 1440 974 1474
rect 1008 1440 1048 1474
rect 1082 1440 1122 1474
rect 1156 1440 1196 1474
rect 1230 1440 1270 1474
rect 1304 1440 1344 1474
rect 1378 1440 1418 1474
rect 1452 1440 1492 1474
rect 1526 1440 1566 1474
rect 1600 1440 1640 1474
rect 1674 1440 1714 1474
rect 1748 1440 1788 1474
rect 1822 1440 1862 1474
rect 1896 1440 1936 1474
rect 1970 1440 2010 1474
rect 2044 1440 2056 1474
rect 230 1402 2056 1440
rect 230 1368 242 1402
rect 276 1368 315 1402
rect 349 1368 388 1402
rect 422 1368 461 1402
rect 495 1368 534 1402
rect 568 1368 607 1402
rect 641 1368 680 1402
rect 714 1368 753 1402
rect 787 1368 826 1402
rect 860 1368 900 1402
rect 934 1368 974 1402
rect 1008 1368 1048 1402
rect 1082 1368 1122 1402
rect 1156 1368 1196 1402
rect 1230 1368 1270 1402
rect 1304 1368 1344 1402
rect 1378 1368 1418 1402
rect 1452 1368 1492 1402
rect 1526 1368 1566 1402
rect 1600 1368 1640 1402
rect 1674 1368 1714 1402
rect 1748 1368 1788 1402
rect 1822 1368 1862 1402
rect 1896 1368 1936 1402
rect 1970 1368 2010 1402
rect 2044 1368 2056 1402
rect 230 1258 2056 1368
tri 230 1145 343 1258 ne
rect 343 1145 1943 1258
tri 1943 1145 2056 1258 nw
rect 214 522 2072 574
rect 215 520 2071 521
rect 214 464 2072 520
rect 215 463 2071 464
rect 214 329 2072 462
rect 214 295 242 329
rect 276 295 315 329
rect 349 295 388 329
rect 422 295 461 329
rect 495 295 534 329
rect 568 295 607 329
rect 641 295 680 329
rect 714 295 753 329
rect 787 295 826 329
rect 860 295 900 329
rect 934 295 974 329
rect 1008 295 1048 329
rect 1082 295 1122 329
rect 1156 295 1196 329
rect 1230 295 1270 329
rect 1304 295 1344 329
rect 1378 295 1418 329
rect 1452 295 1492 329
rect 1526 295 1566 329
rect 1600 295 1640 329
rect 1674 295 1714 329
rect 1748 295 1788 329
rect 1822 295 1862 329
rect 1896 295 1936 329
rect 1970 295 2010 329
rect 2044 295 2072 329
rect 214 257 2072 295
rect 214 223 242 257
rect 276 223 315 257
rect 349 223 388 257
rect 422 223 461 257
rect 495 223 534 257
rect 568 223 607 257
rect 641 223 680 257
rect 714 223 753 257
rect 787 223 826 257
rect 860 223 900 257
rect 934 223 974 257
rect 1008 223 1048 257
rect 1082 223 1122 257
rect 1156 223 1196 257
rect 1230 223 1270 257
rect 1304 223 1344 257
rect 1378 223 1418 257
rect 1452 223 1492 257
rect 1526 223 1566 257
rect 1600 223 1640 257
rect 1674 223 1714 257
rect 1748 223 1788 257
rect 1822 223 1862 257
rect 1896 223 1936 257
rect 1970 223 2010 257
rect 2044 223 2072 257
rect 214 90 2072 223
tri 214 43 261 90 ne
rect 261 43 2025 90
tri 2025 43 2072 90 nw
<< rmetal1 >>
rect 230 2289 2056 2290
rect 230 2288 231 2289
rect 2055 2288 2056 2289
rect 230 2231 231 2232
rect 2055 2231 2056 2232
rect 230 2230 2056 2231
rect 214 521 2072 522
rect 214 520 215 521
rect 2071 520 2072 521
rect 214 463 215 464
rect 2071 463 2072 464
rect 214 462 2072 463
use sky130_fd_io__tk_em1s_CDNS_524688791851594  sky130_fd_io__tk_em1s_CDNS_524688791851594_0
timestamp 1701704242
transform 0 1 230 -1 0 2342
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851596  sky130_fd_io__tk_em1s_CDNS_524688791851596_0
timestamp 1701704242
transform 0 1 214 1 0 410
box 0 0 1 1
<< properties >>
string GDS_END 94823922
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94763772
string path 50.350 92.775 5.100 92.775 
<< end >>
