magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 176 326
<< mvnmos >>
rect 0 0 100 300
<< mvndiff >>
rect -53 250 0 300
rect -53 216 -45 250
rect -11 216 0 250
rect -53 182 0 216
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 100 0 150 300
<< mvndiffc >>
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
<< poly >>
rect 0 300 100 326
rect 0 -26 100 0
<< locali >>
rect -45 250 -11 266
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
use hvDFL1sd_CDNS_52468879185376  hvDFL1sd_CDNS_52468879185376_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
flabel comment s 125 150 125 150 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87730216
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87729442
<< end >>
