magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 322 1066
<< mvpmos >>
rect 0 0 200 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 200 0 250 1000
<< poly >>
rect 0 1000 200 1032
rect 0 -32 200 0
<< locali >>
rect 211 -4 245 946
<< metal1 >>
rect -51 -16 -5 978
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_0
timestamp 1701704242
transform 1 0 200 0 1 0
box -36 -36 92 1036
use hvDFM1sd_CDNS_52468879185165  hvDFM1sd_CDNS_52468879185165_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 481 -28 481 0 FreeSans 300 0 0 0 D
flabel comment s 228 471 228 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85612062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85611044
<< end >>
