magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pdiff >>
rect 14875 1324 14913 1656
rect 14875 1288 15671 1324
<< locali >>
rect 16205 1882 16239 1920
<< viali >>
rect 16205 1920 16239 1954
rect 16205 1848 16239 1882
<< metal1 >>
rect 35159 13541 35479 13587
rect 21351 13052 21671 13098
rect 22660 11377 22980 11425
rect 22572 10959 22892 11007
tri 6158 9331 6198 9371 sw
tri 6158 9290 6159 9291 nw
rect 30784 9103 31104 9149
tri 4001 9007 4055 9061 ne
tri 8144 7574 8183 7613 se
tri 7181 7003 7187 7009 se
tri 7239 7003 7245 7009 sw
tri 12514 6678 12528 6692 sw
rect 12514 6669 12528 6678
tri 12528 6669 12537 6678 sw
rect 16834 6672 18250 6678
rect 16886 6626 18250 6672
rect 16886 6624 16928 6626
tri 16928 6624 16930 6626 nw
rect 16886 6620 16894 6624
tri 12514 6594 12537 6617 nw
rect 14030 6590 14038 6618
tri 14038 6590 14066 6618 nw
rect 16834 6608 16894 6620
tri 14030 6582 14038 6590 nw
rect 16886 6590 16894 6608
tri 16894 6590 16928 6624 nw
tri 18723 6590 18757 6624 se
tri 16886 6582 16894 6590 nw
rect 16834 6550 16886 6556
tri 18715 6506 18757 6548 ne
tri 8386 6452 8387 6453 nw
tri 14043 6423 14069 6449 se
tri 14043 6345 14069 6371 ne
rect 18331 5841 18365 5878
rect 27868 5722 28188 5770
rect 36544 5195 36596 5246
tri 5959 5137 5960 5138 ne
tri 6076 5137 6077 5138 nw
rect 15634 2160 15640 2212
rect 15692 2160 15704 2212
rect 15756 2206 15762 2212
tri 15762 2206 15768 2212 sw
rect 15756 2160 15778 2206
rect 16199 1954 16245 1966
rect 16199 1920 16205 1954
rect 16239 1920 16245 1954
rect 16199 1882 16245 1920
rect 16199 1848 16205 1882
rect 16239 1848 16245 1882
rect 16199 1836 16245 1848
rect 11610 1562 11616 1614
rect 11668 1562 11680 1614
rect 11732 1562 12012 1614
rect 12064 1562 12076 1614
rect 12128 1562 12134 1614
rect 11690 -190 11696 -138
rect 11748 -190 11760 -138
rect 11812 -190 16689 -138
rect 16741 -190 16753 -138
rect 16805 -190 16811 -138
rect 11516 -355 11522 -303
rect 11574 -355 11586 -303
rect 11638 -355 15365 -303
rect 15417 -355 15429 -303
rect 15481 -355 15487 -303
<< via1 >>
rect 16834 6620 16886 6672
rect 16834 6556 16886 6608
rect 15640 2160 15692 2212
rect 15704 2160 15756 2212
rect 11616 1562 11668 1614
rect 11680 1562 11732 1614
rect 12012 1562 12064 1614
rect 12076 1562 12128 1614
rect 11696 -190 11748 -138
rect 11760 -190 11812 -138
rect 16689 -190 16741 -138
rect 16753 -190 16805 -138
rect 11522 -355 11574 -303
rect 11586 -355 11638 -303
rect 15365 -355 15417 -303
rect 15429 -355 15481 -303
<< metal2 >>
rect 34708 10540 34907 10583
rect 36187 10540 36537 10583
rect 18990 8764 19310 8810
rect 19466 8764 19786 8810
rect 19814 8765 20221 8810
rect 23221 8122 23577 8158
tri 15494 7998 15522 8026 ne
tri 15574 8001 15599 8026 nw
rect 6738 7441 6790 7478
tri 15863 6947 15904 6988 se
tri 16136 6803 16140 6807 sw
rect 16834 6672 16886 6678
rect 18505 6644 18707 6670
rect 16834 6608 16886 6620
rect 16834 6550 16886 6556
tri 16834 6538 16846 6550 ne
rect 12166 5109 12218 5455
rect 5550 5068 5602 5109
rect 10466 5060 10518 5109
rect 10546 5060 10598 5109
rect 11766 5062 11818 5109
rect 12501 5062 12553 5109
rect 12581 5062 12645 5109
rect 13703 5062 13755 5109
rect 13958 5062 13994 5109
rect 14166 5056 14474 5109
rect 14750 5062 14802 5109
rect 14910 5056 15226 5108
rect 16762 5058 16814 5109
rect 3890 4894 4006 4949
rect 5054 4895 6603 4925
rect 5054 4839 5063 4895
rect 5119 4839 5145 4895
rect 5201 4839 5227 4895
rect 5283 4839 5309 4895
rect 5365 4839 5391 4895
rect 5447 4839 5473 4895
rect 5529 4839 5555 4895
rect 5611 4839 5637 4895
rect 5693 4839 5719 4895
rect 5775 4839 5801 4895
rect 5857 4839 5883 4895
rect 5939 4839 5965 4895
rect 6021 4839 6047 4895
rect 6103 4839 6129 4895
rect 6185 4839 6211 4895
rect 6267 4839 6293 4895
rect 6349 4839 6375 4895
rect 6431 4839 6457 4895
rect 6513 4839 6538 4895
rect 6594 4839 6603 4895
rect 5054 4809 6603 4839
rect 15030 4454 15081 4491
rect 12678 4223 12910 4232
rect 12678 4167 12686 4223
rect 12742 4167 12766 4223
rect 12822 4167 12846 4223
rect 12902 4167 12910 4223
rect 12678 4122 12910 4167
rect 12678 4066 12686 4122
rect 12742 4066 12766 4122
rect 12822 4066 12846 4122
rect 12902 4066 12910 4122
rect 12678 4021 12910 4066
rect 12678 3965 12686 4021
rect 12742 3965 12766 4021
rect 12822 3965 12846 4021
rect 12902 3965 12910 4021
rect 12678 3956 12910 3965
rect 4526 3894 6313 3910
rect 4526 3838 4535 3894
rect 4591 3838 4617 3894
rect 4673 3838 4699 3894
rect 4755 3838 4781 3894
rect 4837 3838 4863 3894
rect 4919 3838 4945 3894
rect 5001 3838 5027 3894
rect 5083 3838 5109 3894
rect 5165 3838 5191 3894
rect 5247 3838 5273 3894
rect 5329 3838 5355 3894
rect 5411 3838 5437 3894
rect 5493 3838 5519 3894
rect 5575 3838 5600 3894
rect 5656 3838 5681 3894
rect 5737 3838 5762 3894
rect 5818 3838 5843 3894
rect 5899 3838 5924 3894
rect 5980 3838 6005 3894
rect 6061 3838 6086 3894
rect 6142 3838 6167 3894
rect 6223 3838 6248 3894
rect 6304 3838 6313 3894
rect 4526 3814 6313 3838
rect 4526 3758 4535 3814
rect 4591 3758 4617 3814
rect 4673 3758 4699 3814
rect 4755 3758 4781 3814
rect 4837 3758 4863 3814
rect 4919 3758 4945 3814
rect 5001 3758 5027 3814
rect 5083 3758 5109 3814
rect 5165 3758 5191 3814
rect 5247 3758 5273 3814
rect 5329 3758 5355 3814
rect 5411 3758 5437 3814
rect 5493 3758 5519 3814
rect 5575 3758 5600 3814
rect 5656 3758 5681 3814
rect 5737 3758 5762 3814
rect 5818 3758 5843 3814
rect 5899 3758 5924 3814
rect 5980 3758 6005 3814
rect 6061 3758 6086 3814
rect 6142 3758 6167 3814
rect 6223 3758 6248 3814
rect 6304 3758 6313 3814
rect 4526 3742 6313 3758
tri 12012 2947 12086 3021 se
rect 12086 2999 12138 3913
tri 16788 3177 16846 3235 se
rect 16846 3217 16886 6550
rect 20364 6356 20864 6404
rect 21167 6356 21486 6404
rect 33067 6356 33387 6450
rect 22069 5546 22389 5594
rect 22417 5546 22737 5594
rect 23793 5532 24113 5594
rect 24461 5500 24760 5595
rect 25461 5500 26071 5594
rect 26179 5500 26751 5594
rect 27006 5500 27374 5594
rect 27430 5500 28113 5594
rect 28224 5500 29181 5594
rect 29409 5500 30066 5594
rect 30530 5500 30922 5594
rect 31163 5500 31359 5594
rect 31520 5500 31840 5594
rect 33707 5500 33885 5594
rect 33916 5500 34044 5594
rect 34088 5500 34401 5594
rect 33010 5248 33297 5342
rect 33477 5134 33605 5135
rect 17299 5059 17425 5106
rect 17476 5058 17528 5109
rect 17734 5056 18019 5108
rect 35437 5036 35757 5130
tri 16846 3177 16886 3217 nw
tri 16730 3119 16788 3177 se
tri 16788 3119 16846 3177 nw
tri 16672 3061 16730 3119 se
tri 16730 3061 16788 3119 nw
tri 16614 3003 16672 3061 se
tri 16672 3003 16730 3061 nw
tri 12086 2947 12138 2999 nw
tri 16589 2978 16614 3003 se
rect 16614 2978 16647 3003
tri 16647 2978 16672 3003 nw
tri 12006 2941 12012 2947 se
rect 12012 2941 12080 2947
tri 12080 2941 12086 2947 nw
rect 12006 1614 12058 2941
tri 12058 2919 12080 2941 nw
rect 16589 2496 16629 2978
tri 16629 2960 16647 2978 nw
tri 16629 2496 16647 2514 sw
tri 16589 2438 16647 2496 ne
tri 16647 2474 16669 2496 sw
rect 16647 2438 16669 2474
tri 16669 2438 16705 2474 sw
tri 16647 2416 16669 2438 ne
rect 16669 2434 16705 2438
tri 16705 2434 16709 2438 sw
rect 15634 2160 15640 2212
rect 15692 2160 15704 2212
rect 15756 2160 15762 2212
tri 15560 2005 15634 2079 se
rect 15634 2057 15686 2160
tri 15686 2115 15731 2160 nw
tri 15634 2005 15686 2057 nw
tri 15486 1931 15560 2005 se
tri 15560 1931 15634 2005 nw
tri 15412 1857 15486 1931 se
tri 15486 1857 15560 1931 nw
tri 15397 1842 15412 1857 se
rect 15412 1842 15471 1857
tri 15471 1842 15486 1857 nw
tri 12058 1614 12134 1690 sw
rect 11610 1562 11616 1614
rect 11668 1562 11680 1614
rect 11732 1562 11738 1614
rect 12006 1562 12012 1614
rect 12064 1562 12076 1614
rect 12128 1562 12134 1614
tri 11610 1524 11648 1562 ne
tri 11574 956 11648 1030 se
rect 11648 1008 11700 1562
tri 11700 1524 11738 1562 nw
tri 11648 956 11700 1008 nw
tri 11516 898 11574 956 se
rect 11574 898 11590 956
tri 11590 898 11648 956 nw
rect 10480 -50 10532 -5
rect 10560 -50 10612 -5
rect 11516 -265 11568 898
tri 11568 876 11590 898 nw
tri 11690 716 11766 792 ne
tri 11729 -138 11766 -101 se
rect 11766 -138 11818 792
rect 11690 -190 11696 -138
rect 11748 -190 11760 -138
rect 11812 -190 11818 -138
tri 11568 -265 11606 -227 sw
rect 11516 -303 11606 -265
tri 11606 -303 11644 -265 sw
rect 11516 -355 11522 -303
rect 11574 -355 11586 -303
rect 11638 -355 11644 -303
tri 15359 -303 15397 -265 se
rect 15397 -303 15449 1842
tri 15449 1820 15471 1842 nw
rect 16669 1834 16709 2434
tri 16709 1834 16727 1852 sw
tri 16669 1820 16683 1834 ne
rect 16683 1820 16727 1834
tri 16683 1776 16727 1820 ne
tri 16727 1790 16771 1834 sw
rect 16727 1776 16771 1790
tri 16771 1776 16785 1790 sw
tri 16727 1732 16771 1776 ne
rect 16771 1750 16785 1776
tri 16785 1750 16811 1776 sw
rect 16446 417 16599 495
tri 16728 -138 16771 -95 se
rect 16771 -138 16811 1750
rect 16683 -190 16689 -138
rect 16741 -190 16753 -138
rect 16805 -190 16811 -138
tri 15449 -303 15487 -265 sw
rect 15359 -355 15365 -303
rect 15417 -355 15429 -303
rect 15481 -355 15487 -303
<< via2 >>
rect 5063 4839 5119 4895
rect 5145 4839 5201 4895
rect 5227 4839 5283 4895
rect 5309 4839 5365 4895
rect 5391 4839 5447 4895
rect 5473 4839 5529 4895
rect 5555 4839 5611 4895
rect 5637 4839 5693 4895
rect 5719 4839 5775 4895
rect 5801 4839 5857 4895
rect 5883 4839 5939 4895
rect 5965 4839 6021 4895
rect 6047 4839 6103 4895
rect 6129 4839 6185 4895
rect 6211 4839 6267 4895
rect 6293 4839 6349 4895
rect 6375 4839 6431 4895
rect 6457 4839 6513 4895
rect 6538 4839 6594 4895
rect 12686 4167 12742 4223
rect 12766 4167 12822 4223
rect 12846 4167 12902 4223
rect 12686 4066 12742 4122
rect 12766 4066 12822 4122
rect 12846 4066 12902 4122
rect 12686 3965 12742 4021
rect 12766 3965 12822 4021
rect 12846 3965 12902 4021
rect 4535 3838 4591 3894
rect 4617 3838 4673 3894
rect 4699 3838 4755 3894
rect 4781 3838 4837 3894
rect 4863 3838 4919 3894
rect 4945 3838 5001 3894
rect 5027 3838 5083 3894
rect 5109 3838 5165 3894
rect 5191 3838 5247 3894
rect 5273 3838 5329 3894
rect 5355 3838 5411 3894
rect 5437 3838 5493 3894
rect 5519 3838 5575 3894
rect 5600 3838 5656 3894
rect 5681 3838 5737 3894
rect 5762 3838 5818 3894
rect 5843 3838 5899 3894
rect 5924 3838 5980 3894
rect 6005 3838 6061 3894
rect 6086 3838 6142 3894
rect 6167 3838 6223 3894
rect 6248 3838 6304 3894
rect 4535 3758 4591 3814
rect 4617 3758 4673 3814
rect 4699 3758 4755 3814
rect 4781 3758 4837 3814
rect 4863 3758 4919 3814
rect 4945 3758 5001 3814
rect 5027 3758 5083 3814
rect 5109 3758 5165 3814
rect 5191 3758 5247 3814
rect 5273 3758 5329 3814
rect 5355 3758 5411 3814
rect 5437 3758 5493 3814
rect 5519 3758 5575 3814
rect 5600 3758 5656 3814
rect 5681 3758 5737 3814
rect 5762 3758 5818 3814
rect 5843 3758 5899 3814
rect 5924 3758 5980 3814
rect 6005 3758 6061 3814
rect 6086 3758 6142 3814
rect 6167 3758 6223 3814
rect 6248 3758 6304 3814
<< metal3 >>
rect 32693 6180 35051 7028
rect 5053 5589 12125 5594
tri 12125 5589 12130 5594 sw
tri 12451 5589 12456 5594 se
rect 12456 5589 18919 5594
rect 5053 5564 12130 5589
tri 12130 5564 12155 5589 sw
tri 12426 5564 12451 5589 se
rect 12451 5564 18919 5589
rect 5053 5446 18919 5564
rect 19958 5446 34397 5594
rect 5053 4895 34397 5446
rect 5053 4839 5063 4895
rect 5119 4839 5145 4895
rect 5201 4839 5227 4895
rect 5283 4839 5309 4895
rect 5365 4839 5391 4895
rect 5447 4839 5473 4895
rect 5529 4839 5555 4895
rect 5611 4839 5637 4895
rect 5693 4839 5719 4895
rect 5775 4839 5801 4895
rect 5857 4839 5883 4895
rect 5939 4839 5965 4895
rect 6021 4839 6047 4895
rect 6103 4839 6129 4895
rect 6185 4839 6211 4895
rect 6267 4839 6293 4895
rect 6349 4839 6375 4895
rect 6431 4839 6457 4895
rect 6513 4839 6538 4895
rect 6594 4839 34397 4895
rect 5053 4736 34397 4839
rect 4497 4223 32669 4236
rect 4497 4167 12686 4223
rect 12742 4167 12766 4223
rect 12822 4167 12846 4223
rect 12902 4167 32669 4223
rect 4497 4122 32669 4167
rect 4497 4066 12686 4122
rect 12742 4066 12766 4122
rect 12822 4066 12846 4122
rect 12902 4066 32669 4122
rect 4497 4021 32669 4066
rect 4497 3965 12686 4021
rect 12742 3965 12766 4021
rect 12822 3965 12846 4021
rect 12902 3965 32669 4021
rect 4497 3894 32669 3965
rect 4497 3838 4535 3894
rect 4591 3838 4617 3894
rect 4673 3838 4699 3894
rect 4755 3838 4781 3894
rect 4837 3838 4863 3894
rect 4919 3838 4945 3894
rect 5001 3838 5027 3894
rect 5083 3838 5109 3894
rect 5165 3838 5191 3894
rect 5247 3838 5273 3894
rect 5329 3838 5355 3894
rect 5411 3838 5437 3894
rect 5493 3838 5519 3894
rect 5575 3838 5600 3894
rect 5656 3838 5681 3894
rect 5737 3838 5762 3894
rect 5818 3838 5843 3894
rect 5899 3838 5924 3894
rect 5980 3838 6005 3894
rect 6061 3838 6086 3894
rect 6142 3838 6167 3894
rect 6223 3838 6248 3894
rect 6304 3838 32669 3894
rect 4497 3814 32669 3838
rect 4497 3758 4535 3814
rect 4591 3758 4617 3814
rect 4673 3758 4699 3814
rect 4755 3758 4781 3814
rect 4837 3758 4863 3814
rect 4919 3758 4945 3814
rect 5001 3758 5027 3814
rect 5083 3758 5109 3814
rect 5165 3758 5191 3814
rect 5247 3758 5273 3814
rect 5329 3758 5355 3814
rect 5411 3758 5437 3814
rect 5493 3758 5519 3814
rect 5575 3758 5600 3814
rect 5656 3758 5681 3814
rect 5737 3758 5762 3814
rect 5818 3758 5843 3814
rect 5899 3758 5924 3814
rect 5980 3758 6005 3814
rect 6061 3758 6086 3814
rect 6142 3758 6167 3814
rect 6223 3758 6248 3814
rect 6304 3758 32669 3814
rect 4497 3332 32669 3758
rect 12557 2020 35539 2878
rect 12346 662 19851 1520
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 16239 1 0 1848
box 0 0 1 1
use sky130_fd_io__sio_ibuf_diff_tsg4  sky130_fd_io__sio_ibuf_diff_tsg4_0
timestamp 1701704242
transform 1 0 23031 0 1 -1151
box -6313 647 13870 14823
use sky130_fd_io__sio_ipath_com  sky130_fd_io__sio_ipath_com_0
timestamp 1701704242
transform 1 0 3870 0 1 -50
box 0 -404 14524 7059
<< labels >>
flabel comment s 13479 1139 13479 1139 0 FreeSans 4000 0 0 0 vpb_ka
flabel comment s 13756 2489 13756 2489 0 FreeSans 4000 0 0 0 vpwr_ka
flabel comment s 9956 3811 9956 3811 0 FreeSans 4000 0 0 0 vgnd
flabel comment s 11102 5300 11102 5300 0 FreeSans 1600 0 0 0 vcc_ioq
flabel metal1 s 35159 13541 35479 13587 0 FreeSans 400 0 0 0 vpwr_ka
port 2 nsew
flabel metal1 s 21351 13052 21671 13098 0 FreeSans 400 0 0 0 vpwr_ka
port 2 nsew
flabel metal1 s 30784 9103 31104 9149 0 FreeSans 400 0 0 0 vpwr_ka
port 2 nsew
flabel metal1 s 27868 5722 28188 5770 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal1 s 22660 11377 22980 11425 0 FreeSans 400 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 22572 10959 22892 11007 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal1 s 17829 1457 17829 1457 0 FreeSans 200 0 0 0 out_h_n_einv
flabel metal1 s 17820 830 17820 830 0 FreeSans 200 0 0 0 out_n_einv
flabel metal1 s 18494 6984 18494 6984 0 FreeSans 200 0 0 0 ie_diff_sel_n
flabel metal1 s 18331 5841 18365 5878 7 FreeSans 200 180 0 0 sio_diff_hyst_en_h
port 5 nsew
flabel metal1 s 36544 5195 36596 5246 0 FreeSans 400 180 0 0 vinref
port 6 nsew
flabel metal2 s 12189 5004 12189 5004 0 FreeSans 200 0 0 0 ie_diff_sel_n
flabel metal2 s 18161 2091 18161 2091 0 FreeSans 200 0 0 0 ie_diff_sel_h
flabel metal2 s 18072 2041 18072 2041 0 FreeSans 200 0 0 0 ie_diff_sel_h_n
flabel metal2 s 36187 10540 36537 10583 0 FreeSans 400 0 0 0 vpwr_ka
port 2 nsew
flabel metal2 s 18990 8764 19310 8810 0 FreeSans 400 0 0 0 vpwr_ka
port 2 nsew
flabel metal2 s 19466 8764 19786 8810 0 FreeSans 400 0 0 0 vpb_ka
port 7 nsew
flabel metal2 s 34708 10540 34907 10583 0 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal2 s 23221 8122 23577 8158 0 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal2 s 17476 5058 17528 5109 7 FreeSans 200 90 0 0 inp_dis_h
port 8 nsew
flabel metal2 s 10546 5060 10598 5109 7 FreeSans 200 90 0 0 ibuf_sel_h_n
port 9 nsew
flabel metal2 s 21167 6356 21486 6404 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 35437 5036 35757 5130 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 10466 5060 10518 5109 7 FreeSans 200 90 0 0 ibuf_sel_h
port 10 nsew
flabel metal2 s 12501 5062 12553 5109 7 FreeSans 200 90 0 0 dm_h_n<2>
port 11 nsew
flabel metal2 s 30530 5500 30922 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 29409 5500 30066 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 28224 5500 29181 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 11766 5062 11818 5109 7 FreeSans 200 90 0 0 dm_h_n<1>
port 12 nsew
flabel metal2 s 5550 5068 5602 5109 7 FreeSans 200 90 0 0 dm_h_n<0>
port 13 nsew
flabel metal2 s 27430 5500 28113 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 27006 5500 27374 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 26179 5500 26751 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 25461 5500 26071 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 23793 5532 24113 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 14750 5062 14802 5109 7 FreeSans 200 90 0 0 dm_h<2>
port 14 nsew
flabel metal2 s 22417 5546 22737 5594 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 22069 5546 22389 5594 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 20364 6356 20864 6404 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 34088 5500 34401 5594 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 24461 5500 24760 5595 0 FreeSans 400 180 0 0 vcc_io
port 4 nsew
flabel metal2 s 33010 5248 33297 5342 0 FreeSans 400 180 0 0 vcc_io
port 4 nsew
flabel metal2 s 33916 5500 34044 5594 0 FreeSans 400 180 0 0 pad
port 16 nsew
flabel metal2 s 13958 5062 13994 5109 7 FreeSans 200 90 0 0 vtrip_sel_h_n
port 17 nsew
flabel metal2 s 13703 5062 13755 5109 7 FreeSans 200 90 0 0 vtrip_sel_h
port 18 nsew
flabel metal2 s 14910 5056 15226 5108 0 FreeSans 200 0 0 0 vpwr_ka
port 2 nsew
flabel metal2 s 12581 5062 12645 5109 7 FreeSans 200 90 0 0 dm_h<0>
port 19 nsew
flabel metal2 s 16446 417 16599 495 0 FreeSans 200 0 0 0 vpb_ka
port 7 nsew
flabel metal2 s 33707 5500 33885 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 31520 5500 31840 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 18505 6644 18707 6670 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal2 s 17734 5056 18019 5108 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal2 s 14166 5056 14474 5109 0 FreeSans 200 0 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 3890 4894 4006 4949 0 FreeSans 200 0 0 0 pad
port 16 nsew
flabel metal2 s 10480 -50 10532 -5 3 FreeSans 200 90 0 0 out_h
port 20 nsew
flabel metal2 s 10560 -50 10612 -5 3 FreeSans 200 90 0 0 out
port 21 nsew
flabel metal2 s 16762 5058 16814 5109 7 FreeSans 200 90 0 0 inp_dis_h_n
port 22 nsew
flabel metal2 s 33067 6356 33387 6450 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 6738 7441 6790 7478 3 FreeSans 200 0 0 0 dm_h<1>
port 23 nsew
flabel metal2 s 19814 8765 20221 8810 0 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal2 s 17299 5059 17425 5106 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal2 s 31163 5500 31359 5594 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
<< properties >>
string GDS_END 87511680
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87493114
string path 319.850 99.000 319.850 105.700 
<< end >>
