magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 0 0 1310 647
<< mvpdiff >>
rect 66 434 187 472
rect 66 400 153 434
rect 66 388 187 400
rect 545 434 666 472
rect 579 400 666 434
rect 545 388 666 400
rect 66 112 187 150
rect 66 78 153 112
rect 66 66 187 78
rect 545 112 666 150
rect 579 78 666 112
rect 545 66 666 78
<< mvpdiffc >>
rect 153 400 187 434
rect 545 400 579 434
rect 153 78 187 112
rect 545 78 579 112
<< mvnsubdiff >>
rect 67 546 155 580
rect 189 546 223 580
rect 257 546 291 580
rect 325 546 359 580
rect 393 546 427 580
rect 461 546 495 580
rect 529 546 563 580
rect 597 546 631 580
rect 665 546 699 580
rect 733 546 767 580
rect 801 546 835 580
rect 869 546 903 580
rect 937 546 971 580
rect 1005 546 1039 580
rect 1073 546 1107 580
rect 1141 546 1175 580
rect 1209 546 1243 580
<< mvnsubdiffcont >>
rect 155 546 189 580
rect 223 546 257 580
rect 291 546 325 580
rect 359 546 393 580
rect 427 546 461 580
rect 495 546 529 580
rect 563 546 597 580
rect 631 546 665 580
rect 699 546 733 580
rect 767 546 801 580
rect 835 546 869 580
rect 903 546 937 580
rect 971 546 1005 580
rect 1039 546 1073 580
rect 1107 546 1141 580
rect 1175 546 1209 580
<< poly >>
rect 266 340 466 356
rect 266 306 282 340
rect 316 306 416 340
rect 450 306 466 340
rect 266 290 466 306
rect 266 232 466 248
rect 266 198 282 232
rect 316 198 416 232
rect 450 198 466 232
rect 266 182 466 198
rect 779 84 1035 100
rect 779 50 795 84
rect 829 50 890 84
rect 924 50 985 84
rect 1019 50 1035 84
rect 779 34 1035 50
rect 1091 84 1225 100
rect 1091 50 1107 84
rect 1141 50 1175 84
rect 1209 50 1225 84
rect 1091 34 1225 50
<< polycont >>
rect 282 306 316 340
rect 416 306 450 340
rect 282 198 316 232
rect 416 198 450 232
rect 795 50 829 84
rect 890 50 924 84
rect 985 50 1019 84
rect 1107 50 1141 84
rect 1175 50 1209 84
<< locali >>
rect 101 546 144 580
rect 189 546 221 580
rect 257 546 291 580
rect 331 546 359 580
rect 407 546 427 580
rect 483 546 495 580
rect 559 546 563 580
rect 597 546 601 580
rect 665 546 677 580
rect 733 546 753 580
rect 801 546 829 580
rect 869 546 903 580
rect 939 546 971 580
rect 1015 546 1039 580
rect 1091 546 1107 580
rect 1167 546 1175 580
rect 221 450 255 468
rect 153 434 255 450
rect 504 439 579 450
rect 187 430 255 434
rect 187 400 221 430
rect 153 396 221 400
rect 511 434 549 439
rect 511 405 545 434
rect 504 400 545 405
rect 153 384 238 396
rect 504 384 579 400
rect 734 348 768 398
rect 266 306 282 340
rect 316 339 416 340
rect 450 339 466 340
rect 316 306 377 339
rect 411 306 416 339
rect 411 305 449 306
rect 734 263 768 314
rect 266 198 282 232
rect 316 199 342 232
rect 376 199 414 233
rect 316 198 416 199
rect 450 198 466 232
rect 734 178 768 229
rect 153 116 221 128
rect 153 112 255 116
rect 187 78 255 112
rect 153 62 221 78
rect 890 348 924 398
rect 890 263 924 314
rect 890 178 924 229
rect 1046 348 1080 398
rect 1046 263 1080 314
rect 1046 178 1080 229
rect 1202 348 1236 398
rect 1202 263 1236 314
rect 1202 178 1236 229
rect 511 116 579 128
rect 477 112 579 116
rect 477 78 545 112
rect 511 62 579 78
rect 779 50 795 84
rect 840 50 890 84
rect 924 50 973 84
rect 1019 50 1035 84
rect 1091 50 1100 84
rect 1141 50 1172 84
rect 1209 50 1225 84
<< viali >>
rect 67 546 101 580
rect 144 546 155 580
rect 155 546 178 580
rect 221 546 223 580
rect 223 546 255 580
rect 297 546 325 580
rect 325 546 331 580
rect 373 546 393 580
rect 393 546 407 580
rect 449 546 461 580
rect 461 546 483 580
rect 525 546 529 580
rect 529 546 559 580
rect 601 546 631 580
rect 631 546 635 580
rect 677 546 699 580
rect 699 546 711 580
rect 753 546 767 580
rect 767 546 787 580
rect 829 546 835 580
rect 835 546 863 580
rect 905 546 937 580
rect 937 546 939 580
rect 981 546 1005 580
rect 1005 546 1015 580
rect 1057 546 1073 580
rect 1073 546 1091 580
rect 1133 546 1141 580
rect 1141 546 1167 580
rect 1209 546 1243 580
rect 221 468 255 502
rect 221 396 255 430
rect 477 405 511 439
rect 549 434 583 439
rect 549 405 579 434
rect 579 405 583 434
rect 734 398 768 432
rect 377 305 411 339
rect 449 306 450 339
rect 450 306 483 339
rect 449 305 483 306
rect 734 314 768 348
rect 342 199 376 233
rect 414 232 448 233
rect 414 199 416 232
rect 416 199 448 232
rect 734 229 768 263
rect 221 116 255 150
rect 221 44 255 78
rect 477 116 511 150
rect 734 144 768 178
rect 890 398 924 432
rect 890 314 924 348
rect 890 229 924 263
rect 890 144 924 178
rect 1046 398 1080 432
rect 1046 314 1080 348
rect 1046 229 1080 263
rect 1046 144 1080 178
rect 1202 398 1236 432
rect 1202 314 1236 348
rect 1202 229 1236 263
rect 1202 144 1236 178
rect 477 44 511 78
rect 806 50 829 84
rect 829 50 840 84
rect 890 50 924 84
rect 973 50 985 84
rect 985 50 1007 84
rect 1100 50 1107 84
rect 1107 50 1134 84
rect 1172 50 1175 84
rect 1175 50 1206 84
<< metal1 >>
rect 0 580 1310 647
rect 0 546 67 580
rect 101 546 144 580
rect 178 546 221 580
rect 255 546 297 580
rect 331 546 373 580
rect 407 546 449 580
rect 483 546 525 580
rect 559 546 601 580
rect 635 546 677 580
rect 711 546 753 580
rect 787 546 829 580
rect 863 546 905 580
rect 939 546 981 580
rect 1015 546 1057 580
rect 1091 546 1133 580
rect 1167 546 1209 580
rect 1243 546 1310 580
rect 0 502 1310 546
rect 0 501 221 502
tri 127 468 160 501 ne
rect 160 468 221 501
rect 255 501 1310 502
rect 255 468 261 501
tri 160 467 161 468 ne
rect 161 430 261 468
tri 261 467 295 501 nw
tri 694 467 728 501 ne
rect 161 396 221 430
rect 255 396 261 430
rect 161 150 261 396
rect 289 439 595 445
rect 289 405 477 439
rect 511 405 549 439
rect 583 405 595 439
rect 289 399 595 405
rect 728 432 774 501
tri 774 467 808 501 nw
tri 1006 467 1040 501 ne
rect 289 398 368 399
tri 368 398 369 399 nw
rect 728 398 734 432
rect 768 398 774 432
rect 289 263 335 398
tri 335 365 368 398 nw
rect 728 348 774 398
rect 365 339 540 348
rect 365 305 377 339
rect 411 305 449 339
rect 483 305 540 339
rect 365 296 540 305
tri 454 273 477 296 ne
rect 477 273 540 296
tri 335 263 345 273 sw
tri 477 263 487 273 ne
rect 487 263 540 273
rect 289 239 345 263
tri 345 239 369 263 sw
tri 487 262 488 263 ne
rect 289 233 460 239
rect 289 199 342 233
rect 376 199 414 233
rect 448 199 460 233
rect 289 193 460 199
tri 487 178 488 179 se
rect 488 178 540 263
rect 161 116 221 150
rect 255 116 261 150
rect 161 78 261 116
rect 161 44 221 78
rect 255 44 261 78
rect 161 32 261 44
tri 471 162 487 178 se
rect 487 162 540 178
rect 471 150 540 162
rect 471 116 477 150
rect 511 116 540 150
rect 728 314 734 348
rect 768 314 774 348
rect 728 263 774 314
rect 728 229 734 263
rect 768 229 774 263
rect 728 178 774 229
rect 728 144 734 178
rect 768 144 774 178
rect 728 132 774 144
rect 884 432 930 444
rect 884 398 890 432
rect 924 398 930 432
rect 884 348 930 398
rect 884 314 890 348
rect 924 314 930 348
rect 884 263 930 314
rect 884 229 890 263
rect 924 229 930 263
rect 884 178 930 229
rect 884 144 890 178
rect 924 144 930 178
rect 884 132 930 144
rect 1040 432 1086 501
tri 1086 467 1120 501 nw
rect 1040 398 1046 432
rect 1080 398 1086 432
rect 1040 348 1086 398
rect 1040 314 1046 348
rect 1080 314 1086 348
rect 1040 263 1086 314
rect 1040 229 1046 263
rect 1080 229 1086 263
rect 1040 178 1086 229
rect 1040 144 1046 178
rect 1080 144 1086 178
rect 1040 132 1086 144
rect 1196 432 1242 444
rect 1196 398 1202 432
rect 1236 398 1242 432
rect 1196 348 1242 398
rect 1196 314 1202 348
rect 1236 314 1242 348
rect 1196 263 1242 314
rect 1196 229 1202 263
rect 1236 229 1242 263
rect 1196 178 1242 229
rect 1196 144 1202 178
rect 1236 144 1242 178
rect 1196 132 1242 144
rect 471 90 540 116
tri 540 90 574 124 sw
rect 471 84 1019 90
rect 471 78 806 84
rect 471 44 477 78
rect 511 50 806 78
rect 840 50 890 84
rect 924 50 973 84
rect 1007 50 1019 84
rect 511 44 1019 50
rect 1088 84 1218 90
rect 1088 50 1100 84
rect 1134 50 1172 84
rect 1206 50 1218 84
rect 1088 44 1218 50
rect 471 32 1019 44
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_0
timestamp 1701704242
transform -1 0 195 0 1 66
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_1
timestamp 1701704242
transform 1 0 537 0 1 66
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_2
timestamp 1701704242
transform 1 0 145 0 1 388
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_3
timestamp 1701704242
transform 1 0 537 0 1 388
box 0 0 1 1
use pfet_CDNS_52468879185272  pfet_CDNS_52468879185272_0
timestamp 1701704242
transform 1 0 779 0 1 132
box -119 -66 375 366
use pfet_CDNS_52468879185674  pfet_CDNS_52468879185674_0
timestamp 1701704242
transform 1 0 1091 0 1 132
box -119 -66 219 366
use pfet_CDNS_52468879185675  pfet_CDNS_52468879185675_0
timestamp 1701704242
transform 1 0 266 0 1 388
box -119 -66 319 150
use pfet_CDNS_52468879185675  pfet_CDNS_52468879185675_1
timestamp 1701704242
transform 1 0 266 0 1 66
box -119 -66 319 150
<< properties >>
string GDS_END 7554956
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7544962
string path 31.725 14.075 1.025 14.075 
<< end >>
