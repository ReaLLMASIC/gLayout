magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 100 0 896 391
<< mvpdiff >>
rect 170 66 291 216
rect 705 66 826 216
<< mvnsubdiff >>
rect 167 290 217 324
rect 251 290 285 324
rect 319 290 353 324
rect 387 290 421 324
rect 455 290 489 324
rect 523 290 557 324
rect 591 290 625 324
rect 659 290 693 324
rect 727 290 761 324
rect 795 290 829 324
<< mvnsubdiffcont >>
rect 217 290 251 324
rect 285 290 319 324
rect 353 290 387 324
rect 421 290 455 324
rect 489 290 523 324
rect 557 290 591 324
rect 625 290 659 324
rect 693 290 727 324
rect 761 290 795 324
<< poly >>
rect 336 18 470 34
rect 336 -16 352 18
rect 386 -16 420 18
rect 454 -16 470 18
rect 336 -32 470 -16
rect 526 18 660 34
rect 526 -16 542 18
rect 576 -16 610 18
rect 644 -16 660 18
rect 526 -32 660 -16
<< polycont >>
rect 352 -16 386 18
rect 420 -16 454 18
rect 542 -16 576 18
rect 610 -16 644 18
<< locali >>
rect 201 290 217 324
rect 280 290 285 324
rect 319 290 325 324
rect 387 290 404 324
rect 455 290 483 324
rect 523 290 557 324
rect 595 290 625 324
rect 673 290 693 324
rect 751 290 761 324
rect 325 124 359 162
rect 481 132 515 170
rect 637 108 671 146
rect 336 -16 352 18
rect 393 -16 420 18
rect 465 -16 470 18
rect 526 -16 538 18
rect 576 -16 610 18
rect 644 -16 660 18
<< viali >>
rect 167 290 201 324
rect 246 290 251 324
rect 251 290 280 324
rect 325 290 353 324
rect 353 290 359 324
rect 404 290 421 324
rect 421 290 438 324
rect 483 290 489 324
rect 489 290 517 324
rect 561 290 591 324
rect 591 290 595 324
rect 639 290 659 324
rect 659 290 673 324
rect 717 290 727 324
rect 727 290 751 324
rect 795 290 829 324
rect 325 162 359 196
rect 325 90 359 124
rect 481 170 515 204
rect 481 98 515 132
rect 637 146 671 180
rect 637 74 671 108
rect 359 -16 386 18
rect 386 -16 393 18
rect 431 -16 454 18
rect 454 -16 465 18
rect 538 -16 542 18
rect 542 -16 572 18
rect 610 -16 644 18
<< metal1 >>
rect 155 324 841 391
rect 155 290 167 324
rect 201 290 246 324
rect 280 290 325 324
rect 359 290 404 324
rect 438 290 483 324
rect 517 290 561 324
rect 595 290 639 324
rect 673 290 717 324
rect 751 290 795 324
rect 829 290 841 324
rect 155 264 841 290
tri 441 230 475 264 ne
rect 319 196 368 208
tri 317 162 319 164 se
rect 319 162 325 196
rect 359 162 368 196
tri 301 146 317 162 se
rect 317 146 368 162
tri 287 132 301 146 se
rect 301 132 368 146
tri 285 130 287 132 se
rect 287 130 368 132
rect 240 78 246 130
rect 298 78 310 130
rect 362 78 368 130
rect 475 204 521 264
tri 521 230 555 264 nw
rect 475 170 481 204
rect 515 170 521 204
rect 475 132 521 170
rect 475 98 481 132
rect 515 98 521 132
rect 475 86 521 98
rect 631 180 677 192
rect 631 146 637 180
rect 671 146 677 180
rect 631 108 677 146
rect 631 74 637 108
rect 671 74 677 108
rect 631 62 677 74
rect 347 18 477 24
rect 347 -16 359 18
rect 393 -16 431 18
rect 465 -16 477 18
rect 347 -22 477 -16
rect 526 -25 532 27
rect 584 -25 596 27
rect 648 -25 656 27
<< via1 >>
rect 246 78 298 130
rect 310 124 362 130
rect 310 90 325 124
rect 325 90 359 124
rect 359 90 362 124
rect 310 78 362 90
rect 532 18 584 27
rect 532 -16 538 18
rect 538 -16 572 18
rect 572 -16 584 18
rect 532 -25 584 -16
rect 596 18 648 27
rect 596 -16 610 18
rect 610 -16 644 18
rect 644 -16 648 18
rect 596 -25 648 -16
<< metal2 >>
rect 240 78 246 130
rect 298 78 310 130
rect 362 78 578 130
tri 492 44 526 78 ne
rect 526 27 578 78
rect 526 -25 532 27
rect 584 -25 596 27
rect 648 -25 654 27
use pfet_CDNS_5246887918545  pfet_CDNS_5246887918545_0
timestamp 1701704242
transform 1 0 526 0 1 66
box -119 -66 219 216
use pfet_CDNS_5246887918545  pfet_CDNS_5246887918545_1
timestamp 1701704242
transform 1 0 370 0 1 66
box -119 -66 219 216
<< properties >>
string GDS_END 7541186
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7536114
string path 13.150 0.025 16.350 0.025 
<< end >>
