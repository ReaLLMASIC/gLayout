magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 737 53
<< metal1 >>
rect -6 53 743 56
rect -6 0 0 53
rect 737 0 743 53
rect -6 -3 743 0
<< properties >>
string GDS_END 95632190
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95629370
<< end >>
