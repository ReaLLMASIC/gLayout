magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 2332 781 4322 1654
rect 7321 -314 8420 -202
rect 7321 -480 8448 -314
rect 7321 -1154 8420 -480
rect 10032 -1154 10198 -22
<< pwell >>
rect 10072 -2454 10158 -1294
<< mvpsubdiff >>
rect 10098 -1344 10132 -1320
rect 10098 -1415 10132 -1378
rect 10098 -1486 10132 -1449
rect 10098 -1557 10132 -1520
rect 10098 -1628 10132 -1591
rect 10098 -1699 10132 -1662
rect 10098 -1770 10132 -1733
rect 10098 -1841 10132 -1804
rect 10098 -1912 10132 -1875
rect 10098 -1982 10132 -1946
rect 10098 -2052 10132 -2016
rect 10098 -2122 10132 -2086
rect 10098 -2192 10132 -2156
rect 10098 -2262 10132 -2226
rect 10098 -2428 10132 -2296
<< mvnsubdiff >>
rect 10098 -112 10132 -88
rect 10098 -183 10132 -146
rect 10098 -254 10132 -217
rect 10098 -325 10132 -288
rect 7588 -414 7612 -380
rect 7646 -414 7684 -380
rect 7718 -414 7756 -380
rect 7790 -414 7827 -380
rect 7861 -414 7898 -380
rect 7932 -414 7969 -380
rect 8003 -414 8040 -380
rect 8074 -414 8111 -380
rect 8145 -414 8182 -380
rect 8216 -414 8253 -380
rect 8287 -414 8324 -380
rect 8358 -414 8382 -380
rect 7588 -488 7622 -414
rect 8348 -488 8382 -414
rect 10098 -396 10132 -359
rect 10098 -467 10132 -430
rect 10098 -538 10132 -501
rect 10098 -609 10132 -572
rect 10098 -680 10132 -643
rect 10098 -750 10132 -714
rect 10098 -820 10132 -784
rect 10098 -890 10132 -854
rect 10098 -960 10132 -924
rect 10098 -1030 10132 -994
rect 10098 -1088 10132 -1064
<< mvpsubdiffcont >>
rect 10098 -1378 10132 -1344
rect 10098 -1449 10132 -1415
rect 10098 -1520 10132 -1486
rect 10098 -1591 10132 -1557
rect 10098 -1662 10132 -1628
rect 10098 -1733 10132 -1699
rect 10098 -1804 10132 -1770
rect 10098 -1875 10132 -1841
rect 10098 -1946 10132 -1912
rect 10098 -2016 10132 -1982
rect 10098 -2086 10132 -2052
rect 10098 -2156 10132 -2122
rect 10098 -2226 10132 -2192
rect 10098 -2296 10132 -2262
<< mvnsubdiffcont >>
rect 10098 -146 10132 -112
rect 10098 -217 10132 -183
rect 10098 -288 10132 -254
rect 10098 -359 10132 -325
rect 7612 -414 7646 -380
rect 7684 -414 7718 -380
rect 7756 -414 7790 -380
rect 7827 -414 7861 -380
rect 7898 -414 7932 -380
rect 7969 -414 8003 -380
rect 8040 -414 8074 -380
rect 8111 -414 8145 -380
rect 8182 -414 8216 -380
rect 8253 -414 8287 -380
rect 8324 -414 8358 -380
rect 10098 -430 10132 -396
rect 10098 -501 10132 -467
rect 10098 -572 10132 -538
rect 10098 -643 10132 -609
rect 10098 -714 10132 -680
rect 10098 -784 10132 -750
rect 10098 -854 10132 -820
rect 10098 -924 10132 -890
rect 10098 -994 10132 -960
rect 10098 -1064 10132 -1030
<< locali >>
rect 10098 -112 10132 -88
rect 10098 -183 10132 -146
rect 10098 -254 10132 -217
rect 10098 -325 10132 -288
rect 7588 -414 7612 -380
rect 7646 -414 7684 -380
rect 7718 -414 7756 -380
rect 7790 -414 7827 -380
rect 7861 -414 7898 -380
rect 7932 -414 7969 -380
rect 8003 -414 8040 -380
rect 8074 -414 8111 -380
rect 8145 -414 8182 -380
rect 8216 -414 8253 -380
rect 8287 -414 8324 -380
rect 8358 -414 8382 -380
rect 7588 -488 7622 -414
rect 8348 -488 8382 -414
rect 10098 -396 10132 -359
rect 10098 -467 10132 -430
rect 10098 -538 10132 -501
rect 10098 -609 10132 -572
rect 10098 -680 10132 -643
rect 10098 -750 10132 -714
rect 10098 -812 10132 -784
rect 10098 -884 10132 -854
rect 10098 -956 10132 -924
rect 10098 -1030 10132 -994
rect 7842 -1070 7880 -1036
rect 7989 -1124 8303 -1068
rect 10098 -1088 10132 -1064
rect 7989 -1164 8045 -1124
rect 9078 -1154 9116 -1120
rect 9150 -1154 9188 -1120
rect 9222 -1154 9260 -1120
rect 9294 -1154 9332 -1120
rect 9366 -1154 9404 -1120
rect 9438 -1154 9476 -1120
rect 8149 -1198 8187 -1164
rect 9690 -1170 9728 -1136
rect 8823 -1238 8861 -1204
rect 8789 -1244 8895 -1238
rect 8985 -1238 9023 -1204
rect 9806 -1227 9840 -1197
rect 8951 -1278 9157 -1238
rect 9342 -1278 9425 -1244
rect 10098 -1326 10132 -1320
rect 10092 -1338 10138 -1326
rect 10092 -1378 10098 -1338
rect 10132 -1378 10138 -1338
rect 10092 -1410 10138 -1378
rect 10092 -1449 10098 -1410
rect 10132 -1449 10138 -1410
rect 10092 -1482 10138 -1449
rect 10092 -1520 10098 -1482
rect 10132 -1520 10138 -1482
rect 8056 -1594 8090 -1524
rect 10092 -1528 10138 -1520
rect 10098 -1557 10132 -1528
rect 10098 -1628 10132 -1604
rect 10098 -1699 10132 -1676
rect 10098 -1770 10132 -1748
rect 10098 -1841 10132 -1820
rect 10098 -1912 10132 -1875
rect 8266 -2007 8304 -1973
rect 8232 -2066 8338 -2007
rect 10098 -1982 10132 -1946
rect 10098 -2052 10132 -2016
rect 10092 -2086 10098 -2078
rect 10132 -2086 10138 -2078
rect 10092 -2122 10138 -2086
rect 10092 -2168 10098 -2122
rect 10132 -2168 10138 -2122
rect 10092 -2192 10138 -2168
rect 10092 -2240 10098 -2192
rect 10132 -2240 10138 -2192
rect 10092 -2262 10138 -2240
rect 10092 -2312 10098 -2262
rect 10132 -2312 10138 -2262
rect 10092 -2324 10138 -2312
rect 10098 -2428 10132 -2324
rect 8125 -2500 8163 -2466
rect 8388 -2484 8426 -2450
rect 8670 -2566 8708 -2532
rect 9223 -2566 9261 -2532
rect 9555 -2767 9589 -2729
rect 9083 -2828 9132 -2790
rect 9555 -2839 9589 -2801
rect 8062 -2946 8096 -2908
rect 9555 -2911 9589 -2873
rect 9199 -3235 9233 -3197
<< viali >>
rect 10098 -820 10132 -812
rect 10098 -846 10132 -820
rect 10098 -890 10132 -884
rect 10098 -918 10132 -890
rect 10098 -960 10132 -956
rect 10098 -990 10132 -960
rect 7808 -1070 7842 -1036
rect 7880 -1070 7914 -1036
rect 9044 -1154 9078 -1120
rect 9116 -1154 9150 -1120
rect 9188 -1154 9222 -1120
rect 9260 -1154 9294 -1120
rect 9332 -1154 9366 -1120
rect 9404 -1154 9438 -1120
rect 9476 -1154 9510 -1120
rect 8115 -1198 8149 -1164
rect 8187 -1198 8221 -1164
rect 9656 -1170 9690 -1136
rect 9728 -1170 9762 -1136
rect 8789 -1238 8823 -1204
rect 8861 -1238 8895 -1204
rect 8951 -1238 8985 -1204
rect 9023 -1238 9057 -1204
rect 10098 -1344 10132 -1338
rect 10098 -1372 10132 -1344
rect 10098 -1415 10132 -1410
rect 10098 -1444 10132 -1415
rect 10098 -1486 10132 -1482
rect 10098 -1516 10132 -1486
rect 10098 -1591 10132 -1570
rect 10098 -1604 10132 -1591
rect 10098 -1662 10132 -1642
rect 10098 -1676 10132 -1662
rect 10098 -1733 10132 -1714
rect 10098 -1748 10132 -1733
rect 10098 -1804 10132 -1786
rect 10098 -1820 10132 -1804
rect 8232 -2007 8266 -1973
rect 8304 -2007 8338 -1973
rect 10098 -2156 10132 -2134
rect 10098 -2168 10132 -2156
rect 10098 -2226 10132 -2206
rect 10098 -2240 10132 -2226
rect 10098 -2296 10132 -2278
rect 10098 -2312 10132 -2296
rect 8091 -2500 8125 -2466
rect 8163 -2500 8197 -2466
rect 8354 -2484 8388 -2450
rect 8426 -2484 8460 -2450
rect 8636 -2566 8670 -2532
rect 8708 -2566 8742 -2532
rect 9189 -2566 9223 -2532
rect 9261 -2566 9295 -2532
rect 9555 -2729 9589 -2695
rect 9555 -2801 9589 -2767
rect 9555 -2873 9589 -2839
rect 8062 -2908 8096 -2874
rect 9555 -2945 9589 -2911
rect 8062 -2980 8096 -2946
rect 9199 -3197 9233 -3163
rect 9199 -3269 9233 -3235
<< metal1 >>
tri 9616 -10 9623 -3 ne
rect 9623 -10 9629 42
rect 9681 -10 9693 42
rect 9745 -10 9751 42
tri 9751 -10 9758 -3 nw
tri 8586 -574 8598 -562 se
rect 8598 -574 9032 -562
tri 7684 -598 7708 -574 se
rect 7708 -598 9032 -574
rect 7611 -614 9032 -598
rect 9084 -614 9096 -562
rect 9148 -614 9154 -562
rect 7611 -626 8610 -614
tri 8610 -626 8622 -614 nw
rect 6491 -1002 7545 -800
rect 9560 -812 10364 -800
rect 9560 -846 10098 -812
rect 10132 -846 10364 -812
rect 9560 -884 10364 -846
rect 9560 -918 10098 -884
rect 10132 -918 10364 -884
rect 9560 -956 10364 -918
rect 9560 -990 10098 -956
rect 10132 -990 10364 -956
rect 9560 -1002 10364 -990
rect 7796 -1036 9774 -1030
rect 7796 -1070 7808 -1036
rect 7842 -1070 7880 -1036
rect 7914 -1070 9774 -1036
rect 7796 -1076 9774 -1070
tri 9619 -1101 9644 -1076 ne
tri 8372 -1120 8385 -1107 se
rect 8385 -1120 8391 -1107
tri 8338 -1154 8372 -1120 se
rect 8372 -1154 8391 -1120
tri 8334 -1158 8338 -1154 se
rect 8338 -1158 8391 -1154
rect 8103 -1159 8391 -1158
rect 8443 -1159 8455 -1107
rect 8507 -1114 8939 -1107
tri 8939 -1114 8946 -1107 sw
rect 8507 -1120 8946 -1114
tri 8946 -1120 8952 -1114 sw
rect 9032 -1120 9522 -1114
rect 8507 -1154 8952 -1120
tri 8952 -1154 8986 -1120 sw
rect 9032 -1154 9044 -1120
rect 9078 -1122 9116 -1120
rect 9150 -1122 9188 -1120
rect 9078 -1154 9102 -1122
rect 9154 -1154 9188 -1122
rect 9222 -1154 9260 -1120
rect 9294 -1154 9332 -1120
rect 9366 -1154 9404 -1120
rect 9438 -1154 9476 -1120
rect 9510 -1154 9522 -1120
rect 8507 -1159 8986 -1154
tri 8986 -1159 8991 -1154 sw
rect 8103 -1164 8388 -1159
rect 8103 -1198 8115 -1164
rect 8149 -1198 8187 -1164
rect 8221 -1170 8388 -1164
tri 8388 -1170 8399 -1159 nw
tri 8914 -1170 8925 -1159 ne
rect 8925 -1160 8991 -1159
tri 8991 -1160 8992 -1159 sw
rect 9032 -1160 9102 -1154
rect 8925 -1170 8992 -1160
tri 8992 -1170 9002 -1160 sw
tri 9077 -1170 9087 -1160 ne
rect 9087 -1170 9102 -1160
rect 8221 -1192 8366 -1170
tri 8366 -1192 8388 -1170 nw
tri 8925 -1184 8939 -1170 ne
rect 8939 -1192 9002 -1170
tri 9002 -1192 9024 -1170 sw
tri 9087 -1185 9102 -1170 ne
rect 9154 -1160 9522 -1154
rect 9644 -1136 9774 -1076
rect 9154 -1170 9169 -1160
tri 9169 -1170 9179 -1160 nw
rect 9644 -1170 9656 -1136
rect 9690 -1170 9728 -1136
rect 9762 -1170 9774 -1136
rect 9154 -1174 9163 -1170
rect 9102 -1176 9163 -1174
tri 9163 -1176 9169 -1170 nw
rect 9644 -1176 9774 -1170
rect 9102 -1186 9154 -1176
tri 9154 -1185 9163 -1176 nw
rect 8221 -1198 8354 -1192
rect 8103 -1204 8354 -1198
tri 8354 -1204 8366 -1192 nw
rect 8577 -1244 8707 -1238
rect 8777 -1244 8783 -1192
rect 8835 -1244 8847 -1192
rect 8899 -1244 8907 -1192
rect 8939 -1204 9069 -1192
rect 8939 -1238 8951 -1204
rect 8985 -1238 9023 -1204
rect 9057 -1238 9069 -1204
rect 8939 -1244 9069 -1238
rect 9102 -1244 9154 -1238
rect 8577 -1292 8587 -1244
rect 8639 -1296 8651 -1244
rect 8703 -1292 8707 -1244
tri 8707 -1272 8732 -1247 sw
tri 9175 -1272 9199 -1248 se
rect 9199 -1272 9329 -1248
rect 8587 -1302 8703 -1296
rect 8953 -1302 8994 -1272
rect 9736 -1338 10344 -1326
rect 9736 -1372 10098 -1338
rect 10132 -1372 10344 -1338
rect 9736 -1410 10344 -1372
rect 9736 -1444 10098 -1410
rect 10132 -1444 10344 -1410
rect 9736 -1482 10344 -1444
rect 9736 -1516 10098 -1482
rect 10132 -1516 10344 -1482
rect 9736 -1528 10344 -1516
tri 10053 -1561 10086 -1528 ne
rect 10086 -1570 10144 -1528
tri 10144 -1562 10178 -1528 nw
tri 7544 -1642 7555 -1631 se
rect 7555 -1642 8405 -1588
rect 10086 -1604 10098 -1570
rect 10132 -1604 10144 -1570
tri 8405 -1642 8416 -1631 sw
tri 10075 -1642 10086 -1631 se
rect 10086 -1642 10144 -1604
tri 7530 -1656 7544 -1642 se
rect 7544 -1656 8416 -1642
tri 8416 -1656 8430 -1642 sw
tri 10061 -1656 10075 -1642 se
rect 10075 -1656 10098 -1642
rect 7509 -1708 9629 -1656
rect 9681 -1708 9693 -1656
rect 9745 -1676 10098 -1656
rect 10132 -1676 10144 -1642
rect 9745 -1708 10144 -1676
rect 7509 -1714 10144 -1708
rect 7509 -1722 10098 -1714
tri 10061 -1747 10086 -1722 ne
rect 10086 -1748 10098 -1722
rect 10132 -1748 10144 -1714
rect 10086 -1786 10144 -1748
rect 10086 -1820 10098 -1786
rect 10132 -1820 10144 -1786
rect 10086 -1826 10144 -1820
rect 8050 -1967 8102 -1961
tri 8025 -2038 8050 -2013 ne
rect 8220 -1973 8350 -1961
rect 8220 -2007 8232 -1973
rect 8266 -2007 8304 -1973
rect 8338 -2007 8350 -1973
rect 8220 -2013 8350 -2007
rect 8102 -2018 8122 -2013
tri 8122 -2018 8127 -2013 nw
rect 8540 -2018 8546 -1966
rect 8598 -2018 8610 -1966
rect 8662 -1972 9595 -1966
rect 8662 -2018 9543 -1972
rect 8050 -2031 8102 -2019
tri 8102 -2038 8122 -2018 nw
tri 9518 -2038 9538 -2018 ne
rect 9538 -2024 9543 -2018
rect 9538 -2036 9595 -2024
rect 9538 -2038 9543 -2036
tri 9538 -2043 9543 -2038 ne
rect 8050 -2089 8102 -2083
rect 9543 -2094 9595 -2088
tri 10081 -2094 10086 -2089 se
rect 10086 -2094 10144 -2042
tri 10053 -2122 10081 -2094 se
rect 10081 -2122 10144 -2094
tri 10144 -2122 10178 -2088 sw
rect 9736 -2134 10344 -2122
rect 9736 -2168 10098 -2134
rect 10132 -2168 10344 -2134
rect 9736 -2206 10344 -2168
rect 9736 -2240 10098 -2206
rect 10132 -2240 10344 -2206
rect 9736 -2278 10344 -2240
rect 9736 -2312 10098 -2278
rect 10132 -2312 10344 -2278
rect 9736 -2324 10344 -2312
rect 8342 -2404 8546 -2352
rect 8598 -2404 8610 -2352
rect 8662 -2404 8668 -2352
rect 8342 -2450 8472 -2404
tri 8472 -2429 8497 -2404 nw
rect 9500 -2437 9629 -2385
rect 9681 -2437 9693 -2385
rect 9745 -2437 10030 -2385
rect 10082 -2437 10094 -2385
rect 10146 -2437 10152 -2385
rect 8079 -2466 8209 -2460
rect 8079 -2500 8091 -2466
rect 8125 -2500 8163 -2466
rect 8197 -2500 8209 -2466
rect 8342 -2484 8354 -2450
rect 8388 -2484 8426 -2450
rect 8460 -2484 8472 -2450
rect 8342 -2490 8472 -2484
rect 8079 -2506 8209 -2500
tri 8209 -2506 8221 -2494 sw
rect 8079 -2508 8221 -2506
tri 8221 -2508 8223 -2506 sw
rect 8079 -2519 8223 -2508
tri 8223 -2519 8234 -2508 sw
rect 8540 -2514 9307 -2508
rect 8079 -2571 8283 -2519
rect 8335 -2571 8347 -2519
rect 8399 -2571 8405 -2519
rect 8540 -2532 8699 -2514
rect 8540 -2566 8636 -2532
rect 8670 -2566 8699 -2532
rect 8751 -2566 8763 -2514
rect 8815 -2566 8827 -2514
rect 8879 -2566 8891 -2514
rect 8943 -2566 8955 -2514
rect 9007 -2532 9307 -2514
rect 9007 -2566 9189 -2532
rect 9223 -2566 9261 -2532
rect 9295 -2566 9307 -2532
rect 8540 -2572 9307 -2566
rect 9261 -2788 9298 -2600
rect 9070 -2834 9298 -2788
rect 9543 -2695 9595 -2683
rect 9543 -2707 9555 -2695
rect 9589 -2707 9595 -2695
rect 9543 -2767 9595 -2759
rect 9543 -2771 9555 -2767
rect 9589 -2771 9595 -2767
rect 9543 -2835 9595 -2823
rect 8050 -2868 8102 -2862
rect 8050 -2932 8102 -2920
rect 9543 -2899 9595 -2887
rect 9543 -2957 9595 -2951
rect 8050 -2992 8102 -2984
rect 9971 -3039 10344 -2641
rect 9280 -3118 9314 -3083
tri 9181 -3163 9193 -3151 se
rect 9193 -3163 9239 -3151
tri 9165 -3179 9181 -3163 se
rect 9181 -3179 9199 -3163
rect 8277 -3231 8283 -3179
rect 8335 -3231 8347 -3179
rect 8399 -3197 9199 -3179
rect 9233 -3197 9239 -3163
rect 8399 -3231 9239 -3197
tri 9166 -3235 9170 -3231 ne
rect 9170 -3235 9239 -3231
tri 9170 -3258 9193 -3235 ne
rect 9193 -3269 9199 -3235
rect 9233 -3269 9239 -3235
rect 9193 -3281 9239 -3269
rect 8066 -3288 9060 -3282
rect 8066 -3340 8700 -3288
rect 8752 -3340 8764 -3288
rect 8816 -3340 8828 -3288
rect 8880 -3340 8892 -3288
rect 8944 -3340 8956 -3288
rect 9008 -3340 9060 -3288
rect 8066 -3346 9060 -3340
<< via1 >>
rect 9629 -10 9681 42
rect 9693 -10 9745 42
rect 9032 -614 9084 -562
rect 9096 -614 9148 -562
rect 8391 -1159 8443 -1107
rect 8455 -1159 8507 -1107
rect 9102 -1154 9116 -1122
rect 9116 -1154 9150 -1122
rect 9150 -1154 9154 -1122
rect 9102 -1174 9154 -1154
rect 8783 -1204 8835 -1192
rect 8783 -1238 8789 -1204
rect 8789 -1238 8823 -1204
rect 8823 -1238 8835 -1204
rect 8783 -1244 8835 -1238
rect 8847 -1204 8899 -1192
rect 8847 -1238 8861 -1204
rect 8861 -1238 8895 -1204
rect 8895 -1238 8899 -1204
rect 8847 -1244 8899 -1238
rect 9102 -1238 9154 -1186
rect 8587 -1296 8639 -1244
rect 8651 -1296 8703 -1244
rect 9629 -1708 9681 -1656
rect 9693 -1708 9745 -1656
rect 8050 -2019 8102 -1967
rect 8546 -2018 8598 -1966
rect 8610 -2018 8662 -1966
rect 8050 -2083 8102 -2031
rect 9543 -2024 9595 -1972
rect 9543 -2088 9595 -2036
rect 8546 -2404 8598 -2352
rect 8610 -2404 8662 -2352
rect 9629 -2437 9681 -2385
rect 9693 -2437 9745 -2385
rect 10030 -2437 10082 -2385
rect 10094 -2437 10146 -2385
rect 8283 -2571 8335 -2519
rect 8347 -2571 8399 -2519
rect 8699 -2532 8751 -2514
rect 8699 -2566 8708 -2532
rect 8708 -2566 8742 -2532
rect 8742 -2566 8751 -2532
rect 8763 -2566 8815 -2514
rect 8827 -2566 8879 -2514
rect 8891 -2566 8943 -2514
rect 8955 -2566 9007 -2514
rect 9543 -2729 9555 -2707
rect 9555 -2729 9589 -2707
rect 9589 -2729 9595 -2707
rect 9543 -2759 9595 -2729
rect 9543 -2801 9555 -2771
rect 9555 -2801 9589 -2771
rect 9589 -2801 9595 -2771
rect 9543 -2823 9595 -2801
rect 9543 -2839 9595 -2835
rect 8050 -2874 8102 -2868
rect 8050 -2908 8062 -2874
rect 8062 -2908 8096 -2874
rect 8096 -2908 8102 -2874
rect 8050 -2920 8102 -2908
rect 8050 -2946 8102 -2932
rect 8050 -2980 8062 -2946
rect 8062 -2980 8096 -2946
rect 8096 -2980 8102 -2946
rect 9543 -2873 9555 -2839
rect 9555 -2873 9589 -2839
rect 9589 -2873 9595 -2839
rect 9543 -2887 9595 -2873
rect 9543 -2911 9595 -2899
rect 9543 -2945 9555 -2911
rect 9555 -2945 9589 -2911
rect 9589 -2945 9595 -2911
rect 9543 -2951 9595 -2945
rect 8050 -2984 8102 -2980
rect 8283 -3231 8335 -3179
rect 8347 -3231 8399 -3179
rect 8700 -3340 8752 -3288
rect 8764 -3340 8816 -3288
rect 8828 -3340 8880 -3288
rect 8892 -3340 8944 -3288
rect 8956 -3340 9008 -3288
<< metal2 >>
rect 4335 -20 4378 34
rect 6491 -1059 6807 1763
rect 10024 1761 10344 1762
tri 10024 1745 10040 1761 ne
rect 10040 1745 10344 1761
rect 7235 -2802 7551 1745
rect 8385 -1107 8513 -25
rect 8385 -1159 8391 -1107
rect 8443 -1159 8455 -1107
rect 8507 -1159 8513 -1107
rect 8577 -1244 8705 -472
tri 8795 -1174 8808 -1161 se
rect 8808 -1174 8872 473
rect 9623 42 9751 1745
tri 10040 1726 10059 1745 ne
rect 9623 -10 9629 42
rect 9681 -10 9693 42
rect 9745 -10 9751 42
rect 9026 -614 9032 -562
rect 9084 -614 9096 -562
rect 9148 -614 9154 -562
tri 9026 -690 9102 -614 ne
rect 9102 -1122 9154 -614
tri 8872 -1174 8885 -1161 sw
tri 8783 -1186 8795 -1174 se
rect 8795 -1186 8885 -1174
tri 8885 -1186 8897 -1174 sw
rect 9102 -1186 9154 -1174
tri 8777 -1192 8783 -1186 se
rect 8783 -1192 8897 -1186
tri 8897 -1192 8903 -1186 sw
rect 8777 -1244 8783 -1192
rect 8835 -1244 8847 -1192
rect 8899 -1244 8905 -1192
rect 9102 -1244 9154 -1238
rect 8577 -1296 8587 -1244
rect 8639 -1296 8651 -1244
rect 8703 -1296 8705 -1244
rect 8577 -1302 8705 -1296
rect 9623 -1656 9751 -10
rect 9623 -1708 9629 -1656
rect 9681 -1708 9693 -1656
rect 9745 -1708 9751 -1656
rect 8050 -1967 8102 -1961
rect 8050 -2031 8102 -2019
rect 8050 -2868 8102 -2083
rect 8540 -2018 8546 -1966
rect 8598 -2018 8610 -1966
rect 8662 -2018 8668 -1966
rect 8540 -2352 8668 -2018
rect 9543 -1972 9595 -1966
rect 9543 -2036 9595 -2024
rect 8540 -2404 8546 -2352
rect 8598 -2404 8610 -2352
rect 8662 -2404 8668 -2352
rect 8696 -2514 9012 -2306
rect 8050 -2932 8102 -2920
rect 8050 -2990 8102 -2984
rect 8277 -2571 8283 -2519
rect 8335 -2571 8347 -2519
rect 8399 -2571 8405 -2519
rect -183 -3174 -143 -3128
rect 8277 -3179 8405 -2571
rect 8277 -3231 8283 -3179
rect 8335 -3231 8347 -3179
rect 8399 -3231 8405 -3179
rect 8696 -2566 8699 -2514
rect 8751 -2566 8763 -2514
rect 8815 -2566 8827 -2514
rect 8879 -2566 8891 -2514
rect 8943 -2566 8955 -2514
rect 9007 -2566 9012 -2514
rect 8696 -3288 9012 -2566
rect 9543 -2707 9595 -2088
rect 9623 -2385 9751 -1708
rect 9623 -2437 9629 -2385
rect 9681 -2437 9693 -2385
rect 9745 -2437 9751 -2385
tri 10024 347 10059 382 se
rect 10059 347 10344 1745
rect 10024 -2385 10344 347
rect 10024 -2437 10030 -2385
rect 10082 -2437 10094 -2385
rect 10146 -2437 10344 -2385
rect 10024 -2703 10344 -2437
rect 9543 -2771 9595 -2759
rect 9543 -2835 9595 -2823
rect 9543 -2899 9595 -2887
rect 9543 -2957 9595 -2951
rect 8696 -3340 8700 -3288
rect 8752 -3340 8764 -3288
rect 8816 -3340 8828 -3288
rect 8880 -3340 8892 -3288
rect 8944 -3340 8956 -3288
rect 9008 -3340 9012 -3288
rect 8696 -3346 9012 -3340
rect -183 -3429 -143 -3383
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 9233 -1 0 -3163
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 8096 -1 0 -2874
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 9762 0 1 -1170
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 7914 0 1 -1070
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 9057 0 1 -1238
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform -1 0 8895 0 1 -1238
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform -1 0 8742 0 1 -2566
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform -1 0 9295 0 1 -2566
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform -1 0 8338 0 1 -2007
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform -1 0 8197 0 -1 -2466
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 1 0 8115 0 1 -1198
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 1 0 8354 0 1 -2484
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 10132 -1 0 -812
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1701704242
transform 1 0 7567 0 1 -1628
box -12 -6 838 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1701704242
transform 0 -1 9589 1 0 -2945
box 0 0 1 1
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1701704242
transform 1 0 9512 0 1 -2428
box -12 -6 622 40
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1701704242
transform -1 0 9510 0 1 -1154
box 0 0 1 1
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1701704242
transform -1 0 9048 0 1 -3332
box -12 -6 982 40
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1701704242
transform 1 0 10098 0 -1 -1570
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 9154 -1 0 -1116
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 8102 -1 0 -2862
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 9595 -1 0 -1966
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 1 8050 -1 0 -1961
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform -1 0 8513 0 1 -1159
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform -1 0 8905 0 1 -1244
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform -1 0 8405 0 1 -2571
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform -1 0 8405 0 1 -3231
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 1 0 9623 0 -1 42
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 1 0 9026 0 -1 -562
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 1 0 9623 0 -1 -2385
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 1 0 10024 0 -1 -2385
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 1 0 9623 0 1 -1708
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 1 0 8540 0 1 -2404
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 1 0 8540 0 1 -2018
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1701704242
transform 0 -1 9595 -1 0 -2701
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 0 1 8587 1 0 -1302
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_0
timestamp 1701704242
transform 0 1 8699 -1 0 -2508
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_1
timestamp 1701704242
transform 0 1 8700 1 0 -3346
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1701704242
transform -1 0 10281 0 -1 636
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1701704242
transform -1 0 10281 0 -1 1089
box 0 0 192 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1701704242
transform -1 0 10344 0 -1 -2134
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1701704242
transform -1 0 10344 0 -1 -1336
box 0 0 320 180
use M1M2_CDNS_524688791851176  M1M2_CDNS_524688791851176_0
timestamp 1701704242
transform 0 1 6491 -1 0 -803
box 0 0 256 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_0
timestamp 1701704242
transform 0 1 7239 -1 0 -2605
box 0 0 192 308
use M1M2_CDNS_524688791851200  M1M2_CDNS_524688791851200_0
timestamp 1701704242
transform -1 0 10344 0 -1 -2646
box 0 0 320 372
use sky130_fd_io__sio_com_inbuf_einv  sky130_fd_io__sio_com_inbuf_einv_0
timestamp 1701704242
transform 0 -1 10191 -1 0 -2464
box -27 -66 904 2202
use sky130_fd_io__sio_com_inbuf_einv_hv  sky130_fd_io__sio_com_inbuf_einv_hv_0
timestamp 1701704242
transform -1 0 10024 0 1 -2411
box -128 -43 1634 2389
use sky130_fd_io__sio_gpio_in_buf  sky130_fd_io__sio_gpio_in_buf_0
timestamp 1701704242
transform 1 0 167 0 1 64
box -423 -1390 10151 3581
use sky130_fd_io__sio_inbuf_hvinv_x1  sky130_fd_io__sio_inbuf_hvinv_x1_0
timestamp 1701704242
transform 1 0 8073 0 1 -1548
box -91 -106 403 1126
use sky130_fd_io__sio_inbuf_hvinv_x2  sky130_fd_io__sio_inbuf_hvinv_x2_0
timestamp 1701704242
transform -1 0 8073 0 1 -1548
box -91 -106 579 1126
use sky130_fd_io__sio_inbuf_ls  sky130_fd_io__sio_inbuf_ls_0
timestamp 1701704242
transform -1 0 9369 0 -1 -1228
box -43 -24 1345 1574
<< labels >>
flabel comment s 9383 -1158 9383 -1158 0 FreeSans 400 0 0 0 en_h_n
flabel comment s 9305 -3065 9305 -3065 0 FreeSans 200 0 0 0 ibufmux_out_n
flabel metal1 s 8664 -2690 8664 -2690 0 FreeSans 440 0 0 0 vpwr_ka
flabel metal1 s 8953 -1302 8994 -1272 0 FreeSans 200 180 0 0 en_h
port 2 nsew
flabel metal1 s 7708 -626 7750 -574 3 FreeSans 200 0 0 0 en_h_n
port 3 nsew
flabel metal1 s 8399 -2396 8432 -2363 0 FreeSans 200 0 0 0 en
port 4 nsew
flabel metal1 s 9280 -3118 9314 -3083 0 FreeSans 200 0 0 0 ibufmux_out_n
port 5 nsew
flabel metal1 s 8728 -3327 8756 -3300 0 FreeSans 200 0 0 0 vpb_ka
port 7 nsew
flabel metal1 s 8265 -2008 8304 -1973 0 FreeSans 200 0 0 0 en_n
port 6 nsew
flabel locali s 9806 -1227 9840 -1197 0 FreeSans 200 0 0 0 ibufmux_out_h_n
port 8 nsew
flabel metal2 s 6491 1692 6799 1745 0 FreeSans 200 0 0 0 vcc_io
port 9 nsew
flabel metal2 s 7235 1692 7551 1744 0 FreeSans 200 0 0 0 vpwr_ka
port 10 nsew
flabel metal2 s 10059 1692 10344 1744 0 FreeSans 200 0 0 0 vgnd
port 11 nsew
flabel metal2 s 4335 -20 4378 34 0 FreeSans 200 0 0 0 vtrip_sel_h_n
port 12 nsew
flabel metal2 s -183 -3429 -143 -3383 3 FreeSans 200 0 0 0 in_vt
port 13 nsew
flabel metal2 s -183 -3174 -143 -3128 3 FreeSans 200 0 0 0 in_h
port 14 nsew
<< properties >>
string GDS_END 85791658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85776970
string path 189.050 -9.925 210.200 -9.925 
<< end >>
