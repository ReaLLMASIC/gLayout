magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 15552 2653 15925 3354
<< pwell >>
rect 14668 836 14842 1246
<< psubdiff >>
rect 14694 1196 14816 1220
rect 14728 1162 14782 1196
rect 14694 1104 14816 1162
rect 14728 1070 14782 1104
rect 14694 1012 14816 1070
rect 14728 978 14782 1012
rect 14694 920 14816 978
rect 14728 886 14782 920
rect 14694 862 14816 886
<< psubdiffcont >>
rect 14694 1162 14728 1196
rect 14782 1162 14816 1196
rect 14694 1070 14728 1104
rect 14782 1070 14816 1104
rect 14694 978 14728 1012
rect 14782 978 14816 1012
rect 14694 886 14728 920
rect 14782 886 14816 920
<< locali >>
rect 14694 1196 14816 1220
rect 14728 1162 14782 1196
rect 14694 1104 14816 1162
rect 14728 1070 14782 1104
rect 14694 1012 14816 1070
rect 14728 978 14782 1012
rect 14694 920 14816 978
rect 14728 894 14782 920
rect 14728 860 14776 894
rect 14810 862 14816 886
rect 14694 822 14810 860
rect 14728 788 14776 822
<< viali >>
rect 14694 886 14728 894
rect 14694 860 14728 886
rect 14776 886 14782 894
rect 14782 886 14810 894
rect 14776 860 14810 886
rect 14694 788 14728 822
rect 14776 788 14810 822
<< metal1 >>
rect 2949 3060 3189 3066
rect 2949 3008 3049 3060
rect 3101 3008 3137 3060
rect 2949 2978 3189 3008
rect 2949 2926 3049 2978
rect 3101 2926 3137 2978
rect 2949 2895 3189 2926
rect 2649 2823 2726 2855
rect 2949 2843 3049 2895
rect 3101 2843 3137 2895
rect 2949 2812 3189 2843
rect 2949 2760 3049 2812
rect 3101 2760 3137 2812
rect 2949 2754 3189 2760
tri 14341 2154 14415 2228 se
rect 14415 2222 14940 2228
rect 14415 2176 14888 2222
tri 14415 2154 14437 2176 nw
tri 14856 2154 14878 2176 ne
rect 14878 2170 14888 2176
rect 14878 2158 14940 2170
rect 14878 2154 14888 2158
tri 14336 2149 14341 2154 se
rect 14341 2149 14410 2154
tri 14410 2149 14415 2154 nw
tri 14878 2149 14883 2154 ne
rect 14883 2149 14888 2154
rect 883 2097 889 2149
rect 941 2097 953 2149
rect 1005 2097 2759 2149
rect 2811 2097 2823 2149
rect 2875 2097 5667 2149
rect 5719 2097 5731 2149
rect 5783 2097 6846 2149
rect 6898 2097 6916 2149
rect 6968 2097 9821 2149
rect 9873 2097 9885 2149
rect 9937 2097 13975 2149
rect 14027 2097 14039 2149
rect 14091 2100 14361 2149
tri 14361 2100 14410 2149 nw
tri 14883 2144 14888 2149 ne
rect 14888 2100 14940 2106
rect 14091 2097 14358 2100
tri 14358 2097 14361 2100 nw
rect 2478 2017 2484 2069
rect 2536 2017 2548 2069
rect 2600 2017 2898 2069
rect 2950 2017 2962 2069
rect 3014 2017 5199 2069
rect 5505 2017 5511 2069
rect 5563 2017 5575 2069
rect 5627 2017 6078 2069
rect 6130 2017 6142 2069
rect 6194 2017 6426 2069
rect 6478 2017 6490 2069
rect 6542 2017 6993 2069
rect 7045 2017 7057 2069
rect 7109 2017 9470 2069
rect 9624 2017 9630 2069
rect 9682 2017 9694 2069
rect 9746 2017 10137 2069
rect 10189 2017 10201 2069
rect 10253 2017 13819 2069
rect 13871 2017 13883 2069
rect 13935 2017 14462 2069
rect 14514 2017 14526 2069
rect 14578 2017 14584 2069
rect 14674 2027 14735 2056
rect 2639 1702 2682 1904
rect 10464 1702 12541 1904
rect 2628 1673 2681 1674
rect 2628 1550 2682 1673
rect 3048 1668 3188 1674
rect 3100 1616 3136 1668
rect 3048 1602 3188 1616
rect 3100 1550 3136 1602
rect 2628 1544 2681 1550
rect 3048 1544 3188 1550
rect 5992 1668 6120 1674
rect 6044 1616 6068 1668
rect 5992 1602 6120 1616
rect 6044 1550 6068 1602
rect 5992 1544 6120 1550
rect 6500 1668 6628 1674
rect 6552 1616 6576 1668
rect 6500 1602 6628 1616
rect 6552 1550 6576 1602
rect 6500 1544 6628 1550
rect 10464 1544 12541 1674
rect 3813 1464 3865 1470
tri 3809 1418 3813 1422 se
rect 2753 1412 2812 1418
tri 2727 1346 2753 1372 se
rect 2805 1360 2812 1412
tri 3779 1388 3809 1418 se
rect 3809 1412 3813 1418
rect 4601 1464 4653 1470
tri 3865 1418 3869 1422 sw
tri 4597 1418 4601 1422 se
rect 3865 1412 3869 1418
rect 3809 1400 3869 1412
rect 3809 1388 3813 1400
rect 2753 1346 2812 1360
rect 2280 1342 2812 1346
rect 3865 1388 3869 1400
tri 3869 1388 3899 1418 sw
tri 4567 1388 4597 1418 se
rect 4597 1412 4601 1418
rect 7967 1464 8019 1470
tri 4653 1418 4657 1422 sw
tri 7963 1418 7967 1422 se
rect 4653 1412 4657 1418
rect 4597 1400 4657 1412
rect 4597 1388 4601 1400
rect 3813 1342 3865 1348
rect 4653 1388 4657 1400
tri 4657 1388 4687 1418 sw
rect 5654 1412 5713 1418
rect 4601 1342 4653 1348
rect 5654 1360 5661 1412
rect 5654 1342 5713 1360
rect 6907 1412 6966 1418
rect 6959 1360 6966 1412
tri 7933 1388 7963 1418 se
rect 7963 1412 7967 1418
rect 8755 1464 8807 1470
tri 8019 1418 8023 1422 sw
tri 8751 1418 8755 1422 se
rect 8019 1412 8023 1418
rect 7963 1400 8023 1412
rect 7963 1388 7967 1400
rect 2280 1290 2753 1342
rect 2805 1290 2812 1342
rect 2280 1284 2812 1290
rect 5654 1290 5661 1342
rect 5836 1303 5842 1355
rect 5894 1303 5906 1355
rect 5958 1303 5964 1355
rect 6662 1303 6668 1355
rect 6720 1303 6732 1355
rect 6784 1303 6790 1355
rect 6907 1342 6966 1360
rect 8019 1388 8023 1400
tri 8023 1388 8053 1418 sw
tri 8721 1388 8751 1418 se
rect 8751 1412 8755 1418
rect 12995 1464 13047 1470
tri 8807 1418 8811 1422 sw
tri 12991 1418 12995 1422 se
rect 8807 1412 8811 1418
rect 8751 1400 8811 1412
rect 8751 1388 8755 1400
rect 7967 1342 8019 1348
rect 8807 1388 8811 1400
tri 8811 1388 8841 1418 sw
rect 9808 1412 9867 1418
rect 8755 1342 8807 1348
rect 9808 1360 9815 1412
tri 12961 1388 12991 1418 se
rect 12991 1412 12995 1418
rect 12991 1400 13047 1412
rect 12991 1388 12995 1400
rect 9808 1342 9867 1360
rect 5654 1284 5713 1290
rect 6959 1290 6966 1342
rect 6907 1284 6966 1290
rect 9808 1290 9815 1342
rect 9990 1303 9996 1355
rect 10048 1303 10060 1355
rect 10112 1303 10118 1355
rect 12995 1342 13047 1348
rect 13962 1412 14021 1418
rect 13962 1360 13969 1412
rect 13962 1342 14021 1360
rect 9808 1284 9867 1290
rect 13962 1290 13969 1342
rect 14144 1303 14150 1355
rect 14202 1303 14214 1355
rect 14266 1303 14272 1355
rect 13962 1284 14021 1290
rect 887 1019 893 1071
rect 945 1019 957 1071
rect 1009 1019 1015 1071
tri 1015 1019 1021 1025 nw
rect 3907 1019 3913 1071
rect 3965 1019 3977 1071
rect 4029 1019 4035 1071
rect 4431 1019 4437 1071
rect 4489 1019 4501 1071
rect 4553 1019 4559 1071
rect 8061 1019 8067 1071
rect 8119 1019 8131 1071
rect 8183 1019 8189 1071
rect 8585 1019 8591 1071
rect 8643 1019 8655 1071
rect 8707 1019 8713 1071
rect 12825 1019 12831 1071
rect 12883 1019 12895 1071
rect 12947 1019 12953 1071
rect 2162 707 2205 906
rect 14618 894 14856 906
rect 14618 860 14694 894
rect 14728 860 14776 894
rect 14810 860 14856 894
rect 14618 822 14856 860
rect 14618 788 14694 822
rect 14728 788 14776 822
rect 14810 798 14856 822
tri 14856 798 14964 906 sw
rect 14810 791 15707 798
rect 14810 788 15089 791
rect 14618 739 15089 788
rect 15141 739 15707 791
rect 14618 724 15707 739
tri 14235 680 14262 707 ne
rect 2266 670 2318 676
rect 6148 670 6200 676
rect 2266 606 2318 618
rect 2266 545 2318 554
rect 2689 658 2741 664
rect 2689 594 2741 606
tri 2688 544 2689 545 se
rect 2267 543 2317 544
tri 2687 543 2688 544 se
rect 2688 543 2689 544
tri 2651 507 2687 543 se
rect 2687 542 2689 543
rect 2687 531 2741 542
rect 2687 507 2701 531
rect 2267 506 2317 507
tri 2650 506 2651 507 se
rect 2651 506 2701 507
tri 2649 505 2650 506 se
rect 2650 505 2701 506
rect 2266 453 2318 505
tri 2644 500 2649 505 se
rect 2649 500 2701 505
rect 2466 457 2512 500
tri 2635 491 2644 500 se
rect 2644 491 2701 500
tri 2701 491 2741 531 nw
rect 5725 658 5777 664
rect 5725 594 5777 606
rect 6148 606 6200 618
rect 6148 545 6200 554
rect 5725 536 5777 542
tri 5777 536 5786 545 sw
rect 6149 543 6199 544
rect 6420 670 6472 676
rect 10302 670 10354 676
rect 6420 606 6472 618
rect 6420 545 6472 554
rect 6843 658 6895 664
rect 6843 594 6895 606
tri 6842 544 6843 545 se
rect 6421 543 6471 544
tri 6841 543 6842 544 se
rect 6842 543 6843 544
rect 5725 531 5786 536
tri 5725 491 5765 531 ne
rect 5765 491 5786 531
tri 5786 491 5831 536 sw
rect 6420 507 6472 543
tri 6834 536 6841 543 se
rect 6841 542 6843 543
rect 6841 536 6895 542
tri 6805 507 6834 536 se
rect 6834 531 6895 536
rect 6834 507 6864 531
rect 6149 506 6199 507
tri 2512 457 2546 491 sw
tri 2601 457 2635 491 se
rect 2635 479 2689 491
tri 2689 479 2701 491 nw
tri 5765 479 5777 491 ne
rect 5777 479 5831 491
tri 5831 479 5843 491 sw
tri 5942 479 5954 491 se
rect 5954 479 6000 500
rect 2635 457 2681 479
tri 2681 471 2689 479 nw
tri 5777 471 5785 479 ne
rect 5785 471 5843 479
tri 5843 471 5851 479 sw
tri 5934 471 5942 479 se
rect 5942 471 6000 479
rect 2466 411 2552 457
rect 2554 456 2590 457
rect 2553 412 2591 456
rect 2554 411 2590 412
rect 2592 411 2681 457
rect 5785 457 5851 471
tri 5851 457 5865 471 sw
tri 5920 457 5934 471 se
rect 5934 457 6000 471
rect 5785 411 5874 457
rect 5876 456 5912 457
rect 5875 412 5913 456
rect 5876 411 5912 412
rect 5914 411 6000 457
rect 6148 453 6200 505
rect 6421 506 6471 507
tri 6804 506 6805 507 se
rect 6805 506 6864 507
tri 6803 505 6804 506 se
rect 6804 505 6864 506
rect 6420 453 6472 505
tri 6798 500 6803 505 se
rect 6803 500 6864 505
tri 6864 500 6895 531 nw
rect 9879 658 9931 664
rect 9879 594 9931 606
rect 10302 606 10354 618
rect 10302 545 10354 554
rect 9879 536 9931 542
tri 9931 536 9940 545 sw
rect 10303 543 10353 544
rect 14033 658 14085 664
rect 14262 656 14308 708
rect 14456 707 14508 714
rect 14618 707 15089 724
tri 14308 682 14333 707 nw
tri 14422 682 14447 707 ne
rect 14447 682 14511 707
tri 14511 682 14536 707 nw
tri 14775 682 14800 707 ne
rect 14800 682 15089 707
tri 14447 680 14449 682 ne
rect 14449 680 14509 682
tri 14509 680 14511 682 nw
tri 14800 680 14802 682 ne
rect 14802 680 15089 682
tri 14449 676 14453 680 ne
rect 14453 676 14508 680
tri 14508 679 14509 680 nw
tri 14802 679 14803 680 ne
rect 14803 679 15089 680
tri 14803 676 14806 679 ne
rect 14806 676 15089 679
tri 14453 673 14456 676 ne
rect 14263 654 14307 655
rect 14456 662 14508 676
tri 14806 662 14820 676 ne
rect 14820 672 15089 676
rect 15141 672 15707 724
rect 14820 662 15707 672
tri 14820 661 14821 662 ne
rect 14821 661 15707 662
rect 14457 660 14507 661
tri 14821 660 14822 661 ne
rect 14822 660 15707 661
rect 14456 624 14508 660
tri 14822 624 14858 660 ne
rect 14858 658 15707 660
rect 14858 624 15089 658
rect 14457 623 14507 624
rect 14033 594 14085 606
rect 14263 617 14307 618
rect 14262 564 14308 616
rect 14456 570 14508 622
rect 14731 618 14783 624
tri 14858 600 14882 624 ne
rect 14882 606 15089 624
rect 15141 606 15707 658
rect 14882 600 15707 606
rect 14731 554 14783 566
rect 14033 536 14085 542
tri 14085 536 14094 545 sw
rect 9879 531 9940 536
tri 9879 500 9910 531 ne
rect 9910 500 9940 531
tri 9940 500 9976 536 sw
rect 14033 531 14094 536
tri 14033 507 14057 531 ne
rect 14057 507 14094 531
rect 10303 506 10353 507
tri 14057 506 14058 507 ne
rect 14058 506 14094 507
tri 14058 505 14059 506 ne
rect 14059 505 14094 506
rect 6620 479 6666 500
tri 6789 491 6798 500 se
rect 6798 491 6855 500
tri 6855 491 6864 500 nw
tri 9910 491 9919 500 ne
rect 9919 491 9976 500
tri 9976 491 9985 500 sw
tri 6666 479 6678 491 sw
tri 6777 479 6789 491 se
rect 6789 479 6843 491
tri 6843 479 6855 491 nw
tri 9919 479 9931 491 ne
rect 9931 479 9985 491
rect 6620 471 6678 479
tri 6678 471 6686 479 sw
tri 6769 471 6777 479 se
rect 6777 471 6835 479
tri 6835 471 6843 479 nw
tri 9931 471 9939 479 ne
rect 6620 457 6686 471
tri 6686 457 6700 471 sw
tri 6755 457 6769 471 se
rect 6769 457 6835 471
rect 2266 358 2318 410
rect 2466 398 2533 411
tri 2533 398 2546 411 nw
tri 5920 398 5933 411 ne
rect 5933 398 6000 411
rect 6620 411 6706 457
rect 6707 412 6708 456
rect 6744 412 6745 456
rect 6746 411 6835 457
rect 9939 457 9985 479
tri 9985 457 10019 491 sw
tri 10074 457 10108 491 se
rect 10108 457 10154 500
rect 9939 411 10028 457
rect 10030 456 10066 457
rect 10029 412 10067 456
rect 10030 411 10066 412
rect 10068 411 10154 457
rect 10302 453 10354 505
tri 14059 500 14064 505 ne
rect 14064 500 14094 505
tri 14094 500 14130 536 sw
tri 14064 491 14073 500 ne
rect 14073 491 14130 500
tri 14130 491 14139 500 sw
tri 14073 479 14085 491 ne
rect 14085 479 14139 491
tri 14085 471 14093 479 ne
rect 2466 372 2512 398
tri 2512 377 2533 398 nw
rect 2467 370 2511 371
rect 2267 356 2317 357
rect 2266 320 2318 356
rect 2467 333 2511 334
tri 2462 320 2466 324 se
rect 2466 320 2512 332
rect 2267 319 2317 320
tri 2461 319 2462 320 se
rect 2462 319 2512 320
tri 2460 318 2461 319 se
rect 2461 318 2512 319
rect 2266 290 2318 318
tri 2458 316 2460 318 se
rect 2460 316 2512 318
tri 2318 290 2344 316 sw
tri 2432 290 2458 316 se
rect 2458 290 2512 316
tri 2512 290 2546 324 sw
tri 4176 290 4210 324 se
rect 4210 290 4256 398
tri 5933 377 5954 398 ne
rect 5954 372 6000 398
rect 5955 370 5999 371
rect 6148 358 6200 410
rect 6149 356 6199 357
rect 6420 358 6472 410
rect 6421 356 6471 357
rect 6620 372 6666 411
tri 6666 377 6700 411 nw
tri 10074 398 10087 411 ne
rect 10087 398 10154 411
rect 14093 411 14139 479
tri 14139 411 14169 441 sw
tri 14232 411 14262 441 se
rect 14262 411 14308 500
rect 14456 469 14508 521
rect 14457 467 14507 468
rect 14910 548 14962 600
rect 14911 546 14961 547
rect 15452 520 15523 558
rect 15842 550 15873 608
rect 14731 496 14783 502
rect 6621 370 6665 371
rect 5955 333 5999 334
tri 5920 290 5954 324 se
rect 5954 316 6000 332
tri 6000 316 6008 324 sw
rect 6148 320 6200 356
rect 6620 334 6666 370
rect 6621 333 6665 334
tri 6616 320 6620 324 se
rect 6620 320 6666 332
rect 6149 319 6199 320
rect 5954 290 6008 316
tri 6008 290 6034 316 sw
tri 6122 290 6148 316 se
rect 6148 290 6200 318
rect 6421 319 6471 320
tri 6615 319 6616 320 se
rect 6616 319 6666 320
tri 6614 318 6615 319 se
rect 6615 318 6666 319
tri 6200 290 6226 316 sw
tri 6394 290 6420 316 se
rect 6420 290 6472 318
tri 6612 316 6614 318 se
rect 6614 316 6666 318
tri 6472 290 6498 316 sw
tri 6586 290 6612 316 se
rect 6612 290 6666 316
tri 6666 290 6700 324 sw
rect 8364 290 8410 398
tri 10087 377 10108 398 ne
rect 10108 372 10154 398
rect 10109 370 10153 371
rect 10302 358 10354 410
rect 14093 407 14169 411
tri 14169 407 14173 411 sw
tri 14228 407 14232 411 se
rect 14232 407 14308 411
rect 14093 361 14182 407
rect 14184 406 14220 407
rect 14183 362 14221 406
rect 14184 361 14220 362
rect 14222 361 14308 407
rect 14457 430 14507 431
rect 14456 413 14508 429
rect 14641 413 14693 419
tri 14638 370 14641 373 se
rect 10303 356 10353 357
rect 10109 333 10153 334
tri 8410 290 8444 324 sw
tri 10074 290 10108 324 se
rect 10108 290 10154 332
tri 10154 290 10188 324 sw
rect 10302 320 10354 356
rect 10303 319 10353 320
tri 10276 290 10302 316 se
rect 10302 290 10354 318
rect 14456 349 14508 361
tri 14508 343 14535 370 sw
tri 14611 343 14638 370 se
rect 14638 361 14641 370
rect 14638 349 14693 361
rect 14638 343 14641 349
rect 14508 297 14641 343
rect 14456 291 14693 297
rect 2266 238 4256 290
rect 4346 238 7881 290
rect 8364 238 10354 290
rect 2162 9 2205 210
rect 10464 9 12534 210
rect 14731 134 14777 496
tri 14777 490 14783 496 nw
rect 14911 509 14961 510
rect 14910 467 14962 508
rect 14910 403 14962 415
rect 14734 12 14774 64
rect 14910 -26 14962 351
rect 15081 102 15133 104
rect 15253 -33 15305 -24
<< rmetal1 >>
rect 2266 544 2318 545
rect 2266 543 2267 544
rect 2317 543 2318 544
rect 2266 506 2267 507
rect 2317 506 2318 507
rect 2266 505 2318 506
rect 6148 544 6200 545
rect 6148 543 6149 544
rect 6199 543 6200 544
rect 6420 544 6472 545
rect 6420 543 6421 544
rect 6471 543 6472 544
rect 6148 506 6149 507
rect 6199 506 6200 507
rect 6148 505 6200 506
rect 2552 456 2554 457
rect 2590 456 2592 457
rect 2552 412 2553 456
rect 2591 412 2592 456
rect 2552 411 2554 412
rect 2590 411 2592 412
rect 5874 456 5876 457
rect 5912 456 5914 457
rect 5874 412 5875 456
rect 5913 412 5914 456
rect 5874 411 5876 412
rect 5912 411 5914 412
rect 6420 506 6421 507
rect 6471 506 6472 507
rect 6420 505 6472 506
rect 10302 544 10354 545
rect 10302 543 10303 544
rect 10353 543 10354 544
rect 14262 655 14308 656
rect 14262 654 14263 655
rect 14307 654 14308 655
rect 14456 661 14508 662
rect 14456 660 14457 661
rect 14507 660 14508 661
rect 14456 623 14457 624
rect 14507 623 14508 624
rect 14456 622 14508 623
rect 14262 617 14263 618
rect 14307 617 14308 618
rect 14262 616 14308 617
rect 10302 506 10303 507
rect 10353 506 10354 507
rect 10302 505 10354 506
rect 6706 456 6708 457
rect 6706 412 6707 456
rect 6706 411 6708 412
rect 6744 456 6746 457
rect 6745 412 6746 456
rect 6744 411 6746 412
rect 10028 456 10030 457
rect 10066 456 10068 457
rect 10028 412 10029 456
rect 10067 412 10068 456
rect 10028 411 10030 412
rect 10066 411 10068 412
rect 2466 371 2512 372
rect 2466 370 2467 371
rect 2511 370 2512 371
rect 2266 357 2318 358
rect 2266 356 2267 357
rect 2317 356 2318 357
rect 2466 333 2467 334
rect 2511 333 2512 334
rect 2466 332 2512 333
rect 2266 319 2267 320
rect 2317 319 2318 320
rect 2266 318 2318 319
rect 5954 371 6000 372
rect 5954 370 5955 371
rect 5999 370 6000 371
rect 6148 357 6200 358
rect 6148 356 6149 357
rect 6199 356 6200 357
rect 6420 357 6472 358
rect 6420 356 6421 357
rect 6471 356 6472 357
rect 14456 468 14508 469
rect 14456 467 14457 468
rect 14507 467 14508 468
rect 14910 547 14962 548
rect 14910 546 14911 547
rect 14961 546 14962 547
rect 6620 371 6666 372
rect 6620 370 6621 371
rect 6665 370 6666 371
rect 5954 333 5955 334
rect 5999 333 6000 334
rect 5954 332 6000 333
rect 6620 333 6621 334
rect 6665 333 6666 334
rect 6620 332 6666 333
rect 6148 319 6149 320
rect 6199 319 6200 320
rect 6148 318 6200 319
rect 6420 319 6421 320
rect 6471 319 6472 320
rect 6420 318 6472 319
rect 10108 371 10154 372
rect 10108 370 10109 371
rect 10153 370 10154 371
rect 14182 406 14184 407
rect 14220 406 14222 407
rect 14182 362 14183 406
rect 14221 362 14222 406
rect 14182 361 14184 362
rect 14220 361 14222 362
rect 14456 430 14457 431
rect 14507 430 14508 431
rect 14456 429 14508 430
rect 10302 357 10354 358
rect 10302 356 10303 357
rect 10353 356 10354 357
rect 10108 333 10109 334
rect 10153 333 10154 334
rect 10108 332 10154 333
rect 10302 319 10303 320
rect 10353 319 10354 320
rect 10302 318 10354 319
rect 14910 509 14911 510
rect 14961 509 14962 510
rect 14910 508 14962 509
<< via1 >>
rect 3049 3008 3101 3060
rect 3137 3008 3189 3060
rect 3049 2926 3101 2978
rect 3137 2926 3189 2978
rect 3049 2843 3101 2895
rect 3137 2843 3189 2895
rect 3049 2760 3101 2812
rect 3137 2760 3189 2812
rect 14888 2170 14940 2222
rect 889 2097 941 2149
rect 953 2097 1005 2149
rect 2759 2097 2811 2149
rect 2823 2097 2875 2149
rect 5667 2097 5719 2149
rect 5731 2097 5783 2149
rect 6846 2097 6898 2149
rect 6916 2097 6968 2149
rect 9821 2097 9873 2149
rect 9885 2097 9937 2149
rect 13975 2097 14027 2149
rect 14039 2097 14091 2149
rect 14888 2106 14940 2158
rect 2484 2017 2536 2069
rect 2548 2017 2600 2069
rect 2898 2017 2950 2069
rect 2962 2017 3014 2069
rect 5511 2017 5563 2069
rect 5575 2017 5627 2069
rect 6078 2017 6130 2069
rect 6142 2017 6194 2069
rect 6426 2017 6478 2069
rect 6490 2017 6542 2069
rect 6993 2017 7045 2069
rect 7057 2017 7109 2069
rect 9630 2017 9682 2069
rect 9694 2017 9746 2069
rect 10137 2017 10189 2069
rect 10201 2017 10253 2069
rect 13819 2017 13871 2069
rect 13883 2017 13935 2069
rect 14462 2017 14514 2069
rect 14526 2017 14578 2069
rect 3048 1616 3100 1668
rect 3136 1616 3188 1668
rect 3048 1550 3100 1602
rect 3136 1550 3188 1602
rect 5992 1616 6044 1668
rect 6068 1616 6120 1668
rect 5992 1550 6044 1602
rect 6068 1550 6120 1602
rect 6500 1616 6552 1668
rect 6576 1616 6628 1668
rect 6500 1550 6552 1602
rect 6576 1550 6628 1602
rect 2753 1360 2805 1412
rect 3813 1412 3865 1464
rect 3813 1348 3865 1400
rect 4601 1412 4653 1464
rect 4601 1348 4653 1400
rect 5661 1360 5713 1412
rect 6907 1360 6959 1412
rect 7967 1412 8019 1464
rect 2753 1290 2805 1342
rect 5661 1290 5713 1342
rect 5842 1303 5894 1355
rect 5906 1303 5958 1355
rect 6668 1303 6720 1355
rect 6732 1303 6784 1355
rect 7967 1348 8019 1400
rect 8755 1412 8807 1464
rect 8755 1348 8807 1400
rect 9815 1360 9867 1412
rect 12995 1412 13047 1464
rect 6907 1290 6959 1342
rect 9815 1290 9867 1342
rect 9996 1303 10048 1355
rect 10060 1303 10112 1355
rect 12995 1348 13047 1400
rect 13969 1360 14021 1412
rect 13969 1290 14021 1342
rect 14150 1303 14202 1355
rect 14214 1303 14266 1355
rect 893 1019 945 1071
rect 957 1019 1009 1071
rect 3913 1019 3965 1071
rect 3977 1019 4029 1071
rect 4437 1019 4489 1071
rect 4501 1019 4553 1071
rect 8067 1019 8119 1071
rect 8131 1019 8183 1071
rect 8591 1019 8643 1071
rect 8655 1019 8707 1071
rect 12831 1019 12883 1071
rect 12895 1019 12947 1071
rect 15089 739 15141 791
rect 2266 618 2318 670
rect 2266 554 2318 606
rect 2689 606 2741 658
rect 2689 542 2741 594
rect 5725 606 5777 658
rect 5725 542 5777 594
rect 6148 618 6200 670
rect 6148 554 6200 606
rect 6420 618 6472 670
rect 6420 554 6472 606
rect 6843 606 6895 658
rect 6843 542 6895 594
rect 9879 606 9931 658
rect 9879 542 9931 594
rect 10302 618 10354 670
rect 10302 554 10354 606
rect 14033 606 14085 658
rect 15089 672 15141 724
rect 14033 542 14085 594
rect 14731 566 14783 618
rect 15089 606 15141 658
rect 14731 502 14783 554
rect 14456 361 14508 413
rect 14456 297 14508 349
rect 14641 361 14693 413
rect 14641 297 14693 349
rect 14910 415 14962 467
rect 14910 351 14962 403
<< metal2 >>
rect 3048 3060 3189 3066
rect 3048 3008 3049 3060
rect 3101 3008 3137 3060
rect 3048 2978 3189 3008
rect 3048 2926 3049 2978
rect 3101 2926 3137 2978
rect 3048 2895 3189 2926
rect 3048 2843 3049 2895
rect 3101 2843 3137 2895
rect 3048 2812 3189 2843
rect 3048 2760 3049 2812
rect 3101 2760 3137 2812
rect 883 2097 889 2149
rect 941 2097 953 2149
rect 1005 2097 1011 2149
tri 883 2069 911 2097 ne
rect 911 2069 983 2097
tri 983 2069 1011 2097 nw
rect 2753 2097 2759 2149
rect 2811 2097 2823 2149
rect 2875 2097 2881 2149
rect 2753 2069 2811 2097
tri 2811 2069 2839 2097 nw
tri 911 2059 921 2069 ne
tri 887 1071 921 1105 se
rect 921 1071 973 2069
tri 973 2059 983 2069 nw
rect 2478 2017 2484 2069
rect 2536 2017 2548 2069
rect 2600 2017 2606 2069
tri 2474 1284 2478 1288 se
rect 2478 1284 2530 2017
tri 2530 1983 2564 2017 nw
rect 2753 1412 2805 2069
tri 2805 2063 2811 2069 nw
rect 2892 2017 2898 2069
rect 2950 2017 2962 2069
rect 3014 2017 3020 2069
rect 2753 1342 2805 1360
rect 2753 1284 2805 1290
tri 2833 1813 2892 1872 se
rect 2892 1850 2944 2017
tri 2944 1983 2978 2017 nw
rect 2892 1813 2907 1850
tri 2907 1813 2944 1850 nw
tri 2443 1253 2474 1284 se
rect 2474 1266 2530 1284
rect 2474 1253 2517 1266
tri 2517 1253 2530 1266 nw
rect 2443 1188 2498 1253
tri 2498 1234 2517 1253 nw
tri 973 1071 1015 1113 sw
rect 887 1019 893 1071
rect 945 1019 957 1071
rect 1009 1019 1015 1071
rect 2443 1079 2484 1188
tri 2484 1174 2498 1188 nw
tri 2484 1079 2498 1093 sw
tri 2441 889 2443 891 se
rect 2443 889 2498 1079
tri 2799 889 2833 923 se
rect 2833 889 2885 1813
tri 2885 1791 2907 1813 nw
rect 3048 1668 3189 2760
rect 14888 2222 14940 2228
rect 14888 2158 14940 2170
rect 5661 2097 5667 2149
rect 5719 2097 5731 2149
rect 5783 2097 5789 2149
rect 6840 2097 6846 2149
rect 6898 2097 6916 2149
rect 6968 2097 6974 2149
rect 5661 2069 5761 2097
tri 5761 2069 5789 2097 nw
tri 6867 2069 6895 2097 ne
rect 6895 2069 6959 2097
tri 6959 2082 6974 2097 nw
rect 9815 2097 9821 2149
rect 9873 2097 9885 2149
rect 9937 2097 9943 2149
rect 9815 2082 9928 2097
tri 9928 2082 9943 2097 nw
rect 13969 2097 13975 2149
rect 14027 2097 14039 2149
rect 14091 2097 14097 2149
rect 9815 2069 9915 2082
tri 9915 2069 9928 2082 nw
rect 13969 2069 14069 2097
tri 14069 2069 14097 2097 nw
rect 5505 2017 5511 2069
rect 5563 2017 5575 2069
rect 5627 2017 5633 2069
tri 5547 1983 5581 2017 ne
rect 3100 1616 3136 1668
rect 3188 1616 3189 1668
rect 3048 1602 3189 1616
rect 3100 1550 3136 1602
rect 3188 1550 3189 1602
rect 3048 1544 3189 1550
tri 2369 817 2441 889 se
rect 2441 872 2498 889
rect 2441 817 2443 872
tri 2443 817 2498 872 nw
tri 2689 847 2731 889 se
rect 2731 862 2885 889
rect 2731 847 2870 862
tri 2870 847 2885 862 nw
rect 3813 1464 3865 1470
rect 3813 1400 3865 1412
rect 2689 837 2860 847
tri 2860 837 2870 847 nw
tri 2343 791 2369 817 se
rect 2369 791 2417 817
tri 2417 791 2443 817 nw
tri 2295 743 2343 791 se
rect 2343 743 2369 791
tri 2369 743 2417 791 nw
tri 2291 739 2295 743 se
rect 2295 739 2365 743
tri 2365 739 2369 743 nw
tri 2276 724 2291 739 se
rect 2291 724 2350 739
tri 2350 724 2365 739 nw
tri 2266 714 2276 724 se
rect 2276 714 2340 724
tri 2340 714 2350 724 nw
rect 2266 670 2318 714
tri 2318 692 2340 714 nw
rect 2266 606 2318 618
rect 2266 548 2318 554
rect 2689 658 2741 837
tri 2741 803 2775 837 nw
rect 2689 594 2741 606
rect 2689 536 2741 542
rect 3813 9 3865 1348
rect 4601 1464 4653 1470
rect 4601 1400 4653 1412
rect 3907 1019 3913 1071
rect 3965 1019 3977 1071
rect 4029 1019 4035 1071
rect 4431 1019 4437 1071
rect 4489 1019 4501 1071
rect 4553 1019 4559 1071
rect 3907 9 3959 1019
tri 3959 964 4014 1019 nw
tri 4470 982 4507 1019 ne
rect 4507 9 4559 1019
rect 4601 9 4653 1348
rect 5581 889 5633 2017
rect 5661 1412 5713 2069
tri 5713 2021 5761 2069 nw
rect 6072 2017 6078 2069
rect 6130 2017 6142 2069
rect 6194 2017 6200 2069
tri 6114 1998 6133 2017 ne
rect 6133 1998 6200 2017
tri 5864 1365 5902 1403 se
rect 5902 1365 5954 1998
tri 6133 1983 6148 1998 ne
rect 5992 1668 6120 1674
rect 6044 1616 6068 1668
rect 5992 1602 6120 1616
rect 6044 1550 6068 1602
rect 5992 1514 6120 1550
tri 5859 1360 5864 1365 se
rect 5864 1360 5954 1365
tri 5954 1360 5959 1365 sw
rect 5661 1342 5713 1360
tri 5854 1355 5859 1360 se
rect 5859 1355 5959 1360
tri 5959 1355 5964 1360 sw
rect 5836 1303 5842 1355
rect 5894 1303 5906 1355
rect 5958 1303 5964 1355
rect 5661 1284 5713 1290
tri 5633 889 5667 923 sw
rect 5581 862 5735 889
tri 5581 847 5596 862 ne
rect 5596 847 5735 862
tri 5735 847 5777 889 sw
tri 5596 837 5606 847 ne
rect 5606 837 5777 847
tri 5691 803 5725 837 ne
rect 5725 658 5777 837
rect 5725 594 5777 606
rect 6148 670 6200 1998
rect 6148 606 6200 618
rect 6148 548 6200 554
rect 6420 2017 6426 2069
rect 6478 2017 6490 2069
rect 6542 2017 6548 2069
tri 6895 2057 6907 2069 ne
rect 6420 1998 6487 2017
tri 6487 1998 6506 2017 nw
rect 6420 670 6472 1998
tri 6472 1983 6487 1998 nw
rect 6500 1668 6628 1674
rect 6552 1616 6576 1668
rect 6500 1602 6628 1616
rect 6552 1550 6576 1602
rect 6500 1514 6628 1550
tri 6673 1360 6702 1389 se
rect 6702 1360 6754 1998
rect 6907 1412 6959 2069
tri 6754 1360 6783 1389 sw
tri 6668 1355 6673 1360 se
rect 6673 1355 6783 1360
tri 6783 1355 6788 1360 sw
rect 6662 1303 6668 1355
rect 6720 1303 6732 1355
rect 6784 1303 6790 1355
rect 6907 1342 6959 1360
rect 6907 1284 6959 1290
rect 6987 2017 6993 2069
rect 7045 2017 7057 2069
rect 7109 2017 7115 2069
rect 9624 2017 9630 2069
rect 9682 2017 9694 2069
rect 9746 2017 9752 2069
tri 6953 889 6987 923 se
rect 6987 889 7039 2017
tri 7039 1983 7073 2017 nw
tri 9642 1993 9666 2017 ne
rect 9666 1993 9728 2017
tri 9728 1993 9752 2017 nw
tri 9666 1983 9676 1993 ne
rect 9676 1850 9728 1993
tri 9676 1813 9713 1850 ne
rect 9713 1813 9728 1850
tri 9728 1813 9787 1872 sw
tri 9713 1798 9728 1813 ne
rect 9728 1798 9787 1813
tri 9728 1791 9735 1798 ne
rect 6420 606 6472 618
rect 6420 548 6472 554
tri 6843 847 6885 889 se
rect 6885 862 7039 889
rect 6885 847 7024 862
tri 7024 847 7039 862 nw
rect 7967 1464 8019 1470
rect 7967 1400 8019 1412
rect 6843 837 7014 847
tri 7014 837 7024 847 nw
rect 6843 658 6895 837
tri 6895 803 6929 837 nw
rect 6843 594 6895 606
rect 5725 536 5777 542
rect 6843 536 6895 542
rect 7967 9 8019 1348
rect 8755 1464 8807 1470
rect 8755 1400 8807 1412
rect 8061 1019 8067 1071
rect 8119 1019 8131 1071
rect 8183 1019 8189 1071
rect 8585 1019 8591 1071
rect 8643 1019 8655 1071
rect 8707 1019 8713 1071
rect 8061 9 8113 1019
tri 8113 965 8167 1019 nw
tri 8603 965 8657 1019 ne
rect 8657 965 8713 1019
tri 8657 961 8661 965 ne
rect 8661 9 8713 965
rect 8755 9 8807 1348
rect 9735 889 9787 1798
rect 9815 1412 9867 2069
tri 9867 2021 9915 2069 nw
rect 10131 2017 10137 2069
rect 10189 2017 10201 2069
rect 10253 2017 10259 2069
rect 13813 2017 13819 2069
rect 13871 2017 13883 2069
rect 13935 2017 13941 2069
tri 10131 2010 10138 2017 ne
rect 10138 2010 10259 2017
tri 10138 1998 10150 2010 ne
rect 10150 1998 10232 2010
rect 9815 1342 9867 1360
tri 9997 1355 10031 1389 se
rect 10031 1355 10083 1998
tri 10150 1983 10165 1998 ne
rect 10165 1983 10232 1998
tri 10232 1983 10259 2010 nw
tri 13855 1983 13889 2017 ne
tri 10165 1968 10180 1983 ne
rect 10180 1703 10232 1983
tri 10180 1677 10206 1703 ne
rect 10206 1677 10232 1703
tri 10232 1677 10280 1725 sw
tri 10206 1651 10232 1677 ne
rect 10232 1651 10280 1677
tri 10232 1603 10280 1651 ne
tri 10280 1603 10354 1677 sw
tri 10280 1581 10302 1603 ne
tri 10083 1355 10117 1389 sw
rect 9990 1303 9996 1355
rect 10048 1303 10060 1355
rect 10112 1303 10118 1355
rect 9815 1284 9867 1290
tri 9787 889 9821 923 sw
rect 9735 862 9889 889
tri 9735 847 9750 862 ne
rect 9750 847 9889 862
tri 9889 847 9931 889 sw
tri 9750 837 9760 847 ne
rect 9760 837 9931 847
tri 9845 803 9879 837 ne
rect 9879 658 9931 837
rect 9879 594 9931 606
rect 10302 670 10354 1603
rect 12995 1464 13047 1470
rect 12995 1400 13047 1412
rect 12825 1019 12831 1071
rect 12883 1019 12895 1071
rect 12947 1019 12953 1071
tri 12837 955 12901 1019 ne
rect 10302 606 10354 618
rect 10302 548 10354 554
rect 9879 536 9931 542
rect 12901 9 12953 1019
rect 12995 9 13047 1348
rect 13889 889 13941 2017
rect 13969 2063 14063 2069
tri 14063 2063 14069 2069 nw
rect 13969 2022 14022 2063
tri 14022 2022 14063 2063 nw
rect 13969 1412 14021 2022
tri 14021 2021 14022 2022 nw
rect 14456 2017 14462 2069
rect 14514 2017 14526 2069
rect 14578 2017 14584 2069
tri 14181 1391 14184 1394 se
rect 14184 1391 14236 1998
rect 13969 1342 14021 1360
tri 14145 1355 14181 1391 se
rect 14181 1355 14236 1391
tri 14236 1355 14272 1391 sw
rect 14144 1303 14150 1355
rect 14202 1303 14214 1355
rect 14266 1303 14272 1355
rect 13969 1284 14021 1290
tri 13941 889 13975 923 sw
rect 13889 862 14043 889
tri 13889 847 13904 862 ne
rect 13904 847 14043 862
tri 14043 847 14085 889 sw
tri 13904 837 13914 847 ne
rect 13914 837 14085 847
tri 13999 803 14033 837 ne
rect 14033 658 14085 837
rect 14033 594 14085 606
rect 14033 536 14085 542
rect 14456 413 14508 2017
tri 14508 1983 14542 2017 nw
tri 14883 791 14888 796 se
rect 14888 791 14940 2106
tri 14831 739 14883 791 se
rect 14883 774 14940 791
rect 14883 739 14905 774
tri 14905 739 14940 774 nw
rect 15089 791 15141 797
tri 14816 724 14831 739 se
rect 14831 724 14890 739
tri 14890 724 14905 739 nw
rect 15089 724 15141 739
tri 14814 722 14816 724 se
rect 14816 722 14888 724
tri 14888 722 14890 724 nw
tri 14764 672 14814 722 se
rect 14814 672 14838 722
tri 14838 672 14888 722 nw
tri 14750 658 14764 672 se
rect 14764 658 14824 672
tri 14824 658 14838 672 nw
rect 15089 658 15141 672
tri 14740 648 14750 658 se
rect 14750 648 14814 658
tri 14814 648 14824 658 nw
tri 14731 639 14740 648 se
rect 14740 639 14805 648
tri 14805 639 14814 648 nw
rect 14731 624 14790 639
tri 14790 624 14805 639 nw
rect 14731 618 14783 624
tri 14783 617 14790 624 nw
rect 14731 554 14783 566
rect 14731 496 14783 502
tri 14904 467 14910 473 se
rect 14910 467 14962 473
tri 14898 461 14904 467 se
rect 14904 461 14910 467
rect 14456 349 14508 361
rect 14456 291 14508 297
rect 14641 413 14798 461
rect 14800 460 14836 461
rect 14693 409 14798 413
rect 14799 410 14837 460
rect 14838 415 14910 461
rect 14800 409 14836 410
rect 14838 409 14962 415
rect 14693 403 14735 409
tri 14735 403 14741 409 nw
tri 14880 403 14886 409 ne
rect 14886 403 14962 409
tri 14693 361 14735 403 nw
tri 14886 379 14910 403 ne
rect 14641 349 14693 361
rect 14910 345 14962 351
rect 15089 367 15141 606
rect 15090 365 15140 366
rect 14641 229 14693 297
rect 15089 329 15141 365
rect 15090 328 15140 329
tri 14693 229 14695 231 sw
rect 14641 209 14695 229
tri 14641 155 14695 209 ne
tri 14695 155 14769 229 sw
tri 15057 155 15089 187 se
rect 15089 155 15141 327
tri 14695 103 14747 155 ne
rect 14747 103 14989 155
rect 14990 104 14991 154
rect 15027 104 15028 154
rect 15029 141 15141 155
rect 15029 103 15133 141
tri 15133 133 15141 141 nw
tri 15056 78 15081 103 ne
rect 15081 102 15133 103
rect 14820 9 14949 54
tri 14949 9 14994 54 sw
rect 14820 2 14994 9
tri 14994 2 15001 9 sw
tri 14927 -72 15001 2 ne
tri 15001 -17 15020 2 sw
rect 15001 -39 15020 -17
tri 15020 -39 15042 -17 sw
tri 15231 -39 15253 -17 se
rect 15253 -39 15305 -24
rect 15001 -49 15042 -39
tri 15042 -49 15052 -39 sw
tri 15221 -49 15231 -39 se
rect 15231 -49 15295 -39
tri 15295 -49 15305 -39 nw
rect 15001 -71 15052 -49
tri 15052 -71 15074 -49 sw
tri 15199 -71 15221 -49 se
rect 15221 -71 15272 -49
rect 15001 -72 15272 -71
tri 15272 -72 15295 -49 nw
tri 15001 -123 15052 -72 ne
rect 15052 -123 15221 -72
tri 15221 -123 15272 -72 nw
<< rmetal2 >>
rect 14798 460 14800 461
rect 14836 460 14838 461
rect 14798 410 14799 460
rect 14837 410 14838 460
rect 14798 409 14800 410
rect 14836 409 14838 410
rect 15089 366 15141 367
rect 15089 365 15090 366
rect 15140 365 15141 366
rect 15089 328 15090 329
rect 15140 328 15141 329
rect 15089 327 15141 328
rect 14989 154 14991 155
rect 14989 104 14990 154
rect 14989 103 14991 104
rect 15027 154 15029 155
rect 15028 104 15029 154
rect 15027 103 15029 104
use sky130_fd_io__com_ctl_ls_1v2  sky130_fd_io__com_ctl_ls_1v2_0
timestamp 1701704242
transform 1 0 12541 0 -1 2028
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_en_1_v2  sky130_fd_io__com_ctl_ls_en_1_v2_0
timestamp 1701704242
transform -1 0 4233 0 -1 2028
box -71 -1302 2077 2019
use sky130_fd_io__com_ctl_ls_v2  sky130_fd_io__com_ctl_ls_v2_0
timestamp 1701704242
transform 1 0 8387 0 -1 2028
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_v2  sky130_fd_io__com_ctl_ls_v2_1
timestamp 1701704242
transform -1 0 8387 0 -1 2028
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_v2  sky130_fd_io__com_ctl_ls_v2_2
timestamp 1701704242
transform 1 0 4233 0 -1 2028
box -71 10 2077 2019
use sky130_fd_io__com_ctl_lsv2  sky130_fd_io__com_ctl_lsv2_0
timestamp 1701704242
transform -1 0 20585 0 -1 2028
box 4577 -1281 6166 3353
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_0
timestamp 1701704242
transform 0 -1 14308 -1 0 708
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_1
timestamp 1701704242
transform 1 0 6654 0 1 411
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_2
timestamp 1701704242
transform 0 1 10108 1 0 280
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_3
timestamp 1701704242
transform 0 1 5954 1 0 280
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_4
timestamp 1701704242
transform 0 -1 2512 1 0 280
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1701704242
transform 0 -1 14508 1 0 377
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1701704242
transform 0 1 14910 -1 0 600
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_2
timestamp 1701704242
transform 0 1 6420 -1 0 410
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_3
timestamp 1701704242
transform 0 -1 10354 -1 0 597
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_4
timestamp 1701704242
transform 0 -1 6200 -1 0 597
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_5
timestamp 1701704242
transform 0 1 2266 -1 0 597
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1701704242
transform 1 0 14130 0 1 361
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_1
timestamp 1701704242
transform 0 -1 6666 1 0 280
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_2
timestamp 1701704242
transform -1 0 10120 0 1 411
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_3
timestamp 1701704242
transform -1 0 5966 0 1 411
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_4
timestamp 1701704242
transform 1 0 2500 0 1 411
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1701704242
transform 0 1 6420 -1 0 597
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1701704242
transform 0 -1 10354 -1 0 410
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_2
timestamp 1701704242
transform 0 -1 6200 -1 0 410
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_3
timestamp 1701704242
transform 0 1 2266 -1 0 410
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_4
timestamp 1701704242
transform 0 -1 14508 -1 0 714
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808439  sky130_fd_io__tk_em2o_cdns_55959141808439_0
timestamp 1701704242
transform 1 0 14937 0 -1 155
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808438  sky130_fd_io__tk_em2s_cdns_55959141808438_0
timestamp 1701704242
transform -1 0 14890 0 -1 461
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808438  sky130_fd_io__tk_em2s_cdns_55959141808438_1
timestamp 1701704242
transform 0 -1 15141 1 0 275
box 0 0 1 1
<< labels >>
flabel metal2 s 12995 9 13047 61 3 FreeSans 520 90 0 0 VTRIP_SEL_H
port 2 nsew
flabel metal2 s 14184 1946 14236 1998 3 FreeSans 520 270 0 0 VTRIP_SEL
port 3 nsew
flabel metal2 s 12901 9 12953 61 3 FreeSans 520 90 0 0 VTRIP_SEL_H_N
port 4 nsew
flabel metal2 s 6702 1946 6754 1998 3 FreeSans 520 270 0 0 INP_DIS
port 5 nsew
flabel metal2 s 7967 9 8019 61 3 FreeSans 520 90 0 0 INP_DIS_H
port 6 nsew
flabel metal2 s 8061 9 8113 61 3 FreeSans 520 90 0 0 INP_DIS_H_N
port 7 nsew
flabel metal2 s 5902 1946 5954 1998 3 FreeSans 520 270 0 0 DM[0]
port 8 nsew
flabel metal2 s 4601 9 4653 61 3 FreeSans 520 90 0 0 DM_H[0]
port 9 nsew
flabel metal2 s 4507 9 4559 61 3 FreeSans 520 90 0 0 DM_H_N[0]
port 10 nsew
flabel metal2 s 3813 9 3865 61 3 FreeSans 520 90 0 0 DM_H[1]
port 11 nsew
flabel metal2 s 3907 9 3959 61 3 FreeSans 520 90 0 0 DM_H_N[1]
port 12 nsew
flabel metal2 s 10031 1946 10083 1998 3 FreeSans 520 270 0 0 DM[2]
port 13 nsew
flabel metal2 s 8755 9 8807 61 3 FreeSans 520 90 0 0 DM_H[2]
port 14 nsew
flabel metal2 s 8661 9 8713 61 3 FreeSans 520 90 0 0 DM_H_N[2]
port 15 nsew
flabel metal1 s 2639 1550 2682 1673 3 FreeSans 520 0 0 0 VPWR
port 17 nsew
flabel metal1 s 2649 2823 2726 2855 3 FreeSans 520 0 0 0 DM[1]
port 19 nsew
flabel metal1 s 2162 9 2205 210 3 FreeSans 520 0 0 0 VPWR
port 17 nsew
flabel metal1 s 2639 1702 2682 1904 3 FreeSans 520 0 0 0 VCC_IO
port 18 nsew
flabel metal1 s 2638 1544 2681 1674 3 FreeSans 520 0 0 0 VPWR
port 17 nsew
flabel metal1 s 4346 238 4430 286 3 FreeSans 520 0 0 0 STARTUP_ST_H
port 20 nsew
flabel metal1 s 2162 707 2205 906 3 FreeSans 520 0 0 0 VGND
port 21 nsew
flabel metal1 s 9377 2017 9470 2069 3 FreeSans 520 0 0 0 STARTUP_RST_H
port 22 nsew
flabel metal1 s 14191 2103 14243 2143 3 FreeSans 520 180 0 0 HLD_I_H_N
port 16 nsew
flabel metal1 s 14110 2025 14173 2062 3 FreeSans 520 0 0 0 OD_I_H
port 23 nsew
flabel metal1 s 15452 520 15523 558 3 FreeSans 520 270 0 0 IB_MODE_SEL_H_N
port 24 nsew
flabel metal1 s 15842 550 15873 608 3 FreeSans 520 180 0 0 IB_MODE_SEL_H
port 25 nsew
flabel metal1 s 14674 2027 14735 2056 3 FreeSans 520 0 0 0 IB_MODE_SEL
port 26 nsew
flabel metal1 s 14734 12 14774 64 3 FreeSans 520 270 0 0 HLD_I_H_N
port 16 nsew
<< properties >>
string GDS_END 21520892
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21489116
<< end >>
