magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect 0 2192 1504 2312
rect 4 2142 1500 2192
rect 4 1280 1500 1330
rect 0 1032 1504 1280
rect 4 982 1500 1032
rect 4 120 1500 170
rect 0 0 1504 120
<< mvndiff >>
rect 26 2278 92 2286
rect 26 2244 42 2278
rect 76 2244 92 2278
rect 26 2218 92 2244
rect 152 2278 218 2286
rect 152 2244 168 2278
rect 202 2244 218 2278
rect 152 2218 218 2244
rect 278 2278 344 2286
rect 278 2244 294 2278
rect 328 2244 344 2278
rect 278 2218 344 2244
rect 404 2278 470 2286
rect 404 2244 420 2278
rect 454 2244 470 2278
rect 404 2218 470 2244
rect 530 2278 596 2286
rect 530 2244 546 2278
rect 580 2244 596 2278
rect 530 2218 596 2244
rect 656 2278 722 2286
rect 656 2244 672 2278
rect 706 2244 722 2278
rect 656 2218 722 2244
rect 782 2278 848 2286
rect 782 2244 798 2278
rect 832 2244 848 2278
rect 782 2218 848 2244
rect 908 2278 974 2286
rect 908 2244 924 2278
rect 958 2244 974 2278
rect 908 2218 974 2244
rect 1034 2278 1100 2286
rect 1034 2244 1050 2278
rect 1084 2244 1100 2278
rect 1034 2218 1100 2244
rect 1160 2278 1226 2286
rect 1160 2244 1176 2278
rect 1210 2244 1226 2278
rect 1160 2218 1226 2244
rect 1286 2278 1352 2286
rect 1286 2244 1302 2278
rect 1336 2244 1352 2278
rect 1286 2218 1352 2244
rect 1412 2278 1478 2286
rect 1412 2244 1428 2278
rect 1462 2244 1478 2278
rect 1412 2218 1478 2244
rect 30 2210 88 2218
rect 30 2176 42 2210
rect 76 2176 88 2210
rect 30 2168 88 2176
rect 156 2210 214 2218
rect 156 2176 168 2210
rect 202 2176 214 2210
rect 156 2168 214 2176
rect 282 2210 340 2218
rect 282 2176 294 2210
rect 328 2176 340 2210
rect 282 2168 340 2176
rect 408 2210 466 2218
rect 408 2176 420 2210
rect 454 2176 466 2210
rect 408 2168 466 2176
rect 534 2210 592 2218
rect 534 2176 546 2210
rect 580 2176 592 2210
rect 534 2168 592 2176
rect 660 2210 718 2218
rect 660 2176 672 2210
rect 706 2176 718 2210
rect 660 2168 718 2176
rect 786 2210 844 2218
rect 786 2176 798 2210
rect 832 2176 844 2210
rect 786 2168 844 2176
rect 912 2210 970 2218
rect 912 2176 924 2210
rect 958 2176 970 2210
rect 912 2168 970 2176
rect 1038 2210 1096 2218
rect 1038 2176 1050 2210
rect 1084 2176 1096 2210
rect 1038 2168 1096 2176
rect 1164 2210 1222 2218
rect 1164 2176 1176 2210
rect 1210 2176 1222 2210
rect 1164 2168 1222 2176
rect 1290 2210 1348 2218
rect 1290 2176 1302 2210
rect 1336 2176 1348 2210
rect 1290 2168 1348 2176
rect 1416 2210 1474 2218
rect 1416 2176 1428 2210
rect 1462 2176 1474 2210
rect 1416 2168 1474 2176
rect 30 1296 88 1304
rect 30 1262 42 1296
rect 76 1262 88 1296
rect 30 1254 88 1262
rect 156 1296 214 1304
rect 156 1262 168 1296
rect 202 1262 214 1296
rect 156 1254 214 1262
rect 282 1296 340 1304
rect 282 1262 294 1296
rect 328 1262 340 1296
rect 282 1254 340 1262
rect 408 1296 466 1304
rect 408 1262 420 1296
rect 454 1262 466 1296
rect 408 1254 466 1262
rect 534 1296 592 1304
rect 534 1262 546 1296
rect 580 1262 592 1296
rect 534 1254 592 1262
rect 660 1296 718 1304
rect 660 1262 672 1296
rect 706 1262 718 1296
rect 660 1254 718 1262
rect 786 1296 844 1304
rect 786 1262 798 1296
rect 832 1262 844 1296
rect 786 1254 844 1262
rect 912 1296 970 1304
rect 912 1262 924 1296
rect 958 1262 970 1296
rect 912 1254 970 1262
rect 1038 1296 1096 1304
rect 1038 1262 1050 1296
rect 1084 1262 1096 1296
rect 1038 1254 1096 1262
rect 1164 1296 1222 1304
rect 1164 1262 1176 1296
rect 1210 1262 1222 1296
rect 1164 1254 1222 1262
rect 1290 1296 1348 1304
rect 1290 1262 1302 1296
rect 1336 1262 1348 1296
rect 1290 1254 1348 1262
rect 1416 1296 1474 1304
rect 1416 1262 1428 1296
rect 1462 1262 1474 1296
rect 1416 1254 1474 1262
rect 26 1228 92 1254
rect 26 1194 42 1228
rect 76 1194 92 1228
rect 26 1186 92 1194
rect 152 1228 218 1254
rect 152 1194 168 1228
rect 202 1194 218 1228
rect 152 1186 218 1194
rect 278 1228 344 1254
rect 278 1194 294 1228
rect 328 1194 344 1228
rect 278 1186 344 1194
rect 404 1228 470 1254
rect 404 1194 420 1228
rect 454 1194 470 1228
rect 404 1186 470 1194
rect 530 1228 596 1254
rect 530 1194 546 1228
rect 580 1194 596 1228
rect 530 1186 596 1194
rect 656 1228 722 1254
rect 656 1194 672 1228
rect 706 1194 722 1228
rect 656 1186 722 1194
rect 782 1228 848 1254
rect 782 1194 798 1228
rect 832 1194 848 1228
rect 782 1186 848 1194
rect 908 1228 974 1254
rect 908 1194 924 1228
rect 958 1194 974 1228
rect 908 1186 974 1194
rect 1034 1228 1100 1254
rect 1034 1194 1050 1228
rect 1084 1194 1100 1228
rect 1034 1186 1100 1194
rect 1160 1228 1226 1254
rect 1160 1194 1176 1228
rect 1210 1194 1226 1228
rect 1160 1186 1226 1194
rect 1286 1228 1352 1254
rect 1286 1194 1302 1228
rect 1336 1194 1352 1228
rect 1286 1186 1352 1194
rect 1412 1228 1478 1254
rect 1412 1194 1428 1228
rect 1462 1194 1478 1228
rect 1412 1186 1478 1194
rect 26 1118 92 1126
rect 26 1084 42 1118
rect 76 1084 92 1118
rect 26 1058 92 1084
rect 152 1118 218 1126
rect 152 1084 168 1118
rect 202 1084 218 1118
rect 152 1058 218 1084
rect 278 1118 344 1126
rect 278 1084 294 1118
rect 328 1084 344 1118
rect 278 1058 344 1084
rect 404 1118 470 1126
rect 404 1084 420 1118
rect 454 1084 470 1118
rect 404 1058 470 1084
rect 530 1118 596 1126
rect 530 1084 546 1118
rect 580 1084 596 1118
rect 530 1058 596 1084
rect 656 1118 722 1126
rect 656 1084 672 1118
rect 706 1084 722 1118
rect 656 1058 722 1084
rect 782 1118 848 1126
rect 782 1084 798 1118
rect 832 1084 848 1118
rect 782 1058 848 1084
rect 908 1118 974 1126
rect 908 1084 924 1118
rect 958 1084 974 1118
rect 908 1058 974 1084
rect 1034 1118 1100 1126
rect 1034 1084 1050 1118
rect 1084 1084 1100 1118
rect 1034 1058 1100 1084
rect 1160 1118 1226 1126
rect 1160 1084 1176 1118
rect 1210 1084 1226 1118
rect 1160 1058 1226 1084
rect 1286 1118 1352 1126
rect 1286 1084 1302 1118
rect 1336 1084 1352 1118
rect 1286 1058 1352 1084
rect 1412 1118 1478 1126
rect 1412 1084 1428 1118
rect 1462 1084 1478 1118
rect 1412 1058 1478 1084
rect 30 1050 88 1058
rect 30 1016 42 1050
rect 76 1016 88 1050
rect 30 1008 88 1016
rect 156 1050 214 1058
rect 156 1016 168 1050
rect 202 1016 214 1050
rect 156 1008 214 1016
rect 282 1050 340 1058
rect 282 1016 294 1050
rect 328 1016 340 1050
rect 282 1008 340 1016
rect 408 1050 466 1058
rect 408 1016 420 1050
rect 454 1016 466 1050
rect 408 1008 466 1016
rect 534 1050 592 1058
rect 534 1016 546 1050
rect 580 1016 592 1050
rect 534 1008 592 1016
rect 660 1050 718 1058
rect 660 1016 672 1050
rect 706 1016 718 1050
rect 660 1008 718 1016
rect 786 1050 844 1058
rect 786 1016 798 1050
rect 832 1016 844 1050
rect 786 1008 844 1016
rect 912 1050 970 1058
rect 912 1016 924 1050
rect 958 1016 970 1050
rect 912 1008 970 1016
rect 1038 1050 1096 1058
rect 1038 1016 1050 1050
rect 1084 1016 1096 1050
rect 1038 1008 1096 1016
rect 1164 1050 1222 1058
rect 1164 1016 1176 1050
rect 1210 1016 1222 1050
rect 1164 1008 1222 1016
rect 1290 1050 1348 1058
rect 1290 1016 1302 1050
rect 1336 1016 1348 1050
rect 1290 1008 1348 1016
rect 1416 1050 1474 1058
rect 1416 1016 1428 1050
rect 1462 1016 1474 1050
rect 1416 1008 1474 1016
rect 30 136 88 144
rect 30 102 42 136
rect 76 102 88 136
rect 30 94 88 102
rect 156 136 214 144
rect 156 102 168 136
rect 202 102 214 136
rect 156 94 214 102
rect 282 136 340 144
rect 282 102 294 136
rect 328 102 340 136
rect 282 94 340 102
rect 408 136 466 144
rect 408 102 420 136
rect 454 102 466 136
rect 408 94 466 102
rect 534 136 592 144
rect 534 102 546 136
rect 580 102 592 136
rect 534 94 592 102
rect 660 136 718 144
rect 660 102 672 136
rect 706 102 718 136
rect 660 94 718 102
rect 786 136 844 144
rect 786 102 798 136
rect 832 102 844 136
rect 786 94 844 102
rect 912 136 970 144
rect 912 102 924 136
rect 958 102 970 136
rect 912 94 970 102
rect 1038 136 1096 144
rect 1038 102 1050 136
rect 1084 102 1096 136
rect 1038 94 1096 102
rect 1164 136 1222 144
rect 1164 102 1176 136
rect 1210 102 1222 136
rect 1164 94 1222 102
rect 1290 136 1348 144
rect 1290 102 1302 136
rect 1336 102 1348 136
rect 1290 94 1348 102
rect 1416 136 1474 144
rect 1416 102 1428 136
rect 1462 102 1474 136
rect 1416 94 1474 102
rect 26 68 92 94
rect 26 34 42 68
rect 76 34 92 68
rect 26 26 92 34
rect 152 68 218 94
rect 152 34 168 68
rect 202 34 218 68
rect 152 26 218 34
rect 278 68 344 94
rect 278 34 294 68
rect 328 34 344 68
rect 278 26 344 34
rect 404 68 470 94
rect 404 34 420 68
rect 454 34 470 68
rect 404 26 470 34
rect 530 68 596 94
rect 530 34 546 68
rect 580 34 596 68
rect 530 26 596 34
rect 656 68 722 94
rect 656 34 672 68
rect 706 34 722 68
rect 656 26 722 34
rect 782 68 848 94
rect 782 34 798 68
rect 832 34 848 68
rect 782 26 848 34
rect 908 68 974 94
rect 908 34 924 68
rect 958 34 974 68
rect 908 26 974 34
rect 1034 68 1100 94
rect 1034 34 1050 68
rect 1084 34 1100 68
rect 1034 26 1100 34
rect 1160 68 1226 94
rect 1160 34 1176 68
rect 1210 34 1226 68
rect 1160 26 1226 34
rect 1286 68 1352 94
rect 1286 34 1302 68
rect 1336 34 1352 68
rect 1286 26 1352 34
rect 1412 68 1478 94
rect 1412 34 1428 68
rect 1462 34 1478 68
rect 1412 26 1478 34
<< ndiffc >>
rect 42 2176 76 2210
rect 168 2176 202 2210
rect 294 2176 328 2210
rect 420 2176 454 2210
rect 546 2176 580 2210
rect 672 2176 706 2210
rect 798 2176 832 2210
rect 924 2176 958 2210
rect 1050 2176 1084 2210
rect 1176 2176 1210 2210
rect 1302 2176 1336 2210
rect 1428 2176 1462 2210
rect 42 1262 76 1296
rect 168 1262 202 1296
rect 294 1262 328 1296
rect 420 1262 454 1296
rect 546 1262 580 1296
rect 672 1262 706 1296
rect 798 1262 832 1296
rect 924 1262 958 1296
rect 1050 1262 1084 1296
rect 1176 1262 1210 1296
rect 1302 1262 1336 1296
rect 1428 1262 1462 1296
rect 42 1016 76 1050
rect 168 1016 202 1050
rect 294 1016 328 1050
rect 420 1016 454 1050
rect 546 1016 580 1050
rect 672 1016 706 1050
rect 798 1016 832 1050
rect 924 1016 958 1050
rect 1050 1016 1084 1050
rect 1176 1016 1210 1050
rect 1302 1016 1336 1050
rect 1428 1016 1462 1050
rect 42 102 76 136
rect 168 102 202 136
rect 294 102 328 136
rect 420 102 454 136
rect 546 102 580 136
rect 672 102 706 136
rect 798 102 832 136
rect 924 102 958 136
rect 1050 102 1084 136
rect 1176 102 1210 136
rect 1302 102 1336 136
rect 1428 102 1462 136
<< mvndiffc >>
rect 42 2244 76 2278
rect 168 2244 202 2278
rect 294 2244 328 2278
rect 420 2244 454 2278
rect 546 2244 580 2278
rect 672 2244 706 2278
rect 798 2244 832 2278
rect 924 2244 958 2278
rect 1050 2244 1084 2278
rect 1176 2244 1210 2278
rect 1302 2244 1336 2278
rect 1428 2244 1462 2278
rect 42 1194 76 1228
rect 168 1194 202 1228
rect 294 1194 328 1228
rect 420 1194 454 1228
rect 546 1194 580 1228
rect 672 1194 706 1228
rect 798 1194 832 1228
rect 924 1194 958 1228
rect 1050 1194 1084 1228
rect 1176 1194 1210 1228
rect 1302 1194 1336 1228
rect 1428 1194 1462 1228
rect 42 1084 76 1118
rect 168 1084 202 1118
rect 294 1084 328 1118
rect 420 1084 454 1118
rect 546 1084 580 1118
rect 672 1084 706 1118
rect 798 1084 832 1118
rect 924 1084 958 1118
rect 1050 1084 1084 1118
rect 1176 1084 1210 1118
rect 1302 1084 1336 1118
rect 1428 1084 1462 1118
rect 42 34 76 68
rect 168 34 202 68
rect 294 34 328 68
rect 420 34 454 68
rect 546 34 580 68
rect 672 34 706 68
rect 798 34 832 68
rect 924 34 958 68
rect 1050 34 1084 68
rect 1176 34 1210 68
rect 1302 34 1336 68
rect 1428 34 1462 68
<< locali >>
rect 20 2278 58 2311
rect 20 2277 42 2278
rect 26 2244 42 2277
rect 76 2244 92 2277
rect 26 2176 92 2244
rect 152 2244 168 2278
rect 202 2244 294 2278
rect 328 2244 344 2278
rect 412 2278 450 2311
rect 412 2277 420 2278
rect 484 2277 546 2278
rect 152 2176 344 2244
rect 404 2244 420 2277
rect 454 2244 546 2277
rect 580 2244 596 2278
rect 404 2176 596 2244
rect 656 2244 672 2278
rect 706 2244 798 2278
rect 832 2244 848 2278
rect 916 2278 954 2311
rect 1446 2278 1484 2311
rect 916 2277 924 2278
rect 988 2277 1050 2278
rect 656 2176 848 2244
rect 908 2244 924 2277
rect 958 2244 1050 2277
rect 1084 2244 1100 2278
rect 908 2176 1100 2244
rect 1160 2244 1176 2278
rect 1210 2244 1302 2278
rect 1336 2244 1352 2278
rect 1160 2176 1352 2244
rect 1462 2277 1484 2278
rect 1412 2244 1428 2277
rect 1462 2244 1478 2277
rect 1412 2176 1478 2244
rect 26 1228 92 1296
rect 26 1194 42 1228
rect 76 1194 92 1228
rect 26 1118 92 1194
rect 26 1084 42 1118
rect 76 1084 92 1118
rect 26 1016 92 1084
rect 152 1228 218 1296
rect 152 1194 168 1228
rect 202 1194 218 1228
rect 152 1118 218 1194
rect 152 1084 168 1118
rect 202 1084 218 1118
rect 152 1016 218 1084
rect 278 1228 344 1296
rect 278 1194 294 1228
rect 328 1194 344 1228
rect 278 1118 344 1194
rect 278 1084 294 1118
rect 328 1084 344 1118
rect 278 1016 344 1084
rect 404 1228 470 1296
rect 404 1194 420 1228
rect 454 1194 470 1228
rect 404 1118 470 1194
rect 404 1084 420 1118
rect 454 1084 470 1118
rect 404 1016 470 1084
rect 530 1228 596 1296
rect 530 1194 546 1228
rect 580 1194 596 1228
rect 530 1118 596 1194
rect 530 1084 546 1118
rect 580 1084 596 1118
rect 530 1016 596 1084
rect 656 1228 722 1296
rect 656 1194 672 1228
rect 706 1194 722 1228
rect 656 1118 722 1194
rect 656 1084 672 1118
rect 706 1084 722 1118
rect 656 1016 722 1084
rect 782 1228 848 1296
rect 782 1194 798 1228
rect 832 1194 848 1228
rect 782 1118 848 1194
rect 782 1084 798 1118
rect 832 1084 848 1118
rect 782 1016 848 1084
rect 908 1228 974 1296
rect 908 1194 924 1228
rect 958 1194 974 1228
rect 908 1118 974 1194
rect 908 1084 924 1118
rect 958 1084 974 1118
rect 908 1016 974 1084
rect 1034 1228 1100 1296
rect 1034 1194 1050 1228
rect 1084 1194 1100 1228
rect 1034 1118 1100 1194
rect 1034 1084 1050 1118
rect 1084 1084 1100 1118
rect 1034 1016 1100 1084
rect 1160 1228 1226 1296
rect 1160 1194 1176 1228
rect 1210 1194 1226 1228
rect 1160 1118 1226 1194
rect 1160 1084 1176 1118
rect 1210 1084 1226 1118
rect 1160 1016 1226 1084
rect 1286 1228 1352 1296
rect 1286 1194 1302 1228
rect 1336 1194 1352 1228
rect 1286 1118 1352 1194
rect 1286 1084 1302 1118
rect 1336 1084 1352 1118
rect 1286 1016 1352 1084
rect 1412 1228 1478 1296
rect 1412 1194 1428 1228
rect 1462 1194 1478 1228
rect 1412 1118 1478 1194
rect 1412 1084 1428 1118
rect 1462 1084 1478 1118
rect 1412 1016 1478 1084
rect 26 68 218 136
rect 26 34 42 68
rect 76 34 168 68
rect 202 34 218 68
rect 278 68 470 136
rect 278 34 294 68
rect 328 34 420 68
rect 454 34 470 68
rect 530 68 722 136
rect 530 34 546 68
rect 580 34 672 68
rect 706 34 722 68
rect 782 68 974 136
rect 782 34 798 68
rect 832 34 924 68
rect 958 34 974 68
rect 1034 68 1226 136
rect 1034 34 1050 68
rect 1084 34 1176 68
rect 1210 34 1226 68
rect 1286 68 1478 136
rect 1286 34 1302 68
rect 1336 34 1428 68
rect 1462 34 1478 68
<< viali >>
rect -14 2277 20 2311
rect 58 2278 92 2311
rect 58 2277 76 2278
rect 76 2277 92 2278
rect 378 2277 412 2311
rect 450 2278 484 2311
rect 450 2277 454 2278
rect 454 2277 484 2278
rect 882 2277 916 2311
rect 954 2278 988 2311
rect 1412 2278 1446 2311
rect 954 2277 958 2278
rect 958 2277 988 2278
rect 1412 2277 1428 2278
rect 1428 2277 1446 2278
rect 1484 2277 1518 2311
<< metal1 >>
rect -26 2311 108 2317
rect -26 2277 -14 2311
rect 20 2277 58 2311
rect 92 2277 108 2311
rect -26 2271 108 2277
rect 109 2272 110 2316
rect 146 2272 147 2316
rect 148 2311 500 2317
rect 148 2277 378 2311
rect 412 2277 450 2311
rect 484 2277 500 2311
rect 148 2271 500 2277
rect 501 2272 502 2316
rect 538 2272 539 2316
rect 540 2311 1001 2317
rect 540 2277 882 2311
rect 916 2277 954 2311
rect 988 2277 1001 2311
rect 540 2271 1001 2277
rect 1002 2272 1003 2316
rect 1039 2272 1040 2316
rect 1041 2311 1530 2317
rect 1041 2277 1412 2311
rect 1446 2277 1484 2311
rect 1518 2277 1530 2311
rect 1041 2271 1530 2277
<< rmetal1 >>
rect 108 2316 110 2317
rect 108 2272 109 2316
rect 108 2271 110 2272
rect 146 2316 148 2317
rect 147 2272 148 2316
rect 500 2316 502 2317
rect 146 2271 148 2272
rect 500 2272 501 2316
rect 500 2271 502 2272
rect 538 2316 540 2317
rect 539 2272 540 2316
rect 1001 2316 1003 2317
rect 538 2271 540 2272
rect 1001 2272 1002 2316
rect 1001 2271 1003 2272
rect 1039 2316 1041 2317
rect 1040 2272 1041 2316
rect 1039 2271 1041 2272
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_0
timestamp 1701704242
transform 0 -1 88 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_1
timestamp 1701704242
transform 0 -1 214 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_2
timestamp 1701704242
transform 0 -1 214 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_3
timestamp 1701704242
transform 0 -1 88 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_4
timestamp 1701704242
transform 0 -1 466 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_5
timestamp 1701704242
transform 0 -1 340 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_6
timestamp 1701704242
transform 0 -1 466 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_7
timestamp 1701704242
transform 0 -1 340 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_8
timestamp 1701704242
transform 0 -1 844 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_9
timestamp 1701704242
transform 0 -1 970 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_10
timestamp 1701704242
transform 0 -1 844 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_11
timestamp 1701704242
transform 0 -1 970 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_12
timestamp 1701704242
transform 0 -1 718 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_13
timestamp 1701704242
transform 0 -1 592 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_14
timestamp 1701704242
transform 0 -1 718 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_15
timestamp 1701704242
transform 0 -1 592 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_16
timestamp 1701704242
transform 0 -1 1348 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_17
timestamp 1701704242
transform 0 -1 1474 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_18
timestamp 1701704242
transform 0 -1 1348 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_19
timestamp 1701704242
transform 0 -1 1474 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_20
timestamp 1701704242
transform 0 -1 1222 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_21
timestamp 1701704242
transform 0 -1 1096 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_22
timestamp 1701704242
transform 0 -1 1222 -1 0 1304
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_23
timestamp 1701704242
transform 0 -1 1096 -1 0 144
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_24
timestamp 1701704242
transform 0 -1 214 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_25
timestamp 1701704242
transform 0 -1 214 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_26
timestamp 1701704242
transform 0 -1 88 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_27
timestamp 1701704242
transform 0 -1 88 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_28
timestamp 1701704242
transform 0 -1 466 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_29
timestamp 1701704242
transform 0 -1 466 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_30
timestamp 1701704242
transform 0 -1 340 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_31
timestamp 1701704242
transform 0 -1 340 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_32
timestamp 1701704242
transform 0 -1 844 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_33
timestamp 1701704242
transform 0 -1 844 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_34
timestamp 1701704242
transform 0 -1 970 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_35
timestamp 1701704242
transform 0 -1 970 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_36
timestamp 1701704242
transform 0 -1 718 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_37
timestamp 1701704242
transform 0 -1 718 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_38
timestamp 1701704242
transform 0 -1 592 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_39
timestamp 1701704242
transform 0 -1 592 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_40
timestamp 1701704242
transform 0 -1 1348 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_41
timestamp 1701704242
transform 0 -1 1348 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_42
timestamp 1701704242
transform 0 -1 1474 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_43
timestamp 1701704242
transform 0 -1 1474 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_44
timestamp 1701704242
transform 0 -1 1222 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_45
timestamp 1701704242
transform 0 -1 1222 1 0 2168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_46
timestamp 1701704242
transform 0 -1 1096 1 0 1008
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_47
timestamp 1701704242
transform 0 -1 1096 1 0 2168
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 92 0 -1 2311
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 1518 0 -1 2311
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 484 0 -1 2311
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 988 0 -1 2311
box 0 0 1 1
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_0
timestamp 1701704242
transform 0 -1 92 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_1
timestamp 1701704242
transform 0 -1 92 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_2
timestamp 1701704242
transform 0 -1 218 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_3
timestamp 1701704242
transform 0 -1 218 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_4
timestamp 1701704242
transform 0 -1 974 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_5
timestamp 1701704242
transform 0 -1 470 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_6
timestamp 1701704242
transform 0 -1 470 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_7
timestamp 1701704242
transform 0 -1 344 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_8
timestamp 1701704242
transform 0 -1 344 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_9
timestamp 1701704242
transform 0 -1 848 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_10
timestamp 1701704242
transform 0 -1 848 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_11
timestamp 1701704242
transform 0 -1 974 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_12
timestamp 1701704242
transform 0 -1 722 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_13
timestamp 1701704242
transform 0 -1 722 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_14
timestamp 1701704242
transform 0 -1 596 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_15
timestamp 1701704242
transform 0 -1 596 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_16
timestamp 1701704242
transform 0 -1 1352 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_17
timestamp 1701704242
transform 0 -1 1352 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_18
timestamp 1701704242
transform 0 -1 1478 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_19
timestamp 1701704242
transform 0 -1 1478 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_20
timestamp 1701704242
transform 0 -1 1226 1 0 136
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_21
timestamp 1701704242
transform 0 -1 1226 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_22
timestamp 1701704242
transform 0 -1 1100 1 0 1296
box -68 -26 948 92
use nDFres_CDNS_524688791851650  nDFres_CDNS_524688791851650_23
timestamp 1701704242
transform 0 -1 1100 1 0 136
box -68 -26 948 92
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1701704242
transform -1 0 1093 0 -1 2317
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_1
timestamp 1701704242
transform -1 0 200 0 -1 2317
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_2
timestamp 1701704242
transform 1 0 448 0 -1 2317
box 0 0 1 1
<< labels >>
flabel metal1 s 20 2277 58 2311 0 FreeSans 400 0 0 0 r1
port 1 nsew
flabel metal1 s 1446 2277 1484 2311 0 FreeSans 400 0 0 0 r2
port 2 nsew
<< properties >>
string GDS_END 97488464
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97474920
<< end >>
