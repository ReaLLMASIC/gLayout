magic
tech sky130B
timestamp 1701704242
<< pwell >>
rect -13 -13 54 1206
<< psubdiff >>
rect 0 1181 41 1193
rect 0 1164 12 1181
rect 29 1164 41 1181
rect 0 1145 41 1164
rect 0 1128 12 1145
rect 29 1128 41 1145
rect 0 1109 41 1128
rect 0 1092 12 1109
rect 29 1092 41 1109
rect 0 1073 41 1092
rect 0 1056 12 1073
rect 29 1056 41 1073
rect 0 1037 41 1056
rect 0 1020 12 1037
rect 29 1020 41 1037
rect 0 1001 41 1020
rect 0 984 12 1001
rect 29 984 41 1001
rect 0 965 41 984
rect 0 948 12 965
rect 29 948 41 965
rect 0 929 41 948
rect 0 912 12 929
rect 29 912 41 929
rect 0 893 41 912
rect 0 876 12 893
rect 29 876 41 893
rect 0 857 41 876
rect 0 840 12 857
rect 29 840 41 857
rect 0 821 41 840
rect 0 804 12 821
rect 29 804 41 821
rect 0 785 41 804
rect 0 768 12 785
rect 29 768 41 785
rect 0 749 41 768
rect 0 732 12 749
rect 29 732 41 749
rect 0 713 41 732
rect 0 696 12 713
rect 29 696 41 713
rect 0 677 41 696
rect 0 660 12 677
rect 29 660 41 677
rect 0 641 41 660
rect 0 624 12 641
rect 29 624 41 641
rect 0 605 41 624
rect 0 588 12 605
rect 29 588 41 605
rect 0 569 41 588
rect 0 552 12 569
rect 29 552 41 569
rect 0 533 41 552
rect 0 516 12 533
rect 29 516 41 533
rect 0 497 41 516
rect 0 480 12 497
rect 29 480 41 497
rect 0 461 41 480
rect 0 444 12 461
rect 29 444 41 461
rect 0 425 41 444
rect 0 408 12 425
rect 29 408 41 425
rect 0 389 41 408
rect 0 372 12 389
rect 29 372 41 389
rect 0 353 41 372
rect 0 336 12 353
rect 29 336 41 353
rect 0 317 41 336
rect 0 300 12 317
rect 29 300 41 317
rect 0 281 41 300
rect 0 264 12 281
rect 29 264 41 281
rect 0 245 41 264
rect 0 228 12 245
rect 29 228 41 245
rect 0 209 41 228
rect 0 192 12 209
rect 29 192 41 209
rect 0 173 41 192
rect 0 156 12 173
rect 29 156 41 173
rect 0 137 41 156
rect 0 120 12 137
rect 29 120 41 137
rect 0 101 41 120
rect 0 84 12 101
rect 29 84 41 101
rect 0 65 41 84
rect 0 48 12 65
rect 29 48 41 65
rect 0 29 41 48
rect 0 12 12 29
rect 29 12 41 29
rect 0 0 41 12
<< psubdiffcont >>
rect 12 1164 29 1181
rect 12 1128 29 1145
rect 12 1092 29 1109
rect 12 1056 29 1073
rect 12 1020 29 1037
rect 12 984 29 1001
rect 12 948 29 965
rect 12 912 29 929
rect 12 876 29 893
rect 12 840 29 857
rect 12 804 29 821
rect 12 768 29 785
rect 12 732 29 749
rect 12 696 29 713
rect 12 660 29 677
rect 12 624 29 641
rect 12 588 29 605
rect 12 552 29 569
rect 12 516 29 533
rect 12 480 29 497
rect 12 444 29 461
rect 12 408 29 425
rect 12 372 29 389
rect 12 336 29 353
rect 12 300 29 317
rect 12 264 29 281
rect 12 228 29 245
rect 12 192 29 209
rect 12 156 29 173
rect 12 120 29 137
rect 12 84 29 101
rect 12 48 29 65
rect 12 12 29 29
<< locali >>
rect 12 1181 29 1189
rect 12 1145 29 1164
rect 12 1109 29 1128
rect 12 1073 29 1092
rect 12 1037 29 1056
rect 12 1001 29 1020
rect 12 965 29 984
rect 12 929 29 948
rect 12 893 29 912
rect 12 857 29 876
rect 12 821 29 840
rect 12 785 29 804
rect 12 749 29 768
rect 12 713 29 732
rect 12 677 29 696
rect 12 641 29 660
rect 12 605 29 624
rect 12 569 29 588
rect 12 533 29 552
rect 12 497 29 516
rect 12 461 29 480
rect 12 425 29 444
rect 12 389 29 408
rect 12 353 29 372
rect 12 317 29 336
rect 12 281 29 300
rect 12 245 29 264
rect 12 209 29 228
rect 12 173 29 192
rect 12 137 29 156
rect 12 101 29 120
rect 12 65 29 84
rect 12 29 29 48
rect 12 4 29 12
<< properties >>
string GDS_END 88593092
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88590784
<< end >>
