magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 138 900 1592 2140
<< pwell >>
rect -108 86 -22 760
rect -108 0 1620 86
<< psubdiff >>
rect -82 710 -48 734
rect -82 641 -48 676
rect -82 572 -48 607
rect -82 503 -48 538
rect -82 434 -48 469
rect -82 364 -48 400
rect -82 294 -48 330
rect -82 224 -48 260
rect -82 154 -48 190
rect -82 84 -48 120
rect -48 50 -10 60
rect -82 26 -10 50
<< mvpsubdiff >>
rect -10 26 50 60
rect 84 26 121 60
rect 155 26 192 60
rect 226 26 263 60
rect 297 26 334 60
rect 368 26 405 60
rect 439 26 476 60
rect 510 26 547 60
rect 581 26 618 60
rect 652 26 689 60
rect 723 26 760 60
rect 794 26 831 60
rect 865 26 902 60
rect 936 26 973 60
rect 1007 26 1044 60
rect 1078 26 1115 60
rect 1149 26 1186 60
rect 1220 26 1256 60
rect 1290 26 1326 60
rect 1360 26 1396 60
rect 1430 26 1466 60
rect 1500 26 1536 60
rect 1570 26 1594 60
<< mvnsubdiff >>
rect 204 2040 228 2074
rect 262 2040 297 2074
rect 331 2040 366 2074
rect 400 2040 435 2074
rect 469 2040 504 2074
rect 538 2040 573 2074
rect 607 2040 642 2074
rect 676 2040 711 2074
rect 745 2040 780 2074
rect 814 2040 849 2074
rect 883 2040 918 2074
rect 952 2040 987 2074
rect 1021 2040 1056 2074
rect 1090 2040 1125 2074
rect 1159 2040 1194 2074
rect 1228 2040 1263 2074
rect 1297 2040 1332 2074
rect 1366 2040 1400 2074
rect 1434 2050 1526 2074
rect 1434 2040 1492 2050
rect 204 1982 238 2040
rect 204 1914 238 1948
rect 204 1846 238 1880
rect 204 1778 238 1812
rect 204 1710 238 1744
rect 204 1642 238 1676
rect 204 1574 238 1608
rect 204 1506 238 1540
rect 204 1438 238 1472
rect 204 1369 238 1404
rect 204 1300 238 1335
rect 204 1231 238 1266
rect 204 1162 238 1197
rect 204 1093 238 1128
rect 204 1024 238 1059
rect 204 966 238 990
rect 1492 1981 1526 2016
rect 1492 1912 1526 1947
rect 1492 1843 1526 1878
rect 1492 1774 1526 1809
rect 1492 1705 1526 1740
rect 1492 1636 1526 1671
rect 1492 1568 1526 1602
rect 1492 1500 1526 1534
rect 1492 1432 1526 1466
rect 1492 1364 1526 1398
rect 1492 1296 1526 1330
rect 1492 1228 1526 1262
rect 1492 1160 1526 1194
rect 1492 1092 1526 1126
rect 1492 1024 1526 1058
rect 1492 966 1526 990
<< psubdiffcont >>
rect -82 676 -48 710
rect -82 607 -48 641
rect -82 538 -48 572
rect -82 469 -48 503
rect -82 400 -48 434
rect -82 330 -48 364
rect -82 260 -48 294
rect -82 190 -48 224
rect -82 120 -48 154
rect -82 50 -48 84
<< mvpsubdiffcont >>
rect 50 26 84 60
rect 121 26 155 60
rect 192 26 226 60
rect 263 26 297 60
rect 334 26 368 60
rect 405 26 439 60
rect 476 26 510 60
rect 547 26 581 60
rect 618 26 652 60
rect 689 26 723 60
rect 760 26 794 60
rect 831 26 865 60
rect 902 26 936 60
rect 973 26 1007 60
rect 1044 26 1078 60
rect 1115 26 1149 60
rect 1186 26 1220 60
rect 1256 26 1290 60
rect 1326 26 1360 60
rect 1396 26 1430 60
rect 1466 26 1500 60
rect 1536 26 1570 60
<< mvnsubdiffcont >>
rect 228 2040 262 2074
rect 297 2040 331 2074
rect 366 2040 400 2074
rect 435 2040 469 2074
rect 504 2040 538 2074
rect 573 2040 607 2074
rect 642 2040 676 2074
rect 711 2040 745 2074
rect 780 2040 814 2074
rect 849 2040 883 2074
rect 918 2040 952 2074
rect 987 2040 1021 2074
rect 1056 2040 1090 2074
rect 1125 2040 1159 2074
rect 1194 2040 1228 2074
rect 1263 2040 1297 2074
rect 1332 2040 1366 2074
rect 1400 2040 1434 2074
rect 204 1948 238 1982
rect 204 1880 238 1914
rect 204 1812 238 1846
rect 204 1744 238 1778
rect 204 1676 238 1710
rect 204 1608 238 1642
rect 204 1540 238 1574
rect 204 1472 238 1506
rect 204 1404 238 1438
rect 204 1335 238 1369
rect 204 1266 238 1300
rect 204 1197 238 1231
rect 204 1128 238 1162
rect 204 1059 238 1093
rect 204 990 238 1024
rect 1492 2016 1526 2050
rect 1492 1947 1526 1981
rect 1492 1878 1526 1912
rect 1492 1809 1526 1843
rect 1492 1740 1526 1774
rect 1492 1671 1526 1705
rect 1492 1602 1526 1636
rect 1492 1534 1526 1568
rect 1492 1466 1526 1500
rect 1492 1398 1526 1432
rect 1492 1330 1526 1364
rect 1492 1262 1526 1296
rect 1492 1194 1526 1228
rect 1492 1126 1526 1160
rect 1492 1058 1526 1092
rect 1492 990 1526 1024
<< poly >>
rect 365 934 485 940
rect 541 934 661 940
rect 717 934 837 940
rect 893 934 1013 940
rect 1069 934 1189 940
rect 365 918 1189 934
rect 365 884 428 918
rect 462 884 496 918
rect 530 884 564 918
rect 598 884 1189 918
rect 365 868 1189 884
rect 79 760 727 868
rect 1245 826 1365 940
rect 893 810 1541 826
rect 893 776 956 810
rect 990 776 1024 810
rect 1058 776 1092 810
rect 1126 776 1301 810
rect 1335 776 1369 810
rect 1403 776 1437 810
rect 1471 776 1541 810
rect 893 760 1541 776
<< polycont >>
rect 428 884 462 918
rect 496 884 530 918
rect 564 884 598 918
rect 956 776 990 810
rect 1024 776 1058 810
rect 1092 776 1126 810
rect 1301 776 1335 810
rect 1369 776 1403 810
rect 1437 776 1471 810
<< locali >>
rect 204 2040 228 2074
rect 262 2040 297 2074
rect 331 2040 366 2074
rect 400 2040 435 2074
rect 469 2040 504 2074
rect 538 2040 573 2074
rect 607 2040 642 2074
rect 676 2040 711 2074
rect 745 2040 780 2074
rect 814 2040 849 2074
rect 883 2040 918 2074
rect 952 2040 987 2074
rect 1021 2040 1056 2074
rect 1090 2040 1125 2074
rect 1159 2040 1194 2074
rect 1228 2040 1263 2074
rect 1297 2040 1332 2074
rect 1366 2040 1400 2074
rect 1434 2050 1526 2074
rect 1434 2040 1492 2050
rect 204 1982 238 2040
rect 204 1914 238 1948
rect 496 1881 530 2040
rect 848 1892 882 2040
rect 1200 1892 1234 2040
rect 1492 1981 1526 2016
rect 1492 1912 1526 1947
rect 204 1846 238 1880
rect 204 1778 238 1812
rect 204 1710 238 1744
rect 1492 1843 1526 1878
rect 1492 1774 1526 1809
rect 354 1676 392 1710
rect 670 1676 708 1710
rect 1022 1676 1060 1710
rect 1338 1676 1376 1710
rect 1492 1705 1526 1740
rect 204 1642 238 1676
rect 204 1574 238 1608
rect 204 1506 238 1540
rect 204 1438 238 1472
rect 1492 1636 1526 1671
rect 1492 1568 1526 1602
rect 1492 1500 1526 1534
rect 1492 1432 1526 1466
rect 204 1369 238 1374
rect 204 1300 238 1302
rect 204 1264 238 1266
rect 496 1336 530 1374
rect 496 1264 530 1302
rect 848 1336 882 1374
rect 848 1264 882 1302
rect 1200 1336 1234 1374
rect 1200 1264 1234 1302
rect 1492 1364 1526 1374
rect 1492 1296 1526 1302
rect 204 1162 238 1197
rect 204 1093 238 1128
rect 204 1024 238 1059
rect 1492 1228 1526 1230
rect 1492 1160 1526 1194
rect 1492 1092 1526 1126
rect 204 966 238 990
rect 320 823 354 1045
rect 672 928 706 1025
rect 1024 928 1058 1028
rect 1376 928 1410 1036
rect 1492 1024 1526 1058
rect 1492 966 1526 990
rect 412 884 428 918
rect 462 884 496 918
rect 530 884 564 918
rect 598 884 614 918
rect 672 894 1410 928
rect 672 823 706 894
rect -82 739 -48 777
rect 210 772 706 823
rect 210 738 244 772
rect 562 738 596 772
rect 848 739 882 777
rect 940 776 956 810
rect 990 776 1024 810
rect 1058 776 1092 810
rect 1126 776 1142 810
rect 1200 739 1234 777
rect 1285 776 1301 810
rect 1335 776 1369 810
rect 1403 776 1437 810
rect 1471 776 1487 810
rect 1552 739 1586 777
rect -82 641 -48 676
rect -82 572 -48 607
rect -82 503 -48 538
rect -82 434 -48 469
rect -82 364 -48 400
rect -82 294 -48 330
rect -82 224 -48 260
rect 68 241 106 275
rect 384 241 422 275
rect 700 241 738 275
rect 1022 241 1060 275
rect 1374 241 1412 275
rect -82 154 -48 161
rect -82 84 -48 89
rect 848 195 882 196
rect 848 123 882 161
rect 848 60 882 89
rect 1200 195 1234 196
rect 1200 123 1234 161
rect 1200 60 1234 89
rect 1552 195 1586 196
rect 1552 123 1586 161
rect 1552 60 1586 89
rect -48 50 50 60
rect -82 26 50 50
rect 84 26 121 60
rect 155 26 192 60
rect 226 26 263 60
rect 297 26 334 60
rect 368 26 405 60
rect 439 26 476 60
rect 510 26 547 60
rect 581 26 618 60
rect 652 26 689 60
rect 723 26 760 60
rect 794 26 831 60
rect 865 26 902 60
rect 947 26 973 60
rect 1019 26 1044 60
rect 1091 26 1115 60
rect 1163 26 1186 60
rect 1220 26 1256 60
rect 1294 26 1326 60
rect 1366 26 1396 60
rect 1438 26 1466 60
rect 1510 26 1536 60
rect 1570 26 1594 60
<< viali >>
rect 320 1676 354 1710
rect 392 1676 426 1710
rect 636 1676 670 1710
rect 708 1676 742 1710
rect 988 1676 1022 1710
rect 1060 1676 1094 1710
rect 1304 1676 1338 1710
rect 1376 1676 1410 1710
rect 204 1404 238 1408
rect 204 1374 238 1404
rect 204 1335 238 1336
rect 204 1302 238 1335
rect 204 1231 238 1264
rect 204 1230 238 1231
rect 496 1374 530 1408
rect 496 1302 530 1336
rect 496 1230 530 1264
rect 848 1374 882 1408
rect 848 1302 882 1336
rect 848 1230 882 1264
rect 1200 1374 1234 1408
rect 1200 1302 1234 1336
rect 1200 1230 1234 1264
rect 1492 1398 1526 1408
rect 1492 1374 1526 1398
rect 1492 1330 1526 1336
rect 1492 1302 1526 1330
rect 1492 1262 1526 1264
rect 1492 1230 1526 1262
rect -82 777 -48 811
rect -82 710 -48 739
rect 848 777 882 811
rect 1200 777 1234 811
rect -82 705 -48 710
rect 848 705 882 739
rect 1552 777 1586 811
rect 1200 705 1234 739
rect 1552 705 1586 739
rect 34 241 68 275
rect 106 241 140 275
rect 350 241 384 275
rect 422 241 456 275
rect 666 241 700 275
rect 738 241 772 275
rect 988 241 1022 275
rect 1060 241 1094 275
rect 1340 241 1374 275
rect 1412 241 1446 275
rect -82 190 -48 195
rect -82 161 -48 190
rect -82 120 -48 123
rect -82 89 -48 120
rect 848 161 882 195
rect 848 89 882 123
rect 1200 161 1234 195
rect 1200 89 1234 123
rect 1552 161 1586 195
rect 1552 89 1586 123
rect 913 26 936 60
rect 936 26 947 60
rect 985 26 1007 60
rect 1007 26 1019 60
rect 1057 26 1078 60
rect 1078 26 1091 60
rect 1129 26 1149 60
rect 1149 26 1163 60
rect 1260 26 1290 60
rect 1290 26 1294 60
rect 1332 26 1360 60
rect 1360 26 1366 60
rect 1404 26 1430 60
rect 1430 26 1438 60
rect 1476 26 1500 60
rect 1500 26 1510 60
<< metal1 >>
rect 308 1710 1422 1716
rect 308 1676 320 1710
rect 354 1676 392 1710
rect 426 1676 636 1710
rect 670 1676 708 1710
rect 742 1676 988 1710
rect 1022 1676 1060 1710
rect 1094 1676 1304 1710
rect 1338 1676 1376 1710
rect 1410 1676 1422 1710
rect 308 1670 1422 1676
rect 198 1408 1592 1420
rect 198 1374 204 1408
rect 238 1374 496 1408
rect 530 1374 848 1408
rect 882 1374 1200 1408
rect 1234 1374 1492 1408
rect 1526 1374 1592 1408
rect 198 1336 1592 1374
rect 198 1302 204 1336
rect 238 1302 496 1336
rect 530 1302 848 1336
rect 882 1302 1200 1336
rect 1234 1302 1492 1336
rect 1526 1302 1592 1336
rect 198 1264 1592 1302
rect 198 1230 204 1264
rect 238 1230 496 1264
rect 530 1230 848 1264
rect 882 1230 1200 1264
rect 1234 1230 1492 1264
rect 1526 1230 1592 1264
rect 198 1218 1592 1230
rect -88 811 1592 823
rect -88 777 -82 811
rect -48 777 848 811
rect 882 777 1200 811
rect 1234 777 1552 811
rect 1586 777 1592 811
rect -88 739 1592 777
rect -88 705 -82 739
rect -48 705 848 739
rect 882 705 1200 739
rect 1234 705 1552 739
rect 1586 705 1592 739
rect -88 693 1592 705
rect 22 275 1458 281
rect 22 241 34 275
rect 68 241 106 275
rect 140 241 350 275
rect 384 241 422 275
rect 456 241 666 275
rect 700 241 738 275
rect 772 241 988 275
rect 1022 241 1060 275
rect 1094 241 1340 275
rect 1374 241 1412 275
rect 1446 241 1458 275
rect 22 235 1458 241
rect -88 195 1592 207
rect -88 161 -82 195
rect -48 161 848 195
rect 882 161 1200 195
rect 1234 161 1552 195
rect 1586 161 1592 195
rect -88 123 1592 161
rect -88 89 -82 123
rect -48 89 848 123
rect 882 89 1200 123
rect 1234 89 1552 123
rect 1586 89 1592 123
rect -88 77 1592 89
tri 66 66 77 77 ne
rect 77 66 1592 77
tri 77 60 83 66 ne
rect 83 60 1592 66
tri 83 26 117 60 ne
rect 117 26 913 60
rect 947 26 985 60
rect 1019 26 1057 60
rect 1091 26 1129 60
rect 1163 26 1260 60
rect 1294 26 1332 60
rect 1366 26 1404 60
rect 1438 26 1476 60
rect 1510 26 1592 60
tri 117 20 123 26 ne
rect 123 20 1592 26
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 1234 -1 0 195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 882 -1 0 195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 -1 -48 -1 0 195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 1 1552 1 0 705
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 0 1 848 1 0 705
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 1 1200 1 0 705
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 1 -82 1 0 705
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 -1 1586 1 0 89
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 1 0 34 0 -1 275
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 1 0 350 0 -1 275
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 1 0 666 0 -1 275
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 1 0 988 0 -1 275
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 1 0 1340 0 -1 275
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 1 0 636 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 1 0 320 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform 1 0 988 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1701704242
transform 1 0 1304 0 1 1676
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 530 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 882 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 1234 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 -1 1526 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1701704242
transform 0 -1 238 -1 0 1408
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1701704242
transform 1 0 913 0 1 26
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1701704242
transform 1 0 1260 0 1 26
box 0 0 1 1
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1701704242
transform 1 0 135 0 1 26
box -12 -6 694 40
use nfet_CDNS_52468879185450  nfet_CDNS_52468879185450_0
timestamp 1701704242
transform 1 0 893 0 -1 734
box -79 -26 727 626
use nfet_CDNS_52468879185450  nfet_CDNS_52468879185450_1
timestamp 1701704242
transform 1 0 79 0 -1 734
box -79 -26 727 626
use pfet_CDNS_52468879185313  pfet_CDNS_52468879185313_0
timestamp 1701704242
transform 1 0 1245 0 -1 1966
box -119 -66 239 1066
use pfet_CDNS_524688791851430  pfet_CDNS_524688791851430_0
timestamp 1701704242
transform -1 0 1189 0 -1 1966
box -119 -66 943 1066
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 -1 614 1 0 868
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1701704242
transform 0 -1 1142 1 0 760
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1701704242
transform 0 -1 1487 1 0 760
box 0 0 1 1
<< labels >>
flabel metal1 s 1546 20 1571 207 7 FreeSans 200 0 0 0 vgnd_io
port 1 nsew
flabel metal1 s 913 1670 963 1716 0 FreeSans 200 0 0 0 pu_h_n
port 3 nsew
flabel metal1 s 267 1218 301 1420 3 FreeSans 300 0 0 0 vcc_io
port 2 nsew
flabel locali s 496 884 530 918 0 FreeSans 400 0 0 0 drvhi_h
port 5 nsew
flabel locali s 1024 776 1058 810 0 FreeSans 400 0 0 0 puen_h
port 6 nsew
<< properties >>
string GDS_END 88142084
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88131948
string path 5.525 23.500 5.525 51.425 37.725 51.425 37.725 23.500 
<< end >>
