magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 89 197
<< metal1 >>
rect -6 197 95 200
rect -6 0 0 197
rect 89 0 95 197
rect -6 -3 95 0
<< properties >>
string GDS_END 86914536
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86913252
<< end >>
