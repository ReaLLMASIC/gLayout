magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 209 394 375 1126
<< pwell >>
rect -26 -106 401 -20
<< mvpsubdiff >>
rect 0 -80 34 -46
rect 68 -80 103 -46
rect 137 -80 171 -46
rect 205 -80 239 -46
rect 273 -80 307 -46
rect 341 -80 375 -46
<< mvnsubdiff >>
rect 275 1026 309 1060
rect 275 954 309 992
rect 275 883 309 920
rect 275 812 309 849
rect 275 741 309 778
rect 275 670 309 707
rect 275 599 309 636
rect 275 528 309 565
rect 275 460 309 494
<< mvpsubdiffcont >>
rect 34 -80 68 -46
rect 103 -80 137 -46
rect 171 -80 205 -46
rect 239 -80 273 -46
rect 307 -80 341 -46
<< mvnsubdiffcont >>
rect 275 992 309 1026
rect 275 920 309 954
rect 275 849 309 883
rect 275 778 309 812
rect 275 707 309 741
rect 275 636 309 670
rect 275 565 309 599
rect 275 494 309 528
<< poly >>
rect 28 400 148 437
rect 28 384 162 400
rect 28 350 44 384
rect 78 350 112 384
rect 146 357 162 384
rect 146 350 324 357
rect 28 254 324 350
<< polycont >>
rect 44 350 78 384
rect 112 350 146 384
<< locali >>
rect 275 1026 309 1060
rect 275 954 309 992
rect 275 883 309 920
rect 275 812 309 849
rect 275 741 309 778
rect -17 664 17 702
rect -17 592 17 630
rect 275 670 309 702
rect 275 599 309 630
rect 275 528 309 558
rect 159 446 241 522
rect 275 460 309 494
rect 196 434 241 446
rect 28 350 44 384
rect 78 350 112 384
rect 146 350 162 384
rect 196 281 252 434
rect 159 225 252 281
rect -17 138 17 176
rect -17 66 17 104
rect 335 138 369 176
rect 335 66 369 104
rect 0 -80 34 -46
rect 68 -80 103 -46
rect 137 -80 171 -46
rect 205 -80 239 -46
rect 273 -80 307 -46
rect 341 -80 375 -46
<< viali >>
rect -17 702 17 736
rect -17 630 17 664
rect -17 558 17 592
rect 275 707 309 736
rect 275 702 309 707
rect 275 636 309 664
rect 275 630 309 636
rect 275 565 309 592
rect 275 558 309 565
rect -17 176 17 210
rect -17 104 17 138
rect -17 32 17 66
rect 335 176 369 210
rect 335 104 369 138
rect 335 32 369 66
<< metal1 >>
rect -23 736 375 748
rect -23 702 -17 736
rect 17 702 275 736
rect 309 702 375 736
rect -23 664 375 702
rect -23 630 -17 664
rect 17 630 275 664
rect 309 630 375 664
rect -23 592 375 630
rect -23 558 -17 592
rect 17 558 275 592
rect 309 558 375 592
rect -23 546 375 558
rect -23 210 375 222
rect -23 176 -17 210
rect 17 176 335 210
rect 369 176 375 210
rect -23 138 375 176
rect -23 104 -17 138
rect 17 104 335 138
rect 369 104 375 138
rect -23 66 375 104
rect -23 32 -17 66
rect 17 32 335 66
rect 369 32 375 66
rect -23 20 375 32
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 17 -1 0 210
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 369 -1 0 210
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 309 1 0 558
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 -1 17 1 0 558
box 0 0 1 1
use nfet_CDNS_52468879185131  nfet_CDNS_52468879185131_0
timestamp 1701704242
transform 1 0 28 0 1 28
box -79 -26 375 226
use pfet_CDNS_52468879185134  pfet_CDNS_52468879185134_0
timestamp 1701704242
transform 1 0 28 0 -1 1060
box -119 -66 239 666
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 28 1 0 334
box 0 0 1 1
<< labels >>
flabel metal1 s -23 546 0 748 3 FreeSans 400 0 0 0 vcc_io
port 1 nsew
flabel metal1 s -23 20 0 222 3 FreeSans 400 0 0 0 vgnd
port 2 nsew
flabel locali s 196 350 232 384 0 FreeSans 200 0 0 0 out
port 4 nsew
flabel locali s 78 350 112 384 0 FreeSans 600 0 0 0 in
port 5 nsew
<< properties >>
string GDS_END 85584338
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85581502
string path 7.300 27.150 7.300 10.850 
<< end >>
