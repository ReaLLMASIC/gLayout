magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 506
rect 413 0 416 506
<< via1 >>
rect 3 0 413 506
<< metal2 >>
rect 0 0 3 506
rect 413 0 416 506
<< properties >>
string GDS_END 88493224
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88479780
<< end >>
