magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -36 679 404 1471
<< pwell >>
rect 232 25 334 159
<< psubdiff >>
rect 258 109 308 133
rect 258 75 266 109
rect 300 75 308 109
rect 258 51 308 75
<< nsubdiff >>
rect 258 1339 308 1363
rect 258 1305 266 1339
rect 300 1305 308 1339
rect 258 1281 308 1305
<< psubdiffcont >>
rect 266 75 300 109
<< nsubdiffcont >>
rect 266 1305 300 1339
<< poly >>
rect 114 724 144 937
rect 48 708 144 724
rect 48 674 64 708
rect 98 674 144 708
rect 48 658 144 674
rect 114 413 144 658
<< polycont >>
rect 64 674 98 708
<< locali >>
rect 0 1397 368 1431
rect 62 1130 96 1397
rect 266 1339 300 1397
rect 266 1289 300 1305
rect 64 708 98 724
rect 64 658 98 674
rect 162 708 196 1196
rect 162 674 213 708
rect 162 186 196 674
rect 62 17 96 186
rect 266 109 300 125
rect 266 17 300 75
rect 0 -17 368 17
use contact_12  contact_12_0
timestamp 1701704242
transform 1 0 48 0 1 658
box 0 0 1 1
use contact_23  contact_23_0
timestamp 1701704242
transform 1 0 258 0 1 1281
box 0 0 1 1
use contact_24  contact_24_0
timestamp 1701704242
transform 1 0 258 0 1 51
box 0 0 1 1
use nmos_m7_w1_680_sli_dli_da_p  nmos_m7_w1_680_sli_dli_da_p_0
timestamp 1701704242
transform 1 0 54 0 1 51
box -26 -26 176 362
use pmos_m7_w2_000_sli_dli_da_p  pmos_m7_w2_000_sli_dli_da_p_0
timestamp 1701704242
transform 1 0 54 0 1 963
box -59 -54 209 454
<< labels >>
rlabel locali s 196 691 196 691 4 Z
port 2 nsew
rlabel locali s 81 691 81 691 4 A
port 1 nsew
rlabel locali s 184 1414 184 1414 4 vdd
port 3 nsew
rlabel locali s 184 0 184 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1414
string GDS_END 48928
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 47210
<< end >>
