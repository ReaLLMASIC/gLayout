magic
tech sky130B
magscale 1 2
timestamp 1701807570
<< obsli1 >>
rect 1830 39689 14025 39939
rect 14469 39876 14535 39884
rect 14449 39842 14555 39876
rect 1830 33880 2080 39689
rect 2220 39367 13631 39545
rect 2220 34083 2398 39367
rect 3156 39074 3298 39108
rect 3558 39074 3700 39108
rect 4076 39074 4218 39108
rect 4478 39074 4620 39108
rect 4996 39074 5138 39108
rect 5398 39074 5540 39108
rect 5916 39074 6058 39108
rect 6318 39074 6460 39108
rect 6836 39074 6978 39108
rect 7238 39074 7380 39108
rect 7756 39074 7898 39108
rect 8158 39074 8300 39108
rect 8676 39074 8818 39108
rect 9078 39074 9220 39108
rect 9596 39074 9738 39108
rect 9998 39074 10140 39108
rect 10516 39074 10658 39108
rect 10918 39074 11060 39108
rect 11436 39074 11578 39108
rect 11838 39074 11980 39108
rect 12356 39074 12498 39108
rect 12758 39074 12900 39108
rect 2877 37032 3087 39037
rect 3373 37105 3479 39011
rect 3797 39002 3975 39015
rect 3377 37065 3479 37105
rect 3769 37032 4007 39002
rect 4293 37105 4399 39011
rect 4717 39002 4895 39006
rect 4297 37065 4399 37105
rect 4689 37032 4927 39002
rect 5213 37105 5319 39011
rect 5637 39002 5815 39006
rect 5217 37065 5319 37105
rect 5609 37032 5847 39002
rect 6133 37105 6239 39011
rect 6557 39002 6735 39006
rect 6137 37065 6239 37105
rect 6529 37032 6767 39002
rect 7053 37105 7159 39011
rect 7477 39002 7655 39006
rect 7057 37065 7159 37105
rect 7449 37032 7687 39002
rect 7973 37105 8079 39011
rect 8397 39002 8575 39006
rect 7977 37065 8079 37105
rect 8369 37032 8607 39002
rect 8893 37105 8999 39011
rect 9317 39002 9495 39006
rect 8897 37065 8999 37105
rect 9289 37032 9527 39002
rect 9813 37105 9919 39011
rect 10237 39002 10415 39006
rect 9817 37065 9919 37105
rect 10209 37032 10447 39002
rect 10733 37105 10839 39011
rect 11157 39002 11335 39028
rect 10737 37065 10839 37105
rect 11129 37032 11367 39002
rect 11653 37105 11759 39011
rect 12077 39002 12255 39028
rect 11657 37065 11759 37105
rect 12049 37032 12287 39002
rect 12573 37105 12679 39011
rect 12577 37065 12679 37105
rect 12969 37032 13175 39036
rect 2566 36514 13337 36998
rect 3156 36468 13337 36514
rect 2225 33981 2395 34083
rect 1834 33830 2072 33880
rect 1702 32531 2072 33830
rect 2154 32531 2395 33981
rect 1834 26908 2072 32531
rect 2225 31783 2395 32531
rect 2877 32432 3087 36386
rect 3377 36139 3479 36407
rect 3373 32505 3479 36139
rect 3377 32465 3479 32505
rect 3769 32432 4007 36374
rect 4297 36139 4399 36407
rect 4293 32505 4399 36139
rect 4297 32465 4399 32505
rect 4689 32432 4927 36374
rect 5217 36139 5319 36407
rect 5213 32505 5319 36139
rect 5217 32465 5319 32505
rect 5609 32432 5847 36374
rect 6137 36139 6239 36407
rect 6133 32505 6239 36139
rect 6137 32465 6239 32505
rect 6529 32432 6767 36374
rect 7057 36139 7159 36407
rect 7053 32505 7159 36139
rect 7057 32465 7159 32505
rect 7449 32432 7687 36374
rect 7977 36139 8079 36407
rect 7973 32505 8079 36139
rect 7977 32465 8079 32505
rect 8369 32432 8607 36374
rect 8897 36139 8999 36407
rect 8893 32505 8999 36139
rect 8897 32465 8999 32505
rect 9289 32432 9527 36374
rect 9817 36139 9919 36407
rect 9813 32505 9919 36139
rect 9817 32465 9919 32505
rect 10209 32432 10447 36374
rect 10737 36139 10839 36407
rect 10733 32505 10839 36139
rect 10737 32465 10839 32505
rect 11129 32432 11367 36374
rect 11657 36139 11759 36407
rect 11653 32505 11759 36139
rect 11657 32465 11759 32505
rect 12049 32432 12287 36374
rect 12577 36139 12679 36407
rect 12573 32505 12679 36139
rect 12577 32465 12679 32505
rect 12969 32432 13175 36386
rect 13453 33209 13631 39367
rect 13458 33129 13628 33209
rect 2480 31911 12900 32398
rect 3156 31868 12900 31911
rect 2225 27233 2420 31783
rect 2877 27832 3087 31786
rect 3377 31539 3479 31807
rect 3373 27905 3479 31539
rect 3377 27865 3479 27905
rect 3769 27832 4007 31774
rect 4297 31539 4399 31807
rect 4293 27905 4399 31539
rect 4297 27865 4399 27905
rect 4689 27832 4927 31774
rect 5217 31539 5319 31807
rect 5213 27905 5319 31539
rect 5217 27865 5319 27905
rect 5609 27832 5847 31774
rect 6137 31539 6239 31807
rect 6133 27905 6239 31539
rect 6137 27865 6239 27905
rect 6529 27832 6767 31774
rect 7057 31539 7159 31807
rect 7053 27905 7159 31539
rect 7057 27865 7159 27905
rect 7449 27832 7687 31774
rect 7977 31539 8079 31807
rect 7973 27905 8079 31539
rect 7977 27865 8079 27905
rect 8369 27832 8607 31774
rect 8897 31539 8999 31807
rect 8893 27905 8999 31539
rect 8897 27865 8999 27905
rect 9289 27832 9527 31774
rect 9817 31539 9919 31807
rect 9813 27905 9919 31539
rect 9817 27865 9919 27905
rect 10209 27832 10447 31774
rect 10737 31539 10839 31807
rect 10733 27905 10839 31539
rect 10737 27865 10839 27905
rect 11129 27832 11367 31774
rect 11657 31539 11759 31807
rect 11653 27905 11759 31539
rect 11657 27865 11759 27905
rect 12049 27832 12287 31774
rect 12577 31539 12679 31807
rect 12573 27905 12679 31539
rect 12577 27865 12679 27905
rect 12969 27832 13175 31786
rect 3156 27308 12900 27798
rect 4996 27274 12900 27308
rect 5134 27268 12900 27274
rect 2225 27063 4532 27233
rect 1834 26670 4198 26908
rect 1840 26641 2838 26670
rect 3567 26629 4198 26670
rect 3913 19500 4198 26629
rect 3960 19379 4198 19500
rect 4362 19490 4532 27063
rect 4717 23232 4927 27186
rect 5217 26939 5319 27207
rect 5213 23305 5319 26939
rect 5217 23265 5319 23305
rect 5609 23232 5847 27174
rect 6137 26939 6239 27207
rect 6133 23305 6239 26939
rect 6137 23265 6239 23305
rect 6529 23232 6767 27174
rect 7057 26939 7159 27207
rect 7053 23305 7159 26939
rect 7057 23265 7159 23305
rect 7449 23232 7687 27174
rect 7977 26939 8079 27207
rect 7973 23305 8079 26939
rect 7977 23265 8079 23305
rect 8369 23232 8607 27174
rect 8897 26939 8999 27207
rect 8893 23305 8999 26939
rect 8897 23265 8999 23305
rect 9289 23232 9527 27174
rect 9817 26939 9919 27207
rect 9813 23305 9919 26939
rect 9817 23265 9919 23305
rect 10209 23232 10447 27174
rect 10737 26939 10839 27207
rect 10733 23305 10839 26939
rect 10737 23265 10839 23305
rect 11129 23232 11367 27174
rect 11657 26939 11759 27207
rect 11653 23305 11759 26939
rect 11657 23265 11759 23305
rect 12049 23232 12287 27174
rect 12577 26939 12679 27207
rect 12573 23305 12679 26939
rect 12577 23265 12679 23305
rect 12969 23232 13175 27186
rect 4611 22668 12900 23198
rect 3682 14874 3748 14877
rect 1900 14870 1966 14871
rect 1881 14836 1987 14870
rect 3682 14840 3800 14874
rect 3682 14837 3748 14840
rect 3960 14564 4217 19379
rect 1827 14314 4217 14564
rect 1827 8951 2077 14314
rect 4358 14173 4536 19490
rect 4717 18632 4927 22586
rect 5217 22339 5319 22607
rect 5213 18705 5319 22339
rect 5217 18665 5319 18705
rect 5609 18632 5847 22574
rect 6137 22339 6239 22607
rect 6133 18705 6239 22339
rect 6137 18665 6239 18705
rect 6529 18632 6767 22574
rect 7057 22339 7159 22607
rect 7053 18705 7159 22339
rect 7057 18665 7159 18705
rect 7449 18632 7687 22574
rect 7977 22339 8079 22607
rect 7973 18705 8079 22339
rect 7977 18665 8079 18705
rect 8369 18632 8607 22574
rect 8897 22339 8999 22607
rect 8893 18705 8999 22339
rect 8897 18665 8999 18705
rect 9289 18632 9527 22574
rect 9817 22339 9919 22607
rect 9813 18705 9919 22339
rect 9817 18665 9919 18705
rect 10209 18632 10447 22574
rect 10737 22339 10839 22607
rect 10733 18705 10839 22339
rect 10737 18665 10839 18705
rect 11129 18632 11367 22574
rect 11657 22339 11759 22607
rect 11653 18705 11759 22339
rect 11657 18665 11759 18705
rect 12049 18632 12287 22574
rect 12577 22339 12679 22607
rect 12573 18705 12679 22339
rect 12577 18665 12679 18705
rect 12969 18632 13175 22587
rect 13458 20342 13631 33129
rect 13458 20263 13628 20342
rect 4605 18099 12900 18598
rect 4996 18074 12900 18099
rect 5134 18068 12900 18074
rect 2221 13995 4536 14173
rect 4717 14032 4927 17986
rect 5217 17739 5319 18007
rect 5213 14105 5319 17739
rect 5217 14065 5319 14105
rect 5609 14032 5847 17974
rect 6137 17739 6239 18007
rect 6133 14105 6239 17739
rect 6137 14065 6239 14105
rect 6529 14032 6767 17974
rect 7057 17739 7159 18007
rect 7053 14105 7159 17739
rect 7057 14065 7159 14105
rect 7449 14032 7687 17974
rect 7977 17739 8079 18007
rect 7973 14105 8079 17739
rect 7977 14065 8079 14105
rect 8369 14032 8607 17974
rect 8897 17739 8999 18007
rect 8893 14105 8999 17739
rect 8897 14065 8999 14105
rect 9289 14032 9527 17974
rect 9817 17739 9919 18007
rect 9813 14105 9919 17739
rect 9817 14065 9919 14105
rect 10209 14032 10447 17974
rect 10737 17739 10839 18007
rect 10733 14105 10839 17739
rect 10737 14065 10839 14105
rect 11129 14032 11367 17974
rect 11657 17739 11759 18007
rect 11653 14105 11759 17739
rect 11657 14065 11759 14105
rect 12049 14032 12287 17974
rect 12577 17739 12679 18007
rect 12573 14105 12679 17739
rect 12577 14065 12679 14105
rect 12969 14032 13175 17986
rect 2221 9270 2399 13995
rect 4702 13799 12900 13998
rect 2617 9398 2651 13593
rect 3141 13468 12900 13799
rect 2877 9432 3087 13386
rect 3377 13139 3479 13407
rect 3373 9505 3479 13139
rect 3377 9465 3479 9505
rect 3769 9432 4007 13374
rect 4297 13139 4399 13407
rect 4293 9505 4399 13139
rect 4297 9465 4399 9505
rect 4689 9432 4927 13374
rect 5217 13139 5319 13407
rect 5213 9505 5319 13139
rect 5217 9465 5319 9505
rect 5609 9432 5847 13374
rect 6137 13139 6239 13407
rect 6133 9505 6239 13139
rect 6137 9465 6239 9505
rect 6529 9432 6767 13374
rect 7057 13139 7159 13407
rect 7053 9505 7159 13139
rect 7057 9465 7159 9505
rect 7449 9432 7687 13374
rect 7977 13139 8079 13407
rect 7973 9505 8079 13139
rect 7977 9465 8079 9505
rect 8369 9432 8607 13374
rect 8897 13139 8999 13407
rect 8893 9505 8999 13139
rect 8897 9465 8999 9505
rect 9289 9432 9527 13374
rect 9817 13139 9919 13407
rect 9813 9505 9919 13139
rect 9817 9465 9919 9505
rect 10209 9432 10447 13374
rect 10737 13139 10839 13407
rect 10733 9505 10839 13139
rect 10737 9465 10839 9505
rect 11129 9432 11367 13374
rect 11657 13139 11759 13407
rect 11653 9505 11759 13139
rect 11657 9465 11759 9505
rect 12049 9432 12287 13374
rect 12577 13139 12679 13407
rect 12573 9505 12679 13139
rect 12577 9465 12679 9505
rect 12969 9432 13175 13386
rect 2617 9363 12900 9398
rect 2618 9348 12900 9363
rect 13453 9270 13631 20263
rect 2221 9092 13631 9270
rect 13775 9237 14025 39689
rect 13781 9199 14019 9237
rect 13775 8951 14025 9199
rect 229 8688 263 8762
rect 1827 8701 14025 8951
rect 214 8654 280 8688
rect 1610 8654 1738 8688
rect 14145 8598 14211 8603
rect 14094 8564 14211 8598
rect 14145 8547 14211 8564
rect 10464 8291 13773 8499
rect 626 7913 9640 7917
rect 620 7739 9640 7913
rect 620 5606 804 7739
rect 947 7485 9191 7519
rect 947 5886 981 7485
rect 1268 7394 9012 7446
rect 1223 5956 1257 7314
rect 1379 5955 1413 7314
rect 1535 5956 1569 7314
rect 1691 5954 1725 7314
rect 1847 5956 1881 7314
rect 2003 5955 2037 7314
rect 2159 5956 2193 7314
rect 2315 5954 2349 7314
rect 2471 5956 2505 7314
rect 2627 5955 2661 7314
rect 2783 5956 2817 7314
rect 2939 5954 2973 7314
rect 3095 5956 3129 7314
rect 3251 5954 3285 7314
rect 3407 5956 3441 7314
rect 3563 5954 3597 7314
rect 3719 5956 3753 7314
rect 3875 5955 3909 7314
rect 4031 5956 4065 7314
rect 4187 5954 4221 7314
rect 4343 5956 4377 7314
rect 4499 5955 4533 7314
rect 4655 5956 4689 7314
rect 4811 5954 4845 7314
rect 4967 5956 5001 7314
rect 5123 5955 5157 7314
rect 5279 5956 5313 7314
rect 5435 5954 5469 7314
rect 5591 5956 5625 7314
rect 5747 5955 5781 7314
rect 5903 5956 5937 7314
rect 6059 5954 6093 7314
rect 6215 5956 6249 7314
rect 6371 5955 6405 7314
rect 6527 5956 6561 7314
rect 6683 5954 6717 7314
rect 6839 5956 6873 7314
rect 6995 5955 7029 7314
rect 7151 5956 7185 7314
rect 7307 5954 7341 7314
rect 7463 5956 7497 7314
rect 7619 5955 7653 7314
rect 7775 5956 7809 7314
rect 7931 5954 7965 7314
rect 8087 5956 8121 7314
rect 8243 5954 8277 7314
rect 8399 5956 8433 7314
rect 8555 5955 8589 7314
rect 8711 5956 8745 7314
rect 8867 5954 8901 7314
rect 9023 5956 9057 7314
rect 9151 5886 9191 7485
rect 9462 5905 9640 7739
rect 10464 6212 10642 8291
rect 13595 8263 13773 8291
rect 10792 8082 13428 8116
rect 13600 8096 13766 8263
rect 10792 6401 10826 8082
rect 10988 7954 13267 7988
rect 10938 7858 10972 7870
rect 10938 7238 10973 7858
rect 10938 6512 10972 7238
rect 11094 7154 11128 7870
rect 11093 6524 11128 7154
rect 11094 6512 11128 6524
rect 11250 7858 11284 7870
rect 11250 7238 11285 7858
rect 11250 6512 11284 7238
rect 11406 7154 11440 7870
rect 11405 6524 11440 7154
rect 11406 6512 11440 6524
rect 11562 7858 11596 7870
rect 11562 7238 11597 7858
rect 11562 6512 11596 7238
rect 11718 7154 11752 7870
rect 11717 6524 11752 7154
rect 11718 6512 11752 6524
rect 11874 7858 11908 7870
rect 11874 7238 11909 7858
rect 11874 6512 11908 7238
rect 12030 7154 12064 7870
rect 12029 6524 12064 7154
rect 12030 6512 12064 6524
rect 12186 7858 12220 7870
rect 12186 7238 12221 7858
rect 12186 6512 12220 7238
rect 12342 7154 12376 7870
rect 12341 6524 12376 7154
rect 12342 6512 12376 6524
rect 12498 7858 12532 7870
rect 12498 7238 12533 7858
rect 12498 6512 12532 7238
rect 12654 7154 12688 7870
rect 12653 6524 12688 7154
rect 12654 6512 12688 6524
rect 12810 7858 12844 7870
rect 12810 7238 12845 7858
rect 12810 6512 12844 7238
rect 12966 7154 13000 7870
rect 12965 6524 13000 7154
rect 12966 6512 13000 6524
rect 13122 7858 13156 7870
rect 13122 7238 13157 7858
rect 13122 6512 13156 7238
rect 13278 7154 13312 7870
rect 13387 7255 13428 8082
rect 13394 7213 13428 7255
rect 13277 6524 13312 7154
rect 13278 6512 13312 6524
rect 13387 6401 13428 7213
rect 10792 6367 13428 6401
rect 13595 6212 13773 8096
rect 947 5846 9191 5886
rect 9466 5843 9636 5905
rect 10464 5860 13773 6212
rect 9462 5606 9640 5843
rect 620 5432 9640 5606
rect 626 5428 9640 5432
rect 11043 5669 14126 5860
rect 11043 4648 11221 5669
rect 11364 5497 13714 5543
rect 11364 4696 11410 5497
rect 11518 5286 11552 5433
rect 12374 5286 12408 5433
rect 11511 4696 11557 5286
rect 12370 4696 12416 5286
rect 12516 4696 12562 5497
rect 12670 5286 12704 5433
rect 13526 5286 13560 5433
rect 12663 4696 12709 5286
rect 13522 4696 13568 5286
rect 13668 4696 13714 5497
rect 2413 4470 11221 4648
rect 2413 4446 11217 4470
rect 2413 378 2609 4446
rect 11370 4299 11404 4696
rect 11518 4483 11552 4696
rect 12374 4483 12408 4696
rect 11563 4347 12363 4393
rect 12522 4299 12556 4696
rect 12670 4483 12704 4696
rect 13526 4483 13560 4696
rect 12715 4347 13515 4393
rect 13674 4299 13708 4696
rect 13948 4504 14126 5669
rect 2756 4253 13714 4299
rect 2756 3452 2802 4253
rect 2910 4042 2944 4189
rect 3766 4042 3800 4189
rect 2903 3452 2949 4042
rect 3762 3452 3808 4042
rect 3908 3452 3954 4253
rect 4062 4042 4096 4189
rect 5718 4042 5752 4189
rect 4055 3452 4101 4042
rect 5714 3452 5760 4042
rect 5860 3452 5906 4253
rect 6014 4042 6048 4189
rect 7670 4042 7704 4189
rect 6007 3452 6053 4042
rect 7666 3452 7712 4042
rect 7812 3452 7858 4253
rect 7966 4042 8000 4189
rect 9622 4042 9656 4189
rect 7959 3452 8005 4042
rect 9618 3452 9664 4042
rect 9764 3452 9810 4253
rect 9918 4042 9952 4189
rect 11574 4042 11608 4189
rect 9911 3452 9957 4042
rect 11570 3452 11616 4042
rect 11716 3452 11762 4253
rect 11870 4042 11904 4189
rect 13526 4042 13560 4189
rect 11863 3452 11909 4042
rect 13522 3452 13568 4042
rect 13668 3452 13714 4253
rect 13956 4247 14126 4504
rect 2762 3055 2796 3452
rect 2910 3239 2944 3452
rect 3766 3239 3800 3452
rect 2955 3103 3755 3149
rect 3914 3055 3948 3452
rect 4062 3239 4096 3452
rect 5718 3239 5752 3452
rect 4107 3103 5707 3149
rect 5866 3055 5900 3452
rect 6014 3239 6048 3452
rect 7670 3239 7704 3452
rect 6059 3103 7659 3149
rect 7818 3055 7852 3452
rect 7966 3239 8000 3452
rect 9622 3239 9656 3452
rect 8011 3103 9611 3149
rect 9770 3055 9804 3452
rect 9918 3239 9952 3452
rect 11574 3239 11608 3452
rect 9963 3103 11563 3149
rect 11722 3055 11756 3452
rect 11870 3239 11904 3452
rect 13526 3239 13560 3452
rect 11915 3103 13515 3149
rect 13674 3055 13708 3452
rect 13953 3233 14126 4247
rect 2756 3009 13714 3055
rect 2756 2208 2802 3009
rect 2910 2798 2944 2945
rect 3766 2798 3800 2945
rect 2903 2208 2949 2798
rect 3762 2208 3808 2798
rect 3908 2208 3954 3009
rect 4062 2798 4096 2945
rect 5718 2798 5752 2945
rect 4055 2208 4101 2798
rect 5714 2208 5760 2798
rect 5860 2208 5906 3009
rect 6014 2798 6048 2945
rect 7670 2798 7704 2945
rect 6007 2208 6053 2798
rect 7666 2208 7712 2798
rect 7812 2208 7858 3009
rect 7966 2798 8000 2945
rect 9622 2798 9656 2945
rect 7959 2208 8005 2798
rect 9618 2208 9664 2798
rect 9764 2208 9810 3009
rect 9918 2798 9952 2945
rect 11574 2798 11608 2945
rect 9911 2208 9957 2798
rect 11570 2208 11616 2798
rect 11716 2208 11762 3009
rect 11870 2798 11904 2945
rect 13526 2798 13560 2945
rect 11863 2208 11909 2798
rect 13522 2208 13568 2798
rect 13668 2208 13714 3009
rect 13956 2983 14126 3233
rect 2762 1811 2796 2208
rect 2910 1995 2944 2208
rect 3766 1995 3800 2208
rect 2955 1859 3755 1905
rect 3914 1811 3948 2208
rect 4062 1995 4096 2208
rect 5718 1995 5752 2208
rect 4107 1859 5707 1905
rect 5866 1811 5900 2208
rect 6014 1995 6048 2208
rect 7670 1995 7704 2208
rect 6059 1859 7659 1905
rect 7818 1811 7852 2208
rect 7966 1995 8000 2208
rect 9622 1995 9656 2208
rect 8011 1859 9611 1905
rect 9770 1811 9804 2208
rect 9918 1995 9952 2208
rect 11574 1995 11608 2208
rect 9963 1859 11563 1905
rect 11722 1811 11756 2208
rect 11870 1995 11904 2208
rect 13526 1995 13560 2208
rect 11915 1859 13515 1905
rect 13674 1811 13708 2208
rect 13953 1969 14126 2983
rect 2756 1765 13714 1811
rect 13956 1783 14126 1969
rect 2756 964 2802 1765
rect 2910 1554 2944 1701
rect 3766 1554 3800 1701
rect 2903 964 2949 1554
rect 3762 964 3808 1554
rect 3908 964 3954 1765
rect 4062 1554 4096 1701
rect 5718 1554 5752 1701
rect 4055 964 4101 1554
rect 5714 964 5760 1554
rect 5860 964 5906 1765
rect 6014 1554 6048 1701
rect 7670 1554 7704 1701
rect 6007 964 6053 1554
rect 7666 964 7712 1554
rect 7812 964 7858 1765
rect 7966 1554 8000 1701
rect 9622 1554 9656 1701
rect 7959 964 8005 1554
rect 9618 964 9664 1554
rect 9764 964 9810 1765
rect 9918 1554 9952 1701
rect 11574 1554 11608 1701
rect 9911 964 9957 1554
rect 11570 964 11616 1554
rect 11716 964 11762 1765
rect 11870 1554 11904 1701
rect 13526 1554 13560 1701
rect 11863 964 11909 1554
rect 13522 964 13568 1554
rect 13668 964 13714 1765
rect 2762 567 2796 964
rect 2910 751 2944 964
rect 3766 751 3800 964
rect 2955 615 3755 661
rect 3914 567 3948 964
rect 4062 751 4096 964
rect 5718 751 5752 964
rect 4107 615 5707 661
rect 5866 567 5900 964
rect 6014 751 6048 964
rect 7670 751 7704 964
rect 6059 615 7659 661
rect 7818 567 7852 964
rect 7966 751 8000 964
rect 9622 751 9656 964
rect 8011 615 9611 661
rect 9770 567 9804 964
rect 9918 751 9952 964
rect 11574 751 11608 964
rect 9963 615 11563 661
rect 11722 567 11756 964
rect 11870 751 11904 964
rect 13526 751 13560 964
rect 11915 615 13515 661
rect 13674 567 13708 964
rect 13953 769 14126 1783
rect 2762 527 13708 567
rect 13956 554 14126 769
rect 2796 521 3914 527
rect 3948 521 5866 527
rect 5900 521 7818 527
rect 7852 521 9770 527
rect 9804 521 11722 527
rect 11756 521 13674 527
rect 13952 378 14130 554
rect 2413 200 14130 378
<< obsm1 >>
rect 0 0 15000 40000
<< metal2 >>
rect 201 38112 13440 39015
rect 201 38099 3006 38112
rect 201 38085 2992 38099
rect 201 38071 2978 38085
rect 201 38057 2964 38071
rect 201 38043 2950 38057
rect 201 38031 2936 38043
rect 201 37973 2880 38031
rect 201 37959 2866 37973
rect 201 37945 2852 37959
rect 201 37931 2838 37945
rect 201 37010 2824 37931
rect 3124 37059 14858 38003
rect 11746 37052 14858 37059
rect 11760 37038 14858 37052
rect 201 36996 2825 37010
rect 11774 37024 14858 37038
rect 11788 37010 14858 37024
rect 201 36982 2839 36996
rect 11802 36996 14858 37010
rect 201 36968 2853 36982
rect 11816 36982 14858 36996
rect 201 36954 2867 36968
rect 11830 36968 14858 36982
rect 201 36940 2881 36954
rect 11844 36954 14858 36968
rect 201 36926 2895 36940
rect 11858 36940 14858 36954
rect 201 36912 2909 36926
rect 11872 36926 14858 36940
rect 201 36898 2923 36912
rect 11886 36912 14858 36926
rect 201 36884 2937 36898
rect 11900 36898 14858 36912
rect 201 36870 2951 36884
rect 11914 36884 14858 36898
rect 201 36856 2965 36870
rect 11928 36870 14858 36884
rect 201 36842 2979 36856
rect 11942 36856 14858 36870
rect 201 36828 2993 36842
rect 11956 36842 14858 36856
rect 201 36814 3007 36828
rect 11970 36828 14858 36842
rect 201 36800 3021 36814
rect 11984 36814 14858 36828
rect 201 36786 3035 36800
rect 11998 36800 14858 36814
rect 201 36772 3049 36786
rect 12012 36786 14858 36800
rect 201 36758 3063 36772
rect 12026 36772 14858 36786
rect 201 36744 3077 36758
rect 12040 36758 14858 36772
rect 201 36730 3091 36744
rect 12054 36744 14858 36758
rect 201 36716 3105 36730
rect 12068 36730 14858 36744
rect 201 36702 3119 36716
rect 12082 36716 14858 36730
rect 201 36688 3133 36702
rect 12096 36702 14858 36716
rect 201 36674 3147 36688
rect 12110 36688 14858 36702
rect 201 36660 3161 36674
rect 12124 36674 14858 36688
rect 201 36646 3175 36660
rect 12138 36660 14858 36674
rect 201 36632 3189 36646
rect 12152 36646 14858 36660
rect 201 36618 3203 36632
rect 12166 36632 14858 36646
rect 201 36604 3217 36618
rect 12180 36618 14858 36632
rect 201 36590 3231 36604
rect 12194 36604 14858 36618
rect 201 36576 3245 36590
rect 12208 36590 14858 36604
rect 201 36562 3259 36576
rect 201 36548 3273 36562
rect 201 36534 3287 36548
rect 201 36520 3301 36534
rect 201 36506 3315 36520
rect 201 36492 3329 36506
rect 201 36478 3343 36492
rect 201 36464 3357 36478
rect 201 36450 3371 36464
rect 201 36436 3385 36450
rect 201 36422 3399 36436
rect 201 36408 3413 36422
rect 201 36394 3427 36408
rect 201 36380 3441 36394
rect 201 36366 3455 36380
rect 201 36352 3469 36366
rect 201 36338 3483 36352
rect 201 36324 3497 36338
rect 201 36310 3511 36324
rect 201 36296 3525 36310
rect 201 34556 11592 36296
rect 201 34544 3524 34556
rect 201 34530 3510 34544
rect 201 34516 3496 34530
rect 201 34502 3482 34516
rect 201 34500 3468 34502
rect 12222 34931 14858 36590
rect 12213 34917 14858 34931
rect 12199 34903 14858 34917
rect 12194 34500 14858 34903
rect 201 34348 3318 34500
rect 201 34334 3314 34348
rect 201 34320 3300 34334
rect 201 34306 3286 34320
rect 201 34292 3272 34306
rect 201 34278 3258 34292
rect 201 34264 3244 34278
rect 201 34259 3230 34264
rect 11793 34497 14858 34500
rect 11779 34483 14858 34497
rect 11765 34469 14858 34483
rect 11751 34455 14858 34469
rect 11742 34259 14858 34455
rect 201 33900 2880 34259
rect 201 33886 2866 33900
rect 201 33872 2852 33886
rect 201 33858 2838 33872
rect 201 32410 2824 33858
rect 11541 34245 14858 34259
rect 11527 34231 14858 34245
rect 3361 32491 14858 34231
rect 11508 32488 14858 32491
rect 11522 32474 14858 32488
rect 11536 32460 14858 32474
rect 11550 32446 14858 32460
rect 11564 32432 14858 32446
rect 11578 32418 14858 32432
rect 201 32396 2830 32410
rect 11592 32404 14858 32418
rect 201 32382 2844 32396
rect 11606 32390 14858 32404
rect 201 32368 2858 32382
rect 11620 32376 14858 32390
rect 201 32354 2872 32368
rect 11634 32362 14858 32376
rect 201 32340 2886 32354
rect 11648 32348 14858 32362
rect 201 32326 2900 32340
rect 11662 32334 14858 32348
rect 201 32312 2914 32326
rect 11676 32320 14858 32334
rect 201 32298 2928 32312
rect 11690 32306 14858 32320
rect 201 32284 2942 32298
rect 11704 32292 14858 32306
rect 201 32270 2956 32284
rect 11718 32278 14858 32292
rect 201 32256 2970 32270
rect 11732 32264 14858 32278
rect 201 32242 2984 32256
rect 11746 32250 14858 32264
rect 201 32228 2998 32242
rect 11760 32236 14858 32250
rect 201 32214 3012 32228
rect 11774 32222 14858 32236
rect 201 32200 3026 32214
rect 11788 32208 14858 32222
rect 201 32186 3040 32200
rect 11802 32194 14858 32208
rect 201 32172 3054 32186
rect 11816 32180 14858 32194
rect 201 32158 3068 32172
rect 11830 32166 14858 32180
rect 201 32144 3082 32158
rect 11844 32152 14858 32166
rect 201 32130 3096 32144
rect 11858 32138 14858 32152
rect 201 32116 3110 32130
rect 11872 32124 14858 32138
rect 201 32102 3124 32116
rect 11886 32110 14858 32124
rect 201 32088 3138 32102
rect 11900 32096 14858 32110
rect 201 32074 3152 32088
rect 11914 32082 14858 32096
rect 201 32060 3166 32074
rect 11928 32068 14858 32082
rect 201 32046 3180 32060
rect 11942 32054 14858 32068
rect 201 32032 3194 32046
rect 11956 32040 14858 32054
rect 201 32018 3208 32032
rect 11970 32026 14858 32040
rect 201 32004 3222 32018
rect 11984 32012 14858 32026
rect 201 31990 3236 32004
rect 11998 31998 14858 32012
rect 201 31976 3250 31990
rect 12012 31984 14858 31998
rect 201 31962 3264 31976
rect 12026 31970 14858 31984
rect 201 31948 3278 31962
rect 12040 31956 14858 31970
rect 201 31934 3292 31948
rect 12054 31942 14858 31956
rect 201 31920 3306 31934
rect 12068 31928 14858 31942
rect 201 31906 3320 31920
rect 12082 31914 14858 31928
rect 201 31892 3334 31906
rect 12096 31900 14858 31914
rect 201 31878 3348 31892
rect 12110 31886 14858 31900
rect 201 31864 3362 31878
rect 12124 31872 14858 31886
rect 201 31850 3376 31864
rect 12138 31858 14858 31872
rect 201 31836 3390 31850
rect 12152 31844 14858 31858
rect 201 31822 3404 31836
rect 12166 31830 14858 31844
rect 201 31808 3418 31822
rect 12180 31816 14858 31830
rect 201 31794 3432 31808
rect 12194 31802 14858 31816
rect 201 31780 3446 31794
rect 12208 31788 14858 31802
rect 201 31766 3460 31780
rect 201 31752 3474 31766
rect 201 31738 3488 31752
rect 201 31724 3502 31738
rect 201 31710 3516 31724
rect 201 31696 3530 31710
rect 201 29956 11341 31696
rect 201 29943 3524 29956
rect 201 29929 3510 29943
rect 201 29915 3496 29929
rect 201 29901 3482 29915
rect 201 29900 3468 29901
rect 12222 30345 14858 31788
rect 12211 30331 14858 30345
rect 12197 30317 14858 30331
rect 12194 29900 14858 30317
rect 201 29747 3319 29900
rect 201 29733 3314 29747
rect 201 29719 3300 29733
rect 201 29705 3286 29719
rect 201 29691 3272 29705
rect 201 29677 3258 29691
rect 201 29663 3244 29677
rect 201 29659 3230 29663
rect 11777 29897 14858 29900
rect 11763 29883 14858 29897
rect 11749 29869 14858 29883
rect 11735 29855 14858 29869
rect 11726 29659 14858 29855
rect 201 29439 3014 29659
rect 201 29425 3006 29439
rect 201 29411 2992 29425
rect 201 29397 2978 29411
rect 201 29383 2964 29397
rect 201 29369 2950 29383
rect 201 29355 2936 29369
rect 201 29354 2922 29355
rect 11525 29645 14858 29659
rect 11511 29631 14858 29645
rect 3650 29622 14858 29631
rect 3641 29608 14858 29622
rect 3638 29354 14858 29608
rect 201 29299 2880 29354
rect 201 29285 2866 29299
rect 201 29271 2852 29285
rect 201 29257 2838 29271
rect 201 27824 2824 29257
rect 3375 29342 14858 29354
rect 3361 27891 14858 29342
rect 11508 27885 14858 27891
rect 11522 27871 14858 27885
rect 11536 27857 14858 27871
rect 11550 27843 14858 27857
rect 11564 27829 14858 27843
rect 201 27810 2834 27824
rect 11578 27815 14858 27829
rect 201 27796 2848 27810
rect 11592 27801 14858 27815
rect 201 27782 2862 27796
rect 11606 27787 14858 27801
rect 201 27768 2876 27782
rect 11620 27773 14858 27787
rect 201 27754 2890 27768
rect 11634 27759 14858 27773
rect 201 27740 2904 27754
rect 11648 27745 14858 27759
rect 201 27726 2918 27740
rect 11662 27731 14858 27745
rect 201 27712 2932 27726
rect 11676 27717 14858 27731
rect 201 27698 2946 27712
rect 11690 27703 14858 27717
rect 201 27684 2960 27698
rect 11704 27689 14858 27703
rect 201 27670 2974 27684
rect 11718 27675 14858 27689
rect 201 27656 2988 27670
rect 11732 27661 14858 27675
rect 201 27642 3002 27656
rect 11746 27647 14858 27661
rect 201 27628 3016 27642
rect 11760 27633 14858 27647
rect 201 27614 3030 27628
rect 11774 27619 14858 27633
rect 201 27600 3044 27614
rect 11788 27605 14858 27619
rect 201 27586 3058 27600
rect 11802 27591 14858 27605
rect 201 27572 3072 27586
rect 11816 27577 14858 27591
rect 201 27558 3086 27572
rect 11830 27563 14858 27577
rect 201 27544 3100 27558
rect 11844 27549 14858 27563
rect 201 27530 3114 27544
rect 11858 27535 14858 27549
rect 201 27516 3128 27530
rect 11872 27521 14858 27535
rect 201 27502 3142 27516
rect 11886 27507 14858 27521
rect 201 27488 3156 27502
rect 11900 27493 14858 27507
rect 201 27474 3170 27488
rect 11914 27479 14858 27493
rect 201 27460 3184 27474
rect 11928 27465 14858 27479
rect 201 27446 3198 27460
rect 11942 27451 14858 27465
rect 201 27432 3212 27446
rect 11956 27437 14858 27451
rect 201 27418 3226 27432
rect 11970 27423 14858 27437
rect 201 27404 3240 27418
rect 11984 27409 14858 27423
rect 201 27390 3254 27404
rect 11998 27395 14858 27409
rect 201 27376 3268 27390
rect 12012 27381 14858 27395
rect 201 27362 3282 27376
rect 12026 27367 14858 27381
rect 201 27348 3296 27362
rect 12040 27353 14858 27367
rect 201 27334 3310 27348
rect 12054 27339 14858 27353
rect 201 27320 3324 27334
rect 12068 27325 14858 27339
rect 201 27306 3338 27320
rect 12082 27311 14858 27325
rect 201 27292 3352 27306
rect 12096 27297 14858 27311
rect 201 27278 3366 27292
rect 12110 27283 14858 27297
rect 201 27264 3380 27278
rect 12124 27269 14858 27283
rect 201 27250 3394 27264
rect 12138 27255 14858 27269
rect 201 27236 3408 27250
rect 12152 27241 14858 27255
rect 201 27222 3422 27236
rect 12166 27227 14858 27241
rect 201 27208 3436 27222
rect 12180 27213 14858 27227
rect 201 27194 3450 27208
rect 12194 27199 14858 27213
rect 201 27180 3464 27194
rect 12208 27185 14858 27199
rect 201 27166 3478 27180
rect 201 27152 3492 27166
rect 201 27138 3506 27152
rect 201 27124 3520 27138
rect 201 27110 3534 27124
rect 201 27096 3548 27110
rect 201 25356 11341 27096
rect 201 25343 3538 25356
rect 201 25329 3524 25343
rect 201 25315 3510 25329
rect 201 25301 3496 25315
rect 201 25300 3482 25301
rect 12222 25731 14858 27185
rect 12211 25717 14858 25731
rect 12197 25703 14858 25717
rect 12194 25300 14858 25703
rect 201 25147 3333 25300
rect 201 25133 3328 25147
rect 201 25119 3314 25133
rect 201 25105 3300 25119
rect 201 25091 3286 25105
rect 201 25077 3272 25091
rect 201 25063 3258 25077
rect 201 25059 3244 25063
rect 11791 25297 14858 25300
rect 11777 25283 14858 25297
rect 11763 25269 14858 25283
rect 11749 25255 14858 25269
rect 11740 25059 14858 25255
rect 201 24685 2880 25059
rect 201 24671 2866 24685
rect 201 24657 2852 24671
rect 201 24643 2838 24657
rect 201 23210 2824 24643
rect 11539 25045 14858 25059
rect 11525 25031 14858 25045
rect 4964 23291 14858 25031
rect 11508 23278 14858 23291
rect 11522 23264 14858 23278
rect 11536 23250 14858 23264
rect 11550 23236 14858 23250
rect 11564 23222 14858 23236
rect 201 23196 2827 23210
rect 11578 23208 14858 23222
rect 201 23182 2841 23196
rect 11592 23194 14858 23208
rect 201 23168 2855 23182
rect 11606 23180 14858 23194
rect 201 23154 2869 23168
rect 11620 23166 14858 23180
rect 201 23140 2883 23154
rect 11634 23152 14858 23166
rect 201 23126 2897 23140
rect 11648 23138 14858 23152
rect 201 23112 2911 23126
rect 11662 23124 14858 23138
rect 201 23098 2925 23112
rect 11676 23110 14858 23124
rect 201 23084 2939 23098
rect 11690 23096 14858 23110
rect 201 23070 2953 23084
rect 11704 23082 14858 23096
rect 201 23056 2967 23070
rect 11718 23068 14858 23082
rect 201 23042 2981 23056
rect 11732 23054 14858 23068
rect 201 23028 2995 23042
rect 11746 23040 14858 23054
rect 201 23014 3009 23028
rect 11760 23026 14858 23040
rect 201 23000 3023 23014
rect 11774 23012 14858 23026
rect 201 22986 3037 23000
rect 11788 22998 14858 23012
rect 201 22972 3051 22986
rect 11802 22984 14858 22998
rect 201 22958 3065 22972
rect 11816 22970 14858 22984
rect 201 22944 3079 22958
rect 11830 22956 14858 22970
rect 201 22930 3093 22944
rect 11844 22942 14858 22956
rect 201 22916 3107 22930
rect 11858 22928 14858 22942
rect 201 22902 3121 22916
rect 11872 22914 14858 22928
rect 201 22888 3135 22902
rect 11886 22900 14858 22914
rect 201 22874 3149 22888
rect 11900 22886 14858 22900
rect 201 22860 3163 22874
rect 11914 22872 14858 22886
rect 201 22846 3177 22860
rect 11928 22858 14858 22872
rect 201 22832 3191 22846
rect 11942 22844 14858 22858
rect 201 22818 3205 22832
rect 11956 22830 14858 22844
rect 201 22804 3219 22818
rect 11970 22816 14858 22830
rect 201 22790 3233 22804
rect 11984 22802 14858 22816
rect 201 22776 3247 22790
rect 11998 22788 14858 22802
rect 201 22762 3261 22776
rect 12012 22774 14858 22788
rect 201 22748 3275 22762
rect 12026 22760 14858 22774
rect 201 22734 3289 22748
rect 12040 22746 14858 22760
rect 201 22720 3303 22734
rect 12054 22732 14858 22746
rect 201 22706 3317 22720
rect 12068 22718 14858 22732
rect 201 22692 3331 22706
rect 12082 22704 14858 22718
rect 201 22678 3345 22692
rect 12096 22690 14858 22704
rect 201 22664 3359 22678
rect 12110 22676 14858 22690
rect 201 22650 3373 22664
rect 12124 22662 14858 22676
rect 201 22636 3387 22650
rect 12138 22648 14858 22662
rect 201 22622 3401 22636
rect 12152 22634 14858 22648
rect 201 22608 3415 22622
rect 12166 22620 14858 22634
rect 201 22594 3429 22608
rect 12180 22606 14858 22620
rect 201 22580 3443 22594
rect 12194 22592 14858 22606
rect 201 22566 3457 22580
rect 12208 22578 14858 22592
rect 201 22552 3471 22566
rect 201 22538 3485 22552
rect 201 22524 3499 22538
rect 201 22510 3513 22524
rect 201 22496 3527 22510
rect 201 20756 11341 22496
rect 201 20748 3524 20756
rect 201 20734 3510 20748
rect 201 20720 3496 20734
rect 201 20706 3482 20720
rect 201 20700 3468 20706
rect 12222 21131 14858 22578
rect 12211 21117 14858 21131
rect 12197 21103 14858 21117
rect 12194 20700 14858 21103
rect 201 20538 3314 20700
rect 201 20524 3300 20538
rect 201 20510 3286 20524
rect 201 20496 3272 20510
rect 201 20482 3258 20496
rect 201 20468 3244 20482
rect 201 20459 3230 20468
rect 11791 20697 14858 20700
rect 11777 20683 14858 20697
rect 11763 20669 14858 20683
rect 11749 20655 14858 20669
rect 11740 20459 14858 20655
rect 201 20104 2880 20459
rect 201 20090 2866 20104
rect 201 20076 2852 20090
rect 201 20062 2838 20076
rect 201 18596 2824 20062
rect 11539 20445 14858 20459
rect 11525 20431 14858 20445
rect 4964 18691 14858 20431
rect 11522 18682 14858 18691
rect 11536 18668 14858 18682
rect 11550 18654 14858 18668
rect 11564 18640 14858 18654
rect 11578 18626 14858 18640
rect 11592 18612 14858 18626
rect 201 18582 2833 18596
rect 11606 18598 14858 18612
rect 201 18568 2847 18582
rect 11620 18584 14858 18598
rect 201 18554 2861 18568
rect 11634 18570 14858 18584
rect 201 18540 2875 18554
rect 11648 18556 14858 18570
rect 201 18526 2889 18540
rect 11662 18542 14858 18556
rect 201 18512 2903 18526
rect 11676 18528 14858 18542
rect 201 18498 2917 18512
rect 11690 18514 14858 18528
rect 201 18484 2931 18498
rect 11704 18500 14858 18514
rect 201 18470 2945 18484
rect 11718 18486 14858 18500
rect 201 18456 2959 18470
rect 11732 18472 14858 18486
rect 201 18442 2973 18456
rect 11746 18458 14858 18472
rect 201 18428 2987 18442
rect 11760 18444 14858 18458
rect 201 18414 3001 18428
rect 11774 18430 14858 18444
rect 201 18400 3015 18414
rect 11788 18416 14858 18430
rect 201 18386 3029 18400
rect 11802 18402 14858 18416
rect 201 18372 3043 18386
rect 11816 18388 14858 18402
rect 201 18358 3057 18372
rect 11830 18374 14858 18388
rect 201 18344 3071 18358
rect 11844 18360 14858 18374
rect 201 18330 3085 18344
rect 11858 18346 14858 18360
rect 201 18316 3099 18330
rect 11872 18332 14858 18346
rect 201 18302 3113 18316
rect 11886 18318 14858 18332
rect 201 18288 3127 18302
rect 11900 18304 14858 18318
rect 201 18274 3141 18288
rect 11914 18290 14858 18304
rect 201 18260 3155 18274
rect 11928 18276 14858 18290
rect 201 18246 3169 18260
rect 11942 18262 14858 18276
rect 201 18232 3183 18246
rect 11956 18248 14858 18262
rect 201 18218 3197 18232
rect 11970 18234 14858 18248
rect 201 18204 3211 18218
rect 11984 18220 14858 18234
rect 201 18190 3225 18204
rect 11998 18206 14858 18220
rect 201 18176 3239 18190
rect 12012 18192 14858 18206
rect 201 18162 3253 18176
rect 12026 18178 14858 18192
rect 201 18148 3267 18162
rect 12040 18164 14858 18178
rect 201 18134 3281 18148
rect 12054 18150 14858 18164
rect 201 18120 3295 18134
rect 12068 18136 14858 18150
rect 201 18106 3309 18120
rect 12082 18122 14858 18136
rect 201 18092 3323 18106
rect 12096 18108 14858 18122
rect 201 18078 3337 18092
rect 12110 18094 14858 18108
rect 201 18064 3351 18078
rect 12124 18080 14858 18094
rect 201 18050 3365 18064
rect 12138 18066 14858 18080
rect 201 18036 3379 18050
rect 12152 18052 14858 18066
rect 201 18022 3393 18036
rect 12166 18038 14858 18052
rect 201 18008 3407 18022
rect 12180 18024 14858 18038
rect 201 17994 3421 18008
rect 12194 18010 14858 18024
rect 201 17980 3435 17994
rect 12208 17996 14858 18010
rect 201 17966 3449 17980
rect 201 17952 3463 17966
rect 201 17938 3477 17952
rect 201 17924 3491 17938
rect 201 17910 3505 17924
rect 201 17896 3519 17910
rect 201 16156 11341 17896
rect 201 16148 3524 16156
rect 201 16134 3510 16148
rect 201 16120 3496 16134
rect 201 16106 3482 16120
rect 201 16100 3468 16106
rect 12222 16531 14858 17996
rect 12211 16517 14858 16531
rect 12197 16503 14858 16517
rect 12194 16100 14858 16503
rect 201 15938 3314 16100
rect 201 15924 3300 15938
rect 201 15910 3286 15924
rect 201 15896 3272 15910
rect 201 15882 3258 15896
rect 201 15868 3244 15882
rect 201 15859 3230 15868
rect 11791 16097 14858 16100
rect 11777 16083 14858 16097
rect 11763 16069 14858 16083
rect 11749 16055 14858 16069
rect 11740 15859 14858 16055
rect 201 15504 2880 15859
rect 201 15490 2866 15504
rect 201 15476 2852 15490
rect 201 15462 2838 15476
rect 201 13996 2824 15462
rect 11539 15845 14858 15859
rect 11525 15831 14858 15845
rect 4964 15121 14858 15831
rect 4962 15107 14858 15121
rect 4948 15093 14858 15107
rect 4936 14911 14858 15093
rect 4752 14897 14858 14911
rect 4738 14883 14858 14897
rect 3682 14831 14858 14883
rect 4740 14821 14858 14831
rect 4754 14807 14858 14821
rect 4768 14793 14858 14807
rect 4782 14779 14858 14793
rect 4796 14765 14858 14779
rect 4810 14751 14858 14765
rect 4824 14737 14858 14751
rect 4838 14723 14858 14737
rect 4852 14709 14858 14723
rect 4866 14695 14858 14709
rect 4880 14681 14858 14695
rect 4894 14667 14858 14681
rect 4908 14653 14858 14667
rect 4922 14639 14858 14653
rect 4936 14625 14858 14639
rect 4950 14611 14858 14625
rect 4964 14091 14858 14611
rect 11508 14084 14858 14091
rect 11522 14070 14858 14084
rect 11536 14056 14858 14070
rect 11550 14042 14858 14056
rect 11564 14028 14858 14042
rect 11578 14014 14858 14028
rect 11592 14000 14858 14014
rect 201 13982 2833 13996
rect 11606 13986 14858 14000
rect 201 13968 2847 13982
rect 11620 13972 14858 13986
rect 201 13954 2861 13968
rect 11634 13958 14858 13972
rect 201 13940 2875 13954
rect 11648 13944 14858 13958
rect 201 13926 2889 13940
rect 11662 13930 14858 13944
rect 201 13912 2903 13926
rect 11676 13916 14858 13930
rect 201 13898 2917 13912
rect 11690 13902 14858 13916
rect 201 13884 2931 13898
rect 11704 13888 14858 13902
rect 201 13870 2945 13884
rect 11718 13874 14858 13888
rect 201 13856 2959 13870
rect 11732 13860 14858 13874
rect 201 13842 2973 13856
rect 11746 13846 14858 13860
rect 201 13828 2987 13842
rect 11760 13832 14858 13846
rect 201 13814 3001 13828
rect 11774 13818 14858 13832
rect 201 13800 3015 13814
rect 11788 13804 14858 13818
rect 201 13786 3029 13800
rect 11802 13790 14858 13804
rect 201 13772 3043 13786
rect 11816 13776 14858 13790
rect 201 13758 3057 13772
rect 11830 13762 14858 13776
rect 201 13744 3071 13758
rect 11844 13748 14858 13762
rect 201 13730 3085 13744
rect 11858 13734 14858 13748
rect 201 13716 3099 13730
rect 11872 13720 14858 13734
rect 201 13702 3113 13716
rect 11886 13706 14858 13720
rect 201 13688 3127 13702
rect 11900 13692 14858 13706
rect 201 13674 3141 13688
rect 11914 13678 14858 13692
rect 201 13660 3155 13674
rect 11928 13664 14858 13678
rect 201 13646 3169 13660
rect 11942 13650 14858 13664
rect 201 13632 3183 13646
rect 11956 13636 14858 13650
rect 201 13618 3197 13632
rect 11970 13622 14858 13636
rect 201 13604 3211 13618
rect 11984 13608 14858 13622
rect 201 13590 3225 13604
rect 11998 13594 14858 13608
rect 201 13576 3239 13590
rect 12012 13580 14858 13594
rect 201 13562 3253 13576
rect 12026 13566 14858 13580
rect 201 13548 3267 13562
rect 12040 13552 14858 13566
rect 201 13534 3281 13548
rect 12054 13538 14858 13552
rect 201 13520 3295 13534
rect 12068 13524 14858 13538
rect 201 13506 3309 13520
rect 12082 13510 14858 13524
rect 201 13492 3323 13506
rect 12096 13496 14858 13510
rect 201 13478 3337 13492
rect 12110 13482 14858 13496
rect 201 13464 3351 13478
rect 12124 13468 14858 13482
rect 201 13450 3365 13464
rect 12138 13454 14858 13468
rect 201 13436 3379 13450
rect 12152 13440 14858 13454
rect 201 13422 3393 13436
rect 12166 13426 14858 13440
rect 201 13408 3407 13422
rect 12180 13412 14858 13426
rect 201 13394 3421 13408
rect 12194 13398 14858 13412
rect 201 13380 3435 13394
rect 12208 13384 14858 13398
rect 201 13366 3449 13380
rect 201 13352 3463 13366
rect 201 13338 3477 13352
rect 201 13324 3491 13338
rect 201 13310 3505 13324
rect 201 13296 3519 13310
rect 201 11556 11342 13296
rect 201 11543 3524 11556
rect 201 11529 3510 11543
rect 201 11515 3496 11529
rect 201 11501 3482 11515
rect 201 11500 3468 11501
rect 12222 11945 14858 13384
rect 12219 11931 14858 11945
rect 12205 11917 14858 11931
rect 12194 11500 14858 11917
rect 201 11347 3319 11500
rect 201 11333 3314 11347
rect 201 11319 3300 11333
rect 201 11305 3286 11319
rect 201 11291 3272 11305
rect 201 11277 3258 11291
rect 201 11263 3244 11277
rect 201 11259 3230 11263
rect 11785 11497 14858 11500
rect 11771 11483 14858 11497
rect 11757 11469 14858 11483
rect 11743 11455 14858 11469
rect 11734 11259 14858 11455
rect 201 11067 3041 11259
rect 201 11053 3034 11067
rect 201 11039 3020 11053
rect 201 11025 3006 11039
rect 201 11011 2992 11025
rect 201 10997 2978 11011
rect 201 10983 2964 10997
rect 201 10981 2950 10983
rect 11533 11245 14858 11259
rect 11519 11231 14858 11245
rect 3770 11219 14858 11231
rect 3758 10981 14858 11219
rect 201 10899 2880 10981
rect 201 10885 2866 10899
rect 201 10871 2852 10885
rect 201 10857 2838 10871
rect 201 9420 2824 10857
rect 202 9419 2824 9420
rect 210 9411 2824 9419
rect 218 9050 2824 9411
rect 3520 10967 14858 10981
rect 3506 10953 14858 10967
rect 3361 9491 14858 10953
rect 11508 9478 14858 9491
rect 11522 9464 14858 9478
rect 11536 9450 14858 9464
rect 11550 9436 14858 9450
rect 11564 9422 14858 9436
rect 11578 9408 14858 9422
rect 11592 9394 14858 9408
rect 11606 9380 14858 9394
rect 11620 9366 14858 9380
rect 11634 9352 14858 9366
rect 11648 9338 14858 9352
rect 11662 9324 14858 9338
rect 11676 9310 14858 9324
rect 11690 9296 14858 9310
rect 11704 9282 14858 9296
rect 11718 9268 14858 9282
rect 11732 9254 14858 9268
rect 11746 9240 14858 9254
rect 11760 9226 14858 9240
rect 11774 9212 14858 9226
rect 11788 9198 14858 9212
rect 11802 9184 14858 9198
rect 11816 9170 14858 9184
rect 11830 9156 14858 9170
rect 11844 9142 14858 9156
rect 11858 9128 14858 9142
rect 11872 9114 14858 9128
rect 11886 9100 14858 9114
rect 11900 9086 14858 9100
rect 11914 9072 14858 9086
rect 218 9036 2837 9050
rect 11928 9058 14858 9072
rect 218 9022 2851 9036
rect 11942 9044 14858 9058
rect 218 9008 2865 9022
rect 11956 9030 14858 9044
rect 218 8994 2879 9008
rect 11970 9016 14858 9030
rect 218 8980 2893 8994
rect 11984 9002 14858 9016
rect 218 8966 2907 8980
rect 11998 8988 14858 9002
rect 218 8952 2921 8966
rect 12012 8974 14858 8988
rect 218 8938 2935 8952
rect 12026 8960 14858 8974
rect 218 8924 2949 8938
rect 12040 8946 14858 8960
rect 218 8910 2963 8924
rect 12054 8932 14858 8946
rect 218 8896 2977 8910
rect 12068 8918 14858 8932
rect 218 8882 2991 8896
rect 12082 8904 14858 8918
rect 218 8868 3005 8882
rect 12096 8890 14858 8904
rect 218 8854 3019 8868
rect 12110 8876 14858 8890
rect 218 8840 3033 8854
rect 12124 8862 14858 8876
rect 218 8826 3047 8840
rect 12138 8848 14858 8862
rect 218 8812 3061 8826
rect 12152 8834 14858 8848
rect 218 8798 3075 8812
rect 12166 8820 14858 8834
rect 218 8784 3089 8798
rect 12180 8806 14858 8820
rect 218 8770 3103 8784
rect 12194 8792 14858 8806
rect 218 8756 3117 8770
rect 12208 8778 14858 8792
rect 218 8742 3131 8756
rect 218 8728 3145 8742
rect 218 8714 3159 8728
rect 218 8700 3173 8714
rect 218 8686 3187 8700
rect 218 8672 3201 8686
rect 218 8658 3215 8672
rect 218 8644 3229 8658
rect 218 8630 3243 8644
rect 218 8616 3257 8630
rect 218 8602 3271 8616
rect 218 8588 3285 8602
rect 218 8574 3299 8588
rect 218 8560 3313 8574
rect 218 8546 3327 8560
rect 218 8532 3341 8546
rect 218 8518 3355 8532
rect 218 8504 3369 8518
rect 218 8490 3383 8504
rect 218 8476 3397 8490
rect 218 8462 10840 8476
rect 218 8448 10854 8462
rect 218 8434 10868 8448
rect 218 8420 10882 8434
rect 218 8406 10896 8420
rect 218 8392 10910 8406
rect 218 8378 10924 8392
rect 218 8364 10938 8378
rect 218 8350 10952 8364
rect 218 8336 10966 8350
rect 218 8322 10980 8336
rect 218 8308 10994 8322
rect 218 8294 11008 8308
rect 218 8280 11022 8294
rect 218 8266 11036 8280
rect 218 8252 11050 8266
rect 218 8238 11064 8252
rect 218 8224 11078 8238
rect 218 8210 11092 8224
rect 218 8196 11106 8210
rect 218 8182 11120 8196
rect 218 8168 11134 8182
rect 218 8154 11148 8168
rect 218 8140 11162 8154
rect 218 8126 11176 8140
rect 218 8112 11190 8126
rect 218 8098 11204 8112
rect 218 8084 11218 8098
rect 218 8070 11232 8084
rect 218 8060 3968 8070
rect 218 8046 3954 8060
rect 10526 8059 11246 8070
rect 218 8032 3940 8046
rect 10540 8045 11257 8059
rect 218 8018 3926 8032
rect 218 8014 3912 8018
rect 10554 8031 11271 8045
rect 10568 8017 11285 8031
rect 218 7724 3627 8014
rect 10582 8003 11299 8017
rect 10596 7989 11313 8003
rect 10610 7975 11327 7989
rect 10624 7961 11341 7975
rect 10638 7947 11355 7961
rect 10652 7933 11369 7947
rect 10654 7931 11383 7933
rect 10668 7917 11383 7931
rect 10682 7903 11383 7917
rect 10696 7889 11383 7903
rect 10710 7875 11383 7889
rect 10724 7861 11383 7875
rect 10738 7847 11383 7861
rect 10752 7833 11383 7847
rect 10766 7819 11383 7833
rect 10780 7805 11383 7819
rect 10794 7791 11383 7805
rect 10808 7777 11383 7791
rect 10822 7763 11383 7777
rect 10836 7749 11383 7763
rect 10850 7735 11383 7749
rect 218 7710 3618 7724
rect 10864 7721 11383 7735
rect 218 7696 3604 7710
rect 10878 7707 11383 7721
rect 218 7682 3590 7696
rect 10892 7693 11383 7707
rect 218 7668 3576 7682
rect 10906 7679 11383 7693
rect 218 7654 3562 7668
rect 10920 7665 11383 7679
rect 218 7640 3548 7654
rect 218 7639 3534 7640
rect 218 7387 3182 7639
rect 217 7379 3182 7387
rect 209 7371 3182 7379
rect 201 7287 3182 7371
rect 201 7273 3181 7287
rect 201 7259 3167 7273
rect 201 7245 3153 7259
rect 201 7231 3139 7245
rect 201 7217 3125 7231
rect 201 7203 3111 7217
rect 201 7189 3097 7203
rect 10934 7223 11383 7665
rect 201 7175 3083 7189
rect 201 7161 3069 7175
rect 201 7147 3055 7161
rect 201 5854 3041 7147
rect 12222 6182 14858 8778
rect 12213 6168 14858 6182
rect 12199 6154 14858 6168
rect 12194 5886 14858 6154
rect 11919 5874 14858 5886
rect 11905 5860 14858 5874
rect 201 5840 3050 5854
rect 11891 5846 14858 5860
rect 201 5826 3064 5840
rect 201 5812 3078 5826
rect 201 5798 3092 5812
rect 201 5784 3106 5798
rect 201 5770 3120 5784
rect 201 5756 3134 5770
rect 201 5742 3148 5756
rect 201 5728 3162 5742
rect 201 5714 3176 5728
rect 201 5700 3190 5714
rect 201 5686 3204 5700
rect 201 5672 3218 5686
rect 201 5658 3232 5672
rect 201 5644 3246 5658
rect 201 5630 3260 5644
rect 201 5616 3274 5630
rect 201 5602 3288 5616
rect 201 5588 3302 5602
rect 201 5574 3316 5588
rect 201 5560 3330 5574
rect 201 5546 3344 5560
rect 201 5532 3358 5546
rect 201 5518 3372 5532
rect 201 5504 3386 5518
rect 201 5490 3400 5504
rect 201 5476 3414 5490
rect 201 5462 3428 5476
rect 201 5448 3442 5462
rect 201 5434 3456 5448
rect 201 5420 3470 5434
rect 201 5406 3484 5420
rect 201 5392 3498 5406
rect 201 5378 3512 5392
rect 201 5364 3526 5378
rect 201 5350 3540 5364
rect 201 5336 3554 5350
rect 201 5322 3568 5336
rect 201 5308 3582 5322
rect 201 5294 3596 5308
rect 201 5280 3610 5294
rect 201 5266 3624 5280
rect 201 5252 3638 5266
rect 201 5238 3652 5252
rect 201 5224 3666 5238
rect 201 5210 3680 5224
rect 201 5196 3694 5210
rect 11878 5196 14858 5846
rect 201 5182 3708 5196
rect 201 5168 3722 5182
rect 201 5154 3736 5168
rect 11233 5188 14858 5196
rect 11219 5174 14858 5188
rect 11205 5160 14858 5174
rect 201 5140 3750 5154
rect 201 2480 7379 5140
rect 201 2475 5635 2480
rect 201 2461 5621 2475
rect 201 2447 5607 2461
rect 201 2433 5593 2447
rect 201 2424 5579 2433
rect 11191 5146 14858 5160
rect 11177 5132 14858 5146
rect 7578 2459 14858 5132
rect 9350 2453 14858 2459
rect 9364 2439 14858 2453
rect 9378 2425 14858 2439
rect 201 1803 4953 2424
rect 9392 2411 14858 2425
rect 9406 2397 14858 2411
rect 9420 2383 14858 2397
rect 9434 2369 14858 2383
rect 9448 2355 14858 2369
rect 9462 2341 14858 2355
rect 9476 2327 14858 2341
rect 9490 2313 14858 2327
rect 9504 2299 14858 2313
rect 9518 2285 14858 2299
rect 9532 2271 14858 2285
rect 9546 2257 14858 2271
rect 9560 2243 14858 2257
rect 9574 2229 14858 2243
rect 9588 2215 14858 2229
rect 9602 2201 14858 2215
rect 9616 2187 14858 2201
rect 9630 2173 14858 2187
rect 9644 2159 14858 2173
rect 9658 2145 14858 2159
rect 9672 2131 14858 2145
rect 9686 2117 14858 2131
rect 9700 2103 14858 2117
rect 9714 2089 14858 2103
rect 9728 2075 14858 2089
rect 9742 2061 14858 2075
rect 9756 2047 14858 2061
rect 9770 2033 14858 2047
rect 9784 2019 14858 2033
rect 9798 2005 14858 2019
rect 9812 1991 14858 2005
rect 9826 1977 14858 1991
rect 9840 1963 14858 1977
rect 9854 1949 14858 1963
rect 9868 1935 14858 1949
rect 9882 1921 14858 1935
rect 9896 1907 14858 1921
rect 9910 1893 14858 1907
rect 9924 1879 14858 1893
rect 9938 1865 14858 1879
rect 9952 1851 14858 1865
rect 9966 1837 14858 1851
rect 9980 1823 14858 1837
rect 201 1789 4949 1803
rect 9994 1809 14858 1823
rect 201 1775 4935 1789
rect 10008 1795 14858 1809
rect 201 1761 4921 1775
rect 10022 1781 14858 1795
rect 201 1747 4907 1761
rect 10036 1767 14858 1781
rect 201 1733 4893 1747
rect 10050 1753 14858 1767
rect 201 509 4879 1733
rect 10064 1739 14858 1753
rect 197 495 4879 509
rect 183 481 4879 495
rect 169 467 4879 481
rect 155 453 4879 467
rect 145 434 4879 453
rect 127 425 4879 434
rect 113 411 4879 425
rect 99 0 4879 411
rect 5179 0 5579 107
rect 10078 0 14858 1739
<< obsm2 >>
rect 0 39071 15000 40000
rect 0 9396 145 39071
rect 13496 38056 15000 39071
rect 3017 38031 15000 38056
rect 2880 37034 3096 38031
rect 2883 37031 3096 37034
rect 2897 37017 3068 37031
rect 2911 37003 3068 37017
rect 3350 37003 11727 37031
rect 2913 37001 11727 37003
rect 2927 36987 11727 37001
rect 2941 36973 11732 36987
rect 2955 36959 11746 36973
rect 2969 36945 11760 36959
rect 2983 36931 11774 36945
rect 2997 36917 11788 36931
rect 3011 36903 11802 36917
rect 3025 36889 11816 36903
rect 3039 36875 11830 36889
rect 3053 36861 11844 36875
rect 3067 36847 11858 36861
rect 3081 36833 11872 36847
rect 3095 36819 11886 36833
rect 3109 36805 11900 36819
rect 3123 36791 11914 36805
rect 3137 36777 11928 36791
rect 3151 36763 11942 36777
rect 3165 36749 11956 36763
rect 3179 36735 11970 36749
rect 3193 36721 11984 36735
rect 3207 36707 11998 36721
rect 3221 36693 12012 36707
rect 3235 36679 12026 36693
rect 3249 36665 12040 36679
rect 3263 36651 12054 36665
rect 3277 36637 12068 36651
rect 3291 36623 12082 36637
rect 3305 36609 12096 36623
rect 3319 36595 12110 36609
rect 3333 36581 12124 36595
rect 3347 36567 12138 36581
rect 3350 36564 12152 36567
rect 3361 36553 12194 36564
rect 3366 36548 12194 36553
rect 3380 36534 12194 36548
rect 3394 36520 12194 36534
rect 3408 36506 12194 36520
rect 3422 36492 12194 36506
rect 3436 36478 12194 36492
rect 3450 36464 12194 36478
rect 3464 36450 12194 36464
rect 3478 36436 12194 36450
rect 3492 36422 12194 36436
rect 3506 36408 12194 36422
rect 3520 36394 12194 36408
rect 3534 36380 12194 36394
rect 3548 36366 12194 36380
rect 3562 36352 12194 36366
rect 11648 34500 12194 36352
rect 3318 34259 11742 34500
rect 2880 32463 3333 34259
rect 2880 32439 11493 32463
rect 2882 32437 3305 32439
rect 2884 32435 3305 32437
rect 3557 32435 11517 32439
rect 2895 32424 11517 32435
rect 2909 32410 11517 32424
rect 2923 32396 11517 32410
rect 2937 32382 11521 32396
rect 2951 32368 11535 32382
rect 2965 32354 11549 32368
rect 2979 32340 11563 32354
rect 2993 32326 11577 32340
rect 3007 32312 11591 32326
rect 3021 32298 11605 32312
rect 3035 32284 11619 32298
rect 3049 32270 11633 32284
rect 3063 32256 11647 32270
rect 3077 32242 11661 32256
rect 3091 32228 11675 32242
rect 3105 32214 11689 32228
rect 3119 32200 11703 32214
rect 3133 32186 11717 32200
rect 3147 32172 11731 32186
rect 3161 32158 11745 32172
rect 3175 32144 11759 32158
rect 3189 32130 11773 32144
rect 3203 32116 11787 32130
rect 3217 32102 11801 32116
rect 3231 32088 11815 32102
rect 3245 32074 11829 32088
rect 3259 32060 11843 32074
rect 3273 32046 11857 32060
rect 3287 32032 11871 32046
rect 3301 32018 11885 32032
rect 3315 32004 11899 32018
rect 3329 31990 11913 32004
rect 3343 31976 11927 31990
rect 3357 31962 11941 31976
rect 3371 31948 11955 31962
rect 3385 31934 11969 31948
rect 3399 31920 11983 31934
rect 3413 31906 11997 31920
rect 3427 31892 12011 31906
rect 3441 31878 12025 31892
rect 3455 31864 12039 31878
rect 3469 31850 12053 31864
rect 3483 31836 12067 31850
rect 3497 31822 12081 31836
rect 3511 31808 12095 31822
rect 3525 31794 12109 31808
rect 3539 31780 12123 31794
rect 3553 31766 12137 31780
rect 3557 31762 12151 31766
rect 3567 31752 12194 31762
rect 11397 29900 12194 31752
rect 3319 29659 11726 29900
rect 3014 29354 3638 29659
rect 2880 27863 3333 29354
rect 2880 27857 11490 27863
rect 2891 27846 3305 27857
rect 2902 27835 3305 27846
rect 3578 27835 11496 27857
rect 2913 27824 11496 27835
rect 2927 27810 11496 27824
rect 2941 27796 11504 27810
rect 2955 27782 11518 27796
rect 2969 27768 11532 27782
rect 2983 27754 11546 27768
rect 2997 27740 11560 27754
rect 3011 27726 11574 27740
rect 3025 27712 11588 27726
rect 3039 27698 11602 27712
rect 3053 27684 11616 27698
rect 3067 27670 11630 27684
rect 3081 27656 11644 27670
rect 3095 27642 11658 27656
rect 3109 27628 11672 27642
rect 3123 27614 11686 27628
rect 3137 27600 11700 27614
rect 3151 27586 11714 27600
rect 3165 27572 11728 27586
rect 3179 27558 11742 27572
rect 3193 27544 11756 27558
rect 3207 27530 11770 27544
rect 3221 27516 11784 27530
rect 3235 27502 11798 27516
rect 3249 27488 11812 27502
rect 3263 27474 11826 27488
rect 3277 27460 11840 27474
rect 3291 27446 11854 27460
rect 3305 27432 11868 27446
rect 3319 27418 11882 27432
rect 3333 27404 11896 27418
rect 3347 27390 11910 27404
rect 3361 27376 11924 27390
rect 3375 27362 11938 27376
rect 3389 27348 11952 27362
rect 3403 27334 11966 27348
rect 3417 27320 11980 27334
rect 3431 27306 11994 27320
rect 3445 27292 12008 27306
rect 3459 27278 12022 27292
rect 3473 27264 12036 27278
rect 3487 27250 12050 27264
rect 3501 27236 12064 27250
rect 3515 27222 12078 27236
rect 3529 27208 12092 27222
rect 3543 27194 12106 27208
rect 3557 27180 12120 27194
rect 3571 27166 12134 27180
rect 3578 27159 12148 27166
rect 3585 27152 12194 27159
rect 11397 25300 12194 27152
rect 3333 25059 11740 25300
rect 2880 23263 4936 25059
rect 2880 23236 11483 23263
rect 2881 23235 11510 23236
rect 2892 23224 11510 23235
rect 2906 23210 11510 23224
rect 2920 23196 11510 23210
rect 2934 23182 11511 23196
rect 2948 23168 11525 23182
rect 2962 23154 11539 23168
rect 2976 23140 11553 23154
rect 2990 23126 11567 23140
rect 3004 23112 11581 23126
rect 3018 23098 11595 23112
rect 3032 23084 11609 23098
rect 3046 23070 11623 23084
rect 3060 23056 11637 23070
rect 3074 23042 11651 23056
rect 3088 23028 11665 23042
rect 3102 23014 11679 23028
rect 3116 23000 11693 23014
rect 3130 22986 11707 23000
rect 3144 22972 11721 22986
rect 3158 22958 11735 22972
rect 3172 22944 11749 22958
rect 3186 22930 11763 22944
rect 3200 22916 11777 22930
rect 3214 22902 11791 22916
rect 3228 22888 11805 22902
rect 3242 22874 11819 22888
rect 3256 22860 11833 22874
rect 3270 22846 11847 22860
rect 3284 22832 11861 22846
rect 3298 22818 11875 22832
rect 3312 22804 11889 22818
rect 3326 22790 11903 22804
rect 3340 22776 11917 22790
rect 3354 22762 11931 22776
rect 3368 22748 11945 22762
rect 3382 22734 11959 22748
rect 3396 22720 11973 22734
rect 3410 22706 11987 22720
rect 3424 22692 12001 22706
rect 3438 22678 12015 22692
rect 3452 22664 12029 22678
rect 3466 22650 12043 22664
rect 3480 22636 12057 22650
rect 3494 22622 12071 22636
rect 3508 22608 12085 22622
rect 3522 22594 12099 22608
rect 3536 22580 12113 22594
rect 3550 22566 12127 22580
rect 3564 22552 12141 22566
rect 11397 20700 12194 22552
rect 3314 20459 11740 20700
rect 2880 18663 4936 20459
rect 2880 18628 11501 18663
rect 2891 18617 11536 18628
rect 2905 18603 11536 18617
rect 2919 18589 11536 18603
rect 2933 18575 11536 18589
rect 2947 18561 11550 18575
rect 2961 18547 11564 18561
rect 2975 18533 11578 18547
rect 2989 18519 11592 18533
rect 3003 18505 11606 18519
rect 3017 18491 11620 18505
rect 3031 18477 11634 18491
rect 3045 18463 11648 18477
rect 3059 18449 11662 18463
rect 3073 18435 11676 18449
rect 3087 18421 11690 18435
rect 3101 18407 11704 18421
rect 3115 18393 11718 18407
rect 3129 18379 11732 18393
rect 3143 18365 11746 18379
rect 3157 18351 11760 18365
rect 3171 18337 11774 18351
rect 3185 18323 11788 18337
rect 3199 18309 11802 18323
rect 3213 18295 11816 18309
rect 3227 18281 11830 18295
rect 3241 18267 11844 18281
rect 3255 18253 11858 18267
rect 3269 18239 11872 18253
rect 3283 18225 11886 18239
rect 3297 18211 11900 18225
rect 3311 18197 11914 18211
rect 3325 18183 11928 18197
rect 3339 18169 11942 18183
rect 3353 18155 11956 18169
rect 3367 18141 11970 18155
rect 3381 18127 11984 18141
rect 3395 18113 11998 18127
rect 3409 18099 12012 18113
rect 3423 18085 12026 18099
rect 3437 18071 12040 18085
rect 3451 18057 12054 18071
rect 3465 18043 12068 18057
rect 3479 18029 12082 18043
rect 3493 18015 12096 18029
rect 3507 18001 12110 18015
rect 3521 17987 12124 18001
rect 3535 17973 12138 17987
rect 3538 17970 12152 17973
rect 3549 17959 12194 17970
rect 3550 17958 12194 17959
rect 3553 17955 12194 17958
rect 3556 17952 12194 17955
rect 11397 16100 12194 17952
rect 3314 15859 11740 16100
rect 2880 14911 4936 15859
rect 2880 14803 3654 14911
rect 2880 14756 4718 14803
rect 2880 14742 4726 14756
rect 2880 14728 4740 14742
rect 2880 14714 4754 14728
rect 2880 14700 4768 14714
rect 2880 14686 4782 14700
rect 2880 14672 4796 14686
rect 2880 14658 4810 14672
rect 2880 14644 4824 14658
rect 2880 14630 4838 14644
rect 2880 14616 4852 14630
rect 2880 14602 4866 14616
rect 2880 14588 4880 14602
rect 2880 14585 4894 14588
rect 2880 14063 4936 14585
rect 2880 14028 11489 14063
rect 2884 14024 11524 14028
rect 2898 14010 11524 14024
rect 2912 13996 11524 14010
rect 2926 13982 11524 13996
rect 2940 13968 11531 13982
rect 2954 13954 11545 13968
rect 2968 13940 11559 13954
rect 2982 13926 11573 13940
rect 2996 13912 11587 13926
rect 3010 13898 11601 13912
rect 3024 13884 11615 13898
rect 3038 13870 11629 13884
rect 3052 13856 11643 13870
rect 3066 13842 11657 13856
rect 3080 13828 11671 13842
rect 3094 13814 11685 13828
rect 3108 13800 11699 13814
rect 3122 13786 11713 13800
rect 3136 13772 11727 13786
rect 3150 13758 11741 13772
rect 3164 13744 11755 13758
rect 3178 13730 11769 13744
rect 3192 13716 11783 13730
rect 3206 13702 11797 13716
rect 3220 13688 11811 13702
rect 3234 13674 11825 13688
rect 3248 13660 11839 13674
rect 3262 13646 11853 13660
rect 3276 13632 11867 13646
rect 3290 13618 11881 13632
rect 3304 13604 11895 13618
rect 3318 13590 11909 13604
rect 3332 13576 11923 13590
rect 3346 13562 11937 13576
rect 3360 13548 11951 13562
rect 3374 13534 11965 13548
rect 3388 13520 11979 13534
rect 3402 13506 11993 13520
rect 3416 13492 12007 13506
rect 3430 13478 12021 13492
rect 3444 13464 12035 13478
rect 3458 13450 12049 13464
rect 3472 13436 12063 13450
rect 3486 13422 12077 13436
rect 3500 13408 12091 13422
rect 3514 13394 12105 13408
rect 3528 13380 12119 13394
rect 3542 13366 12133 13380
rect 3550 13358 12147 13366
rect 3556 13352 12194 13358
rect 11398 11500 12194 13352
rect 3319 11259 11734 11500
rect 3041 10981 3758 11259
rect 0 9388 146 9396
rect 0 9380 154 9388
rect 0 7394 162 9380
rect 2880 9463 3333 10981
rect 2880 9422 11483 9463
rect 2880 9408 11485 9422
rect 2880 9394 11499 9408
rect 2880 9380 11513 9394
rect 2880 9366 11527 9380
rect 2880 9352 11541 9366
rect 2880 9338 11555 9352
rect 2880 9324 11569 9338
rect 2880 9310 11583 9324
rect 2880 9296 11597 9310
rect 2880 9282 11611 9296
rect 2880 9268 11625 9282
rect 2880 9254 11639 9268
rect 2880 9240 11653 9254
rect 2880 9226 11667 9240
rect 2880 9212 11681 9226
rect 2880 9198 11695 9212
rect 2880 9184 11709 9198
rect 2880 9170 11723 9184
rect 2880 9156 11737 9170
rect 2880 9142 11751 9156
rect 2880 9128 11765 9142
rect 2880 9114 11779 9128
rect 2880 9100 11793 9114
rect 2880 9086 11807 9100
rect 2889 9077 11860 9086
rect 2903 9063 11860 9077
rect 2917 9049 11860 9063
rect 2931 9035 11860 9049
rect 2945 9021 11872 9035
rect 2959 9007 11886 9021
rect 2973 8993 11900 9007
rect 2987 8979 11914 8993
rect 3001 8965 11928 8979
rect 3015 8951 11942 8965
rect 3029 8937 11956 8951
rect 3043 8923 11970 8937
rect 3057 8909 11984 8923
rect 3071 8895 11998 8909
rect 3085 8881 12012 8895
rect 3099 8867 12026 8881
rect 3113 8853 12040 8867
rect 3127 8839 12054 8853
rect 3141 8825 12068 8839
rect 3155 8811 12082 8825
rect 3169 8797 12096 8811
rect 3183 8783 12110 8797
rect 3197 8769 12124 8783
rect 3211 8755 12138 8769
rect 3214 8752 12152 8755
rect 3225 8741 12194 8752
rect 3238 8728 12194 8741
rect 3252 8714 12194 8728
rect 3266 8700 12194 8714
rect 3280 8686 12194 8700
rect 3294 8672 12194 8686
rect 3308 8658 12194 8672
rect 3322 8644 12194 8658
rect 3336 8630 12194 8644
rect 3350 8616 12194 8630
rect 3364 8602 12194 8616
rect 3378 8588 12194 8602
rect 3392 8574 12194 8588
rect 3406 8560 12194 8574
rect 3420 8546 12194 8560
rect 3434 8532 12194 8546
rect 4570 8504 12194 8532
rect 10893 8502 12194 8504
rect 10907 8488 12194 8502
rect 10921 8474 12194 8488
rect 10935 8460 12194 8474
rect 10949 8446 12194 8460
rect 10963 8432 12194 8446
rect 10977 8418 12194 8432
rect 10991 8404 12194 8418
rect 11005 8390 12194 8404
rect 11019 8376 12194 8390
rect 11033 8362 12194 8376
rect 11047 8348 12194 8362
rect 11061 8334 12194 8348
rect 11075 8320 12194 8334
rect 11089 8306 12194 8320
rect 11103 8292 12194 8306
rect 11117 8278 12194 8292
rect 11131 8264 12194 8278
rect 11145 8250 12194 8264
rect 11159 8236 12194 8250
rect 11173 8222 12194 8236
rect 11187 8208 12194 8222
rect 11201 8194 12194 8208
rect 11215 8180 12194 8194
rect 11229 8166 12194 8180
rect 11243 8152 12194 8166
rect 11257 8138 12194 8152
rect 11271 8124 12194 8138
rect 11285 8110 12194 8124
rect 11299 8096 12194 8110
rect 11313 8082 12194 8096
rect 11327 8068 12194 8082
rect 11341 8054 12194 8068
rect 4080 8014 10503 8042
rect 11355 8040 12194 8054
rect 11369 8026 12194 8040
rect 3627 7964 10531 8014
rect 11383 8012 12194 8026
rect 11397 7998 12194 8012
rect 3627 7950 10542 7964
rect 3627 7936 10556 7950
rect 3627 7922 10570 7936
rect 3627 7908 10584 7922
rect 3627 7894 10598 7908
rect 3627 7880 10612 7894
rect 3627 7866 10626 7880
rect 3627 7852 10640 7866
rect 3627 7838 10654 7852
rect 3627 7824 10668 7838
rect 3627 7810 10682 7824
rect 3627 7796 10696 7810
rect 3627 7782 10710 7796
rect 3627 7768 10724 7782
rect 3627 7754 10738 7768
rect 3627 7740 10752 7754
rect 3627 7726 10766 7740
rect 3627 7712 10780 7726
rect 3627 7698 10794 7712
rect 3627 7684 10808 7698
rect 3627 7670 10822 7684
rect 3627 7656 10836 7670
rect 3627 7642 10850 7656
rect 3627 7639 10864 7642
rect 0 434 145 7394
rect 3182 7195 10906 7639
rect 11411 7195 12194 7998
rect 3097 5886 12194 7195
rect 3101 5882 11878 5886
rect 3115 5868 11878 5882
rect 3129 5854 11878 5868
rect 3143 5840 11878 5854
rect 3157 5826 11878 5840
rect 3171 5812 11878 5826
rect 3185 5798 11878 5812
rect 3199 5784 11878 5798
rect 3213 5770 11878 5784
rect 3227 5756 11878 5770
rect 3241 5742 11878 5756
rect 3255 5728 11878 5742
rect 3269 5714 11878 5728
rect 3283 5700 11878 5714
rect 3297 5686 11878 5700
rect 3311 5672 11878 5686
rect 3325 5658 11878 5672
rect 3339 5644 11878 5658
rect 3353 5630 11878 5644
rect 3367 5616 11878 5630
rect 3381 5602 11878 5616
rect 3395 5588 11878 5602
rect 3409 5574 11878 5588
rect 3423 5560 11878 5574
rect 3437 5546 11878 5560
rect 3451 5532 11878 5546
rect 3465 5518 11878 5532
rect 3479 5504 11878 5518
rect 3493 5490 11878 5504
rect 3507 5476 11878 5490
rect 3521 5462 11878 5476
rect 3535 5448 11878 5462
rect 3549 5434 11878 5448
rect 3563 5420 11878 5434
rect 3577 5406 11878 5420
rect 3591 5392 11878 5406
rect 3605 5378 11878 5392
rect 3619 5364 11878 5378
rect 3633 5350 11878 5364
rect 3647 5336 11878 5350
rect 3661 5322 11878 5336
rect 3675 5308 11878 5322
rect 3689 5294 11878 5308
rect 3703 5280 11878 5294
rect 3717 5266 11878 5280
rect 3731 5252 11878 5266
rect 3745 5238 11878 5252
rect 3759 5224 11878 5238
rect 3773 5210 11878 5224
rect 3787 5196 11878 5210
rect 7435 5160 11187 5196
rect 7435 2431 7550 5160
rect 7435 2424 9332 2431
rect 4953 2374 9339 2424
rect 4953 2360 9350 2374
rect 4953 2346 9364 2360
rect 4953 2332 9378 2346
rect 4953 2318 9392 2332
rect 4953 2304 9406 2318
rect 4953 2290 9420 2304
rect 4953 2276 9434 2290
rect 4953 2262 9448 2276
rect 4953 2248 9462 2262
rect 4953 2234 9476 2248
rect 4953 2220 9490 2234
rect 4953 2206 9504 2220
rect 4953 2192 9518 2206
rect 4953 2178 9532 2192
rect 4953 2164 9546 2178
rect 4953 2150 9560 2164
rect 4953 2136 9574 2150
rect 4953 2122 9588 2136
rect 4953 2108 9602 2122
rect 4953 2094 9616 2108
rect 4953 2080 9630 2094
rect 4953 2066 9644 2080
rect 4953 2052 9658 2066
rect 4953 2038 9672 2052
rect 4953 2024 9686 2038
rect 4953 2010 9700 2024
rect 4953 1996 9714 2010
rect 4953 1982 9728 1996
rect 4953 1968 9742 1982
rect 4953 1954 9756 1968
rect 4953 1940 9770 1954
rect 4953 1926 9784 1940
rect 4953 1912 9798 1926
rect 4953 1898 9812 1912
rect 4953 1884 9826 1898
rect 4953 1870 9840 1884
rect 4953 1856 9854 1870
rect 4953 1842 9868 1856
rect 4953 1828 9882 1842
rect 4953 1814 9896 1828
rect 4953 1800 9910 1814
rect 4953 1786 9924 1800
rect 4953 1772 9938 1786
rect 4953 1758 9952 1772
rect 4953 1744 9966 1758
rect 4953 1730 9980 1744
rect 4953 1716 9994 1730
rect 4953 1713 10008 1716
rect 0 0 43 434
rect 4935 135 10050 1713
rect 4935 0 5151 135
rect 5607 0 10050 135
rect 14886 0 15000 38031
<< metal3 >>
rect 632 37072 5002 40000
rect 640 37064 5002 37072
rect 670 37034 5002 37064
rect 700 37004 5002 37034
rect 730 36974 5002 37004
rect 760 36944 5002 36974
rect 790 36914 5002 36944
rect 820 36884 5002 36914
rect 850 36854 5002 36884
rect 880 36824 5002 36854
rect 910 36794 5002 36824
rect 940 36764 5002 36794
rect 970 36734 5002 36764
rect 1000 36704 5002 36734
rect 1030 36674 5002 36704
rect 1060 36644 5002 36674
rect 1090 36614 5002 36644
rect 1120 36584 5002 36614
rect 1150 36554 5002 36584
rect 1180 36524 5002 36554
rect 1210 36494 5002 36524
rect 1240 36464 5002 36494
rect 1270 36434 5002 36464
rect 1300 36404 5002 36434
rect 1330 36374 5002 36404
rect 1360 36344 5002 36374
rect 1390 36314 5002 36344
rect 1420 36284 5002 36314
rect 1450 36254 5002 36284
rect 1480 36224 5002 36254
rect 1510 36194 5002 36224
rect 1540 36164 5002 36194
rect 1570 36134 5002 36164
rect 1600 36104 5002 36134
rect 1630 36074 5002 36104
rect 1660 36044 5002 36074
rect 1690 36014 5002 36044
rect 1720 35984 5002 36014
rect 1750 35954 5002 35984
rect 1780 35924 5002 35954
rect 1810 35894 5002 35924
rect 1840 35864 5002 35894
rect 1870 35834 5002 35864
rect 1900 35804 5002 35834
rect 1930 35774 5002 35804
rect 1960 35744 5002 35774
rect 1990 35714 5002 35744
rect 2020 35684 5002 35714
rect 2050 35654 5002 35684
rect 2080 35624 5002 35654
rect 2110 35594 5002 35624
rect 2140 35564 5002 35594
rect 2170 35534 5002 35564
rect 2200 35504 5002 35534
rect 2230 35474 5002 35504
rect 2260 35444 5002 35474
rect 2290 35414 5002 35444
rect 2320 35384 5002 35414
rect 2350 35354 5002 35384
rect 2380 35324 5002 35354
rect 2410 35294 5002 35324
rect 2440 35264 5002 35294
rect 2470 35234 5002 35264
rect 2500 35204 5002 35234
rect 2530 35174 5002 35204
rect 2560 35144 5002 35174
rect 2590 35114 5002 35144
rect 2620 35084 5002 35114
rect 2650 35054 5002 35084
rect 2680 35024 5002 35054
rect 2710 34994 5002 35024
rect 2740 34964 5002 34994
rect 2770 34934 5002 34964
rect 2800 34904 5002 34934
rect 2830 34874 5002 34904
rect 2860 34844 5002 34874
rect 2890 34814 5002 34844
rect 2920 34784 5002 34814
rect 2950 34754 5002 34784
rect 2980 34724 5002 34754
rect 3010 34694 5002 34724
rect 3040 34664 5002 34694
rect 3070 34634 5002 34664
rect 3100 34528 5002 34634
rect 3100 34516 4990 34528
rect 3100 34495 4960 34516
rect 3100 33916 4380 34495
rect 3100 33886 4360 33916
rect 3100 33856 4330 33886
rect 3100 20920 4300 33856
rect 3100 20890 4316 20920
rect 3100 20860 4346 20890
rect 3100 20830 4376 20860
rect 3100 20800 4406 20830
rect 3100 20770 4436 20800
rect 3100 20740 4466 20770
rect 3100 20710 4496 20740
rect 3100 20680 4526 20710
rect 3100 20650 4556 20680
rect 3100 20620 4586 20650
rect 3100 20590 4616 20620
rect 3100 20560 4646 20590
rect 3100 20530 4676 20560
rect 3100 20500 4706 20530
rect 3100 20470 4736 20500
rect 5186 35070 7364 40000
rect 5186 35052 7346 35070
rect 5186 35037 7316 35052
rect 7593 35070 9771 38004
rect 7611 35052 9771 35070
rect 7641 35037 9771 35052
rect 5186 34182 6466 35037
rect 5186 34152 6446 34182
rect 5186 34122 6416 34152
rect 5186 20958 6386 34122
rect 8491 34182 9771 35037
rect 8511 34152 9771 34182
rect 8541 34122 9771 34152
rect 8571 22110 9771 34122
rect 8557 22080 9771 22110
rect 8527 22050 9771 22080
rect 8497 22020 9771 22050
rect 8491 21630 9771 22020
rect 9955 37072 14325 38008
rect 9955 37064 14317 37072
rect 9955 37039 14287 37064
rect 9955 34844 12090 37039
rect 9955 34814 12067 34844
rect 9955 34784 12037 34814
rect 9955 34754 12007 34784
rect 9955 34724 11977 34754
rect 9955 34694 11937 34724
rect 9955 34664 11917 34694
rect 9955 34634 11887 34664
rect 9955 34529 11857 34634
rect 9967 34517 11857 34529
rect 9997 34487 11857 34517
rect 10027 34457 11857 34487
rect 10057 34427 11857 34457
rect 10087 34397 11857 34427
rect 10117 34367 11857 34397
rect 10147 34337 11857 34367
rect 10177 34307 11857 34337
rect 10207 34277 11857 34307
rect 10237 34247 11857 34277
rect 10267 34217 11857 34247
rect 10297 34187 11857 34217
rect 10327 34157 11857 34187
rect 10357 34127 11857 34157
rect 10387 34097 11857 34127
rect 10417 34067 11857 34097
rect 10447 34037 11857 34067
rect 10477 34007 11857 34037
rect 10507 33977 11857 34007
rect 10537 33947 11857 33977
rect 10567 33917 11857 33947
rect 10597 33887 11857 33917
rect 10627 33857 11857 33887
rect 8491 21611 9752 21630
rect 8491 21597 9722 21611
rect 10657 22072 11857 33857
rect 10641 22042 11857 22072
rect 10611 22012 11857 22042
rect 10581 21982 11857 22012
rect 10577 21597 11857 21982
rect 8491 21164 8770 21597
rect 5186 20928 6400 20958
rect 5186 20898 6430 20928
rect 5186 20868 6460 20898
rect 5186 20478 6466 20868
rect 3100 20440 4766 20470
rect 5205 20459 6466 20478
rect 3129 20411 4796 20440
rect 5235 20429 6466 20459
rect 3159 20381 4825 20411
rect 5265 20399 6466 20429
rect 3189 20351 4855 20381
rect 5295 20369 6466 20399
rect 3219 20321 4885 20351
rect 5325 20339 6466 20369
rect 3249 20291 4915 20321
rect 5355 20309 6466 20339
rect 3279 20261 4945 20291
rect 5385 20279 6466 20309
rect 3309 20231 4975 20261
rect 5415 20249 6466 20279
rect 3339 20201 5005 20231
rect 5445 20219 6466 20249
rect 3369 20171 5035 20201
rect 5475 20189 6466 20219
rect 3399 20141 5065 20171
rect 5505 20159 6466 20189
rect 3429 20111 5095 20141
rect 5535 20129 6466 20159
rect 3459 20081 5125 20111
rect 5565 20099 6466 20129
rect 3489 20051 5155 20081
rect 5595 20069 6466 20099
rect 3519 20021 5185 20051
rect 5625 20039 6466 20069
rect 3549 19991 5215 20021
rect 5655 20009 6466 20039
rect 3579 19961 5245 19991
rect 5685 19979 6466 20009
rect 5699 19973 6466 19979
rect 7638 21161 8770 21164
rect 7608 21131 8770 21161
rect 5699 19965 7379 19973
rect 3609 19931 5275 19961
rect 5729 19935 7379 19965
rect 3639 19901 5305 19931
rect 5759 19905 7379 19935
rect 3669 19871 5335 19901
rect 5789 19875 7379 19905
rect 3699 19841 5365 19871
rect 5819 19845 7379 19875
rect 3729 19811 5395 19841
rect 5849 19815 7379 19845
rect 3759 19781 5425 19811
rect 5879 19785 7379 19815
rect 3789 19751 5455 19781
rect 5909 19755 7379 19785
rect 3819 19721 5485 19751
rect 5939 19725 7379 19755
rect 3849 19691 5515 19721
rect 5969 19695 7379 19725
rect 3879 19661 5545 19691
rect 5999 19665 7379 19695
rect 3909 19631 5575 19661
rect 6029 19635 7379 19665
rect 3939 19601 5605 19631
rect 6059 19605 7379 19635
rect 3969 19571 5635 19601
rect 6089 19575 7379 19605
rect 3999 19541 5665 19571
rect 6119 19545 7379 19575
rect 4029 19511 5695 19541
rect 6149 19515 7379 19545
rect 4059 19481 5725 19511
rect 6179 19485 7379 19515
rect 4089 19451 5755 19481
rect 6209 19455 7379 19485
rect 4119 19421 5785 19451
rect 6239 19425 7379 19455
rect 4149 19391 5815 19421
rect 6269 19395 7379 19425
rect 4179 19361 5845 19391
rect 6299 19365 7379 19395
rect 4209 19331 5875 19361
rect 6329 19335 7379 19365
rect 4239 19301 5905 19331
rect 4269 19271 5905 19301
rect 4299 19241 5905 19271
rect 4329 19211 5905 19241
rect 4359 19181 5905 19211
rect 4389 19151 5905 19181
rect 4419 19121 5905 19151
rect 4449 19091 5905 19121
rect 4479 19061 5905 19091
rect 4509 19031 5905 19061
rect 4539 19001 5905 19031
rect 4569 18971 5905 19001
rect 4599 18941 5905 18971
rect 4629 18911 5905 18941
rect 4659 18881 5905 18911
rect 4689 18851 5905 18881
rect 4719 18821 5905 18851
rect 4749 18598 5905 18821
rect 6359 19305 7379 19335
rect 4749 18568 5927 18598
rect 6389 18598 7379 19305
rect 4749 18538 5957 18568
rect 6367 18568 7379 18598
rect 6337 18538 7379 18568
rect 4749 18508 5987 18538
rect 6307 18508 7379 18538
rect 4764 18493 6017 18508
rect 4779 18478 6032 18493
rect 6277 18478 7379 18508
rect 4789 18468 7379 18478
rect 4819 18438 7379 18468
rect 4849 18408 7379 18438
rect 4879 18378 7379 18408
rect 4909 18348 7379 18378
rect 4939 18318 7379 18348
rect 4969 18288 7379 18318
rect 4999 18258 7379 18288
rect 5029 18228 7379 18258
rect 5059 18198 7379 18228
rect 5089 18168 7379 18198
rect 5119 18138 7379 18168
rect 5149 18108 7379 18138
rect 99 0 4879 7302
rect 5179 0 7379 18108
rect 7578 20637 8770 21131
rect 7578 20607 8748 20637
rect 7578 20577 8718 20607
rect 7578 20547 8688 20577
rect 7578 20517 8658 20547
rect 7578 20487 8628 20517
rect 10191 21592 11857 21597
rect 10161 21563 11828 21592
rect 10132 21559 11798 21563
rect 10132 21533 10662 21559
rect 10102 21503 10662 21533
rect 10072 21473 10662 21503
rect 10053 20516 10662 21473
rect 7578 20457 8598 20487
rect 7578 20021 8568 20457
rect 9112 20513 10662 20516
rect 9082 20483 10662 20513
rect 7578 19991 8590 20021
rect 9052 20403 10662 20483
rect 9052 20373 10638 20403
rect 9052 20343 10608 20373
rect 9052 20313 10578 20343
rect 9052 20284 10548 20313
rect 9052 20033 10288 20284
rect 7578 19961 8620 19991
rect 9042 20003 10268 20033
rect 9012 19973 10238 20003
rect 7578 19931 8650 19961
rect 8982 19943 10208 19973
rect 7578 19901 8680 19931
rect 8952 19922 10208 19943
rect 8931 19901 10208 19922
rect 7578 19660 10208 19901
rect 7578 19650 10198 19660
rect 7578 19627 10168 19650
rect 7578 19320 9858 19627
rect 7578 19290 9838 19320
rect 7578 19260 9808 19290
rect 7578 0 9778 19260
rect 10078 0 14858 10000
<< obsm3 >>
rect 0 37021 552 40000
rect 0 36991 570 37021
rect 0 36961 600 36991
rect 0 36931 630 36961
rect 0 36901 660 36931
rect 0 36871 690 36901
rect 0 36841 720 36871
rect 0 36811 750 36841
rect 0 36781 780 36811
rect 0 36751 810 36781
rect 0 36721 840 36751
rect 0 36691 870 36721
rect 0 36661 900 36691
rect 0 36631 930 36661
rect 0 36601 960 36631
rect 0 36571 990 36601
rect 0 36541 1020 36571
rect 0 36511 1050 36541
rect 0 36481 1080 36511
rect 0 36451 1110 36481
rect 0 36421 1140 36451
rect 0 36391 1170 36421
rect 0 36361 1200 36391
rect 0 36331 1230 36361
rect 0 36301 1260 36331
rect 0 36271 1290 36301
rect 0 36241 1320 36271
rect 0 36211 1350 36241
rect 0 36181 1380 36211
rect 0 36151 1410 36181
rect 0 36121 1440 36151
rect 0 36091 1470 36121
rect 0 36061 1500 36091
rect 0 36031 1530 36061
rect 0 36001 1560 36031
rect 0 35971 1590 36001
rect 0 35941 1620 35971
rect 0 35911 1650 35941
rect 0 35881 1680 35911
rect 0 35851 1710 35881
rect 0 35821 1740 35851
rect 0 35791 1770 35821
rect 0 35761 1800 35791
rect 0 35731 1830 35761
rect 0 35701 1860 35731
rect 0 35671 1890 35701
rect 0 35641 1920 35671
rect 0 35611 1950 35641
rect 0 35581 1980 35611
rect 0 35551 2010 35581
rect 0 35521 2040 35551
rect 0 35491 2070 35521
rect 0 35461 2100 35491
rect 0 35431 2130 35461
rect 0 35401 2160 35431
rect 0 35371 2190 35401
rect 0 35341 2220 35371
rect 0 35311 2250 35341
rect 0 35281 2280 35311
rect 0 35251 2310 35281
rect 0 35221 2340 35251
rect 0 35191 2370 35221
rect 0 35161 2400 35191
rect 0 35131 2430 35161
rect 0 35101 2460 35131
rect 0 35071 2490 35101
rect 0 35041 2520 35071
rect 0 35011 2550 35041
rect 0 34981 2580 35011
rect 0 34951 2610 34981
rect 0 34921 2640 34951
rect 0 34891 2670 34921
rect 0 34861 2700 34891
rect 0 34831 2730 34861
rect 0 34801 2760 34831
rect 0 34771 2790 34801
rect 0 34741 2820 34771
rect 0 34711 2850 34741
rect 0 34691 552 34711
rect 2780 34691 2880 34711
rect 0 9326 39 34691
rect 2760 34661 2900 34691
rect 2760 34631 2930 34661
rect 2760 34601 2960 34631
rect 2760 34571 2990 34601
rect 2760 20402 3020 34571
rect 5082 34495 5106 40000
rect 4380 20969 5106 34495
rect 4394 20955 5106 20969
rect 4424 20925 5106 20955
rect 4454 20895 5106 20925
rect 4484 20865 5106 20895
rect 4514 20835 5106 20865
rect 4544 20805 5106 20835
rect 4574 20775 5106 20805
rect 4604 20745 5106 20775
rect 4634 20715 5106 20745
rect 4664 20685 5106 20715
rect 4694 20655 5106 20685
rect 4724 20625 5106 20655
rect 4754 20595 5106 20625
rect 4784 20565 5106 20595
rect 4814 20535 5106 20565
rect 4844 20505 5106 20535
rect 4874 20475 5106 20505
rect 7444 38088 15000 40000
rect 7444 38084 9875 38088
rect 7444 35037 7513 38084
rect 6466 21164 8491 35037
rect 9851 34484 9875 38084
rect 14405 37039 15000 38088
rect 12090 34724 15000 37039
rect 9851 34454 9887 34484
rect 9851 34424 9917 34454
rect 9851 34394 9947 34424
rect 9851 34364 9977 34394
rect 9851 34334 10007 34364
rect 9851 34304 10037 34334
rect 9851 34274 10067 34304
rect 9851 34244 10097 34274
rect 9851 34214 10127 34244
rect 9851 34184 10157 34214
rect 9851 34154 10187 34184
rect 9851 34124 10217 34154
rect 9851 34094 10247 34124
rect 9851 34064 10277 34094
rect 9851 34034 10307 34064
rect 9851 34004 10337 34034
rect 9851 33974 10367 34004
rect 9851 33944 10397 33974
rect 9851 33914 10427 33944
rect 9851 33884 10457 33914
rect 9851 33854 10487 33884
rect 9851 33824 10517 33854
rect 9851 33794 10547 33824
rect 9851 21597 10577 33794
rect 4904 20445 5106 20475
rect 4905 20444 5106 20445
rect 4935 20414 5107 20444
rect 2760 20372 3025 20402
rect 4965 20384 5137 20414
rect 2760 20342 3055 20372
rect 4995 20354 5167 20384
rect 2760 20312 3085 20342
rect 5025 20324 5197 20354
rect 2760 20304 3115 20312
rect 2804 20288 3115 20304
rect 5055 20294 5227 20324
rect 2834 20258 3139 20288
rect 5085 20264 5257 20294
rect 2864 20228 3169 20258
rect 5115 20234 5287 20264
rect 2894 20198 3199 20228
rect 5145 20204 5317 20234
rect 2924 20168 3229 20198
rect 5175 20174 5347 20204
rect 2954 20138 3259 20168
rect 5205 20144 5377 20174
rect 2984 20108 3289 20138
rect 5235 20114 5407 20144
rect 3014 20078 3319 20108
rect 5265 20084 5437 20114
rect 3044 20048 3349 20078
rect 5295 20054 5467 20084
rect 3074 20018 3379 20048
rect 5325 20024 5497 20054
rect 3104 19988 3409 20018
rect 5355 19994 5527 20024
rect 3134 19958 3439 19988
rect 5385 19964 5557 19994
rect 6466 19973 7498 21164
rect 3164 19928 3469 19958
rect 5415 19934 5587 19964
rect 3194 19898 3499 19928
rect 5445 19904 5617 19934
rect 3224 19868 3529 19898
rect 5475 19874 5647 19904
rect 3254 19838 3559 19868
rect 5505 19844 5677 19874
rect 3284 19808 3589 19838
rect 5535 19814 5707 19844
rect 3314 19778 3619 19808
rect 5565 19784 5737 19814
rect 3344 19748 3649 19778
rect 5595 19754 5767 19784
rect 3374 19718 3679 19748
rect 5625 19724 5797 19754
rect 3404 19688 3709 19718
rect 5655 19694 5827 19724
rect 3434 19658 3739 19688
rect 5685 19664 5857 19694
rect 3464 19628 3769 19658
rect 5715 19634 5887 19664
rect 3494 19598 3799 19628
rect 5745 19604 5917 19634
rect 3524 19568 3829 19598
rect 5775 19574 5947 19604
rect 3554 19538 3859 19568
rect 5805 19544 5977 19574
rect 3584 19508 3889 19538
rect 5835 19514 6007 19544
rect 3614 19478 3919 19508
rect 5865 19484 6037 19514
rect 3644 19448 3949 19478
rect 5895 19454 6067 19484
rect 3674 19418 3979 19448
rect 5925 19424 6097 19454
rect 3704 19388 4009 19418
rect 5955 19394 6127 19424
rect 3734 19358 4039 19388
rect 5985 19364 6157 19394
rect 5985 19362 6187 19364
rect 3764 19328 4069 19358
rect 5985 19332 6189 19362
rect 3794 19298 4099 19328
rect 3824 19268 4129 19298
rect 3854 19238 4159 19268
rect 3884 19208 4189 19238
rect 3914 19178 4219 19208
rect 3944 19148 4249 19178
rect 3974 19118 4279 19148
rect 4004 19088 4309 19118
rect 4034 19058 4339 19088
rect 4064 19028 4369 19058
rect 4094 18998 4399 19028
rect 4124 18968 4429 18998
rect 4154 18938 4459 18968
rect 4184 18908 4489 18938
rect 4214 18878 4519 18908
rect 4244 18848 4549 18878
rect 4274 18818 4579 18848
rect 4304 18788 4609 18818
rect 4334 18758 4639 18788
rect 4339 18753 4669 18758
rect 4369 18723 4669 18753
rect 4399 18693 4669 18723
rect 4429 18663 4669 18693
rect 4459 18633 4669 18663
rect 4489 18603 4669 18633
rect 4519 18573 4669 18603
rect 4549 18543 4669 18573
rect 4579 18513 4669 18543
rect 4589 18475 4669 18513
rect 5985 19302 6219 19332
rect 5985 19272 6249 19302
rect 5985 19242 6279 19272
rect 5985 18653 6309 19242
rect 5990 18648 6309 18653
rect 6020 18618 6309 18648
rect 6050 18588 6309 18618
rect 6080 18558 6309 18588
rect 4639 18453 4669 18475
rect 4959 18135 4979 18165
rect 4959 18125 5009 18135
rect 4939 18105 5019 18125
rect 4939 18075 5039 18105
rect 4939 18045 5069 18075
rect 0 9296 52 9326
rect 0 9266 82 9296
rect 0 9244 112 9266
rect 0 7327 162 9244
rect 0 0 39 7327
rect 4939 0 5099 18045
rect 7459 0 7498 19973
rect 8770 20516 10053 21597
rect 11937 21559 12240 34724
rect 8648 20076 8972 20516
rect 8653 20071 8972 20076
rect 8683 20041 8972 20071
rect 8713 20011 8972 20041
rect 10662 20284 12240 21559
rect 8743 19981 8972 20011
rect 10288 19910 12240 20284
rect 10288 19627 11866 19910
rect 9858 19197 11583 19627
rect 9858 18062 11153 19197
rect 9858 0 10018 18062
rect 14918 0 15000 34724
<< metal4 >>
rect 0 35157 15000 40000
rect 0 14007 15000 19000
rect 0 12817 15000 13707
rect 0 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 15000 9247
rect 0 7347 15000 8037
rect 0 6377 15000 7067
rect 0 5167 15000 6097
rect 0 3957 15000 4887
rect 0 2987 15000 3677
rect 0 1777 15000 2707
rect 0 407 15000 1497
<< obsm4 >>
rect 2266 34590 12734 34620
rect 2236 34560 12764 34590
rect 2206 34530 12794 34560
rect 2176 34500 12824 34530
rect 2146 34473 12854 34500
rect 2122 34470 12876 34473
rect 2116 34440 12884 34470
rect 2086 34410 12914 34440
rect 2056 34380 12944 34410
rect 2026 34350 12974 34380
rect 1996 34320 13004 34350
rect 1966 34290 13034 34320
rect 1936 34260 13064 34290
rect 1906 34230 13094 34260
rect 1876 34215 13124 34230
rect 1864 34200 13134 34215
rect 1846 34170 13154 34200
rect 1816 34140 13184 34170
rect 1786 34110 13214 34140
rect 1756 34080 13244 34110
rect 1726 34064 2474 34080
rect 12526 34064 13274 34080
rect 1710 34034 2444 34064
rect 12556 34034 13290 34064
rect 1680 34004 2414 34034
rect 12586 34004 13320 34034
rect 1650 33974 2384 34004
rect 12616 33974 13350 34004
rect 1620 33944 2354 33974
rect 12646 33944 13380 33974
rect 1590 33918 2324 33944
rect 1575 33914 2324 33918
rect 12676 33918 13410 33944
rect 12676 33914 13423 33918
rect 1560 33911 2303 33914
rect 12695 33911 13440 33914
rect 1560 33884 2294 33911
rect 12706 33884 13440 33911
rect 1530 33854 2264 33884
rect 12736 33854 13470 33884
rect 1500 33824 2234 33854
rect 12766 33824 13500 33854
rect 1470 33794 2204 33824
rect 12796 33794 13530 33824
rect 1440 33764 2174 33794
rect 12826 33764 13560 33794
rect 1410 33734 2144 33764
rect 12856 33734 13590 33764
rect 1380 33704 2114 33734
rect 12886 33704 13620 33734
rect 1350 33674 2084 33704
rect 12916 33674 13650 33704
rect 1320 33644 2054 33674
rect 12946 33644 13680 33674
rect 1290 33614 2024 33644
rect 12976 33614 13710 33644
rect 1260 33590 1994 33614
rect 1247 33584 1994 33590
rect 13006 33590 13740 33614
rect 13006 33584 13751 33590
rect 1230 33554 1964 33584
rect 13036 33554 13770 33584
rect 1200 33524 1934 33554
rect 13066 33524 13800 33554
rect 1170 33494 1904 33524
rect 13096 33494 13830 33524
rect 1140 33464 1874 33494
rect 13126 33464 13860 33494
rect 1110 33435 1844 33464
rect 1094 33434 1844 33435
rect 13156 33435 13890 33464
rect 13156 33434 13904 33435
rect 1080 33404 1814 33434
rect 13186 33404 13920 33434
rect 1050 33374 1784 33404
rect 13216 33374 13950 33404
rect 1020 33344 1754 33374
rect 13246 33344 13980 33374
rect 990 33314 1724 33344
rect 13276 33314 14010 33344
rect 960 33300 1710 33314
rect 13290 33300 14006 33314
rect 960 33270 1680 33300
rect 13320 33270 13934 33300
rect 14006 33270 14040 33300
rect 960 33240 1650 33270
rect 13350 33240 13904 33270
rect 13934 33240 14040 33270
rect 960 33210 1620 33240
rect 13380 33210 14040 33240
rect 960 33180 1590 33210
rect 13410 33180 14040 33210
rect 960 33150 1560 33180
rect 13440 33150 14040 33180
rect 960 33120 1530 33150
rect 13470 33135 14040 33150
rect 13470 33120 13572 33135
rect 13645 33120 14040 33135
rect 960 21070 1500 33120
rect 13572 33109 14040 33120
rect 13506 33090 14040 33109
rect 960 21056 1492 21070
rect 13500 21056 14040 33090
rect 960 21026 1514 21056
rect 13486 21026 14040 21056
rect 960 20996 1544 21026
rect 13456 20996 14040 21026
rect 960 20971 1574 20996
rect 13426 20971 14040 20996
rect 960 20966 1587 20971
rect 13411 20966 14040 20971
rect 960 20936 1604 20966
rect 13396 20936 14040 20966
rect 960 20906 1634 20936
rect 13366 20906 14040 20936
rect 960 20876 1664 20906
rect 13336 20876 14040 20906
rect 968 20853 1694 20876
rect 1032 20846 1694 20853
rect 13306 20846 14040 20876
rect 976 20830 1724 20846
rect 13276 20830 14024 20846
rect 1006 20800 1740 20830
rect 13260 20800 13994 20830
rect 1036 20770 1770 20800
rect 13230 20770 13964 20800
rect 1066 20740 1800 20770
rect 13200 20740 13934 20770
rect 1096 20710 1830 20740
rect 13170 20718 13907 20740
rect 13170 20710 13904 20718
rect 1126 20680 1860 20710
rect 13140 20680 13874 20710
rect 1156 20650 1890 20680
rect 13110 20650 13844 20680
rect 1186 20620 1920 20650
rect 13080 20646 13834 20650
rect 13080 20620 13814 20646
rect 1216 20590 1950 20620
rect 13050 20590 13784 20620
rect 1246 20560 1980 20590
rect 13020 20560 13754 20590
rect 1276 20530 2010 20560
rect 12990 20530 13724 20560
rect 1302 20526 2040 20530
rect 1306 20506 2040 20526
rect 12960 20526 13696 20530
rect 12960 20506 13694 20526
rect 1306 20500 2047 20506
rect 12951 20500 13694 20506
rect 1336 20470 2070 20500
rect 12930 20470 13664 20500
rect 1366 20440 2100 20470
rect 12900 20440 13634 20470
rect 1396 20410 2130 20440
rect 12870 20410 13604 20440
rect 1426 20380 2160 20410
rect 12840 20380 13574 20410
rect 1455 20371 2190 20380
rect 1456 20350 2190 20371
rect 12810 20350 13544 20380
rect 1486 20320 2220 20350
rect 12780 20320 13514 20350
rect 1516 20290 2250 20320
rect 12750 20290 13484 20320
rect 1546 20260 2280 20290
rect 12720 20260 13454 20290
rect 1576 20230 2310 20260
rect 12690 20230 13424 20260
rect 1606 20200 2340 20230
rect 12660 20200 13394 20230
rect 1636 20182 2370 20200
rect 12630 20182 13364 20200
rect 1636 20170 2371 20182
rect 12627 20170 13364 20182
rect 1666 20140 2400 20170
rect 12600 20140 13334 20170
rect 1696 20110 2430 20140
rect 12570 20110 13304 20140
rect 1726 20080 2460 20110
rect 12540 20080 13274 20110
rect 1756 20070 12510 20080
rect 12522 20070 13244 20080
rect 1756 20050 13244 20070
rect 1783 20043 13215 20050
rect 1786 20020 13214 20043
rect 1816 19990 13184 20020
rect 1846 19960 12552 19990
rect 12560 19960 13154 19990
rect 1876 19930 12560 19960
rect 12572 19930 13124 19960
rect 1906 19900 12572 19930
rect 12585 19900 13094 19930
rect 1936 19870 12585 19900
rect 12597 19870 13064 19900
rect 1966 19845 12597 19870
rect 12610 19845 13034 19870
rect 1966 19840 13034 19845
rect 1996 19810 13004 19840
rect 2026 19780 12974 19810
rect 2056 19750 12944 19780
rect 2086 19720 12914 19750
rect 2116 19690 12884 19720
rect 2146 19660 12854 19690
rect 2176 19630 12824 19660
rect 2206 19600 12794 19630
rect 2236 19570 12715 19600
rect 12722 19570 12764 19600
rect 2266 19540 12722 19570
<< metal5 >>
rect 0 35157 15000 40000
rect 2266 34594 12734 34620
rect 2240 34514 12760 34594
rect 2160 34434 12840 34514
rect 2080 34354 12920 34434
rect 2000 34274 13000 34354
rect 1920 34194 13080 34274
rect 1840 34114 13160 34194
rect 1760 34034 13240 34114
rect 1680 33954 13320 34034
rect 1600 33874 13400 33954
rect 1520 33794 13480 33874
rect 1440 33714 13560 33794
rect 1360 33634 13640 33714
rect 1280 33554 13720 33634
rect 1200 33474 13800 33554
rect 1120 33394 13880 33474
rect 1040 33314 13960 33394
rect 960 20846 14040 33314
rect 986 20820 14014 20846
rect 1066 20740 13934 20820
rect 1146 20660 13854 20740
rect 1226 20580 13774 20660
rect 1306 20500 13694 20580
rect 1386 20420 13614 20500
rect 1466 20340 13534 20420
rect 1546 20260 13454 20340
rect 1626 20180 13374 20260
rect 1706 20100 13294 20180
rect 1786 20020 13214 20100
rect 1866 19940 13134 20020
rect 1946 19860 13054 19940
rect 2026 19780 12974 19860
rect 2106 19700 12894 19780
rect 2186 19620 12814 19700
rect 2266 19540 12734 19620
rect 0 14007 15000 18997
rect 0 12837 15000 13687
rect 0 11667 15000 12517
rect 0 9547 15000 11347
rect 0 8337 15000 9227
rect 0 7367 15000 8017
rect 0 6397 15000 7047
rect 0 5187 15000 6077
rect 0 3977 15000 4867
rect 0 3007 15000 3657
rect 0 1797 15000 2687
rect 0 427 15000 1477
<< labels >>
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 2266 34594 12734 34620 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2266 19540 12734 19620 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2240 34514 12760 34594 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2186 19620 12814 19700 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2160 34434 12840 34514 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2106 19700 12894 19780 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2080 34354 12920 34434 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2026 19780 12974 19860 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 2000 34274 13000 34354 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1946 19860 13054 19940 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1920 34194 13080 34274 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1866 19940 13134 20020 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1840 34114 13160 34194 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1786 20020 13214 20100 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1760 34034 13240 34114 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1706 20100 13294 20180 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1680 33954 13320 34034 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1626 20180 13374 20260 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1600 33874 13400 33954 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1546 20260 13454 20340 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1520 33794 13480 33874 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1466 20340 13534 20420 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1440 33714 13560 33794 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1386 20420 13614 20500 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1360 33634 13640 33714 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1306 20500 13694 20580 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1280 33554 13720 33634 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1226 20580 13774 20660 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1200 33474 13800 33554 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1146 20660 13854 20740 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1120 33394 13880 33474 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1066 20740 13934 20820 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 1040 33314 13960 33394 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 986 20820 14014 20846 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal5 s 960 20846 14040 33314 6 P_PAD
port 3 nsew signal bidirectional
rlabel metal2 s 12222 36576 14858 36590 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 34940 14858 36576 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 34931 14858 34940 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 31774 14858 31788 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 30356 14858 31774 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 30345 14858 30356 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 27171 14858 27185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 25742 14858 27171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 25731 14858 25742 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 22564 14858 22578 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 21142 14858 22564 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 21131 14858 21142 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 17982 14858 17996 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 16542 14858 17982 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 16531 14858 16542 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 13370 14858 13384 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 11948 14858 13370 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 11945 14858 11948 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 8764 14858 8778 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 6191 14858 8764 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12222 6182 14858 6191 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12219 11931 14858 11945 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12213 34917 14858 34931 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12213 6168 14858 6182 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12211 30331 14858 30345 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12211 25717 14858 25731 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12211 21117 14858 21131 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12211 16517 14858 16531 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 36590 14858 36604 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 31788 14858 31802 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 27185 14858 27199 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 22578 14858 22592 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 17996 14858 18010 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 13384 14858 13398 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12208 8778 14858 8792 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12205 11917 14858 11931 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12199 34903 14858 34917 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12199 6154 14858 6168 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12197 30317 14858 30331 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12197 25703 14858 25717 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12197 21103 14858 21117 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12197 16503 14858 16517 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 36604 14858 36618 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 31802 14858 31816 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 27199 14858 27213 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 22592 14858 22606 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 18010 14858 18024 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 13398 14858 13412 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12194 8792 14858 8806 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12191 11903 14858 11917 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12185 34889 14858 34903 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12185 6140 14858 6154 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12183 30303 14858 30317 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12183 25689 14858 25703 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12183 21089 14858 21103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12183 16489 14858 16503 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 36618 14858 36632 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 31816 14858 31830 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 27213 14858 27227 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 22606 14858 22620 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 18024 14858 18038 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 13412 14858 13426 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12180 8806 14858 8820 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12177 11889 14858 11903 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12171 34875 14858 34889 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12171 6126 14858 6140 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12169 30289 14858 30303 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12169 25675 14858 25689 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12169 21075 14858 21089 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12169 16475 14858 16489 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 36632 14858 36646 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 31830 14858 31844 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 27227 14858 27241 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 22620 14858 22634 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 18038 14858 18052 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 13426 14858 13440 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12166 8820 14858 8834 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12163 11875 14858 11889 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12157 34861 14858 34875 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12157 6112 14858 6126 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12155 30275 14858 30289 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12155 25661 14858 25675 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12155 21061 14858 21075 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12155 16461 14858 16475 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 36646 14858 36660 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 31844 14858 31858 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 27241 14858 27255 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 22634 14858 22648 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 18052 14858 18066 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 13440 14858 13454 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12152 8834 14858 8848 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12149 11861 14858 11875 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12143 34847 14858 34861 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12143 6098 14858 6112 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12141 30261 14858 30275 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12141 25647 14858 25661 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12141 21047 14858 21061 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12141 16447 14858 16461 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 36660 14858 36674 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 31858 14858 31872 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 27255 14858 27269 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 22648 14858 22662 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 18066 14858 18080 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 13454 14858 13468 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12138 8848 14858 8862 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12135 11847 14858 11861 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12129 34833 14858 34847 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12129 6084 14858 6098 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12127 30247 14858 30261 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12127 25633 14858 25647 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12127 21033 14858 21047 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12127 16433 14858 16447 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 36674 14858 36688 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 31872 14858 31886 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 27269 14858 27283 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 22662 14858 22676 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 18080 14858 18094 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 13468 14858 13482 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12124 8862 14858 8876 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12121 11833 14858 11847 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12115 34819 14858 34833 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12115 6070 14858 6084 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12113 30233 14858 30247 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12113 25619 14858 25633 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12113 21019 14858 21033 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12113 16419 14858 16433 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 36688 14858 36702 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 31886 14858 31900 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 27283 14858 27297 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 22676 14858 22690 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 18094 14858 18108 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 13482 14858 13496 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12110 8876 14858 8890 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12107 11819 14858 11833 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12101 34805 14858 34819 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12101 6056 14858 6070 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12099 30219 14858 30233 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12099 25605 14858 25619 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12099 21005 14858 21019 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12099 16405 14858 16419 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 36702 14858 36716 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 31900 14858 31914 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 27297 14858 27311 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 22690 14858 22704 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 18108 14858 18122 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 13496 14858 13510 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12096 8890 14858 8904 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12093 11805 14858 11819 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12087 34791 14858 34805 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12087 6042 14858 6056 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12085 30205 14858 30219 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12085 25591 14858 25605 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12085 20991 14858 21005 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12085 16391 14858 16405 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 36716 14858 36730 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 31914 14858 31928 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 27311 14858 27325 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 22704 14858 22718 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 18122 14858 18136 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 13510 14858 13524 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12082 8904 14858 8918 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12079 11791 14858 11805 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12073 34777 14858 34791 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12073 6028 14858 6042 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12071 30191 14858 30205 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12071 25577 14858 25591 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12071 20977 14858 20991 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12071 16377 14858 16391 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 36730 14858 36744 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 31928 14858 31942 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 27325 14858 27339 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 22718 14858 22732 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 18136 14858 18150 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 13524 14858 13538 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12068 8918 14858 8932 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12065 11777 14858 11791 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12059 34763 14858 34777 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12059 6014 14858 6028 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12057 30177 14858 30191 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12057 25563 14858 25577 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12057 20963 14858 20977 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12057 16363 14858 16377 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 36744 14858 36758 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 31942 14858 31956 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 27339 14858 27353 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 22732 14858 22746 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 18150 14858 18164 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 13538 14858 13552 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12054 8932 14858 8946 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12051 11763 14858 11777 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12045 34749 14858 34763 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12045 6000 14858 6014 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12043 30163 14858 30177 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12043 25549 14858 25563 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12043 20949 14858 20963 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12043 16349 14858 16363 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 36758 14858 36772 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 31956 14858 31970 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 27353 14858 27367 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 22746 14858 22760 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 18164 14858 18178 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 13552 14858 13566 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12040 8946 14858 8960 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12037 11749 14858 11763 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12031 34735 14858 34749 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12031 5986 14858 6000 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12029 30149 14858 30163 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12029 25535 14858 25549 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12029 20935 14858 20949 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12029 16335 14858 16349 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 36772 14858 36786 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 31970 14858 31984 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 27367 14858 27381 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 22760 14858 22774 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 18178 14858 18192 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 13566 14858 13580 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12026 8960 14858 8974 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12023 11735 14858 11749 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12017 34721 14858 34735 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12017 5972 14858 5986 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12015 30135 14858 30149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12015 25521 14858 25535 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12015 20921 14858 20935 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12015 16321 14858 16335 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 36786 14858 36800 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 31984 14858 31998 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 27381 14858 27395 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 22774 14858 22788 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 18192 14858 18206 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 13580 14858 13594 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12012 8974 14858 8988 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12009 11721 14858 11735 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12003 34707 14858 34721 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12003 5958 14858 5972 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12001 30121 14858 30135 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12001 25507 14858 25521 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12001 20907 14858 20921 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 12001 16307 14858 16321 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 36800 14858 36814 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 31998 14858 32012 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 27395 14858 27409 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 22788 14858 22802 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 18206 14858 18220 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 13594 14858 13608 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11998 8988 14858 9002 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11995 11707 14858 11721 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11989 34693 14858 34707 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11989 5944 14858 5958 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11987 30107 14858 30121 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11987 25493 14858 25507 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11987 20893 14858 20907 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11987 16293 14858 16307 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 36814 14858 36828 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 32012 14858 32026 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 27409 14858 27423 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 22802 14858 22816 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 18220 14858 18234 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 13608 14858 13622 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11984 9002 14858 9016 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11981 11693 14858 11707 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11975 34679 14858 34693 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11975 5930 14858 5944 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11973 30093 14858 30107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11973 25479 14858 25493 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11973 20879 14858 20893 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11973 16279 14858 16293 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 36828 14858 36842 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 32026 14858 32040 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 27423 14858 27437 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 22816 14858 22830 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 18234 14858 18248 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 13622 14858 13636 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11970 9016 14858 9030 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11967 11679 14858 11693 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11961 34665 14858 34679 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11961 5916 14858 5930 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11959 30079 14858 30093 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11959 25465 14858 25479 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11959 20865 14858 20879 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11959 16265 14858 16279 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 36842 14858 36856 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 32040 14858 32054 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 27437 14858 27451 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 22830 14858 22844 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 18248 14858 18262 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 13636 14858 13650 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11956 9030 14858 9044 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11953 11665 14858 11679 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11947 34651 14858 34665 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11947 5902 14858 5916 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11945 30065 14858 30079 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11945 25451 14858 25465 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11945 20851 14858 20865 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11945 16251 14858 16265 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 36856 14858 36870 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 32054 14858 32068 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 27451 14858 27465 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 22844 14858 22858 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 18262 14858 18276 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 13650 14858 13664 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11942 9044 14858 9058 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11939 11651 14858 11665 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11933 34637 14858 34651 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11933 5888 14858 5902 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11931 30051 14858 30065 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11931 25437 14858 25451 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11931 20837 14858 20851 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11931 16237 14858 16251 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 36870 14858 36884 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 32068 14858 32082 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 27465 14858 27479 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 22858 14858 22872 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 18276 14858 18290 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 13664 14858 13678 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11928 9058 14858 9072 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11925 11637 14858 11651 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11919 34623 14858 34637 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11919 5874 14858 5888 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11917 30037 14858 30051 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11917 25423 14858 25437 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11917 20823 14858 20837 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11917 16223 14858 16237 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 36884 14858 36898 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 32082 14858 32096 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 27479 14858 27493 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 22872 14858 22886 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 18290 14858 18304 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 13678 14858 13692 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11914 9072 14858 9086 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11911 11623 14858 11637 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11905 34609 14858 34623 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11905 5860 14858 5874 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11903 30023 14858 30037 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11903 25409 14858 25423 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11903 20809 14858 20823 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11903 16209 14858 16223 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 36898 14858 36912 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 32096 14858 32110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 27493 14858 27507 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 22886 14858 22900 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 18304 14858 18318 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 13692 14858 13706 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11900 9086 14858 9100 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11897 11609 14858 11623 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11891 34595 14858 34609 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11891 5846 14858 5860 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11889 30009 14858 30023 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11889 25395 14858 25409 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11889 20795 14858 20809 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11889 16195 14858 16209 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 36912 14858 36926 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 32110 14858 32124 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 27507 14858 27521 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 22900 14858 22914 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 18318 14858 18332 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 13706 14858 13720 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11886 9100 14858 9114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11883 11595 14858 11609 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11877 34581 14858 34595 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11877 5832 14858 5846 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11875 29995 14858 30009 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11875 25381 14858 25395 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11875 20781 14858 20795 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11875 16181 14858 16195 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 36926 14858 36940 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 32124 14858 32138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 27521 14858 27535 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 22914 14858 22928 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 18332 14858 18346 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 13720 14858 13734 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11872 9114 14858 9128 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11869 11581 14858 11595 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11863 34567 14858 34581 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11863 5818 14858 5832 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11861 29981 14858 29995 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11861 25367 14858 25381 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11861 20767 14858 20781 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11861 16167 14858 16181 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 36940 14858 36954 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 32138 14858 32152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 27535 14858 27549 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 22928 14858 22942 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 18346 14858 18360 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 13734 14858 13748 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11858 9128 14858 9142 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11855 11567 14858 11581 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11849 34553 14858 34567 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11849 5804 14858 5818 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11847 29967 14858 29981 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11847 25353 14858 25367 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11847 20753 14858 20767 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11847 16153 14858 16167 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 36954 14858 36968 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 32152 14858 32166 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 27549 14858 27563 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 22942 14858 22956 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 18360 14858 18374 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 13748 14858 13762 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11844 9142 14858 9156 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11841 11553 14858 11567 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11835 34539 14858 34553 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11835 5790 14858 5804 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11833 29953 14858 29967 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11833 25339 14858 25353 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11833 20739 14858 20753 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11833 16139 14858 16153 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 36968 14858 36982 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 32166 14858 32180 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 27563 14858 27577 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 22956 14858 22970 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 18374 14858 18388 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 13762 14858 13776 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11830 9156 14858 9170 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11827 11539 14858 11553 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11821 34525 14858 34539 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11821 5776 14858 5790 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11819 29939 14858 29953 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11819 25325 14858 25339 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11819 20725 14858 20739 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11819 16125 14858 16139 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 36982 14858 36996 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 32180 14858 32194 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 27577 14858 27591 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 22970 14858 22984 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 18388 14858 18402 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 13776 14858 13790 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11816 9170 14858 9184 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11813 11525 14858 11539 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11807 34511 14858 34525 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11807 5762 14858 5776 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11805 29925 14858 29939 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11805 25311 14858 25325 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11805 20711 14858 20725 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11805 16111 14858 16125 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 36996 14858 37010 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 32194 14858 32208 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 27591 14858 27605 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 22984 14858 22998 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 18402 14858 18416 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 13790 14858 13804 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11802 9184 14858 9198 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11799 11511 14858 11525 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11793 34497 14858 34511 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11793 5748 14858 5762 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11791 29911 14858 29925 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11791 25297 14858 25311 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11791 20697 14858 20711 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11791 16097 14858 16111 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 37010 14858 37024 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 32208 14858 32222 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 27605 14858 27619 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 22998 14858 23012 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 18416 14858 18430 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 13804 14858 13818 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11788 9198 14858 9212 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11785 11497 14858 11511 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11779 34483 14858 34497 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11779 5734 14858 5748 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11777 29897 14858 29911 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11777 25283 14858 25297 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11777 20683 14858 20697 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11777 16083 14858 16097 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 37024 14858 37038 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 32222 14858 32236 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 27619 14858 27633 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 23012 14858 23026 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 18430 14858 18444 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 13818 14858 13832 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11774 9212 14858 9226 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11771 11483 14858 11497 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11765 34469 14858 34483 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11765 5720 14858 5734 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11763 29883 14858 29897 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11763 25269 14858 25283 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11763 20669 14858 20683 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11763 16069 14858 16083 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 37038 14858 37052 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 32236 14858 32250 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 27633 14858 27647 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 23026 14858 23040 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 18444 14858 18458 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 13832 14858 13846 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11760 9226 14858 9240 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11757 11469 14858 11483 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11751 34455 14858 34469 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11751 5706 14858 5720 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11749 29869 14858 29883 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11749 25255 14858 25269 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11749 20655 14858 20669 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11749 16055 14858 16069 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 37052 14858 37059 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 32250 14858 32264 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 27647 14858 27661 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 23040 14858 23054 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 18458 14858 18472 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 13846 14858 13860 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11746 9240 14858 9254 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11743 11455 14858 11469 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11737 34441 14858 34455 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11737 5692 14858 5706 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11735 29855 14858 29869 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11735 25241 14858 25255 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11735 20641 14858 20655 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11735 16041 14858 16055 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11732 32264 14858 32278 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11732 27661 14858 27675 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11732 23054 14858 23068 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11732 18472 14858 18486 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11732 13860 14858 13874 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11732 9254 14858 9268 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11729 11441 14858 11455 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11723 34427 14858 34441 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11723 5678 14858 5692 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11721 29841 14858 29855 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11721 25227 14858 25241 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11721 20627 14858 20641 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11721 16027 14858 16041 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11718 32278 14858 32292 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11718 27675 14858 27689 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11718 23068 14858 23082 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11718 18486 14858 18500 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11718 13874 14858 13888 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11718 9268 14858 9282 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11715 11427 14858 11441 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11709 34413 14858 34427 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11709 5664 14858 5678 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11707 29827 14858 29841 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11707 25213 14858 25227 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11707 20613 14858 20627 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11707 16013 14858 16027 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11704 32292 14858 32306 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11704 27689 14858 27703 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11704 23082 14858 23096 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11704 18500 14858 18514 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11704 13888 14858 13902 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11704 9282 14858 9296 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11701 11413 14858 11427 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11695 34399 14858 34413 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11695 5650 14858 5664 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11693 29813 14858 29827 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11693 25199 14858 25213 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11693 20599 14858 20613 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11693 15999 14858 16013 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11690 32306 14858 32320 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11690 27703 14858 27717 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11690 23096 14858 23110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11690 18514 14858 18528 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11690 13902 14858 13916 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11690 9296 14858 9310 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11687 11399 14858 11413 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11681 34385 14858 34399 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11681 5636 14858 5650 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11679 29799 14858 29813 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11679 25185 14858 25199 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11679 20585 14858 20599 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11679 15985 14858 15999 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11676 32320 14858 32334 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11676 27717 14858 27731 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11676 23110 14858 23124 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11676 18528 14858 18542 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11676 13916 14858 13930 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11676 9310 14858 9324 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11673 11385 14858 11399 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11667 34371 14858 34385 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11667 5622 14858 5636 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11665 29785 14858 29799 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11665 25171 14858 25185 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11665 20571 14858 20585 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11665 15971 14858 15985 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11662 32334 14858 32348 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11662 27731 14858 27745 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11662 23124 14858 23138 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11662 18542 14858 18556 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11662 13930 14858 13944 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11662 9324 14858 9338 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11659 11371 14858 11385 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11653 34357 14858 34371 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11653 5608 14858 5622 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11651 29771 14858 29785 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11651 25157 14858 25171 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11651 20557 14858 20571 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11651 15957 14858 15971 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11648 32348 14858 32362 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11648 27745 14858 27759 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11648 23138 14858 23152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11648 18556 14858 18570 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11648 13944 14858 13958 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11648 9338 14858 9352 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11645 11357 14858 11371 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11639 34343 14858 34357 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11639 5594 14858 5608 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11637 29757 14858 29771 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11637 25143 14858 25157 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11637 20543 14858 20557 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11637 15943 14858 15957 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11634 32362 14858 32376 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11634 27759 14858 27773 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11634 23152 14858 23166 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11634 18570 14858 18584 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11634 13958 14858 13972 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11634 9352 14858 9366 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11631 11343 14858 11357 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11625 34329 14858 34343 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11625 5580 14858 5594 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11623 29743 14858 29757 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11623 25129 14858 25143 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11623 20529 14858 20543 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11623 15929 14858 15943 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11620 32376 14858 32390 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11620 27773 14858 27787 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11620 23166 14858 23180 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11620 18584 14858 18598 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11620 13972 14858 13986 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11620 9366 14858 9380 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11617 11329 14858 11343 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11611 34315 14858 34329 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11611 5566 14858 5580 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11609 29729 14858 29743 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11609 25115 14858 25129 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11609 20515 14858 20529 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11609 15915 14858 15929 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11606 32390 14858 32404 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11606 27787 14858 27801 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11606 23180 14858 23194 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11606 18598 14858 18612 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11606 13986 14858 14000 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11606 9380 14858 9394 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11603 11315 14858 11329 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11597 34301 14858 34315 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11597 5552 14858 5566 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11595 29715 14858 29729 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11595 25101 14858 25115 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11595 20501 14858 20515 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11595 15901 14858 15915 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11592 32404 14858 32418 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11592 27801 14858 27815 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11592 23194 14858 23208 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11592 18612 14858 18626 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11592 14000 14858 14014 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11592 9394 14858 9408 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11589 11301 14858 11315 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11583 34287 14858 34301 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11583 5538 14858 5552 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11581 29701 14858 29715 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11581 25087 14858 25101 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11581 20487 14858 20501 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11581 15887 14858 15901 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11578 32418 14858 32432 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11578 27815 14858 27829 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11578 23208 14858 23222 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11578 18626 14858 18640 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11578 14014 14858 14028 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11578 9408 14858 9422 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11575 11287 14858 11301 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11569 34273 14858 34287 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11569 5524 14858 5538 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11567 29687 14858 29701 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11567 25073 14858 25087 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11567 20473 14858 20487 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11567 15873 14858 15887 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11564 32432 14858 32446 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11564 27829 14858 27843 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11564 23222 14858 23236 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11564 18640 14858 18654 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11564 14028 14858 14042 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11564 9422 14858 9436 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11561 11273 14858 11287 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11555 34259 14858 34273 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11555 5510 14858 5524 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11553 29673 14858 29687 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11553 25059 14858 25073 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11553 20459 14858 20473 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11553 15859 14858 15873 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11550 32446 14858 32460 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11550 27843 14858 27857 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11550 23236 14858 23250 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11550 18654 14858 18668 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11550 14042 14858 14056 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11550 9436 14858 9450 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11547 11259 14858 11273 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11541 34245 14858 34259 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11541 5496 14858 5510 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11539 29659 14858 29673 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11539 25045 14858 25059 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11539 20445 14858 20459 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11539 15845 14858 15859 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11536 32460 14858 32474 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11536 27857 14858 27871 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11536 23250 14858 23264 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11536 18668 14858 18682 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11536 14056 14858 14070 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11536 9450 14858 9464 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11533 11245 14858 11259 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11527 34231 14858 34245 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11527 5482 14858 5496 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11525 29645 14858 29659 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11525 25031 14858 25045 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11525 20431 14858 20445 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11525 15831 14858 15845 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11522 32474 14858 32488 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11522 27871 14858 27885 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11522 23264 14858 23278 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11522 18682 14858 18691 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11522 14070 14858 14084 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11522 9464 14858 9478 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11519 11231 14858 11245 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11513 5468 14858 5482 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11511 29631 14858 29645 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11508 32488 14858 32491 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11508 27885 14858 27891 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11508 23278 14858 23291 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11508 14084 14858 14091 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11508 9478 14858 9491 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11499 5454 14858 5468 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11485 5440 14858 5454 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11471 5426 14858 5440 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11457 5412 14858 5426 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11443 5398 14858 5412 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11429 5384 14858 5398 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11415 5370 14858 5384 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11401 5356 14858 5370 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11387 5342 14858 5356 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11373 5328 14858 5342 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11359 5314 14858 5328 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11345 5300 14858 5314 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11331 5286 14858 5300 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11317 5272 14858 5286 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11303 5258 14858 5272 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11289 5244 14858 5258 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11275 5230 14858 5244 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11261 5216 14858 5230 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11247 5202 14858 5216 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11233 5188 14858 5202 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11219 5174 14858 5188 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11205 5160 14858 5174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11191 5146 14858 5160 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 11177 5132 14858 5146 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10078 1725 14858 1739 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10078 0 14858 1725 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10064 1739 14858 1753 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10050 1753 14858 1767 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10036 1767 14858 1781 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10022 1781 14858 1795 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 10008 1795 14858 1809 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9994 1809 14858 1823 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9980 1823 14858 1837 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9966 1837 14858 1851 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9952 1851 14858 1865 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9938 1865 14858 1879 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9924 1879 14858 1893 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9910 1893 14858 1907 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9896 1907 14858 1921 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9882 1921 14858 1935 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9868 1935 14858 1949 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9854 1949 14858 1963 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9840 1963 14858 1977 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9826 1977 14858 1991 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9812 1991 14858 2005 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9798 2005 14858 2019 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9784 2019 14858 2033 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9770 2033 14858 2047 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9756 2047 14858 2061 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9742 2061 14858 2075 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9728 2075 14858 2089 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9714 2089 14858 2103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9700 2103 14858 2117 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9686 2117 14858 2131 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9672 2131 14858 2145 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9658 2145 14858 2159 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9644 2159 14858 2173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9630 2173 14858 2187 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9616 2187 14858 2201 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9602 2201 14858 2215 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9588 2215 14858 2229 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9574 2229 14858 2243 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9560 2243 14858 2257 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9546 2257 14858 2271 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9532 2271 14858 2285 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9518 2285 14858 2299 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9504 2299 14858 2313 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9490 2313 14858 2327 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9476 2327 14858 2341 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9462 2341 14858 2355 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9448 2355 14858 2369 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9434 2369 14858 2383 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9420 2383 14858 2397 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9406 2397 14858 2411 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9392 2411 14858 2425 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9378 2425 14858 2439 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9364 2439 14858 2453 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 9350 2453 14858 2459 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 7578 2459 14858 5132 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4964 23291 14858 25031 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4964 18691 14858 20431 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4964 15123 14858 15831 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4964 15121 14858 15123 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4964 14597 14858 14611 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4964 14091 14858 14597 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4962 15107 14858 15121 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4950 14611 14858 14625 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4948 15093 14858 15107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4936 14625 14858 14639 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4934 15079 14858 15093 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4922 14639 14858 14653 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4920 15065 14858 15079 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4908 14653 14858 14667 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4906 15051 14858 15065 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4894 14667 14858 14681 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4892 15037 14858 15051 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4880 14681 14858 14695 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4878 15023 14858 15037 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4866 14695 14858 14709 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4864 15009 14858 15023 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4852 14709 14858 14723 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4850 14995 14858 15009 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4838 14723 14858 14737 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4836 14981 14858 14995 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4824 14737 14858 14751 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4822 14967 14858 14981 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4810 14751 14858 14765 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4808 14953 14858 14967 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4796 14765 14858 14779 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4794 14939 14858 14953 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4782 14779 14858 14793 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4780 14925 14858 14939 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4768 14793 14858 14807 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4766 14911 14858 14925 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4754 14807 14858 14821 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4752 14897 14858 14911 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4740 14821 14858 14831 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 4738 14883 14858 14897 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3770 11219 14858 11231 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3758 11205 14858 11219 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3744 11191 14858 11205 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3730 11177 14858 11191 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3716 11163 14858 11177 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3702 11149 14858 11163 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3688 11135 14858 11149 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3682 14831 14858 14883 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3674 11121 14858 11135 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3660 11107 14858 11121 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3650 29622 14858 29631 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3646 11093 14858 11107 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3641 29608 14858 29622 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3632 11079 14858 11093 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3627 29594 14858 29608 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3618 11065 14858 11079 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3613 29580 14858 29594 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3604 11051 14858 11065 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3599 29566 14858 29580 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3590 11037 14858 11051 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3585 29552 14858 29566 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3576 11023 14858 11037 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3571 29538 14858 29552 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3562 11009 14858 11023 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3557 29524 14858 29538 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3548 10995 14858 11009 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3543 29510 14858 29524 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3534 10981 14858 10995 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3529 29496 14858 29510 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3520 10967 14858 10981 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3515 29482 14858 29496 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3506 10953 14858 10967 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3501 29468 14858 29482 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3487 29454 14858 29468 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3473 29440 14858 29454 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3459 29426 14858 29440 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3445 29412 14858 29426 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3431 29398 14858 29412 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3417 29384 14858 29398 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3403 29370 14858 29384 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3389 29356 14858 29370 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3375 29342 14858 29356 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3361 32491 14858 34231 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3361 27891 14858 29342 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3361 9491 14858 10953 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 3124 37059 14858 38003 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 33827 11857 33857 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 22088 11857 33827 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 22072 11857 22088 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10641 22042 11857 22072 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10627 33857 11857 33887 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10611 22012 11857 22042 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10597 33887 11857 33917 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10581 21982 11857 22012 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10567 33917 11857 33947 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10551 21952 11857 21982 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10537 33947 11857 33977 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10521 21922 11857 21952 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10507 33977 11857 34007 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10491 21892 11857 21922 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10477 34007 11857 34037 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10461 21862 11857 21892 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10447 34037 11857 34067 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10431 21832 11857 21862 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10417 34067 11857 34097 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10401 21802 11857 21832 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10387 34097 11857 34127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10371 21772 11857 21802 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10357 34127 11857 34157 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10341 21742 11857 21772 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10327 34157 11857 34187 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10311 21712 11857 21742 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10297 34187 11857 34217 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10281 21682 11857 21712 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10267 34217 11857 34247 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10251 21652 11857 21682 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10237 34247 11857 34277 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10221 21622 11857 21652 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10207 34277 11857 34307 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10191 21592 11857 21622 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10177 34307 11857 34337 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10161 21563 11828 21592 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10147 34337 11857 34367 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10132 21533 11798 21563 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10117 34367 11857 34397 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10102 21503 11768 21533 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10087 34397 11857 34427 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10072 21473 11738 21503 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10057 34427 11857 34457 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10042 21443 11708 21473 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10027 34457 11857 34487 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10012 21413 11678 21443 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9997 34487 11857 34517 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9982 21383 11648 21413 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9967 34517 11857 34529 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37072 14325 38008 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37064 14317 37072 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37034 14287 37064 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37004 14257 37034 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36974 14227 37004 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36944 14197 36974 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36914 14167 36944 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36884 14137 36914 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36854 14107 36884 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36824 14077 36854 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36794 14047 36824 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36764 14017 36794 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36734 13987 36764 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36704 13957 36734 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36674 13927 36704 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36644 13897 36674 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36614 13867 36644 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36584 13837 36614 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36554 13807 36584 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36524 13777 36554 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36494 13747 36524 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36464 13717 36494 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36434 13687 36464 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36404 13657 36434 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36374 13627 36404 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36344 13597 36374 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36314 13567 36344 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36284 13537 36314 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36254 13507 36284 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36224 13477 36254 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36194 13447 36224 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36164 13417 36194 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36134 13387 36164 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36104 13357 36134 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36074 13327 36104 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36044 13297 36074 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36014 13267 36044 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35984 13237 36014 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35954 13207 35984 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35924 13177 35954 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35894 13147 35924 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35864 13117 35894 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35834 13087 35864 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35804 13057 35834 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35774 13027 35804 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35744 12997 35774 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35714 12967 35744 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35684 12937 35714 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35654 12907 35684 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35624 12877 35654 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35594 12847 35624 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35564 12817 35594 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35534 12787 35564 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35504 12757 35534 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35474 12727 35504 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35444 12697 35474 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35414 12667 35444 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35384 12637 35414 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35354 12607 35384 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35324 12577 35354 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35294 12547 35324 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35264 12517 35294 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35234 12487 35264 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35204 12457 35234 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35174 12427 35204 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35144 12397 35174 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35114 12367 35144 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35084 12337 35114 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35054 12307 35084 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35024 12277 35054 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34994 12247 35024 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34964 12217 34994 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34934 12187 34964 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34904 12157 34934 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34874 12127 34904 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34844 12097 34874 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34814 12067 34844 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34784 12037 34814 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34754 12007 34784 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34724 11977 34754 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34694 11947 34724 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34664 11917 34694 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34634 11887 34664 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34604 11857 34634 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34529 11857 34604 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9952 21353 11618 21383 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9922 21323 11588 21353 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9892 21293 11558 21323 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9862 21263 11528 21293 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9832 21233 11498 21263 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9802 21203 11468 21233 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9772 21173 11438 21203 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9742 21143 11408 21173 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9712 21113 11378 21143 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9682 21083 11348 21113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9652 21053 11318 21083 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9622 21023 11288 21053 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9592 20993 11258 21023 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9562 20963 11228 20993 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9532 20933 11198 20963 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9502 20903 11168 20933 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9472 20873 11138 20903 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9442 20843 11108 20873 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9412 20813 11078 20843 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9382 20783 11048 20813 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9352 20753 11018 20783 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9322 20723 10988 20753 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9292 20693 10958 20723 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9262 20663 10928 20693 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9232 20633 10898 20663 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9202 20603 10868 20633 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9172 20573 10838 20603 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9142 20543 10808 20573 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9112 20513 10778 20543 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9082 20483 10748 20513 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20463 10728 20483 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20433 10698 20463 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20403 10668 20433 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20373 10638 20403 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20343 10608 20373 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20313 10578 20343 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20283 10548 20313 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20253 10518 20283 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20223 10488 20253 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20193 10458 20223 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20163 10428 20193 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20133 10398 20163 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20103 10368 20133 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20073 10338 20103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20043 10308 20073 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20033 10298 20043 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9042 20003 10268 20033 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9012 19973 10238 20003 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8982 19943 10208 19973 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8952 19922 10208 19943 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8931 19901 10208 19922 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 34092 9771 34122 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 22124 9771 34092 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 22110 9771 22124 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8557 22080 9771 22110 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8541 34122 9771 34152 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8527 22050 9771 22080 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8511 34152 9771 34182 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8497 22020 9771 22050 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8481 34182 9771 34212 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8467 21990 9771 22020 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8451 34212 9771 34242 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8437 21960 9771 21990 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8421 34242 9771 34272 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8407 21930 9771 21960 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8391 34272 9771 34302 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8377 21900 9771 21930 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8361 34302 9771 34332 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8347 21870 9771 21900 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8331 34332 9771 34362 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8317 21840 9771 21870 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8301 34362 9771 34392 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8287 21810 9771 21840 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8271 34392 9771 34422 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8257 21780 9771 21810 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8241 34422 9771 34452 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8227 21750 9771 21780 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8211 34452 9771 34482 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8197 21720 9771 21750 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8181 34482 9771 34512 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8167 21690 9771 21720 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8151 34512 9771 34542 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8137 21660 9771 21690 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8121 34542 9771 34572 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8107 21630 9771 21660 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8091 34572 9771 34602 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8077 21611 9752 21630 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8061 34602 9771 34632 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8058 21581 9722 21611 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8031 34632 9771 34662 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8028 21551 9692 21581 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8001 34662 9771 34692 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7998 21521 9662 21551 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7971 34692 9771 34722 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7968 21491 9632 21521 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7941 34722 9771 34752 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7938 21461 9602 21491 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7911 34752 9771 34782 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7908 21431 9572 21461 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7881 34782 9771 34812 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7878 21401 9542 21431 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7851 34812 9771 34842 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7848 21371 9512 21401 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7821 34842 9771 34872 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7818 21341 9482 21371 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7791 34872 9771 34902 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7788 21311 9452 21341 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7761 34902 9771 34932 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7758 21281 9422 21311 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7731 34932 9771 34962 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7728 21251 9392 21281 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7701 34962 9771 34992 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7698 21221 9362 21251 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7671 34992 9771 35022 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7668 21191 9332 21221 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7641 35022 9771 35052 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7638 21161 9302 21191 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7611 35052 9771 35070 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7608 21131 9272 21161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7593 35070 9771 38004 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21117 9258 21131 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21087 9228 21117 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21057 9198 21087 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21027 9168 21057 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20997 9138 21027 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20967 9108 20997 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20937 9078 20967 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20907 9048 20937 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20877 9018 20907 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20847 8988 20877 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20817 8958 20847 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20787 8928 20817 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20757 8898 20787 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20727 8868 20757 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20697 8838 20727 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20667 8808 20697 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20637 8778 20667 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20607 8748 20637 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20577 8718 20607 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20547 8688 20577 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20517 8658 20547 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20487 8628 20517 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20457 8598 20487 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20427 8568 20457 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20043 8568 20427 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20021 8568 20043 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19991 8590 20021 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19961 8620 19991 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19931 8650 19961 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19901 8680 19931 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19660 10208 19901 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19650 10198 19660 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19620 10168 19650 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19590 10138 19620 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19560 10108 19590 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19530 10078 19560 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19500 10048 19530 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19470 10018 19500 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19440 9988 19470 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19410 9958 19440 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19380 9928 19410 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19350 9898 19380 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19320 9868 19350 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19290 9838 19320 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19260 9808 19290 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19230 9778 19260 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 0 9778 19230 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal2 s 5179 0 5579 107 6 OGC_HVC
port 5 nsew power bidirectional
rlabel metal3 s 99 0 4879 7302 6 P_CORE
port 6 nsew power bidirectional
rlabel metal3 s 10078 0 14858 10000 6 P_CORE
port 6 nsew power bidirectional
rlabel metal2 s 10934 7651 11383 7665 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10934 7223 11383 7651 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10920 7665 11383 7679 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10906 7679 11383 7693 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10892 7693 11383 7707 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10878 7707 11383 7721 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10864 7721 11383 7735 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10850 7735 11383 7749 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10836 7749 11383 7763 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10822 7763 11383 7777 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10808 7777 11383 7791 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10794 7791 11383 7805 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10780 7805 11383 7819 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10766 7819 11383 7833 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10752 7833 11383 7847 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10738 7847 11383 7861 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10724 7861 11383 7875 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10710 7875 11383 7889 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10696 7889 11383 7903 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10682 7903 11383 7917 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10668 7917 11383 7931 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10654 7931 11383 7933 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10652 7933 11369 7947 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10638 7947 11355 7961 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10624 7961 11341 7975 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10610 7975 11327 7989 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10596 7989 11313 8003 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10582 8003 11299 8017 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10568 8017 11285 8031 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10554 8031 11271 8045 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10540 8045 11257 8059 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 10526 8059 11246 8070 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 9403 2824 9411 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 9063 2824 9403 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 9050 2824 9063 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 9036 2837 9050 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 9022 2851 9036 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 9008 2865 9022 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8994 2879 9008 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8980 2893 8994 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8966 2907 8980 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8952 2921 8966 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8938 2935 8952 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8924 2949 8938 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8910 2963 8924 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8896 2977 8910 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8882 2991 8896 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8868 3005 8882 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8854 3019 8868 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8840 3033 8854 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8826 3047 8840 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8812 3061 8826 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8798 3075 8812 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8784 3089 8798 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8770 3103 8784 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8756 3117 8770 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8742 3131 8756 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8728 3145 8742 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8714 3159 8728 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8700 3173 8714 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8686 3187 8700 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8672 3201 8686 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8658 3215 8672 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8644 3229 8658 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8630 3243 8644 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8616 3257 8630 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8602 3271 8616 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8588 3285 8602 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8574 3299 8588 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8560 3313 8574 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8546 3327 8560 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8532 3341 8546 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8518 3355 8532 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8504 3369 8518 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8490 3383 8504 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8476 3397 8490 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8462 10840 8476 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8448 10854 8462 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8434 10868 8448 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8420 10882 8434 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8406 10896 8420 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8392 10910 8406 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8378 10924 8392 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8364 10938 8378 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8350 10952 8364 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8336 10966 8350 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8322 10980 8336 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8308 10994 8322 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8294 11008 8308 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8280 11022 8294 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8266 11036 8280 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8252 11050 8266 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8238 11064 8252 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8224 11078 8238 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8210 11092 8224 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8196 11106 8210 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8182 11120 8196 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8168 11134 8182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8154 11148 8168 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8140 11162 8154 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8126 11176 8140 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8112 11190 8126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8098 11204 8112 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8084 11218 8098 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8070 11232 8084 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8060 3968 8070 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8046 3954 8060 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8032 3940 8046 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8018 3926 8032 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 8004 3912 8018 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7990 3898 8004 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7976 3884 7990 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7962 3870 7976 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7948 3856 7962 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7934 3842 7948 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7920 3828 7934 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7906 3814 7920 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7892 3800 7906 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7878 3786 7892 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7864 3772 7878 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7850 3758 7864 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7836 3744 7850 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7822 3730 7836 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7808 3716 7822 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7794 3702 7808 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7780 3688 7794 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7766 3674 7780 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7752 3660 7766 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7738 3646 7752 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7724 3632 7738 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7710 3618 7724 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7696 3604 7710 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7682 3590 7696 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7668 3576 7682 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7654 3562 7668 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7640 3548 7654 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7626 3534 7640 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7612 3520 7626 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7598 3506 7612 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7584 3492 7598 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7570 3478 7584 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7556 3464 7570 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7542 3450 7556 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7528 3436 7542 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7514 3422 7528 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7500 3408 7514 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7486 3394 7500 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7472 3380 7486 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7458 3366 7472 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7444 3352 7458 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7430 3338 7444 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7416 3324 7430 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7402 3310 7416 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7388 3296 7402 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 218 7387 3295 7388 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 217 7379 3287 7387 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 210 9411 2824 9419 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 209 7371 3279 7379 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 202 9419 2824 9420 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38112 13440 39015 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38099 3006 38112 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38085 2992 38099 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38071 2978 38085 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38057 2964 38071 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38043 2950 38057 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38029 2936 38043 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38015 2922 38029 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 38001 2908 38015 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37987 2894 38001 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37973 2880 37987 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37959 2866 37973 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37945 2852 37959 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37931 2838 37945 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37917 2824 37931 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37011 2824 37917 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 37010 2824 37011 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36996 2825 37010 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36982 2839 36996 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36968 2853 36982 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36954 2867 36968 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36940 2881 36954 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36926 2895 36940 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36912 2909 36926 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36898 2923 36912 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36884 2937 36898 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36870 2951 36884 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36856 2965 36870 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36842 2979 36856 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36828 2993 36842 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36814 3007 36828 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36800 3021 36814 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36786 3035 36800 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36772 3049 36786 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36758 3063 36772 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36744 3077 36758 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36730 3091 36744 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36716 3105 36730 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36702 3119 36716 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36688 3133 36702 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36674 3147 36688 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36660 3161 36674 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36646 3175 36660 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36632 3189 36646 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36618 3203 36632 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36604 3217 36618 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36590 3231 36604 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36576 3245 36590 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36562 3259 36576 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36548 3273 36562 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36534 3287 36548 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36520 3301 36534 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36506 3315 36520 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36492 3329 36506 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36478 3343 36492 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36464 3357 36478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36450 3371 36464 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36436 3385 36450 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36422 3399 36436 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36408 3413 36422 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36394 3427 36408 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36380 3441 36394 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36366 3455 36380 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36352 3469 36366 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36338 3483 36352 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36324 3497 36338 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36310 3511 36324 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 36296 3525 36310 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34556 11592 36296 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34544 3524 34556 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34530 3510 34544 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34516 3496 34530 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34502 3482 34516 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34488 3468 34502 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34474 3454 34488 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34460 3440 34474 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34446 3426 34460 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34432 3412 34446 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34418 3398 34432 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34404 3384 34418 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34390 3370 34404 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34376 3356 34390 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34362 3342 34376 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34348 3328 34362 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34334 3314 34348 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34320 3300 34334 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34306 3286 34320 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34292 3272 34306 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34278 3258 34292 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34264 3244 34278 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34250 3230 34264 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34236 3216 34250 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34222 3202 34236 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34208 3188 34222 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34194 3174 34208 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34180 3160 34194 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34166 3146 34180 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34152 3132 34166 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34138 3118 34152 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34124 3104 34138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34110 3090 34124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34096 3076 34110 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34082 3062 34096 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34068 3048 34082 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34054 3034 34068 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34040 3020 34054 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34026 3006 34040 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 34012 2992 34026 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33998 2978 34012 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33984 2964 33998 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33970 2950 33984 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33956 2936 33970 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33942 2922 33956 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33928 2908 33942 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33914 2894 33928 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33900 2880 33914 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33886 2866 33900 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33872 2852 33886 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33858 2838 33872 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 33844 2824 33858 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32416 2824 33844 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32410 2824 32416 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32396 2830 32410 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32382 2844 32396 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32368 2858 32382 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32354 2872 32368 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32340 2886 32354 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32326 2900 32340 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32312 2914 32326 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32298 2928 32312 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32284 2942 32298 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32270 2956 32284 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32256 2970 32270 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32242 2984 32256 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32228 2998 32242 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32214 3012 32228 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32200 3026 32214 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32186 3040 32200 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32172 3054 32186 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32158 3068 32172 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32144 3082 32158 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32130 3096 32144 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32116 3110 32130 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32102 3124 32116 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32088 3138 32102 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32074 3152 32088 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32060 3166 32074 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32046 3180 32060 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32032 3194 32046 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32018 3208 32032 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 32004 3222 32018 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31990 3236 32004 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31976 3250 31990 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31962 3264 31976 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31948 3278 31962 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31934 3292 31948 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31920 3306 31934 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31906 3320 31920 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31892 3334 31906 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31878 3348 31892 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31864 3362 31878 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31850 3376 31864 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31836 3390 31850 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31822 3404 31836 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31808 3418 31822 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31794 3432 31808 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31780 3446 31794 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31766 3460 31780 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31752 3474 31766 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31738 3488 31752 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31724 3502 31738 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31710 3516 31724 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 31696 3530 31710 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29956 11341 31696 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29943 3524 29956 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29929 3510 29943 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29915 3496 29929 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29901 3482 29915 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29887 3468 29901 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29873 3454 29887 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29859 3440 29873 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29845 3426 29859 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29831 3412 29845 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29817 3398 29831 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29803 3384 29817 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29789 3370 29803 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29775 3356 29789 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29761 3342 29775 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29747 3328 29761 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29733 3314 29747 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29719 3300 29733 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29705 3286 29719 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29691 3272 29705 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29677 3258 29691 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29663 3244 29677 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29649 3230 29663 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29635 3216 29649 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29621 3202 29635 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29607 3188 29621 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29593 3174 29607 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29579 3160 29593 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29565 3146 29579 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29551 3132 29565 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29537 3118 29551 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29523 3104 29537 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29509 3090 29523 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29495 3076 29509 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29481 3062 29495 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29467 3048 29481 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29453 3034 29467 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29439 3020 29453 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29425 3006 29439 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29411 2992 29425 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29397 2978 29411 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29383 2964 29397 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29369 2950 29383 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29355 2936 29369 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29341 2922 29355 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29327 2908 29341 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29313 2894 29327 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29299 2880 29313 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29285 2866 29299 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29271 2852 29285 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29257 2838 29271 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 29243 2824 29257 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27834 2824 29243 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27824 2824 27834 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27810 2834 27824 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27796 2848 27810 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27782 2862 27796 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27768 2876 27782 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27754 2890 27768 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27740 2904 27754 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27726 2918 27740 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27712 2932 27726 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27698 2946 27712 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27684 2960 27698 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27670 2974 27684 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27656 2988 27670 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27642 3002 27656 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27628 3016 27642 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27614 3030 27628 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27600 3044 27614 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27586 3058 27600 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27572 3072 27586 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27558 3086 27572 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27544 3100 27558 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27530 3114 27544 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27516 3128 27530 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27502 3142 27516 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27488 3156 27502 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27474 3170 27488 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27460 3184 27474 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27446 3198 27460 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27432 3212 27446 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27418 3226 27432 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27404 3240 27418 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27390 3254 27404 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27376 3268 27390 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27362 3282 27376 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27348 3296 27362 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27334 3310 27348 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27320 3324 27334 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27306 3338 27320 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27292 3352 27306 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27278 3366 27292 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27264 3380 27278 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27250 3394 27264 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27236 3408 27250 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27222 3422 27236 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27208 3436 27222 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27194 3450 27208 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27180 3464 27194 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27166 3478 27180 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27152 3492 27166 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27138 3506 27152 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27124 3520 27138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27110 3534 27124 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 27096 3548 27110 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25356 11341 27096 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25343 3538 25356 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25329 3524 25343 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25315 3510 25329 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25301 3496 25315 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25287 3482 25301 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25273 3468 25287 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25259 3454 25273 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25245 3440 25259 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25231 3426 25245 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25217 3412 25231 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25203 3398 25217 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25189 3384 25203 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25175 3370 25189 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25161 3356 25175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25147 3342 25161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25133 3328 25147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25119 3314 25133 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25105 3300 25119 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25091 3286 25105 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25077 3272 25091 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25063 3258 25077 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25049 3244 25063 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25035 3230 25049 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25021 3216 25035 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 25007 3202 25021 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24993 3188 25007 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24979 3174 24993 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24965 3160 24979 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24951 3146 24965 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24937 3132 24951 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24923 3118 24937 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24909 3104 24923 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24895 3090 24909 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24881 3076 24895 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24867 3062 24881 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24853 3048 24867 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24839 3034 24853 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24825 3020 24839 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24811 3006 24825 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24797 2992 24811 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24783 2978 24797 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24769 2964 24783 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24755 2950 24769 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24741 2936 24755 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24727 2922 24741 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24713 2908 24727 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24699 2894 24713 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24685 2880 24699 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24671 2866 24685 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24657 2852 24671 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24643 2838 24657 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 24629 2824 24643 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23213 2824 24629 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23210 2824 23213 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23196 2827 23210 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23182 2841 23196 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23168 2855 23182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23154 2869 23168 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23140 2883 23154 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23126 2897 23140 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23112 2911 23126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23098 2925 23112 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23084 2939 23098 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23070 2953 23084 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23056 2967 23070 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23042 2981 23056 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23028 2995 23042 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23014 3009 23028 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 23000 3023 23014 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22986 3037 23000 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22972 3051 22986 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22958 3065 22972 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22944 3079 22958 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22930 3093 22944 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22916 3107 22930 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22902 3121 22916 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22888 3135 22902 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22874 3149 22888 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22860 3163 22874 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22846 3177 22860 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22832 3191 22846 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22818 3205 22832 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22804 3219 22818 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22790 3233 22804 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22776 3247 22790 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22762 3261 22776 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22748 3275 22762 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22734 3289 22748 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22720 3303 22734 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22706 3317 22720 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22692 3331 22706 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22678 3345 22692 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22664 3359 22678 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22650 3373 22664 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22636 3387 22650 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22622 3401 22636 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22608 3415 22622 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22594 3429 22608 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22580 3443 22594 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22566 3457 22580 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22552 3471 22566 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22538 3485 22552 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22524 3499 22538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22510 3513 22524 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 22496 3527 22510 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20756 11341 22496 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20748 3524 20756 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20734 3510 20748 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20720 3496 20734 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20706 3482 20720 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20692 3468 20706 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20678 3454 20692 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20664 3440 20678 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20650 3426 20664 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20636 3412 20650 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20622 3398 20636 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20608 3384 20622 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20594 3370 20608 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20580 3356 20594 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20566 3342 20580 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20552 3328 20566 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20538 3314 20552 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20524 3300 20538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20510 3286 20524 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20496 3272 20510 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20482 3258 20496 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20468 3244 20482 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20454 3230 20468 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20440 3216 20454 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20426 3202 20440 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20412 3188 20426 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20398 3174 20412 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20384 3160 20398 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20370 3146 20384 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20356 3132 20370 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20342 3118 20356 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20328 3104 20342 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20314 3090 20328 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20300 3076 20314 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20286 3062 20300 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20272 3048 20286 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20258 3034 20272 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20244 3020 20258 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20230 3006 20244 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20216 2992 20230 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20202 2978 20216 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20188 2964 20202 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20174 2950 20188 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20160 2936 20174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20146 2922 20160 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20132 2908 20146 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20118 2894 20132 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20104 2880 20118 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20090 2866 20104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20076 2852 20090 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20062 2838 20076 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 20048 2824 20062 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18605 2824 20048 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18596 2824 18605 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18582 2833 18596 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18568 2847 18582 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18554 2861 18568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18540 2875 18554 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18526 2889 18540 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18512 2903 18526 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18498 2917 18512 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18484 2931 18498 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18470 2945 18484 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18456 2959 18470 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18442 2973 18456 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18428 2987 18442 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18414 3001 18428 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18400 3015 18414 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18386 3029 18400 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18372 3043 18386 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18358 3057 18372 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18344 3071 18358 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18330 3085 18344 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18316 3099 18330 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18302 3113 18316 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18288 3127 18302 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18274 3141 18288 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18260 3155 18274 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18246 3169 18260 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18232 3183 18246 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18218 3197 18232 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18204 3211 18218 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18190 3225 18204 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18176 3239 18190 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18162 3253 18176 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18148 3267 18162 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18134 3281 18148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18120 3295 18134 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18106 3309 18120 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18092 3323 18106 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18078 3337 18092 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18064 3351 18078 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18050 3365 18064 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18036 3379 18050 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18022 3393 18036 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 18008 3407 18022 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17994 3421 18008 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17980 3435 17994 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17966 3449 17980 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17952 3463 17966 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17938 3477 17952 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17924 3491 17938 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17910 3505 17924 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 17896 3519 17910 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16156 11341 17896 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16148 3524 16156 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16134 3510 16148 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16120 3496 16134 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16106 3482 16120 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16092 3468 16106 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16078 3454 16092 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16064 3440 16078 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16050 3426 16064 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16036 3412 16050 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16022 3398 16036 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 16008 3384 16022 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15994 3370 16008 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15980 3356 15994 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15966 3342 15980 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15952 3328 15966 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15938 3314 15952 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15924 3300 15938 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15910 3286 15924 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15896 3272 15910 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15882 3258 15896 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15868 3244 15882 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15854 3230 15868 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15840 3216 15854 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15826 3202 15840 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15812 3188 15826 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15798 3174 15812 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15784 3160 15798 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15770 3146 15784 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15756 3132 15770 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15742 3118 15756 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15728 3104 15742 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15714 3090 15728 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15700 3076 15714 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15686 3062 15700 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15672 3048 15686 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15658 3034 15672 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15644 3020 15658 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15630 3006 15644 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15616 2992 15630 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15602 2978 15616 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15588 2964 15602 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15574 2950 15588 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15560 2936 15574 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15546 2922 15560 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15532 2908 15546 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15518 2894 15532 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15504 2880 15518 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15490 2866 15504 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15476 2852 15490 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15462 2838 15476 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 15448 2824 15462 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 14005 2824 15448 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13996 2824 14005 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13982 2833 13996 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13968 2847 13982 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13954 2861 13968 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13940 2875 13954 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13926 2889 13940 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13912 2903 13926 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13898 2917 13912 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13884 2931 13898 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13870 2945 13884 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13856 2959 13870 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13842 2973 13856 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13828 2987 13842 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13814 3001 13828 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13800 3015 13814 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13786 3029 13800 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13772 3043 13786 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13758 3057 13772 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13744 3071 13758 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13730 3085 13744 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13716 3099 13730 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13702 3113 13716 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13688 3127 13702 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13674 3141 13688 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13660 3155 13674 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13646 3169 13660 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13632 3183 13646 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13618 3197 13632 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13604 3211 13618 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13590 3225 13604 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13576 3239 13590 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13562 3253 13576 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13548 3267 13562 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13534 3281 13548 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13520 3295 13534 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13506 3309 13520 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13492 3323 13506 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13478 3337 13492 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13464 3351 13478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13450 3365 13464 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13436 3379 13450 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13422 3393 13436 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13408 3407 13422 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13394 3421 13408 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13380 3435 13394 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13366 3449 13380 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13352 3463 13366 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13338 3477 13352 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13324 3491 13338 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13310 3505 13324 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 13296 3519 13310 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11556 11342 13296 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11543 3524 11556 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11529 3510 11543 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11515 3496 11529 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11501 3482 11515 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11487 3468 11501 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11473 3454 11487 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11459 3440 11473 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11445 3426 11459 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11431 3412 11445 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11417 3398 11431 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11403 3384 11417 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11389 3370 11403 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11375 3356 11389 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11361 3342 11375 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11347 3328 11361 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11333 3314 11347 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11319 3300 11333 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11305 3286 11319 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11291 3272 11305 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11277 3258 11291 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11263 3244 11277 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11249 3230 11263 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11235 3216 11249 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11221 3202 11235 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11207 3188 11221 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11193 3174 11207 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11179 3160 11193 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11165 3146 11179 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11151 3132 11165 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11137 3118 11151 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11123 3104 11137 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11109 3090 11123 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11095 3076 11109 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11081 3062 11095 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11067 3048 11081 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11053 3034 11067 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11039 3020 11053 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11025 3006 11039 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 11011 2992 11025 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10997 2978 11011 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10983 2964 10997 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10969 2950 10983 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10955 2936 10969 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10941 2922 10955 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10927 2908 10941 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10913 2894 10927 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10899 2880 10913 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10885 2866 10899 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10871 2852 10885 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10857 2838 10871 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 10843 2824 10857 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 9420 2824 10843 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7357 3265 7371 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7343 3251 7357 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7329 3237 7343 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7315 3223 7329 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7301 3209 7315 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7287 3195 7301 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7273 3181 7287 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7259 3167 7273 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7245 3153 7259 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7231 3139 7245 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7217 3125 7231 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7203 3111 7217 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7189 3097 7203 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7175 3083 7189 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7161 3069 7175 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7147 3055 7161 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 7133 3041 7147 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5863 3041 7133 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5854 3041 5863 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5840 3050 5854 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5826 3064 5840 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5812 3078 5826 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5798 3092 5812 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5784 3106 5798 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5770 3120 5784 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5756 3134 5770 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5742 3148 5756 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5728 3162 5742 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5714 3176 5728 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5700 3190 5714 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5686 3204 5700 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5672 3218 5686 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5658 3232 5672 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5644 3246 5658 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5630 3260 5644 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5616 3274 5630 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5602 3288 5616 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5588 3302 5602 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5574 3316 5588 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5560 3330 5574 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5546 3344 5560 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5532 3358 5546 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5518 3372 5532 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5504 3386 5518 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5490 3400 5504 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5476 3414 5490 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5462 3428 5476 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5448 3442 5462 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5434 3456 5448 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5420 3470 5434 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5406 3484 5420 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5392 3498 5406 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5378 3512 5392 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5364 3526 5378 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5350 3540 5364 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5336 3554 5350 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5322 3568 5336 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5308 3582 5322 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5294 3596 5308 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5280 3610 5294 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5266 3624 5280 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5252 3638 5266 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5238 3652 5252 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5224 3666 5238 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5210 3680 5224 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5196 3694 5210 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5182 3708 5196 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5168 3722 5182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5154 3736 5168 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 5140 3750 5154 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2480 7379 5140 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2475 5635 2480 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2461 5621 2475 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2447 5607 2461 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2433 5593 2447 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2419 5579 2433 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2405 5565 2419 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2391 5551 2405 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2377 5537 2391 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2363 5523 2377 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2349 5509 2363 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2335 5495 2349 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2321 5481 2335 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2307 5467 2321 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2293 5453 2307 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2279 5439 2293 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2265 5425 2279 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2251 5411 2265 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2237 5397 2251 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2223 5383 2237 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2209 5369 2223 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2195 5355 2209 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2181 5341 2195 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2167 5327 2181 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2153 5313 2167 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2139 5299 2153 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2125 5285 2139 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2111 5271 2125 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2097 5257 2111 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2083 5243 2097 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2069 5229 2083 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2055 5215 2069 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2041 5201 2055 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2027 5187 2041 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 2013 5173 2027 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1999 5159 2013 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1985 5145 1999 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1971 5131 1985 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1957 5117 1971 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1943 5103 1957 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1929 5089 1943 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1915 5075 1929 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1901 5061 1915 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1887 5047 1901 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1873 5033 1887 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1859 5019 1873 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1845 5005 1859 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1831 4991 1845 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1817 4977 1831 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1803 4963 1817 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1789 4949 1803 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1775 4935 1789 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1761 4921 1775 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1747 4907 1761 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1733 4893 1747 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 1719 4879 1733 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 513 4879 1719 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 201 509 4879 513 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 197 495 4879 509 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 183 481 4879 495 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 169 467 4879 481 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 155 453 4879 467 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 141 439 4879 453 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 127 425 4879 439 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 113 411 4879 425 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal2 s 99 0 4879 411 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6389 19275 7379 19305 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6389 18620 7379 19275 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6389 18598 7379 18620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6367 18568 7379 18598 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6359 19305 7379 19335 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6337 18538 7379 18568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6329 19335 7379 19365 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6307 18508 7379 18538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6299 19365 7379 19395 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6277 18478 7379 18508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6269 19395 7379 19425 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6239 19425 7379 19455 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6209 19455 7379 19485 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6179 19485 7379 19515 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6149 19515 7379 19545 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6119 19545 7379 19575 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6089 19575 7379 19605 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6059 19605 7379 19635 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6029 19635 7379 19665 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5999 19665 7379 19695 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5969 19695 7379 19725 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5939 19725 7379 19755 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5909 19755 7379 19785 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5879 19785 7379 19815 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5849 19815 7379 19845 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5819 19845 7379 19875 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5789 19875 7379 19905 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5759 19905 7379 19935 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5729 19935 7379 19965 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5699 19965 7379 19979 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5685 19979 7349 20009 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5655 20009 7319 20039 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5625 20039 7289 20069 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5595 20069 7259 20099 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5565 20099 7229 20129 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5535 20129 7199 20159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5505 20159 7169 20189 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5475 20189 7139 20219 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5445 20219 7109 20249 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5415 20249 7079 20279 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5385 20279 7049 20309 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5355 20309 7019 20339 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5325 20339 6989 20369 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5295 20369 6959 20399 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5265 20399 6929 20429 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5235 20429 6899 20459 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5205 20459 6880 20478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 35070 7364 40000 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 35052 7346 35070 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 35022 7316 35052 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34992 7286 35022 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34962 7256 34992 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34932 7226 34962 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34902 7196 34932 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34872 7166 34902 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34842 7136 34872 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34812 7106 34842 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34782 7076 34812 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34752 7046 34782 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34722 7016 34752 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34692 6986 34722 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34662 6956 34692 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34632 6926 34662 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34602 6896 34632 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34572 6866 34602 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34542 6836 34572 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34512 6806 34542 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34482 6776 34512 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34452 6746 34482 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34422 6716 34452 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34392 6686 34422 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34362 6656 34392 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34332 6626 34362 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34302 6596 34332 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34272 6566 34302 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34242 6536 34272 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34212 6506 34242 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34182 6476 34212 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34152 6446 34182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34122 6416 34152 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34092 6386 34122 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20972 6386 34092 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20958 6386 20972 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20928 6400 20958 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20898 6430 20928 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20868 6460 20898 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20838 6490 20868 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20808 6520 20838 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20778 6550 20808 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20748 6580 20778 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20718 6610 20748 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20688 6640 20718 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20658 6670 20688 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20628 6700 20658 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20598 6730 20628 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20568 6760 20598 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20538 6790 20568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20508 6820 20538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20478 6850 20508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5179 18078 7379 18108 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5179 0 7379 18078 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5149 18108 7379 18138 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5119 18138 7379 18168 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5089 18168 7379 18198 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5059 18198 7379 18228 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5029 18228 7379 18258 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4999 18258 7379 18288 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4969 18288 7379 18318 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4939 18318 7379 18348 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4909 18348 7379 18378 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4879 18378 7379 18408 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4849 18408 7379 18438 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4819 18438 7379 18468 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4789 18468 7379 18478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4779 18478 6032 18493 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4764 18493 6017 18508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18791 5905 18821 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18620 5905 18791 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18598 5905 18620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18568 5927 18598 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18538 5957 18568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18508 5987 18538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4719 18821 5905 18851 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4689 18851 5905 18881 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4659 18881 5905 18911 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4629 18911 5905 18941 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4599 18941 5905 18971 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4569 18971 5905 19001 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4539 19001 5905 19031 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4509 19031 5905 19061 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4479 19061 5905 19091 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4449 19091 5905 19121 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4419 19121 5905 19151 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4389 19151 5905 19181 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4359 19181 5905 19211 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4329 19211 5905 19241 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4299 19241 5905 19271 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4269 19271 5905 19301 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4239 19301 5905 19331 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4209 19331 5875 19361 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4179 19361 5845 19391 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4149 19391 5815 19421 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4119 19421 5785 19451 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4089 19451 5755 19481 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4059 19481 5725 19511 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4029 19511 5695 19541 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3999 19541 5665 19571 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3969 19571 5635 19601 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3939 19601 5605 19631 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3909 19631 5575 19661 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3879 19661 5545 19691 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3849 19691 5515 19721 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3819 19721 5485 19751 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3789 19751 5455 19781 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3759 19781 5425 19811 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3729 19811 5395 19841 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3699 19841 5365 19871 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3669 19871 5335 19901 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3639 19901 5305 19931 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3609 19931 5275 19961 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3579 19961 5245 19991 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3549 19991 5215 20021 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3519 20021 5185 20051 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3489 20051 5155 20081 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3459 20081 5125 20111 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3429 20111 5095 20141 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3399 20141 5065 20171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3369 20171 5035 20201 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3339 20201 5005 20231 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3309 20231 4975 20261 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3279 20261 4945 20291 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3249 20291 4915 20321 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3219 20321 4885 20351 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3189 20351 4855 20381 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3159 20381 4825 20411 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3129 20411 4796 20440 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34604 5002 34634 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34528 5002 34604 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34516 4990 34528 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34486 4960 34516 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34456 4930 34486 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34426 4900 34456 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34396 4870 34426 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34366 4840 34396 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34336 4810 34366 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34306 4780 34336 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34276 4750 34306 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34246 4720 34276 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34216 4690 34246 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34186 4660 34216 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34156 4630 34186 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34126 4600 34156 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34096 4570 34126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34066 4540 34096 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34036 4510 34066 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34006 4480 34036 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33976 4450 34006 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33946 4420 33976 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33916 4390 33946 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33886 4360 33916 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33856 4330 33886 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33826 4300 33856 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20936 4300 33826 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20920 4300 20936 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20890 4316 20920 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20860 4346 20890 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20830 4376 20860 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20800 4406 20830 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20770 4436 20800 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20740 4466 20770 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20710 4496 20740 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20680 4526 20710 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20650 4556 20680 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20620 4586 20650 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20590 4616 20620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20560 4646 20590 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20530 4676 20560 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20500 4706 20530 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20470 4736 20500 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20440 4766 20470 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3070 34634 5002 34664 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3040 34664 5002 34694 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3010 34694 5002 34724 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2980 34724 5002 34754 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2950 34754 5002 34784 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2920 34784 5002 34814 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2890 34814 5002 34844 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2860 34844 5002 34874 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2830 34874 5002 34904 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2800 34904 5002 34934 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2770 34934 5002 34964 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2740 34964 5002 34994 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2710 34994 5002 35024 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2680 35024 5002 35054 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2650 35054 5002 35084 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2620 35084 5002 35114 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2590 35114 5002 35144 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2560 35144 5002 35174 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2530 35174 5002 35204 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2500 35204 5002 35234 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2470 35234 5002 35264 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2440 35264 5002 35294 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2410 35294 5002 35324 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2380 35324 5002 35354 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2350 35354 5002 35384 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2320 35384 5002 35414 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2290 35414 5002 35444 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2260 35444 5002 35474 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2230 35474 5002 35504 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2200 35504 5002 35534 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2170 35534 5002 35564 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2140 35564 5002 35594 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2110 35594 5002 35624 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2080 35624 5002 35654 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2050 35654 5002 35684 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2020 35684 5002 35714 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1990 35714 5002 35744 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1960 35744 5002 35774 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1930 35774 5002 35804 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1900 35804 5002 35834 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1870 35834 5002 35864 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1840 35864 5002 35894 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1810 35894 5002 35924 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1780 35924 5002 35954 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1750 35954 5002 35984 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1720 35984 5002 36014 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1690 36014 5002 36044 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1660 36044 5002 36074 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1630 36074 5002 36104 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1600 36104 5002 36134 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1570 36134 5002 36164 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1540 36164 5002 36194 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1510 36194 5002 36224 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1480 36224 5002 36254 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1450 36254 5002 36284 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1420 36284 5002 36314 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1390 36314 5002 36344 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1360 36344 5002 36374 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1330 36374 5002 36404 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1300 36404 5002 36434 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1270 36434 5002 36464 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1240 36464 5002 36494 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1210 36494 5002 36524 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1180 36524 5002 36554 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1150 36554 5002 36584 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1120 36584 5002 36614 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1090 36614 5002 36644 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1060 36644 5002 36674 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1030 36674 5002 36704 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 1000 36704 5002 36734 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 970 36734 5002 36764 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 940 36764 5002 36794 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 910 36794 5002 36824 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 880 36824 5002 36854 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 850 36854 5002 36884 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 820 36884 5002 36914 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 790 36914 5002 36944 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 760 36944 5002 36974 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 730 36974 5002 37004 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 700 37004 5002 37034 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 670 37034 5002 37064 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 640 37064 5002 37072 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 632 37072 5002 40000 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal4 s 0 1777 15000 2707 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 0 1797 15000 2687 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 0 407 15000 1497 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 0 427 15000 1477 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal4 s 0 2987 15000 3677 6 VDDA
port 10 nsew power bidirectional
rlabel metal5 s 0 3007 15000 3657 6 VDDA
port 10 nsew power bidirectional
rlabel metal4 s 0 3957 15000 4887 6 VDDIO
port 11 nsew power bidirectional
rlabel metal4 s 0 14007 15000 19000 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 0 3977 15000 4867 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 0 14007 15000 18997 6 VDDIO
port 11 nsew power bidirectional
rlabel metal4 s 0 12817 15000 13707 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel metal5 s 0 12837 15000 13687 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel metal4 s 0 7347 15000 8037 6 VSSA
port 13 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 13 nsew ground bidirectional
rlabel metal4 s 0 10329 15000 10565 6 VSSA
port 13 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 13 nsew ground bidirectional
rlabel metal5 s 0 7367 15000 8017 6 VSSA
port 13 nsew ground bidirectional
rlabel metal5 s 0 9547 15000 11347 6 VSSA
port 13 nsew ground bidirectional
rlabel metal4 s 0 8317 15000 9247 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 0 8337 15000 9227 6 VSSD
port 14 nsew ground bidirectional
rlabel metal4 s 0 35157 15000 40000 6 VSSIO
port 15 nsew ground bidirectional
rlabel metal4 s 0 5167 15000 6097 6 VSSIO
port 15 nsew ground bidirectional
rlabel metal5 s 0 35157 15000 40000 6 VSSIO
port 15 nsew ground bidirectional
rlabel metal5 s 0 5187 15000 6077 6 VSSIO
port 15 nsew ground bidirectional
rlabel metal4 s 0 11647 15000 12537 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal5 s 0 11667 15000 12517 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal4 s 0 6377 15000 7067 6 VSWITCH
port 17 nsew power bidirectional
rlabel metal5 s 0 6397 15000 7047 6 VSWITCH
port 17 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
