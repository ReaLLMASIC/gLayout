magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 967 226
<< mvnnmos >>
rect 0 0 180 200
rect 236 0 416 200
rect 472 0 652 200
rect 708 0 888 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 180 182 236 200
rect 180 148 191 182
rect 225 148 236 182
rect 180 114 236 148
rect 180 80 191 114
rect 225 80 236 114
rect 180 46 236 80
rect 180 12 191 46
rect 225 12 236 46
rect 180 0 236 12
rect 416 182 472 200
rect 416 148 427 182
rect 461 148 472 182
rect 416 114 472 148
rect 416 80 427 114
rect 461 80 472 114
rect 416 46 472 80
rect 416 12 427 46
rect 461 12 472 46
rect 416 0 472 12
rect 652 182 708 200
rect 652 148 663 182
rect 697 148 708 182
rect 652 114 708 148
rect 652 80 663 114
rect 697 80 708 114
rect 652 46 708 80
rect 652 12 663 46
rect 697 12 708 46
rect 652 0 708 12
rect 888 182 941 200
rect 888 148 899 182
rect 933 148 941 182
rect 888 114 941 148
rect 888 80 899 114
rect 933 80 941 114
rect 888 46 941 80
rect 888 12 899 46
rect 933 12 941 46
rect 888 0 941 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 191 148 225 182
rect 191 80 225 114
rect 191 12 225 46
rect 427 148 461 182
rect 427 80 461 114
rect 427 12 461 46
rect 663 148 697 182
rect 663 80 697 114
rect 663 12 697 46
rect 899 148 933 182
rect 899 80 933 114
rect 899 12 933 46
<< poly >>
rect 0 200 180 232
rect 236 200 416 232
rect 472 200 652 232
rect 708 200 888 232
rect 0 -32 180 0
rect 236 -32 416 0
rect 472 -32 652 0
rect 708 -32 888 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 191 182 225 198
rect 191 114 225 148
rect 191 46 225 80
rect 191 -4 225 12
rect 427 182 461 198
rect 427 114 461 148
rect 427 46 461 80
rect 427 -4 461 12
rect 663 182 697 198
rect 663 114 697 148
rect 663 46 697 80
rect 663 -4 697 12
rect 899 182 933 198
rect 899 114 933 148
rect 899 46 933 80
rect 899 -4 933 12
use DFL1sd2_CDNS_5595914180816  DFL1sd2_CDNS_5595914180816_0
timestamp 1701704242
transform 1 0 180 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_5595914180816  DFL1sd2_CDNS_5595914180816_1
timestamp 1701704242
transform 1 0 416 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_5595914180816  DFL1sd2_CDNS_5595914180816_2
timestamp 1701704242
transform 1 0 652 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5595914180815  DFL1sd_CDNS_5595914180815_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5595914180815  DFL1sd_CDNS_5595914180815_1
timestamp 1701704242
transform 1 0 888 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 916 97 916 97 0 FreeSans 300 0 0 0 S
flabel comment s 680 97 680 97 0 FreeSans 300 0 0 0 D
flabel comment s 444 97 444 97 0 FreeSans 300 0 0 0 S
flabel comment s 208 97 208 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 652088
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 649650
<< end >>
