magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 190 1034 2613 1767
rect 2161 994 2613 1034
<< poly >>
rect 309 1782 565 1798
rect 309 1748 357 1782
rect 391 1748 425 1782
rect 459 1748 493 1782
rect 527 1748 565 1782
rect 309 1726 565 1748
rect 621 1782 877 1798
rect 621 1748 669 1782
rect 703 1748 737 1782
rect 771 1748 805 1782
rect 839 1748 877 1782
rect 621 1726 877 1748
rect 1043 1782 1499 1798
rect 1043 1748 1087 1782
rect 1121 1748 1155 1782
rect 1189 1748 1223 1782
rect 1257 1748 1291 1782
rect 1325 1748 1359 1782
rect 1393 1748 1427 1782
rect 1461 1748 1499 1782
rect 1043 1700 1499 1748
rect 1555 1782 2011 1798
rect 1555 1748 1599 1782
rect 1633 1748 1667 1782
rect 1701 1748 1735 1782
rect 1769 1748 1803 1782
rect 1837 1748 1871 1782
rect 1905 1748 1939 1782
rect 1973 1748 2011 1782
rect 1555 1700 2011 1748
rect 2294 1736 2494 1752
rect 2294 1702 2310 1736
rect 2344 1702 2444 1736
rect 2478 1702 2494 1736
rect 2294 1686 2494 1702
rect 2280 1000 2480 1016
rect 2280 966 2296 1000
rect 2330 966 2430 1000
rect 2464 966 2480 1000
rect 2280 950 2480 966
rect 1164 802 1230 818
rect 1164 768 1180 802
rect 1214 768 1230 802
rect 1164 734 1230 768
rect 1164 700 1180 734
rect 1214 700 1230 734
rect 1164 684 1230 700
rect 1164 612 1230 628
rect 1164 578 1180 612
rect 1214 578 1230 612
rect 1164 531 1230 578
rect 1164 497 1180 531
rect 1214 497 1230 531
rect 1164 450 1230 497
rect 1164 416 1180 450
rect 1214 416 1230 450
rect 1164 369 1230 416
rect 1164 335 1180 369
rect 1214 335 1230 369
rect 1164 288 1230 335
rect 1164 254 1180 288
rect 1214 254 1230 288
rect 1164 206 1230 254
rect 1164 172 1180 206
rect 1214 172 1230 206
rect 1164 156 1230 172
<< polycont >>
rect 357 1748 391 1782
rect 425 1748 459 1782
rect 493 1748 527 1782
rect 669 1748 703 1782
rect 737 1748 771 1782
rect 805 1748 839 1782
rect 1087 1748 1121 1782
rect 1155 1748 1189 1782
rect 1223 1748 1257 1782
rect 1291 1748 1325 1782
rect 1359 1748 1393 1782
rect 1427 1748 1461 1782
rect 1599 1748 1633 1782
rect 1667 1748 1701 1782
rect 1735 1748 1769 1782
rect 1803 1748 1837 1782
rect 1871 1748 1905 1782
rect 1939 1748 1973 1782
rect 2310 1702 2344 1736
rect 2444 1702 2478 1736
rect 2296 966 2330 1000
rect 2430 966 2464 1000
rect 1180 768 1214 802
rect 1180 700 1214 734
rect 1180 578 1214 612
rect 1180 497 1214 531
rect 1180 416 1214 450
rect 1180 335 1214 369
rect 1180 254 1214 288
rect 1180 172 1214 206
<< locali >>
rect 341 1786 854 1788
rect 341 1782 615 1786
rect 341 1748 357 1782
rect 391 1748 425 1782
rect 459 1748 493 1782
rect 527 1752 615 1782
rect 649 1782 690 1786
rect 724 1782 764 1786
rect 798 1782 854 1786
rect 1117 1782 1170 1784
rect 1204 1782 1257 1784
rect 649 1752 669 1782
rect 724 1752 737 1782
rect 798 1752 805 1782
rect 527 1748 669 1752
rect 703 1748 737 1752
rect 771 1748 805 1752
rect 839 1748 855 1782
rect 1071 1750 1083 1782
rect 1071 1748 1087 1750
rect 1121 1748 1155 1782
rect 1204 1750 1223 1782
rect 1189 1748 1223 1750
rect 1291 1782 1344 1784
rect 1378 1782 1431 1784
rect 1629 1782 1682 1784
rect 1716 1782 1769 1784
rect 1257 1748 1291 1750
rect 1325 1750 1344 1782
rect 1325 1748 1359 1750
rect 1393 1748 1427 1782
rect 1465 1750 1477 1782
rect 1461 1748 1477 1750
rect 1583 1750 1595 1782
rect 1583 1748 1599 1750
rect 1633 1748 1667 1782
rect 1716 1750 1735 1782
rect 1701 1748 1735 1750
rect 1803 1782 1856 1784
rect 1890 1782 1943 1784
rect 1769 1748 1803 1750
rect 1837 1750 1856 1782
rect 1837 1748 1871 1750
rect 1905 1748 1939 1782
rect 1977 1750 1989 1782
rect 1973 1748 1989 1750
rect 2294 1735 2310 1736
rect 2110 1702 2310 1735
rect 2344 1702 2444 1736
rect 2478 1702 2494 1736
rect 2110 1696 2494 1702
rect 726 1629 764 1663
rect 1765 1629 1803 1663
rect 998 1475 1032 1529
rect 1510 1475 1544 1529
rect 2022 1475 2056 1529
rect 418 1339 456 1373
rect 1248 1339 1286 1373
rect 264 1182 298 1236
rect 576 1182 610 1236
rect 888 1182 922 1236
rect 2110 1087 2177 1696
rect 1149 1053 1161 1087
rect 1195 1053 1233 1087
rect 2093 1053 2131 1087
rect 2165 1053 2177 1087
rect 2223 1056 2303 1658
rect 2505 1475 2539 1529
rect 2491 1182 2525 1236
rect 180 815 227 849
rect 261 815 308 849
rect 342 815 389 849
rect 423 815 469 849
rect 503 815 549 849
rect 583 815 629 849
rect 663 815 709 849
rect 743 815 789 849
rect 1149 802 1214 1053
rect 2326 1000 2434 1018
rect 1149 768 1180 802
rect 1149 734 1214 768
rect 1149 700 1180 734
rect 1149 684 1214 700
rect 1282 955 1320 989
rect 2280 984 2292 1000
rect 2280 966 2296 984
rect 2330 966 2430 1000
rect 2468 984 2480 1000
rect 2464 966 2480 984
rect 419 638 462 672
rect 496 638 539 672
rect 573 638 616 672
rect 650 638 693 672
rect 727 638 770 672
rect 804 638 847 672
rect 881 638 924 672
rect 958 638 1001 672
rect 1035 638 1078 672
rect 1248 628 1293 955
rect 1180 612 1293 628
rect 1214 578 1293 612
rect 1180 531 1293 578
rect 1214 497 1293 531
rect 674 463 712 497
rect 746 463 784 497
rect 1180 450 1293 497
rect 1214 416 1293 450
rect 1180 369 1293 416
rect 1214 335 1293 369
rect 392 286 430 320
rect 464 286 502 320
rect 536 286 574 320
rect 608 286 646 320
rect 680 286 718 320
rect 752 286 790 320
rect 824 286 862 320
rect 896 286 934 320
rect 968 286 1006 320
rect 1040 286 1078 320
rect 1180 288 1293 335
rect 1214 254 1293 288
rect 1180 206 1293 254
rect 1214 172 1293 206
rect 1180 156 1293 172
rect 180 111 221 145
rect 255 111 296 145
rect 330 111 371 145
rect 405 111 446 145
rect 480 111 520 145
rect 554 111 594 145
rect 628 111 668 145
rect 702 111 742 145
rect 776 111 816 145
rect 850 111 890 145
rect 924 111 964 145
rect 998 111 1038 145
<< viali >>
rect 615 1752 649 1786
rect 690 1782 724 1786
rect 764 1782 798 1786
rect 1083 1782 1117 1784
rect 1170 1782 1204 1784
rect 690 1752 703 1782
rect 703 1752 724 1782
rect 764 1752 771 1782
rect 771 1752 798 1782
rect 1083 1750 1087 1782
rect 1087 1750 1117 1782
rect 1170 1750 1189 1782
rect 1189 1750 1204 1782
rect 1257 1750 1291 1784
rect 1344 1782 1378 1784
rect 1431 1782 1465 1784
rect 1595 1782 1629 1784
rect 1682 1782 1716 1784
rect 1344 1750 1359 1782
rect 1359 1750 1378 1782
rect 1431 1750 1461 1782
rect 1461 1750 1465 1782
rect 1595 1750 1599 1782
rect 1599 1750 1629 1782
rect 1682 1750 1701 1782
rect 1701 1750 1716 1782
rect 1769 1750 1803 1784
rect 1856 1782 1890 1784
rect 1943 1782 1977 1784
rect 1856 1750 1871 1782
rect 1871 1750 1890 1782
rect 1943 1750 1973 1782
rect 1973 1750 1977 1782
rect 692 1629 726 1663
rect 764 1629 798 1663
rect 1731 1629 1765 1663
rect 1803 1629 1837 1663
rect 998 1529 1032 1563
rect 998 1441 1032 1475
rect 1510 1529 1544 1563
rect 1510 1441 1544 1475
rect 2022 1529 2056 1563
rect 2022 1441 2056 1475
rect 384 1339 418 1373
rect 456 1339 490 1373
rect 1214 1339 1248 1373
rect 1286 1339 1320 1373
rect 264 1236 298 1270
rect 264 1148 298 1182
rect 576 1236 610 1270
rect 576 1148 610 1182
rect 888 1236 922 1270
rect 888 1148 922 1182
rect 1161 1053 1195 1087
rect 1233 1053 1267 1087
rect 2059 1053 2093 1087
rect 2131 1053 2165 1087
rect 2505 1529 2539 1563
rect 2505 1441 2539 1475
rect 2491 1236 2525 1270
rect 2491 1148 2525 1182
rect 146 815 180 849
rect 227 815 261 849
rect 308 815 342 849
rect 389 815 423 849
rect 469 815 503 849
rect 549 815 583 849
rect 629 815 663 849
rect 709 815 743 849
rect 789 815 823 849
rect 2292 1000 2326 1018
rect 2434 1000 2468 1018
rect 1248 955 1282 989
rect 1320 955 1354 989
rect 2292 984 2296 1000
rect 2296 984 2326 1000
rect 2434 984 2464 1000
rect 2464 984 2468 1000
rect 385 638 419 672
rect 462 638 496 672
rect 539 638 573 672
rect 616 638 650 672
rect 693 638 727 672
rect 770 638 804 672
rect 847 638 881 672
rect 924 638 958 672
rect 1001 638 1035 672
rect 1078 638 1112 672
rect 640 463 674 497
rect 712 463 746 497
rect 784 463 818 497
rect 358 286 392 320
rect 430 286 464 320
rect 502 286 536 320
rect 574 286 608 320
rect 646 286 680 320
rect 718 286 752 320
rect 790 286 824 320
rect 862 286 896 320
rect 934 286 968 320
rect 1006 286 1040 320
rect 1078 286 1112 320
rect 146 111 180 145
rect 221 111 255 145
rect 296 111 330 145
rect 371 111 405 145
rect 446 111 480 145
rect 520 111 554 145
rect 594 111 628 145
rect 668 111 702 145
rect 742 111 776 145
rect 816 111 850 145
rect 890 111 924 145
rect 964 111 998 145
rect 1038 111 1072 145
<< metal1 >>
rect 678 1792 684 1795
rect 603 1786 684 1792
rect 603 1752 615 1786
rect 649 1752 684 1786
rect 603 1746 684 1752
rect 678 1743 684 1746
rect 736 1743 750 1795
rect 802 1792 808 1795
rect 802 1746 810 1792
rect 1071 1784 1477 1790
rect 1071 1750 1083 1784
rect 1117 1750 1170 1784
rect 1204 1750 1257 1784
rect 1291 1750 1344 1784
rect 1378 1750 1431 1784
rect 1465 1750 1477 1784
rect 802 1743 808 1746
rect 1071 1744 1477 1750
rect 1583 1784 1989 1790
rect 1583 1750 1595 1784
rect 1629 1750 1682 1784
rect 1716 1750 1769 1784
rect 1803 1750 1856 1784
rect 1890 1750 1943 1784
rect 1977 1750 1989 1784
rect 1583 1744 1989 1750
rect 679 1663 1849 1688
rect 679 1629 692 1663
rect 726 1629 764 1663
rect 798 1629 1731 1663
rect 1765 1629 1803 1663
rect 1837 1629 1849 1663
rect 679 1604 1849 1629
rect 990 1563 2546 1575
rect 990 1529 998 1563
rect 1032 1529 1510 1563
rect 1544 1529 2022 1563
rect 2056 1529 2505 1563
rect 2539 1529 2546 1563
rect 990 1475 2546 1529
rect 990 1441 998 1475
rect 1032 1441 1510 1475
rect 1544 1441 2022 1475
rect 2056 1441 2505 1475
rect 2539 1441 2546 1475
rect 990 1429 2546 1441
rect 371 1373 1332 1398
rect 371 1339 384 1373
rect 418 1339 456 1373
rect 490 1339 1214 1373
rect 1248 1339 1286 1373
rect 1320 1339 1332 1373
rect 371 1314 1332 1339
rect 258 1270 2534 1282
rect 258 1236 264 1270
rect 298 1236 576 1270
rect 610 1236 888 1270
rect 922 1236 2491 1270
rect 2525 1236 2534 1270
rect 258 1182 2534 1236
rect 258 1148 264 1182
rect 298 1148 576 1182
rect 610 1148 888 1182
rect 922 1148 2491 1182
rect 2525 1148 2534 1182
rect 258 1136 2534 1148
tri 555 1097 594 1136 ne
rect 594 1101 676 1136
tri 676 1101 711 1136 nw
tri 555 855 594 894 se
rect 594 855 672 1101
tri 672 1097 676 1101 nw
rect 1149 1087 2180 1101
rect 701 1014 707 1066
rect 759 1014 782 1066
rect 834 1053 1032 1066
tri 1032 1053 1045 1066 sw
rect 1149 1053 1161 1087
rect 1195 1053 1233 1087
rect 1267 1053 2059 1087
rect 2093 1053 2131 1087
rect 2165 1053 2180 1087
rect 834 1040 1045 1053
tri 1045 1040 1058 1053 sw
rect 1149 1040 2180 1053
rect 834 1024 1058 1040
tri 1058 1024 1074 1040 sw
rect 834 1018 1074 1024
tri 1074 1018 1080 1024 sw
tri 2274 1018 2280 1024 se
rect 2280 1018 2480 1024
rect 834 1014 1080 1018
tri 1080 1014 1084 1018 sw
tri 2270 1014 2274 1018 se
rect 2274 1014 2292 1018
tri 1004 1001 1017 1014 ne
rect 1017 1001 1084 1014
tri 1084 1001 1097 1014 sw
tri 2257 1001 2270 1014 se
rect 2270 1001 2292 1014
tri 1017 995 1023 1001 ne
rect 1023 995 2292 1001
tri 1023 989 1029 995 ne
rect 1029 989 2292 995
tri 1029 986 1032 989 ne
rect 1032 986 1248 989
tri 1032 955 1063 986 ne
rect 1063 955 1248 986
rect 1282 955 1320 989
rect 1354 984 2292 989
rect 2326 984 2434 1018
rect 2468 984 2480 1018
rect 1354 955 2480 984
tri 1063 949 1069 955 ne
rect 1069 949 2480 955
tri 672 855 711 894 sw
rect 134 849 679 855
rect 731 849 743 855
rect 795 849 835 855
rect 134 815 146 849
rect 180 815 227 849
rect 261 815 308 849
rect 342 815 389 849
rect 423 815 469 849
rect 503 815 549 849
rect 583 815 629 849
rect 663 815 679 849
rect 823 815 835 849
rect 134 809 679 815
rect 673 803 679 809
rect 731 803 743 815
rect 795 809 835 815
rect 795 803 801 809
rect 373 672 1124 678
rect 373 638 385 672
rect 419 638 462 672
rect 496 638 539 672
rect 573 638 616 672
rect 650 638 693 672
rect 727 638 770 672
rect 804 638 847 672
rect 881 638 924 672
rect 958 638 1001 672
rect 1035 638 1078 672
rect 1112 638 1124 672
rect 373 632 1124 638
rect 673 503 679 506
rect 628 497 679 503
rect 731 497 743 506
rect 795 503 801 506
rect 795 497 830 503
rect 628 463 640 497
rect 674 463 679 497
rect 818 463 830 497
rect 628 457 679 463
rect 673 454 679 457
rect 731 454 743 463
rect 795 457 830 463
rect 795 454 801 457
rect 871 326 1124 632
rect 346 320 1124 326
rect 346 286 358 320
rect 392 286 430 320
rect 464 286 502 320
rect 536 286 574 320
rect 608 286 646 320
rect 680 286 718 320
rect 752 286 790 320
rect 824 286 862 320
rect 896 286 934 320
rect 968 286 1006 320
rect 1040 286 1078 320
rect 1112 286 1124 320
rect 346 280 1124 286
rect 673 151 679 154
rect 134 145 679 151
rect 731 145 743 154
rect 795 151 801 154
rect 795 145 1084 151
rect 134 111 146 145
rect 180 111 221 145
rect 255 111 296 145
rect 330 111 371 145
rect 405 111 446 145
rect 480 111 520 145
rect 554 111 594 145
rect 628 111 668 145
rect 731 111 742 145
rect 795 111 816 145
rect 850 111 890 145
rect 924 111 964 145
rect 998 111 1038 145
rect 1072 111 1084 145
rect 134 105 679 111
rect 673 102 679 105
rect 731 102 743 111
rect 795 105 1084 111
rect 795 102 801 105
<< via1 >>
rect 684 1786 736 1795
rect 684 1752 690 1786
rect 690 1752 724 1786
rect 724 1752 736 1786
rect 684 1743 736 1752
rect 750 1786 802 1795
rect 750 1752 764 1786
rect 764 1752 798 1786
rect 798 1752 802 1786
rect 750 1743 802 1752
rect 707 1014 759 1066
rect 782 1014 834 1066
rect 679 849 731 855
rect 743 849 795 855
rect 679 815 709 849
rect 709 815 731 849
rect 743 815 789 849
rect 789 815 795 849
rect 679 803 731 815
rect 743 803 795 815
rect 679 497 731 506
rect 743 497 795 506
rect 679 463 712 497
rect 712 463 731 497
rect 743 463 746 497
rect 746 463 784 497
rect 784 463 795 497
rect 679 454 731 463
rect 743 454 795 463
rect 679 145 731 154
rect 743 145 795 154
rect 679 111 702 145
rect 702 111 731 145
rect 743 111 776 145
rect 776 111 795 145
rect 679 102 731 111
rect 743 102 795 111
<< metal2 >>
rect 678 1743 684 1795
rect 736 1743 750 1795
rect 802 1743 808 1795
rect 701 1066 768 1743
tri 768 1066 818 1116 sw
rect 701 1014 707 1066
rect 759 1014 782 1066
rect 834 1014 840 1066
tri 1608 862 1630 884 sw
rect 673 803 679 855
rect 731 803 743 855
rect 795 803 801 855
rect 673 506 801 803
rect 673 454 679 506
rect 731 454 743 506
rect 795 454 801 506
rect 673 154 801 454
rect 673 102 679 154
rect 731 102 743 154
rect 795 102 801 154
use nfet_CDNS_524688791851405  nfet_CDNS_524688791851405_0
timestamp 1701704242
transform 0 1 138 -1 0 804
box -79 -26 727 1026
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_0
timestamp 1701704242
transform -1 0 565 0 -1 1700
box -119 -66 375 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_1
timestamp 1701704242
transform 1 0 621 0 -1 1700
box -119 -66 375 666
use pfet_CDNS_524688791851406  pfet_CDNS_524688791851406_0
timestamp 1701704242
transform 1 0 2280 0 1 1048
box -119 -66 319 366
use pfet_CDNS_524688791851407  pfet_CDNS_524688791851407_0
timestamp 1701704242
transform -1 0 2494 0 -1 1654
box -119 -66 319 266
use pfet_CDNS_524688791851408  pfet_CDNS_524688791851408_0
timestamp 1701704242
transform -1 0 1499 0 -1 1674
box -119 -66 575 666
use pfet_CDNS_524688791851408  pfet_CDNS_524688791851408_1
timestamp 1701704242
transform 1 0 1555 0 -1 1674
box -119 -66 575 666
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1701704242
transform 0 -1 855 -1 0 1798
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1701704242
transform 0 -1 543 -1 0 1798
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1701704242
transform 0 -1 1477 -1 0 1798
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_1
timestamp 1701704242
transform 0 -1 1989 -1 0 1798
box 0 0 1 1
<< labels >>
flabel metal1 s 2380 1204 2429 1248 3 FreeSans 300 0 0 0 pd_h
port 1 nsew
flabel metal1 s 951 446 997 485 3 FreeSans 300 0 0 0 vgnd_io
port 2 nsew
flabel metal1 s 1315 1472 1391 1542 3 FreeSans 300 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 1250 1044 1308 1096 3 FreeSans 300 0 0 0 pden_h_n
port 4 nsew
flabel metal1 s 1733 1748 1809 1782 3 FreeSans 300 0 0 0 en_fast_n<1>
port 5 nsew
flabel metal1 s 1256 1748 1323 1782 3 FreeSans 300 0 0 0 en_fast_n<0>
port 6 nsew
flabel metal1 s 769 1014 835 1066 3 FreeSans 300 0 0 0 drvlo_h_n
port 7 nsew
<< properties >>
string GDS_END 87842474
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87828236
string path 16.825 3.200 20.025 3.200 
<< end >>
