magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 59 800 865 1568
<< pwell >>
rect 278 76 732 728
<< mvnmos >>
rect 357 102 477 702
rect 533 102 653 702
<< mvpmos >>
rect 178 866 278 1466
rect 334 866 434 1466
rect 490 866 590 1466
rect 646 866 746 1466
<< mvndiff >>
rect 304 624 357 702
rect 304 590 312 624
rect 346 590 357 624
rect 304 556 357 590
rect 304 522 312 556
rect 346 522 357 556
rect 304 488 357 522
rect 304 454 312 488
rect 346 454 357 488
rect 304 420 357 454
rect 304 386 312 420
rect 346 386 357 420
rect 304 352 357 386
rect 304 318 312 352
rect 346 318 357 352
rect 304 284 357 318
rect 304 250 312 284
rect 346 250 357 284
rect 304 216 357 250
rect 304 182 312 216
rect 346 182 357 216
rect 304 148 357 182
rect 304 114 312 148
rect 346 114 357 148
rect 304 102 357 114
rect 477 624 533 702
rect 477 590 488 624
rect 522 590 533 624
rect 477 556 533 590
rect 477 522 488 556
rect 522 522 533 556
rect 477 488 533 522
rect 477 454 488 488
rect 522 454 533 488
rect 477 420 533 454
rect 477 386 488 420
rect 522 386 533 420
rect 477 352 533 386
rect 477 318 488 352
rect 522 318 533 352
rect 477 284 533 318
rect 477 250 488 284
rect 522 250 533 284
rect 477 216 533 250
rect 477 182 488 216
rect 522 182 533 216
rect 477 148 533 182
rect 477 114 488 148
rect 522 114 533 148
rect 477 102 533 114
rect 653 624 706 702
rect 653 590 664 624
rect 698 590 706 624
rect 653 556 706 590
rect 653 522 664 556
rect 698 522 706 556
rect 653 488 706 522
rect 653 454 664 488
rect 698 454 706 488
rect 653 420 706 454
rect 653 386 664 420
rect 698 386 706 420
rect 653 352 706 386
rect 653 318 664 352
rect 698 318 706 352
rect 653 284 706 318
rect 653 250 664 284
rect 698 250 706 284
rect 653 216 706 250
rect 653 182 664 216
rect 698 182 706 216
rect 653 148 706 182
rect 653 114 664 148
rect 698 114 706 148
rect 653 102 706 114
<< mvpdiff >>
rect 125 1454 178 1466
rect 125 1420 133 1454
rect 167 1420 178 1454
rect 125 1386 178 1420
rect 125 1352 133 1386
rect 167 1352 178 1386
rect 125 1318 178 1352
rect 125 1284 133 1318
rect 167 1284 178 1318
rect 125 1250 178 1284
rect 125 1216 133 1250
rect 167 1216 178 1250
rect 125 1182 178 1216
rect 125 1148 133 1182
rect 167 1148 178 1182
rect 125 1114 178 1148
rect 125 1080 133 1114
rect 167 1080 178 1114
rect 125 1046 178 1080
rect 125 1012 133 1046
rect 167 1012 178 1046
rect 125 978 178 1012
rect 125 944 133 978
rect 167 944 178 978
rect 125 866 178 944
rect 278 1454 334 1466
rect 278 1420 289 1454
rect 323 1420 334 1454
rect 278 1386 334 1420
rect 278 1352 289 1386
rect 323 1352 334 1386
rect 278 1318 334 1352
rect 278 1284 289 1318
rect 323 1284 334 1318
rect 278 1250 334 1284
rect 278 1216 289 1250
rect 323 1216 334 1250
rect 278 1182 334 1216
rect 278 1148 289 1182
rect 323 1148 334 1182
rect 278 1114 334 1148
rect 278 1080 289 1114
rect 323 1080 334 1114
rect 278 1046 334 1080
rect 278 1012 289 1046
rect 323 1012 334 1046
rect 278 978 334 1012
rect 278 944 289 978
rect 323 944 334 978
rect 278 866 334 944
rect 434 1454 490 1466
rect 434 1420 445 1454
rect 479 1420 490 1454
rect 434 1386 490 1420
rect 434 1352 445 1386
rect 479 1352 490 1386
rect 434 1318 490 1352
rect 434 1284 445 1318
rect 479 1284 490 1318
rect 434 1250 490 1284
rect 434 1216 445 1250
rect 479 1216 490 1250
rect 434 1182 490 1216
rect 434 1148 445 1182
rect 479 1148 490 1182
rect 434 1114 490 1148
rect 434 1080 445 1114
rect 479 1080 490 1114
rect 434 1046 490 1080
rect 434 1012 445 1046
rect 479 1012 490 1046
rect 434 978 490 1012
rect 434 944 445 978
rect 479 944 490 978
rect 434 866 490 944
rect 590 1454 646 1466
rect 590 1420 601 1454
rect 635 1420 646 1454
rect 590 1386 646 1420
rect 590 1352 601 1386
rect 635 1352 646 1386
rect 590 1318 646 1352
rect 590 1284 601 1318
rect 635 1284 646 1318
rect 590 1250 646 1284
rect 590 1216 601 1250
rect 635 1216 646 1250
rect 590 1182 646 1216
rect 590 1148 601 1182
rect 635 1148 646 1182
rect 590 1114 646 1148
rect 590 1080 601 1114
rect 635 1080 646 1114
rect 590 1046 646 1080
rect 590 1012 601 1046
rect 635 1012 646 1046
rect 590 978 646 1012
rect 590 944 601 978
rect 635 944 646 978
rect 590 866 646 944
rect 746 1454 799 1466
rect 746 1420 757 1454
rect 791 1420 799 1454
rect 746 1386 799 1420
rect 746 1352 757 1386
rect 791 1352 799 1386
rect 746 1318 799 1352
rect 746 1284 757 1318
rect 791 1284 799 1318
rect 746 1250 799 1284
rect 746 1216 757 1250
rect 791 1216 799 1250
rect 746 1182 799 1216
rect 746 1148 757 1182
rect 791 1148 799 1182
rect 746 1114 799 1148
rect 746 1080 757 1114
rect 791 1080 799 1114
rect 746 1046 799 1080
rect 746 1012 757 1046
rect 791 1012 799 1046
rect 746 978 799 1012
rect 746 944 757 978
rect 791 944 799 978
rect 746 866 799 944
<< mvndiffc >>
rect 312 590 346 624
rect 312 522 346 556
rect 312 454 346 488
rect 312 386 346 420
rect 312 318 346 352
rect 312 250 346 284
rect 312 182 346 216
rect 312 114 346 148
rect 488 590 522 624
rect 488 522 522 556
rect 488 454 522 488
rect 488 386 522 420
rect 488 318 522 352
rect 488 250 522 284
rect 488 182 522 216
rect 488 114 522 148
rect 664 590 698 624
rect 664 522 698 556
rect 664 454 698 488
rect 664 386 698 420
rect 664 318 698 352
rect 664 250 698 284
rect 664 182 698 216
rect 664 114 698 148
<< mvpdiffc >>
rect 133 1420 167 1454
rect 133 1352 167 1386
rect 133 1284 167 1318
rect 133 1216 167 1250
rect 133 1148 167 1182
rect 133 1080 167 1114
rect 133 1012 167 1046
rect 133 944 167 978
rect 289 1420 323 1454
rect 289 1352 323 1386
rect 289 1284 323 1318
rect 289 1216 323 1250
rect 289 1148 323 1182
rect 289 1080 323 1114
rect 289 1012 323 1046
rect 289 944 323 978
rect 445 1420 479 1454
rect 445 1352 479 1386
rect 445 1284 479 1318
rect 445 1216 479 1250
rect 445 1148 479 1182
rect 445 1080 479 1114
rect 445 1012 479 1046
rect 445 944 479 978
rect 601 1420 635 1454
rect 601 1352 635 1386
rect 601 1284 635 1318
rect 601 1216 635 1250
rect 601 1148 635 1182
rect 601 1080 635 1114
rect 601 1012 635 1046
rect 601 944 635 978
rect 757 1420 791 1454
rect 757 1352 791 1386
rect 757 1284 791 1318
rect 757 1216 791 1250
rect 757 1148 791 1182
rect 757 1080 791 1114
rect 757 1012 791 1046
rect 757 944 791 978
<< poly >>
rect 178 1548 434 1568
rect 178 1514 233 1548
rect 267 1514 301 1548
rect 335 1514 369 1548
rect 403 1514 434 1548
rect 178 1492 434 1514
rect 178 1466 278 1492
rect 334 1466 434 1492
rect 490 1548 746 1568
rect 490 1514 526 1548
rect 560 1514 594 1548
rect 628 1514 662 1548
rect 696 1514 746 1548
rect 490 1492 746 1514
rect 490 1466 590 1492
rect 646 1466 746 1492
rect 178 840 278 866
rect 334 840 434 866
rect 490 840 590 866
rect 646 840 746 866
rect 117 785 434 840
rect 117 751 137 785
rect 171 751 205 785
rect 239 751 434 785
rect 117 728 434 751
rect 533 785 746 840
rect 533 751 553 785
rect 587 751 621 785
rect 655 751 689 785
rect 723 751 746 785
rect 533 728 746 751
rect 357 702 477 728
rect 533 702 653 728
rect 357 76 477 102
rect 335 54 477 76
rect 335 20 355 54
rect 389 20 423 54
rect 457 20 477 54
rect 335 0 477 20
rect 533 76 653 102
rect 533 54 677 76
rect 533 20 555 54
rect 589 20 623 54
rect 657 20 677 54
rect 533 0 677 20
<< polycont >>
rect 233 1514 267 1548
rect 301 1514 335 1548
rect 369 1514 403 1548
rect 526 1514 560 1548
rect 594 1514 628 1548
rect 662 1514 696 1548
rect 137 751 171 785
rect 205 751 239 785
rect 553 751 587 785
rect 621 751 655 785
rect 689 751 723 785
rect 355 20 389 54
rect 423 20 457 54
rect 555 20 589 54
rect 623 20 657 54
<< locali >>
rect 217 1514 233 1548
rect 267 1514 301 1548
rect 335 1514 369 1548
rect 403 1514 419 1548
rect 510 1514 526 1548
rect 560 1514 594 1548
rect 628 1514 662 1548
rect 696 1514 712 1548
rect 133 1454 167 1470
rect 133 1386 167 1420
rect 289 1454 323 1470
rect 289 1386 323 1420
rect 133 1318 167 1352
rect 285 1352 289 1374
rect 445 1454 479 1470
rect 445 1386 479 1420
rect 285 1340 323 1352
rect 133 1250 167 1284
rect 133 1182 167 1216
rect 289 1318 323 1340
rect 289 1250 323 1284
rect 289 1182 323 1216
rect 133 1142 149 1148
rect 183 1142 221 1176
rect 445 1318 479 1352
rect 445 1250 479 1284
rect 445 1182 479 1216
rect 133 1114 167 1142
rect 133 1046 167 1080
rect 133 978 167 1012
rect 133 928 167 944
rect 289 1114 323 1148
rect 443 1148 445 1176
rect 601 1454 635 1470
rect 601 1386 635 1420
rect 601 1318 635 1352
rect 601 1250 635 1284
rect 601 1182 635 1216
rect 479 1148 481 1176
rect 443 1142 481 1148
rect 757 1454 791 1470
rect 757 1386 791 1420
rect 757 1318 791 1352
rect 757 1250 791 1284
rect 757 1182 791 1216
rect 289 1046 323 1080
rect 289 978 323 1012
rect 121 751 137 785
rect 171 751 205 785
rect 239 751 255 785
rect 289 708 323 944
rect 445 1114 479 1142
rect 445 1046 479 1080
rect 445 978 479 1012
rect 445 928 479 944
rect 601 1114 635 1148
rect 703 1142 741 1176
rect 775 1142 791 1148
rect 601 1046 635 1056
rect 601 978 635 984
rect 757 1114 791 1142
rect 757 1046 791 1080
rect 757 978 791 1012
rect 757 928 791 944
rect 537 751 553 785
rect 587 751 621 785
rect 655 751 689 785
rect 723 751 739 785
rect 289 674 522 708
rect 312 624 346 640
rect 312 576 346 590
rect 312 504 346 522
rect 312 432 346 454
rect 312 352 346 386
rect 312 284 346 318
rect 312 216 346 250
rect 312 148 346 182
rect 312 98 346 114
rect 488 624 522 674
rect 488 556 522 590
rect 488 488 522 522
rect 488 420 522 454
rect 488 352 522 386
rect 488 284 522 318
rect 488 216 522 250
rect 488 148 522 182
rect 488 98 522 114
rect 664 624 698 640
rect 664 576 698 590
rect 664 504 698 522
rect 664 432 698 454
rect 664 352 698 386
rect 664 284 698 318
rect 664 216 698 250
rect 664 148 698 182
rect 664 98 698 114
rect 339 20 355 54
rect 389 20 423 54
rect 457 20 473 54
rect 539 20 555 54
rect 589 20 623 54
rect 657 20 673 54
<< viali >>
rect 251 1340 285 1374
rect 323 1340 357 1374
rect 149 1148 167 1176
rect 167 1148 183 1176
rect 149 1142 183 1148
rect 221 1142 255 1176
rect 409 1142 443 1176
rect 481 1142 515 1176
rect 669 1142 703 1176
rect 741 1148 757 1176
rect 757 1148 775 1176
rect 741 1142 775 1148
rect 601 1080 635 1090
rect 601 1056 635 1080
rect 601 1012 635 1018
rect 601 984 635 1012
rect 601 944 635 946
rect 601 912 635 944
rect 312 556 346 576
rect 312 542 346 556
rect 312 488 346 504
rect 312 470 346 488
rect 312 420 346 432
rect 312 398 346 420
rect 664 556 698 576
rect 664 542 698 556
rect 664 488 698 504
rect 664 470 698 488
rect 664 420 698 432
rect 664 398 698 420
<< metal1 >>
rect 239 1374 369 1380
rect 239 1340 251 1374
rect 285 1340 323 1374
rect 357 1340 369 1374
rect 239 1334 369 1340
rect 137 1176 787 1182
rect 137 1142 149 1176
rect 183 1142 221 1176
rect 255 1142 409 1176
rect 443 1142 481 1176
rect 515 1142 669 1176
rect 703 1142 741 1176
rect 775 1142 787 1176
rect 137 1136 787 1142
rect 0 1090 872 1108
rect 0 1056 601 1090
rect 635 1056 872 1090
rect 0 1018 872 1056
rect 0 984 601 1018
rect 635 984 872 1018
rect 0 946 872 984
rect 0 912 601 946
rect 635 912 872 946
rect 0 906 872 912
rect 0 576 872 582
rect 0 542 312 576
rect 346 542 664 576
rect 698 542 872 576
rect 0 504 872 542
rect 0 470 312 504
rect 346 470 664 504
rect 698 470 872 504
rect 0 432 872 470
rect 0 398 312 432
rect 346 398 664 432
rect 698 398 872 432
rect 0 380 872 398
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_0
timestamp 1701704242
transform 1 0 357 0 1 102
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_1
timestamp 1701704242
transform -1 0 653 0 1 102
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808364  sky130_fd_pr__pfet_01v8__example_55959141808364_0
timestamp 1701704242
transform 1 0 490 0 -1 1466
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808364  sky130_fd_pr__pfet_01v8__example_55959141808364_1
timestamp 1701704242
transform 1 0 178 0 -1 1466
box -1 0 257 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1701704242
transform 1 0 251 0 1 1340
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1701704242
transform -1 0 255 0 1 1142
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1701704242
transform -1 0 515 0 1 1142
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1701704242
transform -1 0 775 0 1 1142
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1701704242
transform 1 0 312 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1701704242
transform 1 0 664 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_2
timestamp 1701704242
transform 1 0 601 0 1 912
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1701704242
transform 0 1 121 1 0 735
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1701704242
transform 0 -1 673 1 0 4
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1701704242
transform 0 -1 473 1 0 4
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1701704242
transform 0 1 537 1 0 735
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_1
timestamp 1701704242
transform 0 1 510 -1 0 1564
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_2
timestamp 1701704242
transform 0 1 217 1 0 1498
box 0 0 1 1
<< labels >>
flabel locali s 133 751 167 785 3 FreeSans 300 0 0 0 DRVLO_H_N
port 1 nsew
flabel locali s 705 751 739 785 3 FreeSans 300 180 0 0 PDEN_H_N
port 2 nsew
flabel metal1 s 0 906 42 1108 6 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 0 380 42 582 7 FreeSans 300 0 0 0 VGND_IO
port 4 nsew
flabel metal1 s 830 906 872 1108 7 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 830 380 872 582 7 FreeSans 300 180 0 0 VGND_IO
port 4 nsew
flabel metal1 s 239 1334 285 1380 7 FreeSans 300 0 0 0 PD_H
port 5 nsew
flabel comment s 544 1164 544 1164 0 FreeSans 200 0 0 0 INT
<< properties >>
string GDS_END 67939712
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 67936156
<< end >>
