magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -36 -36 89 4036
<< pdiff >>
rect 0 3922 53 4000
rect 0 3888 11 3922
rect 45 3888 53 3922
rect 0 3854 53 3888
rect 0 3820 11 3854
rect 45 3820 53 3854
rect 0 3786 53 3820
rect 0 3752 11 3786
rect 45 3752 53 3786
rect 0 3718 53 3752
rect 0 3684 11 3718
rect 45 3684 53 3718
rect 0 3650 53 3684
rect 0 3616 11 3650
rect 45 3616 53 3650
rect 0 3582 53 3616
rect 0 3548 11 3582
rect 45 3548 53 3582
rect 0 3514 53 3548
rect 0 3480 11 3514
rect 45 3480 53 3514
rect 0 3446 53 3480
rect 0 3412 11 3446
rect 45 3412 53 3446
rect 0 3378 53 3412
rect 0 3344 11 3378
rect 45 3344 53 3378
rect 0 3310 53 3344
rect 0 3276 11 3310
rect 45 3276 53 3310
rect 0 3242 53 3276
rect 0 3208 11 3242
rect 45 3208 53 3242
rect 0 3174 53 3208
rect 0 3140 11 3174
rect 45 3140 53 3174
rect 0 3106 53 3140
rect 0 3072 11 3106
rect 45 3072 53 3106
rect 0 3038 53 3072
rect 0 3004 11 3038
rect 45 3004 53 3038
rect 0 2970 53 3004
rect 0 2936 11 2970
rect 45 2936 53 2970
rect 0 2902 53 2936
rect 0 2868 11 2902
rect 45 2868 53 2902
rect 0 2834 53 2868
rect 0 2800 11 2834
rect 45 2800 53 2834
rect 0 2766 53 2800
rect 0 2732 11 2766
rect 45 2732 53 2766
rect 0 2698 53 2732
rect 0 2664 11 2698
rect 45 2664 53 2698
rect 0 2630 53 2664
rect 0 2596 11 2630
rect 45 2596 53 2630
rect 0 2562 53 2596
rect 0 2528 11 2562
rect 45 2528 53 2562
rect 0 2494 53 2528
rect 0 2460 11 2494
rect 45 2460 53 2494
rect 0 2426 53 2460
rect 0 2392 11 2426
rect 45 2392 53 2426
rect 0 2358 53 2392
rect 0 2324 11 2358
rect 45 2324 53 2358
rect 0 2290 53 2324
rect 0 2256 11 2290
rect 45 2256 53 2290
rect 0 2222 53 2256
rect 0 2188 11 2222
rect 45 2188 53 2222
rect 0 2154 53 2188
rect 0 2120 11 2154
rect 45 2120 53 2154
rect 0 2086 53 2120
rect 0 2052 11 2086
rect 45 2052 53 2086
rect 0 2018 53 2052
rect 0 1984 11 2018
rect 45 1984 53 2018
rect 0 1950 53 1984
rect 0 1916 11 1950
rect 45 1916 53 1950
rect 0 1882 53 1916
rect 0 1848 11 1882
rect 45 1848 53 1882
rect 0 1814 53 1848
rect 0 1780 11 1814
rect 45 1780 53 1814
rect 0 1746 53 1780
rect 0 1712 11 1746
rect 45 1712 53 1746
rect 0 1678 53 1712
rect 0 1644 11 1678
rect 45 1644 53 1678
rect 0 1610 53 1644
rect 0 1576 11 1610
rect 45 1576 53 1610
rect 0 1542 53 1576
rect 0 1508 11 1542
rect 45 1508 53 1542
rect 0 1474 53 1508
rect 0 1440 11 1474
rect 45 1440 53 1474
rect 0 1406 53 1440
rect 0 1372 11 1406
rect 45 1372 53 1406
rect 0 1338 53 1372
rect 0 1304 11 1338
rect 45 1304 53 1338
rect 0 1270 53 1304
rect 0 1236 11 1270
rect 45 1236 53 1270
rect 0 1202 53 1236
rect 0 1168 11 1202
rect 45 1168 53 1202
rect 0 1134 53 1168
rect 0 1100 11 1134
rect 45 1100 53 1134
rect 0 1066 53 1100
rect 0 1032 11 1066
rect 45 1032 53 1066
rect 0 998 53 1032
rect 0 964 11 998
rect 45 964 53 998
rect 0 930 53 964
rect 0 896 11 930
rect 45 896 53 930
rect 0 862 53 896
rect 0 828 11 862
rect 45 828 53 862
rect 0 794 53 828
rect 0 760 11 794
rect 45 760 53 794
rect 0 726 53 760
rect 0 692 11 726
rect 45 692 53 726
rect 0 658 53 692
rect 0 624 11 658
rect 45 624 53 658
rect 0 590 53 624
rect 0 556 11 590
rect 45 556 53 590
rect 0 522 53 556
rect 0 488 11 522
rect 45 488 53 522
rect 0 454 53 488
rect 0 420 11 454
rect 45 420 53 454
rect 0 386 53 420
rect 0 352 11 386
rect 45 352 53 386
rect 0 318 53 352
rect 0 284 11 318
rect 45 284 53 318
rect 0 250 53 284
rect 0 216 11 250
rect 45 216 53 250
rect 0 182 53 216
rect 0 148 11 182
rect 45 148 53 182
rect 0 114 53 148
rect 0 80 11 114
rect 45 80 53 114
rect 0 46 53 80
rect 0 12 11 46
rect 45 12 53 46
rect 0 0 53 12
<< pdiffc >>
rect 11 3888 45 3922
rect 11 3820 45 3854
rect 11 3752 45 3786
rect 11 3684 45 3718
rect 11 3616 45 3650
rect 11 3548 45 3582
rect 11 3480 45 3514
rect 11 3412 45 3446
rect 11 3344 45 3378
rect 11 3276 45 3310
rect 11 3208 45 3242
rect 11 3140 45 3174
rect 11 3072 45 3106
rect 11 3004 45 3038
rect 11 2936 45 2970
rect 11 2868 45 2902
rect 11 2800 45 2834
rect 11 2732 45 2766
rect 11 2664 45 2698
rect 11 2596 45 2630
rect 11 2528 45 2562
rect 11 2460 45 2494
rect 11 2392 45 2426
rect 11 2324 45 2358
rect 11 2256 45 2290
rect 11 2188 45 2222
rect 11 2120 45 2154
rect 11 2052 45 2086
rect 11 1984 45 2018
rect 11 1916 45 1950
rect 11 1848 45 1882
rect 11 1780 45 1814
rect 11 1712 45 1746
rect 11 1644 45 1678
rect 11 1576 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1474
rect 11 1372 45 1406
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 3922 45 3938
rect 11 3854 45 3888
rect 11 3786 45 3820
rect 11 3718 45 3752
rect 11 3650 45 3684
rect 11 3582 45 3616
rect 11 3514 45 3548
rect 11 3446 45 3480
rect 11 3378 45 3412
rect 11 3310 45 3344
rect 11 3242 45 3276
rect 11 3174 45 3208
rect 11 3106 45 3140
rect 11 3038 45 3072
rect 11 2970 45 3004
rect 11 2902 45 2936
rect 11 2834 45 2868
rect 11 2766 45 2800
rect 11 2698 45 2732
rect 11 2630 45 2664
rect 11 2562 45 2596
rect 11 2494 45 2528
rect 11 2426 45 2460
rect 11 2358 45 2392
rect 11 2290 45 2324
rect 11 2222 45 2256
rect 11 2154 45 2188
rect 11 2086 45 2120
rect 11 2018 45 2052
rect 11 1950 45 1984
rect 11 1882 45 1916
rect 11 1814 45 1848
rect 11 1746 45 1780
rect 11 1678 45 1712
rect 11 1610 45 1644
rect 11 1542 45 1576
rect 11 1474 45 1508
rect 11 1406 45 1440
rect 11 1338 45 1372
rect 11 1270 45 1304
rect 11 1202 45 1236
rect 11 1134 45 1168
rect 11 1066 45 1100
rect 11 998 45 1032
rect 11 930 45 964
rect 11 862 45 896
rect 11 794 45 828
rect 11 726 45 760
rect 11 658 45 692
rect 11 590 45 624
rect 11 522 45 556
rect 11 454 45 488
rect 11 386 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 216
rect 11 114 45 148
rect 11 46 45 80
rect 11 -4 45 12
<< properties >>
string GDS_END 95600970
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95596998
<< end >>
