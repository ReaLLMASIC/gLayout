magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal2 >>
rect -1157 428 1157 437
rect -1157 -428 -1148 428
rect 1148 -428 1157 428
rect -1157 -437 1157 -428
<< via2 >>
rect -1148 -428 1148 428
<< metal3 >>
rect -1153 428 1153 433
rect -1153 -428 -1148 428
rect 1148 -428 1153 428
rect -1153 -433 1153 -428
<< properties >>
string GDS_END 34505700
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34485152
<< end >>
