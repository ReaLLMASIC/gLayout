magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 3375 266
<< mvpmos >>
rect 0 0 1600 200
rect 1656 0 3256 200
<< mvpdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 1600 182 1656 200
rect 1600 148 1611 182
rect 1645 148 1656 182
rect 1600 114 1656 148
rect 1600 80 1611 114
rect 1645 80 1656 114
rect 1600 46 1656 80
rect 1600 12 1611 46
rect 1645 12 1656 46
rect 1600 0 1656 12
rect 3256 182 3309 200
rect 3256 148 3267 182
rect 3301 148 3309 182
rect 3256 114 3309 148
rect 3256 80 3267 114
rect 3301 80 3309 114
rect 3256 46 3309 80
rect 3256 12 3267 46
rect 3301 12 3309 46
rect 3256 0 3309 12
<< mvpdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 1611 148 1645 182
rect 1611 80 1645 114
rect 1611 12 1645 46
rect 3267 148 3301 182
rect 3267 80 3301 114
rect 3267 12 3301 46
<< poly >>
rect 0 200 1600 232
rect 1656 200 3256 232
rect 0 -32 1600 0
rect 1656 -32 3256 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 1611 182 1645 198
rect 1611 114 1645 148
rect 1611 46 1645 80
rect 1611 -4 1645 12
rect 3267 182 3301 198
rect 3267 114 3301 148
rect 3267 46 3301 80
rect 3267 -4 3301 12
use DFL1sd2_CDNS_52468879185419  DFL1sd2_CDNS_52468879185419_0
timestamp 1701704242
transform 1 0 1600 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_1
timestamp 1701704242
transform 1 0 3256 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 1628 97 1628 97 0 FreeSans 300 0 0 0 D
flabel comment s 3284 97 3284 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 6079304
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6077792
<< end >>
