magic
tech sky130B
timestamp 1701704242
<< nwell >>
rect -18 -18 535 59
<< nsubdiff >>
rect 0 29 517 41
rect 0 12 12 29
rect 29 12 46 29
rect 63 12 80 29
rect 97 12 114 29
rect 131 12 148 29
rect 165 12 182 29
rect 199 12 216 29
rect 233 12 250 29
rect 267 12 284 29
rect 301 12 318 29
rect 335 12 352 29
rect 369 12 386 29
rect 403 12 420 29
rect 437 12 454 29
rect 471 12 488 29
rect 505 12 517 29
rect 0 0 517 12
<< nsubdiffcont >>
rect 12 12 29 29
rect 46 12 63 29
rect 80 12 97 29
rect 114 12 131 29
rect 148 12 165 29
rect 182 12 199 29
rect 216 12 233 29
rect 250 12 267 29
rect 284 12 301 29
rect 318 12 335 29
rect 352 12 369 29
rect 386 12 403 29
rect 420 12 437 29
rect 454 12 471 29
rect 488 12 505 29
<< locali >>
rect 12 29 505 37
rect 29 12 46 29
rect 63 12 80 29
rect 97 12 114 29
rect 131 12 148 29
rect 165 12 182 29
rect 199 12 216 29
rect 233 12 250 29
rect 267 12 284 29
rect 301 12 318 29
rect 335 12 352 29
rect 369 12 386 29
rect 403 12 420 29
rect 437 12 454 29
rect 471 12 488 29
rect 12 4 505 12
<< properties >>
string GDS_END 85830430
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85829210
<< end >>
