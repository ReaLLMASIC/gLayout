magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1513 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 166 47 196 177
rect 252 47 282 177
rect 338 47 368 177
rect 424 47 454 177
rect 510 47 540 177
rect 596 47 626 177
rect 684 47 714 177
rect 776 47 806 177
rect 862 47 892 177
rect 948 47 978 177
rect 1032 47 1062 177
rect 1116 47 1146 177
rect 1200 47 1230 177
rect 1284 47 1314 177
rect 1378 47 1408 177
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 252 297 282 497
rect 338 297 368 497
rect 424 297 454 497
rect 510 297 540 497
rect 596 297 626 497
rect 682 297 712 497
rect 776 297 806 497
rect 862 297 892 497
rect 948 297 978 497
rect 1032 297 1062 497
rect 1116 297 1146 497
rect 1200 297 1230 497
rect 1284 297 1314 497
rect 1368 297 1398 497
<< ndiff >>
rect 27 157 80 177
rect 27 123 35 157
rect 69 123 80 157
rect 27 47 80 123
rect 110 89 166 177
rect 110 55 121 89
rect 155 55 166 89
rect 110 47 166 55
rect 196 159 252 177
rect 196 125 207 159
rect 241 125 252 159
rect 196 47 252 125
rect 282 89 338 177
rect 282 55 293 89
rect 327 55 338 89
rect 282 47 338 55
rect 368 159 424 177
rect 368 125 379 159
rect 413 125 424 159
rect 368 47 424 125
rect 454 89 510 177
rect 454 55 465 89
rect 499 55 510 89
rect 454 47 510 55
rect 540 159 596 177
rect 540 125 551 159
rect 585 125 596 159
rect 540 47 596 125
rect 626 89 684 177
rect 626 55 637 89
rect 671 55 684 89
rect 626 47 684 55
rect 714 116 776 177
rect 714 82 727 116
rect 761 82 776 116
rect 714 47 776 82
rect 806 163 862 177
rect 806 129 817 163
rect 851 129 862 163
rect 806 47 862 129
rect 892 90 948 177
rect 892 56 903 90
rect 937 56 948 90
rect 892 47 948 56
rect 978 47 1032 177
rect 1062 90 1116 177
rect 1062 56 1072 90
rect 1106 56 1116 90
rect 1062 47 1116 56
rect 1146 162 1200 177
rect 1146 128 1156 162
rect 1190 128 1200 162
rect 1146 47 1200 128
rect 1230 90 1284 177
rect 1230 56 1240 90
rect 1274 56 1284 90
rect 1230 47 1284 56
rect 1314 47 1378 177
rect 1408 96 1487 177
rect 1408 62 1419 96
rect 1453 62 1487 96
rect 1408 47 1487 62
<< pdiff >>
rect 27 485 80 497
rect 27 451 35 485
rect 69 451 80 485
rect 27 383 80 451
rect 27 349 35 383
rect 69 349 80 383
rect 27 297 80 349
rect 110 422 166 497
rect 110 388 121 422
rect 155 388 166 422
rect 110 297 166 388
rect 196 489 252 497
rect 196 455 207 489
rect 241 455 252 489
rect 196 297 252 455
rect 282 449 338 497
rect 282 415 293 449
rect 327 415 338 449
rect 282 297 338 415
rect 368 405 424 497
rect 368 371 379 405
rect 413 371 424 405
rect 368 297 424 371
rect 454 489 510 497
rect 454 455 465 489
rect 499 455 510 489
rect 454 297 510 455
rect 540 405 596 497
rect 540 371 551 405
rect 585 371 596 405
rect 540 297 596 371
rect 626 489 682 497
rect 626 455 637 489
rect 671 455 682 489
rect 626 297 682 455
rect 712 489 776 497
rect 712 455 727 489
rect 761 455 776 489
rect 712 297 776 455
rect 806 405 862 497
rect 806 371 817 405
rect 851 371 862 405
rect 806 297 862 371
rect 892 489 948 497
rect 892 455 903 489
rect 937 455 948 489
rect 892 297 948 455
rect 978 405 1032 497
rect 978 371 988 405
rect 1022 371 1032 405
rect 978 297 1032 371
rect 1062 489 1116 497
rect 1062 455 1072 489
rect 1106 455 1116 489
rect 1062 297 1116 455
rect 1146 405 1200 497
rect 1146 371 1156 405
rect 1190 371 1200 405
rect 1146 297 1200 371
rect 1230 489 1284 497
rect 1230 455 1240 489
rect 1274 455 1284 489
rect 1230 297 1284 455
rect 1314 405 1368 497
rect 1314 371 1324 405
rect 1358 371 1368 405
rect 1314 297 1368 371
rect 1398 489 1533 497
rect 1398 455 1487 489
rect 1521 455 1533 489
rect 1398 297 1533 455
<< ndiffc >>
rect 35 123 69 157
rect 121 55 155 89
rect 207 125 241 159
rect 293 55 327 89
rect 379 125 413 159
rect 465 55 499 89
rect 551 125 585 159
rect 637 55 671 89
rect 727 82 761 116
rect 817 129 851 163
rect 903 56 937 90
rect 1072 56 1106 90
rect 1156 128 1190 162
rect 1240 56 1274 90
rect 1419 62 1453 96
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 121 388 155 422
rect 207 455 241 489
rect 293 415 327 449
rect 379 371 413 405
rect 465 455 499 489
rect 551 371 585 405
rect 637 455 671 489
rect 727 455 761 489
rect 817 371 851 405
rect 903 455 937 489
rect 988 371 1022 405
rect 1072 455 1106 489
rect 1156 371 1190 405
rect 1240 455 1274 489
rect 1324 371 1358 405
rect 1487 455 1521 489
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 252 497 282 523
rect 338 497 368 523
rect 424 497 454 523
rect 510 497 540 523
rect 596 497 626 523
rect 682 497 712 523
rect 776 497 806 523
rect 862 497 892 523
rect 948 497 978 523
rect 1032 497 1062 523
rect 1116 497 1146 523
rect 1200 497 1230 523
rect 1284 497 1314 523
rect 1368 497 1398 523
rect 80 265 110 297
rect 166 265 196 297
rect 252 265 282 297
rect 80 249 282 265
rect 80 215 96 249
rect 130 215 164 249
rect 198 215 232 249
rect 266 215 282 249
rect 80 199 282 215
rect 80 177 110 199
rect 166 177 196 199
rect 252 177 282 199
rect 338 275 368 297
rect 424 275 454 297
rect 510 275 540 297
rect 596 275 626 297
rect 338 249 626 275
rect 682 265 712 297
rect 776 265 806 297
rect 862 265 892 297
rect 948 265 978 297
rect 338 215 357 249
rect 391 215 425 249
rect 459 215 493 249
rect 527 215 561 249
rect 595 215 626 249
rect 338 199 626 215
rect 668 249 734 265
rect 668 215 684 249
rect 718 215 734 249
rect 668 199 734 215
rect 776 249 978 265
rect 776 215 792 249
rect 826 215 860 249
rect 894 215 928 249
rect 962 215 978 249
rect 776 199 978 215
rect 338 177 368 199
rect 424 177 454 199
rect 510 177 540 199
rect 596 177 626 199
rect 684 177 714 199
rect 776 177 806 199
rect 862 177 892 199
rect 948 177 978 199
rect 1032 265 1062 297
rect 1116 265 1146 297
rect 1200 265 1230 297
rect 1284 265 1314 297
rect 1368 265 1398 297
rect 1032 249 1314 265
rect 1032 215 1102 249
rect 1136 215 1170 249
rect 1204 215 1238 249
rect 1272 215 1314 249
rect 1032 199 1314 215
rect 1356 249 1410 265
rect 1356 215 1366 249
rect 1400 215 1410 249
rect 1356 199 1410 215
rect 1032 177 1062 199
rect 1116 177 1146 199
rect 1200 177 1230 199
rect 1284 177 1314 199
rect 1378 177 1408 199
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 684 21 714 47
rect 776 21 806 47
rect 862 21 892 47
rect 948 21 978 47
rect 1032 21 1062 47
rect 1116 21 1146 47
rect 1200 21 1230 47
rect 1284 21 1314 47
rect 1378 21 1408 47
<< polycont >>
rect 96 215 130 249
rect 164 215 198 249
rect 232 215 266 249
rect 357 215 391 249
rect 425 215 459 249
rect 493 215 527 249
rect 561 215 595 249
rect 684 215 718 249
rect 792 215 826 249
rect 860 215 894 249
rect 928 215 962 249
rect 1102 215 1136 249
rect 1170 215 1204 249
rect 1238 215 1272 249
rect 1366 215 1400 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 485 77 527
rect 18 451 35 485
rect 69 451 77 485
rect 191 489 257 527
rect 191 455 207 489
rect 241 455 257 489
rect 291 489 687 493
rect 291 455 465 489
rect 499 455 637 489
rect 671 455 687 489
rect 723 489 777 527
rect 723 455 727 489
rect 761 455 777 489
rect 887 489 953 527
rect 887 455 903 489
rect 937 455 953 489
rect 1056 489 1122 527
rect 1056 455 1072 489
rect 1106 455 1122 489
rect 1224 489 1291 527
rect 1224 455 1240 489
rect 1274 455 1291 489
rect 1471 489 1537 527
rect 1471 455 1487 489
rect 1521 455 1537 489
rect 18 383 77 451
rect 291 449 327 455
rect 18 349 35 383
rect 69 349 77 383
rect 111 422 155 438
rect 111 388 121 422
rect 291 421 293 449
rect 155 415 293 421
rect 723 439 777 455
rect 155 388 327 415
rect 111 387 327 388
rect 361 405 694 421
rect 809 405 1536 421
rect 111 372 155 387
rect 361 371 379 405
rect 413 371 551 405
rect 585 371 817 405
rect 851 371 988 405
rect 1022 371 1156 405
rect 1190 371 1324 405
rect 1358 371 1536 405
rect 18 333 77 349
rect 193 303 726 337
rect 193 266 282 303
rect 80 249 282 266
rect 80 215 96 249
rect 130 215 164 249
rect 198 215 232 249
rect 266 215 282 249
rect 341 249 636 269
rect 341 215 357 249
rect 391 215 425 249
rect 459 215 493 249
rect 527 215 561 249
rect 595 215 636 249
rect 670 249 726 303
rect 852 303 1400 337
rect 852 282 995 303
rect 670 215 684 249
rect 718 215 726 249
rect 670 199 726 215
rect 760 249 995 282
rect 760 215 792 249
rect 826 215 860 249
rect 894 215 928 249
rect 962 215 995 249
rect 1074 249 1288 269
rect 1074 215 1102 249
rect 1136 215 1170 249
rect 1204 215 1238 249
rect 1272 215 1288 249
rect 1366 249 1400 303
rect 760 199 995 215
rect 1366 199 1400 215
rect 1434 268 1536 371
rect 31 173 359 181
rect 31 159 626 173
rect 1434 165 1470 268
rect 31 157 207 159
rect 31 123 35 157
rect 69 125 207 157
rect 241 139 379 159
rect 241 125 248 139
rect 355 125 379 139
rect 413 125 551 159
rect 585 125 767 159
rect 801 129 817 163
rect 851 162 1234 163
rect 851 129 1156 162
rect 801 128 1156 129
rect 1190 128 1234 162
rect 801 127 1234 128
rect 1313 131 1470 165
rect 69 123 71 125
rect 31 107 71 123
rect 205 119 248 125
rect 105 55 121 89
rect 155 55 171 89
rect 205 85 214 119
rect 721 116 767 125
rect 293 89 327 105
rect 105 17 171 55
rect 293 17 327 55
rect 449 55 465 89
rect 499 55 515 89
rect 449 17 515 55
rect 621 55 637 89
rect 671 55 687 89
rect 621 17 687 55
rect 721 82 727 116
rect 761 91 767 116
rect 761 90 984 91
rect 1313 90 1347 131
rect 761 82 903 90
rect 721 56 903 82
rect 937 56 984 90
rect 721 51 984 56
rect 1056 56 1072 90
rect 1106 56 1240 90
rect 1274 56 1347 90
rect 1396 62 1419 96
rect 1453 85 1502 96
rect 1453 62 1536 85
rect 1056 54 1347 56
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 214 85 248 119
rect 1502 85 1536 119
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 202 119 260 125
rect 202 85 214 119
rect 248 116 260 119
rect 1490 119 1548 125
rect 1490 116 1502 119
rect 248 88 1502 116
rect 248 85 260 88
rect 202 79 260 85
rect 1490 85 1502 88
rect 1536 85 1548 119
rect 1490 79 1548 85
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 214 289 248 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 950 289 984 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1226 221 1260 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1502 357 1536 391 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o211ai_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 793882
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 783862
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 7.820 0.000 
<< end >>
