magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -79 -26 179 176
<< mvnmos >>
rect 0 0 100 150
<< mvndiff >>
rect -53 114 0 150
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 100 114 153 150
rect 100 80 111 114
rect 145 80 153 114
rect 100 46 153 80
rect 100 12 111 46
rect 145 12 153 46
rect 100 0 153 12
<< mvndiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 150 100 182
rect 0 -32 100 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 80
rect -45 -4 -11 12
rect 111 114 145 130
rect 111 46 145 80
rect 111 -4 145 12
use DFL1sd_CDNS_52468879185245  DFL1sd_CDNS_52468879185245_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185245  DFL1sd_CDNS_52468879185245_1
timestamp 1701704242
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
flabel comment s 128 63 128 63 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 7563920
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7563034
<< end >>
