magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -68 -26 1068 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 1000 50 1042 66
rect 1034 16 1042 50
rect 1000 0 1042 16
<< ndiffc >>
rect -34 16 0 50
rect 1000 16 1034 50
<< ndiffres >>
rect 0 0 1000 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 1000 50 1034 66
rect 1000 0 1034 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 1 0 992 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 96448098
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96447596
<< end >>
