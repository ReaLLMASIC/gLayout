magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< poly >>
rect 0 4594 11146 4610
rect 0 4560 34 4594
rect 68 4560 102 4594
rect 136 4560 170 4594
rect 204 4560 238 4594
rect 272 4560 306 4594
rect 340 4560 374 4594
rect 408 4560 442 4594
rect 476 4560 510 4594
rect 544 4560 578 4594
rect 612 4560 646 4594
rect 680 4560 714 4594
rect 748 4560 782 4594
rect 816 4560 850 4594
rect 884 4560 918 4594
rect 952 4560 986 4594
rect 1020 4560 1054 4594
rect 1088 4560 1122 4594
rect 1156 4560 1190 4594
rect 1224 4560 1258 4594
rect 1292 4560 1326 4594
rect 1360 4560 1394 4594
rect 1428 4560 1462 4594
rect 1496 4560 1530 4594
rect 1564 4560 1598 4594
rect 1632 4560 1666 4594
rect 1700 4560 1734 4594
rect 1768 4560 1802 4594
rect 1836 4560 1870 4594
rect 1904 4560 1938 4594
rect 1972 4560 2006 4594
rect 2040 4560 2074 4594
rect 2108 4560 2142 4594
rect 2176 4560 2210 4594
rect 2244 4560 2278 4594
rect 2312 4560 2346 4594
rect 2380 4560 2414 4594
rect 2448 4560 2482 4594
rect 2516 4560 2550 4594
rect 2584 4560 2618 4594
rect 2652 4560 2686 4594
rect 2720 4560 2754 4594
rect 2788 4560 2822 4594
rect 2856 4560 2890 4594
rect 2924 4560 2958 4594
rect 2992 4560 3026 4594
rect 3060 4560 3094 4594
rect 3128 4560 3162 4594
rect 3196 4560 3230 4594
rect 3264 4560 3298 4594
rect 3332 4560 3366 4594
rect 3400 4560 3434 4594
rect 3468 4560 3502 4594
rect 3536 4560 3570 4594
rect 3604 4560 3638 4594
rect 3672 4560 3706 4594
rect 3740 4560 3774 4594
rect 3808 4560 3842 4594
rect 3876 4560 3910 4594
rect 3944 4560 3978 4594
rect 4012 4560 4046 4594
rect 4080 4560 4114 4594
rect 4148 4560 4182 4594
rect 4216 4560 4250 4594
rect 4284 4560 4318 4594
rect 4352 4560 4386 4594
rect 4420 4560 4454 4594
rect 4488 4560 4522 4594
rect 4556 4560 4590 4594
rect 4624 4560 4658 4594
rect 4692 4560 4726 4594
rect 4760 4560 4794 4594
rect 4828 4560 4862 4594
rect 4896 4560 4930 4594
rect 4964 4560 4998 4594
rect 5032 4560 5066 4594
rect 5100 4560 5134 4594
rect 5168 4560 5202 4594
rect 5236 4560 5270 4594
rect 5304 4560 5338 4594
rect 5372 4560 5406 4594
rect 5440 4560 5474 4594
rect 5508 4560 5542 4594
rect 5576 4560 5610 4594
rect 5644 4560 5678 4594
rect 5712 4560 5746 4594
rect 5780 4560 5814 4594
rect 5848 4560 5882 4594
rect 5916 4560 5950 4594
rect 5984 4560 6018 4594
rect 6052 4560 6086 4594
rect 6120 4560 6154 4594
rect 6188 4560 6222 4594
rect 6256 4560 6290 4594
rect 6324 4560 6358 4594
rect 6392 4560 6426 4594
rect 6460 4560 6494 4594
rect 6528 4560 6562 4594
rect 6596 4560 6630 4594
rect 6664 4560 6698 4594
rect 6732 4560 6766 4594
rect 6800 4560 6834 4594
rect 6868 4560 6902 4594
rect 6936 4560 6970 4594
rect 7004 4560 7038 4594
rect 7072 4560 7106 4594
rect 7140 4560 7174 4594
rect 7208 4560 7242 4594
rect 7276 4560 7310 4594
rect 7344 4560 7378 4594
rect 7412 4560 7446 4594
rect 7480 4560 7514 4594
rect 7548 4560 7582 4594
rect 7616 4560 7650 4594
rect 7684 4560 7718 4594
rect 7752 4560 7786 4594
rect 7820 4560 7854 4594
rect 7888 4560 7922 4594
rect 7956 4560 7990 4594
rect 8024 4560 8058 4594
rect 8092 4560 8126 4594
rect 8160 4560 8194 4594
rect 8228 4560 8262 4594
rect 8296 4560 8330 4594
rect 8364 4560 8398 4594
rect 8432 4560 8466 4594
rect 8500 4560 8534 4594
rect 8568 4560 8602 4594
rect 8636 4560 8670 4594
rect 8704 4560 8738 4594
rect 8772 4560 8806 4594
rect 8840 4560 8874 4594
rect 8908 4560 8942 4594
rect 8976 4560 9010 4594
rect 9044 4560 9078 4594
rect 9112 4560 9146 4594
rect 9180 4560 9214 4594
rect 9248 4560 9282 4594
rect 9316 4560 9350 4594
rect 9384 4560 9418 4594
rect 9452 4560 9486 4594
rect 9520 4560 9554 4594
rect 9588 4560 9622 4594
rect 9656 4560 9690 4594
rect 9724 4560 9758 4594
rect 9792 4560 9826 4594
rect 9860 4560 9894 4594
rect 9928 4560 9962 4594
rect 9996 4560 10030 4594
rect 10064 4560 10098 4594
rect 10132 4560 10166 4594
rect 10200 4560 10234 4594
rect 10268 4560 10302 4594
rect 10336 4560 10370 4594
rect 10404 4560 10438 4594
rect 10472 4560 10506 4594
rect 10540 4560 10574 4594
rect 10608 4560 10642 4594
rect 10676 4560 10710 4594
rect 10744 4560 10778 4594
rect 10812 4560 10846 4594
rect 10880 4560 10914 4594
rect 10948 4560 10982 4594
rect 11016 4560 11050 4594
rect 11084 4560 11146 4594
rect 0 4544 11146 4560
rect 0 108 30 4544
rect 72 66 102 4502
rect 144 108 174 4544
rect 216 66 246 4502
rect 288 108 318 4544
rect 360 66 390 4502
rect 432 108 462 4544
rect 504 66 534 4502
rect 576 108 606 4544
rect 648 66 678 4502
rect 720 108 750 4544
rect 792 66 822 4502
rect 864 108 894 4544
rect 936 66 966 4502
rect 1008 108 1038 4544
rect 1080 66 1110 4502
rect 1152 108 1182 4544
rect 1224 66 1254 4502
rect 1296 108 1326 4544
rect 1368 66 1398 4502
rect 1440 108 1470 4544
rect 1512 66 1542 4502
rect 1584 108 1614 4544
rect 1656 66 1686 4502
rect 1728 108 1758 4544
rect 1800 66 1830 4502
rect 1872 108 1902 4544
rect 1944 66 1974 4502
rect 2016 108 2046 4544
rect 2088 66 2118 4502
rect 2160 108 2190 4544
rect 2232 66 2262 4502
rect 2304 108 2334 4544
rect 2376 66 2406 4502
rect 2448 108 2478 4544
rect 2520 66 2550 4502
rect 2592 108 2622 4544
rect 2664 66 2694 4502
rect 2736 108 2766 4544
rect 2808 66 2838 4502
rect 2880 108 2910 4544
rect 2952 66 2982 4502
rect 3024 108 3054 4544
rect 3096 66 3126 4502
rect 3168 108 3198 4544
rect 3240 66 3270 4502
rect 3312 108 3342 4544
rect 3384 66 3414 4502
rect 3456 108 3486 4544
rect 3528 66 3558 4502
rect 3600 108 3630 4544
rect 3672 66 3702 4502
rect 3744 108 3774 4544
rect 3816 66 3846 4502
rect 3888 108 3918 4544
rect 3960 66 3990 4502
rect 4032 108 4062 4544
rect 4104 66 4134 4502
rect 4176 108 4206 4544
rect 4248 66 4278 4502
rect 4320 108 4350 4544
rect 4392 66 4422 4502
rect 4464 108 4494 4544
rect 4536 66 4566 4502
rect 4608 108 4638 4544
rect 4680 66 4710 4502
rect 4752 108 4782 4544
rect 4824 66 4854 4502
rect 4896 108 4926 4544
rect 4968 66 4998 4502
rect 5040 108 5070 4544
rect 5112 66 5142 4502
rect 5184 108 5214 4544
rect 5256 66 5286 4502
rect 5328 108 5358 4544
rect 5400 66 5430 4502
rect 5472 108 5502 4544
rect 5544 66 5574 4502
rect 5616 108 5646 4544
rect 5688 66 5718 4502
rect 5760 108 5790 4544
rect 5832 66 5862 4502
rect 5904 108 5934 4544
rect 5976 66 6006 4502
rect 6048 108 6078 4544
rect 6120 66 6150 4502
rect 6192 108 6222 4544
rect 6264 66 6294 4502
rect 6336 108 6366 4544
rect 6408 66 6438 4502
rect 6480 108 6510 4544
rect 6552 66 6582 4502
rect 6624 108 6654 4544
rect 6696 66 6726 4502
rect 6768 108 6798 4544
rect 6840 66 6870 4502
rect 6912 108 6942 4544
rect 6984 66 7014 4502
rect 7056 108 7086 4544
rect 7128 66 7158 4502
rect 7200 108 7230 4544
rect 7272 66 7302 4502
rect 7344 108 7374 4544
rect 7416 66 7446 4502
rect 7488 108 7518 4544
rect 7560 66 7590 4502
rect 7632 108 7662 4544
rect 7704 66 7734 4502
rect 7776 108 7806 4544
rect 7848 66 7878 4502
rect 7920 108 7950 4544
rect 7992 66 8022 4502
rect 8064 108 8094 4544
rect 8136 66 8166 4502
rect 8208 108 8238 4544
rect 8280 66 8310 4502
rect 8352 108 8382 4544
rect 8424 66 8454 4502
rect 8496 108 8526 4544
rect 8568 66 8598 4502
rect 8640 108 8670 4544
rect 8712 66 8742 4502
rect 8784 108 8814 4544
rect 8856 66 8886 4502
rect 8928 108 8958 4544
rect 9000 66 9030 4502
rect 9072 108 9102 4544
rect 9144 66 9174 4502
rect 9216 108 9246 4544
rect 9288 66 9318 4502
rect 9360 108 9390 4544
rect 9432 66 9462 4502
rect 9504 108 9534 4544
rect 9576 66 9606 4502
rect 9648 108 9678 4544
rect 9720 66 9750 4502
rect 9792 108 9822 4544
rect 9864 66 9894 4502
rect 9936 108 9966 4544
rect 10008 66 10038 4502
rect 10080 108 10110 4544
rect 10152 66 10182 4502
rect 10224 108 10254 4544
rect 10296 66 10326 4502
rect 10368 108 10398 4544
rect 10440 66 10470 4502
rect 10512 108 10542 4544
rect 10584 66 10614 4502
rect 10656 108 10686 4544
rect 10728 66 10758 4502
rect 10800 108 10830 4544
rect 10872 66 10902 4502
rect 10944 108 10974 4544
rect 11016 66 11046 4502
rect 11088 108 11146 4544
rect 0 50 11146 66
rect 0 16 34 50
rect 68 16 102 50
rect 136 16 170 50
rect 204 16 238 50
rect 272 16 306 50
rect 340 16 374 50
rect 408 16 442 50
rect 476 16 510 50
rect 544 16 578 50
rect 612 16 646 50
rect 680 16 714 50
rect 748 16 782 50
rect 816 16 850 50
rect 884 16 918 50
rect 952 16 986 50
rect 1020 16 1054 50
rect 1088 16 1122 50
rect 1156 16 1190 50
rect 1224 16 1258 50
rect 1292 16 1326 50
rect 1360 16 1394 50
rect 1428 16 1462 50
rect 1496 16 1530 50
rect 1564 16 1598 50
rect 1632 16 1666 50
rect 1700 16 1734 50
rect 1768 16 1802 50
rect 1836 16 1870 50
rect 1904 16 1938 50
rect 1972 16 2006 50
rect 2040 16 2074 50
rect 2108 16 2142 50
rect 2176 16 2210 50
rect 2244 16 2278 50
rect 2312 16 2346 50
rect 2380 16 2414 50
rect 2448 16 2482 50
rect 2516 16 2550 50
rect 2584 16 2618 50
rect 2652 16 2686 50
rect 2720 16 2754 50
rect 2788 16 2822 50
rect 2856 16 2890 50
rect 2924 16 2958 50
rect 2992 16 3026 50
rect 3060 16 3094 50
rect 3128 16 3162 50
rect 3196 16 3230 50
rect 3264 16 3298 50
rect 3332 16 3366 50
rect 3400 16 3434 50
rect 3468 16 3502 50
rect 3536 16 3570 50
rect 3604 16 3638 50
rect 3672 16 3706 50
rect 3740 16 3774 50
rect 3808 16 3842 50
rect 3876 16 3910 50
rect 3944 16 3978 50
rect 4012 16 4046 50
rect 4080 16 4114 50
rect 4148 16 4182 50
rect 4216 16 4250 50
rect 4284 16 4318 50
rect 4352 16 4386 50
rect 4420 16 4454 50
rect 4488 16 4522 50
rect 4556 16 4590 50
rect 4624 16 4658 50
rect 4692 16 4726 50
rect 4760 16 4794 50
rect 4828 16 4862 50
rect 4896 16 4930 50
rect 4964 16 4998 50
rect 5032 16 5066 50
rect 5100 16 5134 50
rect 5168 16 5202 50
rect 5236 16 5270 50
rect 5304 16 5338 50
rect 5372 16 5406 50
rect 5440 16 5474 50
rect 5508 16 5542 50
rect 5576 16 5610 50
rect 5644 16 5678 50
rect 5712 16 5746 50
rect 5780 16 5814 50
rect 5848 16 5882 50
rect 5916 16 5950 50
rect 5984 16 6018 50
rect 6052 16 6086 50
rect 6120 16 6154 50
rect 6188 16 6222 50
rect 6256 16 6290 50
rect 6324 16 6358 50
rect 6392 16 6426 50
rect 6460 16 6494 50
rect 6528 16 6562 50
rect 6596 16 6630 50
rect 6664 16 6698 50
rect 6732 16 6766 50
rect 6800 16 6834 50
rect 6868 16 6902 50
rect 6936 16 6970 50
rect 7004 16 7038 50
rect 7072 16 7106 50
rect 7140 16 7174 50
rect 7208 16 7242 50
rect 7276 16 7310 50
rect 7344 16 7378 50
rect 7412 16 7446 50
rect 7480 16 7514 50
rect 7548 16 7582 50
rect 7616 16 7650 50
rect 7684 16 7718 50
rect 7752 16 7786 50
rect 7820 16 7854 50
rect 7888 16 7922 50
rect 7956 16 7990 50
rect 8024 16 8058 50
rect 8092 16 8126 50
rect 8160 16 8194 50
rect 8228 16 8262 50
rect 8296 16 8330 50
rect 8364 16 8398 50
rect 8432 16 8466 50
rect 8500 16 8534 50
rect 8568 16 8602 50
rect 8636 16 8670 50
rect 8704 16 8738 50
rect 8772 16 8806 50
rect 8840 16 8874 50
rect 8908 16 8942 50
rect 8976 16 9010 50
rect 9044 16 9078 50
rect 9112 16 9146 50
rect 9180 16 9214 50
rect 9248 16 9282 50
rect 9316 16 9350 50
rect 9384 16 9418 50
rect 9452 16 9486 50
rect 9520 16 9554 50
rect 9588 16 9622 50
rect 9656 16 9690 50
rect 9724 16 9758 50
rect 9792 16 9826 50
rect 9860 16 9894 50
rect 9928 16 9962 50
rect 9996 16 10030 50
rect 10064 16 10098 50
rect 10132 16 10166 50
rect 10200 16 10234 50
rect 10268 16 10302 50
rect 10336 16 10370 50
rect 10404 16 10438 50
rect 10472 16 10506 50
rect 10540 16 10574 50
rect 10608 16 10642 50
rect 10676 16 10710 50
rect 10744 16 10778 50
rect 10812 16 10846 50
rect 10880 16 10914 50
rect 10948 16 10982 50
rect 11016 16 11050 50
rect 11084 16 11146 50
rect 0 0 11146 16
<< polycont >>
rect 34 4560 68 4594
rect 102 4560 136 4594
rect 170 4560 204 4594
rect 238 4560 272 4594
rect 306 4560 340 4594
rect 374 4560 408 4594
rect 442 4560 476 4594
rect 510 4560 544 4594
rect 578 4560 612 4594
rect 646 4560 680 4594
rect 714 4560 748 4594
rect 782 4560 816 4594
rect 850 4560 884 4594
rect 918 4560 952 4594
rect 986 4560 1020 4594
rect 1054 4560 1088 4594
rect 1122 4560 1156 4594
rect 1190 4560 1224 4594
rect 1258 4560 1292 4594
rect 1326 4560 1360 4594
rect 1394 4560 1428 4594
rect 1462 4560 1496 4594
rect 1530 4560 1564 4594
rect 1598 4560 1632 4594
rect 1666 4560 1700 4594
rect 1734 4560 1768 4594
rect 1802 4560 1836 4594
rect 1870 4560 1904 4594
rect 1938 4560 1972 4594
rect 2006 4560 2040 4594
rect 2074 4560 2108 4594
rect 2142 4560 2176 4594
rect 2210 4560 2244 4594
rect 2278 4560 2312 4594
rect 2346 4560 2380 4594
rect 2414 4560 2448 4594
rect 2482 4560 2516 4594
rect 2550 4560 2584 4594
rect 2618 4560 2652 4594
rect 2686 4560 2720 4594
rect 2754 4560 2788 4594
rect 2822 4560 2856 4594
rect 2890 4560 2924 4594
rect 2958 4560 2992 4594
rect 3026 4560 3060 4594
rect 3094 4560 3128 4594
rect 3162 4560 3196 4594
rect 3230 4560 3264 4594
rect 3298 4560 3332 4594
rect 3366 4560 3400 4594
rect 3434 4560 3468 4594
rect 3502 4560 3536 4594
rect 3570 4560 3604 4594
rect 3638 4560 3672 4594
rect 3706 4560 3740 4594
rect 3774 4560 3808 4594
rect 3842 4560 3876 4594
rect 3910 4560 3944 4594
rect 3978 4560 4012 4594
rect 4046 4560 4080 4594
rect 4114 4560 4148 4594
rect 4182 4560 4216 4594
rect 4250 4560 4284 4594
rect 4318 4560 4352 4594
rect 4386 4560 4420 4594
rect 4454 4560 4488 4594
rect 4522 4560 4556 4594
rect 4590 4560 4624 4594
rect 4658 4560 4692 4594
rect 4726 4560 4760 4594
rect 4794 4560 4828 4594
rect 4862 4560 4896 4594
rect 4930 4560 4964 4594
rect 4998 4560 5032 4594
rect 5066 4560 5100 4594
rect 5134 4560 5168 4594
rect 5202 4560 5236 4594
rect 5270 4560 5304 4594
rect 5338 4560 5372 4594
rect 5406 4560 5440 4594
rect 5474 4560 5508 4594
rect 5542 4560 5576 4594
rect 5610 4560 5644 4594
rect 5678 4560 5712 4594
rect 5746 4560 5780 4594
rect 5814 4560 5848 4594
rect 5882 4560 5916 4594
rect 5950 4560 5984 4594
rect 6018 4560 6052 4594
rect 6086 4560 6120 4594
rect 6154 4560 6188 4594
rect 6222 4560 6256 4594
rect 6290 4560 6324 4594
rect 6358 4560 6392 4594
rect 6426 4560 6460 4594
rect 6494 4560 6528 4594
rect 6562 4560 6596 4594
rect 6630 4560 6664 4594
rect 6698 4560 6732 4594
rect 6766 4560 6800 4594
rect 6834 4560 6868 4594
rect 6902 4560 6936 4594
rect 6970 4560 7004 4594
rect 7038 4560 7072 4594
rect 7106 4560 7140 4594
rect 7174 4560 7208 4594
rect 7242 4560 7276 4594
rect 7310 4560 7344 4594
rect 7378 4560 7412 4594
rect 7446 4560 7480 4594
rect 7514 4560 7548 4594
rect 7582 4560 7616 4594
rect 7650 4560 7684 4594
rect 7718 4560 7752 4594
rect 7786 4560 7820 4594
rect 7854 4560 7888 4594
rect 7922 4560 7956 4594
rect 7990 4560 8024 4594
rect 8058 4560 8092 4594
rect 8126 4560 8160 4594
rect 8194 4560 8228 4594
rect 8262 4560 8296 4594
rect 8330 4560 8364 4594
rect 8398 4560 8432 4594
rect 8466 4560 8500 4594
rect 8534 4560 8568 4594
rect 8602 4560 8636 4594
rect 8670 4560 8704 4594
rect 8738 4560 8772 4594
rect 8806 4560 8840 4594
rect 8874 4560 8908 4594
rect 8942 4560 8976 4594
rect 9010 4560 9044 4594
rect 9078 4560 9112 4594
rect 9146 4560 9180 4594
rect 9214 4560 9248 4594
rect 9282 4560 9316 4594
rect 9350 4560 9384 4594
rect 9418 4560 9452 4594
rect 9486 4560 9520 4594
rect 9554 4560 9588 4594
rect 9622 4560 9656 4594
rect 9690 4560 9724 4594
rect 9758 4560 9792 4594
rect 9826 4560 9860 4594
rect 9894 4560 9928 4594
rect 9962 4560 9996 4594
rect 10030 4560 10064 4594
rect 10098 4560 10132 4594
rect 10166 4560 10200 4594
rect 10234 4560 10268 4594
rect 10302 4560 10336 4594
rect 10370 4560 10404 4594
rect 10438 4560 10472 4594
rect 10506 4560 10540 4594
rect 10574 4560 10608 4594
rect 10642 4560 10676 4594
rect 10710 4560 10744 4594
rect 10778 4560 10812 4594
rect 10846 4560 10880 4594
rect 10914 4560 10948 4594
rect 10982 4560 11016 4594
rect 11050 4560 11084 4594
rect 34 16 68 50
rect 102 16 136 50
rect 170 16 204 50
rect 238 16 272 50
rect 306 16 340 50
rect 374 16 408 50
rect 442 16 476 50
rect 510 16 544 50
rect 578 16 612 50
rect 646 16 680 50
rect 714 16 748 50
rect 782 16 816 50
rect 850 16 884 50
rect 918 16 952 50
rect 986 16 1020 50
rect 1054 16 1088 50
rect 1122 16 1156 50
rect 1190 16 1224 50
rect 1258 16 1292 50
rect 1326 16 1360 50
rect 1394 16 1428 50
rect 1462 16 1496 50
rect 1530 16 1564 50
rect 1598 16 1632 50
rect 1666 16 1700 50
rect 1734 16 1768 50
rect 1802 16 1836 50
rect 1870 16 1904 50
rect 1938 16 1972 50
rect 2006 16 2040 50
rect 2074 16 2108 50
rect 2142 16 2176 50
rect 2210 16 2244 50
rect 2278 16 2312 50
rect 2346 16 2380 50
rect 2414 16 2448 50
rect 2482 16 2516 50
rect 2550 16 2584 50
rect 2618 16 2652 50
rect 2686 16 2720 50
rect 2754 16 2788 50
rect 2822 16 2856 50
rect 2890 16 2924 50
rect 2958 16 2992 50
rect 3026 16 3060 50
rect 3094 16 3128 50
rect 3162 16 3196 50
rect 3230 16 3264 50
rect 3298 16 3332 50
rect 3366 16 3400 50
rect 3434 16 3468 50
rect 3502 16 3536 50
rect 3570 16 3604 50
rect 3638 16 3672 50
rect 3706 16 3740 50
rect 3774 16 3808 50
rect 3842 16 3876 50
rect 3910 16 3944 50
rect 3978 16 4012 50
rect 4046 16 4080 50
rect 4114 16 4148 50
rect 4182 16 4216 50
rect 4250 16 4284 50
rect 4318 16 4352 50
rect 4386 16 4420 50
rect 4454 16 4488 50
rect 4522 16 4556 50
rect 4590 16 4624 50
rect 4658 16 4692 50
rect 4726 16 4760 50
rect 4794 16 4828 50
rect 4862 16 4896 50
rect 4930 16 4964 50
rect 4998 16 5032 50
rect 5066 16 5100 50
rect 5134 16 5168 50
rect 5202 16 5236 50
rect 5270 16 5304 50
rect 5338 16 5372 50
rect 5406 16 5440 50
rect 5474 16 5508 50
rect 5542 16 5576 50
rect 5610 16 5644 50
rect 5678 16 5712 50
rect 5746 16 5780 50
rect 5814 16 5848 50
rect 5882 16 5916 50
rect 5950 16 5984 50
rect 6018 16 6052 50
rect 6086 16 6120 50
rect 6154 16 6188 50
rect 6222 16 6256 50
rect 6290 16 6324 50
rect 6358 16 6392 50
rect 6426 16 6460 50
rect 6494 16 6528 50
rect 6562 16 6596 50
rect 6630 16 6664 50
rect 6698 16 6732 50
rect 6766 16 6800 50
rect 6834 16 6868 50
rect 6902 16 6936 50
rect 6970 16 7004 50
rect 7038 16 7072 50
rect 7106 16 7140 50
rect 7174 16 7208 50
rect 7242 16 7276 50
rect 7310 16 7344 50
rect 7378 16 7412 50
rect 7446 16 7480 50
rect 7514 16 7548 50
rect 7582 16 7616 50
rect 7650 16 7684 50
rect 7718 16 7752 50
rect 7786 16 7820 50
rect 7854 16 7888 50
rect 7922 16 7956 50
rect 7990 16 8024 50
rect 8058 16 8092 50
rect 8126 16 8160 50
rect 8194 16 8228 50
rect 8262 16 8296 50
rect 8330 16 8364 50
rect 8398 16 8432 50
rect 8466 16 8500 50
rect 8534 16 8568 50
rect 8602 16 8636 50
rect 8670 16 8704 50
rect 8738 16 8772 50
rect 8806 16 8840 50
rect 8874 16 8908 50
rect 8942 16 8976 50
rect 9010 16 9044 50
rect 9078 16 9112 50
rect 9146 16 9180 50
rect 9214 16 9248 50
rect 9282 16 9316 50
rect 9350 16 9384 50
rect 9418 16 9452 50
rect 9486 16 9520 50
rect 9554 16 9588 50
rect 9622 16 9656 50
rect 9690 16 9724 50
rect 9758 16 9792 50
rect 9826 16 9860 50
rect 9894 16 9928 50
rect 9962 16 9996 50
rect 10030 16 10064 50
rect 10098 16 10132 50
rect 10166 16 10200 50
rect 10234 16 10268 50
rect 10302 16 10336 50
rect 10370 16 10404 50
rect 10438 16 10472 50
rect 10506 16 10540 50
rect 10574 16 10608 50
rect 10642 16 10676 50
rect 10710 16 10744 50
rect 10778 16 10812 50
rect 10846 16 10880 50
rect 10914 16 10948 50
rect 10982 16 11016 50
rect 11050 16 11084 50
<< locali >>
rect 0 4594 11146 4610
rect 0 4560 34 4594
rect 72 4560 102 4594
rect 144 4560 170 4594
rect 216 4560 238 4594
rect 288 4560 306 4594
rect 360 4560 374 4594
rect 432 4560 442 4594
rect 504 4560 510 4594
rect 576 4560 578 4594
rect 612 4560 614 4594
rect 680 4560 686 4594
rect 748 4560 758 4594
rect 816 4560 830 4594
rect 884 4560 902 4594
rect 952 4560 974 4594
rect 1020 4560 1046 4594
rect 1088 4560 1118 4594
rect 1156 4560 1190 4594
rect 1224 4560 1258 4594
rect 1296 4560 1326 4594
rect 1368 4560 1394 4594
rect 1440 4560 1462 4594
rect 1512 4560 1530 4594
rect 1584 4560 1598 4594
rect 1656 4560 1666 4594
rect 1728 4560 1734 4594
rect 1800 4560 1802 4594
rect 1836 4560 1838 4594
rect 1904 4560 1910 4594
rect 1972 4560 1982 4594
rect 2040 4560 2054 4594
rect 2108 4560 2126 4594
rect 2176 4560 2198 4594
rect 2244 4560 2270 4594
rect 2312 4560 2342 4594
rect 2380 4560 2414 4594
rect 2448 4560 2482 4594
rect 2520 4560 2550 4594
rect 2592 4560 2618 4594
rect 2664 4560 2686 4594
rect 2736 4560 2754 4594
rect 2808 4560 2822 4594
rect 2880 4560 2890 4594
rect 2952 4560 2958 4594
rect 3024 4560 3026 4594
rect 3060 4560 3062 4594
rect 3128 4560 3134 4594
rect 3196 4560 3206 4594
rect 3264 4560 3278 4594
rect 3332 4560 3350 4594
rect 3400 4560 3422 4594
rect 3468 4560 3494 4594
rect 3536 4560 3566 4594
rect 3604 4560 3638 4594
rect 3672 4560 3706 4594
rect 3744 4560 3774 4594
rect 3816 4560 3842 4594
rect 3888 4560 3910 4594
rect 3960 4560 3978 4594
rect 4032 4560 4046 4594
rect 4104 4560 4114 4594
rect 4176 4560 4182 4594
rect 4248 4560 4250 4594
rect 4284 4560 4286 4594
rect 4352 4560 4358 4594
rect 4420 4560 4430 4594
rect 4488 4560 4502 4594
rect 4556 4560 4574 4594
rect 4624 4560 4646 4594
rect 4692 4560 4718 4594
rect 4760 4560 4790 4594
rect 4828 4560 4862 4594
rect 4896 4560 4930 4594
rect 4968 4560 4998 4594
rect 5040 4560 5066 4594
rect 5112 4560 5134 4594
rect 5184 4560 5202 4594
rect 5256 4560 5270 4594
rect 5328 4560 5338 4594
rect 5400 4560 5406 4594
rect 5472 4560 5474 4594
rect 5508 4560 5510 4594
rect 5576 4560 5582 4594
rect 5644 4560 5654 4594
rect 5712 4560 5726 4594
rect 5780 4560 5798 4594
rect 5848 4560 5870 4594
rect 5916 4560 5942 4594
rect 5984 4560 6014 4594
rect 6052 4560 6086 4594
rect 6120 4560 6154 4594
rect 6192 4560 6222 4594
rect 6264 4560 6290 4594
rect 6336 4560 6358 4594
rect 6408 4560 6426 4594
rect 6480 4560 6494 4594
rect 6552 4560 6562 4594
rect 6624 4560 6630 4594
rect 6696 4560 6698 4594
rect 6732 4560 6734 4594
rect 6800 4560 6806 4594
rect 6868 4560 6878 4594
rect 6936 4560 6950 4594
rect 7004 4560 7022 4594
rect 7072 4560 7094 4594
rect 7140 4560 7166 4594
rect 7208 4560 7238 4594
rect 7276 4560 7310 4594
rect 7344 4560 7378 4594
rect 7416 4560 7446 4594
rect 7488 4560 7514 4594
rect 7560 4560 7582 4594
rect 7632 4560 7650 4594
rect 7704 4560 7718 4594
rect 7776 4560 7786 4594
rect 7848 4560 7854 4594
rect 7920 4560 7922 4594
rect 7956 4560 7958 4594
rect 8024 4560 8030 4594
rect 8092 4560 8102 4594
rect 8160 4560 8174 4594
rect 8228 4560 8246 4594
rect 8296 4560 8318 4594
rect 8364 4560 8390 4594
rect 8432 4560 8462 4594
rect 8500 4560 8534 4594
rect 8568 4560 8602 4594
rect 8640 4560 8670 4594
rect 8712 4560 8738 4594
rect 8784 4560 8806 4594
rect 8856 4560 8874 4594
rect 8928 4560 8942 4594
rect 9000 4560 9010 4594
rect 9072 4560 9078 4594
rect 9144 4560 9146 4594
rect 9180 4560 9182 4594
rect 9248 4560 9254 4594
rect 9316 4560 9326 4594
rect 9384 4560 9398 4594
rect 9452 4560 9470 4594
rect 9520 4560 9542 4594
rect 9588 4560 9614 4594
rect 9656 4560 9686 4594
rect 9724 4560 9758 4594
rect 9792 4560 9826 4594
rect 9864 4560 9894 4594
rect 9936 4560 9962 4594
rect 10008 4560 10030 4594
rect 10080 4560 10098 4594
rect 10152 4560 10166 4594
rect 10224 4560 10234 4594
rect 10296 4560 10302 4594
rect 10368 4560 10370 4594
rect 10404 4560 10406 4594
rect 10472 4560 10478 4594
rect 10540 4560 10550 4594
rect 10608 4560 10622 4594
rect 10676 4560 10694 4594
rect 10744 4560 10766 4594
rect 10812 4560 10838 4594
rect 10880 4560 10910 4594
rect 10948 4560 10982 4594
rect 11016 4560 11050 4594
rect 11088 4560 11146 4594
rect 0 4544 11146 4560
rect 0 66 28 4516
rect 56 94 84 4544
rect 112 66 140 4516
rect 168 94 196 4544
rect 224 66 252 4516
rect 280 94 308 4544
rect 336 66 364 4516
rect 392 94 420 4544
rect 448 66 476 4516
rect 504 94 532 4544
rect 560 66 588 4516
rect 616 94 644 4544
rect 672 66 700 4516
rect 728 94 756 4544
rect 784 66 812 4516
rect 840 94 868 4544
rect 896 66 924 4516
rect 952 94 980 4544
rect 1008 66 1036 4516
rect 1064 94 1092 4544
rect 1120 66 1148 4516
rect 1176 94 1204 4544
rect 1232 66 1260 4516
rect 1288 94 1316 4544
rect 1344 66 1372 4516
rect 1400 94 1428 4544
rect 1456 66 1484 4516
rect 1512 94 1540 4544
rect 1568 66 1596 4516
rect 1624 94 1652 4544
rect 1680 66 1708 4516
rect 1736 94 1764 4544
rect 1792 66 1820 4516
rect 1848 94 1876 4544
rect 1904 66 1932 4516
rect 1960 94 1988 4544
rect 2016 66 2044 4516
rect 2072 94 2100 4544
rect 2128 66 2156 4516
rect 2184 94 2212 4544
rect 2240 66 2268 4516
rect 2296 94 2324 4544
rect 2352 66 2380 4516
rect 2408 94 2436 4544
rect 2464 66 2492 4516
rect 2520 94 2548 4544
rect 2576 66 2604 4516
rect 2632 94 2660 4544
rect 2688 66 2716 4516
rect 2744 94 2772 4544
rect 2800 66 2828 4516
rect 2856 94 2884 4544
rect 2912 66 2940 4516
rect 2968 94 2996 4544
rect 3024 66 3052 4516
rect 3080 94 3108 4544
rect 3136 66 3164 4516
rect 3192 94 3220 4544
rect 3248 66 3276 4516
rect 3304 94 3332 4544
rect 3360 66 3388 4516
rect 3416 94 3444 4544
rect 3472 66 3500 4516
rect 3528 94 3556 4544
rect 3584 66 3612 4516
rect 3640 94 3668 4544
rect 3696 66 3724 4516
rect 3752 94 3780 4544
rect 3808 66 3836 4516
rect 3864 94 3892 4544
rect 3920 66 3948 4516
rect 3976 94 4004 4544
rect 4032 66 4060 4516
rect 4088 94 4116 4544
rect 4144 66 4172 4516
rect 4200 94 4228 4544
rect 4256 66 4284 4516
rect 4312 94 4340 4544
rect 4368 66 4396 4516
rect 4424 94 4452 4544
rect 4480 66 4508 4516
rect 4536 94 4564 4544
rect 4592 66 4620 4516
rect 4648 94 4676 4544
rect 4704 66 4732 4516
rect 4760 94 4788 4544
rect 4816 66 4844 4516
rect 4872 94 4900 4544
rect 4928 66 4956 4516
rect 4984 94 5012 4544
rect 5040 66 5068 4516
rect 5096 94 5124 4544
rect 5152 66 5180 4516
rect 5208 94 5236 4544
rect 5264 66 5292 4516
rect 5320 94 5348 4544
rect 5376 66 5404 4516
rect 5432 94 5460 4544
rect 5488 66 5516 4516
rect 5544 94 5572 4544
rect 5600 66 5628 4516
rect 5656 94 5684 4544
rect 5712 66 5740 4516
rect 5768 94 5796 4544
rect 5824 66 5852 4516
rect 5880 94 5908 4544
rect 5936 66 5964 4516
rect 5992 94 6020 4544
rect 6048 66 6076 4516
rect 6104 94 6132 4544
rect 6160 66 6188 4516
rect 6216 94 6244 4544
rect 6272 66 6300 4516
rect 6328 94 6356 4544
rect 6384 66 6412 4516
rect 6440 94 6468 4544
rect 6496 66 6524 4516
rect 6552 94 6580 4544
rect 6608 66 6636 4516
rect 6664 94 6692 4544
rect 6720 66 6748 4516
rect 6776 94 6804 4544
rect 6832 66 6860 4516
rect 6888 94 6916 4544
rect 6944 66 6972 4516
rect 7000 94 7028 4544
rect 7056 66 7084 4516
rect 7112 94 7140 4544
rect 7168 66 7196 4516
rect 7224 94 7252 4544
rect 7280 66 7308 4516
rect 7336 94 7364 4544
rect 7392 66 7420 4516
rect 7448 94 7476 4544
rect 7504 66 7532 4516
rect 7560 94 7588 4544
rect 7616 66 7644 4516
rect 7672 94 7700 4544
rect 7728 66 7756 4516
rect 7784 94 7812 4544
rect 7840 66 7868 4516
rect 7896 94 7924 4544
rect 7952 66 7980 4516
rect 8008 94 8036 4544
rect 8064 66 8092 4516
rect 8120 94 8148 4544
rect 8176 66 8204 4516
rect 8232 94 8260 4544
rect 8288 66 8316 4516
rect 8344 94 8372 4544
rect 8400 66 8428 4516
rect 8456 94 8484 4544
rect 8512 66 8540 4516
rect 8568 94 8596 4544
rect 8624 66 8652 4516
rect 8680 94 8708 4544
rect 8736 66 8764 4516
rect 8792 94 8820 4544
rect 8848 66 8876 4516
rect 8904 94 8932 4544
rect 8960 66 8988 4516
rect 9016 94 9044 4544
rect 9072 66 9100 4516
rect 9128 94 9156 4544
rect 9184 66 9212 4516
rect 9240 94 9268 4544
rect 9296 66 9324 4516
rect 9352 94 9380 4544
rect 9408 66 9436 4516
rect 9464 94 9492 4544
rect 9520 66 9548 4516
rect 9576 94 9604 4544
rect 9632 66 9660 4516
rect 9688 94 9716 4544
rect 9744 66 9772 4516
rect 9800 94 9828 4544
rect 9856 66 9884 4516
rect 9912 94 9940 4544
rect 9968 66 9996 4516
rect 10024 94 10052 4544
rect 10080 66 10108 4516
rect 10136 94 10164 4544
rect 10192 66 10220 4516
rect 10248 94 10276 4544
rect 10304 66 10332 4516
rect 10360 94 10388 4544
rect 10416 66 10444 4516
rect 10472 94 10500 4544
rect 10528 66 10556 4516
rect 10584 94 10612 4544
rect 10640 66 10668 4516
rect 10696 94 10724 4544
rect 10752 66 10780 4516
rect 10808 94 10836 4544
rect 10864 66 10892 4516
rect 10920 94 10948 4544
rect 10976 66 11004 4516
rect 11032 94 11060 4544
rect 11088 66 11146 4516
rect 0 50 11146 66
rect 0 16 34 50
rect 72 16 102 50
rect 144 16 170 50
rect 216 16 238 50
rect 288 16 306 50
rect 360 16 374 50
rect 432 16 442 50
rect 504 16 510 50
rect 576 16 578 50
rect 612 16 614 50
rect 680 16 686 50
rect 748 16 758 50
rect 816 16 830 50
rect 884 16 902 50
rect 952 16 974 50
rect 1020 16 1046 50
rect 1088 16 1118 50
rect 1156 16 1190 50
rect 1224 16 1258 50
rect 1296 16 1326 50
rect 1368 16 1394 50
rect 1440 16 1462 50
rect 1512 16 1530 50
rect 1584 16 1598 50
rect 1656 16 1666 50
rect 1728 16 1734 50
rect 1800 16 1802 50
rect 1836 16 1838 50
rect 1904 16 1910 50
rect 1972 16 1982 50
rect 2040 16 2054 50
rect 2108 16 2126 50
rect 2176 16 2198 50
rect 2244 16 2270 50
rect 2312 16 2342 50
rect 2380 16 2414 50
rect 2448 16 2482 50
rect 2520 16 2550 50
rect 2592 16 2618 50
rect 2664 16 2686 50
rect 2736 16 2754 50
rect 2808 16 2822 50
rect 2880 16 2890 50
rect 2952 16 2958 50
rect 3024 16 3026 50
rect 3060 16 3062 50
rect 3128 16 3134 50
rect 3196 16 3206 50
rect 3264 16 3278 50
rect 3332 16 3350 50
rect 3400 16 3422 50
rect 3468 16 3494 50
rect 3536 16 3566 50
rect 3604 16 3638 50
rect 3672 16 3706 50
rect 3744 16 3774 50
rect 3816 16 3842 50
rect 3888 16 3910 50
rect 3960 16 3978 50
rect 4032 16 4046 50
rect 4104 16 4114 50
rect 4176 16 4182 50
rect 4248 16 4250 50
rect 4284 16 4286 50
rect 4352 16 4358 50
rect 4420 16 4430 50
rect 4488 16 4502 50
rect 4556 16 4574 50
rect 4624 16 4646 50
rect 4692 16 4718 50
rect 4760 16 4790 50
rect 4828 16 4862 50
rect 4896 16 4930 50
rect 4968 16 4998 50
rect 5040 16 5066 50
rect 5112 16 5134 50
rect 5184 16 5202 50
rect 5256 16 5270 50
rect 5328 16 5338 50
rect 5400 16 5406 50
rect 5472 16 5474 50
rect 5508 16 5510 50
rect 5576 16 5582 50
rect 5644 16 5654 50
rect 5712 16 5726 50
rect 5780 16 5798 50
rect 5848 16 5870 50
rect 5916 16 5942 50
rect 5984 16 6014 50
rect 6052 16 6086 50
rect 6120 16 6154 50
rect 6192 16 6222 50
rect 6264 16 6290 50
rect 6336 16 6358 50
rect 6408 16 6426 50
rect 6480 16 6494 50
rect 6552 16 6562 50
rect 6624 16 6630 50
rect 6696 16 6698 50
rect 6732 16 6734 50
rect 6800 16 6806 50
rect 6868 16 6878 50
rect 6936 16 6950 50
rect 7004 16 7022 50
rect 7072 16 7094 50
rect 7140 16 7166 50
rect 7208 16 7238 50
rect 7276 16 7310 50
rect 7344 16 7378 50
rect 7416 16 7446 50
rect 7488 16 7514 50
rect 7560 16 7582 50
rect 7632 16 7650 50
rect 7704 16 7718 50
rect 7776 16 7786 50
rect 7848 16 7854 50
rect 7920 16 7922 50
rect 7956 16 7958 50
rect 8024 16 8030 50
rect 8092 16 8102 50
rect 8160 16 8174 50
rect 8228 16 8246 50
rect 8296 16 8318 50
rect 8364 16 8390 50
rect 8432 16 8462 50
rect 8500 16 8534 50
rect 8568 16 8602 50
rect 8640 16 8670 50
rect 8712 16 8738 50
rect 8784 16 8806 50
rect 8856 16 8874 50
rect 8928 16 8942 50
rect 9000 16 9010 50
rect 9072 16 9078 50
rect 9144 16 9146 50
rect 9180 16 9182 50
rect 9248 16 9254 50
rect 9316 16 9326 50
rect 9384 16 9398 50
rect 9452 16 9470 50
rect 9520 16 9542 50
rect 9588 16 9614 50
rect 9656 16 9686 50
rect 9724 16 9758 50
rect 9792 16 9826 50
rect 9864 16 9894 50
rect 9936 16 9962 50
rect 10008 16 10030 50
rect 10080 16 10098 50
rect 10152 16 10166 50
rect 10224 16 10234 50
rect 10296 16 10302 50
rect 10368 16 10370 50
rect 10404 16 10406 50
rect 10472 16 10478 50
rect 10540 16 10550 50
rect 10608 16 10622 50
rect 10676 16 10694 50
rect 10744 16 10766 50
rect 10812 16 10838 50
rect 10880 16 10910 50
rect 10948 16 10982 50
rect 11016 16 11050 50
rect 11088 16 11146 50
rect 0 0 11146 16
<< viali >>
rect 38 4560 68 4594
rect 68 4560 72 4594
rect 110 4560 136 4594
rect 136 4560 144 4594
rect 182 4560 204 4594
rect 204 4560 216 4594
rect 254 4560 272 4594
rect 272 4560 288 4594
rect 326 4560 340 4594
rect 340 4560 360 4594
rect 398 4560 408 4594
rect 408 4560 432 4594
rect 470 4560 476 4594
rect 476 4560 504 4594
rect 542 4560 544 4594
rect 544 4560 576 4594
rect 614 4560 646 4594
rect 646 4560 648 4594
rect 686 4560 714 4594
rect 714 4560 720 4594
rect 758 4560 782 4594
rect 782 4560 792 4594
rect 830 4560 850 4594
rect 850 4560 864 4594
rect 902 4560 918 4594
rect 918 4560 936 4594
rect 974 4560 986 4594
rect 986 4560 1008 4594
rect 1046 4560 1054 4594
rect 1054 4560 1080 4594
rect 1118 4560 1122 4594
rect 1122 4560 1152 4594
rect 1190 4560 1224 4594
rect 1262 4560 1292 4594
rect 1292 4560 1296 4594
rect 1334 4560 1360 4594
rect 1360 4560 1368 4594
rect 1406 4560 1428 4594
rect 1428 4560 1440 4594
rect 1478 4560 1496 4594
rect 1496 4560 1512 4594
rect 1550 4560 1564 4594
rect 1564 4560 1584 4594
rect 1622 4560 1632 4594
rect 1632 4560 1656 4594
rect 1694 4560 1700 4594
rect 1700 4560 1728 4594
rect 1766 4560 1768 4594
rect 1768 4560 1800 4594
rect 1838 4560 1870 4594
rect 1870 4560 1872 4594
rect 1910 4560 1938 4594
rect 1938 4560 1944 4594
rect 1982 4560 2006 4594
rect 2006 4560 2016 4594
rect 2054 4560 2074 4594
rect 2074 4560 2088 4594
rect 2126 4560 2142 4594
rect 2142 4560 2160 4594
rect 2198 4560 2210 4594
rect 2210 4560 2232 4594
rect 2270 4560 2278 4594
rect 2278 4560 2304 4594
rect 2342 4560 2346 4594
rect 2346 4560 2376 4594
rect 2414 4560 2448 4594
rect 2486 4560 2516 4594
rect 2516 4560 2520 4594
rect 2558 4560 2584 4594
rect 2584 4560 2592 4594
rect 2630 4560 2652 4594
rect 2652 4560 2664 4594
rect 2702 4560 2720 4594
rect 2720 4560 2736 4594
rect 2774 4560 2788 4594
rect 2788 4560 2808 4594
rect 2846 4560 2856 4594
rect 2856 4560 2880 4594
rect 2918 4560 2924 4594
rect 2924 4560 2952 4594
rect 2990 4560 2992 4594
rect 2992 4560 3024 4594
rect 3062 4560 3094 4594
rect 3094 4560 3096 4594
rect 3134 4560 3162 4594
rect 3162 4560 3168 4594
rect 3206 4560 3230 4594
rect 3230 4560 3240 4594
rect 3278 4560 3298 4594
rect 3298 4560 3312 4594
rect 3350 4560 3366 4594
rect 3366 4560 3384 4594
rect 3422 4560 3434 4594
rect 3434 4560 3456 4594
rect 3494 4560 3502 4594
rect 3502 4560 3528 4594
rect 3566 4560 3570 4594
rect 3570 4560 3600 4594
rect 3638 4560 3672 4594
rect 3710 4560 3740 4594
rect 3740 4560 3744 4594
rect 3782 4560 3808 4594
rect 3808 4560 3816 4594
rect 3854 4560 3876 4594
rect 3876 4560 3888 4594
rect 3926 4560 3944 4594
rect 3944 4560 3960 4594
rect 3998 4560 4012 4594
rect 4012 4560 4032 4594
rect 4070 4560 4080 4594
rect 4080 4560 4104 4594
rect 4142 4560 4148 4594
rect 4148 4560 4176 4594
rect 4214 4560 4216 4594
rect 4216 4560 4248 4594
rect 4286 4560 4318 4594
rect 4318 4560 4320 4594
rect 4358 4560 4386 4594
rect 4386 4560 4392 4594
rect 4430 4560 4454 4594
rect 4454 4560 4464 4594
rect 4502 4560 4522 4594
rect 4522 4560 4536 4594
rect 4574 4560 4590 4594
rect 4590 4560 4608 4594
rect 4646 4560 4658 4594
rect 4658 4560 4680 4594
rect 4718 4560 4726 4594
rect 4726 4560 4752 4594
rect 4790 4560 4794 4594
rect 4794 4560 4824 4594
rect 4862 4560 4896 4594
rect 4934 4560 4964 4594
rect 4964 4560 4968 4594
rect 5006 4560 5032 4594
rect 5032 4560 5040 4594
rect 5078 4560 5100 4594
rect 5100 4560 5112 4594
rect 5150 4560 5168 4594
rect 5168 4560 5184 4594
rect 5222 4560 5236 4594
rect 5236 4560 5256 4594
rect 5294 4560 5304 4594
rect 5304 4560 5328 4594
rect 5366 4560 5372 4594
rect 5372 4560 5400 4594
rect 5438 4560 5440 4594
rect 5440 4560 5472 4594
rect 5510 4560 5542 4594
rect 5542 4560 5544 4594
rect 5582 4560 5610 4594
rect 5610 4560 5616 4594
rect 5654 4560 5678 4594
rect 5678 4560 5688 4594
rect 5726 4560 5746 4594
rect 5746 4560 5760 4594
rect 5798 4560 5814 4594
rect 5814 4560 5832 4594
rect 5870 4560 5882 4594
rect 5882 4560 5904 4594
rect 5942 4560 5950 4594
rect 5950 4560 5976 4594
rect 6014 4560 6018 4594
rect 6018 4560 6048 4594
rect 6086 4560 6120 4594
rect 6158 4560 6188 4594
rect 6188 4560 6192 4594
rect 6230 4560 6256 4594
rect 6256 4560 6264 4594
rect 6302 4560 6324 4594
rect 6324 4560 6336 4594
rect 6374 4560 6392 4594
rect 6392 4560 6408 4594
rect 6446 4560 6460 4594
rect 6460 4560 6480 4594
rect 6518 4560 6528 4594
rect 6528 4560 6552 4594
rect 6590 4560 6596 4594
rect 6596 4560 6624 4594
rect 6662 4560 6664 4594
rect 6664 4560 6696 4594
rect 6734 4560 6766 4594
rect 6766 4560 6768 4594
rect 6806 4560 6834 4594
rect 6834 4560 6840 4594
rect 6878 4560 6902 4594
rect 6902 4560 6912 4594
rect 6950 4560 6970 4594
rect 6970 4560 6984 4594
rect 7022 4560 7038 4594
rect 7038 4560 7056 4594
rect 7094 4560 7106 4594
rect 7106 4560 7128 4594
rect 7166 4560 7174 4594
rect 7174 4560 7200 4594
rect 7238 4560 7242 4594
rect 7242 4560 7272 4594
rect 7310 4560 7344 4594
rect 7382 4560 7412 4594
rect 7412 4560 7416 4594
rect 7454 4560 7480 4594
rect 7480 4560 7488 4594
rect 7526 4560 7548 4594
rect 7548 4560 7560 4594
rect 7598 4560 7616 4594
rect 7616 4560 7632 4594
rect 7670 4560 7684 4594
rect 7684 4560 7704 4594
rect 7742 4560 7752 4594
rect 7752 4560 7776 4594
rect 7814 4560 7820 4594
rect 7820 4560 7848 4594
rect 7886 4560 7888 4594
rect 7888 4560 7920 4594
rect 7958 4560 7990 4594
rect 7990 4560 7992 4594
rect 8030 4560 8058 4594
rect 8058 4560 8064 4594
rect 8102 4560 8126 4594
rect 8126 4560 8136 4594
rect 8174 4560 8194 4594
rect 8194 4560 8208 4594
rect 8246 4560 8262 4594
rect 8262 4560 8280 4594
rect 8318 4560 8330 4594
rect 8330 4560 8352 4594
rect 8390 4560 8398 4594
rect 8398 4560 8424 4594
rect 8462 4560 8466 4594
rect 8466 4560 8496 4594
rect 8534 4560 8568 4594
rect 8606 4560 8636 4594
rect 8636 4560 8640 4594
rect 8678 4560 8704 4594
rect 8704 4560 8712 4594
rect 8750 4560 8772 4594
rect 8772 4560 8784 4594
rect 8822 4560 8840 4594
rect 8840 4560 8856 4594
rect 8894 4560 8908 4594
rect 8908 4560 8928 4594
rect 8966 4560 8976 4594
rect 8976 4560 9000 4594
rect 9038 4560 9044 4594
rect 9044 4560 9072 4594
rect 9110 4560 9112 4594
rect 9112 4560 9144 4594
rect 9182 4560 9214 4594
rect 9214 4560 9216 4594
rect 9254 4560 9282 4594
rect 9282 4560 9288 4594
rect 9326 4560 9350 4594
rect 9350 4560 9360 4594
rect 9398 4560 9418 4594
rect 9418 4560 9432 4594
rect 9470 4560 9486 4594
rect 9486 4560 9504 4594
rect 9542 4560 9554 4594
rect 9554 4560 9576 4594
rect 9614 4560 9622 4594
rect 9622 4560 9648 4594
rect 9686 4560 9690 4594
rect 9690 4560 9720 4594
rect 9758 4560 9792 4594
rect 9830 4560 9860 4594
rect 9860 4560 9864 4594
rect 9902 4560 9928 4594
rect 9928 4560 9936 4594
rect 9974 4560 9996 4594
rect 9996 4560 10008 4594
rect 10046 4560 10064 4594
rect 10064 4560 10080 4594
rect 10118 4560 10132 4594
rect 10132 4560 10152 4594
rect 10190 4560 10200 4594
rect 10200 4560 10224 4594
rect 10262 4560 10268 4594
rect 10268 4560 10296 4594
rect 10334 4560 10336 4594
rect 10336 4560 10368 4594
rect 10406 4560 10438 4594
rect 10438 4560 10440 4594
rect 10478 4560 10506 4594
rect 10506 4560 10512 4594
rect 10550 4560 10574 4594
rect 10574 4560 10584 4594
rect 10622 4560 10642 4594
rect 10642 4560 10656 4594
rect 10694 4560 10710 4594
rect 10710 4560 10728 4594
rect 10766 4560 10778 4594
rect 10778 4560 10800 4594
rect 10838 4560 10846 4594
rect 10846 4560 10872 4594
rect 10910 4560 10914 4594
rect 10914 4560 10944 4594
rect 10982 4560 11016 4594
rect 11054 4560 11084 4594
rect 11084 4560 11088 4594
rect 38 16 68 50
rect 68 16 72 50
rect 110 16 136 50
rect 136 16 144 50
rect 182 16 204 50
rect 204 16 216 50
rect 254 16 272 50
rect 272 16 288 50
rect 326 16 340 50
rect 340 16 360 50
rect 398 16 408 50
rect 408 16 432 50
rect 470 16 476 50
rect 476 16 504 50
rect 542 16 544 50
rect 544 16 576 50
rect 614 16 646 50
rect 646 16 648 50
rect 686 16 714 50
rect 714 16 720 50
rect 758 16 782 50
rect 782 16 792 50
rect 830 16 850 50
rect 850 16 864 50
rect 902 16 918 50
rect 918 16 936 50
rect 974 16 986 50
rect 986 16 1008 50
rect 1046 16 1054 50
rect 1054 16 1080 50
rect 1118 16 1122 50
rect 1122 16 1152 50
rect 1190 16 1224 50
rect 1262 16 1292 50
rect 1292 16 1296 50
rect 1334 16 1360 50
rect 1360 16 1368 50
rect 1406 16 1428 50
rect 1428 16 1440 50
rect 1478 16 1496 50
rect 1496 16 1512 50
rect 1550 16 1564 50
rect 1564 16 1584 50
rect 1622 16 1632 50
rect 1632 16 1656 50
rect 1694 16 1700 50
rect 1700 16 1728 50
rect 1766 16 1768 50
rect 1768 16 1800 50
rect 1838 16 1870 50
rect 1870 16 1872 50
rect 1910 16 1938 50
rect 1938 16 1944 50
rect 1982 16 2006 50
rect 2006 16 2016 50
rect 2054 16 2074 50
rect 2074 16 2088 50
rect 2126 16 2142 50
rect 2142 16 2160 50
rect 2198 16 2210 50
rect 2210 16 2232 50
rect 2270 16 2278 50
rect 2278 16 2304 50
rect 2342 16 2346 50
rect 2346 16 2376 50
rect 2414 16 2448 50
rect 2486 16 2516 50
rect 2516 16 2520 50
rect 2558 16 2584 50
rect 2584 16 2592 50
rect 2630 16 2652 50
rect 2652 16 2664 50
rect 2702 16 2720 50
rect 2720 16 2736 50
rect 2774 16 2788 50
rect 2788 16 2808 50
rect 2846 16 2856 50
rect 2856 16 2880 50
rect 2918 16 2924 50
rect 2924 16 2952 50
rect 2990 16 2992 50
rect 2992 16 3024 50
rect 3062 16 3094 50
rect 3094 16 3096 50
rect 3134 16 3162 50
rect 3162 16 3168 50
rect 3206 16 3230 50
rect 3230 16 3240 50
rect 3278 16 3298 50
rect 3298 16 3312 50
rect 3350 16 3366 50
rect 3366 16 3384 50
rect 3422 16 3434 50
rect 3434 16 3456 50
rect 3494 16 3502 50
rect 3502 16 3528 50
rect 3566 16 3570 50
rect 3570 16 3600 50
rect 3638 16 3672 50
rect 3710 16 3740 50
rect 3740 16 3744 50
rect 3782 16 3808 50
rect 3808 16 3816 50
rect 3854 16 3876 50
rect 3876 16 3888 50
rect 3926 16 3944 50
rect 3944 16 3960 50
rect 3998 16 4012 50
rect 4012 16 4032 50
rect 4070 16 4080 50
rect 4080 16 4104 50
rect 4142 16 4148 50
rect 4148 16 4176 50
rect 4214 16 4216 50
rect 4216 16 4248 50
rect 4286 16 4318 50
rect 4318 16 4320 50
rect 4358 16 4386 50
rect 4386 16 4392 50
rect 4430 16 4454 50
rect 4454 16 4464 50
rect 4502 16 4522 50
rect 4522 16 4536 50
rect 4574 16 4590 50
rect 4590 16 4608 50
rect 4646 16 4658 50
rect 4658 16 4680 50
rect 4718 16 4726 50
rect 4726 16 4752 50
rect 4790 16 4794 50
rect 4794 16 4824 50
rect 4862 16 4896 50
rect 4934 16 4964 50
rect 4964 16 4968 50
rect 5006 16 5032 50
rect 5032 16 5040 50
rect 5078 16 5100 50
rect 5100 16 5112 50
rect 5150 16 5168 50
rect 5168 16 5184 50
rect 5222 16 5236 50
rect 5236 16 5256 50
rect 5294 16 5304 50
rect 5304 16 5328 50
rect 5366 16 5372 50
rect 5372 16 5400 50
rect 5438 16 5440 50
rect 5440 16 5472 50
rect 5510 16 5542 50
rect 5542 16 5544 50
rect 5582 16 5610 50
rect 5610 16 5616 50
rect 5654 16 5678 50
rect 5678 16 5688 50
rect 5726 16 5746 50
rect 5746 16 5760 50
rect 5798 16 5814 50
rect 5814 16 5832 50
rect 5870 16 5882 50
rect 5882 16 5904 50
rect 5942 16 5950 50
rect 5950 16 5976 50
rect 6014 16 6018 50
rect 6018 16 6048 50
rect 6086 16 6120 50
rect 6158 16 6188 50
rect 6188 16 6192 50
rect 6230 16 6256 50
rect 6256 16 6264 50
rect 6302 16 6324 50
rect 6324 16 6336 50
rect 6374 16 6392 50
rect 6392 16 6408 50
rect 6446 16 6460 50
rect 6460 16 6480 50
rect 6518 16 6528 50
rect 6528 16 6552 50
rect 6590 16 6596 50
rect 6596 16 6624 50
rect 6662 16 6664 50
rect 6664 16 6696 50
rect 6734 16 6766 50
rect 6766 16 6768 50
rect 6806 16 6834 50
rect 6834 16 6840 50
rect 6878 16 6902 50
rect 6902 16 6912 50
rect 6950 16 6970 50
rect 6970 16 6984 50
rect 7022 16 7038 50
rect 7038 16 7056 50
rect 7094 16 7106 50
rect 7106 16 7128 50
rect 7166 16 7174 50
rect 7174 16 7200 50
rect 7238 16 7242 50
rect 7242 16 7272 50
rect 7310 16 7344 50
rect 7382 16 7412 50
rect 7412 16 7416 50
rect 7454 16 7480 50
rect 7480 16 7488 50
rect 7526 16 7548 50
rect 7548 16 7560 50
rect 7598 16 7616 50
rect 7616 16 7632 50
rect 7670 16 7684 50
rect 7684 16 7704 50
rect 7742 16 7752 50
rect 7752 16 7776 50
rect 7814 16 7820 50
rect 7820 16 7848 50
rect 7886 16 7888 50
rect 7888 16 7920 50
rect 7958 16 7990 50
rect 7990 16 7992 50
rect 8030 16 8058 50
rect 8058 16 8064 50
rect 8102 16 8126 50
rect 8126 16 8136 50
rect 8174 16 8194 50
rect 8194 16 8208 50
rect 8246 16 8262 50
rect 8262 16 8280 50
rect 8318 16 8330 50
rect 8330 16 8352 50
rect 8390 16 8398 50
rect 8398 16 8424 50
rect 8462 16 8466 50
rect 8466 16 8496 50
rect 8534 16 8568 50
rect 8606 16 8636 50
rect 8636 16 8640 50
rect 8678 16 8704 50
rect 8704 16 8712 50
rect 8750 16 8772 50
rect 8772 16 8784 50
rect 8822 16 8840 50
rect 8840 16 8856 50
rect 8894 16 8908 50
rect 8908 16 8928 50
rect 8966 16 8976 50
rect 8976 16 9000 50
rect 9038 16 9044 50
rect 9044 16 9072 50
rect 9110 16 9112 50
rect 9112 16 9144 50
rect 9182 16 9214 50
rect 9214 16 9216 50
rect 9254 16 9282 50
rect 9282 16 9288 50
rect 9326 16 9350 50
rect 9350 16 9360 50
rect 9398 16 9418 50
rect 9418 16 9432 50
rect 9470 16 9486 50
rect 9486 16 9504 50
rect 9542 16 9554 50
rect 9554 16 9576 50
rect 9614 16 9622 50
rect 9622 16 9648 50
rect 9686 16 9690 50
rect 9690 16 9720 50
rect 9758 16 9792 50
rect 9830 16 9860 50
rect 9860 16 9864 50
rect 9902 16 9928 50
rect 9928 16 9936 50
rect 9974 16 9996 50
rect 9996 16 10008 50
rect 10046 16 10064 50
rect 10064 16 10080 50
rect 10118 16 10132 50
rect 10132 16 10152 50
rect 10190 16 10200 50
rect 10200 16 10224 50
rect 10262 16 10268 50
rect 10268 16 10296 50
rect 10334 16 10336 50
rect 10336 16 10368 50
rect 10406 16 10438 50
rect 10438 16 10440 50
rect 10478 16 10506 50
rect 10506 16 10512 50
rect 10550 16 10574 50
rect 10574 16 10584 50
rect 10622 16 10642 50
rect 10642 16 10656 50
rect 10694 16 10710 50
rect 10710 16 10728 50
rect 10766 16 10778 50
rect 10778 16 10800 50
rect 10838 16 10846 50
rect 10846 16 10872 50
rect 10910 16 10914 50
rect 10914 16 10944 50
rect 10982 16 11016 50
rect 11054 16 11084 50
rect 11084 16 11088 50
<< metal1 >>
rect 0 4603 11146 4610
rect 0 4594 68 4603
rect 120 4594 132 4603
rect 184 4594 292 4603
rect 344 4594 356 4603
rect 408 4594 516 4603
rect 568 4594 580 4603
rect 632 4594 740 4603
rect 0 4560 38 4594
rect 216 4560 254 4594
rect 288 4560 292 4594
rect 432 4560 470 4594
rect 504 4560 516 4594
rect 576 4560 580 4594
rect 648 4560 686 4594
rect 720 4560 740 4594
rect 0 4551 68 4560
rect 120 4551 132 4560
rect 184 4551 292 4560
rect 344 4551 356 4560
rect 408 4551 516 4560
rect 568 4551 580 4560
rect 632 4551 740 4560
rect 792 4551 804 4603
rect 856 4594 964 4603
rect 864 4560 902 4594
rect 936 4560 964 4594
rect 856 4551 964 4560
rect 1016 4551 1028 4603
rect 1080 4594 1188 4603
rect 1080 4560 1118 4594
rect 1152 4560 1188 4594
rect 1080 4551 1188 4560
rect 1240 4551 1252 4603
rect 1304 4594 1412 4603
rect 1304 4560 1334 4594
rect 1368 4560 1406 4594
rect 1304 4551 1412 4560
rect 1464 4551 1476 4603
rect 1528 4594 1636 4603
rect 1688 4594 1700 4603
rect 1752 4594 1860 4603
rect 1912 4594 1924 4603
rect 1976 4594 2084 4603
rect 2136 4594 2148 4603
rect 2200 4594 2308 4603
rect 2360 4594 2372 4603
rect 2424 4594 2532 4603
rect 2584 4594 2596 4603
rect 2648 4594 2756 4603
rect 1528 4560 1550 4594
rect 1584 4560 1622 4594
rect 1688 4560 1694 4594
rect 1752 4560 1766 4594
rect 1800 4560 1838 4594
rect 1976 4560 1982 4594
rect 2016 4560 2054 4594
rect 2232 4560 2270 4594
rect 2304 4560 2308 4594
rect 2448 4560 2486 4594
rect 2520 4560 2532 4594
rect 2592 4560 2596 4594
rect 2664 4560 2702 4594
rect 2736 4560 2756 4594
rect 1528 4551 1636 4560
rect 1688 4551 1700 4560
rect 1752 4551 1860 4560
rect 1912 4551 1924 4560
rect 1976 4551 2084 4560
rect 2136 4551 2148 4560
rect 2200 4551 2308 4560
rect 2360 4551 2372 4560
rect 2424 4551 2532 4560
rect 2584 4551 2596 4560
rect 2648 4551 2756 4560
rect 2808 4551 2820 4603
rect 2872 4594 2980 4603
rect 2880 4560 2918 4594
rect 2952 4560 2980 4594
rect 2872 4551 2980 4560
rect 3032 4551 3044 4603
rect 3096 4594 3204 4603
rect 3096 4560 3134 4594
rect 3168 4560 3204 4594
rect 3096 4551 3204 4560
rect 3256 4551 3268 4603
rect 3320 4594 3428 4603
rect 3320 4560 3350 4594
rect 3384 4560 3422 4594
rect 3320 4551 3428 4560
rect 3480 4551 3492 4603
rect 3544 4594 3652 4603
rect 3704 4594 3716 4603
rect 3768 4594 3876 4603
rect 3928 4594 3940 4603
rect 3992 4594 4100 4603
rect 4152 4594 4164 4603
rect 4216 4594 4324 4603
rect 4376 4594 4388 4603
rect 4440 4594 4548 4603
rect 4600 4594 4612 4603
rect 4664 4594 4772 4603
rect 3544 4560 3566 4594
rect 3600 4560 3638 4594
rect 3704 4560 3710 4594
rect 3768 4560 3782 4594
rect 3816 4560 3854 4594
rect 3992 4560 3998 4594
rect 4032 4560 4070 4594
rect 4248 4560 4286 4594
rect 4320 4560 4324 4594
rect 4464 4560 4502 4594
rect 4536 4560 4548 4594
rect 4608 4560 4612 4594
rect 4680 4560 4718 4594
rect 4752 4560 4772 4594
rect 3544 4551 3652 4560
rect 3704 4551 3716 4560
rect 3768 4551 3876 4560
rect 3928 4551 3940 4560
rect 3992 4551 4100 4560
rect 4152 4551 4164 4560
rect 4216 4551 4324 4560
rect 4376 4551 4388 4560
rect 4440 4551 4548 4560
rect 4600 4551 4612 4560
rect 4664 4551 4772 4560
rect 4824 4551 4836 4603
rect 4888 4594 4996 4603
rect 4896 4560 4934 4594
rect 4968 4560 4996 4594
rect 4888 4551 4996 4560
rect 5048 4551 5060 4603
rect 5112 4594 5220 4603
rect 5112 4560 5150 4594
rect 5184 4560 5220 4594
rect 5112 4551 5220 4560
rect 5272 4551 5284 4603
rect 5336 4594 5444 4603
rect 5336 4560 5366 4594
rect 5400 4560 5438 4594
rect 5336 4551 5444 4560
rect 5496 4551 5508 4603
rect 5560 4594 5668 4603
rect 5720 4594 5732 4603
rect 5784 4594 5892 4603
rect 5944 4594 5956 4603
rect 6008 4594 6116 4603
rect 6168 4594 6180 4603
rect 6232 4594 6340 4603
rect 6392 4594 6404 4603
rect 6456 4594 6564 4603
rect 6616 4594 6628 4603
rect 6680 4594 6788 4603
rect 5560 4560 5582 4594
rect 5616 4560 5654 4594
rect 5720 4560 5726 4594
rect 5784 4560 5798 4594
rect 5832 4560 5870 4594
rect 6008 4560 6014 4594
rect 6048 4560 6086 4594
rect 6264 4560 6302 4594
rect 6336 4560 6340 4594
rect 6480 4560 6518 4594
rect 6552 4560 6564 4594
rect 6624 4560 6628 4594
rect 6696 4560 6734 4594
rect 6768 4560 6788 4594
rect 5560 4551 5668 4560
rect 5720 4551 5732 4560
rect 5784 4551 5892 4560
rect 5944 4551 5956 4560
rect 6008 4551 6116 4560
rect 6168 4551 6180 4560
rect 6232 4551 6340 4560
rect 6392 4551 6404 4560
rect 6456 4551 6564 4560
rect 6616 4551 6628 4560
rect 6680 4551 6788 4560
rect 6840 4551 6852 4603
rect 6904 4594 7012 4603
rect 6912 4560 6950 4594
rect 6984 4560 7012 4594
rect 6904 4551 7012 4560
rect 7064 4551 7076 4603
rect 7128 4594 7236 4603
rect 7128 4560 7166 4594
rect 7200 4560 7236 4594
rect 7128 4551 7236 4560
rect 7288 4551 7300 4603
rect 7352 4594 7460 4603
rect 7352 4560 7382 4594
rect 7416 4560 7454 4594
rect 7352 4551 7460 4560
rect 7512 4551 7524 4603
rect 7576 4594 7684 4603
rect 7736 4594 7748 4603
rect 7800 4594 7908 4603
rect 7960 4594 7972 4603
rect 8024 4594 8132 4603
rect 8184 4594 8196 4603
rect 8248 4594 8356 4603
rect 8408 4594 8420 4603
rect 8472 4594 8580 4603
rect 8632 4594 8644 4603
rect 8696 4594 8804 4603
rect 7576 4560 7598 4594
rect 7632 4560 7670 4594
rect 7736 4560 7742 4594
rect 7800 4560 7814 4594
rect 7848 4560 7886 4594
rect 8024 4560 8030 4594
rect 8064 4560 8102 4594
rect 8280 4560 8318 4594
rect 8352 4560 8356 4594
rect 8496 4560 8534 4594
rect 8568 4560 8580 4594
rect 8640 4560 8644 4594
rect 8712 4560 8750 4594
rect 8784 4560 8804 4594
rect 7576 4551 7684 4560
rect 7736 4551 7748 4560
rect 7800 4551 7908 4560
rect 7960 4551 7972 4560
rect 8024 4551 8132 4560
rect 8184 4551 8196 4560
rect 8248 4551 8356 4560
rect 8408 4551 8420 4560
rect 8472 4551 8580 4560
rect 8632 4551 8644 4560
rect 8696 4551 8804 4560
rect 8856 4551 8868 4603
rect 8920 4594 9028 4603
rect 8928 4560 8966 4594
rect 9000 4560 9028 4594
rect 8920 4551 9028 4560
rect 9080 4551 9092 4603
rect 9144 4594 9252 4603
rect 9144 4560 9182 4594
rect 9216 4560 9252 4594
rect 9144 4551 9252 4560
rect 9304 4551 9316 4603
rect 9368 4594 9476 4603
rect 9368 4560 9398 4594
rect 9432 4560 9470 4594
rect 9368 4551 9476 4560
rect 9528 4551 9540 4603
rect 9592 4594 9700 4603
rect 9752 4594 9764 4603
rect 9816 4594 9924 4603
rect 9976 4594 9988 4603
rect 10040 4594 10148 4603
rect 10200 4594 10212 4603
rect 10264 4594 10372 4603
rect 10424 4594 10436 4603
rect 10488 4594 10596 4603
rect 10648 4594 10660 4603
rect 10712 4594 10820 4603
rect 9592 4560 9614 4594
rect 9648 4560 9686 4594
rect 9752 4560 9758 4594
rect 9816 4560 9830 4594
rect 9864 4560 9902 4594
rect 10040 4560 10046 4594
rect 10080 4560 10118 4594
rect 10296 4560 10334 4594
rect 10368 4560 10372 4594
rect 10512 4560 10550 4594
rect 10584 4560 10596 4594
rect 10656 4560 10660 4594
rect 10728 4560 10766 4594
rect 10800 4560 10820 4594
rect 9592 4551 9700 4560
rect 9752 4551 9764 4560
rect 9816 4551 9924 4560
rect 9976 4551 9988 4560
rect 10040 4551 10148 4560
rect 10200 4551 10212 4560
rect 10264 4551 10372 4560
rect 10424 4551 10436 4560
rect 10488 4551 10596 4560
rect 10648 4551 10660 4560
rect 10712 4551 10820 4560
rect 10872 4551 10884 4603
rect 10936 4594 11146 4603
rect 10944 4560 10982 4594
rect 11016 4560 11054 4594
rect 11088 4560 11146 4594
rect 10936 4551 11146 4560
rect 0 4544 11146 4551
rect 0 94 28 4544
rect 56 66 84 4516
rect 112 94 140 4544
rect 168 66 196 4516
rect 224 94 252 4544
rect 280 66 308 4516
rect 336 94 364 4544
rect 392 66 420 4516
rect 448 94 476 4544
rect 504 66 532 4516
rect 560 94 588 4544
rect 616 66 644 4516
rect 672 94 700 4544
rect 728 66 756 4516
rect 784 94 812 4544
rect 840 66 868 4516
rect 896 94 924 4544
rect 952 66 980 4516
rect 1008 94 1036 4544
rect 1064 66 1092 4516
rect 1120 94 1148 4544
rect 1176 66 1204 4516
rect 1232 94 1260 4544
rect 1288 66 1316 4516
rect 1344 94 1372 4544
rect 1400 66 1428 4516
rect 1456 94 1484 4544
rect 1512 66 1540 4516
rect 1568 94 1596 4544
rect 1624 66 1652 4516
rect 1680 94 1708 4544
rect 1736 66 1764 4516
rect 1792 94 1820 4544
rect 1848 66 1876 4516
rect 1904 94 1932 4544
rect 1960 66 1988 4516
rect 2016 94 2044 4544
rect 2072 66 2100 4516
rect 2128 94 2156 4544
rect 2184 66 2212 4516
rect 2240 94 2268 4544
rect 2296 66 2324 4516
rect 2352 94 2380 4544
rect 2408 66 2436 4516
rect 2464 94 2492 4544
rect 2520 66 2548 4516
rect 2576 94 2604 4544
rect 2632 66 2660 4516
rect 2688 94 2716 4544
rect 2744 66 2772 4516
rect 2800 94 2828 4544
rect 2856 66 2884 4516
rect 2912 94 2940 4544
rect 2968 66 2996 4516
rect 3024 94 3052 4544
rect 3080 66 3108 4516
rect 3136 94 3164 4544
rect 3192 66 3220 4516
rect 3248 94 3276 4544
rect 3304 66 3332 4516
rect 3360 94 3388 4544
rect 3416 66 3444 4516
rect 3472 94 3500 4544
rect 3528 66 3556 4516
rect 3584 94 3612 4544
rect 3640 66 3668 4516
rect 3696 94 3724 4544
rect 3752 66 3780 4516
rect 3808 94 3836 4544
rect 3864 66 3892 4516
rect 3920 94 3948 4544
rect 3976 66 4004 4516
rect 4032 94 4060 4544
rect 4088 66 4116 4516
rect 4144 94 4172 4544
rect 4200 66 4228 4516
rect 4256 94 4284 4544
rect 4312 66 4340 4516
rect 4368 94 4396 4544
rect 4424 66 4452 4516
rect 4480 94 4508 4544
rect 4536 66 4564 4516
rect 4592 94 4620 4544
rect 4648 66 4676 4516
rect 4704 94 4732 4544
rect 4760 66 4788 4516
rect 4816 94 4844 4544
rect 4872 66 4900 4516
rect 4928 94 4956 4544
rect 4984 66 5012 4516
rect 5040 94 5068 4544
rect 5096 66 5124 4516
rect 5152 94 5180 4544
rect 5208 66 5236 4516
rect 5264 94 5292 4544
rect 5320 66 5348 4516
rect 5376 94 5404 4544
rect 5432 66 5460 4516
rect 5488 94 5516 4544
rect 5544 66 5572 4516
rect 5600 94 5628 4544
rect 5656 66 5684 4516
rect 5712 94 5740 4544
rect 5768 66 5796 4516
rect 5824 94 5852 4544
rect 5880 66 5908 4516
rect 5936 94 5964 4544
rect 5992 66 6020 4516
rect 6048 94 6076 4544
rect 6104 66 6132 4516
rect 6160 94 6188 4544
rect 6216 66 6244 4516
rect 6272 94 6300 4544
rect 6328 66 6356 4516
rect 6384 94 6412 4544
rect 6440 66 6468 4516
rect 6496 94 6524 4544
rect 6552 66 6580 4516
rect 6608 94 6636 4544
rect 6664 66 6692 4516
rect 6720 94 6748 4544
rect 6776 66 6804 4516
rect 6832 94 6860 4544
rect 6888 66 6916 4516
rect 6944 94 6972 4544
rect 7000 66 7028 4516
rect 7056 94 7084 4544
rect 7112 66 7140 4516
rect 7168 94 7196 4544
rect 7224 66 7252 4516
rect 7280 94 7308 4544
rect 7336 66 7364 4516
rect 7392 94 7420 4544
rect 7448 66 7476 4516
rect 7504 94 7532 4544
rect 7560 66 7588 4516
rect 7616 94 7644 4544
rect 7672 66 7700 4516
rect 7728 94 7756 4544
rect 7784 66 7812 4516
rect 7840 94 7868 4544
rect 7896 66 7924 4516
rect 7952 94 7980 4544
rect 8008 66 8036 4516
rect 8064 94 8092 4544
rect 8120 66 8148 4516
rect 8176 94 8204 4544
rect 8232 66 8260 4516
rect 8288 94 8316 4544
rect 8344 66 8372 4516
rect 8400 94 8428 4544
rect 8456 66 8484 4516
rect 8512 94 8540 4544
rect 8568 66 8596 4516
rect 8624 94 8652 4544
rect 8680 66 8708 4516
rect 8736 94 8764 4544
rect 8792 66 8820 4516
rect 8848 94 8876 4544
rect 8904 66 8932 4516
rect 8960 94 8988 4544
rect 9016 66 9044 4516
rect 9072 94 9100 4544
rect 9128 66 9156 4516
rect 9184 94 9212 4544
rect 9240 66 9268 4516
rect 9296 94 9324 4544
rect 9352 66 9380 4516
rect 9408 94 9436 4544
rect 9464 66 9492 4516
rect 9520 94 9548 4544
rect 9576 66 9604 4516
rect 9632 94 9660 4544
rect 9688 66 9716 4516
rect 9744 94 9772 4544
rect 9800 66 9828 4516
rect 9856 94 9884 4544
rect 9912 66 9940 4516
rect 9968 94 9996 4544
rect 10024 66 10052 4516
rect 10080 94 10108 4544
rect 10136 66 10164 4516
rect 10192 94 10220 4544
rect 10248 66 10276 4516
rect 10304 94 10332 4544
rect 10360 66 10388 4516
rect 10416 94 10444 4544
rect 10472 66 10500 4516
rect 10528 94 10556 4544
rect 10584 66 10612 4516
rect 10640 94 10668 4544
rect 10696 66 10724 4516
rect 10752 94 10780 4544
rect 10808 66 10836 4516
rect 10864 94 10892 4544
rect 10920 66 10948 4516
rect 10976 94 11004 4544
rect 11032 66 11060 4516
rect 11088 94 11146 4544
rect 0 59 11146 66
rect 0 7 24 59
rect 76 7 88 59
rect 140 50 236 59
rect 144 16 182 50
rect 216 16 236 50
rect 140 7 236 16
rect 288 7 300 59
rect 352 50 460 59
rect 360 16 398 50
rect 432 16 460 50
rect 352 7 460 16
rect 512 7 524 59
rect 576 50 684 59
rect 576 16 614 50
rect 648 16 684 50
rect 576 7 684 16
rect 736 7 748 59
rect 800 50 908 59
rect 800 16 830 50
rect 864 16 902 50
rect 800 7 908 16
rect 960 7 972 59
rect 1024 50 1132 59
rect 1184 50 1196 59
rect 1248 50 1356 59
rect 1408 50 1420 59
rect 1472 50 1580 59
rect 1632 50 1644 59
rect 1696 50 1804 59
rect 1856 50 1868 59
rect 1920 50 2028 59
rect 2080 50 2092 59
rect 2144 50 2252 59
rect 1024 16 1046 50
rect 1080 16 1118 50
rect 1184 16 1190 50
rect 1248 16 1262 50
rect 1296 16 1334 50
rect 1472 16 1478 50
rect 1512 16 1550 50
rect 1728 16 1766 50
rect 1800 16 1804 50
rect 1944 16 1982 50
rect 2016 16 2028 50
rect 2088 16 2092 50
rect 2160 16 2198 50
rect 2232 16 2252 50
rect 1024 7 1132 16
rect 1184 7 1196 16
rect 1248 7 1356 16
rect 1408 7 1420 16
rect 1472 7 1580 16
rect 1632 7 1644 16
rect 1696 7 1804 16
rect 1856 7 1868 16
rect 1920 7 2028 16
rect 2080 7 2092 16
rect 2144 7 2252 16
rect 2304 7 2316 59
rect 2368 50 2476 59
rect 2376 16 2414 50
rect 2448 16 2476 50
rect 2368 7 2476 16
rect 2528 7 2540 59
rect 2592 50 2700 59
rect 2592 16 2630 50
rect 2664 16 2700 50
rect 2592 7 2700 16
rect 2752 7 2764 59
rect 2816 50 2924 59
rect 2816 16 2846 50
rect 2880 16 2918 50
rect 2816 7 2924 16
rect 2976 7 2988 59
rect 3040 50 3148 59
rect 3200 50 3212 59
rect 3264 50 3372 59
rect 3424 50 3436 59
rect 3488 50 3596 59
rect 3648 50 3660 59
rect 3712 50 3820 59
rect 3872 50 3884 59
rect 3936 50 4044 59
rect 4096 50 4108 59
rect 4160 50 4268 59
rect 3040 16 3062 50
rect 3096 16 3134 50
rect 3200 16 3206 50
rect 3264 16 3278 50
rect 3312 16 3350 50
rect 3488 16 3494 50
rect 3528 16 3566 50
rect 3744 16 3782 50
rect 3816 16 3820 50
rect 3960 16 3998 50
rect 4032 16 4044 50
rect 4104 16 4108 50
rect 4176 16 4214 50
rect 4248 16 4268 50
rect 3040 7 3148 16
rect 3200 7 3212 16
rect 3264 7 3372 16
rect 3424 7 3436 16
rect 3488 7 3596 16
rect 3648 7 3660 16
rect 3712 7 3820 16
rect 3872 7 3884 16
rect 3936 7 4044 16
rect 4096 7 4108 16
rect 4160 7 4268 16
rect 4320 7 4332 59
rect 4384 50 4492 59
rect 4392 16 4430 50
rect 4464 16 4492 50
rect 4384 7 4492 16
rect 4544 7 4556 59
rect 4608 50 4716 59
rect 4608 16 4646 50
rect 4680 16 4716 50
rect 4608 7 4716 16
rect 4768 7 4780 59
rect 4832 50 4940 59
rect 4832 16 4862 50
rect 4896 16 4934 50
rect 4832 7 4940 16
rect 4992 7 5004 59
rect 5056 50 5164 59
rect 5216 50 5228 59
rect 5280 50 5388 59
rect 5440 50 5452 59
rect 5504 50 5612 59
rect 5664 50 5676 59
rect 5728 50 5836 59
rect 5888 50 5900 59
rect 5952 50 6060 59
rect 6112 50 6124 59
rect 6176 50 6284 59
rect 5056 16 5078 50
rect 5112 16 5150 50
rect 5216 16 5222 50
rect 5280 16 5294 50
rect 5328 16 5366 50
rect 5504 16 5510 50
rect 5544 16 5582 50
rect 5760 16 5798 50
rect 5832 16 5836 50
rect 5976 16 6014 50
rect 6048 16 6060 50
rect 6120 16 6124 50
rect 6192 16 6230 50
rect 6264 16 6284 50
rect 5056 7 5164 16
rect 5216 7 5228 16
rect 5280 7 5388 16
rect 5440 7 5452 16
rect 5504 7 5612 16
rect 5664 7 5676 16
rect 5728 7 5836 16
rect 5888 7 5900 16
rect 5952 7 6060 16
rect 6112 7 6124 16
rect 6176 7 6284 16
rect 6336 7 6348 59
rect 6400 50 6508 59
rect 6408 16 6446 50
rect 6480 16 6508 50
rect 6400 7 6508 16
rect 6560 7 6572 59
rect 6624 50 6732 59
rect 6624 16 6662 50
rect 6696 16 6732 50
rect 6624 7 6732 16
rect 6784 7 6796 59
rect 6848 50 6956 59
rect 6848 16 6878 50
rect 6912 16 6950 50
rect 6848 7 6956 16
rect 7008 7 7020 59
rect 7072 50 7180 59
rect 7232 50 7244 59
rect 7296 50 7404 59
rect 7456 50 7468 59
rect 7520 50 7628 59
rect 7680 50 7692 59
rect 7744 50 7852 59
rect 7904 50 7916 59
rect 7968 50 8076 59
rect 8128 50 8140 59
rect 8192 50 8300 59
rect 7072 16 7094 50
rect 7128 16 7166 50
rect 7232 16 7238 50
rect 7296 16 7310 50
rect 7344 16 7382 50
rect 7520 16 7526 50
rect 7560 16 7598 50
rect 7776 16 7814 50
rect 7848 16 7852 50
rect 7992 16 8030 50
rect 8064 16 8076 50
rect 8136 16 8140 50
rect 8208 16 8246 50
rect 8280 16 8300 50
rect 7072 7 7180 16
rect 7232 7 7244 16
rect 7296 7 7404 16
rect 7456 7 7468 16
rect 7520 7 7628 16
rect 7680 7 7692 16
rect 7744 7 7852 16
rect 7904 7 7916 16
rect 7968 7 8076 16
rect 8128 7 8140 16
rect 8192 7 8300 16
rect 8352 7 8364 59
rect 8416 50 8524 59
rect 8424 16 8462 50
rect 8496 16 8524 50
rect 8416 7 8524 16
rect 8576 7 8588 59
rect 8640 50 8748 59
rect 8640 16 8678 50
rect 8712 16 8748 50
rect 8640 7 8748 16
rect 8800 7 8812 59
rect 8864 50 8972 59
rect 8864 16 8894 50
rect 8928 16 8966 50
rect 8864 7 8972 16
rect 9024 7 9036 59
rect 9088 50 9196 59
rect 9248 50 9260 59
rect 9312 50 9420 59
rect 9472 50 9484 59
rect 9536 50 9644 59
rect 9696 50 9708 59
rect 9760 50 9868 59
rect 9920 50 9932 59
rect 9984 50 10092 59
rect 10144 50 10156 59
rect 10208 50 10316 59
rect 9088 16 9110 50
rect 9144 16 9182 50
rect 9248 16 9254 50
rect 9312 16 9326 50
rect 9360 16 9398 50
rect 9536 16 9542 50
rect 9576 16 9614 50
rect 9792 16 9830 50
rect 9864 16 9868 50
rect 10008 16 10046 50
rect 10080 16 10092 50
rect 10152 16 10156 50
rect 10224 16 10262 50
rect 10296 16 10316 50
rect 9088 7 9196 16
rect 9248 7 9260 16
rect 9312 7 9420 16
rect 9472 7 9484 16
rect 9536 7 9644 16
rect 9696 7 9708 16
rect 9760 7 9868 16
rect 9920 7 9932 16
rect 9984 7 10092 16
rect 10144 7 10156 16
rect 10208 7 10316 16
rect 10368 7 10380 59
rect 10432 50 10540 59
rect 10440 16 10478 50
rect 10512 16 10540 50
rect 10432 7 10540 16
rect 10592 7 10604 59
rect 10656 50 10764 59
rect 10656 16 10694 50
rect 10728 16 10764 50
rect 10656 7 10764 16
rect 10816 7 10828 59
rect 10880 50 10988 59
rect 10880 16 10910 50
rect 10944 16 10982 50
rect 10880 7 10988 16
rect 11040 7 11052 59
rect 11104 7 11146 59
rect 0 0 11146 7
<< via1 >>
rect 68 4594 120 4603
rect 132 4594 184 4603
rect 292 4594 344 4603
rect 356 4594 408 4603
rect 516 4594 568 4603
rect 580 4594 632 4603
rect 740 4594 792 4603
rect 68 4560 72 4594
rect 72 4560 110 4594
rect 110 4560 120 4594
rect 132 4560 144 4594
rect 144 4560 182 4594
rect 182 4560 184 4594
rect 292 4560 326 4594
rect 326 4560 344 4594
rect 356 4560 360 4594
rect 360 4560 398 4594
rect 398 4560 408 4594
rect 516 4560 542 4594
rect 542 4560 568 4594
rect 580 4560 614 4594
rect 614 4560 632 4594
rect 740 4560 758 4594
rect 758 4560 792 4594
rect 68 4551 120 4560
rect 132 4551 184 4560
rect 292 4551 344 4560
rect 356 4551 408 4560
rect 516 4551 568 4560
rect 580 4551 632 4560
rect 740 4551 792 4560
rect 804 4594 856 4603
rect 964 4594 1016 4603
rect 804 4560 830 4594
rect 830 4560 856 4594
rect 964 4560 974 4594
rect 974 4560 1008 4594
rect 1008 4560 1016 4594
rect 804 4551 856 4560
rect 964 4551 1016 4560
rect 1028 4594 1080 4603
rect 1188 4594 1240 4603
rect 1028 4560 1046 4594
rect 1046 4560 1080 4594
rect 1188 4560 1190 4594
rect 1190 4560 1224 4594
rect 1224 4560 1240 4594
rect 1028 4551 1080 4560
rect 1188 4551 1240 4560
rect 1252 4594 1304 4603
rect 1412 4594 1464 4603
rect 1252 4560 1262 4594
rect 1262 4560 1296 4594
rect 1296 4560 1304 4594
rect 1412 4560 1440 4594
rect 1440 4560 1464 4594
rect 1252 4551 1304 4560
rect 1412 4551 1464 4560
rect 1476 4594 1528 4603
rect 1636 4594 1688 4603
rect 1700 4594 1752 4603
rect 1860 4594 1912 4603
rect 1924 4594 1976 4603
rect 2084 4594 2136 4603
rect 2148 4594 2200 4603
rect 2308 4594 2360 4603
rect 2372 4594 2424 4603
rect 2532 4594 2584 4603
rect 2596 4594 2648 4603
rect 2756 4594 2808 4603
rect 1476 4560 1478 4594
rect 1478 4560 1512 4594
rect 1512 4560 1528 4594
rect 1636 4560 1656 4594
rect 1656 4560 1688 4594
rect 1700 4560 1728 4594
rect 1728 4560 1752 4594
rect 1860 4560 1872 4594
rect 1872 4560 1910 4594
rect 1910 4560 1912 4594
rect 1924 4560 1944 4594
rect 1944 4560 1976 4594
rect 2084 4560 2088 4594
rect 2088 4560 2126 4594
rect 2126 4560 2136 4594
rect 2148 4560 2160 4594
rect 2160 4560 2198 4594
rect 2198 4560 2200 4594
rect 2308 4560 2342 4594
rect 2342 4560 2360 4594
rect 2372 4560 2376 4594
rect 2376 4560 2414 4594
rect 2414 4560 2424 4594
rect 2532 4560 2558 4594
rect 2558 4560 2584 4594
rect 2596 4560 2630 4594
rect 2630 4560 2648 4594
rect 2756 4560 2774 4594
rect 2774 4560 2808 4594
rect 1476 4551 1528 4560
rect 1636 4551 1688 4560
rect 1700 4551 1752 4560
rect 1860 4551 1912 4560
rect 1924 4551 1976 4560
rect 2084 4551 2136 4560
rect 2148 4551 2200 4560
rect 2308 4551 2360 4560
rect 2372 4551 2424 4560
rect 2532 4551 2584 4560
rect 2596 4551 2648 4560
rect 2756 4551 2808 4560
rect 2820 4594 2872 4603
rect 2980 4594 3032 4603
rect 2820 4560 2846 4594
rect 2846 4560 2872 4594
rect 2980 4560 2990 4594
rect 2990 4560 3024 4594
rect 3024 4560 3032 4594
rect 2820 4551 2872 4560
rect 2980 4551 3032 4560
rect 3044 4594 3096 4603
rect 3204 4594 3256 4603
rect 3044 4560 3062 4594
rect 3062 4560 3096 4594
rect 3204 4560 3206 4594
rect 3206 4560 3240 4594
rect 3240 4560 3256 4594
rect 3044 4551 3096 4560
rect 3204 4551 3256 4560
rect 3268 4594 3320 4603
rect 3428 4594 3480 4603
rect 3268 4560 3278 4594
rect 3278 4560 3312 4594
rect 3312 4560 3320 4594
rect 3428 4560 3456 4594
rect 3456 4560 3480 4594
rect 3268 4551 3320 4560
rect 3428 4551 3480 4560
rect 3492 4594 3544 4603
rect 3652 4594 3704 4603
rect 3716 4594 3768 4603
rect 3876 4594 3928 4603
rect 3940 4594 3992 4603
rect 4100 4594 4152 4603
rect 4164 4594 4216 4603
rect 4324 4594 4376 4603
rect 4388 4594 4440 4603
rect 4548 4594 4600 4603
rect 4612 4594 4664 4603
rect 4772 4594 4824 4603
rect 3492 4560 3494 4594
rect 3494 4560 3528 4594
rect 3528 4560 3544 4594
rect 3652 4560 3672 4594
rect 3672 4560 3704 4594
rect 3716 4560 3744 4594
rect 3744 4560 3768 4594
rect 3876 4560 3888 4594
rect 3888 4560 3926 4594
rect 3926 4560 3928 4594
rect 3940 4560 3960 4594
rect 3960 4560 3992 4594
rect 4100 4560 4104 4594
rect 4104 4560 4142 4594
rect 4142 4560 4152 4594
rect 4164 4560 4176 4594
rect 4176 4560 4214 4594
rect 4214 4560 4216 4594
rect 4324 4560 4358 4594
rect 4358 4560 4376 4594
rect 4388 4560 4392 4594
rect 4392 4560 4430 4594
rect 4430 4560 4440 4594
rect 4548 4560 4574 4594
rect 4574 4560 4600 4594
rect 4612 4560 4646 4594
rect 4646 4560 4664 4594
rect 4772 4560 4790 4594
rect 4790 4560 4824 4594
rect 3492 4551 3544 4560
rect 3652 4551 3704 4560
rect 3716 4551 3768 4560
rect 3876 4551 3928 4560
rect 3940 4551 3992 4560
rect 4100 4551 4152 4560
rect 4164 4551 4216 4560
rect 4324 4551 4376 4560
rect 4388 4551 4440 4560
rect 4548 4551 4600 4560
rect 4612 4551 4664 4560
rect 4772 4551 4824 4560
rect 4836 4594 4888 4603
rect 4996 4594 5048 4603
rect 4836 4560 4862 4594
rect 4862 4560 4888 4594
rect 4996 4560 5006 4594
rect 5006 4560 5040 4594
rect 5040 4560 5048 4594
rect 4836 4551 4888 4560
rect 4996 4551 5048 4560
rect 5060 4594 5112 4603
rect 5220 4594 5272 4603
rect 5060 4560 5078 4594
rect 5078 4560 5112 4594
rect 5220 4560 5222 4594
rect 5222 4560 5256 4594
rect 5256 4560 5272 4594
rect 5060 4551 5112 4560
rect 5220 4551 5272 4560
rect 5284 4594 5336 4603
rect 5444 4594 5496 4603
rect 5284 4560 5294 4594
rect 5294 4560 5328 4594
rect 5328 4560 5336 4594
rect 5444 4560 5472 4594
rect 5472 4560 5496 4594
rect 5284 4551 5336 4560
rect 5444 4551 5496 4560
rect 5508 4594 5560 4603
rect 5668 4594 5720 4603
rect 5732 4594 5784 4603
rect 5892 4594 5944 4603
rect 5956 4594 6008 4603
rect 6116 4594 6168 4603
rect 6180 4594 6232 4603
rect 6340 4594 6392 4603
rect 6404 4594 6456 4603
rect 6564 4594 6616 4603
rect 6628 4594 6680 4603
rect 6788 4594 6840 4603
rect 5508 4560 5510 4594
rect 5510 4560 5544 4594
rect 5544 4560 5560 4594
rect 5668 4560 5688 4594
rect 5688 4560 5720 4594
rect 5732 4560 5760 4594
rect 5760 4560 5784 4594
rect 5892 4560 5904 4594
rect 5904 4560 5942 4594
rect 5942 4560 5944 4594
rect 5956 4560 5976 4594
rect 5976 4560 6008 4594
rect 6116 4560 6120 4594
rect 6120 4560 6158 4594
rect 6158 4560 6168 4594
rect 6180 4560 6192 4594
rect 6192 4560 6230 4594
rect 6230 4560 6232 4594
rect 6340 4560 6374 4594
rect 6374 4560 6392 4594
rect 6404 4560 6408 4594
rect 6408 4560 6446 4594
rect 6446 4560 6456 4594
rect 6564 4560 6590 4594
rect 6590 4560 6616 4594
rect 6628 4560 6662 4594
rect 6662 4560 6680 4594
rect 6788 4560 6806 4594
rect 6806 4560 6840 4594
rect 5508 4551 5560 4560
rect 5668 4551 5720 4560
rect 5732 4551 5784 4560
rect 5892 4551 5944 4560
rect 5956 4551 6008 4560
rect 6116 4551 6168 4560
rect 6180 4551 6232 4560
rect 6340 4551 6392 4560
rect 6404 4551 6456 4560
rect 6564 4551 6616 4560
rect 6628 4551 6680 4560
rect 6788 4551 6840 4560
rect 6852 4594 6904 4603
rect 7012 4594 7064 4603
rect 6852 4560 6878 4594
rect 6878 4560 6904 4594
rect 7012 4560 7022 4594
rect 7022 4560 7056 4594
rect 7056 4560 7064 4594
rect 6852 4551 6904 4560
rect 7012 4551 7064 4560
rect 7076 4594 7128 4603
rect 7236 4594 7288 4603
rect 7076 4560 7094 4594
rect 7094 4560 7128 4594
rect 7236 4560 7238 4594
rect 7238 4560 7272 4594
rect 7272 4560 7288 4594
rect 7076 4551 7128 4560
rect 7236 4551 7288 4560
rect 7300 4594 7352 4603
rect 7460 4594 7512 4603
rect 7300 4560 7310 4594
rect 7310 4560 7344 4594
rect 7344 4560 7352 4594
rect 7460 4560 7488 4594
rect 7488 4560 7512 4594
rect 7300 4551 7352 4560
rect 7460 4551 7512 4560
rect 7524 4594 7576 4603
rect 7684 4594 7736 4603
rect 7748 4594 7800 4603
rect 7908 4594 7960 4603
rect 7972 4594 8024 4603
rect 8132 4594 8184 4603
rect 8196 4594 8248 4603
rect 8356 4594 8408 4603
rect 8420 4594 8472 4603
rect 8580 4594 8632 4603
rect 8644 4594 8696 4603
rect 8804 4594 8856 4603
rect 7524 4560 7526 4594
rect 7526 4560 7560 4594
rect 7560 4560 7576 4594
rect 7684 4560 7704 4594
rect 7704 4560 7736 4594
rect 7748 4560 7776 4594
rect 7776 4560 7800 4594
rect 7908 4560 7920 4594
rect 7920 4560 7958 4594
rect 7958 4560 7960 4594
rect 7972 4560 7992 4594
rect 7992 4560 8024 4594
rect 8132 4560 8136 4594
rect 8136 4560 8174 4594
rect 8174 4560 8184 4594
rect 8196 4560 8208 4594
rect 8208 4560 8246 4594
rect 8246 4560 8248 4594
rect 8356 4560 8390 4594
rect 8390 4560 8408 4594
rect 8420 4560 8424 4594
rect 8424 4560 8462 4594
rect 8462 4560 8472 4594
rect 8580 4560 8606 4594
rect 8606 4560 8632 4594
rect 8644 4560 8678 4594
rect 8678 4560 8696 4594
rect 8804 4560 8822 4594
rect 8822 4560 8856 4594
rect 7524 4551 7576 4560
rect 7684 4551 7736 4560
rect 7748 4551 7800 4560
rect 7908 4551 7960 4560
rect 7972 4551 8024 4560
rect 8132 4551 8184 4560
rect 8196 4551 8248 4560
rect 8356 4551 8408 4560
rect 8420 4551 8472 4560
rect 8580 4551 8632 4560
rect 8644 4551 8696 4560
rect 8804 4551 8856 4560
rect 8868 4594 8920 4603
rect 9028 4594 9080 4603
rect 8868 4560 8894 4594
rect 8894 4560 8920 4594
rect 9028 4560 9038 4594
rect 9038 4560 9072 4594
rect 9072 4560 9080 4594
rect 8868 4551 8920 4560
rect 9028 4551 9080 4560
rect 9092 4594 9144 4603
rect 9252 4594 9304 4603
rect 9092 4560 9110 4594
rect 9110 4560 9144 4594
rect 9252 4560 9254 4594
rect 9254 4560 9288 4594
rect 9288 4560 9304 4594
rect 9092 4551 9144 4560
rect 9252 4551 9304 4560
rect 9316 4594 9368 4603
rect 9476 4594 9528 4603
rect 9316 4560 9326 4594
rect 9326 4560 9360 4594
rect 9360 4560 9368 4594
rect 9476 4560 9504 4594
rect 9504 4560 9528 4594
rect 9316 4551 9368 4560
rect 9476 4551 9528 4560
rect 9540 4594 9592 4603
rect 9700 4594 9752 4603
rect 9764 4594 9816 4603
rect 9924 4594 9976 4603
rect 9988 4594 10040 4603
rect 10148 4594 10200 4603
rect 10212 4594 10264 4603
rect 10372 4594 10424 4603
rect 10436 4594 10488 4603
rect 10596 4594 10648 4603
rect 10660 4594 10712 4603
rect 10820 4594 10872 4603
rect 9540 4560 9542 4594
rect 9542 4560 9576 4594
rect 9576 4560 9592 4594
rect 9700 4560 9720 4594
rect 9720 4560 9752 4594
rect 9764 4560 9792 4594
rect 9792 4560 9816 4594
rect 9924 4560 9936 4594
rect 9936 4560 9974 4594
rect 9974 4560 9976 4594
rect 9988 4560 10008 4594
rect 10008 4560 10040 4594
rect 10148 4560 10152 4594
rect 10152 4560 10190 4594
rect 10190 4560 10200 4594
rect 10212 4560 10224 4594
rect 10224 4560 10262 4594
rect 10262 4560 10264 4594
rect 10372 4560 10406 4594
rect 10406 4560 10424 4594
rect 10436 4560 10440 4594
rect 10440 4560 10478 4594
rect 10478 4560 10488 4594
rect 10596 4560 10622 4594
rect 10622 4560 10648 4594
rect 10660 4560 10694 4594
rect 10694 4560 10712 4594
rect 10820 4560 10838 4594
rect 10838 4560 10872 4594
rect 9540 4551 9592 4560
rect 9700 4551 9752 4560
rect 9764 4551 9816 4560
rect 9924 4551 9976 4560
rect 9988 4551 10040 4560
rect 10148 4551 10200 4560
rect 10212 4551 10264 4560
rect 10372 4551 10424 4560
rect 10436 4551 10488 4560
rect 10596 4551 10648 4560
rect 10660 4551 10712 4560
rect 10820 4551 10872 4560
rect 10884 4594 10936 4603
rect 10884 4560 10910 4594
rect 10910 4560 10936 4594
rect 10884 4551 10936 4560
rect 24 50 76 59
rect 24 16 38 50
rect 38 16 72 50
rect 72 16 76 50
rect 24 7 76 16
rect 88 50 140 59
rect 236 50 288 59
rect 88 16 110 50
rect 110 16 140 50
rect 236 16 254 50
rect 254 16 288 50
rect 88 7 140 16
rect 236 7 288 16
rect 300 50 352 59
rect 460 50 512 59
rect 300 16 326 50
rect 326 16 352 50
rect 460 16 470 50
rect 470 16 504 50
rect 504 16 512 50
rect 300 7 352 16
rect 460 7 512 16
rect 524 50 576 59
rect 684 50 736 59
rect 524 16 542 50
rect 542 16 576 50
rect 684 16 686 50
rect 686 16 720 50
rect 720 16 736 50
rect 524 7 576 16
rect 684 7 736 16
rect 748 50 800 59
rect 908 50 960 59
rect 748 16 758 50
rect 758 16 792 50
rect 792 16 800 50
rect 908 16 936 50
rect 936 16 960 50
rect 748 7 800 16
rect 908 7 960 16
rect 972 50 1024 59
rect 1132 50 1184 59
rect 1196 50 1248 59
rect 1356 50 1408 59
rect 1420 50 1472 59
rect 1580 50 1632 59
rect 1644 50 1696 59
rect 1804 50 1856 59
rect 1868 50 1920 59
rect 2028 50 2080 59
rect 2092 50 2144 59
rect 2252 50 2304 59
rect 972 16 974 50
rect 974 16 1008 50
rect 1008 16 1024 50
rect 1132 16 1152 50
rect 1152 16 1184 50
rect 1196 16 1224 50
rect 1224 16 1248 50
rect 1356 16 1368 50
rect 1368 16 1406 50
rect 1406 16 1408 50
rect 1420 16 1440 50
rect 1440 16 1472 50
rect 1580 16 1584 50
rect 1584 16 1622 50
rect 1622 16 1632 50
rect 1644 16 1656 50
rect 1656 16 1694 50
rect 1694 16 1696 50
rect 1804 16 1838 50
rect 1838 16 1856 50
rect 1868 16 1872 50
rect 1872 16 1910 50
rect 1910 16 1920 50
rect 2028 16 2054 50
rect 2054 16 2080 50
rect 2092 16 2126 50
rect 2126 16 2144 50
rect 2252 16 2270 50
rect 2270 16 2304 50
rect 972 7 1024 16
rect 1132 7 1184 16
rect 1196 7 1248 16
rect 1356 7 1408 16
rect 1420 7 1472 16
rect 1580 7 1632 16
rect 1644 7 1696 16
rect 1804 7 1856 16
rect 1868 7 1920 16
rect 2028 7 2080 16
rect 2092 7 2144 16
rect 2252 7 2304 16
rect 2316 50 2368 59
rect 2476 50 2528 59
rect 2316 16 2342 50
rect 2342 16 2368 50
rect 2476 16 2486 50
rect 2486 16 2520 50
rect 2520 16 2528 50
rect 2316 7 2368 16
rect 2476 7 2528 16
rect 2540 50 2592 59
rect 2700 50 2752 59
rect 2540 16 2558 50
rect 2558 16 2592 50
rect 2700 16 2702 50
rect 2702 16 2736 50
rect 2736 16 2752 50
rect 2540 7 2592 16
rect 2700 7 2752 16
rect 2764 50 2816 59
rect 2924 50 2976 59
rect 2764 16 2774 50
rect 2774 16 2808 50
rect 2808 16 2816 50
rect 2924 16 2952 50
rect 2952 16 2976 50
rect 2764 7 2816 16
rect 2924 7 2976 16
rect 2988 50 3040 59
rect 3148 50 3200 59
rect 3212 50 3264 59
rect 3372 50 3424 59
rect 3436 50 3488 59
rect 3596 50 3648 59
rect 3660 50 3712 59
rect 3820 50 3872 59
rect 3884 50 3936 59
rect 4044 50 4096 59
rect 4108 50 4160 59
rect 4268 50 4320 59
rect 2988 16 2990 50
rect 2990 16 3024 50
rect 3024 16 3040 50
rect 3148 16 3168 50
rect 3168 16 3200 50
rect 3212 16 3240 50
rect 3240 16 3264 50
rect 3372 16 3384 50
rect 3384 16 3422 50
rect 3422 16 3424 50
rect 3436 16 3456 50
rect 3456 16 3488 50
rect 3596 16 3600 50
rect 3600 16 3638 50
rect 3638 16 3648 50
rect 3660 16 3672 50
rect 3672 16 3710 50
rect 3710 16 3712 50
rect 3820 16 3854 50
rect 3854 16 3872 50
rect 3884 16 3888 50
rect 3888 16 3926 50
rect 3926 16 3936 50
rect 4044 16 4070 50
rect 4070 16 4096 50
rect 4108 16 4142 50
rect 4142 16 4160 50
rect 4268 16 4286 50
rect 4286 16 4320 50
rect 2988 7 3040 16
rect 3148 7 3200 16
rect 3212 7 3264 16
rect 3372 7 3424 16
rect 3436 7 3488 16
rect 3596 7 3648 16
rect 3660 7 3712 16
rect 3820 7 3872 16
rect 3884 7 3936 16
rect 4044 7 4096 16
rect 4108 7 4160 16
rect 4268 7 4320 16
rect 4332 50 4384 59
rect 4492 50 4544 59
rect 4332 16 4358 50
rect 4358 16 4384 50
rect 4492 16 4502 50
rect 4502 16 4536 50
rect 4536 16 4544 50
rect 4332 7 4384 16
rect 4492 7 4544 16
rect 4556 50 4608 59
rect 4716 50 4768 59
rect 4556 16 4574 50
rect 4574 16 4608 50
rect 4716 16 4718 50
rect 4718 16 4752 50
rect 4752 16 4768 50
rect 4556 7 4608 16
rect 4716 7 4768 16
rect 4780 50 4832 59
rect 4940 50 4992 59
rect 4780 16 4790 50
rect 4790 16 4824 50
rect 4824 16 4832 50
rect 4940 16 4968 50
rect 4968 16 4992 50
rect 4780 7 4832 16
rect 4940 7 4992 16
rect 5004 50 5056 59
rect 5164 50 5216 59
rect 5228 50 5280 59
rect 5388 50 5440 59
rect 5452 50 5504 59
rect 5612 50 5664 59
rect 5676 50 5728 59
rect 5836 50 5888 59
rect 5900 50 5952 59
rect 6060 50 6112 59
rect 6124 50 6176 59
rect 6284 50 6336 59
rect 5004 16 5006 50
rect 5006 16 5040 50
rect 5040 16 5056 50
rect 5164 16 5184 50
rect 5184 16 5216 50
rect 5228 16 5256 50
rect 5256 16 5280 50
rect 5388 16 5400 50
rect 5400 16 5438 50
rect 5438 16 5440 50
rect 5452 16 5472 50
rect 5472 16 5504 50
rect 5612 16 5616 50
rect 5616 16 5654 50
rect 5654 16 5664 50
rect 5676 16 5688 50
rect 5688 16 5726 50
rect 5726 16 5728 50
rect 5836 16 5870 50
rect 5870 16 5888 50
rect 5900 16 5904 50
rect 5904 16 5942 50
rect 5942 16 5952 50
rect 6060 16 6086 50
rect 6086 16 6112 50
rect 6124 16 6158 50
rect 6158 16 6176 50
rect 6284 16 6302 50
rect 6302 16 6336 50
rect 5004 7 5056 16
rect 5164 7 5216 16
rect 5228 7 5280 16
rect 5388 7 5440 16
rect 5452 7 5504 16
rect 5612 7 5664 16
rect 5676 7 5728 16
rect 5836 7 5888 16
rect 5900 7 5952 16
rect 6060 7 6112 16
rect 6124 7 6176 16
rect 6284 7 6336 16
rect 6348 50 6400 59
rect 6508 50 6560 59
rect 6348 16 6374 50
rect 6374 16 6400 50
rect 6508 16 6518 50
rect 6518 16 6552 50
rect 6552 16 6560 50
rect 6348 7 6400 16
rect 6508 7 6560 16
rect 6572 50 6624 59
rect 6732 50 6784 59
rect 6572 16 6590 50
rect 6590 16 6624 50
rect 6732 16 6734 50
rect 6734 16 6768 50
rect 6768 16 6784 50
rect 6572 7 6624 16
rect 6732 7 6784 16
rect 6796 50 6848 59
rect 6956 50 7008 59
rect 6796 16 6806 50
rect 6806 16 6840 50
rect 6840 16 6848 50
rect 6956 16 6984 50
rect 6984 16 7008 50
rect 6796 7 6848 16
rect 6956 7 7008 16
rect 7020 50 7072 59
rect 7180 50 7232 59
rect 7244 50 7296 59
rect 7404 50 7456 59
rect 7468 50 7520 59
rect 7628 50 7680 59
rect 7692 50 7744 59
rect 7852 50 7904 59
rect 7916 50 7968 59
rect 8076 50 8128 59
rect 8140 50 8192 59
rect 8300 50 8352 59
rect 7020 16 7022 50
rect 7022 16 7056 50
rect 7056 16 7072 50
rect 7180 16 7200 50
rect 7200 16 7232 50
rect 7244 16 7272 50
rect 7272 16 7296 50
rect 7404 16 7416 50
rect 7416 16 7454 50
rect 7454 16 7456 50
rect 7468 16 7488 50
rect 7488 16 7520 50
rect 7628 16 7632 50
rect 7632 16 7670 50
rect 7670 16 7680 50
rect 7692 16 7704 50
rect 7704 16 7742 50
rect 7742 16 7744 50
rect 7852 16 7886 50
rect 7886 16 7904 50
rect 7916 16 7920 50
rect 7920 16 7958 50
rect 7958 16 7968 50
rect 8076 16 8102 50
rect 8102 16 8128 50
rect 8140 16 8174 50
rect 8174 16 8192 50
rect 8300 16 8318 50
rect 8318 16 8352 50
rect 7020 7 7072 16
rect 7180 7 7232 16
rect 7244 7 7296 16
rect 7404 7 7456 16
rect 7468 7 7520 16
rect 7628 7 7680 16
rect 7692 7 7744 16
rect 7852 7 7904 16
rect 7916 7 7968 16
rect 8076 7 8128 16
rect 8140 7 8192 16
rect 8300 7 8352 16
rect 8364 50 8416 59
rect 8524 50 8576 59
rect 8364 16 8390 50
rect 8390 16 8416 50
rect 8524 16 8534 50
rect 8534 16 8568 50
rect 8568 16 8576 50
rect 8364 7 8416 16
rect 8524 7 8576 16
rect 8588 50 8640 59
rect 8748 50 8800 59
rect 8588 16 8606 50
rect 8606 16 8640 50
rect 8748 16 8750 50
rect 8750 16 8784 50
rect 8784 16 8800 50
rect 8588 7 8640 16
rect 8748 7 8800 16
rect 8812 50 8864 59
rect 8972 50 9024 59
rect 8812 16 8822 50
rect 8822 16 8856 50
rect 8856 16 8864 50
rect 8972 16 9000 50
rect 9000 16 9024 50
rect 8812 7 8864 16
rect 8972 7 9024 16
rect 9036 50 9088 59
rect 9196 50 9248 59
rect 9260 50 9312 59
rect 9420 50 9472 59
rect 9484 50 9536 59
rect 9644 50 9696 59
rect 9708 50 9760 59
rect 9868 50 9920 59
rect 9932 50 9984 59
rect 10092 50 10144 59
rect 10156 50 10208 59
rect 10316 50 10368 59
rect 9036 16 9038 50
rect 9038 16 9072 50
rect 9072 16 9088 50
rect 9196 16 9216 50
rect 9216 16 9248 50
rect 9260 16 9288 50
rect 9288 16 9312 50
rect 9420 16 9432 50
rect 9432 16 9470 50
rect 9470 16 9472 50
rect 9484 16 9504 50
rect 9504 16 9536 50
rect 9644 16 9648 50
rect 9648 16 9686 50
rect 9686 16 9696 50
rect 9708 16 9720 50
rect 9720 16 9758 50
rect 9758 16 9760 50
rect 9868 16 9902 50
rect 9902 16 9920 50
rect 9932 16 9936 50
rect 9936 16 9974 50
rect 9974 16 9984 50
rect 10092 16 10118 50
rect 10118 16 10144 50
rect 10156 16 10190 50
rect 10190 16 10208 50
rect 10316 16 10334 50
rect 10334 16 10368 50
rect 9036 7 9088 16
rect 9196 7 9248 16
rect 9260 7 9312 16
rect 9420 7 9472 16
rect 9484 7 9536 16
rect 9644 7 9696 16
rect 9708 7 9760 16
rect 9868 7 9920 16
rect 9932 7 9984 16
rect 10092 7 10144 16
rect 10156 7 10208 16
rect 10316 7 10368 16
rect 10380 50 10432 59
rect 10540 50 10592 59
rect 10380 16 10406 50
rect 10406 16 10432 50
rect 10540 16 10550 50
rect 10550 16 10584 50
rect 10584 16 10592 50
rect 10380 7 10432 16
rect 10540 7 10592 16
rect 10604 50 10656 59
rect 10764 50 10816 59
rect 10604 16 10622 50
rect 10622 16 10656 50
rect 10764 16 10766 50
rect 10766 16 10800 50
rect 10800 16 10816 50
rect 10604 7 10656 16
rect 10764 7 10816 16
rect 10828 50 10880 59
rect 10988 50 11040 59
rect 10828 16 10838 50
rect 10838 16 10872 50
rect 10872 16 10880 50
rect 10988 16 11016 50
rect 11016 16 11040 50
rect 10828 7 10880 16
rect 10988 7 11040 16
rect 11052 50 11104 59
rect 11052 16 11054 50
rect 11054 16 11088 50
rect 11088 16 11104 50
rect 11052 7 11104 16
<< metal2 >>
rect 0 66 28 4610
rect 56 4605 196 4610
rect 56 4603 98 4605
rect 154 4603 196 4605
rect 56 4551 68 4603
rect 184 4551 196 4603
rect 56 4549 98 4551
rect 154 4549 196 4551
rect 56 4544 196 4549
rect 56 94 84 4544
rect 112 66 140 4516
rect 0 61 140 66
rect 0 59 42 61
rect 98 59 140 61
rect 0 7 24 59
rect 0 5 42 7
rect 98 5 140 7
rect 0 0 140 5
rect 168 0 196 4544
rect 224 66 252 4610
rect 280 4605 420 4610
rect 280 4603 322 4605
rect 378 4603 420 4605
rect 280 4551 292 4603
rect 408 4551 420 4603
rect 280 4549 322 4551
rect 378 4549 420 4551
rect 280 4544 420 4549
rect 280 94 308 4544
rect 336 66 364 4516
rect 224 61 364 66
rect 224 59 266 61
rect 322 59 364 61
rect 224 7 236 59
rect 352 7 364 59
rect 224 5 266 7
rect 322 5 364 7
rect 224 0 364 5
rect 392 0 420 4544
rect 448 66 476 4610
rect 504 4605 644 4610
rect 504 4603 546 4605
rect 602 4603 644 4605
rect 504 4551 516 4603
rect 632 4551 644 4603
rect 504 4549 546 4551
rect 602 4549 644 4551
rect 504 4544 644 4549
rect 504 94 532 4544
rect 560 66 588 4516
rect 448 61 588 66
rect 448 59 490 61
rect 546 59 588 61
rect 448 7 460 59
rect 576 7 588 59
rect 448 5 490 7
rect 546 5 588 7
rect 448 0 588 5
rect 616 0 644 4544
rect 672 66 700 4610
rect 728 4605 868 4610
rect 728 4603 770 4605
rect 826 4603 868 4605
rect 728 4551 740 4603
rect 856 4551 868 4603
rect 728 4549 770 4551
rect 826 4549 868 4551
rect 728 4544 868 4549
rect 728 94 756 4544
rect 784 66 812 4516
rect 672 61 812 66
rect 672 59 714 61
rect 770 59 812 61
rect 672 7 684 59
rect 800 7 812 59
rect 672 5 714 7
rect 770 5 812 7
rect 672 0 812 5
rect 840 0 868 4544
rect 896 66 924 4610
rect 952 4605 1092 4610
rect 952 4603 994 4605
rect 1050 4603 1092 4605
rect 952 4551 964 4603
rect 1080 4551 1092 4603
rect 952 4549 994 4551
rect 1050 4549 1092 4551
rect 952 4544 1092 4549
rect 952 94 980 4544
rect 1008 66 1036 4516
rect 896 61 1036 66
rect 896 59 938 61
rect 994 59 1036 61
rect 896 7 908 59
rect 1024 7 1036 59
rect 896 5 938 7
rect 994 5 1036 7
rect 896 0 1036 5
rect 1064 0 1092 4544
rect 1120 66 1148 4610
rect 1176 4605 1316 4610
rect 1176 4603 1218 4605
rect 1274 4603 1316 4605
rect 1176 4551 1188 4603
rect 1304 4551 1316 4603
rect 1176 4549 1218 4551
rect 1274 4549 1316 4551
rect 1176 4544 1316 4549
rect 1176 94 1204 4544
rect 1232 66 1260 4516
rect 1120 61 1260 66
rect 1120 59 1162 61
rect 1218 59 1260 61
rect 1120 7 1132 59
rect 1248 7 1260 59
rect 1120 5 1162 7
rect 1218 5 1260 7
rect 1120 0 1260 5
rect 1288 0 1316 4544
rect 1344 66 1372 4610
rect 1400 4605 1540 4610
rect 1400 4603 1442 4605
rect 1498 4603 1540 4605
rect 1400 4551 1412 4603
rect 1528 4551 1540 4603
rect 1400 4549 1442 4551
rect 1498 4549 1540 4551
rect 1400 4544 1540 4549
rect 1400 94 1428 4544
rect 1456 66 1484 4516
rect 1344 61 1484 66
rect 1344 59 1386 61
rect 1442 59 1484 61
rect 1344 7 1356 59
rect 1472 7 1484 59
rect 1344 5 1386 7
rect 1442 5 1484 7
rect 1344 0 1484 5
rect 1512 0 1540 4544
rect 1568 66 1596 4610
rect 1624 4605 1764 4610
rect 1624 4603 1666 4605
rect 1722 4603 1764 4605
rect 1624 4551 1636 4603
rect 1752 4551 1764 4603
rect 1624 4549 1666 4551
rect 1722 4549 1764 4551
rect 1624 4544 1764 4549
rect 1624 94 1652 4544
rect 1680 66 1708 4516
rect 1568 61 1708 66
rect 1568 59 1610 61
rect 1666 59 1708 61
rect 1568 7 1580 59
rect 1696 7 1708 59
rect 1568 5 1610 7
rect 1666 5 1708 7
rect 1568 0 1708 5
rect 1736 0 1764 4544
rect 1792 66 1820 4610
rect 1848 4605 1988 4610
rect 1848 4603 1890 4605
rect 1946 4603 1988 4605
rect 1848 4551 1860 4603
rect 1976 4551 1988 4603
rect 1848 4549 1890 4551
rect 1946 4549 1988 4551
rect 1848 4544 1988 4549
rect 1848 94 1876 4544
rect 1904 66 1932 4516
rect 1792 61 1932 66
rect 1792 59 1834 61
rect 1890 59 1932 61
rect 1792 7 1804 59
rect 1920 7 1932 59
rect 1792 5 1834 7
rect 1890 5 1932 7
rect 1792 0 1932 5
rect 1960 0 1988 4544
rect 2016 66 2044 4610
rect 2072 4605 2212 4610
rect 2072 4603 2114 4605
rect 2170 4603 2212 4605
rect 2072 4551 2084 4603
rect 2200 4551 2212 4603
rect 2072 4549 2114 4551
rect 2170 4549 2212 4551
rect 2072 4544 2212 4549
rect 2072 94 2100 4544
rect 2128 66 2156 4516
rect 2016 61 2156 66
rect 2016 59 2058 61
rect 2114 59 2156 61
rect 2016 7 2028 59
rect 2144 7 2156 59
rect 2016 5 2058 7
rect 2114 5 2156 7
rect 2016 0 2156 5
rect 2184 0 2212 4544
rect 2240 66 2268 4610
rect 2296 4605 2436 4610
rect 2296 4603 2338 4605
rect 2394 4603 2436 4605
rect 2296 4551 2308 4603
rect 2424 4551 2436 4603
rect 2296 4549 2338 4551
rect 2394 4549 2436 4551
rect 2296 4544 2436 4549
rect 2296 94 2324 4544
rect 2352 66 2380 4516
rect 2240 61 2380 66
rect 2240 59 2282 61
rect 2338 59 2380 61
rect 2240 7 2252 59
rect 2368 7 2380 59
rect 2240 5 2282 7
rect 2338 5 2380 7
rect 2240 0 2380 5
rect 2408 0 2436 4544
rect 2464 66 2492 4610
rect 2520 4605 2660 4610
rect 2520 4603 2562 4605
rect 2618 4603 2660 4605
rect 2520 4551 2532 4603
rect 2648 4551 2660 4603
rect 2520 4549 2562 4551
rect 2618 4549 2660 4551
rect 2520 4544 2660 4549
rect 2520 94 2548 4544
rect 2576 66 2604 4516
rect 2464 61 2604 66
rect 2464 59 2506 61
rect 2562 59 2604 61
rect 2464 7 2476 59
rect 2592 7 2604 59
rect 2464 5 2506 7
rect 2562 5 2604 7
rect 2464 0 2604 5
rect 2632 0 2660 4544
rect 2688 66 2716 4610
rect 2744 4605 2884 4610
rect 2744 4603 2786 4605
rect 2842 4603 2884 4605
rect 2744 4551 2756 4603
rect 2872 4551 2884 4603
rect 2744 4549 2786 4551
rect 2842 4549 2884 4551
rect 2744 4544 2884 4549
rect 2744 94 2772 4544
rect 2800 66 2828 4516
rect 2688 61 2828 66
rect 2688 59 2730 61
rect 2786 59 2828 61
rect 2688 7 2700 59
rect 2816 7 2828 59
rect 2688 5 2730 7
rect 2786 5 2828 7
rect 2688 0 2828 5
rect 2856 0 2884 4544
rect 2912 66 2940 4610
rect 2968 4605 3108 4610
rect 2968 4603 3010 4605
rect 3066 4603 3108 4605
rect 2968 4551 2980 4603
rect 3096 4551 3108 4603
rect 2968 4549 3010 4551
rect 3066 4549 3108 4551
rect 2968 4544 3108 4549
rect 2968 94 2996 4544
rect 3024 66 3052 4516
rect 2912 61 3052 66
rect 2912 59 2954 61
rect 3010 59 3052 61
rect 2912 7 2924 59
rect 3040 7 3052 59
rect 2912 5 2954 7
rect 3010 5 3052 7
rect 2912 0 3052 5
rect 3080 0 3108 4544
rect 3136 66 3164 4610
rect 3192 4605 3332 4610
rect 3192 4603 3234 4605
rect 3290 4603 3332 4605
rect 3192 4551 3204 4603
rect 3320 4551 3332 4603
rect 3192 4549 3234 4551
rect 3290 4549 3332 4551
rect 3192 4544 3332 4549
rect 3192 94 3220 4544
rect 3248 66 3276 4516
rect 3136 61 3276 66
rect 3136 59 3178 61
rect 3234 59 3276 61
rect 3136 7 3148 59
rect 3264 7 3276 59
rect 3136 5 3178 7
rect 3234 5 3276 7
rect 3136 0 3276 5
rect 3304 0 3332 4544
rect 3360 66 3388 4610
rect 3416 4605 3556 4610
rect 3416 4603 3458 4605
rect 3514 4603 3556 4605
rect 3416 4551 3428 4603
rect 3544 4551 3556 4603
rect 3416 4549 3458 4551
rect 3514 4549 3556 4551
rect 3416 4544 3556 4549
rect 3416 94 3444 4544
rect 3472 66 3500 4516
rect 3360 61 3500 66
rect 3360 59 3402 61
rect 3458 59 3500 61
rect 3360 7 3372 59
rect 3488 7 3500 59
rect 3360 5 3402 7
rect 3458 5 3500 7
rect 3360 0 3500 5
rect 3528 0 3556 4544
rect 3584 66 3612 4610
rect 3640 4605 3780 4610
rect 3640 4603 3682 4605
rect 3738 4603 3780 4605
rect 3640 4551 3652 4603
rect 3768 4551 3780 4603
rect 3640 4549 3682 4551
rect 3738 4549 3780 4551
rect 3640 4544 3780 4549
rect 3640 94 3668 4544
rect 3696 66 3724 4516
rect 3584 61 3724 66
rect 3584 59 3626 61
rect 3682 59 3724 61
rect 3584 7 3596 59
rect 3712 7 3724 59
rect 3584 5 3626 7
rect 3682 5 3724 7
rect 3584 0 3724 5
rect 3752 0 3780 4544
rect 3808 66 3836 4610
rect 3864 4605 4004 4610
rect 3864 4603 3906 4605
rect 3962 4603 4004 4605
rect 3864 4551 3876 4603
rect 3992 4551 4004 4603
rect 3864 4549 3906 4551
rect 3962 4549 4004 4551
rect 3864 4544 4004 4549
rect 3864 94 3892 4544
rect 3920 66 3948 4516
rect 3808 61 3948 66
rect 3808 59 3850 61
rect 3906 59 3948 61
rect 3808 7 3820 59
rect 3936 7 3948 59
rect 3808 5 3850 7
rect 3906 5 3948 7
rect 3808 0 3948 5
rect 3976 0 4004 4544
rect 4032 66 4060 4610
rect 4088 4605 4228 4610
rect 4088 4603 4130 4605
rect 4186 4603 4228 4605
rect 4088 4551 4100 4603
rect 4216 4551 4228 4603
rect 4088 4549 4130 4551
rect 4186 4549 4228 4551
rect 4088 4544 4228 4549
rect 4088 94 4116 4544
rect 4144 66 4172 4516
rect 4032 61 4172 66
rect 4032 59 4074 61
rect 4130 59 4172 61
rect 4032 7 4044 59
rect 4160 7 4172 59
rect 4032 5 4074 7
rect 4130 5 4172 7
rect 4032 0 4172 5
rect 4200 0 4228 4544
rect 4256 66 4284 4610
rect 4312 4605 4452 4610
rect 4312 4603 4354 4605
rect 4410 4603 4452 4605
rect 4312 4551 4324 4603
rect 4440 4551 4452 4603
rect 4312 4549 4354 4551
rect 4410 4549 4452 4551
rect 4312 4544 4452 4549
rect 4312 94 4340 4544
rect 4368 66 4396 4516
rect 4256 61 4396 66
rect 4256 59 4298 61
rect 4354 59 4396 61
rect 4256 7 4268 59
rect 4384 7 4396 59
rect 4256 5 4298 7
rect 4354 5 4396 7
rect 4256 0 4396 5
rect 4424 0 4452 4544
rect 4480 66 4508 4610
rect 4536 4605 4676 4610
rect 4536 4603 4578 4605
rect 4634 4603 4676 4605
rect 4536 4551 4548 4603
rect 4664 4551 4676 4603
rect 4536 4549 4578 4551
rect 4634 4549 4676 4551
rect 4536 4544 4676 4549
rect 4536 94 4564 4544
rect 4592 66 4620 4516
rect 4480 61 4620 66
rect 4480 59 4522 61
rect 4578 59 4620 61
rect 4480 7 4492 59
rect 4608 7 4620 59
rect 4480 5 4522 7
rect 4578 5 4620 7
rect 4480 0 4620 5
rect 4648 0 4676 4544
rect 4704 66 4732 4610
rect 4760 4605 4900 4610
rect 4760 4603 4802 4605
rect 4858 4603 4900 4605
rect 4760 4551 4772 4603
rect 4888 4551 4900 4603
rect 4760 4549 4802 4551
rect 4858 4549 4900 4551
rect 4760 4544 4900 4549
rect 4760 94 4788 4544
rect 4816 66 4844 4516
rect 4704 61 4844 66
rect 4704 59 4746 61
rect 4802 59 4844 61
rect 4704 7 4716 59
rect 4832 7 4844 59
rect 4704 5 4746 7
rect 4802 5 4844 7
rect 4704 0 4844 5
rect 4872 0 4900 4544
rect 4928 66 4956 4610
rect 4984 4605 5124 4610
rect 4984 4603 5026 4605
rect 5082 4603 5124 4605
rect 4984 4551 4996 4603
rect 5112 4551 5124 4603
rect 4984 4549 5026 4551
rect 5082 4549 5124 4551
rect 4984 4544 5124 4549
rect 4984 94 5012 4544
rect 5040 66 5068 4516
rect 4928 61 5068 66
rect 4928 59 4970 61
rect 5026 59 5068 61
rect 4928 7 4940 59
rect 5056 7 5068 59
rect 4928 5 4970 7
rect 5026 5 5068 7
rect 4928 0 5068 5
rect 5096 0 5124 4544
rect 5152 66 5180 4610
rect 5208 4605 5348 4610
rect 5208 4603 5250 4605
rect 5306 4603 5348 4605
rect 5208 4551 5220 4603
rect 5336 4551 5348 4603
rect 5208 4549 5250 4551
rect 5306 4549 5348 4551
rect 5208 4544 5348 4549
rect 5208 94 5236 4544
rect 5264 66 5292 4516
rect 5152 61 5292 66
rect 5152 59 5194 61
rect 5250 59 5292 61
rect 5152 7 5164 59
rect 5280 7 5292 59
rect 5152 5 5194 7
rect 5250 5 5292 7
rect 5152 0 5292 5
rect 5320 0 5348 4544
rect 5376 66 5404 4610
rect 5432 4605 5572 4610
rect 5432 4603 5474 4605
rect 5530 4603 5572 4605
rect 5432 4551 5444 4603
rect 5560 4551 5572 4603
rect 5432 4549 5474 4551
rect 5530 4549 5572 4551
rect 5432 4544 5572 4549
rect 5432 94 5460 4544
rect 5488 66 5516 4516
rect 5376 61 5516 66
rect 5376 59 5418 61
rect 5474 59 5516 61
rect 5376 7 5388 59
rect 5504 7 5516 59
rect 5376 5 5418 7
rect 5474 5 5516 7
rect 5376 0 5516 5
rect 5544 0 5572 4544
rect 5600 66 5628 4610
rect 5656 4605 5796 4610
rect 5656 4603 5698 4605
rect 5754 4603 5796 4605
rect 5656 4551 5668 4603
rect 5784 4551 5796 4603
rect 5656 4549 5698 4551
rect 5754 4549 5796 4551
rect 5656 4544 5796 4549
rect 5656 94 5684 4544
rect 5712 66 5740 4516
rect 5600 61 5740 66
rect 5600 59 5642 61
rect 5698 59 5740 61
rect 5600 7 5612 59
rect 5728 7 5740 59
rect 5600 5 5642 7
rect 5698 5 5740 7
rect 5600 0 5740 5
rect 5768 0 5796 4544
rect 5824 66 5852 4610
rect 5880 4605 6020 4610
rect 5880 4603 5922 4605
rect 5978 4603 6020 4605
rect 5880 4551 5892 4603
rect 6008 4551 6020 4603
rect 5880 4549 5922 4551
rect 5978 4549 6020 4551
rect 5880 4544 6020 4549
rect 5880 94 5908 4544
rect 5936 66 5964 4516
rect 5824 61 5964 66
rect 5824 59 5866 61
rect 5922 59 5964 61
rect 5824 7 5836 59
rect 5952 7 5964 59
rect 5824 5 5866 7
rect 5922 5 5964 7
rect 5824 0 5964 5
rect 5992 0 6020 4544
rect 6048 66 6076 4610
rect 6104 4605 6244 4610
rect 6104 4603 6146 4605
rect 6202 4603 6244 4605
rect 6104 4551 6116 4603
rect 6232 4551 6244 4603
rect 6104 4549 6146 4551
rect 6202 4549 6244 4551
rect 6104 4544 6244 4549
rect 6104 94 6132 4544
rect 6160 66 6188 4516
rect 6048 61 6188 66
rect 6048 59 6090 61
rect 6146 59 6188 61
rect 6048 7 6060 59
rect 6176 7 6188 59
rect 6048 5 6090 7
rect 6146 5 6188 7
rect 6048 0 6188 5
rect 6216 0 6244 4544
rect 6272 66 6300 4610
rect 6328 4605 6468 4610
rect 6328 4603 6370 4605
rect 6426 4603 6468 4605
rect 6328 4551 6340 4603
rect 6456 4551 6468 4603
rect 6328 4549 6370 4551
rect 6426 4549 6468 4551
rect 6328 4544 6468 4549
rect 6328 94 6356 4544
rect 6384 66 6412 4516
rect 6272 61 6412 66
rect 6272 59 6314 61
rect 6370 59 6412 61
rect 6272 7 6284 59
rect 6400 7 6412 59
rect 6272 5 6314 7
rect 6370 5 6412 7
rect 6272 0 6412 5
rect 6440 0 6468 4544
rect 6496 66 6524 4610
rect 6552 4605 6692 4610
rect 6552 4603 6594 4605
rect 6650 4603 6692 4605
rect 6552 4551 6564 4603
rect 6680 4551 6692 4603
rect 6552 4549 6594 4551
rect 6650 4549 6692 4551
rect 6552 4544 6692 4549
rect 6552 94 6580 4544
rect 6608 66 6636 4516
rect 6496 61 6636 66
rect 6496 59 6538 61
rect 6594 59 6636 61
rect 6496 7 6508 59
rect 6624 7 6636 59
rect 6496 5 6538 7
rect 6594 5 6636 7
rect 6496 0 6636 5
rect 6664 0 6692 4544
rect 6720 66 6748 4610
rect 6776 4605 6916 4610
rect 6776 4603 6818 4605
rect 6874 4603 6916 4605
rect 6776 4551 6788 4603
rect 6904 4551 6916 4603
rect 6776 4549 6818 4551
rect 6874 4549 6916 4551
rect 6776 4544 6916 4549
rect 6776 94 6804 4544
rect 6832 66 6860 4516
rect 6720 61 6860 66
rect 6720 59 6762 61
rect 6818 59 6860 61
rect 6720 7 6732 59
rect 6848 7 6860 59
rect 6720 5 6762 7
rect 6818 5 6860 7
rect 6720 0 6860 5
rect 6888 0 6916 4544
rect 6944 66 6972 4610
rect 7000 4605 7140 4610
rect 7000 4603 7042 4605
rect 7098 4603 7140 4605
rect 7000 4551 7012 4603
rect 7128 4551 7140 4603
rect 7000 4549 7042 4551
rect 7098 4549 7140 4551
rect 7000 4544 7140 4549
rect 7000 94 7028 4544
rect 7056 66 7084 4516
rect 6944 61 7084 66
rect 6944 59 6986 61
rect 7042 59 7084 61
rect 6944 7 6956 59
rect 7072 7 7084 59
rect 6944 5 6986 7
rect 7042 5 7084 7
rect 6944 0 7084 5
rect 7112 0 7140 4544
rect 7168 66 7196 4610
rect 7224 4605 7364 4610
rect 7224 4603 7266 4605
rect 7322 4603 7364 4605
rect 7224 4551 7236 4603
rect 7352 4551 7364 4603
rect 7224 4549 7266 4551
rect 7322 4549 7364 4551
rect 7224 4544 7364 4549
rect 7224 94 7252 4544
rect 7280 66 7308 4516
rect 7168 61 7308 66
rect 7168 59 7210 61
rect 7266 59 7308 61
rect 7168 7 7180 59
rect 7296 7 7308 59
rect 7168 5 7210 7
rect 7266 5 7308 7
rect 7168 0 7308 5
rect 7336 0 7364 4544
rect 7392 66 7420 4610
rect 7448 4605 7588 4610
rect 7448 4603 7490 4605
rect 7546 4603 7588 4605
rect 7448 4551 7460 4603
rect 7576 4551 7588 4603
rect 7448 4549 7490 4551
rect 7546 4549 7588 4551
rect 7448 4544 7588 4549
rect 7448 94 7476 4544
rect 7504 66 7532 4516
rect 7392 61 7532 66
rect 7392 59 7434 61
rect 7490 59 7532 61
rect 7392 7 7404 59
rect 7520 7 7532 59
rect 7392 5 7434 7
rect 7490 5 7532 7
rect 7392 0 7532 5
rect 7560 0 7588 4544
rect 7616 66 7644 4610
rect 7672 4605 7812 4610
rect 7672 4603 7714 4605
rect 7770 4603 7812 4605
rect 7672 4551 7684 4603
rect 7800 4551 7812 4603
rect 7672 4549 7714 4551
rect 7770 4549 7812 4551
rect 7672 4544 7812 4549
rect 7672 94 7700 4544
rect 7728 66 7756 4516
rect 7616 61 7756 66
rect 7616 59 7658 61
rect 7714 59 7756 61
rect 7616 7 7628 59
rect 7744 7 7756 59
rect 7616 5 7658 7
rect 7714 5 7756 7
rect 7616 0 7756 5
rect 7784 0 7812 4544
rect 7840 66 7868 4610
rect 7896 4605 8036 4610
rect 7896 4603 7938 4605
rect 7994 4603 8036 4605
rect 7896 4551 7908 4603
rect 8024 4551 8036 4603
rect 7896 4549 7938 4551
rect 7994 4549 8036 4551
rect 7896 4544 8036 4549
rect 7896 94 7924 4544
rect 7952 66 7980 4516
rect 7840 61 7980 66
rect 7840 59 7882 61
rect 7938 59 7980 61
rect 7840 7 7852 59
rect 7968 7 7980 59
rect 7840 5 7882 7
rect 7938 5 7980 7
rect 7840 0 7980 5
rect 8008 0 8036 4544
rect 8064 66 8092 4610
rect 8120 4605 8260 4610
rect 8120 4603 8162 4605
rect 8218 4603 8260 4605
rect 8120 4551 8132 4603
rect 8248 4551 8260 4603
rect 8120 4549 8162 4551
rect 8218 4549 8260 4551
rect 8120 4544 8260 4549
rect 8120 94 8148 4544
rect 8176 66 8204 4516
rect 8064 61 8204 66
rect 8064 59 8106 61
rect 8162 59 8204 61
rect 8064 7 8076 59
rect 8192 7 8204 59
rect 8064 5 8106 7
rect 8162 5 8204 7
rect 8064 0 8204 5
rect 8232 0 8260 4544
rect 8288 66 8316 4610
rect 8344 4605 8484 4610
rect 8344 4603 8386 4605
rect 8442 4603 8484 4605
rect 8344 4551 8356 4603
rect 8472 4551 8484 4603
rect 8344 4549 8386 4551
rect 8442 4549 8484 4551
rect 8344 4544 8484 4549
rect 8344 94 8372 4544
rect 8400 66 8428 4516
rect 8288 61 8428 66
rect 8288 59 8330 61
rect 8386 59 8428 61
rect 8288 7 8300 59
rect 8416 7 8428 59
rect 8288 5 8330 7
rect 8386 5 8428 7
rect 8288 0 8428 5
rect 8456 0 8484 4544
rect 8512 66 8540 4610
rect 8568 4605 8708 4610
rect 8568 4603 8610 4605
rect 8666 4603 8708 4605
rect 8568 4551 8580 4603
rect 8696 4551 8708 4603
rect 8568 4549 8610 4551
rect 8666 4549 8708 4551
rect 8568 4544 8708 4549
rect 8568 94 8596 4544
rect 8624 66 8652 4516
rect 8512 61 8652 66
rect 8512 59 8554 61
rect 8610 59 8652 61
rect 8512 7 8524 59
rect 8640 7 8652 59
rect 8512 5 8554 7
rect 8610 5 8652 7
rect 8512 0 8652 5
rect 8680 0 8708 4544
rect 8736 66 8764 4610
rect 8792 4605 8932 4610
rect 8792 4603 8834 4605
rect 8890 4603 8932 4605
rect 8792 4551 8804 4603
rect 8920 4551 8932 4603
rect 8792 4549 8834 4551
rect 8890 4549 8932 4551
rect 8792 4544 8932 4549
rect 8792 94 8820 4544
rect 8848 66 8876 4516
rect 8736 61 8876 66
rect 8736 59 8778 61
rect 8834 59 8876 61
rect 8736 7 8748 59
rect 8864 7 8876 59
rect 8736 5 8778 7
rect 8834 5 8876 7
rect 8736 0 8876 5
rect 8904 0 8932 4544
rect 8960 66 8988 4610
rect 9016 4605 9156 4610
rect 9016 4603 9058 4605
rect 9114 4603 9156 4605
rect 9016 4551 9028 4603
rect 9144 4551 9156 4603
rect 9016 4549 9058 4551
rect 9114 4549 9156 4551
rect 9016 4544 9156 4549
rect 9016 94 9044 4544
rect 9072 66 9100 4516
rect 8960 61 9100 66
rect 8960 59 9002 61
rect 9058 59 9100 61
rect 8960 7 8972 59
rect 9088 7 9100 59
rect 8960 5 9002 7
rect 9058 5 9100 7
rect 8960 0 9100 5
rect 9128 0 9156 4544
rect 9184 66 9212 4610
rect 9240 4605 9380 4610
rect 9240 4603 9282 4605
rect 9338 4603 9380 4605
rect 9240 4551 9252 4603
rect 9368 4551 9380 4603
rect 9240 4549 9282 4551
rect 9338 4549 9380 4551
rect 9240 4544 9380 4549
rect 9240 94 9268 4544
rect 9296 66 9324 4516
rect 9184 61 9324 66
rect 9184 59 9226 61
rect 9282 59 9324 61
rect 9184 7 9196 59
rect 9312 7 9324 59
rect 9184 5 9226 7
rect 9282 5 9324 7
rect 9184 0 9324 5
rect 9352 0 9380 4544
rect 9408 66 9436 4610
rect 9464 4605 9604 4610
rect 9464 4603 9506 4605
rect 9562 4603 9604 4605
rect 9464 4551 9476 4603
rect 9592 4551 9604 4603
rect 9464 4549 9506 4551
rect 9562 4549 9604 4551
rect 9464 4544 9604 4549
rect 9464 94 9492 4544
rect 9520 66 9548 4516
rect 9408 61 9548 66
rect 9408 59 9450 61
rect 9506 59 9548 61
rect 9408 7 9420 59
rect 9536 7 9548 59
rect 9408 5 9450 7
rect 9506 5 9548 7
rect 9408 0 9548 5
rect 9576 0 9604 4544
rect 9632 66 9660 4610
rect 9688 4605 9828 4610
rect 9688 4603 9730 4605
rect 9786 4603 9828 4605
rect 9688 4551 9700 4603
rect 9816 4551 9828 4603
rect 9688 4549 9730 4551
rect 9786 4549 9828 4551
rect 9688 4544 9828 4549
rect 9688 94 9716 4544
rect 9744 66 9772 4516
rect 9632 61 9772 66
rect 9632 59 9674 61
rect 9730 59 9772 61
rect 9632 7 9644 59
rect 9760 7 9772 59
rect 9632 5 9674 7
rect 9730 5 9772 7
rect 9632 0 9772 5
rect 9800 0 9828 4544
rect 9856 66 9884 4610
rect 9912 4605 10052 4610
rect 9912 4603 9954 4605
rect 10010 4603 10052 4605
rect 9912 4551 9924 4603
rect 10040 4551 10052 4603
rect 9912 4549 9954 4551
rect 10010 4549 10052 4551
rect 9912 4544 10052 4549
rect 9912 94 9940 4544
rect 9968 66 9996 4516
rect 9856 61 9996 66
rect 9856 59 9898 61
rect 9954 59 9996 61
rect 9856 7 9868 59
rect 9984 7 9996 59
rect 9856 5 9898 7
rect 9954 5 9996 7
rect 9856 0 9996 5
rect 10024 0 10052 4544
rect 10080 66 10108 4610
rect 10136 4605 10276 4610
rect 10136 4603 10178 4605
rect 10234 4603 10276 4605
rect 10136 4551 10148 4603
rect 10264 4551 10276 4603
rect 10136 4549 10178 4551
rect 10234 4549 10276 4551
rect 10136 4544 10276 4549
rect 10136 94 10164 4544
rect 10192 66 10220 4516
rect 10080 61 10220 66
rect 10080 59 10122 61
rect 10178 59 10220 61
rect 10080 7 10092 59
rect 10208 7 10220 59
rect 10080 5 10122 7
rect 10178 5 10220 7
rect 10080 0 10220 5
rect 10248 0 10276 4544
rect 10304 66 10332 4610
rect 10360 4605 10500 4610
rect 10360 4603 10402 4605
rect 10458 4603 10500 4605
rect 10360 4551 10372 4603
rect 10488 4551 10500 4603
rect 10360 4549 10402 4551
rect 10458 4549 10500 4551
rect 10360 4544 10500 4549
rect 10360 94 10388 4544
rect 10416 66 10444 4516
rect 10304 61 10444 66
rect 10304 59 10346 61
rect 10402 59 10444 61
rect 10304 7 10316 59
rect 10432 7 10444 59
rect 10304 5 10346 7
rect 10402 5 10444 7
rect 10304 0 10444 5
rect 10472 0 10500 4544
rect 10528 66 10556 4610
rect 10584 4605 10724 4610
rect 10584 4603 10626 4605
rect 10682 4603 10724 4605
rect 10584 4551 10596 4603
rect 10712 4551 10724 4603
rect 10584 4549 10626 4551
rect 10682 4549 10724 4551
rect 10584 4544 10724 4549
rect 10584 94 10612 4544
rect 10640 66 10668 4516
rect 10528 61 10668 66
rect 10528 59 10570 61
rect 10626 59 10668 61
rect 10528 7 10540 59
rect 10656 7 10668 59
rect 10528 5 10570 7
rect 10626 5 10668 7
rect 10528 0 10668 5
rect 10696 0 10724 4544
rect 10752 66 10780 4610
rect 10808 4605 11146 4610
rect 10808 4603 10850 4605
rect 10906 4603 11146 4605
rect 10808 4551 10820 4603
rect 10936 4551 11146 4603
rect 10808 4549 10850 4551
rect 10906 4549 11146 4551
rect 10808 4544 11146 4549
rect 10808 94 10836 4544
rect 10864 66 10892 4516
rect 10752 61 10892 66
rect 10752 59 10794 61
rect 10850 59 10892 61
rect 10752 7 10764 59
rect 10880 7 10892 59
rect 10752 5 10794 7
rect 10850 5 10892 7
rect 10752 0 10892 5
rect 10920 0 10948 4544
rect 10976 66 11004 4516
rect 11032 94 11060 4544
rect 11088 66 11146 4516
rect 10976 61 11146 66
rect 10976 59 11018 61
rect 11074 59 11146 61
rect 10976 7 10988 59
rect 11104 7 11146 59
rect 10976 5 11018 7
rect 11074 5 11146 7
rect 10976 0 11146 5
<< via2 >>
rect 98 4603 154 4605
rect 98 4551 120 4603
rect 120 4551 132 4603
rect 132 4551 154 4603
rect 98 4549 154 4551
rect 42 59 98 61
rect 42 7 76 59
rect 76 7 88 59
rect 88 7 98 59
rect 42 5 98 7
rect 322 4603 378 4605
rect 322 4551 344 4603
rect 344 4551 356 4603
rect 356 4551 378 4603
rect 322 4549 378 4551
rect 266 59 322 61
rect 266 7 288 59
rect 288 7 300 59
rect 300 7 322 59
rect 266 5 322 7
rect 546 4603 602 4605
rect 546 4551 568 4603
rect 568 4551 580 4603
rect 580 4551 602 4603
rect 546 4549 602 4551
rect 490 59 546 61
rect 490 7 512 59
rect 512 7 524 59
rect 524 7 546 59
rect 490 5 546 7
rect 770 4603 826 4605
rect 770 4551 792 4603
rect 792 4551 804 4603
rect 804 4551 826 4603
rect 770 4549 826 4551
rect 714 59 770 61
rect 714 7 736 59
rect 736 7 748 59
rect 748 7 770 59
rect 714 5 770 7
rect 994 4603 1050 4605
rect 994 4551 1016 4603
rect 1016 4551 1028 4603
rect 1028 4551 1050 4603
rect 994 4549 1050 4551
rect 938 59 994 61
rect 938 7 960 59
rect 960 7 972 59
rect 972 7 994 59
rect 938 5 994 7
rect 1218 4603 1274 4605
rect 1218 4551 1240 4603
rect 1240 4551 1252 4603
rect 1252 4551 1274 4603
rect 1218 4549 1274 4551
rect 1162 59 1218 61
rect 1162 7 1184 59
rect 1184 7 1196 59
rect 1196 7 1218 59
rect 1162 5 1218 7
rect 1442 4603 1498 4605
rect 1442 4551 1464 4603
rect 1464 4551 1476 4603
rect 1476 4551 1498 4603
rect 1442 4549 1498 4551
rect 1386 59 1442 61
rect 1386 7 1408 59
rect 1408 7 1420 59
rect 1420 7 1442 59
rect 1386 5 1442 7
rect 1666 4603 1722 4605
rect 1666 4551 1688 4603
rect 1688 4551 1700 4603
rect 1700 4551 1722 4603
rect 1666 4549 1722 4551
rect 1610 59 1666 61
rect 1610 7 1632 59
rect 1632 7 1644 59
rect 1644 7 1666 59
rect 1610 5 1666 7
rect 1890 4603 1946 4605
rect 1890 4551 1912 4603
rect 1912 4551 1924 4603
rect 1924 4551 1946 4603
rect 1890 4549 1946 4551
rect 1834 59 1890 61
rect 1834 7 1856 59
rect 1856 7 1868 59
rect 1868 7 1890 59
rect 1834 5 1890 7
rect 2114 4603 2170 4605
rect 2114 4551 2136 4603
rect 2136 4551 2148 4603
rect 2148 4551 2170 4603
rect 2114 4549 2170 4551
rect 2058 59 2114 61
rect 2058 7 2080 59
rect 2080 7 2092 59
rect 2092 7 2114 59
rect 2058 5 2114 7
rect 2338 4603 2394 4605
rect 2338 4551 2360 4603
rect 2360 4551 2372 4603
rect 2372 4551 2394 4603
rect 2338 4549 2394 4551
rect 2282 59 2338 61
rect 2282 7 2304 59
rect 2304 7 2316 59
rect 2316 7 2338 59
rect 2282 5 2338 7
rect 2562 4603 2618 4605
rect 2562 4551 2584 4603
rect 2584 4551 2596 4603
rect 2596 4551 2618 4603
rect 2562 4549 2618 4551
rect 2506 59 2562 61
rect 2506 7 2528 59
rect 2528 7 2540 59
rect 2540 7 2562 59
rect 2506 5 2562 7
rect 2786 4603 2842 4605
rect 2786 4551 2808 4603
rect 2808 4551 2820 4603
rect 2820 4551 2842 4603
rect 2786 4549 2842 4551
rect 2730 59 2786 61
rect 2730 7 2752 59
rect 2752 7 2764 59
rect 2764 7 2786 59
rect 2730 5 2786 7
rect 3010 4603 3066 4605
rect 3010 4551 3032 4603
rect 3032 4551 3044 4603
rect 3044 4551 3066 4603
rect 3010 4549 3066 4551
rect 2954 59 3010 61
rect 2954 7 2976 59
rect 2976 7 2988 59
rect 2988 7 3010 59
rect 2954 5 3010 7
rect 3234 4603 3290 4605
rect 3234 4551 3256 4603
rect 3256 4551 3268 4603
rect 3268 4551 3290 4603
rect 3234 4549 3290 4551
rect 3178 59 3234 61
rect 3178 7 3200 59
rect 3200 7 3212 59
rect 3212 7 3234 59
rect 3178 5 3234 7
rect 3458 4603 3514 4605
rect 3458 4551 3480 4603
rect 3480 4551 3492 4603
rect 3492 4551 3514 4603
rect 3458 4549 3514 4551
rect 3402 59 3458 61
rect 3402 7 3424 59
rect 3424 7 3436 59
rect 3436 7 3458 59
rect 3402 5 3458 7
rect 3682 4603 3738 4605
rect 3682 4551 3704 4603
rect 3704 4551 3716 4603
rect 3716 4551 3738 4603
rect 3682 4549 3738 4551
rect 3626 59 3682 61
rect 3626 7 3648 59
rect 3648 7 3660 59
rect 3660 7 3682 59
rect 3626 5 3682 7
rect 3906 4603 3962 4605
rect 3906 4551 3928 4603
rect 3928 4551 3940 4603
rect 3940 4551 3962 4603
rect 3906 4549 3962 4551
rect 3850 59 3906 61
rect 3850 7 3872 59
rect 3872 7 3884 59
rect 3884 7 3906 59
rect 3850 5 3906 7
rect 4130 4603 4186 4605
rect 4130 4551 4152 4603
rect 4152 4551 4164 4603
rect 4164 4551 4186 4603
rect 4130 4549 4186 4551
rect 4074 59 4130 61
rect 4074 7 4096 59
rect 4096 7 4108 59
rect 4108 7 4130 59
rect 4074 5 4130 7
rect 4354 4603 4410 4605
rect 4354 4551 4376 4603
rect 4376 4551 4388 4603
rect 4388 4551 4410 4603
rect 4354 4549 4410 4551
rect 4298 59 4354 61
rect 4298 7 4320 59
rect 4320 7 4332 59
rect 4332 7 4354 59
rect 4298 5 4354 7
rect 4578 4603 4634 4605
rect 4578 4551 4600 4603
rect 4600 4551 4612 4603
rect 4612 4551 4634 4603
rect 4578 4549 4634 4551
rect 4522 59 4578 61
rect 4522 7 4544 59
rect 4544 7 4556 59
rect 4556 7 4578 59
rect 4522 5 4578 7
rect 4802 4603 4858 4605
rect 4802 4551 4824 4603
rect 4824 4551 4836 4603
rect 4836 4551 4858 4603
rect 4802 4549 4858 4551
rect 4746 59 4802 61
rect 4746 7 4768 59
rect 4768 7 4780 59
rect 4780 7 4802 59
rect 4746 5 4802 7
rect 5026 4603 5082 4605
rect 5026 4551 5048 4603
rect 5048 4551 5060 4603
rect 5060 4551 5082 4603
rect 5026 4549 5082 4551
rect 4970 59 5026 61
rect 4970 7 4992 59
rect 4992 7 5004 59
rect 5004 7 5026 59
rect 4970 5 5026 7
rect 5250 4603 5306 4605
rect 5250 4551 5272 4603
rect 5272 4551 5284 4603
rect 5284 4551 5306 4603
rect 5250 4549 5306 4551
rect 5194 59 5250 61
rect 5194 7 5216 59
rect 5216 7 5228 59
rect 5228 7 5250 59
rect 5194 5 5250 7
rect 5474 4603 5530 4605
rect 5474 4551 5496 4603
rect 5496 4551 5508 4603
rect 5508 4551 5530 4603
rect 5474 4549 5530 4551
rect 5418 59 5474 61
rect 5418 7 5440 59
rect 5440 7 5452 59
rect 5452 7 5474 59
rect 5418 5 5474 7
rect 5698 4603 5754 4605
rect 5698 4551 5720 4603
rect 5720 4551 5732 4603
rect 5732 4551 5754 4603
rect 5698 4549 5754 4551
rect 5642 59 5698 61
rect 5642 7 5664 59
rect 5664 7 5676 59
rect 5676 7 5698 59
rect 5642 5 5698 7
rect 5922 4603 5978 4605
rect 5922 4551 5944 4603
rect 5944 4551 5956 4603
rect 5956 4551 5978 4603
rect 5922 4549 5978 4551
rect 5866 59 5922 61
rect 5866 7 5888 59
rect 5888 7 5900 59
rect 5900 7 5922 59
rect 5866 5 5922 7
rect 6146 4603 6202 4605
rect 6146 4551 6168 4603
rect 6168 4551 6180 4603
rect 6180 4551 6202 4603
rect 6146 4549 6202 4551
rect 6090 59 6146 61
rect 6090 7 6112 59
rect 6112 7 6124 59
rect 6124 7 6146 59
rect 6090 5 6146 7
rect 6370 4603 6426 4605
rect 6370 4551 6392 4603
rect 6392 4551 6404 4603
rect 6404 4551 6426 4603
rect 6370 4549 6426 4551
rect 6314 59 6370 61
rect 6314 7 6336 59
rect 6336 7 6348 59
rect 6348 7 6370 59
rect 6314 5 6370 7
rect 6594 4603 6650 4605
rect 6594 4551 6616 4603
rect 6616 4551 6628 4603
rect 6628 4551 6650 4603
rect 6594 4549 6650 4551
rect 6538 59 6594 61
rect 6538 7 6560 59
rect 6560 7 6572 59
rect 6572 7 6594 59
rect 6538 5 6594 7
rect 6818 4603 6874 4605
rect 6818 4551 6840 4603
rect 6840 4551 6852 4603
rect 6852 4551 6874 4603
rect 6818 4549 6874 4551
rect 6762 59 6818 61
rect 6762 7 6784 59
rect 6784 7 6796 59
rect 6796 7 6818 59
rect 6762 5 6818 7
rect 7042 4603 7098 4605
rect 7042 4551 7064 4603
rect 7064 4551 7076 4603
rect 7076 4551 7098 4603
rect 7042 4549 7098 4551
rect 6986 59 7042 61
rect 6986 7 7008 59
rect 7008 7 7020 59
rect 7020 7 7042 59
rect 6986 5 7042 7
rect 7266 4603 7322 4605
rect 7266 4551 7288 4603
rect 7288 4551 7300 4603
rect 7300 4551 7322 4603
rect 7266 4549 7322 4551
rect 7210 59 7266 61
rect 7210 7 7232 59
rect 7232 7 7244 59
rect 7244 7 7266 59
rect 7210 5 7266 7
rect 7490 4603 7546 4605
rect 7490 4551 7512 4603
rect 7512 4551 7524 4603
rect 7524 4551 7546 4603
rect 7490 4549 7546 4551
rect 7434 59 7490 61
rect 7434 7 7456 59
rect 7456 7 7468 59
rect 7468 7 7490 59
rect 7434 5 7490 7
rect 7714 4603 7770 4605
rect 7714 4551 7736 4603
rect 7736 4551 7748 4603
rect 7748 4551 7770 4603
rect 7714 4549 7770 4551
rect 7658 59 7714 61
rect 7658 7 7680 59
rect 7680 7 7692 59
rect 7692 7 7714 59
rect 7658 5 7714 7
rect 7938 4603 7994 4605
rect 7938 4551 7960 4603
rect 7960 4551 7972 4603
rect 7972 4551 7994 4603
rect 7938 4549 7994 4551
rect 7882 59 7938 61
rect 7882 7 7904 59
rect 7904 7 7916 59
rect 7916 7 7938 59
rect 7882 5 7938 7
rect 8162 4603 8218 4605
rect 8162 4551 8184 4603
rect 8184 4551 8196 4603
rect 8196 4551 8218 4603
rect 8162 4549 8218 4551
rect 8106 59 8162 61
rect 8106 7 8128 59
rect 8128 7 8140 59
rect 8140 7 8162 59
rect 8106 5 8162 7
rect 8386 4603 8442 4605
rect 8386 4551 8408 4603
rect 8408 4551 8420 4603
rect 8420 4551 8442 4603
rect 8386 4549 8442 4551
rect 8330 59 8386 61
rect 8330 7 8352 59
rect 8352 7 8364 59
rect 8364 7 8386 59
rect 8330 5 8386 7
rect 8610 4603 8666 4605
rect 8610 4551 8632 4603
rect 8632 4551 8644 4603
rect 8644 4551 8666 4603
rect 8610 4549 8666 4551
rect 8554 59 8610 61
rect 8554 7 8576 59
rect 8576 7 8588 59
rect 8588 7 8610 59
rect 8554 5 8610 7
rect 8834 4603 8890 4605
rect 8834 4551 8856 4603
rect 8856 4551 8868 4603
rect 8868 4551 8890 4603
rect 8834 4549 8890 4551
rect 8778 59 8834 61
rect 8778 7 8800 59
rect 8800 7 8812 59
rect 8812 7 8834 59
rect 8778 5 8834 7
rect 9058 4603 9114 4605
rect 9058 4551 9080 4603
rect 9080 4551 9092 4603
rect 9092 4551 9114 4603
rect 9058 4549 9114 4551
rect 9002 59 9058 61
rect 9002 7 9024 59
rect 9024 7 9036 59
rect 9036 7 9058 59
rect 9002 5 9058 7
rect 9282 4603 9338 4605
rect 9282 4551 9304 4603
rect 9304 4551 9316 4603
rect 9316 4551 9338 4603
rect 9282 4549 9338 4551
rect 9226 59 9282 61
rect 9226 7 9248 59
rect 9248 7 9260 59
rect 9260 7 9282 59
rect 9226 5 9282 7
rect 9506 4603 9562 4605
rect 9506 4551 9528 4603
rect 9528 4551 9540 4603
rect 9540 4551 9562 4603
rect 9506 4549 9562 4551
rect 9450 59 9506 61
rect 9450 7 9472 59
rect 9472 7 9484 59
rect 9484 7 9506 59
rect 9450 5 9506 7
rect 9730 4603 9786 4605
rect 9730 4551 9752 4603
rect 9752 4551 9764 4603
rect 9764 4551 9786 4603
rect 9730 4549 9786 4551
rect 9674 59 9730 61
rect 9674 7 9696 59
rect 9696 7 9708 59
rect 9708 7 9730 59
rect 9674 5 9730 7
rect 9954 4603 10010 4605
rect 9954 4551 9976 4603
rect 9976 4551 9988 4603
rect 9988 4551 10010 4603
rect 9954 4549 10010 4551
rect 9898 59 9954 61
rect 9898 7 9920 59
rect 9920 7 9932 59
rect 9932 7 9954 59
rect 9898 5 9954 7
rect 10178 4603 10234 4605
rect 10178 4551 10200 4603
rect 10200 4551 10212 4603
rect 10212 4551 10234 4603
rect 10178 4549 10234 4551
rect 10122 59 10178 61
rect 10122 7 10144 59
rect 10144 7 10156 59
rect 10156 7 10178 59
rect 10122 5 10178 7
rect 10402 4603 10458 4605
rect 10402 4551 10424 4603
rect 10424 4551 10436 4603
rect 10436 4551 10458 4603
rect 10402 4549 10458 4551
rect 10346 59 10402 61
rect 10346 7 10368 59
rect 10368 7 10380 59
rect 10380 7 10402 59
rect 10346 5 10402 7
rect 10626 4603 10682 4605
rect 10626 4551 10648 4603
rect 10648 4551 10660 4603
rect 10660 4551 10682 4603
rect 10626 4549 10682 4551
rect 10570 59 10626 61
rect 10570 7 10592 59
rect 10592 7 10604 59
rect 10604 7 10626 59
rect 10570 5 10626 7
rect 10850 4603 10906 4605
rect 10850 4551 10872 4603
rect 10872 4551 10884 4603
rect 10884 4551 10906 4603
rect 10850 4549 10906 4551
rect 10794 59 10850 61
rect 10794 7 10816 59
rect 10816 7 10828 59
rect 10828 7 10850 59
rect 10794 5 10850 7
rect 11018 59 11074 61
rect 11018 7 11040 59
rect 11040 7 11052 59
rect 11052 7 11074 59
rect 11018 5 11074 7
<< metal3 >>
rect 0 4609 11146 4610
rect 0 4545 28 4609
rect 92 4605 108 4609
rect 92 4549 98 4605
rect 92 4545 108 4549
rect 172 4545 188 4609
rect 252 4545 268 4609
rect 332 4605 348 4609
rect 332 4545 348 4549
rect 412 4545 428 4609
rect 492 4545 508 4609
rect 572 4605 588 4609
rect 572 4545 588 4549
rect 652 4545 668 4609
rect 732 4545 748 4609
rect 812 4605 828 4609
rect 826 4549 828 4605
rect 812 4545 828 4549
rect 892 4545 908 4609
rect 972 4545 988 4609
rect 1052 4545 1068 4609
rect 1132 4545 1148 4609
rect 1212 4605 1228 4609
rect 1212 4549 1218 4605
rect 1212 4545 1228 4549
rect 1292 4545 1308 4609
rect 1372 4545 1388 4609
rect 1452 4605 1468 4609
rect 1452 4545 1468 4549
rect 1532 4545 1548 4609
rect 1612 4545 1628 4609
rect 1692 4605 1708 4609
rect 1692 4545 1708 4549
rect 1772 4545 1788 4609
rect 1852 4545 1868 4609
rect 1932 4605 1948 4609
rect 1946 4549 1948 4605
rect 1932 4545 1948 4549
rect 2012 4545 2028 4609
rect 2092 4545 2108 4609
rect 2172 4545 2188 4609
rect 2252 4545 2268 4609
rect 2332 4605 2348 4609
rect 2332 4549 2338 4605
rect 2332 4545 2348 4549
rect 2412 4545 2428 4609
rect 2492 4545 2508 4609
rect 2572 4605 2588 4609
rect 2572 4545 2588 4549
rect 2652 4545 2668 4609
rect 2732 4545 2748 4609
rect 2812 4605 2828 4609
rect 2812 4545 2828 4549
rect 2892 4545 2908 4609
rect 2972 4545 2988 4609
rect 3052 4605 3068 4609
rect 3066 4549 3068 4605
rect 3052 4545 3068 4549
rect 3132 4545 3148 4609
rect 3212 4545 3228 4609
rect 3292 4545 3308 4609
rect 3372 4545 3388 4609
rect 3452 4605 3468 4609
rect 3452 4549 3458 4605
rect 3452 4545 3468 4549
rect 3532 4545 3548 4609
rect 3612 4545 3628 4609
rect 3692 4605 3708 4609
rect 3692 4545 3708 4549
rect 3772 4545 3788 4609
rect 3852 4545 3868 4609
rect 3932 4605 3948 4609
rect 3932 4545 3948 4549
rect 4012 4545 4028 4609
rect 4092 4545 4108 4609
rect 4172 4605 4188 4609
rect 4186 4549 4188 4605
rect 4172 4545 4188 4549
rect 4252 4545 4268 4609
rect 4332 4545 4348 4609
rect 4412 4545 4428 4609
rect 4492 4545 4508 4609
rect 4572 4605 4588 4609
rect 4572 4549 4578 4605
rect 4572 4545 4588 4549
rect 4652 4545 4668 4609
rect 4732 4545 4748 4609
rect 4812 4605 4828 4609
rect 4812 4545 4828 4549
rect 4892 4545 4908 4609
rect 4972 4545 4988 4609
rect 5052 4605 5068 4609
rect 5052 4545 5068 4549
rect 5132 4545 5148 4609
rect 5212 4545 5228 4609
rect 5292 4605 5308 4609
rect 5306 4549 5308 4605
rect 5292 4545 5308 4549
rect 5372 4545 5388 4609
rect 5452 4545 5468 4609
rect 5532 4545 5548 4609
rect 5612 4545 5628 4609
rect 5692 4605 5708 4609
rect 5692 4549 5698 4605
rect 5692 4545 5708 4549
rect 5772 4545 5788 4609
rect 5852 4545 5868 4609
rect 5932 4605 5948 4609
rect 5932 4545 5948 4549
rect 6012 4545 6028 4609
rect 6092 4545 6108 4609
rect 6172 4605 6188 4609
rect 6172 4545 6188 4549
rect 6252 4545 6268 4609
rect 6332 4545 6348 4609
rect 6412 4605 6428 4609
rect 6426 4549 6428 4605
rect 6412 4545 6428 4549
rect 6492 4545 6508 4609
rect 6572 4545 6588 4609
rect 6652 4545 6668 4609
rect 6732 4545 6748 4609
rect 6812 4605 6828 4609
rect 6812 4549 6818 4605
rect 6812 4545 6828 4549
rect 6892 4545 6908 4609
rect 6972 4545 6988 4609
rect 7052 4605 7068 4609
rect 7052 4545 7068 4549
rect 7132 4545 7148 4609
rect 7212 4545 7228 4609
rect 7292 4605 7308 4609
rect 7292 4545 7308 4549
rect 7372 4545 7388 4609
rect 7452 4545 7468 4609
rect 7532 4605 7548 4609
rect 7546 4549 7548 4605
rect 7532 4545 7548 4549
rect 7612 4545 7628 4609
rect 7692 4545 7708 4609
rect 7772 4545 7788 4609
rect 7852 4545 7868 4609
rect 7932 4605 7948 4609
rect 7932 4549 7938 4605
rect 7932 4545 7948 4549
rect 8012 4545 8028 4609
rect 8092 4545 8108 4609
rect 8172 4605 8188 4609
rect 8172 4545 8188 4549
rect 8252 4545 8268 4609
rect 8332 4545 8348 4609
rect 8412 4605 8428 4609
rect 8412 4545 8428 4549
rect 8492 4545 8508 4609
rect 8572 4545 8588 4609
rect 8652 4605 8668 4609
rect 8666 4549 8668 4605
rect 8652 4545 8668 4549
rect 8732 4545 8748 4609
rect 8812 4545 8828 4609
rect 8892 4545 8908 4609
rect 8972 4545 8988 4609
rect 9052 4605 9068 4609
rect 9052 4549 9058 4605
rect 9052 4545 9068 4549
rect 9132 4545 9148 4609
rect 9212 4545 9228 4609
rect 9292 4605 9308 4609
rect 9292 4545 9308 4549
rect 9372 4545 9388 4609
rect 9452 4545 9468 4609
rect 9532 4605 9548 4609
rect 9532 4545 9548 4549
rect 9612 4545 9628 4609
rect 9692 4545 9708 4609
rect 9772 4605 9788 4609
rect 9786 4549 9788 4605
rect 9772 4545 9788 4549
rect 9852 4545 9868 4609
rect 9932 4545 9948 4609
rect 10012 4545 10028 4609
rect 10092 4545 10108 4609
rect 10172 4605 10188 4609
rect 10172 4549 10178 4605
rect 10172 4545 10188 4549
rect 10252 4545 10268 4609
rect 10332 4545 10348 4609
rect 10412 4605 10428 4609
rect 10412 4545 10428 4549
rect 10492 4545 10508 4609
rect 10572 4545 10588 4609
rect 10652 4605 10668 4609
rect 10652 4545 10668 4549
rect 10732 4545 10748 4609
rect 10812 4545 10828 4609
rect 10892 4605 10908 4609
rect 10906 4549 10908 4605
rect 10892 4545 10908 4549
rect 10972 4545 10988 4609
rect 11052 4545 11146 4609
rect 0 4544 11146 4545
rect 0 126 60 4544
rect 120 66 180 4484
rect 240 126 300 4544
rect 360 66 420 4484
rect 480 126 540 4544
rect 600 66 660 4484
rect 720 126 780 4544
rect 840 66 900 4484
rect 960 126 1020 4544
rect 1080 66 1140 4484
rect 1200 126 1260 4544
rect 1320 66 1380 4484
rect 1440 126 1500 4544
rect 1560 66 1620 4484
rect 1680 126 1740 4544
rect 1800 66 1860 4484
rect 1920 126 1980 4544
rect 2040 66 2100 4484
rect 2160 126 2220 4544
rect 2280 66 2340 4484
rect 2400 126 2460 4544
rect 2520 66 2580 4484
rect 2640 126 2700 4544
rect 2760 66 2820 4484
rect 2880 126 2940 4544
rect 3000 66 3060 4484
rect 3120 126 3180 4544
rect 3240 66 3300 4484
rect 3360 126 3420 4544
rect 3480 66 3540 4484
rect 3600 126 3660 4544
rect 3720 66 3780 4484
rect 3840 126 3900 4544
rect 3960 66 4020 4484
rect 4080 126 4140 4544
rect 4200 66 4260 4484
rect 4320 126 4380 4544
rect 4440 66 4500 4484
rect 4560 126 4620 4544
rect 4680 66 4740 4484
rect 4800 126 4860 4544
rect 4920 66 4980 4484
rect 5040 126 5100 4544
rect 5160 66 5220 4484
rect 5280 126 5340 4544
rect 5400 66 5460 4484
rect 5520 126 5580 4544
rect 5640 66 5700 4484
rect 5760 126 5820 4544
rect 5880 66 5940 4484
rect 6000 126 6060 4544
rect 6120 66 6180 4484
rect 6240 126 6300 4544
rect 6360 66 6420 4484
rect 6480 126 6540 4544
rect 6600 66 6660 4484
rect 6720 126 6780 4544
rect 6840 66 6900 4484
rect 6960 126 7020 4544
rect 7080 66 7140 4484
rect 7200 126 7260 4544
rect 7320 66 7380 4484
rect 7440 126 7500 4544
rect 7560 66 7620 4484
rect 7680 126 7740 4544
rect 7800 66 7860 4484
rect 7920 126 7980 4544
rect 8040 66 8100 4484
rect 8160 126 8220 4544
rect 8280 66 8340 4484
rect 8400 126 8460 4544
rect 8520 66 8580 4484
rect 8640 126 8700 4544
rect 8760 66 8820 4484
rect 8880 126 8940 4544
rect 9000 66 9060 4484
rect 9120 126 9180 4544
rect 9240 66 9300 4484
rect 9360 126 9420 4544
rect 9480 66 9540 4484
rect 9600 126 9660 4544
rect 9720 66 9780 4484
rect 9840 126 9900 4544
rect 9960 66 10020 4484
rect 10080 126 10140 4544
rect 10200 66 10260 4484
rect 10320 126 10380 4544
rect 10440 66 10500 4484
rect 10560 126 10620 4544
rect 10680 66 10740 4484
rect 10800 126 10860 4544
rect 10920 66 10980 4484
rect 11040 126 11146 4544
rect 0 65 11146 66
rect 0 1 28 65
rect 92 61 108 65
rect 98 5 108 61
rect 92 1 108 5
rect 172 1 188 65
rect 252 61 268 65
rect 252 5 266 61
rect 252 1 268 5
rect 332 1 348 65
rect 412 1 428 65
rect 492 61 508 65
rect 492 1 508 5
rect 572 1 588 65
rect 652 1 668 65
rect 732 61 748 65
rect 732 1 748 5
rect 812 1 828 65
rect 892 1 908 65
rect 972 61 988 65
rect 972 1 988 5
rect 1052 1 1068 65
rect 1132 1 1148 65
rect 1212 61 1228 65
rect 1218 5 1228 61
rect 1212 1 1228 5
rect 1292 1 1308 65
rect 1372 61 1388 65
rect 1372 5 1386 61
rect 1372 1 1388 5
rect 1452 1 1468 65
rect 1532 1 1548 65
rect 1612 61 1628 65
rect 1612 1 1628 5
rect 1692 1 1708 65
rect 1772 1 1788 65
rect 1852 61 1868 65
rect 1852 1 1868 5
rect 1932 1 1948 65
rect 2012 1 2028 65
rect 2092 61 2108 65
rect 2092 1 2108 5
rect 2172 1 2188 65
rect 2252 1 2268 65
rect 2332 61 2348 65
rect 2338 5 2348 61
rect 2332 1 2348 5
rect 2412 1 2428 65
rect 2492 61 2508 65
rect 2492 5 2506 61
rect 2492 1 2508 5
rect 2572 1 2588 65
rect 2652 1 2668 65
rect 2732 61 2748 65
rect 2732 1 2748 5
rect 2812 1 2828 65
rect 2892 1 2908 65
rect 2972 61 2988 65
rect 2972 1 2988 5
rect 3052 1 3068 65
rect 3132 1 3148 65
rect 3212 61 3228 65
rect 3212 1 3228 5
rect 3292 1 3308 65
rect 3372 1 3388 65
rect 3452 61 3468 65
rect 3458 5 3468 61
rect 3452 1 3468 5
rect 3532 1 3548 65
rect 3612 61 3628 65
rect 3612 5 3626 61
rect 3612 1 3628 5
rect 3692 1 3708 65
rect 3772 1 3788 65
rect 3852 61 3868 65
rect 3852 1 3868 5
rect 3932 1 3948 65
rect 4012 1 4028 65
rect 4092 61 4108 65
rect 4092 1 4108 5
rect 4172 1 4188 65
rect 4252 1 4268 65
rect 4332 61 4348 65
rect 4332 1 4348 5
rect 4412 1 4428 65
rect 4492 1 4508 65
rect 4572 61 4588 65
rect 4578 5 4588 61
rect 4572 1 4588 5
rect 4652 1 4668 65
rect 4732 61 4748 65
rect 4732 5 4746 61
rect 4732 1 4748 5
rect 4812 1 4828 65
rect 4892 1 4908 65
rect 4972 61 4988 65
rect 4972 1 4988 5
rect 5052 1 5068 65
rect 5132 1 5148 65
rect 5212 61 5228 65
rect 5212 1 5228 5
rect 5292 1 5308 65
rect 5372 1 5388 65
rect 5452 61 5468 65
rect 5452 1 5468 5
rect 5532 1 5548 65
rect 5612 1 5628 65
rect 5692 61 5708 65
rect 5698 5 5708 61
rect 5692 1 5708 5
rect 5772 1 5788 65
rect 5852 61 5868 65
rect 5852 5 5866 61
rect 5852 1 5868 5
rect 5932 1 5948 65
rect 6012 1 6028 65
rect 6092 61 6108 65
rect 6092 1 6108 5
rect 6172 1 6188 65
rect 6252 1 6268 65
rect 6332 61 6348 65
rect 6332 1 6348 5
rect 6412 1 6428 65
rect 6492 1 6508 65
rect 6572 61 6588 65
rect 6572 1 6588 5
rect 6652 1 6668 65
rect 6732 1 6748 65
rect 6812 61 6828 65
rect 6818 5 6828 61
rect 6812 1 6828 5
rect 6892 1 6908 65
rect 6972 61 6988 65
rect 6972 5 6986 61
rect 6972 1 6988 5
rect 7052 1 7068 65
rect 7132 1 7148 65
rect 7212 61 7228 65
rect 7212 1 7228 5
rect 7292 1 7308 65
rect 7372 1 7388 65
rect 7452 61 7468 65
rect 7452 1 7468 5
rect 7532 1 7548 65
rect 7612 1 7628 65
rect 7692 61 7708 65
rect 7692 1 7708 5
rect 7772 1 7788 65
rect 7852 1 7868 65
rect 7932 61 7948 65
rect 7938 5 7948 61
rect 7932 1 7948 5
rect 8012 1 8028 65
rect 8092 61 8108 65
rect 8092 5 8106 61
rect 8092 1 8108 5
rect 8172 1 8188 65
rect 8252 1 8268 65
rect 8332 61 8348 65
rect 8332 1 8348 5
rect 8412 1 8428 65
rect 8492 1 8508 65
rect 8572 61 8588 65
rect 8572 1 8588 5
rect 8652 1 8668 65
rect 8732 1 8748 65
rect 8812 61 8828 65
rect 8812 1 8828 5
rect 8892 1 8908 65
rect 8972 1 8988 65
rect 9052 61 9068 65
rect 9058 5 9068 61
rect 9052 1 9068 5
rect 9132 1 9148 65
rect 9212 61 9228 65
rect 9212 5 9226 61
rect 9212 1 9228 5
rect 9292 1 9308 65
rect 9372 1 9388 65
rect 9452 61 9468 65
rect 9452 1 9468 5
rect 9532 1 9548 65
rect 9612 1 9628 65
rect 9692 61 9708 65
rect 9692 1 9708 5
rect 9772 1 9788 65
rect 9852 1 9868 65
rect 9932 61 9948 65
rect 9932 1 9948 5
rect 10012 1 10028 65
rect 10092 1 10108 65
rect 10172 61 10188 65
rect 10178 5 10188 61
rect 10172 1 10188 5
rect 10252 1 10268 65
rect 10332 61 10348 65
rect 10332 5 10346 61
rect 10332 1 10348 5
rect 10412 1 10428 65
rect 10492 1 10508 65
rect 10572 61 10588 65
rect 10572 1 10588 5
rect 10652 1 10668 65
rect 10732 1 10748 65
rect 10812 61 10828 65
rect 10812 1 10828 5
rect 10892 1 10908 65
rect 10972 1 10988 65
rect 11052 61 11146 65
rect 11074 5 11146 61
rect 11052 1 11146 5
rect 0 0 11146 1
<< via3 >>
rect 28 4545 92 4609
rect 108 4605 172 4609
rect 108 4549 154 4605
rect 154 4549 172 4605
rect 108 4545 172 4549
rect 188 4545 252 4609
rect 268 4605 332 4609
rect 348 4605 412 4609
rect 268 4549 322 4605
rect 322 4549 332 4605
rect 348 4549 378 4605
rect 378 4549 412 4605
rect 268 4545 332 4549
rect 348 4545 412 4549
rect 428 4545 492 4609
rect 508 4605 572 4609
rect 588 4605 652 4609
rect 508 4549 546 4605
rect 546 4549 572 4605
rect 588 4549 602 4605
rect 602 4549 652 4605
rect 508 4545 572 4549
rect 588 4545 652 4549
rect 668 4545 732 4609
rect 748 4605 812 4609
rect 748 4549 770 4605
rect 770 4549 812 4605
rect 748 4545 812 4549
rect 828 4545 892 4609
rect 908 4545 972 4609
rect 988 4605 1052 4609
rect 988 4549 994 4605
rect 994 4549 1050 4605
rect 1050 4549 1052 4605
rect 988 4545 1052 4549
rect 1068 4545 1132 4609
rect 1148 4545 1212 4609
rect 1228 4605 1292 4609
rect 1228 4549 1274 4605
rect 1274 4549 1292 4605
rect 1228 4545 1292 4549
rect 1308 4545 1372 4609
rect 1388 4605 1452 4609
rect 1468 4605 1532 4609
rect 1388 4549 1442 4605
rect 1442 4549 1452 4605
rect 1468 4549 1498 4605
rect 1498 4549 1532 4605
rect 1388 4545 1452 4549
rect 1468 4545 1532 4549
rect 1548 4545 1612 4609
rect 1628 4605 1692 4609
rect 1708 4605 1772 4609
rect 1628 4549 1666 4605
rect 1666 4549 1692 4605
rect 1708 4549 1722 4605
rect 1722 4549 1772 4605
rect 1628 4545 1692 4549
rect 1708 4545 1772 4549
rect 1788 4545 1852 4609
rect 1868 4605 1932 4609
rect 1868 4549 1890 4605
rect 1890 4549 1932 4605
rect 1868 4545 1932 4549
rect 1948 4545 2012 4609
rect 2028 4545 2092 4609
rect 2108 4605 2172 4609
rect 2108 4549 2114 4605
rect 2114 4549 2170 4605
rect 2170 4549 2172 4605
rect 2108 4545 2172 4549
rect 2188 4545 2252 4609
rect 2268 4545 2332 4609
rect 2348 4605 2412 4609
rect 2348 4549 2394 4605
rect 2394 4549 2412 4605
rect 2348 4545 2412 4549
rect 2428 4545 2492 4609
rect 2508 4605 2572 4609
rect 2588 4605 2652 4609
rect 2508 4549 2562 4605
rect 2562 4549 2572 4605
rect 2588 4549 2618 4605
rect 2618 4549 2652 4605
rect 2508 4545 2572 4549
rect 2588 4545 2652 4549
rect 2668 4545 2732 4609
rect 2748 4605 2812 4609
rect 2828 4605 2892 4609
rect 2748 4549 2786 4605
rect 2786 4549 2812 4605
rect 2828 4549 2842 4605
rect 2842 4549 2892 4605
rect 2748 4545 2812 4549
rect 2828 4545 2892 4549
rect 2908 4545 2972 4609
rect 2988 4605 3052 4609
rect 2988 4549 3010 4605
rect 3010 4549 3052 4605
rect 2988 4545 3052 4549
rect 3068 4545 3132 4609
rect 3148 4545 3212 4609
rect 3228 4605 3292 4609
rect 3228 4549 3234 4605
rect 3234 4549 3290 4605
rect 3290 4549 3292 4605
rect 3228 4545 3292 4549
rect 3308 4545 3372 4609
rect 3388 4545 3452 4609
rect 3468 4605 3532 4609
rect 3468 4549 3514 4605
rect 3514 4549 3532 4605
rect 3468 4545 3532 4549
rect 3548 4545 3612 4609
rect 3628 4605 3692 4609
rect 3708 4605 3772 4609
rect 3628 4549 3682 4605
rect 3682 4549 3692 4605
rect 3708 4549 3738 4605
rect 3738 4549 3772 4605
rect 3628 4545 3692 4549
rect 3708 4545 3772 4549
rect 3788 4545 3852 4609
rect 3868 4605 3932 4609
rect 3948 4605 4012 4609
rect 3868 4549 3906 4605
rect 3906 4549 3932 4605
rect 3948 4549 3962 4605
rect 3962 4549 4012 4605
rect 3868 4545 3932 4549
rect 3948 4545 4012 4549
rect 4028 4545 4092 4609
rect 4108 4605 4172 4609
rect 4108 4549 4130 4605
rect 4130 4549 4172 4605
rect 4108 4545 4172 4549
rect 4188 4545 4252 4609
rect 4268 4545 4332 4609
rect 4348 4605 4412 4609
rect 4348 4549 4354 4605
rect 4354 4549 4410 4605
rect 4410 4549 4412 4605
rect 4348 4545 4412 4549
rect 4428 4545 4492 4609
rect 4508 4545 4572 4609
rect 4588 4605 4652 4609
rect 4588 4549 4634 4605
rect 4634 4549 4652 4605
rect 4588 4545 4652 4549
rect 4668 4545 4732 4609
rect 4748 4605 4812 4609
rect 4828 4605 4892 4609
rect 4748 4549 4802 4605
rect 4802 4549 4812 4605
rect 4828 4549 4858 4605
rect 4858 4549 4892 4605
rect 4748 4545 4812 4549
rect 4828 4545 4892 4549
rect 4908 4545 4972 4609
rect 4988 4605 5052 4609
rect 5068 4605 5132 4609
rect 4988 4549 5026 4605
rect 5026 4549 5052 4605
rect 5068 4549 5082 4605
rect 5082 4549 5132 4605
rect 4988 4545 5052 4549
rect 5068 4545 5132 4549
rect 5148 4545 5212 4609
rect 5228 4605 5292 4609
rect 5228 4549 5250 4605
rect 5250 4549 5292 4605
rect 5228 4545 5292 4549
rect 5308 4545 5372 4609
rect 5388 4545 5452 4609
rect 5468 4605 5532 4609
rect 5468 4549 5474 4605
rect 5474 4549 5530 4605
rect 5530 4549 5532 4605
rect 5468 4545 5532 4549
rect 5548 4545 5612 4609
rect 5628 4545 5692 4609
rect 5708 4605 5772 4609
rect 5708 4549 5754 4605
rect 5754 4549 5772 4605
rect 5708 4545 5772 4549
rect 5788 4545 5852 4609
rect 5868 4605 5932 4609
rect 5948 4605 6012 4609
rect 5868 4549 5922 4605
rect 5922 4549 5932 4605
rect 5948 4549 5978 4605
rect 5978 4549 6012 4605
rect 5868 4545 5932 4549
rect 5948 4545 6012 4549
rect 6028 4545 6092 4609
rect 6108 4605 6172 4609
rect 6188 4605 6252 4609
rect 6108 4549 6146 4605
rect 6146 4549 6172 4605
rect 6188 4549 6202 4605
rect 6202 4549 6252 4605
rect 6108 4545 6172 4549
rect 6188 4545 6252 4549
rect 6268 4545 6332 4609
rect 6348 4605 6412 4609
rect 6348 4549 6370 4605
rect 6370 4549 6412 4605
rect 6348 4545 6412 4549
rect 6428 4545 6492 4609
rect 6508 4545 6572 4609
rect 6588 4605 6652 4609
rect 6588 4549 6594 4605
rect 6594 4549 6650 4605
rect 6650 4549 6652 4605
rect 6588 4545 6652 4549
rect 6668 4545 6732 4609
rect 6748 4545 6812 4609
rect 6828 4605 6892 4609
rect 6828 4549 6874 4605
rect 6874 4549 6892 4605
rect 6828 4545 6892 4549
rect 6908 4545 6972 4609
rect 6988 4605 7052 4609
rect 7068 4605 7132 4609
rect 6988 4549 7042 4605
rect 7042 4549 7052 4605
rect 7068 4549 7098 4605
rect 7098 4549 7132 4605
rect 6988 4545 7052 4549
rect 7068 4545 7132 4549
rect 7148 4545 7212 4609
rect 7228 4605 7292 4609
rect 7308 4605 7372 4609
rect 7228 4549 7266 4605
rect 7266 4549 7292 4605
rect 7308 4549 7322 4605
rect 7322 4549 7372 4605
rect 7228 4545 7292 4549
rect 7308 4545 7372 4549
rect 7388 4545 7452 4609
rect 7468 4605 7532 4609
rect 7468 4549 7490 4605
rect 7490 4549 7532 4605
rect 7468 4545 7532 4549
rect 7548 4545 7612 4609
rect 7628 4545 7692 4609
rect 7708 4605 7772 4609
rect 7708 4549 7714 4605
rect 7714 4549 7770 4605
rect 7770 4549 7772 4605
rect 7708 4545 7772 4549
rect 7788 4545 7852 4609
rect 7868 4545 7932 4609
rect 7948 4605 8012 4609
rect 7948 4549 7994 4605
rect 7994 4549 8012 4605
rect 7948 4545 8012 4549
rect 8028 4545 8092 4609
rect 8108 4605 8172 4609
rect 8188 4605 8252 4609
rect 8108 4549 8162 4605
rect 8162 4549 8172 4605
rect 8188 4549 8218 4605
rect 8218 4549 8252 4605
rect 8108 4545 8172 4549
rect 8188 4545 8252 4549
rect 8268 4545 8332 4609
rect 8348 4605 8412 4609
rect 8428 4605 8492 4609
rect 8348 4549 8386 4605
rect 8386 4549 8412 4605
rect 8428 4549 8442 4605
rect 8442 4549 8492 4605
rect 8348 4545 8412 4549
rect 8428 4545 8492 4549
rect 8508 4545 8572 4609
rect 8588 4605 8652 4609
rect 8588 4549 8610 4605
rect 8610 4549 8652 4605
rect 8588 4545 8652 4549
rect 8668 4545 8732 4609
rect 8748 4545 8812 4609
rect 8828 4605 8892 4609
rect 8828 4549 8834 4605
rect 8834 4549 8890 4605
rect 8890 4549 8892 4605
rect 8828 4545 8892 4549
rect 8908 4545 8972 4609
rect 8988 4545 9052 4609
rect 9068 4605 9132 4609
rect 9068 4549 9114 4605
rect 9114 4549 9132 4605
rect 9068 4545 9132 4549
rect 9148 4545 9212 4609
rect 9228 4605 9292 4609
rect 9308 4605 9372 4609
rect 9228 4549 9282 4605
rect 9282 4549 9292 4605
rect 9308 4549 9338 4605
rect 9338 4549 9372 4605
rect 9228 4545 9292 4549
rect 9308 4545 9372 4549
rect 9388 4545 9452 4609
rect 9468 4605 9532 4609
rect 9548 4605 9612 4609
rect 9468 4549 9506 4605
rect 9506 4549 9532 4605
rect 9548 4549 9562 4605
rect 9562 4549 9612 4605
rect 9468 4545 9532 4549
rect 9548 4545 9612 4549
rect 9628 4545 9692 4609
rect 9708 4605 9772 4609
rect 9708 4549 9730 4605
rect 9730 4549 9772 4605
rect 9708 4545 9772 4549
rect 9788 4545 9852 4609
rect 9868 4545 9932 4609
rect 9948 4605 10012 4609
rect 9948 4549 9954 4605
rect 9954 4549 10010 4605
rect 10010 4549 10012 4605
rect 9948 4545 10012 4549
rect 10028 4545 10092 4609
rect 10108 4545 10172 4609
rect 10188 4605 10252 4609
rect 10188 4549 10234 4605
rect 10234 4549 10252 4605
rect 10188 4545 10252 4549
rect 10268 4545 10332 4609
rect 10348 4605 10412 4609
rect 10428 4605 10492 4609
rect 10348 4549 10402 4605
rect 10402 4549 10412 4605
rect 10428 4549 10458 4605
rect 10458 4549 10492 4605
rect 10348 4545 10412 4549
rect 10428 4545 10492 4549
rect 10508 4545 10572 4609
rect 10588 4605 10652 4609
rect 10668 4605 10732 4609
rect 10588 4549 10626 4605
rect 10626 4549 10652 4605
rect 10668 4549 10682 4605
rect 10682 4549 10732 4605
rect 10588 4545 10652 4549
rect 10668 4545 10732 4549
rect 10748 4545 10812 4609
rect 10828 4605 10892 4609
rect 10828 4549 10850 4605
rect 10850 4549 10892 4605
rect 10828 4545 10892 4549
rect 10908 4545 10972 4609
rect 10988 4545 11052 4609
rect 28 61 92 65
rect 28 5 42 61
rect 42 5 92 61
rect 28 1 92 5
rect 108 1 172 65
rect 188 1 252 65
rect 268 61 332 65
rect 268 5 322 61
rect 322 5 332 61
rect 268 1 332 5
rect 348 1 412 65
rect 428 61 492 65
rect 508 61 572 65
rect 428 5 490 61
rect 490 5 492 61
rect 508 5 546 61
rect 546 5 572 61
rect 428 1 492 5
rect 508 1 572 5
rect 588 1 652 65
rect 668 61 732 65
rect 748 61 812 65
rect 668 5 714 61
rect 714 5 732 61
rect 748 5 770 61
rect 770 5 812 61
rect 668 1 732 5
rect 748 1 812 5
rect 828 1 892 65
rect 908 61 972 65
rect 988 61 1052 65
rect 908 5 938 61
rect 938 5 972 61
rect 988 5 994 61
rect 994 5 1052 61
rect 908 1 972 5
rect 988 1 1052 5
rect 1068 1 1132 65
rect 1148 61 1212 65
rect 1148 5 1162 61
rect 1162 5 1212 61
rect 1148 1 1212 5
rect 1228 1 1292 65
rect 1308 1 1372 65
rect 1388 61 1452 65
rect 1388 5 1442 61
rect 1442 5 1452 61
rect 1388 1 1452 5
rect 1468 1 1532 65
rect 1548 61 1612 65
rect 1628 61 1692 65
rect 1548 5 1610 61
rect 1610 5 1612 61
rect 1628 5 1666 61
rect 1666 5 1692 61
rect 1548 1 1612 5
rect 1628 1 1692 5
rect 1708 1 1772 65
rect 1788 61 1852 65
rect 1868 61 1932 65
rect 1788 5 1834 61
rect 1834 5 1852 61
rect 1868 5 1890 61
rect 1890 5 1932 61
rect 1788 1 1852 5
rect 1868 1 1932 5
rect 1948 1 2012 65
rect 2028 61 2092 65
rect 2108 61 2172 65
rect 2028 5 2058 61
rect 2058 5 2092 61
rect 2108 5 2114 61
rect 2114 5 2172 61
rect 2028 1 2092 5
rect 2108 1 2172 5
rect 2188 1 2252 65
rect 2268 61 2332 65
rect 2268 5 2282 61
rect 2282 5 2332 61
rect 2268 1 2332 5
rect 2348 1 2412 65
rect 2428 1 2492 65
rect 2508 61 2572 65
rect 2508 5 2562 61
rect 2562 5 2572 61
rect 2508 1 2572 5
rect 2588 1 2652 65
rect 2668 61 2732 65
rect 2748 61 2812 65
rect 2668 5 2730 61
rect 2730 5 2732 61
rect 2748 5 2786 61
rect 2786 5 2812 61
rect 2668 1 2732 5
rect 2748 1 2812 5
rect 2828 1 2892 65
rect 2908 61 2972 65
rect 2988 61 3052 65
rect 2908 5 2954 61
rect 2954 5 2972 61
rect 2988 5 3010 61
rect 3010 5 3052 61
rect 2908 1 2972 5
rect 2988 1 3052 5
rect 3068 1 3132 65
rect 3148 61 3212 65
rect 3228 61 3292 65
rect 3148 5 3178 61
rect 3178 5 3212 61
rect 3228 5 3234 61
rect 3234 5 3292 61
rect 3148 1 3212 5
rect 3228 1 3292 5
rect 3308 1 3372 65
rect 3388 61 3452 65
rect 3388 5 3402 61
rect 3402 5 3452 61
rect 3388 1 3452 5
rect 3468 1 3532 65
rect 3548 1 3612 65
rect 3628 61 3692 65
rect 3628 5 3682 61
rect 3682 5 3692 61
rect 3628 1 3692 5
rect 3708 1 3772 65
rect 3788 61 3852 65
rect 3868 61 3932 65
rect 3788 5 3850 61
rect 3850 5 3852 61
rect 3868 5 3906 61
rect 3906 5 3932 61
rect 3788 1 3852 5
rect 3868 1 3932 5
rect 3948 1 4012 65
rect 4028 61 4092 65
rect 4108 61 4172 65
rect 4028 5 4074 61
rect 4074 5 4092 61
rect 4108 5 4130 61
rect 4130 5 4172 61
rect 4028 1 4092 5
rect 4108 1 4172 5
rect 4188 1 4252 65
rect 4268 61 4332 65
rect 4348 61 4412 65
rect 4268 5 4298 61
rect 4298 5 4332 61
rect 4348 5 4354 61
rect 4354 5 4412 61
rect 4268 1 4332 5
rect 4348 1 4412 5
rect 4428 1 4492 65
rect 4508 61 4572 65
rect 4508 5 4522 61
rect 4522 5 4572 61
rect 4508 1 4572 5
rect 4588 1 4652 65
rect 4668 1 4732 65
rect 4748 61 4812 65
rect 4748 5 4802 61
rect 4802 5 4812 61
rect 4748 1 4812 5
rect 4828 1 4892 65
rect 4908 61 4972 65
rect 4988 61 5052 65
rect 4908 5 4970 61
rect 4970 5 4972 61
rect 4988 5 5026 61
rect 5026 5 5052 61
rect 4908 1 4972 5
rect 4988 1 5052 5
rect 5068 1 5132 65
rect 5148 61 5212 65
rect 5228 61 5292 65
rect 5148 5 5194 61
rect 5194 5 5212 61
rect 5228 5 5250 61
rect 5250 5 5292 61
rect 5148 1 5212 5
rect 5228 1 5292 5
rect 5308 1 5372 65
rect 5388 61 5452 65
rect 5468 61 5532 65
rect 5388 5 5418 61
rect 5418 5 5452 61
rect 5468 5 5474 61
rect 5474 5 5532 61
rect 5388 1 5452 5
rect 5468 1 5532 5
rect 5548 1 5612 65
rect 5628 61 5692 65
rect 5628 5 5642 61
rect 5642 5 5692 61
rect 5628 1 5692 5
rect 5708 1 5772 65
rect 5788 1 5852 65
rect 5868 61 5932 65
rect 5868 5 5922 61
rect 5922 5 5932 61
rect 5868 1 5932 5
rect 5948 1 6012 65
rect 6028 61 6092 65
rect 6108 61 6172 65
rect 6028 5 6090 61
rect 6090 5 6092 61
rect 6108 5 6146 61
rect 6146 5 6172 61
rect 6028 1 6092 5
rect 6108 1 6172 5
rect 6188 1 6252 65
rect 6268 61 6332 65
rect 6348 61 6412 65
rect 6268 5 6314 61
rect 6314 5 6332 61
rect 6348 5 6370 61
rect 6370 5 6412 61
rect 6268 1 6332 5
rect 6348 1 6412 5
rect 6428 1 6492 65
rect 6508 61 6572 65
rect 6588 61 6652 65
rect 6508 5 6538 61
rect 6538 5 6572 61
rect 6588 5 6594 61
rect 6594 5 6652 61
rect 6508 1 6572 5
rect 6588 1 6652 5
rect 6668 1 6732 65
rect 6748 61 6812 65
rect 6748 5 6762 61
rect 6762 5 6812 61
rect 6748 1 6812 5
rect 6828 1 6892 65
rect 6908 1 6972 65
rect 6988 61 7052 65
rect 6988 5 7042 61
rect 7042 5 7052 61
rect 6988 1 7052 5
rect 7068 1 7132 65
rect 7148 61 7212 65
rect 7228 61 7292 65
rect 7148 5 7210 61
rect 7210 5 7212 61
rect 7228 5 7266 61
rect 7266 5 7292 61
rect 7148 1 7212 5
rect 7228 1 7292 5
rect 7308 1 7372 65
rect 7388 61 7452 65
rect 7468 61 7532 65
rect 7388 5 7434 61
rect 7434 5 7452 61
rect 7468 5 7490 61
rect 7490 5 7532 61
rect 7388 1 7452 5
rect 7468 1 7532 5
rect 7548 1 7612 65
rect 7628 61 7692 65
rect 7708 61 7772 65
rect 7628 5 7658 61
rect 7658 5 7692 61
rect 7708 5 7714 61
rect 7714 5 7772 61
rect 7628 1 7692 5
rect 7708 1 7772 5
rect 7788 1 7852 65
rect 7868 61 7932 65
rect 7868 5 7882 61
rect 7882 5 7932 61
rect 7868 1 7932 5
rect 7948 1 8012 65
rect 8028 1 8092 65
rect 8108 61 8172 65
rect 8108 5 8162 61
rect 8162 5 8172 61
rect 8108 1 8172 5
rect 8188 1 8252 65
rect 8268 61 8332 65
rect 8348 61 8412 65
rect 8268 5 8330 61
rect 8330 5 8332 61
rect 8348 5 8386 61
rect 8386 5 8412 61
rect 8268 1 8332 5
rect 8348 1 8412 5
rect 8428 1 8492 65
rect 8508 61 8572 65
rect 8588 61 8652 65
rect 8508 5 8554 61
rect 8554 5 8572 61
rect 8588 5 8610 61
rect 8610 5 8652 61
rect 8508 1 8572 5
rect 8588 1 8652 5
rect 8668 1 8732 65
rect 8748 61 8812 65
rect 8828 61 8892 65
rect 8748 5 8778 61
rect 8778 5 8812 61
rect 8828 5 8834 61
rect 8834 5 8892 61
rect 8748 1 8812 5
rect 8828 1 8892 5
rect 8908 1 8972 65
rect 8988 61 9052 65
rect 8988 5 9002 61
rect 9002 5 9052 61
rect 8988 1 9052 5
rect 9068 1 9132 65
rect 9148 1 9212 65
rect 9228 61 9292 65
rect 9228 5 9282 61
rect 9282 5 9292 61
rect 9228 1 9292 5
rect 9308 1 9372 65
rect 9388 61 9452 65
rect 9468 61 9532 65
rect 9388 5 9450 61
rect 9450 5 9452 61
rect 9468 5 9506 61
rect 9506 5 9532 61
rect 9388 1 9452 5
rect 9468 1 9532 5
rect 9548 1 9612 65
rect 9628 61 9692 65
rect 9708 61 9772 65
rect 9628 5 9674 61
rect 9674 5 9692 61
rect 9708 5 9730 61
rect 9730 5 9772 61
rect 9628 1 9692 5
rect 9708 1 9772 5
rect 9788 1 9852 65
rect 9868 61 9932 65
rect 9948 61 10012 65
rect 9868 5 9898 61
rect 9898 5 9932 61
rect 9948 5 9954 61
rect 9954 5 10012 61
rect 9868 1 9932 5
rect 9948 1 10012 5
rect 10028 1 10092 65
rect 10108 61 10172 65
rect 10108 5 10122 61
rect 10122 5 10172 61
rect 10108 1 10172 5
rect 10188 1 10252 65
rect 10268 1 10332 65
rect 10348 61 10412 65
rect 10348 5 10402 61
rect 10402 5 10412 61
rect 10348 1 10412 5
rect 10428 1 10492 65
rect 10508 61 10572 65
rect 10588 61 10652 65
rect 10508 5 10570 61
rect 10570 5 10572 61
rect 10588 5 10626 61
rect 10626 5 10652 61
rect 10508 1 10572 5
rect 10588 1 10652 5
rect 10668 1 10732 65
rect 10748 61 10812 65
rect 10828 61 10892 65
rect 10748 5 10794 61
rect 10794 5 10812 61
rect 10828 5 10850 61
rect 10850 5 10892 61
rect 10748 1 10812 5
rect 10828 1 10892 5
rect 10908 1 10972 65
rect 10988 61 11052 65
rect 10988 5 11018 61
rect 11018 5 11052 61
rect 10988 1 11052 5
<< metal4 >>
rect 0 4609 11146 4610
rect 0 4545 28 4609
rect 92 4545 108 4609
rect 172 4545 188 4609
rect 252 4545 268 4609
rect 332 4545 348 4609
rect 412 4545 428 4609
rect 492 4545 508 4609
rect 572 4545 588 4609
rect 652 4545 668 4609
rect 732 4545 748 4609
rect 812 4545 828 4609
rect 892 4545 908 4609
rect 972 4545 988 4609
rect 1052 4545 1068 4609
rect 1132 4545 1148 4609
rect 1212 4545 1228 4609
rect 1292 4545 1308 4609
rect 1372 4545 1388 4609
rect 1452 4545 1468 4609
rect 1532 4545 1548 4609
rect 1612 4545 1628 4609
rect 1692 4545 1708 4609
rect 1772 4545 1788 4609
rect 1852 4545 1868 4609
rect 1932 4545 1948 4609
rect 2012 4545 2028 4609
rect 2092 4545 2108 4609
rect 2172 4545 2188 4609
rect 2252 4545 2268 4609
rect 2332 4545 2348 4609
rect 2412 4545 2428 4609
rect 2492 4545 2508 4609
rect 2572 4545 2588 4609
rect 2652 4545 2668 4609
rect 2732 4545 2748 4609
rect 2812 4545 2828 4609
rect 2892 4545 2908 4609
rect 2972 4545 2988 4609
rect 3052 4545 3068 4609
rect 3132 4545 3148 4609
rect 3212 4545 3228 4609
rect 3292 4545 3308 4609
rect 3372 4545 3388 4609
rect 3452 4545 3468 4609
rect 3532 4545 3548 4609
rect 3612 4545 3628 4609
rect 3692 4545 3708 4609
rect 3772 4545 3788 4609
rect 3852 4545 3868 4609
rect 3932 4545 3948 4609
rect 4012 4545 4028 4609
rect 4092 4545 4108 4609
rect 4172 4545 4188 4609
rect 4252 4545 4268 4609
rect 4332 4545 4348 4609
rect 4412 4545 4428 4609
rect 4492 4545 4508 4609
rect 4572 4545 4588 4609
rect 4652 4545 4668 4609
rect 4732 4545 4748 4609
rect 4812 4545 4828 4609
rect 4892 4545 4908 4609
rect 4972 4545 4988 4609
rect 5052 4545 5068 4609
rect 5132 4545 5148 4609
rect 5212 4545 5228 4609
rect 5292 4545 5308 4609
rect 5372 4545 5388 4609
rect 5452 4545 5468 4609
rect 5532 4545 5548 4609
rect 5612 4545 5628 4609
rect 5692 4545 5708 4609
rect 5772 4545 5788 4609
rect 5852 4545 5868 4609
rect 5932 4545 5948 4609
rect 6012 4545 6028 4609
rect 6092 4545 6108 4609
rect 6172 4545 6188 4609
rect 6252 4545 6268 4609
rect 6332 4545 6348 4609
rect 6412 4545 6428 4609
rect 6492 4545 6508 4609
rect 6572 4545 6588 4609
rect 6652 4545 6668 4609
rect 6732 4545 6748 4609
rect 6812 4545 6828 4609
rect 6892 4545 6908 4609
rect 6972 4545 6988 4609
rect 7052 4545 7068 4609
rect 7132 4545 7148 4609
rect 7212 4545 7228 4609
rect 7292 4545 7308 4609
rect 7372 4545 7388 4609
rect 7452 4545 7468 4609
rect 7532 4545 7548 4609
rect 7612 4545 7628 4609
rect 7692 4545 7708 4609
rect 7772 4545 7788 4609
rect 7852 4545 7868 4609
rect 7932 4545 7948 4609
rect 8012 4545 8028 4609
rect 8092 4545 8108 4609
rect 8172 4545 8188 4609
rect 8252 4545 8268 4609
rect 8332 4545 8348 4609
rect 8412 4545 8428 4609
rect 8492 4545 8508 4609
rect 8572 4545 8588 4609
rect 8652 4545 8668 4609
rect 8732 4545 8748 4609
rect 8812 4545 8828 4609
rect 8892 4545 8908 4609
rect 8972 4545 8988 4609
rect 9052 4545 9068 4609
rect 9132 4545 9148 4609
rect 9212 4545 9228 4609
rect 9292 4545 9308 4609
rect 9372 4545 9388 4609
rect 9452 4545 9468 4609
rect 9532 4545 9548 4609
rect 9612 4545 9628 4609
rect 9692 4545 9708 4609
rect 9772 4545 9788 4609
rect 9852 4545 9868 4609
rect 9932 4545 9948 4609
rect 10012 4545 10028 4609
rect 10092 4545 10108 4609
rect 10172 4545 10188 4609
rect 10252 4545 10268 4609
rect 10332 4545 10348 4609
rect 10412 4545 10428 4609
rect 10492 4545 10508 4609
rect 10572 4545 10588 4609
rect 10652 4545 10668 4609
rect 10732 4545 10748 4609
rect 10812 4545 10828 4609
rect 10892 4545 10908 4609
rect 10972 4545 10988 4609
rect 11052 4545 11146 4609
rect 0 4544 11146 4545
rect 120 4535 420 4544
rect 0 66 60 4484
rect 120 4299 152 4535
rect 388 4299 420 4535
rect 120 126 180 4299
rect 240 311 300 4239
rect 360 371 420 4299
rect 480 311 540 4484
rect 240 75 272 311
rect 508 75 540 311
rect 600 126 660 4544
rect 240 66 540 75
rect 720 66 780 4484
rect 840 126 900 4544
rect 960 66 1020 4484
rect 1080 126 1140 4544
rect 1200 66 1260 4484
rect 1320 126 1380 4544
rect 1560 4535 1860 4544
rect 1440 66 1500 4484
rect 1560 4299 1592 4535
rect 1828 4299 1860 4535
rect 1560 126 1620 4299
rect 1680 311 1740 4239
rect 1800 371 1860 4299
rect 1920 311 1980 4484
rect 1680 75 1712 311
rect 1948 75 1980 311
rect 2040 126 2100 4544
rect 1680 66 1980 75
rect 2160 66 2220 4484
rect 2280 126 2340 4544
rect 2400 66 2460 4484
rect 2520 126 2580 4544
rect 2640 66 2700 4484
rect 2760 126 2820 4544
rect 3000 4535 3300 4544
rect 2880 66 2940 4484
rect 3000 4299 3032 4535
rect 3268 4299 3300 4535
rect 3000 126 3060 4299
rect 3120 311 3180 4239
rect 3240 371 3300 4299
rect 3360 311 3420 4484
rect 3120 75 3152 311
rect 3388 75 3420 311
rect 3480 126 3540 4544
rect 3120 66 3420 75
rect 3600 66 3660 4484
rect 3720 126 3780 4544
rect 3840 66 3900 4484
rect 3960 126 4020 4544
rect 4080 66 4140 4484
rect 4200 126 4260 4544
rect 4440 4535 4740 4544
rect 4320 66 4380 4484
rect 4440 4299 4472 4535
rect 4708 4299 4740 4535
rect 4440 126 4500 4299
rect 4560 311 4620 4239
rect 4680 371 4740 4299
rect 4800 311 4860 4484
rect 4560 75 4592 311
rect 4828 75 4860 311
rect 4920 126 4980 4544
rect 4560 66 4860 75
rect 5040 66 5100 4484
rect 5160 126 5220 4544
rect 5280 66 5340 4484
rect 5400 126 5460 4544
rect 5520 66 5580 4484
rect 5640 126 5700 4544
rect 5880 4535 6180 4544
rect 5760 66 5820 4484
rect 5880 4299 5912 4535
rect 6148 4299 6180 4535
rect 5880 126 5940 4299
rect 6000 311 6060 4239
rect 6120 371 6180 4299
rect 6240 311 6300 4484
rect 6000 75 6032 311
rect 6268 75 6300 311
rect 6360 126 6420 4544
rect 6000 66 6300 75
rect 6480 66 6540 4484
rect 6600 126 6660 4544
rect 6720 66 6780 4484
rect 6840 126 6900 4544
rect 6960 66 7020 4484
rect 7080 126 7140 4544
rect 7320 4535 7620 4544
rect 7200 66 7260 4484
rect 7320 4299 7352 4535
rect 7588 4299 7620 4535
rect 7320 126 7380 4299
rect 7440 311 7500 4239
rect 7560 371 7620 4299
rect 7680 311 7740 4484
rect 7440 75 7472 311
rect 7708 75 7740 311
rect 7800 126 7860 4544
rect 7440 66 7740 75
rect 7920 66 7980 4484
rect 8040 126 8100 4544
rect 8160 66 8220 4484
rect 8280 126 8340 4544
rect 8400 66 8460 4484
rect 8520 126 8580 4544
rect 8760 4535 9060 4544
rect 8640 66 8700 4484
rect 8760 4299 8792 4535
rect 9028 4299 9060 4535
rect 8760 126 8820 4299
rect 8880 311 8940 4239
rect 9000 371 9060 4299
rect 9120 311 9180 4484
rect 8880 75 8912 311
rect 9148 75 9180 311
rect 9240 126 9300 4544
rect 8880 66 9180 75
rect 9360 66 9420 4484
rect 9480 126 9540 4544
rect 9600 66 9660 4484
rect 9720 126 9780 4544
rect 9840 66 9900 4484
rect 9960 126 10020 4544
rect 10200 4535 10500 4544
rect 10080 66 10140 4484
rect 10200 4299 10232 4535
rect 10468 4299 10500 4535
rect 10200 126 10260 4299
rect 10320 311 10380 4239
rect 10440 371 10500 4299
rect 10560 311 10620 4484
rect 10320 75 10352 311
rect 10588 75 10620 311
rect 10680 126 10740 4544
rect 10320 66 10620 75
rect 10800 66 10860 4484
rect 10920 126 10980 4544
rect 11040 66 11146 4484
rect 0 65 11146 66
rect 0 1 28 65
rect 92 1 108 65
rect 172 1 188 65
rect 252 1 268 65
rect 332 1 348 65
rect 412 1 428 65
rect 492 1 508 65
rect 572 1 588 65
rect 652 1 668 65
rect 732 1 748 65
rect 812 1 828 65
rect 892 1 908 65
rect 972 1 988 65
rect 1052 1 1068 65
rect 1132 1 1148 65
rect 1212 1 1228 65
rect 1292 1 1308 65
rect 1372 1 1388 65
rect 1452 1 1468 65
rect 1532 1 1548 65
rect 1612 1 1628 65
rect 1692 1 1708 65
rect 1772 1 1788 65
rect 1852 1 1868 65
rect 1932 1 1948 65
rect 2012 1 2028 65
rect 2092 1 2108 65
rect 2172 1 2188 65
rect 2252 1 2268 65
rect 2332 1 2348 65
rect 2412 1 2428 65
rect 2492 1 2508 65
rect 2572 1 2588 65
rect 2652 1 2668 65
rect 2732 1 2748 65
rect 2812 1 2828 65
rect 2892 1 2908 65
rect 2972 1 2988 65
rect 3052 1 3068 65
rect 3132 1 3148 65
rect 3212 1 3228 65
rect 3292 1 3308 65
rect 3372 1 3388 65
rect 3452 1 3468 65
rect 3532 1 3548 65
rect 3612 1 3628 65
rect 3692 1 3708 65
rect 3772 1 3788 65
rect 3852 1 3868 65
rect 3932 1 3948 65
rect 4012 1 4028 65
rect 4092 1 4108 65
rect 4172 1 4188 65
rect 4252 1 4268 65
rect 4332 1 4348 65
rect 4412 1 4428 65
rect 4492 1 4508 65
rect 4572 1 4588 65
rect 4652 1 4668 65
rect 4732 1 4748 65
rect 4812 1 4828 65
rect 4892 1 4908 65
rect 4972 1 4988 65
rect 5052 1 5068 65
rect 5132 1 5148 65
rect 5212 1 5228 65
rect 5292 1 5308 65
rect 5372 1 5388 65
rect 5452 1 5468 65
rect 5532 1 5548 65
rect 5612 1 5628 65
rect 5692 1 5708 65
rect 5772 1 5788 65
rect 5852 1 5868 65
rect 5932 1 5948 65
rect 6012 1 6028 65
rect 6092 1 6108 65
rect 6172 1 6188 65
rect 6252 1 6268 65
rect 6332 1 6348 65
rect 6412 1 6428 65
rect 6492 1 6508 65
rect 6572 1 6588 65
rect 6652 1 6668 65
rect 6732 1 6748 65
rect 6812 1 6828 65
rect 6892 1 6908 65
rect 6972 1 6988 65
rect 7052 1 7068 65
rect 7132 1 7148 65
rect 7212 1 7228 65
rect 7292 1 7308 65
rect 7372 1 7388 65
rect 7452 1 7468 65
rect 7532 1 7548 65
rect 7612 1 7628 65
rect 7692 1 7708 65
rect 7772 1 7788 65
rect 7852 1 7868 65
rect 7932 1 7948 65
rect 8012 1 8028 65
rect 8092 1 8108 65
rect 8172 1 8188 65
rect 8252 1 8268 65
rect 8332 1 8348 65
rect 8412 1 8428 65
rect 8492 1 8508 65
rect 8572 1 8588 65
rect 8652 1 8668 65
rect 8732 1 8748 65
rect 8812 1 8828 65
rect 8892 1 8908 65
rect 8972 1 8988 65
rect 9052 1 9068 65
rect 9132 1 9148 65
rect 9212 1 9228 65
rect 9292 1 9308 65
rect 9372 1 9388 65
rect 9452 1 9468 65
rect 9532 1 9548 65
rect 9612 1 9628 65
rect 9692 1 9708 65
rect 9772 1 9788 65
rect 9852 1 9868 65
rect 9932 1 9948 65
rect 10012 1 10028 65
rect 10092 1 10108 65
rect 10172 1 10188 65
rect 10252 1 10268 65
rect 10332 1 10348 65
rect 10412 1 10428 65
rect 10492 1 10508 65
rect 10572 1 10588 65
rect 10652 1 10668 65
rect 10732 1 10748 65
rect 10812 1 10828 65
rect 10892 1 10908 65
rect 10972 1 10988 65
rect 11052 1 11146 65
rect 0 0 11146 1
<< via4 >>
rect 152 4299 388 4535
rect 272 75 508 311
rect 1592 4299 1828 4535
rect 1712 75 1948 311
rect 3032 4299 3268 4535
rect 3152 75 3388 311
rect 4472 4299 4708 4535
rect 4592 75 4828 311
rect 5912 4299 6148 4535
rect 6032 75 6268 311
rect 7352 4299 7588 4535
rect 7472 75 7708 311
rect 8792 4299 9028 4535
rect 8912 75 9148 311
rect 10232 4299 10468 4535
rect 10352 75 10588 311
<< metal5 >>
rect 0 4535 11146 4610
rect 0 4299 152 4535
rect 388 4299 1592 4535
rect 1828 4299 3032 4535
rect 3268 4299 4472 4535
rect 4708 4299 5912 4535
rect 6148 4299 7352 4535
rect 7588 4299 8792 4535
rect 9028 4299 10232 4535
rect 10468 4299 11146 4535
rect 0 4275 11146 4299
rect 0 655 320 4275
rect 640 335 960 3955
rect 1280 655 1600 4275
rect 1920 335 2240 3955
rect 2560 655 2880 4275
rect 3200 335 3520 3955
rect 3840 655 4160 4275
rect 4480 335 4800 3955
rect 5120 655 5440 4275
rect 5760 335 6080 3955
rect 6400 655 6720 4275
rect 7040 335 7360 3955
rect 7680 655 8000 4275
rect 8320 335 8640 3955
rect 8960 655 9280 4275
rect 9600 335 9920 3955
rect 10240 655 11146 4275
rect 0 311 11146 335
rect 0 75 272 311
rect 508 75 1712 311
rect 1948 75 3152 311
rect 3388 75 4592 311
rect 4828 75 6032 311
rect 6268 75 7472 311
rect 7708 75 8912 311
rect 9148 75 10352 311
rect 10588 75 11146 311
rect 0 0 11146 75
<< properties >>
string GDS_END 5432286
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5276250
<< end >>
