magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 4700 2026
<< mvnmos >>
rect 0 0 100 2000
rect 156 0 256 2000
rect 312 0 412 2000
rect 468 0 568 2000
rect 624 0 724 2000
rect 780 0 880 2000
rect 936 0 1036 2000
rect 1092 0 1192 2000
rect 1248 0 1348 2000
rect 1404 0 1504 2000
rect 1560 0 1660 2000
rect 1716 0 1816 2000
rect 1872 0 1972 2000
rect 2028 0 2128 2000
rect 2184 0 2284 2000
rect 2340 0 2440 2000
rect 2496 0 2596 2000
rect 2652 0 2752 2000
rect 2808 0 2908 2000
rect 2964 0 3064 2000
rect 3120 0 3220 2000
rect 3276 0 3376 2000
rect 3432 0 3532 2000
rect 3588 0 3688 2000
rect 3744 0 3844 2000
rect 3900 0 4000 2000
rect 4056 0 4156 2000
rect 4212 0 4312 2000
rect 4368 0 4468 2000
rect 4524 0 4624 2000
<< mvndiff >>
rect -50 0 0 2000
rect 4624 0 4674 2000
<< poly >>
rect 0 2000 100 2032
rect 0 -32 100 0
rect 156 2000 256 2032
rect 156 -32 256 0
rect 312 2000 412 2032
rect 312 -32 412 0
rect 468 2000 568 2032
rect 468 -32 568 0
rect 624 2000 724 2032
rect 624 -32 724 0
rect 780 2000 880 2032
rect 780 -32 880 0
rect 936 2000 1036 2032
rect 936 -32 1036 0
rect 1092 2000 1192 2032
rect 1092 -32 1192 0
rect 1248 2000 1348 2032
rect 1248 -32 1348 0
rect 1404 2000 1504 2032
rect 1404 -32 1504 0
rect 1560 2000 1660 2032
rect 1560 -32 1660 0
rect 1716 2000 1816 2032
rect 1716 -32 1816 0
rect 1872 2000 1972 2032
rect 1872 -32 1972 0
rect 2028 2000 2128 2032
rect 2028 -32 2128 0
rect 2184 2000 2284 2032
rect 2184 -32 2284 0
rect 2340 2000 2440 2032
rect 2340 -32 2440 0
rect 2496 2000 2596 2032
rect 2496 -32 2596 0
rect 2652 2000 2752 2032
rect 2652 -32 2752 0
rect 2808 2000 2908 2032
rect 2808 -32 2908 0
rect 2964 2000 3064 2032
rect 2964 -32 3064 0
rect 3120 2000 3220 2032
rect 3120 -32 3220 0
rect 3276 2000 3376 2032
rect 3276 -32 3376 0
rect 3432 2000 3532 2032
rect 3432 -32 3532 0
rect 3588 2000 3688 2032
rect 3588 -32 3688 0
rect 3744 2000 3844 2032
rect 3744 -32 3844 0
rect 3900 2000 4000 2032
rect 3900 -32 4000 0
rect 4056 2000 4156 2032
rect 4056 -32 4156 0
rect 4212 2000 4312 2032
rect 4212 -32 4312 0
rect 4368 2000 4468 2032
rect 4368 -32 4468 0
rect 4524 2000 4624 2032
rect 4524 -32 4624 0
<< metal1 >>
rect -51 -16 -5 1986
rect 105 -16 151 1986
rect 261 -16 307 1986
rect 417 -16 463 1986
rect 573 -16 619 1986
rect 729 -16 775 1986
rect 885 -16 931 1986
rect 1041 -16 1087 1986
rect 1197 -16 1243 1986
rect 1353 -16 1399 1986
rect 1509 -16 1555 1986
rect 1665 -16 1711 1986
rect 1821 -16 1867 1986
rect 1977 -16 2023 1986
rect 2133 -16 2179 1986
rect 2289 -16 2335 1986
rect 2445 -16 2491 1986
rect 2601 -16 2647 1986
rect 2757 -16 2803 1986
rect 2913 -16 2959 1986
rect 3069 -16 3115 1986
rect 3225 -16 3271 1986
rect 3381 -16 3427 1986
rect 3537 -16 3583 1986
rect 3693 -16 3739 1986
rect 3849 -16 3895 1986
rect 4005 -16 4051 1986
rect 4161 -16 4207 1986
rect 4317 -16 4363 1986
rect 4473 -16 4519 1986
rect 4629 -16 4675 1986
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_1
timestamp 1701704242
transform 1 0 100 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_2
timestamp 1701704242
transform 1 0 256 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_3
timestamp 1701704242
transform 1 0 412 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_4
timestamp 1701704242
transform 1 0 568 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_5
timestamp 1701704242
transform 1 0 724 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_6
timestamp 1701704242
transform 1 0 880 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_7
timestamp 1701704242
transform 1 0 1036 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_8
timestamp 1701704242
transform 1 0 1192 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_9
timestamp 1701704242
transform 1 0 1348 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_10
timestamp 1701704242
transform 1 0 1504 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_11
timestamp 1701704242
transform 1 0 1660 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_12
timestamp 1701704242
transform 1 0 1816 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_13
timestamp 1701704242
transform 1 0 1972 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_14
timestamp 1701704242
transform 1 0 2128 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_15
timestamp 1701704242
transform 1 0 2284 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_16
timestamp 1701704242
transform 1 0 2440 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_17
timestamp 1701704242
transform 1 0 2596 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_18
timestamp 1701704242
transform 1 0 2752 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_19
timestamp 1701704242
transform 1 0 2908 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_20
timestamp 1701704242
transform 1 0 3064 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_21
timestamp 1701704242
transform 1 0 3220 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_22
timestamp 1701704242
transform 1 0 3376 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_23
timestamp 1701704242
transform 1 0 3532 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_24
timestamp 1701704242
transform 1 0 3688 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_25
timestamp 1701704242
transform 1 0 3844 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_26
timestamp 1701704242
transform 1 0 4000 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_27
timestamp 1701704242
transform 1 0 4156 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_28
timestamp 1701704242
transform 1 0 4312 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_29
timestamp 1701704242
transform 1 0 4468 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5595914180829  hvDFM1sd2_CDNS_5595914180829_30
timestamp 1701704242
transform 1 0 4624 0 1 0
box -26 -26 82 2026
<< labels >>
flabel comment s 4652 985 4652 985 0 FreeSans 300 0 0 0 S
flabel comment s 4496 985 4496 985 0 FreeSans 300 0 0 0 D
flabel comment s 4340 985 4340 985 0 FreeSans 300 0 0 0 S
flabel comment s 4184 985 4184 985 0 FreeSans 300 0 0 0 D
flabel comment s 4028 985 4028 985 0 FreeSans 300 0 0 0 S
flabel comment s 3872 985 3872 985 0 FreeSans 300 0 0 0 D
flabel comment s 3716 985 3716 985 0 FreeSans 300 0 0 0 S
flabel comment s 3560 985 3560 985 0 FreeSans 300 0 0 0 D
flabel comment s 3404 985 3404 985 0 FreeSans 300 0 0 0 S
flabel comment s 3248 985 3248 985 0 FreeSans 300 0 0 0 D
flabel comment s 3092 985 3092 985 0 FreeSans 300 0 0 0 S
flabel comment s 2936 985 2936 985 0 FreeSans 300 0 0 0 D
flabel comment s 2780 985 2780 985 0 FreeSans 300 0 0 0 S
flabel comment s 2624 985 2624 985 0 FreeSans 300 0 0 0 D
flabel comment s 2468 985 2468 985 0 FreeSans 300 0 0 0 S
flabel comment s 2312 985 2312 985 0 FreeSans 300 0 0 0 D
flabel comment s 2156 985 2156 985 0 FreeSans 300 0 0 0 S
flabel comment s 2000 985 2000 985 0 FreeSans 300 0 0 0 D
flabel comment s 1844 985 1844 985 0 FreeSans 300 0 0 0 S
flabel comment s 1688 985 1688 985 0 FreeSans 300 0 0 0 D
flabel comment s 1532 985 1532 985 0 FreeSans 300 0 0 0 S
flabel comment s 1376 985 1376 985 0 FreeSans 300 0 0 0 D
flabel comment s 1220 985 1220 985 0 FreeSans 300 0 0 0 S
flabel comment s 1064 985 1064 985 0 FreeSans 300 0 0 0 D
flabel comment s 908 985 908 985 0 FreeSans 300 0 0 0 S
flabel comment s 752 985 752 985 0 FreeSans 300 0 0 0 D
flabel comment s 596 985 596 985 0 FreeSans 300 0 0 0 S
flabel comment s 440 985 440 985 0 FreeSans 300 0 0 0 D
flabel comment s 284 985 284 985 0 FreeSans 300 0 0 0 S
flabel comment s 128 985 128 985 0 FreeSans 300 0 0 0 D
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 36836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21504
<< end >>
