magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -36 679 404 1471
<< locali >>
rect 0 1397 368 1431
rect 64 674 98 740
rect 179 690 213 724
rect 0 -17 368 17
use pinv_17  pinv_17_0
timestamp 1701704242
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 196 707 196 707 4 Z
port 2 nsew
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 184 1414 184 1414 4 vdd
port 3 nsew
rlabel locali s 184 0 184 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1414
string GDS_END 4087524
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4086684
<< end >>
