magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 88 579 15088 5356
<< nwell >>
rect 0 5150 15173 5493
rect 0 785 362 5150
rect 14811 785 15173 5150
rect 0 423 15173 785
<< pwell >>
rect 529 4760 14693 4982
rect 529 4084 751 4760
rect 14471 4084 14693 4760
rect 529 3032 14693 4084
rect 529 2483 751 3032
rect 1552 2483 1840 3032
rect 2544 2483 2832 3032
rect 3536 2483 3824 3032
rect 4528 2483 4816 3032
rect 5520 2483 5808 3032
rect 6512 2483 6800 3032
rect 7504 2483 7792 3032
rect 8496 2483 8784 3032
rect 9488 2483 9776 3032
rect 10480 2483 10768 3032
rect 11472 2483 11760 3032
rect 12464 2483 12752 3032
rect 13456 2483 13744 3032
rect 14471 2483 14693 3032
rect 529 1431 14693 2483
rect 529 1174 751 1431
rect 14471 1174 14693 1431
rect 529 952 14693 1174
<< mvnmos >>
rect 924 3058 1044 4058
rect 1354 3058 1474 4058
rect 1916 3058 2036 4058
rect 2346 3058 2466 4058
rect 2908 3058 3028 4058
rect 3338 3058 3458 4058
rect 3900 3058 4020 4058
rect 4330 3058 4450 4058
rect 4892 3058 5012 4058
rect 5322 3058 5442 4058
rect 5884 3058 6004 4058
rect 6314 3058 6434 4058
rect 6876 3058 6996 4058
rect 7306 3058 7426 4058
rect 7868 3058 7988 4058
rect 8298 3058 8418 4058
rect 8860 3058 8980 4058
rect 9290 3058 9410 4058
rect 9852 3058 9972 4058
rect 10282 3058 10402 4058
rect 10844 3058 10964 4058
rect 11274 3058 11394 4058
rect 11836 3058 11956 4058
rect 12266 3058 12386 4058
rect 12828 3058 12948 4058
rect 13258 3058 13378 4058
rect 13820 3058 13940 4058
rect 14178 3058 14298 4058
rect 924 1457 1044 2457
rect 1354 1457 1474 2457
rect 1916 1457 2036 2457
rect 2346 1457 2466 2457
rect 2908 1457 3028 2457
rect 3338 1457 3458 2457
rect 3900 1457 4020 2457
rect 4330 1457 4450 2457
rect 4892 1457 5012 2457
rect 5322 1457 5442 2457
rect 5884 1457 6004 2457
rect 6314 1457 6434 2457
rect 6876 1457 6996 2457
rect 7306 1457 7426 2457
rect 7868 1457 7988 2457
rect 8298 1457 8418 2457
rect 8860 1457 8980 2457
rect 9290 1457 9410 2457
rect 9852 1457 9972 2457
rect 10282 1457 10402 2457
rect 10844 1457 10964 2457
rect 11274 1457 11394 2457
rect 11836 1457 11956 2457
rect 12266 1457 12386 2457
rect 12828 1457 12948 2457
rect 13258 1457 13378 2457
rect 13820 1457 13940 2457
rect 14178 1457 14298 2457
<< mvndiff >>
rect 787 4046 924 4058
rect 787 4012 802 4046
rect 836 4012 924 4046
rect 787 3978 924 4012
rect 787 3944 802 3978
rect 836 3944 924 3978
rect 787 3910 924 3944
rect 787 3876 802 3910
rect 836 3876 924 3910
rect 787 3842 924 3876
rect 787 3808 802 3842
rect 836 3808 924 3842
rect 787 3774 924 3808
rect 787 3740 802 3774
rect 836 3740 924 3774
rect 787 3706 924 3740
rect 787 3672 802 3706
rect 836 3672 924 3706
rect 787 3638 924 3672
rect 787 3604 802 3638
rect 836 3604 924 3638
rect 787 3570 924 3604
rect 787 3536 802 3570
rect 836 3536 924 3570
rect 787 3502 924 3536
rect 787 3468 802 3502
rect 836 3468 924 3502
rect 787 3434 924 3468
rect 787 3400 802 3434
rect 836 3400 924 3434
rect 787 3366 924 3400
rect 787 3332 802 3366
rect 836 3332 924 3366
rect 787 3298 924 3332
rect 787 3264 802 3298
rect 836 3264 924 3298
rect 787 3230 924 3264
rect 787 3196 802 3230
rect 836 3196 924 3230
rect 787 3162 924 3196
rect 787 3128 802 3162
rect 836 3128 924 3162
rect 787 3058 924 3128
rect 1044 4046 1354 4058
rect 1044 4012 1146 4046
rect 1180 4012 1218 4046
rect 1252 4012 1354 4046
rect 1044 3978 1354 4012
rect 1044 3944 1146 3978
rect 1180 3944 1218 3978
rect 1252 3944 1354 3978
rect 1044 3910 1354 3944
rect 1044 3876 1146 3910
rect 1180 3876 1218 3910
rect 1252 3876 1354 3910
rect 1044 3842 1354 3876
rect 1044 3808 1146 3842
rect 1180 3808 1218 3842
rect 1252 3808 1354 3842
rect 1044 3774 1354 3808
rect 1044 3740 1146 3774
rect 1180 3740 1218 3774
rect 1252 3740 1354 3774
rect 1044 3706 1354 3740
rect 1044 3672 1146 3706
rect 1180 3672 1218 3706
rect 1252 3672 1354 3706
rect 1044 3638 1354 3672
rect 1044 3604 1146 3638
rect 1180 3604 1218 3638
rect 1252 3604 1354 3638
rect 1044 3570 1354 3604
rect 1044 3536 1146 3570
rect 1180 3536 1218 3570
rect 1252 3536 1354 3570
rect 1044 3502 1354 3536
rect 1044 3468 1146 3502
rect 1180 3468 1218 3502
rect 1252 3468 1354 3502
rect 1044 3434 1354 3468
rect 1044 3400 1146 3434
rect 1180 3400 1218 3434
rect 1252 3400 1354 3434
rect 1044 3366 1354 3400
rect 1044 3332 1146 3366
rect 1180 3332 1218 3366
rect 1252 3332 1354 3366
rect 1044 3298 1354 3332
rect 1044 3264 1146 3298
rect 1180 3264 1218 3298
rect 1252 3264 1354 3298
rect 1044 3230 1354 3264
rect 1044 3196 1146 3230
rect 1180 3196 1218 3230
rect 1252 3196 1354 3230
rect 1044 3162 1354 3196
rect 1044 3128 1146 3162
rect 1180 3128 1218 3162
rect 1252 3128 1354 3162
rect 1044 3058 1354 3128
rect 1474 4046 1625 4058
rect 1765 4046 1916 4058
rect 1474 4012 1576 4046
rect 1610 4012 1625 4046
rect 1765 4012 1780 4046
rect 1814 4012 1916 4046
rect 1474 3978 1625 4012
rect 1765 3978 1916 4012
rect 1474 3944 1576 3978
rect 1610 3944 1625 3978
rect 1765 3944 1780 3978
rect 1814 3944 1916 3978
rect 1474 3910 1625 3944
rect 1765 3910 1916 3944
rect 1474 3876 1576 3910
rect 1610 3876 1625 3910
rect 1765 3876 1780 3910
rect 1814 3876 1916 3910
rect 1474 3842 1625 3876
rect 1765 3842 1916 3876
rect 1474 3808 1576 3842
rect 1610 3808 1625 3842
rect 1765 3808 1780 3842
rect 1814 3808 1916 3842
rect 1474 3774 1625 3808
rect 1765 3774 1916 3808
rect 1474 3740 1576 3774
rect 1610 3740 1625 3774
rect 1765 3740 1780 3774
rect 1814 3740 1916 3774
rect 1474 3706 1625 3740
rect 1765 3706 1916 3740
rect 1474 3672 1576 3706
rect 1610 3672 1625 3706
rect 1765 3672 1780 3706
rect 1814 3672 1916 3706
rect 1474 3638 1625 3672
rect 1765 3638 1916 3672
rect 1474 3604 1576 3638
rect 1610 3604 1625 3638
rect 1765 3604 1780 3638
rect 1814 3604 1916 3638
rect 1474 3570 1625 3604
rect 1765 3570 1916 3604
rect 1474 3536 1576 3570
rect 1610 3536 1625 3570
rect 1765 3536 1780 3570
rect 1814 3536 1916 3570
rect 1474 3502 1625 3536
rect 1765 3502 1916 3536
rect 1474 3468 1576 3502
rect 1610 3468 1625 3502
rect 1765 3468 1780 3502
rect 1814 3468 1916 3502
rect 1474 3434 1625 3468
rect 1765 3434 1916 3468
rect 1474 3400 1576 3434
rect 1610 3400 1625 3434
rect 1765 3400 1780 3434
rect 1814 3400 1916 3434
rect 1474 3366 1625 3400
rect 1765 3366 1916 3400
rect 1474 3332 1576 3366
rect 1610 3332 1625 3366
rect 1765 3332 1780 3366
rect 1814 3332 1916 3366
rect 1474 3298 1625 3332
rect 1765 3298 1916 3332
rect 1474 3264 1576 3298
rect 1610 3264 1625 3298
rect 1765 3264 1780 3298
rect 1814 3264 1916 3298
rect 1474 3230 1625 3264
rect 1765 3230 1916 3264
rect 1474 3196 1576 3230
rect 1610 3196 1625 3230
rect 1765 3196 1780 3230
rect 1814 3196 1916 3230
rect 1474 3162 1625 3196
rect 1765 3162 1916 3196
rect 1474 3128 1576 3162
rect 1610 3128 1625 3162
rect 1765 3128 1780 3162
rect 1814 3128 1916 3162
rect 1474 3058 1625 3128
rect 1765 3058 1916 3128
rect 2036 4046 2346 4058
rect 2036 4012 2138 4046
rect 2172 4012 2210 4046
rect 2244 4012 2346 4046
rect 2036 3978 2346 4012
rect 2036 3944 2138 3978
rect 2172 3944 2210 3978
rect 2244 3944 2346 3978
rect 2036 3910 2346 3944
rect 2036 3876 2138 3910
rect 2172 3876 2210 3910
rect 2244 3876 2346 3910
rect 2036 3842 2346 3876
rect 2036 3808 2138 3842
rect 2172 3808 2210 3842
rect 2244 3808 2346 3842
rect 2036 3774 2346 3808
rect 2036 3740 2138 3774
rect 2172 3740 2210 3774
rect 2244 3740 2346 3774
rect 2036 3706 2346 3740
rect 2036 3672 2138 3706
rect 2172 3672 2210 3706
rect 2244 3672 2346 3706
rect 2036 3638 2346 3672
rect 2036 3604 2138 3638
rect 2172 3604 2210 3638
rect 2244 3604 2346 3638
rect 2036 3570 2346 3604
rect 2036 3536 2138 3570
rect 2172 3536 2210 3570
rect 2244 3536 2346 3570
rect 2036 3502 2346 3536
rect 2036 3468 2138 3502
rect 2172 3468 2210 3502
rect 2244 3468 2346 3502
rect 2036 3434 2346 3468
rect 2036 3400 2138 3434
rect 2172 3400 2210 3434
rect 2244 3400 2346 3434
rect 2036 3366 2346 3400
rect 2036 3332 2138 3366
rect 2172 3332 2210 3366
rect 2244 3332 2346 3366
rect 2036 3298 2346 3332
rect 2036 3264 2138 3298
rect 2172 3264 2210 3298
rect 2244 3264 2346 3298
rect 2036 3230 2346 3264
rect 2036 3196 2138 3230
rect 2172 3196 2210 3230
rect 2244 3196 2346 3230
rect 2036 3162 2346 3196
rect 2036 3128 2138 3162
rect 2172 3128 2210 3162
rect 2244 3128 2346 3162
rect 2036 3058 2346 3128
rect 2466 4046 2617 4058
rect 2757 4046 2908 4058
rect 2466 4012 2568 4046
rect 2602 4012 2617 4046
rect 2757 4012 2772 4046
rect 2806 4012 2908 4046
rect 2466 3978 2617 4012
rect 2757 3978 2908 4012
rect 2466 3944 2568 3978
rect 2602 3944 2617 3978
rect 2757 3944 2772 3978
rect 2806 3944 2908 3978
rect 2466 3910 2617 3944
rect 2757 3910 2908 3944
rect 2466 3876 2568 3910
rect 2602 3876 2617 3910
rect 2757 3876 2772 3910
rect 2806 3876 2908 3910
rect 2466 3842 2617 3876
rect 2757 3842 2908 3876
rect 2466 3808 2568 3842
rect 2602 3808 2617 3842
rect 2757 3808 2772 3842
rect 2806 3808 2908 3842
rect 2466 3774 2617 3808
rect 2757 3774 2908 3808
rect 2466 3740 2568 3774
rect 2602 3740 2617 3774
rect 2757 3740 2772 3774
rect 2806 3740 2908 3774
rect 2466 3706 2617 3740
rect 2757 3706 2908 3740
rect 2466 3672 2568 3706
rect 2602 3672 2617 3706
rect 2757 3672 2772 3706
rect 2806 3672 2908 3706
rect 2466 3638 2617 3672
rect 2757 3638 2908 3672
rect 2466 3604 2568 3638
rect 2602 3604 2617 3638
rect 2757 3604 2772 3638
rect 2806 3604 2908 3638
rect 2466 3570 2617 3604
rect 2757 3570 2908 3604
rect 2466 3536 2568 3570
rect 2602 3536 2617 3570
rect 2757 3536 2772 3570
rect 2806 3536 2908 3570
rect 2466 3502 2617 3536
rect 2757 3502 2908 3536
rect 2466 3468 2568 3502
rect 2602 3468 2617 3502
rect 2757 3468 2772 3502
rect 2806 3468 2908 3502
rect 2466 3434 2617 3468
rect 2757 3434 2908 3468
rect 2466 3400 2568 3434
rect 2602 3400 2617 3434
rect 2757 3400 2772 3434
rect 2806 3400 2908 3434
rect 2466 3366 2617 3400
rect 2757 3366 2908 3400
rect 2466 3332 2568 3366
rect 2602 3332 2617 3366
rect 2757 3332 2772 3366
rect 2806 3332 2908 3366
rect 2466 3298 2617 3332
rect 2757 3298 2908 3332
rect 2466 3264 2568 3298
rect 2602 3264 2617 3298
rect 2757 3264 2772 3298
rect 2806 3264 2908 3298
rect 2466 3230 2617 3264
rect 2757 3230 2908 3264
rect 2466 3196 2568 3230
rect 2602 3196 2617 3230
rect 2757 3196 2772 3230
rect 2806 3196 2908 3230
rect 2466 3162 2617 3196
rect 2757 3162 2908 3196
rect 2466 3128 2568 3162
rect 2602 3128 2617 3162
rect 2757 3128 2772 3162
rect 2806 3128 2908 3162
rect 2466 3058 2617 3128
rect 2757 3058 2908 3128
rect 3028 4046 3338 4058
rect 3028 4012 3130 4046
rect 3164 4012 3202 4046
rect 3236 4012 3338 4046
rect 3028 3978 3338 4012
rect 3028 3944 3130 3978
rect 3164 3944 3202 3978
rect 3236 3944 3338 3978
rect 3028 3910 3338 3944
rect 3028 3876 3130 3910
rect 3164 3876 3202 3910
rect 3236 3876 3338 3910
rect 3028 3842 3338 3876
rect 3028 3808 3130 3842
rect 3164 3808 3202 3842
rect 3236 3808 3338 3842
rect 3028 3774 3338 3808
rect 3028 3740 3130 3774
rect 3164 3740 3202 3774
rect 3236 3740 3338 3774
rect 3028 3706 3338 3740
rect 3028 3672 3130 3706
rect 3164 3672 3202 3706
rect 3236 3672 3338 3706
rect 3028 3638 3338 3672
rect 3028 3604 3130 3638
rect 3164 3604 3202 3638
rect 3236 3604 3338 3638
rect 3028 3570 3338 3604
rect 3028 3536 3130 3570
rect 3164 3536 3202 3570
rect 3236 3536 3338 3570
rect 3028 3502 3338 3536
rect 3028 3468 3130 3502
rect 3164 3468 3202 3502
rect 3236 3468 3338 3502
rect 3028 3434 3338 3468
rect 3028 3400 3130 3434
rect 3164 3400 3202 3434
rect 3236 3400 3338 3434
rect 3028 3366 3338 3400
rect 3028 3332 3130 3366
rect 3164 3332 3202 3366
rect 3236 3332 3338 3366
rect 3028 3298 3338 3332
rect 3028 3264 3130 3298
rect 3164 3264 3202 3298
rect 3236 3264 3338 3298
rect 3028 3230 3338 3264
rect 3028 3196 3130 3230
rect 3164 3196 3202 3230
rect 3236 3196 3338 3230
rect 3028 3162 3338 3196
rect 3028 3128 3130 3162
rect 3164 3128 3202 3162
rect 3236 3128 3338 3162
rect 3028 3058 3338 3128
rect 3458 4046 3609 4058
rect 3749 4046 3900 4058
rect 3458 4012 3560 4046
rect 3594 4012 3609 4046
rect 3749 4012 3764 4046
rect 3798 4012 3900 4046
rect 3458 3978 3609 4012
rect 3749 3978 3900 4012
rect 3458 3944 3560 3978
rect 3594 3944 3609 3978
rect 3749 3944 3764 3978
rect 3798 3944 3900 3978
rect 3458 3910 3609 3944
rect 3749 3910 3900 3944
rect 3458 3876 3560 3910
rect 3594 3876 3609 3910
rect 3749 3876 3764 3910
rect 3798 3876 3900 3910
rect 3458 3842 3609 3876
rect 3749 3842 3900 3876
rect 3458 3808 3560 3842
rect 3594 3808 3609 3842
rect 3749 3808 3764 3842
rect 3798 3808 3900 3842
rect 3458 3774 3609 3808
rect 3749 3774 3900 3808
rect 3458 3740 3560 3774
rect 3594 3740 3609 3774
rect 3749 3740 3764 3774
rect 3798 3740 3900 3774
rect 3458 3706 3609 3740
rect 3749 3706 3900 3740
rect 3458 3672 3560 3706
rect 3594 3672 3609 3706
rect 3749 3672 3764 3706
rect 3798 3672 3900 3706
rect 3458 3638 3609 3672
rect 3749 3638 3900 3672
rect 3458 3604 3560 3638
rect 3594 3604 3609 3638
rect 3749 3604 3764 3638
rect 3798 3604 3900 3638
rect 3458 3570 3609 3604
rect 3749 3570 3900 3604
rect 3458 3536 3560 3570
rect 3594 3536 3609 3570
rect 3749 3536 3764 3570
rect 3798 3536 3900 3570
rect 3458 3502 3609 3536
rect 3749 3502 3900 3536
rect 3458 3468 3560 3502
rect 3594 3468 3609 3502
rect 3749 3468 3764 3502
rect 3798 3468 3900 3502
rect 3458 3434 3609 3468
rect 3749 3434 3900 3468
rect 3458 3400 3560 3434
rect 3594 3400 3609 3434
rect 3749 3400 3764 3434
rect 3798 3400 3900 3434
rect 3458 3366 3609 3400
rect 3749 3366 3900 3400
rect 3458 3332 3560 3366
rect 3594 3332 3609 3366
rect 3749 3332 3764 3366
rect 3798 3332 3900 3366
rect 3458 3298 3609 3332
rect 3749 3298 3900 3332
rect 3458 3264 3560 3298
rect 3594 3264 3609 3298
rect 3749 3264 3764 3298
rect 3798 3264 3900 3298
rect 3458 3230 3609 3264
rect 3749 3230 3900 3264
rect 3458 3196 3560 3230
rect 3594 3196 3609 3230
rect 3749 3196 3764 3230
rect 3798 3196 3900 3230
rect 3458 3162 3609 3196
rect 3749 3162 3900 3196
rect 3458 3128 3560 3162
rect 3594 3128 3609 3162
rect 3749 3128 3764 3162
rect 3798 3128 3900 3162
rect 3458 3058 3609 3128
rect 3749 3058 3900 3128
rect 4020 4046 4330 4058
rect 4020 4012 4122 4046
rect 4156 4012 4194 4046
rect 4228 4012 4330 4046
rect 4020 3978 4330 4012
rect 4020 3944 4122 3978
rect 4156 3944 4194 3978
rect 4228 3944 4330 3978
rect 4020 3910 4330 3944
rect 4020 3876 4122 3910
rect 4156 3876 4194 3910
rect 4228 3876 4330 3910
rect 4020 3842 4330 3876
rect 4020 3808 4122 3842
rect 4156 3808 4194 3842
rect 4228 3808 4330 3842
rect 4020 3774 4330 3808
rect 4020 3740 4122 3774
rect 4156 3740 4194 3774
rect 4228 3740 4330 3774
rect 4020 3706 4330 3740
rect 4020 3672 4122 3706
rect 4156 3672 4194 3706
rect 4228 3672 4330 3706
rect 4020 3638 4330 3672
rect 4020 3604 4122 3638
rect 4156 3604 4194 3638
rect 4228 3604 4330 3638
rect 4020 3570 4330 3604
rect 4020 3536 4122 3570
rect 4156 3536 4194 3570
rect 4228 3536 4330 3570
rect 4020 3502 4330 3536
rect 4020 3468 4122 3502
rect 4156 3468 4194 3502
rect 4228 3468 4330 3502
rect 4020 3434 4330 3468
rect 4020 3400 4122 3434
rect 4156 3400 4194 3434
rect 4228 3400 4330 3434
rect 4020 3366 4330 3400
rect 4020 3332 4122 3366
rect 4156 3332 4194 3366
rect 4228 3332 4330 3366
rect 4020 3298 4330 3332
rect 4020 3264 4122 3298
rect 4156 3264 4194 3298
rect 4228 3264 4330 3298
rect 4020 3230 4330 3264
rect 4020 3196 4122 3230
rect 4156 3196 4194 3230
rect 4228 3196 4330 3230
rect 4020 3162 4330 3196
rect 4020 3128 4122 3162
rect 4156 3128 4194 3162
rect 4228 3128 4330 3162
rect 4020 3058 4330 3128
rect 4450 4046 4601 4058
rect 4741 4046 4892 4058
rect 4450 4012 4552 4046
rect 4586 4012 4601 4046
rect 4741 4012 4756 4046
rect 4790 4012 4892 4046
rect 4450 3978 4601 4012
rect 4741 3978 4892 4012
rect 4450 3944 4552 3978
rect 4586 3944 4601 3978
rect 4741 3944 4756 3978
rect 4790 3944 4892 3978
rect 4450 3910 4601 3944
rect 4741 3910 4892 3944
rect 4450 3876 4552 3910
rect 4586 3876 4601 3910
rect 4741 3876 4756 3910
rect 4790 3876 4892 3910
rect 4450 3842 4601 3876
rect 4741 3842 4892 3876
rect 4450 3808 4552 3842
rect 4586 3808 4601 3842
rect 4741 3808 4756 3842
rect 4790 3808 4892 3842
rect 4450 3774 4601 3808
rect 4741 3774 4892 3808
rect 4450 3740 4552 3774
rect 4586 3740 4601 3774
rect 4741 3740 4756 3774
rect 4790 3740 4892 3774
rect 4450 3706 4601 3740
rect 4741 3706 4892 3740
rect 4450 3672 4552 3706
rect 4586 3672 4601 3706
rect 4741 3672 4756 3706
rect 4790 3672 4892 3706
rect 4450 3638 4601 3672
rect 4741 3638 4892 3672
rect 4450 3604 4552 3638
rect 4586 3604 4601 3638
rect 4741 3604 4756 3638
rect 4790 3604 4892 3638
rect 4450 3570 4601 3604
rect 4741 3570 4892 3604
rect 4450 3536 4552 3570
rect 4586 3536 4601 3570
rect 4741 3536 4756 3570
rect 4790 3536 4892 3570
rect 4450 3502 4601 3536
rect 4741 3502 4892 3536
rect 4450 3468 4552 3502
rect 4586 3468 4601 3502
rect 4741 3468 4756 3502
rect 4790 3468 4892 3502
rect 4450 3434 4601 3468
rect 4741 3434 4892 3468
rect 4450 3400 4552 3434
rect 4586 3400 4601 3434
rect 4741 3400 4756 3434
rect 4790 3400 4892 3434
rect 4450 3366 4601 3400
rect 4741 3366 4892 3400
rect 4450 3332 4552 3366
rect 4586 3332 4601 3366
rect 4741 3332 4756 3366
rect 4790 3332 4892 3366
rect 4450 3298 4601 3332
rect 4741 3298 4892 3332
rect 4450 3264 4552 3298
rect 4586 3264 4601 3298
rect 4741 3264 4756 3298
rect 4790 3264 4892 3298
rect 4450 3230 4601 3264
rect 4741 3230 4892 3264
rect 4450 3196 4552 3230
rect 4586 3196 4601 3230
rect 4741 3196 4756 3230
rect 4790 3196 4892 3230
rect 4450 3162 4601 3196
rect 4741 3162 4892 3196
rect 4450 3128 4552 3162
rect 4586 3128 4601 3162
rect 4741 3128 4756 3162
rect 4790 3128 4892 3162
rect 4450 3058 4601 3128
rect 4741 3058 4892 3128
rect 5012 4046 5322 4058
rect 5012 4012 5114 4046
rect 5148 4012 5186 4046
rect 5220 4012 5322 4046
rect 5012 3978 5322 4012
rect 5012 3944 5114 3978
rect 5148 3944 5186 3978
rect 5220 3944 5322 3978
rect 5012 3910 5322 3944
rect 5012 3876 5114 3910
rect 5148 3876 5186 3910
rect 5220 3876 5322 3910
rect 5012 3842 5322 3876
rect 5012 3808 5114 3842
rect 5148 3808 5186 3842
rect 5220 3808 5322 3842
rect 5012 3774 5322 3808
rect 5012 3740 5114 3774
rect 5148 3740 5186 3774
rect 5220 3740 5322 3774
rect 5012 3706 5322 3740
rect 5012 3672 5114 3706
rect 5148 3672 5186 3706
rect 5220 3672 5322 3706
rect 5012 3638 5322 3672
rect 5012 3604 5114 3638
rect 5148 3604 5186 3638
rect 5220 3604 5322 3638
rect 5012 3570 5322 3604
rect 5012 3536 5114 3570
rect 5148 3536 5186 3570
rect 5220 3536 5322 3570
rect 5012 3502 5322 3536
rect 5012 3468 5114 3502
rect 5148 3468 5186 3502
rect 5220 3468 5322 3502
rect 5012 3434 5322 3468
rect 5012 3400 5114 3434
rect 5148 3400 5186 3434
rect 5220 3400 5322 3434
rect 5012 3366 5322 3400
rect 5012 3332 5114 3366
rect 5148 3332 5186 3366
rect 5220 3332 5322 3366
rect 5012 3298 5322 3332
rect 5012 3264 5114 3298
rect 5148 3264 5186 3298
rect 5220 3264 5322 3298
rect 5012 3230 5322 3264
rect 5012 3196 5114 3230
rect 5148 3196 5186 3230
rect 5220 3196 5322 3230
rect 5012 3162 5322 3196
rect 5012 3128 5114 3162
rect 5148 3128 5186 3162
rect 5220 3128 5322 3162
rect 5012 3058 5322 3128
rect 5442 4046 5593 4058
rect 5733 4046 5884 4058
rect 5442 4012 5544 4046
rect 5578 4012 5593 4046
rect 5733 4012 5748 4046
rect 5782 4012 5884 4046
rect 5442 3978 5593 4012
rect 5733 3978 5884 4012
rect 5442 3944 5544 3978
rect 5578 3944 5593 3978
rect 5733 3944 5748 3978
rect 5782 3944 5884 3978
rect 5442 3910 5593 3944
rect 5733 3910 5884 3944
rect 5442 3876 5544 3910
rect 5578 3876 5593 3910
rect 5733 3876 5748 3910
rect 5782 3876 5884 3910
rect 5442 3842 5593 3876
rect 5733 3842 5884 3876
rect 5442 3808 5544 3842
rect 5578 3808 5593 3842
rect 5733 3808 5748 3842
rect 5782 3808 5884 3842
rect 5442 3774 5593 3808
rect 5733 3774 5884 3808
rect 5442 3740 5544 3774
rect 5578 3740 5593 3774
rect 5733 3740 5748 3774
rect 5782 3740 5884 3774
rect 5442 3706 5593 3740
rect 5733 3706 5884 3740
rect 5442 3672 5544 3706
rect 5578 3672 5593 3706
rect 5733 3672 5748 3706
rect 5782 3672 5884 3706
rect 5442 3638 5593 3672
rect 5733 3638 5884 3672
rect 5442 3604 5544 3638
rect 5578 3604 5593 3638
rect 5733 3604 5748 3638
rect 5782 3604 5884 3638
rect 5442 3570 5593 3604
rect 5733 3570 5884 3604
rect 5442 3536 5544 3570
rect 5578 3536 5593 3570
rect 5733 3536 5748 3570
rect 5782 3536 5884 3570
rect 5442 3502 5593 3536
rect 5733 3502 5884 3536
rect 5442 3468 5544 3502
rect 5578 3468 5593 3502
rect 5733 3468 5748 3502
rect 5782 3468 5884 3502
rect 5442 3434 5593 3468
rect 5733 3434 5884 3468
rect 5442 3400 5544 3434
rect 5578 3400 5593 3434
rect 5733 3400 5748 3434
rect 5782 3400 5884 3434
rect 5442 3366 5593 3400
rect 5733 3366 5884 3400
rect 5442 3332 5544 3366
rect 5578 3332 5593 3366
rect 5733 3332 5748 3366
rect 5782 3332 5884 3366
rect 5442 3298 5593 3332
rect 5733 3298 5884 3332
rect 5442 3264 5544 3298
rect 5578 3264 5593 3298
rect 5733 3264 5748 3298
rect 5782 3264 5884 3298
rect 5442 3230 5593 3264
rect 5733 3230 5884 3264
rect 5442 3196 5544 3230
rect 5578 3196 5593 3230
rect 5733 3196 5748 3230
rect 5782 3196 5884 3230
rect 5442 3162 5593 3196
rect 5733 3162 5884 3196
rect 5442 3128 5544 3162
rect 5578 3128 5593 3162
rect 5733 3128 5748 3162
rect 5782 3128 5884 3162
rect 5442 3058 5593 3128
rect 5733 3058 5884 3128
rect 6004 4046 6314 4058
rect 6004 4012 6106 4046
rect 6140 4012 6178 4046
rect 6212 4012 6314 4046
rect 6004 3978 6314 4012
rect 6004 3944 6106 3978
rect 6140 3944 6178 3978
rect 6212 3944 6314 3978
rect 6004 3910 6314 3944
rect 6004 3876 6106 3910
rect 6140 3876 6178 3910
rect 6212 3876 6314 3910
rect 6004 3842 6314 3876
rect 6004 3808 6106 3842
rect 6140 3808 6178 3842
rect 6212 3808 6314 3842
rect 6004 3774 6314 3808
rect 6004 3740 6106 3774
rect 6140 3740 6178 3774
rect 6212 3740 6314 3774
rect 6004 3706 6314 3740
rect 6004 3672 6106 3706
rect 6140 3672 6178 3706
rect 6212 3672 6314 3706
rect 6004 3638 6314 3672
rect 6004 3604 6106 3638
rect 6140 3604 6178 3638
rect 6212 3604 6314 3638
rect 6004 3570 6314 3604
rect 6004 3536 6106 3570
rect 6140 3536 6178 3570
rect 6212 3536 6314 3570
rect 6004 3502 6314 3536
rect 6004 3468 6106 3502
rect 6140 3468 6178 3502
rect 6212 3468 6314 3502
rect 6004 3434 6314 3468
rect 6004 3400 6106 3434
rect 6140 3400 6178 3434
rect 6212 3400 6314 3434
rect 6004 3366 6314 3400
rect 6004 3332 6106 3366
rect 6140 3332 6178 3366
rect 6212 3332 6314 3366
rect 6004 3298 6314 3332
rect 6004 3264 6106 3298
rect 6140 3264 6178 3298
rect 6212 3264 6314 3298
rect 6004 3230 6314 3264
rect 6004 3196 6106 3230
rect 6140 3196 6178 3230
rect 6212 3196 6314 3230
rect 6004 3162 6314 3196
rect 6004 3128 6106 3162
rect 6140 3128 6178 3162
rect 6212 3128 6314 3162
rect 6004 3058 6314 3128
rect 6434 4046 6585 4058
rect 6725 4046 6876 4058
rect 6434 4012 6536 4046
rect 6570 4012 6585 4046
rect 6725 4012 6740 4046
rect 6774 4012 6876 4046
rect 6434 3978 6585 4012
rect 6725 3978 6876 4012
rect 6434 3944 6536 3978
rect 6570 3944 6585 3978
rect 6725 3944 6740 3978
rect 6774 3944 6876 3978
rect 6434 3910 6585 3944
rect 6725 3910 6876 3944
rect 6434 3876 6536 3910
rect 6570 3876 6585 3910
rect 6725 3876 6740 3910
rect 6774 3876 6876 3910
rect 6434 3842 6585 3876
rect 6725 3842 6876 3876
rect 6434 3808 6536 3842
rect 6570 3808 6585 3842
rect 6725 3808 6740 3842
rect 6774 3808 6876 3842
rect 6434 3774 6585 3808
rect 6725 3774 6876 3808
rect 6434 3740 6536 3774
rect 6570 3740 6585 3774
rect 6725 3740 6740 3774
rect 6774 3740 6876 3774
rect 6434 3706 6585 3740
rect 6725 3706 6876 3740
rect 6434 3672 6536 3706
rect 6570 3672 6585 3706
rect 6725 3672 6740 3706
rect 6774 3672 6876 3706
rect 6434 3638 6585 3672
rect 6725 3638 6876 3672
rect 6434 3604 6536 3638
rect 6570 3604 6585 3638
rect 6725 3604 6740 3638
rect 6774 3604 6876 3638
rect 6434 3570 6585 3604
rect 6725 3570 6876 3604
rect 6434 3536 6536 3570
rect 6570 3536 6585 3570
rect 6725 3536 6740 3570
rect 6774 3536 6876 3570
rect 6434 3502 6585 3536
rect 6725 3502 6876 3536
rect 6434 3468 6536 3502
rect 6570 3468 6585 3502
rect 6725 3468 6740 3502
rect 6774 3468 6876 3502
rect 6434 3434 6585 3468
rect 6725 3434 6876 3468
rect 6434 3400 6536 3434
rect 6570 3400 6585 3434
rect 6725 3400 6740 3434
rect 6774 3400 6876 3434
rect 6434 3366 6585 3400
rect 6725 3366 6876 3400
rect 6434 3332 6536 3366
rect 6570 3332 6585 3366
rect 6725 3332 6740 3366
rect 6774 3332 6876 3366
rect 6434 3298 6585 3332
rect 6725 3298 6876 3332
rect 6434 3264 6536 3298
rect 6570 3264 6585 3298
rect 6725 3264 6740 3298
rect 6774 3264 6876 3298
rect 6434 3230 6585 3264
rect 6725 3230 6876 3264
rect 6434 3196 6536 3230
rect 6570 3196 6585 3230
rect 6725 3196 6740 3230
rect 6774 3196 6876 3230
rect 6434 3162 6585 3196
rect 6725 3162 6876 3196
rect 6434 3128 6536 3162
rect 6570 3128 6585 3162
rect 6725 3128 6740 3162
rect 6774 3128 6876 3162
rect 6434 3058 6585 3128
rect 6725 3058 6876 3128
rect 6996 4046 7306 4058
rect 6996 4012 7098 4046
rect 7132 4012 7170 4046
rect 7204 4012 7306 4046
rect 6996 3978 7306 4012
rect 6996 3944 7098 3978
rect 7132 3944 7170 3978
rect 7204 3944 7306 3978
rect 6996 3910 7306 3944
rect 6996 3876 7098 3910
rect 7132 3876 7170 3910
rect 7204 3876 7306 3910
rect 6996 3842 7306 3876
rect 6996 3808 7098 3842
rect 7132 3808 7170 3842
rect 7204 3808 7306 3842
rect 6996 3774 7306 3808
rect 6996 3740 7098 3774
rect 7132 3740 7170 3774
rect 7204 3740 7306 3774
rect 6996 3706 7306 3740
rect 6996 3672 7098 3706
rect 7132 3672 7170 3706
rect 7204 3672 7306 3706
rect 6996 3638 7306 3672
rect 6996 3604 7098 3638
rect 7132 3604 7170 3638
rect 7204 3604 7306 3638
rect 6996 3570 7306 3604
rect 6996 3536 7098 3570
rect 7132 3536 7170 3570
rect 7204 3536 7306 3570
rect 6996 3502 7306 3536
rect 6996 3468 7098 3502
rect 7132 3468 7170 3502
rect 7204 3468 7306 3502
rect 6996 3434 7306 3468
rect 6996 3400 7098 3434
rect 7132 3400 7170 3434
rect 7204 3400 7306 3434
rect 6996 3366 7306 3400
rect 6996 3332 7098 3366
rect 7132 3332 7170 3366
rect 7204 3332 7306 3366
rect 6996 3298 7306 3332
rect 6996 3264 7098 3298
rect 7132 3264 7170 3298
rect 7204 3264 7306 3298
rect 6996 3230 7306 3264
rect 6996 3196 7098 3230
rect 7132 3196 7170 3230
rect 7204 3196 7306 3230
rect 6996 3162 7306 3196
rect 6996 3128 7098 3162
rect 7132 3128 7170 3162
rect 7204 3128 7306 3162
rect 6996 3058 7306 3128
rect 7426 4046 7577 4058
rect 7717 4046 7868 4058
rect 7426 4012 7528 4046
rect 7562 4012 7577 4046
rect 7717 4012 7732 4046
rect 7766 4012 7868 4046
rect 7426 3978 7577 4012
rect 7717 3978 7868 4012
rect 7426 3944 7528 3978
rect 7562 3944 7577 3978
rect 7717 3944 7732 3978
rect 7766 3944 7868 3978
rect 7426 3910 7577 3944
rect 7717 3910 7868 3944
rect 7426 3876 7528 3910
rect 7562 3876 7577 3910
rect 7717 3876 7732 3910
rect 7766 3876 7868 3910
rect 7426 3842 7577 3876
rect 7717 3842 7868 3876
rect 7426 3808 7528 3842
rect 7562 3808 7577 3842
rect 7717 3808 7732 3842
rect 7766 3808 7868 3842
rect 7426 3774 7577 3808
rect 7717 3774 7868 3808
rect 7426 3740 7528 3774
rect 7562 3740 7577 3774
rect 7717 3740 7732 3774
rect 7766 3740 7868 3774
rect 7426 3706 7577 3740
rect 7717 3706 7868 3740
rect 7426 3672 7528 3706
rect 7562 3672 7577 3706
rect 7717 3672 7732 3706
rect 7766 3672 7868 3706
rect 7426 3638 7577 3672
rect 7717 3638 7868 3672
rect 7426 3604 7528 3638
rect 7562 3604 7577 3638
rect 7717 3604 7732 3638
rect 7766 3604 7868 3638
rect 7426 3570 7577 3604
rect 7717 3570 7868 3604
rect 7426 3536 7528 3570
rect 7562 3536 7577 3570
rect 7717 3536 7732 3570
rect 7766 3536 7868 3570
rect 7426 3502 7577 3536
rect 7717 3502 7868 3536
rect 7426 3468 7528 3502
rect 7562 3468 7577 3502
rect 7717 3468 7732 3502
rect 7766 3468 7868 3502
rect 7426 3434 7577 3468
rect 7717 3434 7868 3468
rect 7426 3400 7528 3434
rect 7562 3400 7577 3434
rect 7717 3400 7732 3434
rect 7766 3400 7868 3434
rect 7426 3366 7577 3400
rect 7717 3366 7868 3400
rect 7426 3332 7528 3366
rect 7562 3332 7577 3366
rect 7717 3332 7732 3366
rect 7766 3332 7868 3366
rect 7426 3298 7577 3332
rect 7717 3298 7868 3332
rect 7426 3264 7528 3298
rect 7562 3264 7577 3298
rect 7717 3264 7732 3298
rect 7766 3264 7868 3298
rect 7426 3230 7577 3264
rect 7717 3230 7868 3264
rect 7426 3196 7528 3230
rect 7562 3196 7577 3230
rect 7717 3196 7732 3230
rect 7766 3196 7868 3230
rect 7426 3162 7577 3196
rect 7717 3162 7868 3196
rect 7426 3128 7528 3162
rect 7562 3128 7577 3162
rect 7717 3128 7732 3162
rect 7766 3128 7868 3162
rect 7426 3058 7577 3128
rect 7717 3058 7868 3128
rect 7988 4046 8298 4058
rect 7988 4012 8090 4046
rect 8124 4012 8162 4046
rect 8196 4012 8298 4046
rect 7988 3978 8298 4012
rect 7988 3944 8090 3978
rect 8124 3944 8162 3978
rect 8196 3944 8298 3978
rect 7988 3910 8298 3944
rect 7988 3876 8090 3910
rect 8124 3876 8162 3910
rect 8196 3876 8298 3910
rect 7988 3842 8298 3876
rect 7988 3808 8090 3842
rect 8124 3808 8162 3842
rect 8196 3808 8298 3842
rect 7988 3774 8298 3808
rect 7988 3740 8090 3774
rect 8124 3740 8162 3774
rect 8196 3740 8298 3774
rect 7988 3706 8298 3740
rect 7988 3672 8090 3706
rect 8124 3672 8162 3706
rect 8196 3672 8298 3706
rect 7988 3638 8298 3672
rect 7988 3604 8090 3638
rect 8124 3604 8162 3638
rect 8196 3604 8298 3638
rect 7988 3570 8298 3604
rect 7988 3536 8090 3570
rect 8124 3536 8162 3570
rect 8196 3536 8298 3570
rect 7988 3502 8298 3536
rect 7988 3468 8090 3502
rect 8124 3468 8162 3502
rect 8196 3468 8298 3502
rect 7988 3434 8298 3468
rect 7988 3400 8090 3434
rect 8124 3400 8162 3434
rect 8196 3400 8298 3434
rect 7988 3366 8298 3400
rect 7988 3332 8090 3366
rect 8124 3332 8162 3366
rect 8196 3332 8298 3366
rect 7988 3298 8298 3332
rect 7988 3264 8090 3298
rect 8124 3264 8162 3298
rect 8196 3264 8298 3298
rect 7988 3230 8298 3264
rect 7988 3196 8090 3230
rect 8124 3196 8162 3230
rect 8196 3196 8298 3230
rect 7988 3162 8298 3196
rect 7988 3128 8090 3162
rect 8124 3128 8162 3162
rect 8196 3128 8298 3162
rect 7988 3058 8298 3128
rect 8418 4046 8569 4058
rect 8709 4046 8860 4058
rect 8418 4012 8520 4046
rect 8554 4012 8569 4046
rect 8709 4012 8724 4046
rect 8758 4012 8860 4046
rect 8418 3978 8569 4012
rect 8709 3978 8860 4012
rect 8418 3944 8520 3978
rect 8554 3944 8569 3978
rect 8709 3944 8724 3978
rect 8758 3944 8860 3978
rect 8418 3910 8569 3944
rect 8709 3910 8860 3944
rect 8418 3876 8520 3910
rect 8554 3876 8569 3910
rect 8709 3876 8724 3910
rect 8758 3876 8860 3910
rect 8418 3842 8569 3876
rect 8709 3842 8860 3876
rect 8418 3808 8520 3842
rect 8554 3808 8569 3842
rect 8709 3808 8724 3842
rect 8758 3808 8860 3842
rect 8418 3774 8569 3808
rect 8709 3774 8860 3808
rect 8418 3740 8520 3774
rect 8554 3740 8569 3774
rect 8709 3740 8724 3774
rect 8758 3740 8860 3774
rect 8418 3706 8569 3740
rect 8709 3706 8860 3740
rect 8418 3672 8520 3706
rect 8554 3672 8569 3706
rect 8709 3672 8724 3706
rect 8758 3672 8860 3706
rect 8418 3638 8569 3672
rect 8709 3638 8860 3672
rect 8418 3604 8520 3638
rect 8554 3604 8569 3638
rect 8709 3604 8724 3638
rect 8758 3604 8860 3638
rect 8418 3570 8569 3604
rect 8709 3570 8860 3604
rect 8418 3536 8520 3570
rect 8554 3536 8569 3570
rect 8709 3536 8724 3570
rect 8758 3536 8860 3570
rect 8418 3502 8569 3536
rect 8709 3502 8860 3536
rect 8418 3468 8520 3502
rect 8554 3468 8569 3502
rect 8709 3468 8724 3502
rect 8758 3468 8860 3502
rect 8418 3434 8569 3468
rect 8709 3434 8860 3468
rect 8418 3400 8520 3434
rect 8554 3400 8569 3434
rect 8709 3400 8724 3434
rect 8758 3400 8860 3434
rect 8418 3366 8569 3400
rect 8709 3366 8860 3400
rect 8418 3332 8520 3366
rect 8554 3332 8569 3366
rect 8709 3332 8724 3366
rect 8758 3332 8860 3366
rect 8418 3298 8569 3332
rect 8709 3298 8860 3332
rect 8418 3264 8520 3298
rect 8554 3264 8569 3298
rect 8709 3264 8724 3298
rect 8758 3264 8860 3298
rect 8418 3230 8569 3264
rect 8709 3230 8860 3264
rect 8418 3196 8520 3230
rect 8554 3196 8569 3230
rect 8709 3196 8724 3230
rect 8758 3196 8860 3230
rect 8418 3162 8569 3196
rect 8709 3162 8860 3196
rect 8418 3128 8520 3162
rect 8554 3128 8569 3162
rect 8709 3128 8724 3162
rect 8758 3128 8860 3162
rect 8418 3058 8569 3128
rect 8709 3058 8860 3128
rect 8980 4046 9290 4058
rect 8980 4012 9082 4046
rect 9116 4012 9154 4046
rect 9188 4012 9290 4046
rect 8980 3978 9290 4012
rect 8980 3944 9082 3978
rect 9116 3944 9154 3978
rect 9188 3944 9290 3978
rect 8980 3910 9290 3944
rect 8980 3876 9082 3910
rect 9116 3876 9154 3910
rect 9188 3876 9290 3910
rect 8980 3842 9290 3876
rect 8980 3808 9082 3842
rect 9116 3808 9154 3842
rect 9188 3808 9290 3842
rect 8980 3774 9290 3808
rect 8980 3740 9082 3774
rect 9116 3740 9154 3774
rect 9188 3740 9290 3774
rect 8980 3706 9290 3740
rect 8980 3672 9082 3706
rect 9116 3672 9154 3706
rect 9188 3672 9290 3706
rect 8980 3638 9290 3672
rect 8980 3604 9082 3638
rect 9116 3604 9154 3638
rect 9188 3604 9290 3638
rect 8980 3570 9290 3604
rect 8980 3536 9082 3570
rect 9116 3536 9154 3570
rect 9188 3536 9290 3570
rect 8980 3502 9290 3536
rect 8980 3468 9082 3502
rect 9116 3468 9154 3502
rect 9188 3468 9290 3502
rect 8980 3434 9290 3468
rect 8980 3400 9082 3434
rect 9116 3400 9154 3434
rect 9188 3400 9290 3434
rect 8980 3366 9290 3400
rect 8980 3332 9082 3366
rect 9116 3332 9154 3366
rect 9188 3332 9290 3366
rect 8980 3298 9290 3332
rect 8980 3264 9082 3298
rect 9116 3264 9154 3298
rect 9188 3264 9290 3298
rect 8980 3230 9290 3264
rect 8980 3196 9082 3230
rect 9116 3196 9154 3230
rect 9188 3196 9290 3230
rect 8980 3162 9290 3196
rect 8980 3128 9082 3162
rect 9116 3128 9154 3162
rect 9188 3128 9290 3162
rect 8980 3058 9290 3128
rect 9410 4046 9561 4058
rect 9701 4046 9852 4058
rect 9410 4012 9512 4046
rect 9546 4012 9561 4046
rect 9701 4012 9716 4046
rect 9750 4012 9852 4046
rect 9410 3978 9561 4012
rect 9701 3978 9852 4012
rect 9410 3944 9512 3978
rect 9546 3944 9561 3978
rect 9701 3944 9716 3978
rect 9750 3944 9852 3978
rect 9410 3910 9561 3944
rect 9701 3910 9852 3944
rect 9410 3876 9512 3910
rect 9546 3876 9561 3910
rect 9701 3876 9716 3910
rect 9750 3876 9852 3910
rect 9410 3842 9561 3876
rect 9701 3842 9852 3876
rect 9410 3808 9512 3842
rect 9546 3808 9561 3842
rect 9701 3808 9716 3842
rect 9750 3808 9852 3842
rect 9410 3774 9561 3808
rect 9701 3774 9852 3808
rect 9410 3740 9512 3774
rect 9546 3740 9561 3774
rect 9701 3740 9716 3774
rect 9750 3740 9852 3774
rect 9410 3706 9561 3740
rect 9701 3706 9852 3740
rect 9410 3672 9512 3706
rect 9546 3672 9561 3706
rect 9701 3672 9716 3706
rect 9750 3672 9852 3706
rect 9410 3638 9561 3672
rect 9701 3638 9852 3672
rect 9410 3604 9512 3638
rect 9546 3604 9561 3638
rect 9701 3604 9716 3638
rect 9750 3604 9852 3638
rect 9410 3570 9561 3604
rect 9701 3570 9852 3604
rect 9410 3536 9512 3570
rect 9546 3536 9561 3570
rect 9701 3536 9716 3570
rect 9750 3536 9852 3570
rect 9410 3502 9561 3536
rect 9701 3502 9852 3536
rect 9410 3468 9512 3502
rect 9546 3468 9561 3502
rect 9701 3468 9716 3502
rect 9750 3468 9852 3502
rect 9410 3434 9561 3468
rect 9701 3434 9852 3468
rect 9410 3400 9512 3434
rect 9546 3400 9561 3434
rect 9701 3400 9716 3434
rect 9750 3400 9852 3434
rect 9410 3366 9561 3400
rect 9701 3366 9852 3400
rect 9410 3332 9512 3366
rect 9546 3332 9561 3366
rect 9701 3332 9716 3366
rect 9750 3332 9852 3366
rect 9410 3298 9561 3332
rect 9701 3298 9852 3332
rect 9410 3264 9512 3298
rect 9546 3264 9561 3298
rect 9701 3264 9716 3298
rect 9750 3264 9852 3298
rect 9410 3230 9561 3264
rect 9701 3230 9852 3264
rect 9410 3196 9512 3230
rect 9546 3196 9561 3230
rect 9701 3196 9716 3230
rect 9750 3196 9852 3230
rect 9410 3162 9561 3196
rect 9701 3162 9852 3196
rect 9410 3128 9512 3162
rect 9546 3128 9561 3162
rect 9701 3128 9716 3162
rect 9750 3128 9852 3162
rect 9410 3058 9561 3128
rect 9701 3058 9852 3128
rect 9972 4046 10282 4058
rect 9972 4012 10074 4046
rect 10108 4012 10146 4046
rect 10180 4012 10282 4046
rect 9972 3978 10282 4012
rect 9972 3944 10074 3978
rect 10108 3944 10146 3978
rect 10180 3944 10282 3978
rect 9972 3910 10282 3944
rect 9972 3876 10074 3910
rect 10108 3876 10146 3910
rect 10180 3876 10282 3910
rect 9972 3842 10282 3876
rect 9972 3808 10074 3842
rect 10108 3808 10146 3842
rect 10180 3808 10282 3842
rect 9972 3774 10282 3808
rect 9972 3740 10074 3774
rect 10108 3740 10146 3774
rect 10180 3740 10282 3774
rect 9972 3706 10282 3740
rect 9972 3672 10074 3706
rect 10108 3672 10146 3706
rect 10180 3672 10282 3706
rect 9972 3638 10282 3672
rect 9972 3604 10074 3638
rect 10108 3604 10146 3638
rect 10180 3604 10282 3638
rect 9972 3570 10282 3604
rect 9972 3536 10074 3570
rect 10108 3536 10146 3570
rect 10180 3536 10282 3570
rect 9972 3502 10282 3536
rect 9972 3468 10074 3502
rect 10108 3468 10146 3502
rect 10180 3468 10282 3502
rect 9972 3434 10282 3468
rect 9972 3400 10074 3434
rect 10108 3400 10146 3434
rect 10180 3400 10282 3434
rect 9972 3366 10282 3400
rect 9972 3332 10074 3366
rect 10108 3332 10146 3366
rect 10180 3332 10282 3366
rect 9972 3298 10282 3332
rect 9972 3264 10074 3298
rect 10108 3264 10146 3298
rect 10180 3264 10282 3298
rect 9972 3230 10282 3264
rect 9972 3196 10074 3230
rect 10108 3196 10146 3230
rect 10180 3196 10282 3230
rect 9972 3162 10282 3196
rect 9972 3128 10074 3162
rect 10108 3128 10146 3162
rect 10180 3128 10282 3162
rect 9972 3058 10282 3128
rect 10402 4046 10553 4058
rect 10693 4046 10844 4058
rect 10402 4012 10504 4046
rect 10538 4012 10553 4046
rect 10693 4012 10708 4046
rect 10742 4012 10844 4046
rect 10402 3978 10553 4012
rect 10693 3978 10844 4012
rect 10402 3944 10504 3978
rect 10538 3944 10553 3978
rect 10693 3944 10708 3978
rect 10742 3944 10844 3978
rect 10402 3910 10553 3944
rect 10693 3910 10844 3944
rect 10402 3876 10504 3910
rect 10538 3876 10553 3910
rect 10693 3876 10708 3910
rect 10742 3876 10844 3910
rect 10402 3842 10553 3876
rect 10693 3842 10844 3876
rect 10402 3808 10504 3842
rect 10538 3808 10553 3842
rect 10693 3808 10708 3842
rect 10742 3808 10844 3842
rect 10402 3774 10553 3808
rect 10693 3774 10844 3808
rect 10402 3740 10504 3774
rect 10538 3740 10553 3774
rect 10693 3740 10708 3774
rect 10742 3740 10844 3774
rect 10402 3706 10553 3740
rect 10693 3706 10844 3740
rect 10402 3672 10504 3706
rect 10538 3672 10553 3706
rect 10693 3672 10708 3706
rect 10742 3672 10844 3706
rect 10402 3638 10553 3672
rect 10693 3638 10844 3672
rect 10402 3604 10504 3638
rect 10538 3604 10553 3638
rect 10693 3604 10708 3638
rect 10742 3604 10844 3638
rect 10402 3570 10553 3604
rect 10693 3570 10844 3604
rect 10402 3536 10504 3570
rect 10538 3536 10553 3570
rect 10693 3536 10708 3570
rect 10742 3536 10844 3570
rect 10402 3502 10553 3536
rect 10693 3502 10844 3536
rect 10402 3468 10504 3502
rect 10538 3468 10553 3502
rect 10693 3468 10708 3502
rect 10742 3468 10844 3502
rect 10402 3434 10553 3468
rect 10693 3434 10844 3468
rect 10402 3400 10504 3434
rect 10538 3400 10553 3434
rect 10693 3400 10708 3434
rect 10742 3400 10844 3434
rect 10402 3366 10553 3400
rect 10693 3366 10844 3400
rect 10402 3332 10504 3366
rect 10538 3332 10553 3366
rect 10693 3332 10708 3366
rect 10742 3332 10844 3366
rect 10402 3298 10553 3332
rect 10693 3298 10844 3332
rect 10402 3264 10504 3298
rect 10538 3264 10553 3298
rect 10693 3264 10708 3298
rect 10742 3264 10844 3298
rect 10402 3230 10553 3264
rect 10693 3230 10844 3264
rect 10402 3196 10504 3230
rect 10538 3196 10553 3230
rect 10693 3196 10708 3230
rect 10742 3196 10844 3230
rect 10402 3162 10553 3196
rect 10693 3162 10844 3196
rect 10402 3128 10504 3162
rect 10538 3128 10553 3162
rect 10693 3128 10708 3162
rect 10742 3128 10844 3162
rect 10402 3058 10553 3128
rect 10693 3058 10844 3128
rect 10964 4046 11274 4058
rect 10964 4012 11066 4046
rect 11100 4012 11138 4046
rect 11172 4012 11274 4046
rect 10964 3978 11274 4012
rect 10964 3944 11066 3978
rect 11100 3944 11138 3978
rect 11172 3944 11274 3978
rect 10964 3910 11274 3944
rect 10964 3876 11066 3910
rect 11100 3876 11138 3910
rect 11172 3876 11274 3910
rect 10964 3842 11274 3876
rect 10964 3808 11066 3842
rect 11100 3808 11138 3842
rect 11172 3808 11274 3842
rect 10964 3774 11274 3808
rect 10964 3740 11066 3774
rect 11100 3740 11138 3774
rect 11172 3740 11274 3774
rect 10964 3706 11274 3740
rect 10964 3672 11066 3706
rect 11100 3672 11138 3706
rect 11172 3672 11274 3706
rect 10964 3638 11274 3672
rect 10964 3604 11066 3638
rect 11100 3604 11138 3638
rect 11172 3604 11274 3638
rect 10964 3570 11274 3604
rect 10964 3536 11066 3570
rect 11100 3536 11138 3570
rect 11172 3536 11274 3570
rect 10964 3502 11274 3536
rect 10964 3468 11066 3502
rect 11100 3468 11138 3502
rect 11172 3468 11274 3502
rect 10964 3434 11274 3468
rect 10964 3400 11066 3434
rect 11100 3400 11138 3434
rect 11172 3400 11274 3434
rect 10964 3366 11274 3400
rect 10964 3332 11066 3366
rect 11100 3332 11138 3366
rect 11172 3332 11274 3366
rect 10964 3298 11274 3332
rect 10964 3264 11066 3298
rect 11100 3264 11138 3298
rect 11172 3264 11274 3298
rect 10964 3230 11274 3264
rect 10964 3196 11066 3230
rect 11100 3196 11138 3230
rect 11172 3196 11274 3230
rect 10964 3162 11274 3196
rect 10964 3128 11066 3162
rect 11100 3128 11138 3162
rect 11172 3128 11274 3162
rect 10964 3058 11274 3128
rect 11394 4046 11545 4058
rect 11685 4046 11836 4058
rect 11394 4012 11496 4046
rect 11530 4012 11545 4046
rect 11685 4012 11700 4046
rect 11734 4012 11836 4046
rect 11394 3978 11545 4012
rect 11685 3978 11836 4012
rect 11394 3944 11496 3978
rect 11530 3944 11545 3978
rect 11685 3944 11700 3978
rect 11734 3944 11836 3978
rect 11394 3910 11545 3944
rect 11685 3910 11836 3944
rect 11394 3876 11496 3910
rect 11530 3876 11545 3910
rect 11685 3876 11700 3910
rect 11734 3876 11836 3910
rect 11394 3842 11545 3876
rect 11685 3842 11836 3876
rect 11394 3808 11496 3842
rect 11530 3808 11545 3842
rect 11685 3808 11700 3842
rect 11734 3808 11836 3842
rect 11394 3774 11545 3808
rect 11685 3774 11836 3808
rect 11394 3740 11496 3774
rect 11530 3740 11545 3774
rect 11685 3740 11700 3774
rect 11734 3740 11836 3774
rect 11394 3706 11545 3740
rect 11685 3706 11836 3740
rect 11394 3672 11496 3706
rect 11530 3672 11545 3706
rect 11685 3672 11700 3706
rect 11734 3672 11836 3706
rect 11394 3638 11545 3672
rect 11685 3638 11836 3672
rect 11394 3604 11496 3638
rect 11530 3604 11545 3638
rect 11685 3604 11700 3638
rect 11734 3604 11836 3638
rect 11394 3570 11545 3604
rect 11685 3570 11836 3604
rect 11394 3536 11496 3570
rect 11530 3536 11545 3570
rect 11685 3536 11700 3570
rect 11734 3536 11836 3570
rect 11394 3502 11545 3536
rect 11685 3502 11836 3536
rect 11394 3468 11496 3502
rect 11530 3468 11545 3502
rect 11685 3468 11700 3502
rect 11734 3468 11836 3502
rect 11394 3434 11545 3468
rect 11685 3434 11836 3468
rect 11394 3400 11496 3434
rect 11530 3400 11545 3434
rect 11685 3400 11700 3434
rect 11734 3400 11836 3434
rect 11394 3366 11545 3400
rect 11685 3366 11836 3400
rect 11394 3332 11496 3366
rect 11530 3332 11545 3366
rect 11685 3332 11700 3366
rect 11734 3332 11836 3366
rect 11394 3298 11545 3332
rect 11685 3298 11836 3332
rect 11394 3264 11496 3298
rect 11530 3264 11545 3298
rect 11685 3264 11700 3298
rect 11734 3264 11836 3298
rect 11394 3230 11545 3264
rect 11685 3230 11836 3264
rect 11394 3196 11496 3230
rect 11530 3196 11545 3230
rect 11685 3196 11700 3230
rect 11734 3196 11836 3230
rect 11394 3162 11545 3196
rect 11685 3162 11836 3196
rect 11394 3128 11496 3162
rect 11530 3128 11545 3162
rect 11685 3128 11700 3162
rect 11734 3128 11836 3162
rect 11394 3058 11545 3128
rect 11685 3058 11836 3128
rect 11956 4046 12266 4058
rect 11956 4012 12058 4046
rect 12092 4012 12130 4046
rect 12164 4012 12266 4046
rect 11956 3978 12266 4012
rect 11956 3944 12058 3978
rect 12092 3944 12130 3978
rect 12164 3944 12266 3978
rect 11956 3910 12266 3944
rect 11956 3876 12058 3910
rect 12092 3876 12130 3910
rect 12164 3876 12266 3910
rect 11956 3842 12266 3876
rect 11956 3808 12058 3842
rect 12092 3808 12130 3842
rect 12164 3808 12266 3842
rect 11956 3774 12266 3808
rect 11956 3740 12058 3774
rect 12092 3740 12130 3774
rect 12164 3740 12266 3774
rect 11956 3706 12266 3740
rect 11956 3672 12058 3706
rect 12092 3672 12130 3706
rect 12164 3672 12266 3706
rect 11956 3638 12266 3672
rect 11956 3604 12058 3638
rect 12092 3604 12130 3638
rect 12164 3604 12266 3638
rect 11956 3570 12266 3604
rect 11956 3536 12058 3570
rect 12092 3536 12130 3570
rect 12164 3536 12266 3570
rect 11956 3502 12266 3536
rect 11956 3468 12058 3502
rect 12092 3468 12130 3502
rect 12164 3468 12266 3502
rect 11956 3434 12266 3468
rect 11956 3400 12058 3434
rect 12092 3400 12130 3434
rect 12164 3400 12266 3434
rect 11956 3366 12266 3400
rect 11956 3332 12058 3366
rect 12092 3332 12130 3366
rect 12164 3332 12266 3366
rect 11956 3298 12266 3332
rect 11956 3264 12058 3298
rect 12092 3264 12130 3298
rect 12164 3264 12266 3298
rect 11956 3230 12266 3264
rect 11956 3196 12058 3230
rect 12092 3196 12130 3230
rect 12164 3196 12266 3230
rect 11956 3162 12266 3196
rect 11956 3128 12058 3162
rect 12092 3128 12130 3162
rect 12164 3128 12266 3162
rect 11956 3058 12266 3128
rect 12386 4046 12537 4058
rect 12677 4046 12828 4058
rect 12386 4012 12488 4046
rect 12522 4012 12537 4046
rect 12677 4012 12692 4046
rect 12726 4012 12828 4046
rect 12386 3978 12537 4012
rect 12677 3978 12828 4012
rect 12386 3944 12488 3978
rect 12522 3944 12537 3978
rect 12677 3944 12692 3978
rect 12726 3944 12828 3978
rect 12386 3910 12537 3944
rect 12677 3910 12828 3944
rect 12386 3876 12488 3910
rect 12522 3876 12537 3910
rect 12677 3876 12692 3910
rect 12726 3876 12828 3910
rect 12386 3842 12537 3876
rect 12677 3842 12828 3876
rect 12386 3808 12488 3842
rect 12522 3808 12537 3842
rect 12677 3808 12692 3842
rect 12726 3808 12828 3842
rect 12386 3774 12537 3808
rect 12677 3774 12828 3808
rect 12386 3740 12488 3774
rect 12522 3740 12537 3774
rect 12677 3740 12692 3774
rect 12726 3740 12828 3774
rect 12386 3706 12537 3740
rect 12677 3706 12828 3740
rect 12386 3672 12488 3706
rect 12522 3672 12537 3706
rect 12677 3672 12692 3706
rect 12726 3672 12828 3706
rect 12386 3638 12537 3672
rect 12677 3638 12828 3672
rect 12386 3604 12488 3638
rect 12522 3604 12537 3638
rect 12677 3604 12692 3638
rect 12726 3604 12828 3638
rect 12386 3570 12537 3604
rect 12677 3570 12828 3604
rect 12386 3536 12488 3570
rect 12522 3536 12537 3570
rect 12677 3536 12692 3570
rect 12726 3536 12828 3570
rect 12386 3502 12537 3536
rect 12677 3502 12828 3536
rect 12386 3468 12488 3502
rect 12522 3468 12537 3502
rect 12677 3468 12692 3502
rect 12726 3468 12828 3502
rect 12386 3434 12537 3468
rect 12677 3434 12828 3468
rect 12386 3400 12488 3434
rect 12522 3400 12537 3434
rect 12677 3400 12692 3434
rect 12726 3400 12828 3434
rect 12386 3366 12537 3400
rect 12677 3366 12828 3400
rect 12386 3332 12488 3366
rect 12522 3332 12537 3366
rect 12677 3332 12692 3366
rect 12726 3332 12828 3366
rect 12386 3298 12537 3332
rect 12677 3298 12828 3332
rect 12386 3264 12488 3298
rect 12522 3264 12537 3298
rect 12677 3264 12692 3298
rect 12726 3264 12828 3298
rect 12386 3230 12537 3264
rect 12677 3230 12828 3264
rect 12386 3196 12488 3230
rect 12522 3196 12537 3230
rect 12677 3196 12692 3230
rect 12726 3196 12828 3230
rect 12386 3162 12537 3196
rect 12677 3162 12828 3196
rect 12386 3128 12488 3162
rect 12522 3128 12537 3162
rect 12677 3128 12692 3162
rect 12726 3128 12828 3162
rect 12386 3058 12537 3128
rect 12677 3058 12828 3128
rect 12948 4046 13258 4058
rect 12948 4012 13050 4046
rect 13084 4012 13122 4046
rect 13156 4012 13258 4046
rect 12948 3978 13258 4012
rect 12948 3944 13050 3978
rect 13084 3944 13122 3978
rect 13156 3944 13258 3978
rect 12948 3910 13258 3944
rect 12948 3876 13050 3910
rect 13084 3876 13122 3910
rect 13156 3876 13258 3910
rect 12948 3842 13258 3876
rect 12948 3808 13050 3842
rect 13084 3808 13122 3842
rect 13156 3808 13258 3842
rect 12948 3774 13258 3808
rect 12948 3740 13050 3774
rect 13084 3740 13122 3774
rect 13156 3740 13258 3774
rect 12948 3706 13258 3740
rect 12948 3672 13050 3706
rect 13084 3672 13122 3706
rect 13156 3672 13258 3706
rect 12948 3638 13258 3672
rect 12948 3604 13050 3638
rect 13084 3604 13122 3638
rect 13156 3604 13258 3638
rect 12948 3570 13258 3604
rect 12948 3536 13050 3570
rect 13084 3536 13122 3570
rect 13156 3536 13258 3570
rect 12948 3502 13258 3536
rect 12948 3468 13050 3502
rect 13084 3468 13122 3502
rect 13156 3468 13258 3502
rect 12948 3434 13258 3468
rect 12948 3400 13050 3434
rect 13084 3400 13122 3434
rect 13156 3400 13258 3434
rect 12948 3366 13258 3400
rect 12948 3332 13050 3366
rect 13084 3332 13122 3366
rect 13156 3332 13258 3366
rect 12948 3298 13258 3332
rect 12948 3264 13050 3298
rect 13084 3264 13122 3298
rect 13156 3264 13258 3298
rect 12948 3230 13258 3264
rect 12948 3196 13050 3230
rect 13084 3196 13122 3230
rect 13156 3196 13258 3230
rect 12948 3162 13258 3196
rect 12948 3128 13050 3162
rect 13084 3128 13122 3162
rect 13156 3128 13258 3162
rect 12948 3058 13258 3128
rect 13378 4046 13529 4058
rect 13669 4046 13820 4058
rect 13378 4012 13480 4046
rect 13514 4012 13529 4046
rect 13669 4012 13684 4046
rect 13718 4012 13820 4046
rect 13378 3978 13529 4012
rect 13669 3978 13820 4012
rect 13378 3944 13480 3978
rect 13514 3944 13529 3978
rect 13669 3944 13684 3978
rect 13718 3944 13820 3978
rect 13378 3910 13529 3944
rect 13669 3910 13820 3944
rect 13378 3876 13480 3910
rect 13514 3876 13529 3910
rect 13669 3876 13684 3910
rect 13718 3876 13820 3910
rect 13378 3842 13529 3876
rect 13669 3842 13820 3876
rect 13378 3808 13480 3842
rect 13514 3808 13529 3842
rect 13669 3808 13684 3842
rect 13718 3808 13820 3842
rect 13378 3774 13529 3808
rect 13669 3774 13820 3808
rect 13378 3740 13480 3774
rect 13514 3740 13529 3774
rect 13669 3740 13684 3774
rect 13718 3740 13820 3774
rect 13378 3706 13529 3740
rect 13669 3706 13820 3740
rect 13378 3672 13480 3706
rect 13514 3672 13529 3706
rect 13669 3672 13684 3706
rect 13718 3672 13820 3706
rect 13378 3638 13529 3672
rect 13669 3638 13820 3672
rect 13378 3604 13480 3638
rect 13514 3604 13529 3638
rect 13669 3604 13684 3638
rect 13718 3604 13820 3638
rect 13378 3570 13529 3604
rect 13669 3570 13820 3604
rect 13378 3536 13480 3570
rect 13514 3536 13529 3570
rect 13669 3536 13684 3570
rect 13718 3536 13820 3570
rect 13378 3502 13529 3536
rect 13669 3502 13820 3536
rect 13378 3468 13480 3502
rect 13514 3468 13529 3502
rect 13669 3468 13684 3502
rect 13718 3468 13820 3502
rect 13378 3434 13529 3468
rect 13669 3434 13820 3468
rect 13378 3400 13480 3434
rect 13514 3400 13529 3434
rect 13669 3400 13684 3434
rect 13718 3400 13820 3434
rect 13378 3366 13529 3400
rect 13669 3366 13820 3400
rect 13378 3332 13480 3366
rect 13514 3332 13529 3366
rect 13669 3332 13684 3366
rect 13718 3332 13820 3366
rect 13378 3298 13529 3332
rect 13669 3298 13820 3332
rect 13378 3264 13480 3298
rect 13514 3264 13529 3298
rect 13669 3264 13684 3298
rect 13718 3264 13820 3298
rect 13378 3230 13529 3264
rect 13669 3230 13820 3264
rect 13378 3196 13480 3230
rect 13514 3196 13529 3230
rect 13669 3196 13684 3230
rect 13718 3196 13820 3230
rect 13378 3162 13529 3196
rect 13669 3162 13820 3196
rect 13378 3128 13480 3162
rect 13514 3128 13529 3162
rect 13669 3128 13684 3162
rect 13718 3128 13820 3162
rect 13378 3058 13529 3128
rect 13669 3058 13820 3128
rect 13940 4046 14178 4058
rect 13940 4012 14042 4046
rect 14076 4012 14178 4046
rect 13940 3978 14178 4012
rect 13940 3944 14042 3978
rect 14076 3944 14178 3978
rect 13940 3910 14178 3944
rect 13940 3876 14042 3910
rect 14076 3876 14178 3910
rect 13940 3842 14178 3876
rect 13940 3808 14042 3842
rect 14076 3808 14178 3842
rect 13940 3774 14178 3808
rect 13940 3740 14042 3774
rect 14076 3740 14178 3774
rect 13940 3706 14178 3740
rect 13940 3672 14042 3706
rect 14076 3672 14178 3706
rect 13940 3638 14178 3672
rect 13940 3604 14042 3638
rect 14076 3604 14178 3638
rect 13940 3570 14178 3604
rect 13940 3536 14042 3570
rect 14076 3536 14178 3570
rect 13940 3502 14178 3536
rect 13940 3468 14042 3502
rect 14076 3468 14178 3502
rect 13940 3434 14178 3468
rect 13940 3400 14042 3434
rect 14076 3400 14178 3434
rect 13940 3366 14178 3400
rect 13940 3332 14042 3366
rect 14076 3332 14178 3366
rect 13940 3298 14178 3332
rect 13940 3264 14042 3298
rect 14076 3264 14178 3298
rect 13940 3230 14178 3264
rect 13940 3196 14042 3230
rect 14076 3196 14178 3230
rect 13940 3162 14178 3196
rect 13940 3128 14042 3162
rect 14076 3128 14178 3162
rect 13940 3058 14178 3128
rect 14298 4046 14435 4058
rect 14298 4012 14386 4046
rect 14420 4012 14435 4046
rect 14298 3978 14435 4012
rect 14298 3944 14386 3978
rect 14420 3944 14435 3978
rect 14298 3910 14435 3944
rect 14298 3876 14386 3910
rect 14420 3876 14435 3910
rect 14298 3842 14435 3876
rect 14298 3808 14386 3842
rect 14420 3808 14435 3842
rect 14298 3774 14435 3808
rect 14298 3740 14386 3774
rect 14420 3740 14435 3774
rect 14298 3706 14435 3740
rect 14298 3672 14386 3706
rect 14420 3672 14435 3706
rect 14298 3638 14435 3672
rect 14298 3604 14386 3638
rect 14420 3604 14435 3638
rect 14298 3570 14435 3604
rect 14298 3536 14386 3570
rect 14420 3536 14435 3570
rect 14298 3502 14435 3536
rect 14298 3468 14386 3502
rect 14420 3468 14435 3502
rect 14298 3434 14435 3468
rect 14298 3400 14386 3434
rect 14420 3400 14435 3434
rect 14298 3366 14435 3400
rect 14298 3332 14386 3366
rect 14420 3332 14435 3366
rect 14298 3298 14435 3332
rect 14298 3264 14386 3298
rect 14420 3264 14435 3298
rect 14298 3230 14435 3264
rect 14298 3196 14386 3230
rect 14420 3196 14435 3230
rect 14298 3162 14435 3196
rect 14298 3128 14386 3162
rect 14420 3128 14435 3162
rect 14298 3058 14435 3128
rect 787 2445 924 2457
rect 787 2411 802 2445
rect 836 2411 924 2445
rect 787 2377 924 2411
rect 787 2343 802 2377
rect 836 2343 924 2377
rect 787 2309 924 2343
rect 787 2275 802 2309
rect 836 2275 924 2309
rect 787 2241 924 2275
rect 787 2207 802 2241
rect 836 2207 924 2241
rect 787 2173 924 2207
rect 787 2139 802 2173
rect 836 2139 924 2173
rect 787 2105 924 2139
rect 787 2071 802 2105
rect 836 2071 924 2105
rect 787 2037 924 2071
rect 787 2003 802 2037
rect 836 2003 924 2037
rect 787 1969 924 2003
rect 787 1935 802 1969
rect 836 1935 924 1969
rect 787 1901 924 1935
rect 787 1867 802 1901
rect 836 1867 924 1901
rect 787 1833 924 1867
rect 787 1799 802 1833
rect 836 1799 924 1833
rect 787 1765 924 1799
rect 787 1731 802 1765
rect 836 1731 924 1765
rect 787 1697 924 1731
rect 787 1663 802 1697
rect 836 1663 924 1697
rect 787 1629 924 1663
rect 787 1595 802 1629
rect 836 1595 924 1629
rect 787 1561 924 1595
rect 787 1527 802 1561
rect 836 1527 924 1561
rect 787 1457 924 1527
rect 1044 2445 1354 2457
rect 1044 2411 1146 2445
rect 1180 2411 1218 2445
rect 1252 2411 1354 2445
rect 1044 2377 1354 2411
rect 1044 2343 1146 2377
rect 1180 2343 1218 2377
rect 1252 2343 1354 2377
rect 1044 2309 1354 2343
rect 1044 2275 1146 2309
rect 1180 2275 1218 2309
rect 1252 2275 1354 2309
rect 1044 2241 1354 2275
rect 1044 2207 1146 2241
rect 1180 2207 1218 2241
rect 1252 2207 1354 2241
rect 1044 2173 1354 2207
rect 1044 2139 1146 2173
rect 1180 2139 1218 2173
rect 1252 2139 1354 2173
rect 1044 2105 1354 2139
rect 1044 2071 1146 2105
rect 1180 2071 1218 2105
rect 1252 2071 1354 2105
rect 1044 2037 1354 2071
rect 1044 2003 1146 2037
rect 1180 2003 1218 2037
rect 1252 2003 1354 2037
rect 1044 1969 1354 2003
rect 1044 1935 1146 1969
rect 1180 1935 1218 1969
rect 1252 1935 1354 1969
rect 1044 1901 1354 1935
rect 1044 1867 1146 1901
rect 1180 1867 1218 1901
rect 1252 1867 1354 1901
rect 1044 1833 1354 1867
rect 1044 1799 1146 1833
rect 1180 1799 1218 1833
rect 1252 1799 1354 1833
rect 1044 1765 1354 1799
rect 1044 1731 1146 1765
rect 1180 1731 1218 1765
rect 1252 1731 1354 1765
rect 1044 1697 1354 1731
rect 1044 1663 1146 1697
rect 1180 1663 1218 1697
rect 1252 1663 1354 1697
rect 1044 1629 1354 1663
rect 1044 1595 1146 1629
rect 1180 1595 1218 1629
rect 1252 1595 1354 1629
rect 1044 1561 1354 1595
rect 1044 1527 1146 1561
rect 1180 1527 1218 1561
rect 1252 1527 1354 1561
rect 1044 1457 1354 1527
rect 1474 2445 1625 2457
rect 1765 2445 1916 2457
rect 1474 2411 1576 2445
rect 1610 2411 1625 2445
rect 1765 2411 1780 2445
rect 1814 2411 1916 2445
rect 1474 2377 1625 2411
rect 1765 2377 1916 2411
rect 1474 2343 1576 2377
rect 1610 2343 1625 2377
rect 1765 2343 1780 2377
rect 1814 2343 1916 2377
rect 1474 2309 1625 2343
rect 1765 2309 1916 2343
rect 1474 2275 1576 2309
rect 1610 2275 1625 2309
rect 1765 2275 1780 2309
rect 1814 2275 1916 2309
rect 1474 2241 1625 2275
rect 1765 2241 1916 2275
rect 1474 2207 1576 2241
rect 1610 2207 1625 2241
rect 1765 2207 1780 2241
rect 1814 2207 1916 2241
rect 1474 2173 1625 2207
rect 1765 2173 1916 2207
rect 1474 2139 1576 2173
rect 1610 2139 1625 2173
rect 1765 2139 1780 2173
rect 1814 2139 1916 2173
rect 1474 2105 1625 2139
rect 1765 2105 1916 2139
rect 1474 2071 1576 2105
rect 1610 2071 1625 2105
rect 1765 2071 1780 2105
rect 1814 2071 1916 2105
rect 1474 2037 1625 2071
rect 1765 2037 1916 2071
rect 1474 2003 1576 2037
rect 1610 2003 1625 2037
rect 1765 2003 1780 2037
rect 1814 2003 1916 2037
rect 1474 1969 1625 2003
rect 1765 1969 1916 2003
rect 1474 1935 1576 1969
rect 1610 1935 1625 1969
rect 1765 1935 1780 1969
rect 1814 1935 1916 1969
rect 1474 1901 1625 1935
rect 1765 1901 1916 1935
rect 1474 1867 1576 1901
rect 1610 1867 1625 1901
rect 1765 1867 1780 1901
rect 1814 1867 1916 1901
rect 1474 1833 1625 1867
rect 1765 1833 1916 1867
rect 1474 1799 1576 1833
rect 1610 1799 1625 1833
rect 1765 1799 1780 1833
rect 1814 1799 1916 1833
rect 1474 1765 1625 1799
rect 1765 1765 1916 1799
rect 1474 1731 1576 1765
rect 1610 1731 1625 1765
rect 1765 1731 1780 1765
rect 1814 1731 1916 1765
rect 1474 1697 1625 1731
rect 1765 1697 1916 1731
rect 1474 1663 1576 1697
rect 1610 1663 1625 1697
rect 1765 1663 1780 1697
rect 1814 1663 1916 1697
rect 1474 1629 1625 1663
rect 1765 1629 1916 1663
rect 1474 1595 1576 1629
rect 1610 1595 1625 1629
rect 1765 1595 1780 1629
rect 1814 1595 1916 1629
rect 1474 1561 1625 1595
rect 1765 1561 1916 1595
rect 1474 1527 1576 1561
rect 1610 1527 1625 1561
rect 1765 1527 1780 1561
rect 1814 1527 1916 1561
rect 1474 1457 1625 1527
rect 1765 1457 1916 1527
rect 2036 2445 2346 2457
rect 2036 2411 2138 2445
rect 2172 2411 2210 2445
rect 2244 2411 2346 2445
rect 2036 2377 2346 2411
rect 2036 2343 2138 2377
rect 2172 2343 2210 2377
rect 2244 2343 2346 2377
rect 2036 2309 2346 2343
rect 2036 2275 2138 2309
rect 2172 2275 2210 2309
rect 2244 2275 2346 2309
rect 2036 2241 2346 2275
rect 2036 2207 2138 2241
rect 2172 2207 2210 2241
rect 2244 2207 2346 2241
rect 2036 2173 2346 2207
rect 2036 2139 2138 2173
rect 2172 2139 2210 2173
rect 2244 2139 2346 2173
rect 2036 2105 2346 2139
rect 2036 2071 2138 2105
rect 2172 2071 2210 2105
rect 2244 2071 2346 2105
rect 2036 2037 2346 2071
rect 2036 2003 2138 2037
rect 2172 2003 2210 2037
rect 2244 2003 2346 2037
rect 2036 1969 2346 2003
rect 2036 1935 2138 1969
rect 2172 1935 2210 1969
rect 2244 1935 2346 1969
rect 2036 1901 2346 1935
rect 2036 1867 2138 1901
rect 2172 1867 2210 1901
rect 2244 1867 2346 1901
rect 2036 1833 2346 1867
rect 2036 1799 2138 1833
rect 2172 1799 2210 1833
rect 2244 1799 2346 1833
rect 2036 1765 2346 1799
rect 2036 1731 2138 1765
rect 2172 1731 2210 1765
rect 2244 1731 2346 1765
rect 2036 1697 2346 1731
rect 2036 1663 2138 1697
rect 2172 1663 2210 1697
rect 2244 1663 2346 1697
rect 2036 1629 2346 1663
rect 2036 1595 2138 1629
rect 2172 1595 2210 1629
rect 2244 1595 2346 1629
rect 2036 1561 2346 1595
rect 2036 1527 2138 1561
rect 2172 1527 2210 1561
rect 2244 1527 2346 1561
rect 2036 1457 2346 1527
rect 2466 2445 2617 2457
rect 2757 2445 2908 2457
rect 2466 2411 2568 2445
rect 2602 2411 2617 2445
rect 2757 2411 2772 2445
rect 2806 2411 2908 2445
rect 2466 2377 2617 2411
rect 2757 2377 2908 2411
rect 2466 2343 2568 2377
rect 2602 2343 2617 2377
rect 2757 2343 2772 2377
rect 2806 2343 2908 2377
rect 2466 2309 2617 2343
rect 2757 2309 2908 2343
rect 2466 2275 2568 2309
rect 2602 2275 2617 2309
rect 2757 2275 2772 2309
rect 2806 2275 2908 2309
rect 2466 2241 2617 2275
rect 2757 2241 2908 2275
rect 2466 2207 2568 2241
rect 2602 2207 2617 2241
rect 2757 2207 2772 2241
rect 2806 2207 2908 2241
rect 2466 2173 2617 2207
rect 2757 2173 2908 2207
rect 2466 2139 2568 2173
rect 2602 2139 2617 2173
rect 2757 2139 2772 2173
rect 2806 2139 2908 2173
rect 2466 2105 2617 2139
rect 2757 2105 2908 2139
rect 2466 2071 2568 2105
rect 2602 2071 2617 2105
rect 2757 2071 2772 2105
rect 2806 2071 2908 2105
rect 2466 2037 2617 2071
rect 2757 2037 2908 2071
rect 2466 2003 2568 2037
rect 2602 2003 2617 2037
rect 2757 2003 2772 2037
rect 2806 2003 2908 2037
rect 2466 1969 2617 2003
rect 2757 1969 2908 2003
rect 2466 1935 2568 1969
rect 2602 1935 2617 1969
rect 2757 1935 2772 1969
rect 2806 1935 2908 1969
rect 2466 1901 2617 1935
rect 2757 1901 2908 1935
rect 2466 1867 2568 1901
rect 2602 1867 2617 1901
rect 2757 1867 2772 1901
rect 2806 1867 2908 1901
rect 2466 1833 2617 1867
rect 2757 1833 2908 1867
rect 2466 1799 2568 1833
rect 2602 1799 2617 1833
rect 2757 1799 2772 1833
rect 2806 1799 2908 1833
rect 2466 1765 2617 1799
rect 2757 1765 2908 1799
rect 2466 1731 2568 1765
rect 2602 1731 2617 1765
rect 2757 1731 2772 1765
rect 2806 1731 2908 1765
rect 2466 1697 2617 1731
rect 2757 1697 2908 1731
rect 2466 1663 2568 1697
rect 2602 1663 2617 1697
rect 2757 1663 2772 1697
rect 2806 1663 2908 1697
rect 2466 1629 2617 1663
rect 2757 1629 2908 1663
rect 2466 1595 2568 1629
rect 2602 1595 2617 1629
rect 2757 1595 2772 1629
rect 2806 1595 2908 1629
rect 2466 1561 2617 1595
rect 2757 1561 2908 1595
rect 2466 1527 2568 1561
rect 2602 1527 2617 1561
rect 2757 1527 2772 1561
rect 2806 1527 2908 1561
rect 2466 1457 2617 1527
rect 2757 1457 2908 1527
rect 3028 2445 3338 2457
rect 3028 2411 3130 2445
rect 3164 2411 3202 2445
rect 3236 2411 3338 2445
rect 3028 2377 3338 2411
rect 3028 2343 3130 2377
rect 3164 2343 3202 2377
rect 3236 2343 3338 2377
rect 3028 2309 3338 2343
rect 3028 2275 3130 2309
rect 3164 2275 3202 2309
rect 3236 2275 3338 2309
rect 3028 2241 3338 2275
rect 3028 2207 3130 2241
rect 3164 2207 3202 2241
rect 3236 2207 3338 2241
rect 3028 2173 3338 2207
rect 3028 2139 3130 2173
rect 3164 2139 3202 2173
rect 3236 2139 3338 2173
rect 3028 2105 3338 2139
rect 3028 2071 3130 2105
rect 3164 2071 3202 2105
rect 3236 2071 3338 2105
rect 3028 2037 3338 2071
rect 3028 2003 3130 2037
rect 3164 2003 3202 2037
rect 3236 2003 3338 2037
rect 3028 1969 3338 2003
rect 3028 1935 3130 1969
rect 3164 1935 3202 1969
rect 3236 1935 3338 1969
rect 3028 1901 3338 1935
rect 3028 1867 3130 1901
rect 3164 1867 3202 1901
rect 3236 1867 3338 1901
rect 3028 1833 3338 1867
rect 3028 1799 3130 1833
rect 3164 1799 3202 1833
rect 3236 1799 3338 1833
rect 3028 1765 3338 1799
rect 3028 1731 3130 1765
rect 3164 1731 3202 1765
rect 3236 1731 3338 1765
rect 3028 1697 3338 1731
rect 3028 1663 3130 1697
rect 3164 1663 3202 1697
rect 3236 1663 3338 1697
rect 3028 1629 3338 1663
rect 3028 1595 3130 1629
rect 3164 1595 3202 1629
rect 3236 1595 3338 1629
rect 3028 1561 3338 1595
rect 3028 1527 3130 1561
rect 3164 1527 3202 1561
rect 3236 1527 3338 1561
rect 3028 1457 3338 1527
rect 3458 2445 3609 2457
rect 3749 2445 3900 2457
rect 3458 2411 3560 2445
rect 3594 2411 3609 2445
rect 3749 2411 3764 2445
rect 3798 2411 3900 2445
rect 3458 2377 3609 2411
rect 3749 2377 3900 2411
rect 3458 2343 3560 2377
rect 3594 2343 3609 2377
rect 3749 2343 3764 2377
rect 3798 2343 3900 2377
rect 3458 2309 3609 2343
rect 3749 2309 3900 2343
rect 3458 2275 3560 2309
rect 3594 2275 3609 2309
rect 3749 2275 3764 2309
rect 3798 2275 3900 2309
rect 3458 2241 3609 2275
rect 3749 2241 3900 2275
rect 3458 2207 3560 2241
rect 3594 2207 3609 2241
rect 3749 2207 3764 2241
rect 3798 2207 3900 2241
rect 3458 2173 3609 2207
rect 3749 2173 3900 2207
rect 3458 2139 3560 2173
rect 3594 2139 3609 2173
rect 3749 2139 3764 2173
rect 3798 2139 3900 2173
rect 3458 2105 3609 2139
rect 3749 2105 3900 2139
rect 3458 2071 3560 2105
rect 3594 2071 3609 2105
rect 3749 2071 3764 2105
rect 3798 2071 3900 2105
rect 3458 2037 3609 2071
rect 3749 2037 3900 2071
rect 3458 2003 3560 2037
rect 3594 2003 3609 2037
rect 3749 2003 3764 2037
rect 3798 2003 3900 2037
rect 3458 1969 3609 2003
rect 3749 1969 3900 2003
rect 3458 1935 3560 1969
rect 3594 1935 3609 1969
rect 3749 1935 3764 1969
rect 3798 1935 3900 1969
rect 3458 1901 3609 1935
rect 3749 1901 3900 1935
rect 3458 1867 3560 1901
rect 3594 1867 3609 1901
rect 3749 1867 3764 1901
rect 3798 1867 3900 1901
rect 3458 1833 3609 1867
rect 3749 1833 3900 1867
rect 3458 1799 3560 1833
rect 3594 1799 3609 1833
rect 3749 1799 3764 1833
rect 3798 1799 3900 1833
rect 3458 1765 3609 1799
rect 3749 1765 3900 1799
rect 3458 1731 3560 1765
rect 3594 1731 3609 1765
rect 3749 1731 3764 1765
rect 3798 1731 3900 1765
rect 3458 1697 3609 1731
rect 3749 1697 3900 1731
rect 3458 1663 3560 1697
rect 3594 1663 3609 1697
rect 3749 1663 3764 1697
rect 3798 1663 3900 1697
rect 3458 1629 3609 1663
rect 3749 1629 3900 1663
rect 3458 1595 3560 1629
rect 3594 1595 3609 1629
rect 3749 1595 3764 1629
rect 3798 1595 3900 1629
rect 3458 1561 3609 1595
rect 3749 1561 3900 1595
rect 3458 1527 3560 1561
rect 3594 1527 3609 1561
rect 3749 1527 3764 1561
rect 3798 1527 3900 1561
rect 3458 1457 3609 1527
rect 3749 1457 3900 1527
rect 4020 2445 4330 2457
rect 4020 2411 4122 2445
rect 4156 2411 4194 2445
rect 4228 2411 4330 2445
rect 4020 2377 4330 2411
rect 4020 2343 4122 2377
rect 4156 2343 4194 2377
rect 4228 2343 4330 2377
rect 4020 2309 4330 2343
rect 4020 2275 4122 2309
rect 4156 2275 4194 2309
rect 4228 2275 4330 2309
rect 4020 2241 4330 2275
rect 4020 2207 4122 2241
rect 4156 2207 4194 2241
rect 4228 2207 4330 2241
rect 4020 2173 4330 2207
rect 4020 2139 4122 2173
rect 4156 2139 4194 2173
rect 4228 2139 4330 2173
rect 4020 2105 4330 2139
rect 4020 2071 4122 2105
rect 4156 2071 4194 2105
rect 4228 2071 4330 2105
rect 4020 2037 4330 2071
rect 4020 2003 4122 2037
rect 4156 2003 4194 2037
rect 4228 2003 4330 2037
rect 4020 1969 4330 2003
rect 4020 1935 4122 1969
rect 4156 1935 4194 1969
rect 4228 1935 4330 1969
rect 4020 1901 4330 1935
rect 4020 1867 4122 1901
rect 4156 1867 4194 1901
rect 4228 1867 4330 1901
rect 4020 1833 4330 1867
rect 4020 1799 4122 1833
rect 4156 1799 4194 1833
rect 4228 1799 4330 1833
rect 4020 1765 4330 1799
rect 4020 1731 4122 1765
rect 4156 1731 4194 1765
rect 4228 1731 4330 1765
rect 4020 1697 4330 1731
rect 4020 1663 4122 1697
rect 4156 1663 4194 1697
rect 4228 1663 4330 1697
rect 4020 1629 4330 1663
rect 4020 1595 4122 1629
rect 4156 1595 4194 1629
rect 4228 1595 4330 1629
rect 4020 1561 4330 1595
rect 4020 1527 4122 1561
rect 4156 1527 4194 1561
rect 4228 1527 4330 1561
rect 4020 1457 4330 1527
rect 4450 2445 4601 2457
rect 4741 2445 4892 2457
rect 4450 2411 4552 2445
rect 4586 2411 4601 2445
rect 4741 2411 4756 2445
rect 4790 2411 4892 2445
rect 4450 2377 4601 2411
rect 4741 2377 4892 2411
rect 4450 2343 4552 2377
rect 4586 2343 4601 2377
rect 4741 2343 4756 2377
rect 4790 2343 4892 2377
rect 4450 2309 4601 2343
rect 4741 2309 4892 2343
rect 4450 2275 4552 2309
rect 4586 2275 4601 2309
rect 4741 2275 4756 2309
rect 4790 2275 4892 2309
rect 4450 2241 4601 2275
rect 4741 2241 4892 2275
rect 4450 2207 4552 2241
rect 4586 2207 4601 2241
rect 4741 2207 4756 2241
rect 4790 2207 4892 2241
rect 4450 2173 4601 2207
rect 4741 2173 4892 2207
rect 4450 2139 4552 2173
rect 4586 2139 4601 2173
rect 4741 2139 4756 2173
rect 4790 2139 4892 2173
rect 4450 2105 4601 2139
rect 4741 2105 4892 2139
rect 4450 2071 4552 2105
rect 4586 2071 4601 2105
rect 4741 2071 4756 2105
rect 4790 2071 4892 2105
rect 4450 2037 4601 2071
rect 4741 2037 4892 2071
rect 4450 2003 4552 2037
rect 4586 2003 4601 2037
rect 4741 2003 4756 2037
rect 4790 2003 4892 2037
rect 4450 1969 4601 2003
rect 4741 1969 4892 2003
rect 4450 1935 4552 1969
rect 4586 1935 4601 1969
rect 4741 1935 4756 1969
rect 4790 1935 4892 1969
rect 4450 1901 4601 1935
rect 4741 1901 4892 1935
rect 4450 1867 4552 1901
rect 4586 1867 4601 1901
rect 4741 1867 4756 1901
rect 4790 1867 4892 1901
rect 4450 1833 4601 1867
rect 4741 1833 4892 1867
rect 4450 1799 4552 1833
rect 4586 1799 4601 1833
rect 4741 1799 4756 1833
rect 4790 1799 4892 1833
rect 4450 1765 4601 1799
rect 4741 1765 4892 1799
rect 4450 1731 4552 1765
rect 4586 1731 4601 1765
rect 4741 1731 4756 1765
rect 4790 1731 4892 1765
rect 4450 1697 4601 1731
rect 4741 1697 4892 1731
rect 4450 1663 4552 1697
rect 4586 1663 4601 1697
rect 4741 1663 4756 1697
rect 4790 1663 4892 1697
rect 4450 1629 4601 1663
rect 4741 1629 4892 1663
rect 4450 1595 4552 1629
rect 4586 1595 4601 1629
rect 4741 1595 4756 1629
rect 4790 1595 4892 1629
rect 4450 1561 4601 1595
rect 4741 1561 4892 1595
rect 4450 1527 4552 1561
rect 4586 1527 4601 1561
rect 4741 1527 4756 1561
rect 4790 1527 4892 1561
rect 4450 1457 4601 1527
rect 4741 1457 4892 1527
rect 5012 2445 5322 2457
rect 5012 2411 5114 2445
rect 5148 2411 5186 2445
rect 5220 2411 5322 2445
rect 5012 2377 5322 2411
rect 5012 2343 5114 2377
rect 5148 2343 5186 2377
rect 5220 2343 5322 2377
rect 5012 2309 5322 2343
rect 5012 2275 5114 2309
rect 5148 2275 5186 2309
rect 5220 2275 5322 2309
rect 5012 2241 5322 2275
rect 5012 2207 5114 2241
rect 5148 2207 5186 2241
rect 5220 2207 5322 2241
rect 5012 2173 5322 2207
rect 5012 2139 5114 2173
rect 5148 2139 5186 2173
rect 5220 2139 5322 2173
rect 5012 2105 5322 2139
rect 5012 2071 5114 2105
rect 5148 2071 5186 2105
rect 5220 2071 5322 2105
rect 5012 2037 5322 2071
rect 5012 2003 5114 2037
rect 5148 2003 5186 2037
rect 5220 2003 5322 2037
rect 5012 1969 5322 2003
rect 5012 1935 5114 1969
rect 5148 1935 5186 1969
rect 5220 1935 5322 1969
rect 5012 1901 5322 1935
rect 5012 1867 5114 1901
rect 5148 1867 5186 1901
rect 5220 1867 5322 1901
rect 5012 1833 5322 1867
rect 5012 1799 5114 1833
rect 5148 1799 5186 1833
rect 5220 1799 5322 1833
rect 5012 1765 5322 1799
rect 5012 1731 5114 1765
rect 5148 1731 5186 1765
rect 5220 1731 5322 1765
rect 5012 1697 5322 1731
rect 5012 1663 5114 1697
rect 5148 1663 5186 1697
rect 5220 1663 5322 1697
rect 5012 1629 5322 1663
rect 5012 1595 5114 1629
rect 5148 1595 5186 1629
rect 5220 1595 5322 1629
rect 5012 1561 5322 1595
rect 5012 1527 5114 1561
rect 5148 1527 5186 1561
rect 5220 1527 5322 1561
rect 5012 1457 5322 1527
rect 5442 2445 5593 2457
rect 5733 2445 5884 2457
rect 5442 2411 5544 2445
rect 5578 2411 5593 2445
rect 5733 2411 5748 2445
rect 5782 2411 5884 2445
rect 5442 2377 5593 2411
rect 5733 2377 5884 2411
rect 5442 2343 5544 2377
rect 5578 2343 5593 2377
rect 5733 2343 5748 2377
rect 5782 2343 5884 2377
rect 5442 2309 5593 2343
rect 5733 2309 5884 2343
rect 5442 2275 5544 2309
rect 5578 2275 5593 2309
rect 5733 2275 5748 2309
rect 5782 2275 5884 2309
rect 5442 2241 5593 2275
rect 5733 2241 5884 2275
rect 5442 2207 5544 2241
rect 5578 2207 5593 2241
rect 5733 2207 5748 2241
rect 5782 2207 5884 2241
rect 5442 2173 5593 2207
rect 5733 2173 5884 2207
rect 5442 2139 5544 2173
rect 5578 2139 5593 2173
rect 5733 2139 5748 2173
rect 5782 2139 5884 2173
rect 5442 2105 5593 2139
rect 5733 2105 5884 2139
rect 5442 2071 5544 2105
rect 5578 2071 5593 2105
rect 5733 2071 5748 2105
rect 5782 2071 5884 2105
rect 5442 2037 5593 2071
rect 5733 2037 5884 2071
rect 5442 2003 5544 2037
rect 5578 2003 5593 2037
rect 5733 2003 5748 2037
rect 5782 2003 5884 2037
rect 5442 1969 5593 2003
rect 5733 1969 5884 2003
rect 5442 1935 5544 1969
rect 5578 1935 5593 1969
rect 5733 1935 5748 1969
rect 5782 1935 5884 1969
rect 5442 1901 5593 1935
rect 5733 1901 5884 1935
rect 5442 1867 5544 1901
rect 5578 1867 5593 1901
rect 5733 1867 5748 1901
rect 5782 1867 5884 1901
rect 5442 1833 5593 1867
rect 5733 1833 5884 1867
rect 5442 1799 5544 1833
rect 5578 1799 5593 1833
rect 5733 1799 5748 1833
rect 5782 1799 5884 1833
rect 5442 1765 5593 1799
rect 5733 1765 5884 1799
rect 5442 1731 5544 1765
rect 5578 1731 5593 1765
rect 5733 1731 5748 1765
rect 5782 1731 5884 1765
rect 5442 1697 5593 1731
rect 5733 1697 5884 1731
rect 5442 1663 5544 1697
rect 5578 1663 5593 1697
rect 5733 1663 5748 1697
rect 5782 1663 5884 1697
rect 5442 1629 5593 1663
rect 5733 1629 5884 1663
rect 5442 1595 5544 1629
rect 5578 1595 5593 1629
rect 5733 1595 5748 1629
rect 5782 1595 5884 1629
rect 5442 1561 5593 1595
rect 5733 1561 5884 1595
rect 5442 1527 5544 1561
rect 5578 1527 5593 1561
rect 5733 1527 5748 1561
rect 5782 1527 5884 1561
rect 5442 1457 5593 1527
rect 5733 1457 5884 1527
rect 6004 2445 6314 2457
rect 6004 2411 6106 2445
rect 6140 2411 6178 2445
rect 6212 2411 6314 2445
rect 6004 2377 6314 2411
rect 6004 2343 6106 2377
rect 6140 2343 6178 2377
rect 6212 2343 6314 2377
rect 6004 2309 6314 2343
rect 6004 2275 6106 2309
rect 6140 2275 6178 2309
rect 6212 2275 6314 2309
rect 6004 2241 6314 2275
rect 6004 2207 6106 2241
rect 6140 2207 6178 2241
rect 6212 2207 6314 2241
rect 6004 2173 6314 2207
rect 6004 2139 6106 2173
rect 6140 2139 6178 2173
rect 6212 2139 6314 2173
rect 6004 2105 6314 2139
rect 6004 2071 6106 2105
rect 6140 2071 6178 2105
rect 6212 2071 6314 2105
rect 6004 2037 6314 2071
rect 6004 2003 6106 2037
rect 6140 2003 6178 2037
rect 6212 2003 6314 2037
rect 6004 1969 6314 2003
rect 6004 1935 6106 1969
rect 6140 1935 6178 1969
rect 6212 1935 6314 1969
rect 6004 1901 6314 1935
rect 6004 1867 6106 1901
rect 6140 1867 6178 1901
rect 6212 1867 6314 1901
rect 6004 1833 6314 1867
rect 6004 1799 6106 1833
rect 6140 1799 6178 1833
rect 6212 1799 6314 1833
rect 6004 1765 6314 1799
rect 6004 1731 6106 1765
rect 6140 1731 6178 1765
rect 6212 1731 6314 1765
rect 6004 1697 6314 1731
rect 6004 1663 6106 1697
rect 6140 1663 6178 1697
rect 6212 1663 6314 1697
rect 6004 1629 6314 1663
rect 6004 1595 6106 1629
rect 6140 1595 6178 1629
rect 6212 1595 6314 1629
rect 6004 1561 6314 1595
rect 6004 1527 6106 1561
rect 6140 1527 6178 1561
rect 6212 1527 6314 1561
rect 6004 1457 6314 1527
rect 6434 2445 6585 2457
rect 6725 2445 6876 2457
rect 6434 2411 6536 2445
rect 6570 2411 6585 2445
rect 6725 2411 6740 2445
rect 6774 2411 6876 2445
rect 6434 2377 6585 2411
rect 6725 2377 6876 2411
rect 6434 2343 6536 2377
rect 6570 2343 6585 2377
rect 6725 2343 6740 2377
rect 6774 2343 6876 2377
rect 6434 2309 6585 2343
rect 6725 2309 6876 2343
rect 6434 2275 6536 2309
rect 6570 2275 6585 2309
rect 6725 2275 6740 2309
rect 6774 2275 6876 2309
rect 6434 2241 6585 2275
rect 6725 2241 6876 2275
rect 6434 2207 6536 2241
rect 6570 2207 6585 2241
rect 6725 2207 6740 2241
rect 6774 2207 6876 2241
rect 6434 2173 6585 2207
rect 6725 2173 6876 2207
rect 6434 2139 6536 2173
rect 6570 2139 6585 2173
rect 6725 2139 6740 2173
rect 6774 2139 6876 2173
rect 6434 2105 6585 2139
rect 6725 2105 6876 2139
rect 6434 2071 6536 2105
rect 6570 2071 6585 2105
rect 6725 2071 6740 2105
rect 6774 2071 6876 2105
rect 6434 2037 6585 2071
rect 6725 2037 6876 2071
rect 6434 2003 6536 2037
rect 6570 2003 6585 2037
rect 6725 2003 6740 2037
rect 6774 2003 6876 2037
rect 6434 1969 6585 2003
rect 6725 1969 6876 2003
rect 6434 1935 6536 1969
rect 6570 1935 6585 1969
rect 6725 1935 6740 1969
rect 6774 1935 6876 1969
rect 6434 1901 6585 1935
rect 6725 1901 6876 1935
rect 6434 1867 6536 1901
rect 6570 1867 6585 1901
rect 6725 1867 6740 1901
rect 6774 1867 6876 1901
rect 6434 1833 6585 1867
rect 6725 1833 6876 1867
rect 6434 1799 6536 1833
rect 6570 1799 6585 1833
rect 6725 1799 6740 1833
rect 6774 1799 6876 1833
rect 6434 1765 6585 1799
rect 6725 1765 6876 1799
rect 6434 1731 6536 1765
rect 6570 1731 6585 1765
rect 6725 1731 6740 1765
rect 6774 1731 6876 1765
rect 6434 1697 6585 1731
rect 6725 1697 6876 1731
rect 6434 1663 6536 1697
rect 6570 1663 6585 1697
rect 6725 1663 6740 1697
rect 6774 1663 6876 1697
rect 6434 1629 6585 1663
rect 6725 1629 6876 1663
rect 6434 1595 6536 1629
rect 6570 1595 6585 1629
rect 6725 1595 6740 1629
rect 6774 1595 6876 1629
rect 6434 1561 6585 1595
rect 6725 1561 6876 1595
rect 6434 1527 6536 1561
rect 6570 1527 6585 1561
rect 6725 1527 6740 1561
rect 6774 1527 6876 1561
rect 6434 1457 6585 1527
rect 6725 1457 6876 1527
rect 6996 2445 7306 2457
rect 6996 2411 7098 2445
rect 7132 2411 7170 2445
rect 7204 2411 7306 2445
rect 6996 2377 7306 2411
rect 6996 2343 7098 2377
rect 7132 2343 7170 2377
rect 7204 2343 7306 2377
rect 6996 2309 7306 2343
rect 6996 2275 7098 2309
rect 7132 2275 7170 2309
rect 7204 2275 7306 2309
rect 6996 2241 7306 2275
rect 6996 2207 7098 2241
rect 7132 2207 7170 2241
rect 7204 2207 7306 2241
rect 6996 2173 7306 2207
rect 6996 2139 7098 2173
rect 7132 2139 7170 2173
rect 7204 2139 7306 2173
rect 6996 2105 7306 2139
rect 6996 2071 7098 2105
rect 7132 2071 7170 2105
rect 7204 2071 7306 2105
rect 6996 2037 7306 2071
rect 6996 2003 7098 2037
rect 7132 2003 7170 2037
rect 7204 2003 7306 2037
rect 6996 1969 7306 2003
rect 6996 1935 7098 1969
rect 7132 1935 7170 1969
rect 7204 1935 7306 1969
rect 6996 1901 7306 1935
rect 6996 1867 7098 1901
rect 7132 1867 7170 1901
rect 7204 1867 7306 1901
rect 6996 1833 7306 1867
rect 6996 1799 7098 1833
rect 7132 1799 7170 1833
rect 7204 1799 7306 1833
rect 6996 1765 7306 1799
rect 6996 1731 7098 1765
rect 7132 1731 7170 1765
rect 7204 1731 7306 1765
rect 6996 1697 7306 1731
rect 6996 1663 7098 1697
rect 7132 1663 7170 1697
rect 7204 1663 7306 1697
rect 6996 1629 7306 1663
rect 6996 1595 7098 1629
rect 7132 1595 7170 1629
rect 7204 1595 7306 1629
rect 6996 1561 7306 1595
rect 6996 1527 7098 1561
rect 7132 1527 7170 1561
rect 7204 1527 7306 1561
rect 6996 1457 7306 1527
rect 7426 2445 7577 2457
rect 7717 2445 7868 2457
rect 7426 2411 7528 2445
rect 7562 2411 7577 2445
rect 7717 2411 7732 2445
rect 7766 2411 7868 2445
rect 7426 2377 7577 2411
rect 7717 2377 7868 2411
rect 7426 2343 7528 2377
rect 7562 2343 7577 2377
rect 7717 2343 7732 2377
rect 7766 2343 7868 2377
rect 7426 2309 7577 2343
rect 7717 2309 7868 2343
rect 7426 2275 7528 2309
rect 7562 2275 7577 2309
rect 7717 2275 7732 2309
rect 7766 2275 7868 2309
rect 7426 2241 7577 2275
rect 7717 2241 7868 2275
rect 7426 2207 7528 2241
rect 7562 2207 7577 2241
rect 7717 2207 7732 2241
rect 7766 2207 7868 2241
rect 7426 2173 7577 2207
rect 7717 2173 7868 2207
rect 7426 2139 7528 2173
rect 7562 2139 7577 2173
rect 7717 2139 7732 2173
rect 7766 2139 7868 2173
rect 7426 2105 7577 2139
rect 7717 2105 7868 2139
rect 7426 2071 7528 2105
rect 7562 2071 7577 2105
rect 7717 2071 7732 2105
rect 7766 2071 7868 2105
rect 7426 2037 7577 2071
rect 7717 2037 7868 2071
rect 7426 2003 7528 2037
rect 7562 2003 7577 2037
rect 7717 2003 7732 2037
rect 7766 2003 7868 2037
rect 7426 1969 7577 2003
rect 7717 1969 7868 2003
rect 7426 1935 7528 1969
rect 7562 1935 7577 1969
rect 7717 1935 7732 1969
rect 7766 1935 7868 1969
rect 7426 1901 7577 1935
rect 7717 1901 7868 1935
rect 7426 1867 7528 1901
rect 7562 1867 7577 1901
rect 7717 1867 7732 1901
rect 7766 1867 7868 1901
rect 7426 1833 7577 1867
rect 7717 1833 7868 1867
rect 7426 1799 7528 1833
rect 7562 1799 7577 1833
rect 7717 1799 7732 1833
rect 7766 1799 7868 1833
rect 7426 1765 7577 1799
rect 7717 1765 7868 1799
rect 7426 1731 7528 1765
rect 7562 1731 7577 1765
rect 7717 1731 7732 1765
rect 7766 1731 7868 1765
rect 7426 1697 7577 1731
rect 7717 1697 7868 1731
rect 7426 1663 7528 1697
rect 7562 1663 7577 1697
rect 7717 1663 7732 1697
rect 7766 1663 7868 1697
rect 7426 1629 7577 1663
rect 7717 1629 7868 1663
rect 7426 1595 7528 1629
rect 7562 1595 7577 1629
rect 7717 1595 7732 1629
rect 7766 1595 7868 1629
rect 7426 1561 7577 1595
rect 7717 1561 7868 1595
rect 7426 1527 7528 1561
rect 7562 1527 7577 1561
rect 7717 1527 7732 1561
rect 7766 1527 7868 1561
rect 7426 1457 7577 1527
rect 7717 1457 7868 1527
rect 7988 2445 8298 2457
rect 7988 2411 8090 2445
rect 8124 2411 8162 2445
rect 8196 2411 8298 2445
rect 7988 2377 8298 2411
rect 7988 2343 8090 2377
rect 8124 2343 8162 2377
rect 8196 2343 8298 2377
rect 7988 2309 8298 2343
rect 7988 2275 8090 2309
rect 8124 2275 8162 2309
rect 8196 2275 8298 2309
rect 7988 2241 8298 2275
rect 7988 2207 8090 2241
rect 8124 2207 8162 2241
rect 8196 2207 8298 2241
rect 7988 2173 8298 2207
rect 7988 2139 8090 2173
rect 8124 2139 8162 2173
rect 8196 2139 8298 2173
rect 7988 2105 8298 2139
rect 7988 2071 8090 2105
rect 8124 2071 8162 2105
rect 8196 2071 8298 2105
rect 7988 2037 8298 2071
rect 7988 2003 8090 2037
rect 8124 2003 8162 2037
rect 8196 2003 8298 2037
rect 7988 1969 8298 2003
rect 7988 1935 8090 1969
rect 8124 1935 8162 1969
rect 8196 1935 8298 1969
rect 7988 1901 8298 1935
rect 7988 1867 8090 1901
rect 8124 1867 8162 1901
rect 8196 1867 8298 1901
rect 7988 1833 8298 1867
rect 7988 1799 8090 1833
rect 8124 1799 8162 1833
rect 8196 1799 8298 1833
rect 7988 1765 8298 1799
rect 7988 1731 8090 1765
rect 8124 1731 8162 1765
rect 8196 1731 8298 1765
rect 7988 1697 8298 1731
rect 7988 1663 8090 1697
rect 8124 1663 8162 1697
rect 8196 1663 8298 1697
rect 7988 1629 8298 1663
rect 7988 1595 8090 1629
rect 8124 1595 8162 1629
rect 8196 1595 8298 1629
rect 7988 1561 8298 1595
rect 7988 1527 8090 1561
rect 8124 1527 8162 1561
rect 8196 1527 8298 1561
rect 7988 1457 8298 1527
rect 8418 2445 8569 2457
rect 8709 2445 8860 2457
rect 8418 2411 8520 2445
rect 8554 2411 8569 2445
rect 8709 2411 8724 2445
rect 8758 2411 8860 2445
rect 8418 2377 8569 2411
rect 8709 2377 8860 2411
rect 8418 2343 8520 2377
rect 8554 2343 8569 2377
rect 8709 2343 8724 2377
rect 8758 2343 8860 2377
rect 8418 2309 8569 2343
rect 8709 2309 8860 2343
rect 8418 2275 8520 2309
rect 8554 2275 8569 2309
rect 8709 2275 8724 2309
rect 8758 2275 8860 2309
rect 8418 2241 8569 2275
rect 8709 2241 8860 2275
rect 8418 2207 8520 2241
rect 8554 2207 8569 2241
rect 8709 2207 8724 2241
rect 8758 2207 8860 2241
rect 8418 2173 8569 2207
rect 8709 2173 8860 2207
rect 8418 2139 8520 2173
rect 8554 2139 8569 2173
rect 8709 2139 8724 2173
rect 8758 2139 8860 2173
rect 8418 2105 8569 2139
rect 8709 2105 8860 2139
rect 8418 2071 8520 2105
rect 8554 2071 8569 2105
rect 8709 2071 8724 2105
rect 8758 2071 8860 2105
rect 8418 2037 8569 2071
rect 8709 2037 8860 2071
rect 8418 2003 8520 2037
rect 8554 2003 8569 2037
rect 8709 2003 8724 2037
rect 8758 2003 8860 2037
rect 8418 1969 8569 2003
rect 8709 1969 8860 2003
rect 8418 1935 8520 1969
rect 8554 1935 8569 1969
rect 8709 1935 8724 1969
rect 8758 1935 8860 1969
rect 8418 1901 8569 1935
rect 8709 1901 8860 1935
rect 8418 1867 8520 1901
rect 8554 1867 8569 1901
rect 8709 1867 8724 1901
rect 8758 1867 8860 1901
rect 8418 1833 8569 1867
rect 8709 1833 8860 1867
rect 8418 1799 8520 1833
rect 8554 1799 8569 1833
rect 8709 1799 8724 1833
rect 8758 1799 8860 1833
rect 8418 1765 8569 1799
rect 8709 1765 8860 1799
rect 8418 1731 8520 1765
rect 8554 1731 8569 1765
rect 8709 1731 8724 1765
rect 8758 1731 8860 1765
rect 8418 1697 8569 1731
rect 8709 1697 8860 1731
rect 8418 1663 8520 1697
rect 8554 1663 8569 1697
rect 8709 1663 8724 1697
rect 8758 1663 8860 1697
rect 8418 1629 8569 1663
rect 8709 1629 8860 1663
rect 8418 1595 8520 1629
rect 8554 1595 8569 1629
rect 8709 1595 8724 1629
rect 8758 1595 8860 1629
rect 8418 1561 8569 1595
rect 8709 1561 8860 1595
rect 8418 1527 8520 1561
rect 8554 1527 8569 1561
rect 8709 1527 8724 1561
rect 8758 1527 8860 1561
rect 8418 1457 8569 1527
rect 8709 1457 8860 1527
rect 8980 2445 9290 2457
rect 8980 2411 9082 2445
rect 9116 2411 9154 2445
rect 9188 2411 9290 2445
rect 8980 2377 9290 2411
rect 8980 2343 9082 2377
rect 9116 2343 9154 2377
rect 9188 2343 9290 2377
rect 8980 2309 9290 2343
rect 8980 2275 9082 2309
rect 9116 2275 9154 2309
rect 9188 2275 9290 2309
rect 8980 2241 9290 2275
rect 8980 2207 9082 2241
rect 9116 2207 9154 2241
rect 9188 2207 9290 2241
rect 8980 2173 9290 2207
rect 8980 2139 9082 2173
rect 9116 2139 9154 2173
rect 9188 2139 9290 2173
rect 8980 2105 9290 2139
rect 8980 2071 9082 2105
rect 9116 2071 9154 2105
rect 9188 2071 9290 2105
rect 8980 2037 9290 2071
rect 8980 2003 9082 2037
rect 9116 2003 9154 2037
rect 9188 2003 9290 2037
rect 8980 1969 9290 2003
rect 8980 1935 9082 1969
rect 9116 1935 9154 1969
rect 9188 1935 9290 1969
rect 8980 1901 9290 1935
rect 8980 1867 9082 1901
rect 9116 1867 9154 1901
rect 9188 1867 9290 1901
rect 8980 1833 9290 1867
rect 8980 1799 9082 1833
rect 9116 1799 9154 1833
rect 9188 1799 9290 1833
rect 8980 1765 9290 1799
rect 8980 1731 9082 1765
rect 9116 1731 9154 1765
rect 9188 1731 9290 1765
rect 8980 1697 9290 1731
rect 8980 1663 9082 1697
rect 9116 1663 9154 1697
rect 9188 1663 9290 1697
rect 8980 1629 9290 1663
rect 8980 1595 9082 1629
rect 9116 1595 9154 1629
rect 9188 1595 9290 1629
rect 8980 1561 9290 1595
rect 8980 1527 9082 1561
rect 9116 1527 9154 1561
rect 9188 1527 9290 1561
rect 8980 1457 9290 1527
rect 9410 2445 9561 2457
rect 9701 2445 9852 2457
rect 9410 2411 9512 2445
rect 9546 2411 9561 2445
rect 9701 2411 9716 2445
rect 9750 2411 9852 2445
rect 9410 2377 9561 2411
rect 9701 2377 9852 2411
rect 9410 2343 9512 2377
rect 9546 2343 9561 2377
rect 9701 2343 9716 2377
rect 9750 2343 9852 2377
rect 9410 2309 9561 2343
rect 9701 2309 9852 2343
rect 9410 2275 9512 2309
rect 9546 2275 9561 2309
rect 9701 2275 9716 2309
rect 9750 2275 9852 2309
rect 9410 2241 9561 2275
rect 9701 2241 9852 2275
rect 9410 2207 9512 2241
rect 9546 2207 9561 2241
rect 9701 2207 9716 2241
rect 9750 2207 9852 2241
rect 9410 2173 9561 2207
rect 9701 2173 9852 2207
rect 9410 2139 9512 2173
rect 9546 2139 9561 2173
rect 9701 2139 9716 2173
rect 9750 2139 9852 2173
rect 9410 2105 9561 2139
rect 9701 2105 9852 2139
rect 9410 2071 9512 2105
rect 9546 2071 9561 2105
rect 9701 2071 9716 2105
rect 9750 2071 9852 2105
rect 9410 2037 9561 2071
rect 9701 2037 9852 2071
rect 9410 2003 9512 2037
rect 9546 2003 9561 2037
rect 9701 2003 9716 2037
rect 9750 2003 9852 2037
rect 9410 1969 9561 2003
rect 9701 1969 9852 2003
rect 9410 1935 9512 1969
rect 9546 1935 9561 1969
rect 9701 1935 9716 1969
rect 9750 1935 9852 1969
rect 9410 1901 9561 1935
rect 9701 1901 9852 1935
rect 9410 1867 9512 1901
rect 9546 1867 9561 1901
rect 9701 1867 9716 1901
rect 9750 1867 9852 1901
rect 9410 1833 9561 1867
rect 9701 1833 9852 1867
rect 9410 1799 9512 1833
rect 9546 1799 9561 1833
rect 9701 1799 9716 1833
rect 9750 1799 9852 1833
rect 9410 1765 9561 1799
rect 9701 1765 9852 1799
rect 9410 1731 9512 1765
rect 9546 1731 9561 1765
rect 9701 1731 9716 1765
rect 9750 1731 9852 1765
rect 9410 1697 9561 1731
rect 9701 1697 9852 1731
rect 9410 1663 9512 1697
rect 9546 1663 9561 1697
rect 9701 1663 9716 1697
rect 9750 1663 9852 1697
rect 9410 1629 9561 1663
rect 9701 1629 9852 1663
rect 9410 1595 9512 1629
rect 9546 1595 9561 1629
rect 9701 1595 9716 1629
rect 9750 1595 9852 1629
rect 9410 1561 9561 1595
rect 9701 1561 9852 1595
rect 9410 1527 9512 1561
rect 9546 1527 9561 1561
rect 9701 1527 9716 1561
rect 9750 1527 9852 1561
rect 9410 1457 9561 1527
rect 9701 1457 9852 1527
rect 9972 2445 10282 2457
rect 9972 2411 10074 2445
rect 10108 2411 10146 2445
rect 10180 2411 10282 2445
rect 9972 2377 10282 2411
rect 9972 2343 10074 2377
rect 10108 2343 10146 2377
rect 10180 2343 10282 2377
rect 9972 2309 10282 2343
rect 9972 2275 10074 2309
rect 10108 2275 10146 2309
rect 10180 2275 10282 2309
rect 9972 2241 10282 2275
rect 9972 2207 10074 2241
rect 10108 2207 10146 2241
rect 10180 2207 10282 2241
rect 9972 2173 10282 2207
rect 9972 2139 10074 2173
rect 10108 2139 10146 2173
rect 10180 2139 10282 2173
rect 9972 2105 10282 2139
rect 9972 2071 10074 2105
rect 10108 2071 10146 2105
rect 10180 2071 10282 2105
rect 9972 2037 10282 2071
rect 9972 2003 10074 2037
rect 10108 2003 10146 2037
rect 10180 2003 10282 2037
rect 9972 1969 10282 2003
rect 9972 1935 10074 1969
rect 10108 1935 10146 1969
rect 10180 1935 10282 1969
rect 9972 1901 10282 1935
rect 9972 1867 10074 1901
rect 10108 1867 10146 1901
rect 10180 1867 10282 1901
rect 9972 1833 10282 1867
rect 9972 1799 10074 1833
rect 10108 1799 10146 1833
rect 10180 1799 10282 1833
rect 9972 1765 10282 1799
rect 9972 1731 10074 1765
rect 10108 1731 10146 1765
rect 10180 1731 10282 1765
rect 9972 1697 10282 1731
rect 9972 1663 10074 1697
rect 10108 1663 10146 1697
rect 10180 1663 10282 1697
rect 9972 1629 10282 1663
rect 9972 1595 10074 1629
rect 10108 1595 10146 1629
rect 10180 1595 10282 1629
rect 9972 1561 10282 1595
rect 9972 1527 10074 1561
rect 10108 1527 10146 1561
rect 10180 1527 10282 1561
rect 9972 1457 10282 1527
rect 10402 2445 10553 2457
rect 10693 2445 10844 2457
rect 10402 2411 10504 2445
rect 10538 2411 10553 2445
rect 10693 2411 10708 2445
rect 10742 2411 10844 2445
rect 10402 2377 10553 2411
rect 10693 2377 10844 2411
rect 10402 2343 10504 2377
rect 10538 2343 10553 2377
rect 10693 2343 10708 2377
rect 10742 2343 10844 2377
rect 10402 2309 10553 2343
rect 10693 2309 10844 2343
rect 10402 2275 10504 2309
rect 10538 2275 10553 2309
rect 10693 2275 10708 2309
rect 10742 2275 10844 2309
rect 10402 2241 10553 2275
rect 10693 2241 10844 2275
rect 10402 2207 10504 2241
rect 10538 2207 10553 2241
rect 10693 2207 10708 2241
rect 10742 2207 10844 2241
rect 10402 2173 10553 2207
rect 10693 2173 10844 2207
rect 10402 2139 10504 2173
rect 10538 2139 10553 2173
rect 10693 2139 10708 2173
rect 10742 2139 10844 2173
rect 10402 2105 10553 2139
rect 10693 2105 10844 2139
rect 10402 2071 10504 2105
rect 10538 2071 10553 2105
rect 10693 2071 10708 2105
rect 10742 2071 10844 2105
rect 10402 2037 10553 2071
rect 10693 2037 10844 2071
rect 10402 2003 10504 2037
rect 10538 2003 10553 2037
rect 10693 2003 10708 2037
rect 10742 2003 10844 2037
rect 10402 1969 10553 2003
rect 10693 1969 10844 2003
rect 10402 1935 10504 1969
rect 10538 1935 10553 1969
rect 10693 1935 10708 1969
rect 10742 1935 10844 1969
rect 10402 1901 10553 1935
rect 10693 1901 10844 1935
rect 10402 1867 10504 1901
rect 10538 1867 10553 1901
rect 10693 1867 10708 1901
rect 10742 1867 10844 1901
rect 10402 1833 10553 1867
rect 10693 1833 10844 1867
rect 10402 1799 10504 1833
rect 10538 1799 10553 1833
rect 10693 1799 10708 1833
rect 10742 1799 10844 1833
rect 10402 1765 10553 1799
rect 10693 1765 10844 1799
rect 10402 1731 10504 1765
rect 10538 1731 10553 1765
rect 10693 1731 10708 1765
rect 10742 1731 10844 1765
rect 10402 1697 10553 1731
rect 10693 1697 10844 1731
rect 10402 1663 10504 1697
rect 10538 1663 10553 1697
rect 10693 1663 10708 1697
rect 10742 1663 10844 1697
rect 10402 1629 10553 1663
rect 10693 1629 10844 1663
rect 10402 1595 10504 1629
rect 10538 1595 10553 1629
rect 10693 1595 10708 1629
rect 10742 1595 10844 1629
rect 10402 1561 10553 1595
rect 10693 1561 10844 1595
rect 10402 1527 10504 1561
rect 10538 1527 10553 1561
rect 10693 1527 10708 1561
rect 10742 1527 10844 1561
rect 10402 1457 10553 1527
rect 10693 1457 10844 1527
rect 10964 2445 11274 2457
rect 10964 2411 11066 2445
rect 11100 2411 11138 2445
rect 11172 2411 11274 2445
rect 10964 2377 11274 2411
rect 10964 2343 11066 2377
rect 11100 2343 11138 2377
rect 11172 2343 11274 2377
rect 10964 2309 11274 2343
rect 10964 2275 11066 2309
rect 11100 2275 11138 2309
rect 11172 2275 11274 2309
rect 10964 2241 11274 2275
rect 10964 2207 11066 2241
rect 11100 2207 11138 2241
rect 11172 2207 11274 2241
rect 10964 2173 11274 2207
rect 10964 2139 11066 2173
rect 11100 2139 11138 2173
rect 11172 2139 11274 2173
rect 10964 2105 11274 2139
rect 10964 2071 11066 2105
rect 11100 2071 11138 2105
rect 11172 2071 11274 2105
rect 10964 2037 11274 2071
rect 10964 2003 11066 2037
rect 11100 2003 11138 2037
rect 11172 2003 11274 2037
rect 10964 1969 11274 2003
rect 10964 1935 11066 1969
rect 11100 1935 11138 1969
rect 11172 1935 11274 1969
rect 10964 1901 11274 1935
rect 10964 1867 11066 1901
rect 11100 1867 11138 1901
rect 11172 1867 11274 1901
rect 10964 1833 11274 1867
rect 10964 1799 11066 1833
rect 11100 1799 11138 1833
rect 11172 1799 11274 1833
rect 10964 1765 11274 1799
rect 10964 1731 11066 1765
rect 11100 1731 11138 1765
rect 11172 1731 11274 1765
rect 10964 1697 11274 1731
rect 10964 1663 11066 1697
rect 11100 1663 11138 1697
rect 11172 1663 11274 1697
rect 10964 1629 11274 1663
rect 10964 1595 11066 1629
rect 11100 1595 11138 1629
rect 11172 1595 11274 1629
rect 10964 1561 11274 1595
rect 10964 1527 11066 1561
rect 11100 1527 11138 1561
rect 11172 1527 11274 1561
rect 10964 1457 11274 1527
rect 11394 2445 11545 2457
rect 11685 2445 11836 2457
rect 11394 2411 11496 2445
rect 11530 2411 11545 2445
rect 11685 2411 11700 2445
rect 11734 2411 11836 2445
rect 11394 2377 11545 2411
rect 11685 2377 11836 2411
rect 11394 2343 11496 2377
rect 11530 2343 11545 2377
rect 11685 2343 11700 2377
rect 11734 2343 11836 2377
rect 11394 2309 11545 2343
rect 11685 2309 11836 2343
rect 11394 2275 11496 2309
rect 11530 2275 11545 2309
rect 11685 2275 11700 2309
rect 11734 2275 11836 2309
rect 11394 2241 11545 2275
rect 11685 2241 11836 2275
rect 11394 2207 11496 2241
rect 11530 2207 11545 2241
rect 11685 2207 11700 2241
rect 11734 2207 11836 2241
rect 11394 2173 11545 2207
rect 11685 2173 11836 2207
rect 11394 2139 11496 2173
rect 11530 2139 11545 2173
rect 11685 2139 11700 2173
rect 11734 2139 11836 2173
rect 11394 2105 11545 2139
rect 11685 2105 11836 2139
rect 11394 2071 11496 2105
rect 11530 2071 11545 2105
rect 11685 2071 11700 2105
rect 11734 2071 11836 2105
rect 11394 2037 11545 2071
rect 11685 2037 11836 2071
rect 11394 2003 11496 2037
rect 11530 2003 11545 2037
rect 11685 2003 11700 2037
rect 11734 2003 11836 2037
rect 11394 1969 11545 2003
rect 11685 1969 11836 2003
rect 11394 1935 11496 1969
rect 11530 1935 11545 1969
rect 11685 1935 11700 1969
rect 11734 1935 11836 1969
rect 11394 1901 11545 1935
rect 11685 1901 11836 1935
rect 11394 1867 11496 1901
rect 11530 1867 11545 1901
rect 11685 1867 11700 1901
rect 11734 1867 11836 1901
rect 11394 1833 11545 1867
rect 11685 1833 11836 1867
rect 11394 1799 11496 1833
rect 11530 1799 11545 1833
rect 11685 1799 11700 1833
rect 11734 1799 11836 1833
rect 11394 1765 11545 1799
rect 11685 1765 11836 1799
rect 11394 1731 11496 1765
rect 11530 1731 11545 1765
rect 11685 1731 11700 1765
rect 11734 1731 11836 1765
rect 11394 1697 11545 1731
rect 11685 1697 11836 1731
rect 11394 1663 11496 1697
rect 11530 1663 11545 1697
rect 11685 1663 11700 1697
rect 11734 1663 11836 1697
rect 11394 1629 11545 1663
rect 11685 1629 11836 1663
rect 11394 1595 11496 1629
rect 11530 1595 11545 1629
rect 11685 1595 11700 1629
rect 11734 1595 11836 1629
rect 11394 1561 11545 1595
rect 11685 1561 11836 1595
rect 11394 1527 11496 1561
rect 11530 1527 11545 1561
rect 11685 1527 11700 1561
rect 11734 1527 11836 1561
rect 11394 1457 11545 1527
rect 11685 1457 11836 1527
rect 11956 2445 12266 2457
rect 11956 2411 12058 2445
rect 12092 2411 12130 2445
rect 12164 2411 12266 2445
rect 11956 2377 12266 2411
rect 11956 2343 12058 2377
rect 12092 2343 12130 2377
rect 12164 2343 12266 2377
rect 11956 2309 12266 2343
rect 11956 2275 12058 2309
rect 12092 2275 12130 2309
rect 12164 2275 12266 2309
rect 11956 2241 12266 2275
rect 11956 2207 12058 2241
rect 12092 2207 12130 2241
rect 12164 2207 12266 2241
rect 11956 2173 12266 2207
rect 11956 2139 12058 2173
rect 12092 2139 12130 2173
rect 12164 2139 12266 2173
rect 11956 2105 12266 2139
rect 11956 2071 12058 2105
rect 12092 2071 12130 2105
rect 12164 2071 12266 2105
rect 11956 2037 12266 2071
rect 11956 2003 12058 2037
rect 12092 2003 12130 2037
rect 12164 2003 12266 2037
rect 11956 1969 12266 2003
rect 11956 1935 12058 1969
rect 12092 1935 12130 1969
rect 12164 1935 12266 1969
rect 11956 1901 12266 1935
rect 11956 1867 12058 1901
rect 12092 1867 12130 1901
rect 12164 1867 12266 1901
rect 11956 1833 12266 1867
rect 11956 1799 12058 1833
rect 12092 1799 12130 1833
rect 12164 1799 12266 1833
rect 11956 1765 12266 1799
rect 11956 1731 12058 1765
rect 12092 1731 12130 1765
rect 12164 1731 12266 1765
rect 11956 1697 12266 1731
rect 11956 1663 12058 1697
rect 12092 1663 12130 1697
rect 12164 1663 12266 1697
rect 11956 1629 12266 1663
rect 11956 1595 12058 1629
rect 12092 1595 12130 1629
rect 12164 1595 12266 1629
rect 11956 1561 12266 1595
rect 11956 1527 12058 1561
rect 12092 1527 12130 1561
rect 12164 1527 12266 1561
rect 11956 1457 12266 1527
rect 12386 2445 12537 2457
rect 12677 2445 12828 2457
rect 12386 2411 12488 2445
rect 12522 2411 12537 2445
rect 12677 2411 12692 2445
rect 12726 2411 12828 2445
rect 12386 2377 12537 2411
rect 12677 2377 12828 2411
rect 12386 2343 12488 2377
rect 12522 2343 12537 2377
rect 12677 2343 12692 2377
rect 12726 2343 12828 2377
rect 12386 2309 12537 2343
rect 12677 2309 12828 2343
rect 12386 2275 12488 2309
rect 12522 2275 12537 2309
rect 12677 2275 12692 2309
rect 12726 2275 12828 2309
rect 12386 2241 12537 2275
rect 12677 2241 12828 2275
rect 12386 2207 12488 2241
rect 12522 2207 12537 2241
rect 12677 2207 12692 2241
rect 12726 2207 12828 2241
rect 12386 2173 12537 2207
rect 12677 2173 12828 2207
rect 12386 2139 12488 2173
rect 12522 2139 12537 2173
rect 12677 2139 12692 2173
rect 12726 2139 12828 2173
rect 12386 2105 12537 2139
rect 12677 2105 12828 2139
rect 12386 2071 12488 2105
rect 12522 2071 12537 2105
rect 12677 2071 12692 2105
rect 12726 2071 12828 2105
rect 12386 2037 12537 2071
rect 12677 2037 12828 2071
rect 12386 2003 12488 2037
rect 12522 2003 12537 2037
rect 12677 2003 12692 2037
rect 12726 2003 12828 2037
rect 12386 1969 12537 2003
rect 12677 1969 12828 2003
rect 12386 1935 12488 1969
rect 12522 1935 12537 1969
rect 12677 1935 12692 1969
rect 12726 1935 12828 1969
rect 12386 1901 12537 1935
rect 12677 1901 12828 1935
rect 12386 1867 12488 1901
rect 12522 1867 12537 1901
rect 12677 1867 12692 1901
rect 12726 1867 12828 1901
rect 12386 1833 12537 1867
rect 12677 1833 12828 1867
rect 12386 1799 12488 1833
rect 12522 1799 12537 1833
rect 12677 1799 12692 1833
rect 12726 1799 12828 1833
rect 12386 1765 12537 1799
rect 12677 1765 12828 1799
rect 12386 1731 12488 1765
rect 12522 1731 12537 1765
rect 12677 1731 12692 1765
rect 12726 1731 12828 1765
rect 12386 1697 12537 1731
rect 12677 1697 12828 1731
rect 12386 1663 12488 1697
rect 12522 1663 12537 1697
rect 12677 1663 12692 1697
rect 12726 1663 12828 1697
rect 12386 1629 12537 1663
rect 12677 1629 12828 1663
rect 12386 1595 12488 1629
rect 12522 1595 12537 1629
rect 12677 1595 12692 1629
rect 12726 1595 12828 1629
rect 12386 1561 12537 1595
rect 12677 1561 12828 1595
rect 12386 1527 12488 1561
rect 12522 1527 12537 1561
rect 12677 1527 12692 1561
rect 12726 1527 12828 1561
rect 12386 1457 12537 1527
rect 12677 1457 12828 1527
rect 12948 2445 13258 2457
rect 12948 2411 13050 2445
rect 13084 2411 13122 2445
rect 13156 2411 13258 2445
rect 12948 2377 13258 2411
rect 12948 2343 13050 2377
rect 13084 2343 13122 2377
rect 13156 2343 13258 2377
rect 12948 2309 13258 2343
rect 12948 2275 13050 2309
rect 13084 2275 13122 2309
rect 13156 2275 13258 2309
rect 12948 2241 13258 2275
rect 12948 2207 13050 2241
rect 13084 2207 13122 2241
rect 13156 2207 13258 2241
rect 12948 2173 13258 2207
rect 12948 2139 13050 2173
rect 13084 2139 13122 2173
rect 13156 2139 13258 2173
rect 12948 2105 13258 2139
rect 12948 2071 13050 2105
rect 13084 2071 13122 2105
rect 13156 2071 13258 2105
rect 12948 2037 13258 2071
rect 12948 2003 13050 2037
rect 13084 2003 13122 2037
rect 13156 2003 13258 2037
rect 12948 1969 13258 2003
rect 12948 1935 13050 1969
rect 13084 1935 13122 1969
rect 13156 1935 13258 1969
rect 12948 1901 13258 1935
rect 12948 1867 13050 1901
rect 13084 1867 13122 1901
rect 13156 1867 13258 1901
rect 12948 1833 13258 1867
rect 12948 1799 13050 1833
rect 13084 1799 13122 1833
rect 13156 1799 13258 1833
rect 12948 1765 13258 1799
rect 12948 1731 13050 1765
rect 13084 1731 13122 1765
rect 13156 1731 13258 1765
rect 12948 1697 13258 1731
rect 12948 1663 13050 1697
rect 13084 1663 13122 1697
rect 13156 1663 13258 1697
rect 12948 1629 13258 1663
rect 12948 1595 13050 1629
rect 13084 1595 13122 1629
rect 13156 1595 13258 1629
rect 12948 1561 13258 1595
rect 12948 1527 13050 1561
rect 13084 1527 13122 1561
rect 13156 1527 13258 1561
rect 12948 1457 13258 1527
rect 13378 2445 13529 2457
rect 13669 2445 13820 2457
rect 13378 2411 13480 2445
rect 13514 2411 13529 2445
rect 13669 2411 13684 2445
rect 13718 2411 13820 2445
rect 13378 2377 13529 2411
rect 13669 2377 13820 2411
rect 13378 2343 13480 2377
rect 13514 2343 13529 2377
rect 13669 2343 13684 2377
rect 13718 2343 13820 2377
rect 13378 2309 13529 2343
rect 13669 2309 13820 2343
rect 13378 2275 13480 2309
rect 13514 2275 13529 2309
rect 13669 2275 13684 2309
rect 13718 2275 13820 2309
rect 13378 2241 13529 2275
rect 13669 2241 13820 2275
rect 13378 2207 13480 2241
rect 13514 2207 13529 2241
rect 13669 2207 13684 2241
rect 13718 2207 13820 2241
rect 13378 2173 13529 2207
rect 13669 2173 13820 2207
rect 13378 2139 13480 2173
rect 13514 2139 13529 2173
rect 13669 2139 13684 2173
rect 13718 2139 13820 2173
rect 13378 2105 13529 2139
rect 13669 2105 13820 2139
rect 13378 2071 13480 2105
rect 13514 2071 13529 2105
rect 13669 2071 13684 2105
rect 13718 2071 13820 2105
rect 13378 2037 13529 2071
rect 13669 2037 13820 2071
rect 13378 2003 13480 2037
rect 13514 2003 13529 2037
rect 13669 2003 13684 2037
rect 13718 2003 13820 2037
rect 13378 1969 13529 2003
rect 13669 1969 13820 2003
rect 13378 1935 13480 1969
rect 13514 1935 13529 1969
rect 13669 1935 13684 1969
rect 13718 1935 13820 1969
rect 13378 1901 13529 1935
rect 13669 1901 13820 1935
rect 13378 1867 13480 1901
rect 13514 1867 13529 1901
rect 13669 1867 13684 1901
rect 13718 1867 13820 1901
rect 13378 1833 13529 1867
rect 13669 1833 13820 1867
rect 13378 1799 13480 1833
rect 13514 1799 13529 1833
rect 13669 1799 13684 1833
rect 13718 1799 13820 1833
rect 13378 1765 13529 1799
rect 13669 1765 13820 1799
rect 13378 1731 13480 1765
rect 13514 1731 13529 1765
rect 13669 1731 13684 1765
rect 13718 1731 13820 1765
rect 13378 1697 13529 1731
rect 13669 1697 13820 1731
rect 13378 1663 13480 1697
rect 13514 1663 13529 1697
rect 13669 1663 13684 1697
rect 13718 1663 13820 1697
rect 13378 1629 13529 1663
rect 13669 1629 13820 1663
rect 13378 1595 13480 1629
rect 13514 1595 13529 1629
rect 13669 1595 13684 1629
rect 13718 1595 13820 1629
rect 13378 1561 13529 1595
rect 13669 1561 13820 1595
rect 13378 1527 13480 1561
rect 13514 1527 13529 1561
rect 13669 1527 13684 1561
rect 13718 1527 13820 1561
rect 13378 1457 13529 1527
rect 13669 1457 13820 1527
rect 13940 2445 14178 2457
rect 13940 2411 14042 2445
rect 14076 2411 14178 2445
rect 13940 2377 14178 2411
rect 13940 2343 14042 2377
rect 14076 2343 14178 2377
rect 13940 2309 14178 2343
rect 13940 2275 14042 2309
rect 14076 2275 14178 2309
rect 13940 2241 14178 2275
rect 13940 2207 14042 2241
rect 14076 2207 14178 2241
rect 13940 2173 14178 2207
rect 13940 2139 14042 2173
rect 14076 2139 14178 2173
rect 13940 2105 14178 2139
rect 13940 2071 14042 2105
rect 14076 2071 14178 2105
rect 13940 2037 14178 2071
rect 13940 2003 14042 2037
rect 14076 2003 14178 2037
rect 13940 1969 14178 2003
rect 13940 1935 14042 1969
rect 14076 1935 14178 1969
rect 13940 1901 14178 1935
rect 13940 1867 14042 1901
rect 14076 1867 14178 1901
rect 13940 1833 14178 1867
rect 13940 1799 14042 1833
rect 14076 1799 14178 1833
rect 13940 1765 14178 1799
rect 13940 1731 14042 1765
rect 14076 1731 14178 1765
rect 13940 1697 14178 1731
rect 13940 1663 14042 1697
rect 14076 1663 14178 1697
rect 13940 1629 14178 1663
rect 13940 1595 14042 1629
rect 14076 1595 14178 1629
rect 13940 1561 14178 1595
rect 13940 1527 14042 1561
rect 14076 1527 14178 1561
rect 13940 1457 14178 1527
rect 14298 2445 14435 2457
rect 14298 2411 14386 2445
rect 14420 2411 14435 2445
rect 14298 2377 14435 2411
rect 14298 2343 14386 2377
rect 14420 2343 14435 2377
rect 14298 2309 14435 2343
rect 14298 2275 14386 2309
rect 14420 2275 14435 2309
rect 14298 2241 14435 2275
rect 14298 2207 14386 2241
rect 14420 2207 14435 2241
rect 14298 2173 14435 2207
rect 14298 2139 14386 2173
rect 14420 2139 14435 2173
rect 14298 2105 14435 2139
rect 14298 2071 14386 2105
rect 14420 2071 14435 2105
rect 14298 2037 14435 2071
rect 14298 2003 14386 2037
rect 14420 2003 14435 2037
rect 14298 1969 14435 2003
rect 14298 1935 14386 1969
rect 14420 1935 14435 1969
rect 14298 1901 14435 1935
rect 14298 1867 14386 1901
rect 14420 1867 14435 1901
rect 14298 1833 14435 1867
rect 14298 1799 14386 1833
rect 14420 1799 14435 1833
rect 14298 1765 14435 1799
rect 14298 1731 14386 1765
rect 14420 1731 14435 1765
rect 14298 1697 14435 1731
rect 14298 1663 14386 1697
rect 14420 1663 14435 1697
rect 14298 1629 14435 1663
rect 14298 1595 14386 1629
rect 14420 1595 14435 1629
rect 14298 1561 14435 1595
rect 14298 1527 14386 1561
rect 14420 1527 14435 1561
rect 14298 1457 14435 1527
<< mvndiffc >>
rect 802 4012 836 4046
rect 802 3944 836 3978
rect 802 3876 836 3910
rect 802 3808 836 3842
rect 802 3740 836 3774
rect 802 3672 836 3706
rect 802 3604 836 3638
rect 802 3536 836 3570
rect 802 3468 836 3502
rect 802 3400 836 3434
rect 802 3332 836 3366
rect 802 3264 836 3298
rect 802 3196 836 3230
rect 802 3128 836 3162
rect 1146 4012 1180 4046
rect 1218 4012 1252 4046
rect 1146 3944 1180 3978
rect 1218 3944 1252 3978
rect 1146 3876 1180 3910
rect 1218 3876 1252 3910
rect 1146 3808 1180 3842
rect 1218 3808 1252 3842
rect 1146 3740 1180 3774
rect 1218 3740 1252 3774
rect 1146 3672 1180 3706
rect 1218 3672 1252 3706
rect 1146 3604 1180 3638
rect 1218 3604 1252 3638
rect 1146 3536 1180 3570
rect 1218 3536 1252 3570
rect 1146 3468 1180 3502
rect 1218 3468 1252 3502
rect 1146 3400 1180 3434
rect 1218 3400 1252 3434
rect 1146 3332 1180 3366
rect 1218 3332 1252 3366
rect 1146 3264 1180 3298
rect 1218 3264 1252 3298
rect 1146 3196 1180 3230
rect 1218 3196 1252 3230
rect 1146 3128 1180 3162
rect 1218 3128 1252 3162
rect 1576 4012 1610 4046
rect 1780 4012 1814 4046
rect 1576 3944 1610 3978
rect 1780 3944 1814 3978
rect 1576 3876 1610 3910
rect 1780 3876 1814 3910
rect 1576 3808 1610 3842
rect 1780 3808 1814 3842
rect 1576 3740 1610 3774
rect 1780 3740 1814 3774
rect 1576 3672 1610 3706
rect 1780 3672 1814 3706
rect 1576 3604 1610 3638
rect 1780 3604 1814 3638
rect 1576 3536 1610 3570
rect 1780 3536 1814 3570
rect 1576 3468 1610 3502
rect 1780 3468 1814 3502
rect 1576 3400 1610 3434
rect 1780 3400 1814 3434
rect 1576 3332 1610 3366
rect 1780 3332 1814 3366
rect 1576 3264 1610 3298
rect 1780 3264 1814 3298
rect 1576 3196 1610 3230
rect 1780 3196 1814 3230
rect 1576 3128 1610 3162
rect 1780 3128 1814 3162
rect 2138 4012 2172 4046
rect 2210 4012 2244 4046
rect 2138 3944 2172 3978
rect 2210 3944 2244 3978
rect 2138 3876 2172 3910
rect 2210 3876 2244 3910
rect 2138 3808 2172 3842
rect 2210 3808 2244 3842
rect 2138 3740 2172 3774
rect 2210 3740 2244 3774
rect 2138 3672 2172 3706
rect 2210 3672 2244 3706
rect 2138 3604 2172 3638
rect 2210 3604 2244 3638
rect 2138 3536 2172 3570
rect 2210 3536 2244 3570
rect 2138 3468 2172 3502
rect 2210 3468 2244 3502
rect 2138 3400 2172 3434
rect 2210 3400 2244 3434
rect 2138 3332 2172 3366
rect 2210 3332 2244 3366
rect 2138 3264 2172 3298
rect 2210 3264 2244 3298
rect 2138 3196 2172 3230
rect 2210 3196 2244 3230
rect 2138 3128 2172 3162
rect 2210 3128 2244 3162
rect 2568 4012 2602 4046
rect 2772 4012 2806 4046
rect 2568 3944 2602 3978
rect 2772 3944 2806 3978
rect 2568 3876 2602 3910
rect 2772 3876 2806 3910
rect 2568 3808 2602 3842
rect 2772 3808 2806 3842
rect 2568 3740 2602 3774
rect 2772 3740 2806 3774
rect 2568 3672 2602 3706
rect 2772 3672 2806 3706
rect 2568 3604 2602 3638
rect 2772 3604 2806 3638
rect 2568 3536 2602 3570
rect 2772 3536 2806 3570
rect 2568 3468 2602 3502
rect 2772 3468 2806 3502
rect 2568 3400 2602 3434
rect 2772 3400 2806 3434
rect 2568 3332 2602 3366
rect 2772 3332 2806 3366
rect 2568 3264 2602 3298
rect 2772 3264 2806 3298
rect 2568 3196 2602 3230
rect 2772 3196 2806 3230
rect 2568 3128 2602 3162
rect 2772 3128 2806 3162
rect 3130 4012 3164 4046
rect 3202 4012 3236 4046
rect 3130 3944 3164 3978
rect 3202 3944 3236 3978
rect 3130 3876 3164 3910
rect 3202 3876 3236 3910
rect 3130 3808 3164 3842
rect 3202 3808 3236 3842
rect 3130 3740 3164 3774
rect 3202 3740 3236 3774
rect 3130 3672 3164 3706
rect 3202 3672 3236 3706
rect 3130 3604 3164 3638
rect 3202 3604 3236 3638
rect 3130 3536 3164 3570
rect 3202 3536 3236 3570
rect 3130 3468 3164 3502
rect 3202 3468 3236 3502
rect 3130 3400 3164 3434
rect 3202 3400 3236 3434
rect 3130 3332 3164 3366
rect 3202 3332 3236 3366
rect 3130 3264 3164 3298
rect 3202 3264 3236 3298
rect 3130 3196 3164 3230
rect 3202 3196 3236 3230
rect 3130 3128 3164 3162
rect 3202 3128 3236 3162
rect 3560 4012 3594 4046
rect 3764 4012 3798 4046
rect 3560 3944 3594 3978
rect 3764 3944 3798 3978
rect 3560 3876 3594 3910
rect 3764 3876 3798 3910
rect 3560 3808 3594 3842
rect 3764 3808 3798 3842
rect 3560 3740 3594 3774
rect 3764 3740 3798 3774
rect 3560 3672 3594 3706
rect 3764 3672 3798 3706
rect 3560 3604 3594 3638
rect 3764 3604 3798 3638
rect 3560 3536 3594 3570
rect 3764 3536 3798 3570
rect 3560 3468 3594 3502
rect 3764 3468 3798 3502
rect 3560 3400 3594 3434
rect 3764 3400 3798 3434
rect 3560 3332 3594 3366
rect 3764 3332 3798 3366
rect 3560 3264 3594 3298
rect 3764 3264 3798 3298
rect 3560 3196 3594 3230
rect 3764 3196 3798 3230
rect 3560 3128 3594 3162
rect 3764 3128 3798 3162
rect 4122 4012 4156 4046
rect 4194 4012 4228 4046
rect 4122 3944 4156 3978
rect 4194 3944 4228 3978
rect 4122 3876 4156 3910
rect 4194 3876 4228 3910
rect 4122 3808 4156 3842
rect 4194 3808 4228 3842
rect 4122 3740 4156 3774
rect 4194 3740 4228 3774
rect 4122 3672 4156 3706
rect 4194 3672 4228 3706
rect 4122 3604 4156 3638
rect 4194 3604 4228 3638
rect 4122 3536 4156 3570
rect 4194 3536 4228 3570
rect 4122 3468 4156 3502
rect 4194 3468 4228 3502
rect 4122 3400 4156 3434
rect 4194 3400 4228 3434
rect 4122 3332 4156 3366
rect 4194 3332 4228 3366
rect 4122 3264 4156 3298
rect 4194 3264 4228 3298
rect 4122 3196 4156 3230
rect 4194 3196 4228 3230
rect 4122 3128 4156 3162
rect 4194 3128 4228 3162
rect 4552 4012 4586 4046
rect 4756 4012 4790 4046
rect 4552 3944 4586 3978
rect 4756 3944 4790 3978
rect 4552 3876 4586 3910
rect 4756 3876 4790 3910
rect 4552 3808 4586 3842
rect 4756 3808 4790 3842
rect 4552 3740 4586 3774
rect 4756 3740 4790 3774
rect 4552 3672 4586 3706
rect 4756 3672 4790 3706
rect 4552 3604 4586 3638
rect 4756 3604 4790 3638
rect 4552 3536 4586 3570
rect 4756 3536 4790 3570
rect 4552 3468 4586 3502
rect 4756 3468 4790 3502
rect 4552 3400 4586 3434
rect 4756 3400 4790 3434
rect 4552 3332 4586 3366
rect 4756 3332 4790 3366
rect 4552 3264 4586 3298
rect 4756 3264 4790 3298
rect 4552 3196 4586 3230
rect 4756 3196 4790 3230
rect 4552 3128 4586 3162
rect 4756 3128 4790 3162
rect 5114 4012 5148 4046
rect 5186 4012 5220 4046
rect 5114 3944 5148 3978
rect 5186 3944 5220 3978
rect 5114 3876 5148 3910
rect 5186 3876 5220 3910
rect 5114 3808 5148 3842
rect 5186 3808 5220 3842
rect 5114 3740 5148 3774
rect 5186 3740 5220 3774
rect 5114 3672 5148 3706
rect 5186 3672 5220 3706
rect 5114 3604 5148 3638
rect 5186 3604 5220 3638
rect 5114 3536 5148 3570
rect 5186 3536 5220 3570
rect 5114 3468 5148 3502
rect 5186 3468 5220 3502
rect 5114 3400 5148 3434
rect 5186 3400 5220 3434
rect 5114 3332 5148 3366
rect 5186 3332 5220 3366
rect 5114 3264 5148 3298
rect 5186 3264 5220 3298
rect 5114 3196 5148 3230
rect 5186 3196 5220 3230
rect 5114 3128 5148 3162
rect 5186 3128 5220 3162
rect 5544 4012 5578 4046
rect 5748 4012 5782 4046
rect 5544 3944 5578 3978
rect 5748 3944 5782 3978
rect 5544 3876 5578 3910
rect 5748 3876 5782 3910
rect 5544 3808 5578 3842
rect 5748 3808 5782 3842
rect 5544 3740 5578 3774
rect 5748 3740 5782 3774
rect 5544 3672 5578 3706
rect 5748 3672 5782 3706
rect 5544 3604 5578 3638
rect 5748 3604 5782 3638
rect 5544 3536 5578 3570
rect 5748 3536 5782 3570
rect 5544 3468 5578 3502
rect 5748 3468 5782 3502
rect 5544 3400 5578 3434
rect 5748 3400 5782 3434
rect 5544 3332 5578 3366
rect 5748 3332 5782 3366
rect 5544 3264 5578 3298
rect 5748 3264 5782 3298
rect 5544 3196 5578 3230
rect 5748 3196 5782 3230
rect 5544 3128 5578 3162
rect 5748 3128 5782 3162
rect 6106 4012 6140 4046
rect 6178 4012 6212 4046
rect 6106 3944 6140 3978
rect 6178 3944 6212 3978
rect 6106 3876 6140 3910
rect 6178 3876 6212 3910
rect 6106 3808 6140 3842
rect 6178 3808 6212 3842
rect 6106 3740 6140 3774
rect 6178 3740 6212 3774
rect 6106 3672 6140 3706
rect 6178 3672 6212 3706
rect 6106 3604 6140 3638
rect 6178 3604 6212 3638
rect 6106 3536 6140 3570
rect 6178 3536 6212 3570
rect 6106 3468 6140 3502
rect 6178 3468 6212 3502
rect 6106 3400 6140 3434
rect 6178 3400 6212 3434
rect 6106 3332 6140 3366
rect 6178 3332 6212 3366
rect 6106 3264 6140 3298
rect 6178 3264 6212 3298
rect 6106 3196 6140 3230
rect 6178 3196 6212 3230
rect 6106 3128 6140 3162
rect 6178 3128 6212 3162
rect 6536 4012 6570 4046
rect 6740 4012 6774 4046
rect 6536 3944 6570 3978
rect 6740 3944 6774 3978
rect 6536 3876 6570 3910
rect 6740 3876 6774 3910
rect 6536 3808 6570 3842
rect 6740 3808 6774 3842
rect 6536 3740 6570 3774
rect 6740 3740 6774 3774
rect 6536 3672 6570 3706
rect 6740 3672 6774 3706
rect 6536 3604 6570 3638
rect 6740 3604 6774 3638
rect 6536 3536 6570 3570
rect 6740 3536 6774 3570
rect 6536 3468 6570 3502
rect 6740 3468 6774 3502
rect 6536 3400 6570 3434
rect 6740 3400 6774 3434
rect 6536 3332 6570 3366
rect 6740 3332 6774 3366
rect 6536 3264 6570 3298
rect 6740 3264 6774 3298
rect 6536 3196 6570 3230
rect 6740 3196 6774 3230
rect 6536 3128 6570 3162
rect 6740 3128 6774 3162
rect 7098 4012 7132 4046
rect 7170 4012 7204 4046
rect 7098 3944 7132 3978
rect 7170 3944 7204 3978
rect 7098 3876 7132 3910
rect 7170 3876 7204 3910
rect 7098 3808 7132 3842
rect 7170 3808 7204 3842
rect 7098 3740 7132 3774
rect 7170 3740 7204 3774
rect 7098 3672 7132 3706
rect 7170 3672 7204 3706
rect 7098 3604 7132 3638
rect 7170 3604 7204 3638
rect 7098 3536 7132 3570
rect 7170 3536 7204 3570
rect 7098 3468 7132 3502
rect 7170 3468 7204 3502
rect 7098 3400 7132 3434
rect 7170 3400 7204 3434
rect 7098 3332 7132 3366
rect 7170 3332 7204 3366
rect 7098 3264 7132 3298
rect 7170 3264 7204 3298
rect 7098 3196 7132 3230
rect 7170 3196 7204 3230
rect 7098 3128 7132 3162
rect 7170 3128 7204 3162
rect 7528 4012 7562 4046
rect 7732 4012 7766 4046
rect 7528 3944 7562 3978
rect 7732 3944 7766 3978
rect 7528 3876 7562 3910
rect 7732 3876 7766 3910
rect 7528 3808 7562 3842
rect 7732 3808 7766 3842
rect 7528 3740 7562 3774
rect 7732 3740 7766 3774
rect 7528 3672 7562 3706
rect 7732 3672 7766 3706
rect 7528 3604 7562 3638
rect 7732 3604 7766 3638
rect 7528 3536 7562 3570
rect 7732 3536 7766 3570
rect 7528 3468 7562 3502
rect 7732 3468 7766 3502
rect 7528 3400 7562 3434
rect 7732 3400 7766 3434
rect 7528 3332 7562 3366
rect 7732 3332 7766 3366
rect 7528 3264 7562 3298
rect 7732 3264 7766 3298
rect 7528 3196 7562 3230
rect 7732 3196 7766 3230
rect 7528 3128 7562 3162
rect 7732 3128 7766 3162
rect 8090 4012 8124 4046
rect 8162 4012 8196 4046
rect 8090 3944 8124 3978
rect 8162 3944 8196 3978
rect 8090 3876 8124 3910
rect 8162 3876 8196 3910
rect 8090 3808 8124 3842
rect 8162 3808 8196 3842
rect 8090 3740 8124 3774
rect 8162 3740 8196 3774
rect 8090 3672 8124 3706
rect 8162 3672 8196 3706
rect 8090 3604 8124 3638
rect 8162 3604 8196 3638
rect 8090 3536 8124 3570
rect 8162 3536 8196 3570
rect 8090 3468 8124 3502
rect 8162 3468 8196 3502
rect 8090 3400 8124 3434
rect 8162 3400 8196 3434
rect 8090 3332 8124 3366
rect 8162 3332 8196 3366
rect 8090 3264 8124 3298
rect 8162 3264 8196 3298
rect 8090 3196 8124 3230
rect 8162 3196 8196 3230
rect 8090 3128 8124 3162
rect 8162 3128 8196 3162
rect 8520 4012 8554 4046
rect 8724 4012 8758 4046
rect 8520 3944 8554 3978
rect 8724 3944 8758 3978
rect 8520 3876 8554 3910
rect 8724 3876 8758 3910
rect 8520 3808 8554 3842
rect 8724 3808 8758 3842
rect 8520 3740 8554 3774
rect 8724 3740 8758 3774
rect 8520 3672 8554 3706
rect 8724 3672 8758 3706
rect 8520 3604 8554 3638
rect 8724 3604 8758 3638
rect 8520 3536 8554 3570
rect 8724 3536 8758 3570
rect 8520 3468 8554 3502
rect 8724 3468 8758 3502
rect 8520 3400 8554 3434
rect 8724 3400 8758 3434
rect 8520 3332 8554 3366
rect 8724 3332 8758 3366
rect 8520 3264 8554 3298
rect 8724 3264 8758 3298
rect 8520 3196 8554 3230
rect 8724 3196 8758 3230
rect 8520 3128 8554 3162
rect 8724 3128 8758 3162
rect 9082 4012 9116 4046
rect 9154 4012 9188 4046
rect 9082 3944 9116 3978
rect 9154 3944 9188 3978
rect 9082 3876 9116 3910
rect 9154 3876 9188 3910
rect 9082 3808 9116 3842
rect 9154 3808 9188 3842
rect 9082 3740 9116 3774
rect 9154 3740 9188 3774
rect 9082 3672 9116 3706
rect 9154 3672 9188 3706
rect 9082 3604 9116 3638
rect 9154 3604 9188 3638
rect 9082 3536 9116 3570
rect 9154 3536 9188 3570
rect 9082 3468 9116 3502
rect 9154 3468 9188 3502
rect 9082 3400 9116 3434
rect 9154 3400 9188 3434
rect 9082 3332 9116 3366
rect 9154 3332 9188 3366
rect 9082 3264 9116 3298
rect 9154 3264 9188 3298
rect 9082 3196 9116 3230
rect 9154 3196 9188 3230
rect 9082 3128 9116 3162
rect 9154 3128 9188 3162
rect 9512 4012 9546 4046
rect 9716 4012 9750 4046
rect 9512 3944 9546 3978
rect 9716 3944 9750 3978
rect 9512 3876 9546 3910
rect 9716 3876 9750 3910
rect 9512 3808 9546 3842
rect 9716 3808 9750 3842
rect 9512 3740 9546 3774
rect 9716 3740 9750 3774
rect 9512 3672 9546 3706
rect 9716 3672 9750 3706
rect 9512 3604 9546 3638
rect 9716 3604 9750 3638
rect 9512 3536 9546 3570
rect 9716 3536 9750 3570
rect 9512 3468 9546 3502
rect 9716 3468 9750 3502
rect 9512 3400 9546 3434
rect 9716 3400 9750 3434
rect 9512 3332 9546 3366
rect 9716 3332 9750 3366
rect 9512 3264 9546 3298
rect 9716 3264 9750 3298
rect 9512 3196 9546 3230
rect 9716 3196 9750 3230
rect 9512 3128 9546 3162
rect 9716 3128 9750 3162
rect 10074 4012 10108 4046
rect 10146 4012 10180 4046
rect 10074 3944 10108 3978
rect 10146 3944 10180 3978
rect 10074 3876 10108 3910
rect 10146 3876 10180 3910
rect 10074 3808 10108 3842
rect 10146 3808 10180 3842
rect 10074 3740 10108 3774
rect 10146 3740 10180 3774
rect 10074 3672 10108 3706
rect 10146 3672 10180 3706
rect 10074 3604 10108 3638
rect 10146 3604 10180 3638
rect 10074 3536 10108 3570
rect 10146 3536 10180 3570
rect 10074 3468 10108 3502
rect 10146 3468 10180 3502
rect 10074 3400 10108 3434
rect 10146 3400 10180 3434
rect 10074 3332 10108 3366
rect 10146 3332 10180 3366
rect 10074 3264 10108 3298
rect 10146 3264 10180 3298
rect 10074 3196 10108 3230
rect 10146 3196 10180 3230
rect 10074 3128 10108 3162
rect 10146 3128 10180 3162
rect 10504 4012 10538 4046
rect 10708 4012 10742 4046
rect 10504 3944 10538 3978
rect 10708 3944 10742 3978
rect 10504 3876 10538 3910
rect 10708 3876 10742 3910
rect 10504 3808 10538 3842
rect 10708 3808 10742 3842
rect 10504 3740 10538 3774
rect 10708 3740 10742 3774
rect 10504 3672 10538 3706
rect 10708 3672 10742 3706
rect 10504 3604 10538 3638
rect 10708 3604 10742 3638
rect 10504 3536 10538 3570
rect 10708 3536 10742 3570
rect 10504 3468 10538 3502
rect 10708 3468 10742 3502
rect 10504 3400 10538 3434
rect 10708 3400 10742 3434
rect 10504 3332 10538 3366
rect 10708 3332 10742 3366
rect 10504 3264 10538 3298
rect 10708 3264 10742 3298
rect 10504 3196 10538 3230
rect 10708 3196 10742 3230
rect 10504 3128 10538 3162
rect 10708 3128 10742 3162
rect 11066 4012 11100 4046
rect 11138 4012 11172 4046
rect 11066 3944 11100 3978
rect 11138 3944 11172 3978
rect 11066 3876 11100 3910
rect 11138 3876 11172 3910
rect 11066 3808 11100 3842
rect 11138 3808 11172 3842
rect 11066 3740 11100 3774
rect 11138 3740 11172 3774
rect 11066 3672 11100 3706
rect 11138 3672 11172 3706
rect 11066 3604 11100 3638
rect 11138 3604 11172 3638
rect 11066 3536 11100 3570
rect 11138 3536 11172 3570
rect 11066 3468 11100 3502
rect 11138 3468 11172 3502
rect 11066 3400 11100 3434
rect 11138 3400 11172 3434
rect 11066 3332 11100 3366
rect 11138 3332 11172 3366
rect 11066 3264 11100 3298
rect 11138 3264 11172 3298
rect 11066 3196 11100 3230
rect 11138 3196 11172 3230
rect 11066 3128 11100 3162
rect 11138 3128 11172 3162
rect 11496 4012 11530 4046
rect 11700 4012 11734 4046
rect 11496 3944 11530 3978
rect 11700 3944 11734 3978
rect 11496 3876 11530 3910
rect 11700 3876 11734 3910
rect 11496 3808 11530 3842
rect 11700 3808 11734 3842
rect 11496 3740 11530 3774
rect 11700 3740 11734 3774
rect 11496 3672 11530 3706
rect 11700 3672 11734 3706
rect 11496 3604 11530 3638
rect 11700 3604 11734 3638
rect 11496 3536 11530 3570
rect 11700 3536 11734 3570
rect 11496 3468 11530 3502
rect 11700 3468 11734 3502
rect 11496 3400 11530 3434
rect 11700 3400 11734 3434
rect 11496 3332 11530 3366
rect 11700 3332 11734 3366
rect 11496 3264 11530 3298
rect 11700 3264 11734 3298
rect 11496 3196 11530 3230
rect 11700 3196 11734 3230
rect 11496 3128 11530 3162
rect 11700 3128 11734 3162
rect 12058 4012 12092 4046
rect 12130 4012 12164 4046
rect 12058 3944 12092 3978
rect 12130 3944 12164 3978
rect 12058 3876 12092 3910
rect 12130 3876 12164 3910
rect 12058 3808 12092 3842
rect 12130 3808 12164 3842
rect 12058 3740 12092 3774
rect 12130 3740 12164 3774
rect 12058 3672 12092 3706
rect 12130 3672 12164 3706
rect 12058 3604 12092 3638
rect 12130 3604 12164 3638
rect 12058 3536 12092 3570
rect 12130 3536 12164 3570
rect 12058 3468 12092 3502
rect 12130 3468 12164 3502
rect 12058 3400 12092 3434
rect 12130 3400 12164 3434
rect 12058 3332 12092 3366
rect 12130 3332 12164 3366
rect 12058 3264 12092 3298
rect 12130 3264 12164 3298
rect 12058 3196 12092 3230
rect 12130 3196 12164 3230
rect 12058 3128 12092 3162
rect 12130 3128 12164 3162
rect 12488 4012 12522 4046
rect 12692 4012 12726 4046
rect 12488 3944 12522 3978
rect 12692 3944 12726 3978
rect 12488 3876 12522 3910
rect 12692 3876 12726 3910
rect 12488 3808 12522 3842
rect 12692 3808 12726 3842
rect 12488 3740 12522 3774
rect 12692 3740 12726 3774
rect 12488 3672 12522 3706
rect 12692 3672 12726 3706
rect 12488 3604 12522 3638
rect 12692 3604 12726 3638
rect 12488 3536 12522 3570
rect 12692 3536 12726 3570
rect 12488 3468 12522 3502
rect 12692 3468 12726 3502
rect 12488 3400 12522 3434
rect 12692 3400 12726 3434
rect 12488 3332 12522 3366
rect 12692 3332 12726 3366
rect 12488 3264 12522 3298
rect 12692 3264 12726 3298
rect 12488 3196 12522 3230
rect 12692 3196 12726 3230
rect 12488 3128 12522 3162
rect 12692 3128 12726 3162
rect 13050 4012 13084 4046
rect 13122 4012 13156 4046
rect 13050 3944 13084 3978
rect 13122 3944 13156 3978
rect 13050 3876 13084 3910
rect 13122 3876 13156 3910
rect 13050 3808 13084 3842
rect 13122 3808 13156 3842
rect 13050 3740 13084 3774
rect 13122 3740 13156 3774
rect 13050 3672 13084 3706
rect 13122 3672 13156 3706
rect 13050 3604 13084 3638
rect 13122 3604 13156 3638
rect 13050 3536 13084 3570
rect 13122 3536 13156 3570
rect 13050 3468 13084 3502
rect 13122 3468 13156 3502
rect 13050 3400 13084 3434
rect 13122 3400 13156 3434
rect 13050 3332 13084 3366
rect 13122 3332 13156 3366
rect 13050 3264 13084 3298
rect 13122 3264 13156 3298
rect 13050 3196 13084 3230
rect 13122 3196 13156 3230
rect 13050 3128 13084 3162
rect 13122 3128 13156 3162
rect 13480 4012 13514 4046
rect 13684 4012 13718 4046
rect 13480 3944 13514 3978
rect 13684 3944 13718 3978
rect 13480 3876 13514 3910
rect 13684 3876 13718 3910
rect 13480 3808 13514 3842
rect 13684 3808 13718 3842
rect 13480 3740 13514 3774
rect 13684 3740 13718 3774
rect 13480 3672 13514 3706
rect 13684 3672 13718 3706
rect 13480 3604 13514 3638
rect 13684 3604 13718 3638
rect 13480 3536 13514 3570
rect 13684 3536 13718 3570
rect 13480 3468 13514 3502
rect 13684 3468 13718 3502
rect 13480 3400 13514 3434
rect 13684 3400 13718 3434
rect 13480 3332 13514 3366
rect 13684 3332 13718 3366
rect 13480 3264 13514 3298
rect 13684 3264 13718 3298
rect 13480 3196 13514 3230
rect 13684 3196 13718 3230
rect 13480 3128 13514 3162
rect 13684 3128 13718 3162
rect 14042 4012 14076 4046
rect 14042 3944 14076 3978
rect 14042 3876 14076 3910
rect 14042 3808 14076 3842
rect 14042 3740 14076 3774
rect 14042 3672 14076 3706
rect 14042 3604 14076 3638
rect 14042 3536 14076 3570
rect 14042 3468 14076 3502
rect 14042 3400 14076 3434
rect 14042 3332 14076 3366
rect 14042 3264 14076 3298
rect 14042 3196 14076 3230
rect 14042 3128 14076 3162
rect 14386 4012 14420 4046
rect 14386 3944 14420 3978
rect 14386 3876 14420 3910
rect 14386 3808 14420 3842
rect 14386 3740 14420 3774
rect 14386 3672 14420 3706
rect 14386 3604 14420 3638
rect 14386 3536 14420 3570
rect 14386 3468 14420 3502
rect 14386 3400 14420 3434
rect 14386 3332 14420 3366
rect 14386 3264 14420 3298
rect 14386 3196 14420 3230
rect 14386 3128 14420 3162
rect 802 2411 836 2445
rect 802 2343 836 2377
rect 802 2275 836 2309
rect 802 2207 836 2241
rect 802 2139 836 2173
rect 802 2071 836 2105
rect 802 2003 836 2037
rect 802 1935 836 1969
rect 802 1867 836 1901
rect 802 1799 836 1833
rect 802 1731 836 1765
rect 802 1663 836 1697
rect 802 1595 836 1629
rect 802 1527 836 1561
rect 1146 2411 1180 2445
rect 1218 2411 1252 2445
rect 1146 2343 1180 2377
rect 1218 2343 1252 2377
rect 1146 2275 1180 2309
rect 1218 2275 1252 2309
rect 1146 2207 1180 2241
rect 1218 2207 1252 2241
rect 1146 2139 1180 2173
rect 1218 2139 1252 2173
rect 1146 2071 1180 2105
rect 1218 2071 1252 2105
rect 1146 2003 1180 2037
rect 1218 2003 1252 2037
rect 1146 1935 1180 1969
rect 1218 1935 1252 1969
rect 1146 1867 1180 1901
rect 1218 1867 1252 1901
rect 1146 1799 1180 1833
rect 1218 1799 1252 1833
rect 1146 1731 1180 1765
rect 1218 1731 1252 1765
rect 1146 1663 1180 1697
rect 1218 1663 1252 1697
rect 1146 1595 1180 1629
rect 1218 1595 1252 1629
rect 1146 1527 1180 1561
rect 1218 1527 1252 1561
rect 1576 2411 1610 2445
rect 1780 2411 1814 2445
rect 1576 2343 1610 2377
rect 1780 2343 1814 2377
rect 1576 2275 1610 2309
rect 1780 2275 1814 2309
rect 1576 2207 1610 2241
rect 1780 2207 1814 2241
rect 1576 2139 1610 2173
rect 1780 2139 1814 2173
rect 1576 2071 1610 2105
rect 1780 2071 1814 2105
rect 1576 2003 1610 2037
rect 1780 2003 1814 2037
rect 1576 1935 1610 1969
rect 1780 1935 1814 1969
rect 1576 1867 1610 1901
rect 1780 1867 1814 1901
rect 1576 1799 1610 1833
rect 1780 1799 1814 1833
rect 1576 1731 1610 1765
rect 1780 1731 1814 1765
rect 1576 1663 1610 1697
rect 1780 1663 1814 1697
rect 1576 1595 1610 1629
rect 1780 1595 1814 1629
rect 1576 1527 1610 1561
rect 1780 1527 1814 1561
rect 2138 2411 2172 2445
rect 2210 2411 2244 2445
rect 2138 2343 2172 2377
rect 2210 2343 2244 2377
rect 2138 2275 2172 2309
rect 2210 2275 2244 2309
rect 2138 2207 2172 2241
rect 2210 2207 2244 2241
rect 2138 2139 2172 2173
rect 2210 2139 2244 2173
rect 2138 2071 2172 2105
rect 2210 2071 2244 2105
rect 2138 2003 2172 2037
rect 2210 2003 2244 2037
rect 2138 1935 2172 1969
rect 2210 1935 2244 1969
rect 2138 1867 2172 1901
rect 2210 1867 2244 1901
rect 2138 1799 2172 1833
rect 2210 1799 2244 1833
rect 2138 1731 2172 1765
rect 2210 1731 2244 1765
rect 2138 1663 2172 1697
rect 2210 1663 2244 1697
rect 2138 1595 2172 1629
rect 2210 1595 2244 1629
rect 2138 1527 2172 1561
rect 2210 1527 2244 1561
rect 2568 2411 2602 2445
rect 2772 2411 2806 2445
rect 2568 2343 2602 2377
rect 2772 2343 2806 2377
rect 2568 2275 2602 2309
rect 2772 2275 2806 2309
rect 2568 2207 2602 2241
rect 2772 2207 2806 2241
rect 2568 2139 2602 2173
rect 2772 2139 2806 2173
rect 2568 2071 2602 2105
rect 2772 2071 2806 2105
rect 2568 2003 2602 2037
rect 2772 2003 2806 2037
rect 2568 1935 2602 1969
rect 2772 1935 2806 1969
rect 2568 1867 2602 1901
rect 2772 1867 2806 1901
rect 2568 1799 2602 1833
rect 2772 1799 2806 1833
rect 2568 1731 2602 1765
rect 2772 1731 2806 1765
rect 2568 1663 2602 1697
rect 2772 1663 2806 1697
rect 2568 1595 2602 1629
rect 2772 1595 2806 1629
rect 2568 1527 2602 1561
rect 2772 1527 2806 1561
rect 3130 2411 3164 2445
rect 3202 2411 3236 2445
rect 3130 2343 3164 2377
rect 3202 2343 3236 2377
rect 3130 2275 3164 2309
rect 3202 2275 3236 2309
rect 3130 2207 3164 2241
rect 3202 2207 3236 2241
rect 3130 2139 3164 2173
rect 3202 2139 3236 2173
rect 3130 2071 3164 2105
rect 3202 2071 3236 2105
rect 3130 2003 3164 2037
rect 3202 2003 3236 2037
rect 3130 1935 3164 1969
rect 3202 1935 3236 1969
rect 3130 1867 3164 1901
rect 3202 1867 3236 1901
rect 3130 1799 3164 1833
rect 3202 1799 3236 1833
rect 3130 1731 3164 1765
rect 3202 1731 3236 1765
rect 3130 1663 3164 1697
rect 3202 1663 3236 1697
rect 3130 1595 3164 1629
rect 3202 1595 3236 1629
rect 3130 1527 3164 1561
rect 3202 1527 3236 1561
rect 3560 2411 3594 2445
rect 3764 2411 3798 2445
rect 3560 2343 3594 2377
rect 3764 2343 3798 2377
rect 3560 2275 3594 2309
rect 3764 2275 3798 2309
rect 3560 2207 3594 2241
rect 3764 2207 3798 2241
rect 3560 2139 3594 2173
rect 3764 2139 3798 2173
rect 3560 2071 3594 2105
rect 3764 2071 3798 2105
rect 3560 2003 3594 2037
rect 3764 2003 3798 2037
rect 3560 1935 3594 1969
rect 3764 1935 3798 1969
rect 3560 1867 3594 1901
rect 3764 1867 3798 1901
rect 3560 1799 3594 1833
rect 3764 1799 3798 1833
rect 3560 1731 3594 1765
rect 3764 1731 3798 1765
rect 3560 1663 3594 1697
rect 3764 1663 3798 1697
rect 3560 1595 3594 1629
rect 3764 1595 3798 1629
rect 3560 1527 3594 1561
rect 3764 1527 3798 1561
rect 4122 2411 4156 2445
rect 4194 2411 4228 2445
rect 4122 2343 4156 2377
rect 4194 2343 4228 2377
rect 4122 2275 4156 2309
rect 4194 2275 4228 2309
rect 4122 2207 4156 2241
rect 4194 2207 4228 2241
rect 4122 2139 4156 2173
rect 4194 2139 4228 2173
rect 4122 2071 4156 2105
rect 4194 2071 4228 2105
rect 4122 2003 4156 2037
rect 4194 2003 4228 2037
rect 4122 1935 4156 1969
rect 4194 1935 4228 1969
rect 4122 1867 4156 1901
rect 4194 1867 4228 1901
rect 4122 1799 4156 1833
rect 4194 1799 4228 1833
rect 4122 1731 4156 1765
rect 4194 1731 4228 1765
rect 4122 1663 4156 1697
rect 4194 1663 4228 1697
rect 4122 1595 4156 1629
rect 4194 1595 4228 1629
rect 4122 1527 4156 1561
rect 4194 1527 4228 1561
rect 4552 2411 4586 2445
rect 4756 2411 4790 2445
rect 4552 2343 4586 2377
rect 4756 2343 4790 2377
rect 4552 2275 4586 2309
rect 4756 2275 4790 2309
rect 4552 2207 4586 2241
rect 4756 2207 4790 2241
rect 4552 2139 4586 2173
rect 4756 2139 4790 2173
rect 4552 2071 4586 2105
rect 4756 2071 4790 2105
rect 4552 2003 4586 2037
rect 4756 2003 4790 2037
rect 4552 1935 4586 1969
rect 4756 1935 4790 1969
rect 4552 1867 4586 1901
rect 4756 1867 4790 1901
rect 4552 1799 4586 1833
rect 4756 1799 4790 1833
rect 4552 1731 4586 1765
rect 4756 1731 4790 1765
rect 4552 1663 4586 1697
rect 4756 1663 4790 1697
rect 4552 1595 4586 1629
rect 4756 1595 4790 1629
rect 4552 1527 4586 1561
rect 4756 1527 4790 1561
rect 5114 2411 5148 2445
rect 5186 2411 5220 2445
rect 5114 2343 5148 2377
rect 5186 2343 5220 2377
rect 5114 2275 5148 2309
rect 5186 2275 5220 2309
rect 5114 2207 5148 2241
rect 5186 2207 5220 2241
rect 5114 2139 5148 2173
rect 5186 2139 5220 2173
rect 5114 2071 5148 2105
rect 5186 2071 5220 2105
rect 5114 2003 5148 2037
rect 5186 2003 5220 2037
rect 5114 1935 5148 1969
rect 5186 1935 5220 1969
rect 5114 1867 5148 1901
rect 5186 1867 5220 1901
rect 5114 1799 5148 1833
rect 5186 1799 5220 1833
rect 5114 1731 5148 1765
rect 5186 1731 5220 1765
rect 5114 1663 5148 1697
rect 5186 1663 5220 1697
rect 5114 1595 5148 1629
rect 5186 1595 5220 1629
rect 5114 1527 5148 1561
rect 5186 1527 5220 1561
rect 5544 2411 5578 2445
rect 5748 2411 5782 2445
rect 5544 2343 5578 2377
rect 5748 2343 5782 2377
rect 5544 2275 5578 2309
rect 5748 2275 5782 2309
rect 5544 2207 5578 2241
rect 5748 2207 5782 2241
rect 5544 2139 5578 2173
rect 5748 2139 5782 2173
rect 5544 2071 5578 2105
rect 5748 2071 5782 2105
rect 5544 2003 5578 2037
rect 5748 2003 5782 2037
rect 5544 1935 5578 1969
rect 5748 1935 5782 1969
rect 5544 1867 5578 1901
rect 5748 1867 5782 1901
rect 5544 1799 5578 1833
rect 5748 1799 5782 1833
rect 5544 1731 5578 1765
rect 5748 1731 5782 1765
rect 5544 1663 5578 1697
rect 5748 1663 5782 1697
rect 5544 1595 5578 1629
rect 5748 1595 5782 1629
rect 5544 1527 5578 1561
rect 5748 1527 5782 1561
rect 6106 2411 6140 2445
rect 6178 2411 6212 2445
rect 6106 2343 6140 2377
rect 6178 2343 6212 2377
rect 6106 2275 6140 2309
rect 6178 2275 6212 2309
rect 6106 2207 6140 2241
rect 6178 2207 6212 2241
rect 6106 2139 6140 2173
rect 6178 2139 6212 2173
rect 6106 2071 6140 2105
rect 6178 2071 6212 2105
rect 6106 2003 6140 2037
rect 6178 2003 6212 2037
rect 6106 1935 6140 1969
rect 6178 1935 6212 1969
rect 6106 1867 6140 1901
rect 6178 1867 6212 1901
rect 6106 1799 6140 1833
rect 6178 1799 6212 1833
rect 6106 1731 6140 1765
rect 6178 1731 6212 1765
rect 6106 1663 6140 1697
rect 6178 1663 6212 1697
rect 6106 1595 6140 1629
rect 6178 1595 6212 1629
rect 6106 1527 6140 1561
rect 6178 1527 6212 1561
rect 6536 2411 6570 2445
rect 6740 2411 6774 2445
rect 6536 2343 6570 2377
rect 6740 2343 6774 2377
rect 6536 2275 6570 2309
rect 6740 2275 6774 2309
rect 6536 2207 6570 2241
rect 6740 2207 6774 2241
rect 6536 2139 6570 2173
rect 6740 2139 6774 2173
rect 6536 2071 6570 2105
rect 6740 2071 6774 2105
rect 6536 2003 6570 2037
rect 6740 2003 6774 2037
rect 6536 1935 6570 1969
rect 6740 1935 6774 1969
rect 6536 1867 6570 1901
rect 6740 1867 6774 1901
rect 6536 1799 6570 1833
rect 6740 1799 6774 1833
rect 6536 1731 6570 1765
rect 6740 1731 6774 1765
rect 6536 1663 6570 1697
rect 6740 1663 6774 1697
rect 6536 1595 6570 1629
rect 6740 1595 6774 1629
rect 6536 1527 6570 1561
rect 6740 1527 6774 1561
rect 7098 2411 7132 2445
rect 7170 2411 7204 2445
rect 7098 2343 7132 2377
rect 7170 2343 7204 2377
rect 7098 2275 7132 2309
rect 7170 2275 7204 2309
rect 7098 2207 7132 2241
rect 7170 2207 7204 2241
rect 7098 2139 7132 2173
rect 7170 2139 7204 2173
rect 7098 2071 7132 2105
rect 7170 2071 7204 2105
rect 7098 2003 7132 2037
rect 7170 2003 7204 2037
rect 7098 1935 7132 1969
rect 7170 1935 7204 1969
rect 7098 1867 7132 1901
rect 7170 1867 7204 1901
rect 7098 1799 7132 1833
rect 7170 1799 7204 1833
rect 7098 1731 7132 1765
rect 7170 1731 7204 1765
rect 7098 1663 7132 1697
rect 7170 1663 7204 1697
rect 7098 1595 7132 1629
rect 7170 1595 7204 1629
rect 7098 1527 7132 1561
rect 7170 1527 7204 1561
rect 7528 2411 7562 2445
rect 7732 2411 7766 2445
rect 7528 2343 7562 2377
rect 7732 2343 7766 2377
rect 7528 2275 7562 2309
rect 7732 2275 7766 2309
rect 7528 2207 7562 2241
rect 7732 2207 7766 2241
rect 7528 2139 7562 2173
rect 7732 2139 7766 2173
rect 7528 2071 7562 2105
rect 7732 2071 7766 2105
rect 7528 2003 7562 2037
rect 7732 2003 7766 2037
rect 7528 1935 7562 1969
rect 7732 1935 7766 1969
rect 7528 1867 7562 1901
rect 7732 1867 7766 1901
rect 7528 1799 7562 1833
rect 7732 1799 7766 1833
rect 7528 1731 7562 1765
rect 7732 1731 7766 1765
rect 7528 1663 7562 1697
rect 7732 1663 7766 1697
rect 7528 1595 7562 1629
rect 7732 1595 7766 1629
rect 7528 1527 7562 1561
rect 7732 1527 7766 1561
rect 8090 2411 8124 2445
rect 8162 2411 8196 2445
rect 8090 2343 8124 2377
rect 8162 2343 8196 2377
rect 8090 2275 8124 2309
rect 8162 2275 8196 2309
rect 8090 2207 8124 2241
rect 8162 2207 8196 2241
rect 8090 2139 8124 2173
rect 8162 2139 8196 2173
rect 8090 2071 8124 2105
rect 8162 2071 8196 2105
rect 8090 2003 8124 2037
rect 8162 2003 8196 2037
rect 8090 1935 8124 1969
rect 8162 1935 8196 1969
rect 8090 1867 8124 1901
rect 8162 1867 8196 1901
rect 8090 1799 8124 1833
rect 8162 1799 8196 1833
rect 8090 1731 8124 1765
rect 8162 1731 8196 1765
rect 8090 1663 8124 1697
rect 8162 1663 8196 1697
rect 8090 1595 8124 1629
rect 8162 1595 8196 1629
rect 8090 1527 8124 1561
rect 8162 1527 8196 1561
rect 8520 2411 8554 2445
rect 8724 2411 8758 2445
rect 8520 2343 8554 2377
rect 8724 2343 8758 2377
rect 8520 2275 8554 2309
rect 8724 2275 8758 2309
rect 8520 2207 8554 2241
rect 8724 2207 8758 2241
rect 8520 2139 8554 2173
rect 8724 2139 8758 2173
rect 8520 2071 8554 2105
rect 8724 2071 8758 2105
rect 8520 2003 8554 2037
rect 8724 2003 8758 2037
rect 8520 1935 8554 1969
rect 8724 1935 8758 1969
rect 8520 1867 8554 1901
rect 8724 1867 8758 1901
rect 8520 1799 8554 1833
rect 8724 1799 8758 1833
rect 8520 1731 8554 1765
rect 8724 1731 8758 1765
rect 8520 1663 8554 1697
rect 8724 1663 8758 1697
rect 8520 1595 8554 1629
rect 8724 1595 8758 1629
rect 8520 1527 8554 1561
rect 8724 1527 8758 1561
rect 9082 2411 9116 2445
rect 9154 2411 9188 2445
rect 9082 2343 9116 2377
rect 9154 2343 9188 2377
rect 9082 2275 9116 2309
rect 9154 2275 9188 2309
rect 9082 2207 9116 2241
rect 9154 2207 9188 2241
rect 9082 2139 9116 2173
rect 9154 2139 9188 2173
rect 9082 2071 9116 2105
rect 9154 2071 9188 2105
rect 9082 2003 9116 2037
rect 9154 2003 9188 2037
rect 9082 1935 9116 1969
rect 9154 1935 9188 1969
rect 9082 1867 9116 1901
rect 9154 1867 9188 1901
rect 9082 1799 9116 1833
rect 9154 1799 9188 1833
rect 9082 1731 9116 1765
rect 9154 1731 9188 1765
rect 9082 1663 9116 1697
rect 9154 1663 9188 1697
rect 9082 1595 9116 1629
rect 9154 1595 9188 1629
rect 9082 1527 9116 1561
rect 9154 1527 9188 1561
rect 9512 2411 9546 2445
rect 9716 2411 9750 2445
rect 9512 2343 9546 2377
rect 9716 2343 9750 2377
rect 9512 2275 9546 2309
rect 9716 2275 9750 2309
rect 9512 2207 9546 2241
rect 9716 2207 9750 2241
rect 9512 2139 9546 2173
rect 9716 2139 9750 2173
rect 9512 2071 9546 2105
rect 9716 2071 9750 2105
rect 9512 2003 9546 2037
rect 9716 2003 9750 2037
rect 9512 1935 9546 1969
rect 9716 1935 9750 1969
rect 9512 1867 9546 1901
rect 9716 1867 9750 1901
rect 9512 1799 9546 1833
rect 9716 1799 9750 1833
rect 9512 1731 9546 1765
rect 9716 1731 9750 1765
rect 9512 1663 9546 1697
rect 9716 1663 9750 1697
rect 9512 1595 9546 1629
rect 9716 1595 9750 1629
rect 9512 1527 9546 1561
rect 9716 1527 9750 1561
rect 10074 2411 10108 2445
rect 10146 2411 10180 2445
rect 10074 2343 10108 2377
rect 10146 2343 10180 2377
rect 10074 2275 10108 2309
rect 10146 2275 10180 2309
rect 10074 2207 10108 2241
rect 10146 2207 10180 2241
rect 10074 2139 10108 2173
rect 10146 2139 10180 2173
rect 10074 2071 10108 2105
rect 10146 2071 10180 2105
rect 10074 2003 10108 2037
rect 10146 2003 10180 2037
rect 10074 1935 10108 1969
rect 10146 1935 10180 1969
rect 10074 1867 10108 1901
rect 10146 1867 10180 1901
rect 10074 1799 10108 1833
rect 10146 1799 10180 1833
rect 10074 1731 10108 1765
rect 10146 1731 10180 1765
rect 10074 1663 10108 1697
rect 10146 1663 10180 1697
rect 10074 1595 10108 1629
rect 10146 1595 10180 1629
rect 10074 1527 10108 1561
rect 10146 1527 10180 1561
rect 10504 2411 10538 2445
rect 10708 2411 10742 2445
rect 10504 2343 10538 2377
rect 10708 2343 10742 2377
rect 10504 2275 10538 2309
rect 10708 2275 10742 2309
rect 10504 2207 10538 2241
rect 10708 2207 10742 2241
rect 10504 2139 10538 2173
rect 10708 2139 10742 2173
rect 10504 2071 10538 2105
rect 10708 2071 10742 2105
rect 10504 2003 10538 2037
rect 10708 2003 10742 2037
rect 10504 1935 10538 1969
rect 10708 1935 10742 1969
rect 10504 1867 10538 1901
rect 10708 1867 10742 1901
rect 10504 1799 10538 1833
rect 10708 1799 10742 1833
rect 10504 1731 10538 1765
rect 10708 1731 10742 1765
rect 10504 1663 10538 1697
rect 10708 1663 10742 1697
rect 10504 1595 10538 1629
rect 10708 1595 10742 1629
rect 10504 1527 10538 1561
rect 10708 1527 10742 1561
rect 11066 2411 11100 2445
rect 11138 2411 11172 2445
rect 11066 2343 11100 2377
rect 11138 2343 11172 2377
rect 11066 2275 11100 2309
rect 11138 2275 11172 2309
rect 11066 2207 11100 2241
rect 11138 2207 11172 2241
rect 11066 2139 11100 2173
rect 11138 2139 11172 2173
rect 11066 2071 11100 2105
rect 11138 2071 11172 2105
rect 11066 2003 11100 2037
rect 11138 2003 11172 2037
rect 11066 1935 11100 1969
rect 11138 1935 11172 1969
rect 11066 1867 11100 1901
rect 11138 1867 11172 1901
rect 11066 1799 11100 1833
rect 11138 1799 11172 1833
rect 11066 1731 11100 1765
rect 11138 1731 11172 1765
rect 11066 1663 11100 1697
rect 11138 1663 11172 1697
rect 11066 1595 11100 1629
rect 11138 1595 11172 1629
rect 11066 1527 11100 1561
rect 11138 1527 11172 1561
rect 11496 2411 11530 2445
rect 11700 2411 11734 2445
rect 11496 2343 11530 2377
rect 11700 2343 11734 2377
rect 11496 2275 11530 2309
rect 11700 2275 11734 2309
rect 11496 2207 11530 2241
rect 11700 2207 11734 2241
rect 11496 2139 11530 2173
rect 11700 2139 11734 2173
rect 11496 2071 11530 2105
rect 11700 2071 11734 2105
rect 11496 2003 11530 2037
rect 11700 2003 11734 2037
rect 11496 1935 11530 1969
rect 11700 1935 11734 1969
rect 11496 1867 11530 1901
rect 11700 1867 11734 1901
rect 11496 1799 11530 1833
rect 11700 1799 11734 1833
rect 11496 1731 11530 1765
rect 11700 1731 11734 1765
rect 11496 1663 11530 1697
rect 11700 1663 11734 1697
rect 11496 1595 11530 1629
rect 11700 1595 11734 1629
rect 11496 1527 11530 1561
rect 11700 1527 11734 1561
rect 12058 2411 12092 2445
rect 12130 2411 12164 2445
rect 12058 2343 12092 2377
rect 12130 2343 12164 2377
rect 12058 2275 12092 2309
rect 12130 2275 12164 2309
rect 12058 2207 12092 2241
rect 12130 2207 12164 2241
rect 12058 2139 12092 2173
rect 12130 2139 12164 2173
rect 12058 2071 12092 2105
rect 12130 2071 12164 2105
rect 12058 2003 12092 2037
rect 12130 2003 12164 2037
rect 12058 1935 12092 1969
rect 12130 1935 12164 1969
rect 12058 1867 12092 1901
rect 12130 1867 12164 1901
rect 12058 1799 12092 1833
rect 12130 1799 12164 1833
rect 12058 1731 12092 1765
rect 12130 1731 12164 1765
rect 12058 1663 12092 1697
rect 12130 1663 12164 1697
rect 12058 1595 12092 1629
rect 12130 1595 12164 1629
rect 12058 1527 12092 1561
rect 12130 1527 12164 1561
rect 12488 2411 12522 2445
rect 12692 2411 12726 2445
rect 12488 2343 12522 2377
rect 12692 2343 12726 2377
rect 12488 2275 12522 2309
rect 12692 2275 12726 2309
rect 12488 2207 12522 2241
rect 12692 2207 12726 2241
rect 12488 2139 12522 2173
rect 12692 2139 12726 2173
rect 12488 2071 12522 2105
rect 12692 2071 12726 2105
rect 12488 2003 12522 2037
rect 12692 2003 12726 2037
rect 12488 1935 12522 1969
rect 12692 1935 12726 1969
rect 12488 1867 12522 1901
rect 12692 1867 12726 1901
rect 12488 1799 12522 1833
rect 12692 1799 12726 1833
rect 12488 1731 12522 1765
rect 12692 1731 12726 1765
rect 12488 1663 12522 1697
rect 12692 1663 12726 1697
rect 12488 1595 12522 1629
rect 12692 1595 12726 1629
rect 12488 1527 12522 1561
rect 12692 1527 12726 1561
rect 13050 2411 13084 2445
rect 13122 2411 13156 2445
rect 13050 2343 13084 2377
rect 13122 2343 13156 2377
rect 13050 2275 13084 2309
rect 13122 2275 13156 2309
rect 13050 2207 13084 2241
rect 13122 2207 13156 2241
rect 13050 2139 13084 2173
rect 13122 2139 13156 2173
rect 13050 2071 13084 2105
rect 13122 2071 13156 2105
rect 13050 2003 13084 2037
rect 13122 2003 13156 2037
rect 13050 1935 13084 1969
rect 13122 1935 13156 1969
rect 13050 1867 13084 1901
rect 13122 1867 13156 1901
rect 13050 1799 13084 1833
rect 13122 1799 13156 1833
rect 13050 1731 13084 1765
rect 13122 1731 13156 1765
rect 13050 1663 13084 1697
rect 13122 1663 13156 1697
rect 13050 1595 13084 1629
rect 13122 1595 13156 1629
rect 13050 1527 13084 1561
rect 13122 1527 13156 1561
rect 13480 2411 13514 2445
rect 13684 2411 13718 2445
rect 13480 2343 13514 2377
rect 13684 2343 13718 2377
rect 13480 2275 13514 2309
rect 13684 2275 13718 2309
rect 13480 2207 13514 2241
rect 13684 2207 13718 2241
rect 13480 2139 13514 2173
rect 13684 2139 13718 2173
rect 13480 2071 13514 2105
rect 13684 2071 13718 2105
rect 13480 2003 13514 2037
rect 13684 2003 13718 2037
rect 13480 1935 13514 1969
rect 13684 1935 13718 1969
rect 13480 1867 13514 1901
rect 13684 1867 13718 1901
rect 13480 1799 13514 1833
rect 13684 1799 13718 1833
rect 13480 1731 13514 1765
rect 13684 1731 13718 1765
rect 13480 1663 13514 1697
rect 13684 1663 13718 1697
rect 13480 1595 13514 1629
rect 13684 1595 13718 1629
rect 13480 1527 13514 1561
rect 13684 1527 13718 1561
rect 14042 2411 14076 2445
rect 14042 2343 14076 2377
rect 14042 2275 14076 2309
rect 14042 2207 14076 2241
rect 14042 2139 14076 2173
rect 14042 2071 14076 2105
rect 14042 2003 14076 2037
rect 14042 1935 14076 1969
rect 14042 1867 14076 1901
rect 14042 1799 14076 1833
rect 14042 1731 14076 1765
rect 14042 1663 14076 1697
rect 14042 1595 14076 1629
rect 14042 1527 14076 1561
rect 14386 2411 14420 2445
rect 14386 2343 14420 2377
rect 14386 2275 14420 2309
rect 14386 2207 14420 2241
rect 14386 2139 14420 2173
rect 14386 2071 14420 2105
rect 14386 2003 14420 2037
rect 14386 1935 14420 1969
rect 14386 1867 14420 1901
rect 14386 1799 14420 1833
rect 14386 1731 14420 1765
rect 14386 1663 14420 1697
rect 14386 1595 14420 1629
rect 14386 1527 14420 1561
<< mvpsubdiff >>
rect 555 4922 657 4956
rect 14495 4922 14530 4956
rect 14564 4922 14599 4956
rect 14633 4922 14667 4956
rect 589 4888 657 4922
rect 14461 4888 14667 4922
rect 555 4854 623 4888
rect 14461 4854 14496 4888
rect 14530 4854 14565 4888
rect 14599 4854 14667 4888
rect 555 4850 691 4854
rect 589 4819 691 4850
rect 589 4816 623 4819
rect 555 4785 623 4816
rect 657 4786 691 4819
rect 14393 4844 14667 4854
rect 14393 4820 14633 4844
rect 14393 4786 14428 4820
rect 14462 4786 14497 4820
rect 14531 4818 14633 4820
rect 14531 4786 14565 4818
rect 657 4785 725 4786
rect 555 4778 725 4785
rect 589 4751 725 4778
rect 589 4750 691 4751
rect 589 4744 623 4750
rect 555 4716 623 4744
rect 657 4717 691 4750
rect 657 4716 725 4717
rect 555 4706 725 4716
rect 589 4682 725 4706
rect 589 4681 691 4682
rect 589 4672 623 4681
rect 555 4647 623 4672
rect 657 4648 691 4681
rect 657 4647 725 4648
rect 555 4634 725 4647
rect 589 4613 725 4634
rect 589 4600 623 4613
rect 555 4563 623 4600
rect 589 4529 623 4563
rect 555 4492 623 4529
rect 589 4458 623 4492
rect 555 4421 623 4458
rect 589 4387 623 4421
rect 555 4350 623 4387
rect 589 4316 623 4350
rect 555 4279 623 4316
rect 589 4245 623 4279
rect 555 4208 623 4245
rect 589 4174 623 4208
rect 555 4137 623 4174
rect 589 4103 623 4137
rect 14497 4784 14565 4786
rect 14599 4810 14633 4818
rect 14599 4784 14667 4810
rect 14497 4771 14667 4784
rect 14497 4750 14633 4771
rect 14531 4748 14633 4750
rect 14531 4716 14565 4748
rect 14497 4714 14565 4716
rect 14599 4737 14633 4748
rect 14599 4714 14667 4737
rect 14497 4698 14667 4714
rect 14497 4680 14633 4698
rect 14531 4678 14633 4680
rect 14531 4646 14565 4678
rect 14497 4644 14565 4646
rect 14599 4664 14633 4678
rect 14599 4644 14667 4664
rect 14497 4625 14667 4644
rect 14497 4610 14633 4625
rect 14531 4608 14633 4610
rect 14531 4576 14565 4608
rect 14497 4574 14565 4576
rect 14599 4591 14633 4608
rect 14599 4574 14667 4591
rect 14497 4552 14667 4574
rect 14497 4540 14633 4552
rect 14531 4538 14633 4540
rect 14531 4506 14565 4538
rect 14497 4504 14565 4506
rect 14599 4518 14633 4538
rect 14599 4504 14667 4518
rect 14497 4479 14667 4504
rect 14497 4470 14633 4479
rect 14531 4468 14633 4470
rect 14531 4436 14565 4468
rect 14497 4434 14565 4436
rect 14599 4445 14633 4468
rect 14599 4434 14667 4445
rect 14497 4406 14667 4434
rect 14497 4399 14633 4406
rect 14531 4398 14633 4399
rect 14531 4365 14565 4398
rect 14497 4364 14565 4365
rect 14599 4372 14633 4398
rect 14599 4364 14667 4372
rect 14497 4333 14667 4364
rect 14497 4328 14633 4333
rect 14531 4294 14565 4328
rect 14599 4299 14633 4328
rect 14599 4294 14667 4299
rect 14497 4260 14667 4294
rect 14497 4257 14633 4260
rect 555 4058 725 4103
rect 14531 4223 14565 4257
rect 14599 4226 14633 4257
rect 14599 4223 14667 4226
rect 14497 4186 14667 4223
rect 14531 4152 14565 4186
rect 14599 4152 14633 4186
rect 14497 4115 14667 4152
rect 14497 4081 14565 4115
rect 14599 4081 14633 4115
rect 14497 4058 14667 4081
rect 555 4041 787 4058
rect 589 4007 623 4041
rect 657 4034 787 4041
rect 657 4007 734 4034
rect 555 4000 734 4007
rect 768 4000 787 4034
rect 555 3970 787 4000
rect 589 3936 623 3970
rect 657 3966 787 3970
rect 657 3936 734 3966
rect 555 3932 734 3936
rect 768 3932 787 3966
rect 555 3898 787 3932
rect 555 3896 734 3898
rect 589 3862 623 3896
rect 657 3864 734 3896
rect 768 3864 787 3898
rect 657 3862 787 3864
rect 555 3830 787 3862
rect 555 3825 734 3830
rect 589 3791 623 3825
rect 657 3796 734 3825
rect 768 3796 787 3830
rect 657 3791 787 3796
rect 555 3762 787 3791
rect 555 3751 734 3762
rect 589 3717 623 3751
rect 657 3728 734 3751
rect 768 3728 787 3762
rect 657 3717 787 3728
rect 555 3694 787 3717
rect 555 3680 734 3694
rect 589 3646 623 3680
rect 657 3660 734 3680
rect 768 3660 787 3694
rect 657 3646 787 3660
rect 555 3626 787 3646
rect 555 3606 734 3626
rect 589 3572 623 3606
rect 657 3592 734 3606
rect 768 3592 787 3626
rect 657 3572 787 3592
rect 555 3558 787 3572
rect 555 3535 734 3558
rect 589 3501 623 3535
rect 657 3524 734 3535
rect 768 3524 787 3558
rect 657 3501 787 3524
rect 555 3490 787 3501
rect 555 3461 734 3490
rect 589 3427 623 3461
rect 657 3456 734 3461
rect 768 3456 787 3490
rect 657 3427 787 3456
rect 555 3422 787 3427
rect 555 3390 734 3422
rect 589 3356 623 3390
rect 657 3388 734 3390
rect 768 3388 787 3422
rect 657 3356 787 3388
rect 555 3354 787 3356
rect 555 3320 734 3354
rect 768 3320 787 3354
rect 555 3316 787 3320
rect 589 3282 623 3316
rect 657 3286 787 3316
rect 657 3282 734 3286
rect 555 3252 734 3282
rect 768 3252 787 3286
rect 555 3245 787 3252
rect 589 3211 623 3245
rect 657 3218 787 3245
rect 657 3211 734 3218
rect 555 3184 734 3211
rect 768 3184 787 3218
rect 555 3151 787 3184
rect 589 3117 623 3151
rect 657 3150 787 3151
rect 657 3117 734 3150
rect 555 3116 734 3117
rect 768 3116 787 3150
rect 555 3081 787 3116
rect 657 3058 787 3081
rect 1625 4046 1765 4058
rect 1625 4012 1678 4046
rect 1712 4012 1765 4046
rect 1625 3978 1765 4012
rect 1625 3944 1678 3978
rect 1712 3944 1765 3978
rect 1625 3910 1765 3944
rect 1625 3876 1678 3910
rect 1712 3876 1765 3910
rect 1625 3842 1765 3876
rect 1625 3808 1678 3842
rect 1712 3808 1765 3842
rect 1625 3774 1765 3808
rect 1625 3740 1678 3774
rect 1712 3740 1765 3774
rect 1625 3706 1765 3740
rect 1625 3672 1678 3706
rect 1712 3672 1765 3706
rect 1625 3638 1765 3672
rect 1625 3604 1678 3638
rect 1712 3604 1765 3638
rect 1625 3570 1765 3604
rect 1625 3536 1678 3570
rect 1712 3536 1765 3570
rect 1625 3502 1765 3536
rect 1625 3468 1678 3502
rect 1712 3468 1765 3502
rect 1625 3434 1765 3468
rect 1625 3400 1678 3434
rect 1712 3400 1765 3434
rect 1625 3366 1765 3400
rect 1625 3332 1678 3366
rect 1712 3332 1765 3366
rect 1625 3298 1765 3332
rect 1625 3264 1678 3298
rect 1712 3264 1765 3298
rect 1625 3230 1765 3264
rect 1625 3196 1678 3230
rect 1712 3196 1765 3230
rect 1625 3162 1765 3196
rect 1625 3128 1678 3162
rect 1712 3128 1765 3162
rect 1625 3058 1765 3128
rect 2617 4046 2757 4058
rect 2617 4012 2670 4046
rect 2704 4012 2757 4046
rect 2617 3978 2757 4012
rect 2617 3944 2670 3978
rect 2704 3944 2757 3978
rect 2617 3910 2757 3944
rect 2617 3876 2670 3910
rect 2704 3876 2757 3910
rect 2617 3842 2757 3876
rect 2617 3808 2670 3842
rect 2704 3808 2757 3842
rect 2617 3774 2757 3808
rect 2617 3740 2670 3774
rect 2704 3740 2757 3774
rect 2617 3706 2757 3740
rect 2617 3672 2670 3706
rect 2704 3672 2757 3706
rect 2617 3638 2757 3672
rect 2617 3604 2670 3638
rect 2704 3604 2757 3638
rect 2617 3570 2757 3604
rect 2617 3536 2670 3570
rect 2704 3536 2757 3570
rect 2617 3502 2757 3536
rect 2617 3468 2670 3502
rect 2704 3468 2757 3502
rect 2617 3434 2757 3468
rect 2617 3400 2670 3434
rect 2704 3400 2757 3434
rect 2617 3366 2757 3400
rect 2617 3332 2670 3366
rect 2704 3332 2757 3366
rect 2617 3298 2757 3332
rect 2617 3264 2670 3298
rect 2704 3264 2757 3298
rect 2617 3230 2757 3264
rect 2617 3196 2670 3230
rect 2704 3196 2757 3230
rect 2617 3162 2757 3196
rect 2617 3128 2670 3162
rect 2704 3128 2757 3162
rect 2617 3058 2757 3128
rect 3609 4046 3749 4058
rect 3609 4012 3662 4046
rect 3696 4012 3749 4046
rect 3609 3978 3749 4012
rect 3609 3944 3662 3978
rect 3696 3944 3749 3978
rect 3609 3910 3749 3944
rect 3609 3876 3662 3910
rect 3696 3876 3749 3910
rect 3609 3842 3749 3876
rect 3609 3808 3662 3842
rect 3696 3808 3749 3842
rect 3609 3774 3749 3808
rect 3609 3740 3662 3774
rect 3696 3740 3749 3774
rect 3609 3706 3749 3740
rect 3609 3672 3662 3706
rect 3696 3672 3749 3706
rect 3609 3638 3749 3672
rect 3609 3604 3662 3638
rect 3696 3604 3749 3638
rect 3609 3570 3749 3604
rect 3609 3536 3662 3570
rect 3696 3536 3749 3570
rect 3609 3502 3749 3536
rect 3609 3468 3662 3502
rect 3696 3468 3749 3502
rect 3609 3434 3749 3468
rect 3609 3400 3662 3434
rect 3696 3400 3749 3434
rect 3609 3366 3749 3400
rect 3609 3332 3662 3366
rect 3696 3332 3749 3366
rect 3609 3298 3749 3332
rect 3609 3264 3662 3298
rect 3696 3264 3749 3298
rect 3609 3230 3749 3264
rect 3609 3196 3662 3230
rect 3696 3196 3749 3230
rect 3609 3162 3749 3196
rect 3609 3128 3662 3162
rect 3696 3128 3749 3162
rect 3609 3058 3749 3128
rect 4601 4046 4741 4058
rect 4601 4012 4654 4046
rect 4688 4012 4741 4046
rect 4601 3978 4741 4012
rect 4601 3944 4654 3978
rect 4688 3944 4741 3978
rect 4601 3910 4741 3944
rect 4601 3876 4654 3910
rect 4688 3876 4741 3910
rect 4601 3842 4741 3876
rect 4601 3808 4654 3842
rect 4688 3808 4741 3842
rect 4601 3774 4741 3808
rect 4601 3740 4654 3774
rect 4688 3740 4741 3774
rect 4601 3706 4741 3740
rect 4601 3672 4654 3706
rect 4688 3672 4741 3706
rect 4601 3638 4741 3672
rect 4601 3604 4654 3638
rect 4688 3604 4741 3638
rect 4601 3570 4741 3604
rect 4601 3536 4654 3570
rect 4688 3536 4741 3570
rect 4601 3502 4741 3536
rect 4601 3468 4654 3502
rect 4688 3468 4741 3502
rect 4601 3434 4741 3468
rect 4601 3400 4654 3434
rect 4688 3400 4741 3434
rect 4601 3366 4741 3400
rect 4601 3332 4654 3366
rect 4688 3332 4741 3366
rect 4601 3298 4741 3332
rect 4601 3264 4654 3298
rect 4688 3264 4741 3298
rect 4601 3230 4741 3264
rect 4601 3196 4654 3230
rect 4688 3196 4741 3230
rect 4601 3162 4741 3196
rect 4601 3128 4654 3162
rect 4688 3128 4741 3162
rect 4601 3058 4741 3128
rect 5593 4046 5733 4058
rect 5593 4012 5646 4046
rect 5680 4012 5733 4046
rect 5593 3978 5733 4012
rect 5593 3944 5646 3978
rect 5680 3944 5733 3978
rect 5593 3910 5733 3944
rect 5593 3876 5646 3910
rect 5680 3876 5733 3910
rect 5593 3842 5733 3876
rect 5593 3808 5646 3842
rect 5680 3808 5733 3842
rect 5593 3774 5733 3808
rect 5593 3740 5646 3774
rect 5680 3740 5733 3774
rect 5593 3706 5733 3740
rect 5593 3672 5646 3706
rect 5680 3672 5733 3706
rect 5593 3638 5733 3672
rect 5593 3604 5646 3638
rect 5680 3604 5733 3638
rect 5593 3570 5733 3604
rect 5593 3536 5646 3570
rect 5680 3536 5733 3570
rect 5593 3502 5733 3536
rect 5593 3468 5646 3502
rect 5680 3468 5733 3502
rect 5593 3434 5733 3468
rect 5593 3400 5646 3434
rect 5680 3400 5733 3434
rect 5593 3366 5733 3400
rect 5593 3332 5646 3366
rect 5680 3332 5733 3366
rect 5593 3298 5733 3332
rect 5593 3264 5646 3298
rect 5680 3264 5733 3298
rect 5593 3230 5733 3264
rect 5593 3196 5646 3230
rect 5680 3196 5733 3230
rect 5593 3162 5733 3196
rect 5593 3128 5646 3162
rect 5680 3128 5733 3162
rect 5593 3058 5733 3128
rect 6585 4046 6725 4058
rect 6585 4012 6638 4046
rect 6672 4012 6725 4046
rect 6585 3978 6725 4012
rect 6585 3944 6638 3978
rect 6672 3944 6725 3978
rect 6585 3910 6725 3944
rect 6585 3876 6638 3910
rect 6672 3876 6725 3910
rect 6585 3842 6725 3876
rect 6585 3808 6638 3842
rect 6672 3808 6725 3842
rect 6585 3774 6725 3808
rect 6585 3740 6638 3774
rect 6672 3740 6725 3774
rect 6585 3706 6725 3740
rect 6585 3672 6638 3706
rect 6672 3672 6725 3706
rect 6585 3638 6725 3672
rect 6585 3604 6638 3638
rect 6672 3604 6725 3638
rect 6585 3570 6725 3604
rect 6585 3536 6638 3570
rect 6672 3536 6725 3570
rect 6585 3502 6725 3536
rect 6585 3468 6638 3502
rect 6672 3468 6725 3502
rect 6585 3434 6725 3468
rect 6585 3400 6638 3434
rect 6672 3400 6725 3434
rect 6585 3366 6725 3400
rect 6585 3332 6638 3366
rect 6672 3332 6725 3366
rect 6585 3298 6725 3332
rect 6585 3264 6638 3298
rect 6672 3264 6725 3298
rect 6585 3230 6725 3264
rect 6585 3196 6638 3230
rect 6672 3196 6725 3230
rect 6585 3162 6725 3196
rect 6585 3128 6638 3162
rect 6672 3128 6725 3162
rect 6585 3058 6725 3128
rect 7577 4046 7717 4058
rect 7577 4012 7630 4046
rect 7664 4012 7717 4046
rect 7577 3978 7717 4012
rect 7577 3944 7630 3978
rect 7664 3944 7717 3978
rect 7577 3910 7717 3944
rect 7577 3876 7630 3910
rect 7664 3876 7717 3910
rect 7577 3842 7717 3876
rect 7577 3808 7630 3842
rect 7664 3808 7717 3842
rect 7577 3774 7717 3808
rect 7577 3740 7630 3774
rect 7664 3740 7717 3774
rect 7577 3706 7717 3740
rect 7577 3672 7630 3706
rect 7664 3672 7717 3706
rect 7577 3638 7717 3672
rect 7577 3604 7630 3638
rect 7664 3604 7717 3638
rect 7577 3570 7717 3604
rect 7577 3536 7630 3570
rect 7664 3536 7717 3570
rect 7577 3502 7717 3536
rect 7577 3468 7630 3502
rect 7664 3468 7717 3502
rect 7577 3434 7717 3468
rect 7577 3400 7630 3434
rect 7664 3400 7717 3434
rect 7577 3366 7717 3400
rect 7577 3332 7630 3366
rect 7664 3332 7717 3366
rect 7577 3298 7717 3332
rect 7577 3264 7630 3298
rect 7664 3264 7717 3298
rect 7577 3230 7717 3264
rect 7577 3196 7630 3230
rect 7664 3196 7717 3230
rect 7577 3162 7717 3196
rect 7577 3128 7630 3162
rect 7664 3128 7717 3162
rect 7577 3058 7717 3128
rect 8569 4046 8709 4058
rect 8569 4012 8622 4046
rect 8656 4012 8709 4046
rect 8569 3978 8709 4012
rect 8569 3944 8622 3978
rect 8656 3944 8709 3978
rect 8569 3910 8709 3944
rect 8569 3876 8622 3910
rect 8656 3876 8709 3910
rect 8569 3842 8709 3876
rect 8569 3808 8622 3842
rect 8656 3808 8709 3842
rect 8569 3774 8709 3808
rect 8569 3740 8622 3774
rect 8656 3740 8709 3774
rect 8569 3706 8709 3740
rect 8569 3672 8622 3706
rect 8656 3672 8709 3706
rect 8569 3638 8709 3672
rect 8569 3604 8622 3638
rect 8656 3604 8709 3638
rect 8569 3570 8709 3604
rect 8569 3536 8622 3570
rect 8656 3536 8709 3570
rect 8569 3502 8709 3536
rect 8569 3468 8622 3502
rect 8656 3468 8709 3502
rect 8569 3434 8709 3468
rect 8569 3400 8622 3434
rect 8656 3400 8709 3434
rect 8569 3366 8709 3400
rect 8569 3332 8622 3366
rect 8656 3332 8709 3366
rect 8569 3298 8709 3332
rect 8569 3264 8622 3298
rect 8656 3264 8709 3298
rect 8569 3230 8709 3264
rect 8569 3196 8622 3230
rect 8656 3196 8709 3230
rect 8569 3162 8709 3196
rect 8569 3128 8622 3162
rect 8656 3128 8709 3162
rect 8569 3058 8709 3128
rect 9561 4046 9701 4058
rect 9561 4012 9614 4046
rect 9648 4012 9701 4046
rect 9561 3978 9701 4012
rect 9561 3944 9614 3978
rect 9648 3944 9701 3978
rect 9561 3910 9701 3944
rect 9561 3876 9614 3910
rect 9648 3876 9701 3910
rect 9561 3842 9701 3876
rect 9561 3808 9614 3842
rect 9648 3808 9701 3842
rect 9561 3774 9701 3808
rect 9561 3740 9614 3774
rect 9648 3740 9701 3774
rect 9561 3706 9701 3740
rect 9561 3672 9614 3706
rect 9648 3672 9701 3706
rect 9561 3638 9701 3672
rect 9561 3604 9614 3638
rect 9648 3604 9701 3638
rect 9561 3570 9701 3604
rect 9561 3536 9614 3570
rect 9648 3536 9701 3570
rect 9561 3502 9701 3536
rect 9561 3468 9614 3502
rect 9648 3468 9701 3502
rect 9561 3434 9701 3468
rect 9561 3400 9614 3434
rect 9648 3400 9701 3434
rect 9561 3366 9701 3400
rect 9561 3332 9614 3366
rect 9648 3332 9701 3366
rect 9561 3298 9701 3332
rect 9561 3264 9614 3298
rect 9648 3264 9701 3298
rect 9561 3230 9701 3264
rect 9561 3196 9614 3230
rect 9648 3196 9701 3230
rect 9561 3162 9701 3196
rect 9561 3128 9614 3162
rect 9648 3128 9701 3162
rect 9561 3058 9701 3128
rect 10553 4046 10693 4058
rect 10553 4012 10606 4046
rect 10640 4012 10693 4046
rect 10553 3978 10693 4012
rect 10553 3944 10606 3978
rect 10640 3944 10693 3978
rect 10553 3910 10693 3944
rect 10553 3876 10606 3910
rect 10640 3876 10693 3910
rect 10553 3842 10693 3876
rect 10553 3808 10606 3842
rect 10640 3808 10693 3842
rect 10553 3774 10693 3808
rect 10553 3740 10606 3774
rect 10640 3740 10693 3774
rect 10553 3706 10693 3740
rect 10553 3672 10606 3706
rect 10640 3672 10693 3706
rect 10553 3638 10693 3672
rect 10553 3604 10606 3638
rect 10640 3604 10693 3638
rect 10553 3570 10693 3604
rect 10553 3536 10606 3570
rect 10640 3536 10693 3570
rect 10553 3502 10693 3536
rect 10553 3468 10606 3502
rect 10640 3468 10693 3502
rect 10553 3434 10693 3468
rect 10553 3400 10606 3434
rect 10640 3400 10693 3434
rect 10553 3366 10693 3400
rect 10553 3332 10606 3366
rect 10640 3332 10693 3366
rect 10553 3298 10693 3332
rect 10553 3264 10606 3298
rect 10640 3264 10693 3298
rect 10553 3230 10693 3264
rect 10553 3196 10606 3230
rect 10640 3196 10693 3230
rect 10553 3162 10693 3196
rect 10553 3128 10606 3162
rect 10640 3128 10693 3162
rect 10553 3058 10693 3128
rect 11545 4046 11685 4058
rect 11545 4012 11598 4046
rect 11632 4012 11685 4046
rect 11545 3978 11685 4012
rect 11545 3944 11598 3978
rect 11632 3944 11685 3978
rect 11545 3910 11685 3944
rect 11545 3876 11598 3910
rect 11632 3876 11685 3910
rect 11545 3842 11685 3876
rect 11545 3808 11598 3842
rect 11632 3808 11685 3842
rect 11545 3774 11685 3808
rect 11545 3740 11598 3774
rect 11632 3740 11685 3774
rect 11545 3706 11685 3740
rect 11545 3672 11598 3706
rect 11632 3672 11685 3706
rect 11545 3638 11685 3672
rect 11545 3604 11598 3638
rect 11632 3604 11685 3638
rect 11545 3570 11685 3604
rect 11545 3536 11598 3570
rect 11632 3536 11685 3570
rect 11545 3502 11685 3536
rect 11545 3468 11598 3502
rect 11632 3468 11685 3502
rect 11545 3434 11685 3468
rect 11545 3400 11598 3434
rect 11632 3400 11685 3434
rect 11545 3366 11685 3400
rect 11545 3332 11598 3366
rect 11632 3332 11685 3366
rect 11545 3298 11685 3332
rect 11545 3264 11598 3298
rect 11632 3264 11685 3298
rect 11545 3230 11685 3264
rect 11545 3196 11598 3230
rect 11632 3196 11685 3230
rect 11545 3162 11685 3196
rect 11545 3128 11598 3162
rect 11632 3128 11685 3162
rect 11545 3058 11685 3128
rect 12537 4046 12677 4058
rect 12537 4012 12590 4046
rect 12624 4012 12677 4046
rect 12537 3978 12677 4012
rect 12537 3944 12590 3978
rect 12624 3944 12677 3978
rect 12537 3910 12677 3944
rect 12537 3876 12590 3910
rect 12624 3876 12677 3910
rect 12537 3842 12677 3876
rect 12537 3808 12590 3842
rect 12624 3808 12677 3842
rect 12537 3774 12677 3808
rect 12537 3740 12590 3774
rect 12624 3740 12677 3774
rect 12537 3706 12677 3740
rect 12537 3672 12590 3706
rect 12624 3672 12677 3706
rect 12537 3638 12677 3672
rect 12537 3604 12590 3638
rect 12624 3604 12677 3638
rect 12537 3570 12677 3604
rect 12537 3536 12590 3570
rect 12624 3536 12677 3570
rect 12537 3502 12677 3536
rect 12537 3468 12590 3502
rect 12624 3468 12677 3502
rect 12537 3434 12677 3468
rect 12537 3400 12590 3434
rect 12624 3400 12677 3434
rect 12537 3366 12677 3400
rect 12537 3332 12590 3366
rect 12624 3332 12677 3366
rect 12537 3298 12677 3332
rect 12537 3264 12590 3298
rect 12624 3264 12677 3298
rect 12537 3230 12677 3264
rect 12537 3196 12590 3230
rect 12624 3196 12677 3230
rect 12537 3162 12677 3196
rect 12537 3128 12590 3162
rect 12624 3128 12677 3162
rect 12537 3058 12677 3128
rect 13529 4046 13669 4058
rect 13529 4012 13582 4046
rect 13616 4012 13669 4046
rect 13529 3978 13669 4012
rect 13529 3944 13582 3978
rect 13616 3944 13669 3978
rect 13529 3910 13669 3944
rect 13529 3876 13582 3910
rect 13616 3876 13669 3910
rect 13529 3842 13669 3876
rect 13529 3808 13582 3842
rect 13616 3808 13669 3842
rect 13529 3774 13669 3808
rect 13529 3740 13582 3774
rect 13616 3740 13669 3774
rect 13529 3706 13669 3740
rect 13529 3672 13582 3706
rect 13616 3672 13669 3706
rect 13529 3638 13669 3672
rect 13529 3604 13582 3638
rect 13616 3604 13669 3638
rect 13529 3570 13669 3604
rect 13529 3536 13582 3570
rect 13616 3536 13669 3570
rect 13529 3502 13669 3536
rect 13529 3468 13582 3502
rect 13616 3468 13669 3502
rect 13529 3434 13669 3468
rect 13529 3400 13582 3434
rect 13616 3400 13669 3434
rect 13529 3366 13669 3400
rect 13529 3332 13582 3366
rect 13616 3332 13669 3366
rect 13529 3298 13669 3332
rect 13529 3264 13582 3298
rect 13616 3264 13669 3298
rect 13529 3230 13669 3264
rect 13529 3196 13582 3230
rect 13616 3196 13669 3230
rect 13529 3162 13669 3196
rect 13529 3128 13582 3162
rect 13616 3128 13669 3162
rect 13529 3058 13669 3128
rect 14435 4041 14667 4058
rect 14435 4034 14565 4041
rect 14435 4000 14454 4034
rect 14488 4007 14565 4034
rect 14599 4007 14633 4041
rect 14488 4000 14667 4007
rect 14435 3970 14667 4000
rect 14435 3966 14565 3970
rect 14435 3932 14454 3966
rect 14488 3936 14565 3966
rect 14599 3936 14633 3970
rect 14488 3932 14667 3936
rect 14435 3898 14667 3932
rect 14435 3864 14454 3898
rect 14488 3896 14667 3898
rect 14488 3864 14565 3896
rect 14435 3862 14565 3864
rect 14599 3862 14633 3896
rect 14435 3830 14667 3862
rect 14435 3796 14454 3830
rect 14488 3825 14667 3830
rect 14488 3796 14565 3825
rect 14435 3791 14565 3796
rect 14599 3791 14633 3825
rect 14435 3762 14667 3791
rect 14435 3728 14454 3762
rect 14488 3751 14667 3762
rect 14488 3728 14565 3751
rect 14435 3717 14565 3728
rect 14599 3717 14633 3751
rect 14435 3694 14667 3717
rect 14435 3660 14454 3694
rect 14488 3680 14667 3694
rect 14488 3660 14565 3680
rect 14435 3646 14565 3660
rect 14599 3646 14633 3680
rect 14435 3626 14667 3646
rect 14435 3592 14454 3626
rect 14488 3606 14667 3626
rect 14488 3592 14565 3606
rect 14435 3572 14565 3592
rect 14599 3572 14633 3606
rect 14435 3558 14667 3572
rect 14435 3524 14454 3558
rect 14488 3535 14667 3558
rect 14488 3524 14565 3535
rect 14435 3501 14565 3524
rect 14599 3501 14633 3535
rect 14435 3490 14667 3501
rect 14435 3456 14454 3490
rect 14488 3461 14667 3490
rect 14488 3456 14565 3461
rect 14435 3427 14565 3456
rect 14599 3427 14633 3461
rect 14435 3422 14667 3427
rect 14435 3388 14454 3422
rect 14488 3390 14667 3422
rect 14488 3388 14565 3390
rect 14435 3356 14565 3388
rect 14599 3356 14633 3390
rect 14435 3354 14667 3356
rect 14435 3320 14454 3354
rect 14488 3320 14667 3354
rect 14435 3316 14667 3320
rect 14435 3286 14565 3316
rect 14435 3252 14454 3286
rect 14488 3282 14565 3286
rect 14599 3282 14633 3316
rect 14488 3252 14667 3282
rect 14435 3245 14667 3252
rect 14435 3218 14565 3245
rect 14435 3184 14454 3218
rect 14488 3211 14565 3218
rect 14599 3211 14633 3245
rect 14488 3184 14667 3211
rect 14435 3151 14667 3184
rect 14435 3150 14565 3151
rect 14435 3116 14454 3150
rect 14488 3117 14565 3150
rect 14599 3117 14633 3151
rect 14488 3116 14667 3117
rect 14435 3066 14667 3116
rect 14435 3058 14565 3066
rect 657 3013 725 3058
rect 657 2457 725 2503
rect 1578 2935 1814 2969
rect 1578 2901 1645 2935
rect 1679 2901 1713 2935
rect 1747 2901 1814 2935
rect 1578 2855 1814 2901
rect 1578 2821 1645 2855
rect 1679 2821 1713 2855
rect 1747 2821 1814 2855
rect 1578 2775 1814 2821
rect 1578 2741 1645 2775
rect 1679 2741 1713 2775
rect 1747 2741 1814 2775
rect 1578 2695 1814 2741
rect 1578 2661 1645 2695
rect 1679 2661 1713 2695
rect 1747 2661 1814 2695
rect 1578 2614 1814 2661
rect 1578 2580 1645 2614
rect 1679 2580 1713 2614
rect 1747 2580 1814 2614
rect 1578 2546 1814 2580
rect 2570 2935 2806 2969
rect 2570 2901 2637 2935
rect 2671 2901 2705 2935
rect 2739 2901 2806 2935
rect 2570 2855 2806 2901
rect 2570 2821 2637 2855
rect 2671 2821 2705 2855
rect 2739 2821 2806 2855
rect 2570 2775 2806 2821
rect 2570 2741 2637 2775
rect 2671 2741 2705 2775
rect 2739 2741 2806 2775
rect 2570 2695 2806 2741
rect 2570 2661 2637 2695
rect 2671 2661 2705 2695
rect 2739 2661 2806 2695
rect 2570 2614 2806 2661
rect 2570 2580 2637 2614
rect 2671 2580 2705 2614
rect 2739 2580 2806 2614
rect 2570 2546 2806 2580
rect 3562 2935 3798 2969
rect 3562 2901 3629 2935
rect 3663 2901 3697 2935
rect 3731 2901 3798 2935
rect 3562 2855 3798 2901
rect 3562 2821 3629 2855
rect 3663 2821 3697 2855
rect 3731 2821 3798 2855
rect 3562 2775 3798 2821
rect 3562 2741 3629 2775
rect 3663 2741 3697 2775
rect 3731 2741 3798 2775
rect 3562 2695 3798 2741
rect 3562 2661 3629 2695
rect 3663 2661 3697 2695
rect 3731 2661 3798 2695
rect 3562 2614 3798 2661
rect 3562 2580 3629 2614
rect 3663 2580 3697 2614
rect 3731 2580 3798 2614
rect 3562 2546 3798 2580
rect 4554 2935 4790 2969
rect 4554 2901 4621 2935
rect 4655 2901 4689 2935
rect 4723 2901 4790 2935
rect 4554 2855 4790 2901
rect 4554 2821 4621 2855
rect 4655 2821 4689 2855
rect 4723 2821 4790 2855
rect 4554 2775 4790 2821
rect 4554 2741 4621 2775
rect 4655 2741 4689 2775
rect 4723 2741 4790 2775
rect 4554 2695 4790 2741
rect 4554 2661 4621 2695
rect 4655 2661 4689 2695
rect 4723 2661 4790 2695
rect 4554 2614 4790 2661
rect 4554 2580 4621 2614
rect 4655 2580 4689 2614
rect 4723 2580 4790 2614
rect 4554 2546 4790 2580
rect 5546 2935 5782 2969
rect 5546 2901 5613 2935
rect 5647 2901 5681 2935
rect 5715 2901 5782 2935
rect 5546 2855 5782 2901
rect 5546 2821 5613 2855
rect 5647 2821 5681 2855
rect 5715 2821 5782 2855
rect 5546 2775 5782 2821
rect 5546 2741 5613 2775
rect 5647 2741 5681 2775
rect 5715 2741 5782 2775
rect 5546 2695 5782 2741
rect 5546 2661 5613 2695
rect 5647 2661 5681 2695
rect 5715 2661 5782 2695
rect 5546 2614 5782 2661
rect 5546 2580 5613 2614
rect 5647 2580 5681 2614
rect 5715 2580 5782 2614
rect 5546 2546 5782 2580
rect 6538 2935 6774 2969
rect 6538 2901 6605 2935
rect 6639 2901 6673 2935
rect 6707 2901 6774 2935
rect 6538 2855 6774 2901
rect 6538 2821 6605 2855
rect 6639 2821 6673 2855
rect 6707 2821 6774 2855
rect 6538 2775 6774 2821
rect 6538 2741 6605 2775
rect 6639 2741 6673 2775
rect 6707 2741 6774 2775
rect 6538 2695 6774 2741
rect 6538 2661 6605 2695
rect 6639 2661 6673 2695
rect 6707 2661 6774 2695
rect 6538 2614 6774 2661
rect 6538 2580 6605 2614
rect 6639 2580 6673 2614
rect 6707 2580 6774 2614
rect 6538 2546 6774 2580
rect 7530 2935 7766 2969
rect 7530 2901 7597 2935
rect 7631 2901 7665 2935
rect 7699 2901 7766 2935
rect 7530 2855 7766 2901
rect 7530 2821 7597 2855
rect 7631 2821 7665 2855
rect 7699 2821 7766 2855
rect 7530 2775 7766 2821
rect 7530 2741 7597 2775
rect 7631 2741 7665 2775
rect 7699 2741 7766 2775
rect 7530 2695 7766 2741
rect 7530 2661 7597 2695
rect 7631 2661 7665 2695
rect 7699 2661 7766 2695
rect 7530 2614 7766 2661
rect 7530 2580 7597 2614
rect 7631 2580 7665 2614
rect 7699 2580 7766 2614
rect 7530 2546 7766 2580
rect 8522 2935 8758 2969
rect 8522 2901 8589 2935
rect 8623 2901 8657 2935
rect 8691 2901 8758 2935
rect 8522 2855 8758 2901
rect 8522 2821 8589 2855
rect 8623 2821 8657 2855
rect 8691 2821 8758 2855
rect 8522 2775 8758 2821
rect 8522 2741 8589 2775
rect 8623 2741 8657 2775
rect 8691 2741 8758 2775
rect 8522 2695 8758 2741
rect 8522 2661 8589 2695
rect 8623 2661 8657 2695
rect 8691 2661 8758 2695
rect 8522 2614 8758 2661
rect 8522 2580 8589 2614
rect 8623 2580 8657 2614
rect 8691 2580 8758 2614
rect 8522 2546 8758 2580
rect 9514 2935 9750 2969
rect 9514 2901 9581 2935
rect 9615 2901 9649 2935
rect 9683 2901 9750 2935
rect 9514 2855 9750 2901
rect 9514 2821 9581 2855
rect 9615 2821 9649 2855
rect 9683 2821 9750 2855
rect 9514 2775 9750 2821
rect 9514 2741 9581 2775
rect 9615 2741 9649 2775
rect 9683 2741 9750 2775
rect 9514 2695 9750 2741
rect 9514 2661 9581 2695
rect 9615 2661 9649 2695
rect 9683 2661 9750 2695
rect 9514 2614 9750 2661
rect 9514 2580 9581 2614
rect 9615 2580 9649 2614
rect 9683 2580 9750 2614
rect 9514 2546 9750 2580
rect 10506 2935 10742 2969
rect 10506 2901 10573 2935
rect 10607 2901 10641 2935
rect 10675 2901 10742 2935
rect 10506 2855 10742 2901
rect 10506 2821 10573 2855
rect 10607 2821 10641 2855
rect 10675 2821 10742 2855
rect 10506 2775 10742 2821
rect 10506 2741 10573 2775
rect 10607 2741 10641 2775
rect 10675 2741 10742 2775
rect 10506 2695 10742 2741
rect 10506 2661 10573 2695
rect 10607 2661 10641 2695
rect 10675 2661 10742 2695
rect 10506 2614 10742 2661
rect 10506 2580 10573 2614
rect 10607 2580 10641 2614
rect 10675 2580 10742 2614
rect 10506 2546 10742 2580
rect 11498 2935 11734 2969
rect 11498 2901 11565 2935
rect 11599 2901 11633 2935
rect 11667 2901 11734 2935
rect 11498 2855 11734 2901
rect 11498 2821 11565 2855
rect 11599 2821 11633 2855
rect 11667 2821 11734 2855
rect 11498 2775 11734 2821
rect 11498 2741 11565 2775
rect 11599 2741 11633 2775
rect 11667 2741 11734 2775
rect 11498 2695 11734 2741
rect 11498 2661 11565 2695
rect 11599 2661 11633 2695
rect 11667 2661 11734 2695
rect 11498 2614 11734 2661
rect 11498 2580 11565 2614
rect 11599 2580 11633 2614
rect 11667 2580 11734 2614
rect 11498 2546 11734 2580
rect 12490 2935 12726 2969
rect 12490 2901 12557 2935
rect 12591 2901 12625 2935
rect 12659 2901 12726 2935
rect 12490 2855 12726 2901
rect 12490 2821 12557 2855
rect 12591 2821 12625 2855
rect 12659 2821 12726 2855
rect 12490 2775 12726 2821
rect 12490 2741 12557 2775
rect 12591 2741 12625 2775
rect 12659 2741 12726 2775
rect 12490 2695 12726 2741
rect 12490 2661 12557 2695
rect 12591 2661 12625 2695
rect 12659 2661 12726 2695
rect 12490 2614 12726 2661
rect 12490 2580 12557 2614
rect 12591 2580 12625 2614
rect 12659 2580 12726 2614
rect 12490 2546 12726 2580
rect 13482 2935 13718 2969
rect 13482 2901 13549 2935
rect 13583 2901 13617 2935
rect 13651 2901 13718 2935
rect 13482 2855 13718 2901
rect 13482 2821 13549 2855
rect 13583 2821 13617 2855
rect 13651 2821 13718 2855
rect 13482 2775 13718 2821
rect 13482 2741 13549 2775
rect 13583 2741 13617 2775
rect 13651 2741 13718 2775
rect 13482 2695 13718 2741
rect 13482 2661 13549 2695
rect 13583 2661 13617 2695
rect 13651 2661 13718 2695
rect 13482 2614 13718 2661
rect 13482 2580 13549 2614
rect 13583 2580 13617 2614
rect 13651 2580 13718 2614
rect 13482 2546 13718 2580
rect 14497 3032 14565 3058
rect 14599 3032 14633 3066
rect 14497 2972 14667 3032
rect 14497 2485 14667 2530
rect 14497 2457 14565 2485
rect 657 2433 787 2457
rect 657 2399 734 2433
rect 768 2399 787 2433
rect 657 2367 787 2399
rect 555 2365 787 2367
rect 555 2331 734 2365
rect 768 2331 787 2365
rect 555 2327 787 2331
rect 589 2293 623 2327
rect 657 2297 787 2327
rect 657 2293 734 2297
rect 555 2263 734 2293
rect 768 2263 787 2297
rect 555 2250 787 2263
rect 589 2216 623 2250
rect 657 2229 787 2250
rect 657 2216 734 2229
rect 555 2195 734 2216
rect 768 2195 787 2229
rect 555 2161 787 2195
rect 555 2156 734 2161
rect 589 2122 623 2156
rect 657 2127 734 2156
rect 768 2127 787 2161
rect 657 2122 787 2127
rect 555 2093 787 2122
rect 555 2085 734 2093
rect 589 2051 623 2085
rect 657 2059 734 2085
rect 768 2059 787 2093
rect 657 2051 787 2059
rect 555 2025 787 2051
rect 555 2011 734 2025
rect 589 1977 623 2011
rect 657 1991 734 2011
rect 768 1991 787 2025
rect 657 1977 787 1991
rect 555 1957 787 1977
rect 555 1940 734 1957
rect 589 1906 623 1940
rect 657 1923 734 1940
rect 768 1923 787 1957
rect 657 1906 787 1923
rect 555 1889 787 1906
rect 555 1866 734 1889
rect 589 1832 623 1866
rect 657 1855 734 1866
rect 768 1855 787 1889
rect 657 1832 787 1855
rect 555 1821 787 1832
rect 555 1795 734 1821
rect 589 1761 623 1795
rect 657 1787 734 1795
rect 768 1787 787 1821
rect 657 1761 787 1787
rect 555 1753 787 1761
rect 555 1721 734 1753
rect 589 1687 623 1721
rect 657 1719 734 1721
rect 768 1719 787 1753
rect 657 1687 787 1719
rect 555 1685 787 1687
rect 555 1651 734 1685
rect 768 1651 787 1685
rect 555 1650 787 1651
rect 589 1616 623 1650
rect 657 1617 787 1650
rect 657 1616 734 1617
rect 555 1583 734 1616
rect 768 1583 787 1617
rect 555 1576 787 1583
rect 589 1542 623 1576
rect 657 1549 787 1576
rect 657 1542 734 1549
rect 555 1515 734 1542
rect 768 1515 787 1549
rect 555 1505 787 1515
rect 589 1471 623 1505
rect 657 1471 787 1505
rect 555 1457 787 1471
rect 1625 2445 1765 2457
rect 1625 2411 1678 2445
rect 1712 2411 1765 2445
rect 1625 2377 1765 2411
rect 1625 2343 1678 2377
rect 1712 2343 1765 2377
rect 1625 2309 1765 2343
rect 1625 2275 1678 2309
rect 1712 2275 1765 2309
rect 1625 2241 1765 2275
rect 1625 2207 1678 2241
rect 1712 2207 1765 2241
rect 1625 2173 1765 2207
rect 1625 2139 1678 2173
rect 1712 2139 1765 2173
rect 1625 2105 1765 2139
rect 1625 2071 1678 2105
rect 1712 2071 1765 2105
rect 1625 2037 1765 2071
rect 1625 2003 1678 2037
rect 1712 2003 1765 2037
rect 1625 1969 1765 2003
rect 1625 1935 1678 1969
rect 1712 1935 1765 1969
rect 1625 1901 1765 1935
rect 1625 1867 1678 1901
rect 1712 1867 1765 1901
rect 1625 1833 1765 1867
rect 1625 1799 1678 1833
rect 1712 1799 1765 1833
rect 1625 1765 1765 1799
rect 1625 1731 1678 1765
rect 1712 1731 1765 1765
rect 1625 1697 1765 1731
rect 1625 1663 1678 1697
rect 1712 1663 1765 1697
rect 1625 1629 1765 1663
rect 1625 1595 1678 1629
rect 1712 1595 1765 1629
rect 1625 1561 1765 1595
rect 1625 1527 1678 1561
rect 1712 1527 1765 1561
rect 1625 1457 1765 1527
rect 2617 2445 2757 2457
rect 2617 2411 2670 2445
rect 2704 2411 2757 2445
rect 2617 2377 2757 2411
rect 2617 2343 2670 2377
rect 2704 2343 2757 2377
rect 2617 2309 2757 2343
rect 2617 2275 2670 2309
rect 2704 2275 2757 2309
rect 2617 2241 2757 2275
rect 2617 2207 2670 2241
rect 2704 2207 2757 2241
rect 2617 2173 2757 2207
rect 2617 2139 2670 2173
rect 2704 2139 2757 2173
rect 2617 2105 2757 2139
rect 2617 2071 2670 2105
rect 2704 2071 2757 2105
rect 2617 2037 2757 2071
rect 2617 2003 2670 2037
rect 2704 2003 2757 2037
rect 2617 1969 2757 2003
rect 2617 1935 2670 1969
rect 2704 1935 2757 1969
rect 2617 1901 2757 1935
rect 2617 1867 2670 1901
rect 2704 1867 2757 1901
rect 2617 1833 2757 1867
rect 2617 1799 2670 1833
rect 2704 1799 2757 1833
rect 2617 1765 2757 1799
rect 2617 1731 2670 1765
rect 2704 1731 2757 1765
rect 2617 1697 2757 1731
rect 2617 1663 2670 1697
rect 2704 1663 2757 1697
rect 2617 1629 2757 1663
rect 2617 1595 2670 1629
rect 2704 1595 2757 1629
rect 2617 1561 2757 1595
rect 2617 1527 2670 1561
rect 2704 1527 2757 1561
rect 2617 1457 2757 1527
rect 3609 2445 3749 2457
rect 3609 2411 3662 2445
rect 3696 2411 3749 2445
rect 3609 2377 3749 2411
rect 3609 2343 3662 2377
rect 3696 2343 3749 2377
rect 3609 2309 3749 2343
rect 3609 2275 3662 2309
rect 3696 2275 3749 2309
rect 3609 2241 3749 2275
rect 3609 2207 3662 2241
rect 3696 2207 3749 2241
rect 3609 2173 3749 2207
rect 3609 2139 3662 2173
rect 3696 2139 3749 2173
rect 3609 2105 3749 2139
rect 3609 2071 3662 2105
rect 3696 2071 3749 2105
rect 3609 2037 3749 2071
rect 3609 2003 3662 2037
rect 3696 2003 3749 2037
rect 3609 1969 3749 2003
rect 3609 1935 3662 1969
rect 3696 1935 3749 1969
rect 3609 1901 3749 1935
rect 3609 1867 3662 1901
rect 3696 1867 3749 1901
rect 3609 1833 3749 1867
rect 3609 1799 3662 1833
rect 3696 1799 3749 1833
rect 3609 1765 3749 1799
rect 3609 1731 3662 1765
rect 3696 1731 3749 1765
rect 3609 1697 3749 1731
rect 3609 1663 3662 1697
rect 3696 1663 3749 1697
rect 3609 1629 3749 1663
rect 3609 1595 3662 1629
rect 3696 1595 3749 1629
rect 3609 1561 3749 1595
rect 3609 1527 3662 1561
rect 3696 1527 3749 1561
rect 3609 1457 3749 1527
rect 4601 2445 4741 2457
rect 4601 2411 4654 2445
rect 4688 2411 4741 2445
rect 4601 2377 4741 2411
rect 4601 2343 4654 2377
rect 4688 2343 4741 2377
rect 4601 2309 4741 2343
rect 4601 2275 4654 2309
rect 4688 2275 4741 2309
rect 4601 2241 4741 2275
rect 4601 2207 4654 2241
rect 4688 2207 4741 2241
rect 4601 2173 4741 2207
rect 4601 2139 4654 2173
rect 4688 2139 4741 2173
rect 4601 2105 4741 2139
rect 4601 2071 4654 2105
rect 4688 2071 4741 2105
rect 4601 2037 4741 2071
rect 4601 2003 4654 2037
rect 4688 2003 4741 2037
rect 4601 1969 4741 2003
rect 4601 1935 4654 1969
rect 4688 1935 4741 1969
rect 4601 1901 4741 1935
rect 4601 1867 4654 1901
rect 4688 1867 4741 1901
rect 4601 1833 4741 1867
rect 4601 1799 4654 1833
rect 4688 1799 4741 1833
rect 4601 1765 4741 1799
rect 4601 1731 4654 1765
rect 4688 1731 4741 1765
rect 4601 1697 4741 1731
rect 4601 1663 4654 1697
rect 4688 1663 4741 1697
rect 4601 1629 4741 1663
rect 4601 1595 4654 1629
rect 4688 1595 4741 1629
rect 4601 1561 4741 1595
rect 4601 1527 4654 1561
rect 4688 1527 4741 1561
rect 4601 1457 4741 1527
rect 5593 2445 5733 2457
rect 5593 2411 5646 2445
rect 5680 2411 5733 2445
rect 5593 2377 5733 2411
rect 5593 2343 5646 2377
rect 5680 2343 5733 2377
rect 5593 2309 5733 2343
rect 5593 2275 5646 2309
rect 5680 2275 5733 2309
rect 5593 2241 5733 2275
rect 5593 2207 5646 2241
rect 5680 2207 5733 2241
rect 5593 2173 5733 2207
rect 5593 2139 5646 2173
rect 5680 2139 5733 2173
rect 5593 2105 5733 2139
rect 5593 2071 5646 2105
rect 5680 2071 5733 2105
rect 5593 2037 5733 2071
rect 5593 2003 5646 2037
rect 5680 2003 5733 2037
rect 5593 1969 5733 2003
rect 5593 1935 5646 1969
rect 5680 1935 5733 1969
rect 5593 1901 5733 1935
rect 5593 1867 5646 1901
rect 5680 1867 5733 1901
rect 5593 1833 5733 1867
rect 5593 1799 5646 1833
rect 5680 1799 5733 1833
rect 5593 1765 5733 1799
rect 5593 1731 5646 1765
rect 5680 1731 5733 1765
rect 5593 1697 5733 1731
rect 5593 1663 5646 1697
rect 5680 1663 5733 1697
rect 5593 1629 5733 1663
rect 5593 1595 5646 1629
rect 5680 1595 5733 1629
rect 5593 1561 5733 1595
rect 5593 1527 5646 1561
rect 5680 1527 5733 1561
rect 5593 1457 5733 1527
rect 6585 2445 6725 2457
rect 6585 2411 6638 2445
rect 6672 2411 6725 2445
rect 6585 2377 6725 2411
rect 6585 2343 6638 2377
rect 6672 2343 6725 2377
rect 6585 2309 6725 2343
rect 6585 2275 6638 2309
rect 6672 2275 6725 2309
rect 6585 2241 6725 2275
rect 6585 2207 6638 2241
rect 6672 2207 6725 2241
rect 6585 2173 6725 2207
rect 6585 2139 6638 2173
rect 6672 2139 6725 2173
rect 6585 2105 6725 2139
rect 6585 2071 6638 2105
rect 6672 2071 6725 2105
rect 6585 2037 6725 2071
rect 6585 2003 6638 2037
rect 6672 2003 6725 2037
rect 6585 1969 6725 2003
rect 6585 1935 6638 1969
rect 6672 1935 6725 1969
rect 6585 1901 6725 1935
rect 6585 1867 6638 1901
rect 6672 1867 6725 1901
rect 6585 1833 6725 1867
rect 6585 1799 6638 1833
rect 6672 1799 6725 1833
rect 6585 1765 6725 1799
rect 6585 1731 6638 1765
rect 6672 1731 6725 1765
rect 6585 1697 6725 1731
rect 6585 1663 6638 1697
rect 6672 1663 6725 1697
rect 6585 1629 6725 1663
rect 6585 1595 6638 1629
rect 6672 1595 6725 1629
rect 6585 1561 6725 1595
rect 6585 1527 6638 1561
rect 6672 1527 6725 1561
rect 6585 1457 6725 1527
rect 7577 2445 7717 2457
rect 7577 2411 7630 2445
rect 7664 2411 7717 2445
rect 7577 2377 7717 2411
rect 7577 2343 7630 2377
rect 7664 2343 7717 2377
rect 7577 2309 7717 2343
rect 7577 2275 7630 2309
rect 7664 2275 7717 2309
rect 7577 2241 7717 2275
rect 7577 2207 7630 2241
rect 7664 2207 7717 2241
rect 7577 2173 7717 2207
rect 7577 2139 7630 2173
rect 7664 2139 7717 2173
rect 7577 2105 7717 2139
rect 7577 2071 7630 2105
rect 7664 2071 7717 2105
rect 7577 2037 7717 2071
rect 7577 2003 7630 2037
rect 7664 2003 7717 2037
rect 7577 1969 7717 2003
rect 7577 1935 7630 1969
rect 7664 1935 7717 1969
rect 7577 1901 7717 1935
rect 7577 1867 7630 1901
rect 7664 1867 7717 1901
rect 7577 1833 7717 1867
rect 7577 1799 7630 1833
rect 7664 1799 7717 1833
rect 7577 1765 7717 1799
rect 7577 1731 7630 1765
rect 7664 1731 7717 1765
rect 7577 1697 7717 1731
rect 7577 1663 7630 1697
rect 7664 1663 7717 1697
rect 7577 1629 7717 1663
rect 7577 1595 7630 1629
rect 7664 1595 7717 1629
rect 7577 1561 7717 1595
rect 7577 1527 7630 1561
rect 7664 1527 7717 1561
rect 7577 1457 7717 1527
rect 8569 2445 8709 2457
rect 8569 2411 8622 2445
rect 8656 2411 8709 2445
rect 8569 2377 8709 2411
rect 8569 2343 8622 2377
rect 8656 2343 8709 2377
rect 8569 2309 8709 2343
rect 8569 2275 8622 2309
rect 8656 2275 8709 2309
rect 8569 2241 8709 2275
rect 8569 2207 8622 2241
rect 8656 2207 8709 2241
rect 8569 2173 8709 2207
rect 8569 2139 8622 2173
rect 8656 2139 8709 2173
rect 8569 2105 8709 2139
rect 8569 2071 8622 2105
rect 8656 2071 8709 2105
rect 8569 2037 8709 2071
rect 8569 2003 8622 2037
rect 8656 2003 8709 2037
rect 8569 1969 8709 2003
rect 8569 1935 8622 1969
rect 8656 1935 8709 1969
rect 8569 1901 8709 1935
rect 8569 1867 8622 1901
rect 8656 1867 8709 1901
rect 8569 1833 8709 1867
rect 8569 1799 8622 1833
rect 8656 1799 8709 1833
rect 8569 1765 8709 1799
rect 8569 1731 8622 1765
rect 8656 1731 8709 1765
rect 8569 1697 8709 1731
rect 8569 1663 8622 1697
rect 8656 1663 8709 1697
rect 8569 1629 8709 1663
rect 8569 1595 8622 1629
rect 8656 1595 8709 1629
rect 8569 1561 8709 1595
rect 8569 1527 8622 1561
rect 8656 1527 8709 1561
rect 8569 1457 8709 1527
rect 9561 2445 9701 2457
rect 9561 2411 9614 2445
rect 9648 2411 9701 2445
rect 9561 2377 9701 2411
rect 9561 2343 9614 2377
rect 9648 2343 9701 2377
rect 9561 2309 9701 2343
rect 9561 2275 9614 2309
rect 9648 2275 9701 2309
rect 9561 2241 9701 2275
rect 9561 2207 9614 2241
rect 9648 2207 9701 2241
rect 9561 2173 9701 2207
rect 9561 2139 9614 2173
rect 9648 2139 9701 2173
rect 9561 2105 9701 2139
rect 9561 2071 9614 2105
rect 9648 2071 9701 2105
rect 9561 2037 9701 2071
rect 9561 2003 9614 2037
rect 9648 2003 9701 2037
rect 9561 1969 9701 2003
rect 9561 1935 9614 1969
rect 9648 1935 9701 1969
rect 9561 1901 9701 1935
rect 9561 1867 9614 1901
rect 9648 1867 9701 1901
rect 9561 1833 9701 1867
rect 9561 1799 9614 1833
rect 9648 1799 9701 1833
rect 9561 1765 9701 1799
rect 9561 1731 9614 1765
rect 9648 1731 9701 1765
rect 9561 1697 9701 1731
rect 9561 1663 9614 1697
rect 9648 1663 9701 1697
rect 9561 1629 9701 1663
rect 9561 1595 9614 1629
rect 9648 1595 9701 1629
rect 9561 1561 9701 1595
rect 9561 1527 9614 1561
rect 9648 1527 9701 1561
rect 9561 1457 9701 1527
rect 10553 2445 10693 2457
rect 10553 2411 10606 2445
rect 10640 2411 10693 2445
rect 10553 2377 10693 2411
rect 10553 2343 10606 2377
rect 10640 2343 10693 2377
rect 10553 2309 10693 2343
rect 10553 2275 10606 2309
rect 10640 2275 10693 2309
rect 10553 2241 10693 2275
rect 10553 2207 10606 2241
rect 10640 2207 10693 2241
rect 10553 2173 10693 2207
rect 10553 2139 10606 2173
rect 10640 2139 10693 2173
rect 10553 2105 10693 2139
rect 10553 2071 10606 2105
rect 10640 2071 10693 2105
rect 10553 2037 10693 2071
rect 10553 2003 10606 2037
rect 10640 2003 10693 2037
rect 10553 1969 10693 2003
rect 10553 1935 10606 1969
rect 10640 1935 10693 1969
rect 10553 1901 10693 1935
rect 10553 1867 10606 1901
rect 10640 1867 10693 1901
rect 10553 1833 10693 1867
rect 10553 1799 10606 1833
rect 10640 1799 10693 1833
rect 10553 1765 10693 1799
rect 10553 1731 10606 1765
rect 10640 1731 10693 1765
rect 10553 1697 10693 1731
rect 10553 1663 10606 1697
rect 10640 1663 10693 1697
rect 10553 1629 10693 1663
rect 10553 1595 10606 1629
rect 10640 1595 10693 1629
rect 10553 1561 10693 1595
rect 10553 1527 10606 1561
rect 10640 1527 10693 1561
rect 10553 1457 10693 1527
rect 11545 2445 11685 2457
rect 11545 2411 11598 2445
rect 11632 2411 11685 2445
rect 11545 2377 11685 2411
rect 11545 2343 11598 2377
rect 11632 2343 11685 2377
rect 11545 2309 11685 2343
rect 11545 2275 11598 2309
rect 11632 2275 11685 2309
rect 11545 2241 11685 2275
rect 11545 2207 11598 2241
rect 11632 2207 11685 2241
rect 11545 2173 11685 2207
rect 11545 2139 11598 2173
rect 11632 2139 11685 2173
rect 11545 2105 11685 2139
rect 11545 2071 11598 2105
rect 11632 2071 11685 2105
rect 11545 2037 11685 2071
rect 11545 2003 11598 2037
rect 11632 2003 11685 2037
rect 11545 1969 11685 2003
rect 11545 1935 11598 1969
rect 11632 1935 11685 1969
rect 11545 1901 11685 1935
rect 11545 1867 11598 1901
rect 11632 1867 11685 1901
rect 11545 1833 11685 1867
rect 11545 1799 11598 1833
rect 11632 1799 11685 1833
rect 11545 1765 11685 1799
rect 11545 1731 11598 1765
rect 11632 1731 11685 1765
rect 11545 1697 11685 1731
rect 11545 1663 11598 1697
rect 11632 1663 11685 1697
rect 11545 1629 11685 1663
rect 11545 1595 11598 1629
rect 11632 1595 11685 1629
rect 11545 1561 11685 1595
rect 11545 1527 11598 1561
rect 11632 1527 11685 1561
rect 11545 1457 11685 1527
rect 12537 2445 12677 2457
rect 12537 2411 12590 2445
rect 12624 2411 12677 2445
rect 12537 2377 12677 2411
rect 12537 2343 12590 2377
rect 12624 2343 12677 2377
rect 12537 2309 12677 2343
rect 12537 2275 12590 2309
rect 12624 2275 12677 2309
rect 12537 2241 12677 2275
rect 12537 2207 12590 2241
rect 12624 2207 12677 2241
rect 12537 2173 12677 2207
rect 12537 2139 12590 2173
rect 12624 2139 12677 2173
rect 12537 2105 12677 2139
rect 12537 2071 12590 2105
rect 12624 2071 12677 2105
rect 12537 2037 12677 2071
rect 12537 2003 12590 2037
rect 12624 2003 12677 2037
rect 12537 1969 12677 2003
rect 12537 1935 12590 1969
rect 12624 1935 12677 1969
rect 12537 1901 12677 1935
rect 12537 1867 12590 1901
rect 12624 1867 12677 1901
rect 12537 1833 12677 1867
rect 12537 1799 12590 1833
rect 12624 1799 12677 1833
rect 12537 1765 12677 1799
rect 12537 1731 12590 1765
rect 12624 1731 12677 1765
rect 12537 1697 12677 1731
rect 12537 1663 12590 1697
rect 12624 1663 12677 1697
rect 12537 1629 12677 1663
rect 12537 1595 12590 1629
rect 12624 1595 12677 1629
rect 12537 1561 12677 1595
rect 12537 1527 12590 1561
rect 12624 1527 12677 1561
rect 12537 1457 12677 1527
rect 13529 2445 13669 2457
rect 13529 2411 13582 2445
rect 13616 2411 13669 2445
rect 13529 2377 13669 2411
rect 13529 2343 13582 2377
rect 13616 2343 13669 2377
rect 13529 2309 13669 2343
rect 13529 2275 13582 2309
rect 13616 2275 13669 2309
rect 13529 2241 13669 2275
rect 13529 2207 13582 2241
rect 13616 2207 13669 2241
rect 13529 2173 13669 2207
rect 13529 2139 13582 2173
rect 13616 2139 13669 2173
rect 13529 2105 13669 2139
rect 13529 2071 13582 2105
rect 13616 2071 13669 2105
rect 13529 2037 13669 2071
rect 13529 2003 13582 2037
rect 13616 2003 13669 2037
rect 13529 1969 13669 2003
rect 13529 1935 13582 1969
rect 13616 1935 13669 1969
rect 13529 1901 13669 1935
rect 13529 1867 13582 1901
rect 13616 1867 13669 1901
rect 13529 1833 13669 1867
rect 13529 1799 13582 1833
rect 13616 1799 13669 1833
rect 13529 1765 13669 1799
rect 13529 1731 13582 1765
rect 13616 1731 13669 1765
rect 13529 1697 13669 1731
rect 13529 1663 13582 1697
rect 13616 1663 13669 1697
rect 13529 1629 13669 1663
rect 13529 1595 13582 1629
rect 13616 1595 13669 1629
rect 13529 1561 13669 1595
rect 13529 1527 13582 1561
rect 13616 1527 13669 1561
rect 13529 1457 13669 1527
rect 14435 2451 14565 2457
rect 14599 2451 14633 2485
rect 14435 2433 14667 2451
rect 14435 2399 14454 2433
rect 14488 2403 14667 2433
rect 14488 2399 14565 2403
rect 14435 2369 14565 2399
rect 14599 2369 14633 2403
rect 14435 2365 14667 2369
rect 14435 2331 14454 2365
rect 14488 2331 14667 2365
rect 14435 2327 14667 2331
rect 14435 2297 14565 2327
rect 14435 2263 14454 2297
rect 14488 2293 14565 2297
rect 14599 2293 14633 2327
rect 14488 2263 14667 2293
rect 14435 2250 14667 2263
rect 14435 2229 14565 2250
rect 14435 2195 14454 2229
rect 14488 2216 14565 2229
rect 14599 2216 14633 2250
rect 14488 2195 14667 2216
rect 14435 2161 14667 2195
rect 14435 2127 14454 2161
rect 14488 2156 14667 2161
rect 14488 2127 14565 2156
rect 14435 2122 14565 2127
rect 14599 2122 14633 2156
rect 14435 2093 14667 2122
rect 14435 2059 14454 2093
rect 14488 2085 14667 2093
rect 14488 2059 14565 2085
rect 14435 2051 14565 2059
rect 14599 2051 14633 2085
rect 14435 2025 14667 2051
rect 14435 1991 14454 2025
rect 14488 2011 14667 2025
rect 14488 1991 14565 2011
rect 14435 1977 14565 1991
rect 14599 1977 14633 2011
rect 14435 1957 14667 1977
rect 14435 1923 14454 1957
rect 14488 1940 14667 1957
rect 14488 1923 14565 1940
rect 14435 1906 14565 1923
rect 14599 1906 14633 1940
rect 14435 1889 14667 1906
rect 14435 1855 14454 1889
rect 14488 1866 14667 1889
rect 14488 1855 14565 1866
rect 14435 1832 14565 1855
rect 14599 1832 14633 1866
rect 14435 1821 14667 1832
rect 14435 1787 14454 1821
rect 14488 1795 14667 1821
rect 14488 1787 14565 1795
rect 14435 1761 14565 1787
rect 14599 1761 14633 1795
rect 14435 1753 14667 1761
rect 14435 1719 14454 1753
rect 14488 1721 14667 1753
rect 14488 1719 14565 1721
rect 14435 1687 14565 1719
rect 14599 1687 14633 1721
rect 14435 1685 14667 1687
rect 14435 1651 14454 1685
rect 14488 1651 14667 1685
rect 14435 1650 14667 1651
rect 14435 1617 14565 1650
rect 14435 1583 14454 1617
rect 14488 1616 14565 1617
rect 14599 1616 14633 1650
rect 14488 1583 14667 1616
rect 14435 1576 14667 1583
rect 14435 1549 14565 1576
rect 14435 1515 14454 1549
rect 14488 1542 14565 1549
rect 14599 1542 14633 1576
rect 14488 1515 14667 1542
rect 14435 1505 14667 1515
rect 14435 1471 14565 1505
rect 14599 1471 14633 1505
rect 14435 1457 14667 1471
rect 555 1375 725 1457
rect 589 1341 623 1375
rect 657 1341 691 1375
rect 555 1221 725 1341
rect 14497 1387 14667 1457
rect 14531 1353 14565 1387
rect 14599 1353 14633 1387
rect 14497 1319 14667 1353
rect 14497 1311 14633 1319
rect 14497 1308 14565 1311
rect 589 1187 623 1221
rect 657 1219 725 1221
rect 657 1187 691 1219
rect 555 1185 691 1187
rect 555 1150 725 1185
rect 555 1140 623 1150
rect 589 1116 623 1140
rect 657 1148 725 1150
rect 14531 1277 14565 1308
rect 14599 1285 14633 1311
rect 14599 1277 14667 1285
rect 14531 1274 14667 1277
rect 14497 1251 14667 1274
rect 14497 1234 14633 1251
rect 14497 1228 14565 1234
rect 14531 1200 14565 1228
rect 14599 1217 14633 1234
rect 14599 1200 14667 1217
rect 14531 1194 14667 1200
rect 14497 1183 14667 1194
rect 14497 1157 14633 1183
rect 14497 1148 14565 1157
rect 657 1116 691 1148
rect 589 1114 691 1116
rect 725 1114 760 1148
rect 794 1114 829 1148
rect 589 1106 829 1114
rect 555 1080 829 1106
rect 14531 1123 14565 1148
rect 14599 1149 14633 1157
rect 14599 1123 14667 1149
rect 14531 1115 14667 1123
rect 14531 1081 14633 1115
rect 14531 1080 14667 1081
rect 555 1046 623 1080
rect 657 1046 692 1080
rect 726 1046 761 1080
rect 14599 1046 14667 1080
rect 555 1012 761 1046
rect 14565 1012 14633 1046
rect 555 978 589 1012
rect 623 978 658 1012
rect 692 978 727 1012
rect 14565 978 14667 1012
<< mvnsubdiff >>
rect 67 5422 15106 5426
rect 67 5303 294 5422
rect 67 5269 71 5303
rect 105 5269 139 5303
rect 173 5269 207 5303
rect 241 5269 294 5303
rect 67 5252 294 5269
rect 10868 5388 10903 5422
rect 10937 5388 10972 5422
rect 11006 5388 11041 5422
rect 11075 5388 11110 5422
rect 11144 5388 11179 5422
rect 11213 5388 11248 5422
rect 11282 5388 11317 5422
rect 11351 5388 11386 5422
rect 11420 5388 11455 5422
rect 11489 5388 11524 5422
rect 11558 5388 11593 5422
rect 11627 5388 11662 5422
rect 11696 5388 11731 5422
rect 11765 5388 11800 5422
rect 11834 5388 11869 5422
rect 11903 5388 11938 5422
rect 11972 5388 12007 5422
rect 12041 5388 12076 5422
rect 12110 5388 12145 5422
rect 12179 5388 12214 5422
rect 12248 5388 12283 5422
rect 12317 5388 12352 5422
rect 12386 5388 12421 5422
rect 12455 5388 12490 5422
rect 12524 5388 12559 5422
rect 12593 5388 12628 5422
rect 12662 5388 12697 5422
rect 12731 5388 12766 5422
rect 12800 5388 12835 5422
rect 12869 5388 12904 5422
rect 12938 5388 12973 5422
rect 13007 5388 13042 5422
rect 13076 5388 13111 5422
rect 13145 5388 13180 5422
rect 13214 5388 13249 5422
rect 13283 5388 13318 5422
rect 13352 5388 13387 5422
rect 13421 5388 13456 5422
rect 13490 5388 13525 5422
rect 13559 5388 13594 5422
rect 13628 5388 13663 5422
rect 13697 5388 13732 5422
rect 13766 5388 13801 5422
rect 13835 5388 13870 5422
rect 13904 5388 13939 5422
rect 13973 5388 14008 5422
rect 14042 5388 14077 5422
rect 14111 5388 14146 5422
rect 14180 5388 14215 5422
rect 14249 5388 14284 5422
rect 14318 5388 14353 5422
rect 14387 5388 14422 5422
rect 14456 5388 14491 5422
rect 14525 5388 14560 5422
rect 14594 5388 14629 5422
rect 14663 5388 14698 5422
rect 14732 5388 14767 5422
rect 14801 5388 14836 5422
rect 14870 5388 15106 5422
rect 10868 5354 15106 5388
rect 10868 5320 10903 5354
rect 10937 5320 10972 5354
rect 11006 5320 11041 5354
rect 11075 5320 11110 5354
rect 11144 5320 11179 5354
rect 11213 5320 11248 5354
rect 11282 5320 11317 5354
rect 11351 5320 11386 5354
rect 11420 5320 11455 5354
rect 11489 5320 11524 5354
rect 11558 5320 11593 5354
rect 11627 5320 11662 5354
rect 11696 5320 11731 5354
rect 11765 5320 11800 5354
rect 11834 5320 11869 5354
rect 11903 5320 11938 5354
rect 11972 5320 12007 5354
rect 12041 5320 12076 5354
rect 12110 5320 12145 5354
rect 12179 5320 12214 5354
rect 12248 5320 12283 5354
rect 12317 5320 12352 5354
rect 12386 5320 12421 5354
rect 12455 5320 12490 5354
rect 12524 5320 12559 5354
rect 12593 5320 12628 5354
rect 12662 5320 12697 5354
rect 12731 5320 12766 5354
rect 12800 5320 12835 5354
rect 12869 5320 12904 5354
rect 12938 5320 12973 5354
rect 13007 5320 13042 5354
rect 13076 5320 13111 5354
rect 13145 5320 13180 5354
rect 13214 5320 13249 5354
rect 13283 5320 13318 5354
rect 13352 5320 13387 5354
rect 13421 5320 13456 5354
rect 13490 5320 13525 5354
rect 13559 5320 13594 5354
rect 13628 5320 13663 5354
rect 13697 5320 13732 5354
rect 13766 5320 13801 5354
rect 13835 5320 13870 5354
rect 13904 5320 13939 5354
rect 13973 5320 14008 5354
rect 14042 5320 14077 5354
rect 14111 5320 14146 5354
rect 14180 5320 14215 5354
rect 14249 5320 14284 5354
rect 14318 5320 14353 5354
rect 14387 5320 14422 5354
rect 14456 5320 14491 5354
rect 14525 5320 14560 5354
rect 14594 5320 14629 5354
rect 14663 5320 14698 5354
rect 14732 5320 14767 5354
rect 14801 5320 14836 5354
rect 14870 5328 15106 5354
rect 14870 5320 14935 5328
rect 10868 5294 14935 5320
rect 14969 5294 15003 5328
rect 15037 5294 15071 5328
rect 15105 5294 15106 5328
rect 10868 5286 15106 5294
rect 10868 5252 10903 5286
rect 10937 5252 10972 5286
rect 11006 5252 11041 5286
rect 11075 5252 11110 5286
rect 11144 5252 11179 5286
rect 11213 5252 11248 5286
rect 11282 5252 11317 5286
rect 11351 5252 11386 5286
rect 11420 5252 11455 5286
rect 11489 5252 11524 5286
rect 11558 5252 11593 5286
rect 11627 5252 11662 5286
rect 11696 5252 11731 5286
rect 11765 5252 11800 5286
rect 11834 5252 11869 5286
rect 11903 5252 11938 5286
rect 11972 5252 12007 5286
rect 12041 5252 12076 5286
rect 12110 5252 12145 5286
rect 12179 5252 12214 5286
rect 12248 5252 12283 5286
rect 12317 5252 12352 5286
rect 12386 5252 12421 5286
rect 12455 5252 12490 5286
rect 12524 5252 12559 5286
rect 12593 5252 12628 5286
rect 12662 5252 12697 5286
rect 12731 5252 12766 5286
rect 12800 5252 12835 5286
rect 12869 5252 12904 5286
rect 12938 5252 12973 5286
rect 13007 5252 13042 5286
rect 13076 5252 13111 5286
rect 13145 5252 13180 5286
rect 13214 5252 13249 5286
rect 13283 5252 13318 5286
rect 13352 5252 13387 5286
rect 13421 5252 13456 5286
rect 13490 5252 13525 5286
rect 13559 5252 13594 5286
rect 13628 5252 13663 5286
rect 13697 5252 13732 5286
rect 13766 5252 13801 5286
rect 13835 5252 13870 5286
rect 13904 5252 13939 5286
rect 13973 5252 14008 5286
rect 14042 5252 14077 5286
rect 14111 5252 14146 5286
rect 14180 5252 14215 5286
rect 14249 5252 14284 5286
rect 14318 5252 14353 5286
rect 14387 5252 14422 5286
rect 14456 5252 14491 5286
rect 14525 5252 14560 5286
rect 14594 5252 14629 5286
rect 14663 5252 14698 5286
rect 14732 5252 14767 5286
rect 14801 5252 14836 5286
rect 14870 5256 15106 5286
rect 14870 5252 14935 5256
rect 67 5248 14935 5252
rect 67 5232 245 5248
rect 67 5198 71 5232
rect 105 5198 139 5232
rect 173 5198 207 5232
rect 241 5198 245 5232
rect 67 5161 245 5198
rect 67 5127 71 5161
rect 105 5127 139 5161
rect 173 5127 207 5161
rect 241 5127 245 5161
rect 67 5090 245 5127
rect 67 5056 71 5090
rect 105 5056 139 5090
rect 173 5056 207 5090
rect 241 5056 245 5090
rect 67 5020 245 5056
rect 67 4986 71 5020
rect 105 4986 139 5020
rect 173 4986 207 5020
rect 241 4986 245 5020
rect 67 4918 245 4986
rect 14928 5222 14935 5248
rect 14969 5222 15003 5256
rect 15037 5222 15071 5256
rect 15105 5222 15106 5256
rect 14928 5184 15106 5222
rect 14928 5150 14935 5184
rect 14969 5150 15003 5184
rect 15037 5150 15071 5184
rect 15105 5150 15106 5184
rect 14928 5112 15106 5150
rect 14928 5078 14935 5112
rect 14969 5078 15003 5112
rect 15037 5078 15071 5112
rect 15105 5078 15106 5112
rect 14928 5040 15106 5078
rect 14928 5006 14935 5040
rect 14969 5006 15003 5040
rect 15037 5006 15071 5040
rect 15105 5006 15106 5040
rect 14928 4968 15106 5006
rect 67 4884 71 4918
rect 105 4884 139 4918
rect 173 4884 207 4918
rect 241 4884 245 4918
rect 67 4849 245 4884
rect 67 4815 71 4849
rect 105 4815 139 4849
rect 173 4815 207 4849
rect 241 4815 245 4849
rect 67 4780 245 4815
rect 67 4746 71 4780
rect 105 4746 139 4780
rect 173 4746 207 4780
rect 241 4746 245 4780
rect 67 4711 245 4746
rect 67 4677 71 4711
rect 105 4677 139 4711
rect 173 4677 207 4711
rect 241 4677 245 4711
rect 67 4642 245 4677
rect 67 4608 71 4642
rect 105 4608 139 4642
rect 173 4608 207 4642
rect 241 4608 245 4642
rect 67 4573 245 4608
rect 67 4539 71 4573
rect 105 4539 139 4573
rect 173 4539 207 4573
rect 241 4539 245 4573
rect 67 4504 245 4539
rect 67 4470 71 4504
rect 105 4470 139 4504
rect 173 4470 207 4504
rect 241 4470 245 4504
rect 67 4435 245 4470
rect 67 4401 71 4435
rect 105 4401 139 4435
rect 173 4401 207 4435
rect 241 4401 245 4435
rect 67 4366 245 4401
rect 67 4332 71 4366
rect 105 4332 139 4366
rect 173 4332 207 4366
rect 241 4332 245 4366
rect 67 4297 245 4332
rect 67 4263 71 4297
rect 105 4263 139 4297
rect 173 4263 207 4297
rect 241 4263 245 4297
rect 67 4228 245 4263
rect 67 4194 71 4228
rect 105 4194 139 4228
rect 173 4194 207 4228
rect 241 4194 245 4228
rect 67 4159 245 4194
rect 67 4125 71 4159
rect 105 4125 139 4159
rect 173 4125 207 4159
rect 241 4125 245 4159
rect 67 4090 245 4125
rect 67 4056 71 4090
rect 105 4056 139 4090
rect 173 4056 207 4090
rect 241 4056 245 4090
rect 67 4021 245 4056
rect 67 3987 71 4021
rect 105 3987 139 4021
rect 173 3987 207 4021
rect 241 3987 245 4021
rect 67 3952 245 3987
rect 67 3918 71 3952
rect 105 3918 139 3952
rect 173 3918 207 3952
rect 241 3918 245 3952
rect 67 3883 245 3918
rect 67 3849 71 3883
rect 105 3849 139 3883
rect 173 3849 207 3883
rect 241 3849 245 3883
rect 67 3814 245 3849
rect 67 3780 71 3814
rect 105 3780 139 3814
rect 173 3780 207 3814
rect 241 3780 245 3814
rect 67 3745 245 3780
rect 67 3711 71 3745
rect 105 3711 139 3745
rect 173 3711 207 3745
rect 241 3711 245 3745
rect 67 3676 245 3711
rect 67 3642 71 3676
rect 105 3642 139 3676
rect 173 3642 207 3676
rect 241 3642 245 3676
rect 67 3607 245 3642
rect 67 3573 71 3607
rect 105 3573 139 3607
rect 173 3573 207 3607
rect 241 3573 245 3607
rect 67 3538 245 3573
rect 67 3504 71 3538
rect 105 3504 139 3538
rect 173 3504 207 3538
rect 241 3504 245 3538
rect 67 3469 245 3504
rect 67 3435 71 3469
rect 105 3435 139 3469
rect 173 3435 207 3469
rect 241 3435 245 3469
rect 67 3400 245 3435
rect 67 3366 71 3400
rect 105 3366 139 3400
rect 173 3366 207 3400
rect 241 3366 245 3400
rect 67 3331 245 3366
rect 67 3297 71 3331
rect 105 3297 139 3331
rect 173 3297 207 3331
rect 241 3297 245 3331
rect 67 3262 245 3297
rect 67 3228 71 3262
rect 105 3228 139 3262
rect 173 3228 207 3262
rect 241 3228 245 3262
rect 67 3193 245 3228
rect 67 3159 71 3193
rect 105 3159 139 3193
rect 173 3159 207 3193
rect 241 3159 245 3193
rect 67 3124 245 3159
rect 67 3090 71 3124
rect 105 3090 139 3124
rect 173 3090 207 3124
rect 241 3090 245 3124
rect 67 3055 245 3090
rect 67 3021 71 3055
rect 105 3021 139 3055
rect 173 3021 207 3055
rect 241 3021 245 3055
rect 67 2986 245 3021
rect 67 2952 71 2986
rect 105 2952 139 2986
rect 173 2952 207 2986
rect 241 2952 245 2986
rect 67 2917 245 2952
rect 67 2883 71 2917
rect 105 2883 139 2917
rect 173 2883 207 2917
rect 241 2883 245 2917
rect 67 2848 245 2883
rect 67 2814 71 2848
rect 105 2814 139 2848
rect 173 2814 207 2848
rect 241 2814 245 2848
rect 67 2779 245 2814
rect 67 2745 71 2779
rect 105 2745 139 2779
rect 173 2745 207 2779
rect 241 2745 245 2779
rect 67 2710 245 2745
rect 67 2676 71 2710
rect 105 2676 139 2710
rect 173 2676 207 2710
rect 241 2676 245 2710
rect 67 2641 245 2676
rect 67 2607 71 2641
rect 105 2607 139 2641
rect 173 2607 207 2641
rect 241 2607 245 2641
rect 67 2572 245 2607
rect 67 2538 71 2572
rect 105 2538 139 2572
rect 173 2538 207 2572
rect 241 2538 245 2572
rect 67 2503 245 2538
rect 67 2469 71 2503
rect 105 2469 139 2503
rect 173 2469 207 2503
rect 241 2469 245 2503
rect 67 2434 245 2469
rect 67 2400 71 2434
rect 105 2400 139 2434
rect 173 2400 207 2434
rect 241 2400 245 2434
rect 67 2365 245 2400
rect 67 2331 71 2365
rect 105 2331 139 2365
rect 173 2331 207 2365
rect 241 2331 245 2365
rect 67 2296 245 2331
rect 67 2262 71 2296
rect 105 2262 139 2296
rect 173 2262 207 2296
rect 241 2262 245 2296
rect 67 2227 245 2262
rect 67 2193 71 2227
rect 105 2193 139 2227
rect 173 2193 207 2227
rect 241 2193 245 2227
rect 67 2158 245 2193
rect 67 2124 71 2158
rect 105 2124 139 2158
rect 173 2124 207 2158
rect 241 2124 245 2158
rect 67 2089 245 2124
rect 67 2055 71 2089
rect 105 2055 139 2089
rect 173 2055 207 2089
rect 241 2055 245 2089
rect 67 2020 245 2055
rect 67 1986 71 2020
rect 105 1986 139 2020
rect 173 1986 207 2020
rect 241 1986 245 2020
rect 67 1951 245 1986
rect 67 1917 71 1951
rect 105 1917 139 1951
rect 173 1917 207 1951
rect 241 1917 245 1951
rect 67 1882 245 1917
rect 67 1848 71 1882
rect 105 1848 139 1882
rect 173 1848 207 1882
rect 241 1848 245 1882
rect 67 1813 245 1848
rect 67 1779 71 1813
rect 105 1779 139 1813
rect 173 1779 207 1813
rect 241 1779 245 1813
rect 67 1744 245 1779
rect 67 1710 71 1744
rect 105 1710 139 1744
rect 173 1710 207 1744
rect 241 1710 245 1744
rect 67 1675 245 1710
rect 67 1641 71 1675
rect 105 1641 139 1675
rect 173 1641 207 1675
rect 241 1641 245 1675
rect 67 1606 245 1641
rect 67 1572 71 1606
rect 105 1572 139 1606
rect 173 1572 207 1606
rect 241 1572 245 1606
rect 67 1537 245 1572
rect 67 1503 71 1537
rect 105 1503 139 1537
rect 173 1503 207 1537
rect 241 1503 245 1537
rect 67 1468 245 1503
rect 67 1434 71 1468
rect 105 1434 139 1468
rect 173 1434 207 1468
rect 241 1434 245 1468
rect 67 1399 245 1434
rect 67 1365 71 1399
rect 105 1365 139 1399
rect 173 1365 207 1399
rect 241 1365 245 1399
rect 67 1330 245 1365
rect 67 1296 71 1330
rect 105 1296 139 1330
rect 173 1296 207 1330
rect 241 1296 245 1330
rect 67 1261 245 1296
rect 67 1227 71 1261
rect 105 1227 139 1261
rect 173 1227 207 1261
rect 241 1227 245 1261
rect 67 1192 245 1227
rect 67 1158 71 1192
rect 105 1158 139 1192
rect 173 1158 207 1192
rect 241 1158 245 1192
rect 67 1123 245 1158
rect 67 545 71 1123
rect 241 668 245 1123
rect 14928 4934 14935 4968
rect 14969 4934 15003 4968
rect 15037 4934 15071 4968
rect 15105 4934 15106 4968
rect 14928 4896 15106 4934
rect 14928 4862 14935 4896
rect 14969 4862 15003 4896
rect 15037 4862 15071 4896
rect 15105 4862 15106 4896
rect 14928 4824 15106 4862
rect 14928 4790 14935 4824
rect 14969 4790 15003 4824
rect 15037 4790 15071 4824
rect 15105 4790 15106 4824
rect 14928 4752 15106 4790
rect 14928 4718 14935 4752
rect 14969 4718 15003 4752
rect 15037 4718 15071 4752
rect 15105 4718 15106 4752
rect 14928 4680 15106 4718
rect 14928 4646 14935 4680
rect 14969 4646 15003 4680
rect 15037 4646 15071 4680
rect 15105 4646 15106 4680
rect 14928 4608 15106 4646
rect 14928 4574 14935 4608
rect 14969 4574 15003 4608
rect 15037 4574 15071 4608
rect 15105 4574 15106 4608
rect 14928 4536 15106 4574
rect 14928 4502 14935 4536
rect 14969 4502 15003 4536
rect 15037 4502 15071 4536
rect 15105 4502 15106 4536
rect 14928 4464 15106 4502
rect 14928 4430 14935 4464
rect 14969 4430 15003 4464
rect 15037 4430 15071 4464
rect 15105 4430 15106 4464
rect 14928 4392 15106 4430
rect 14928 4358 14935 4392
rect 14969 4358 15003 4392
rect 15037 4358 15071 4392
rect 15105 4358 15106 4392
rect 14928 4320 15106 4358
rect 14928 4286 14935 4320
rect 14969 4286 15003 4320
rect 15037 4286 15071 4320
rect 15105 4286 15106 4320
rect 14928 4248 15106 4286
rect 14928 4214 14935 4248
rect 14969 4214 15003 4248
rect 15037 4214 15071 4248
rect 15105 4214 15106 4248
rect 14928 4176 15106 4214
rect 14928 4142 14935 4176
rect 14969 4142 15003 4176
rect 15037 4142 15071 4176
rect 15105 4142 15106 4176
rect 14928 4104 15106 4142
rect 14928 4070 14935 4104
rect 14969 4070 15003 4104
rect 15037 4070 15071 4104
rect 15105 4070 15106 4104
rect 14928 4032 15106 4070
rect 14928 3998 14935 4032
rect 14969 3998 15003 4032
rect 15037 3998 15071 4032
rect 15105 3998 15106 4032
rect 14928 3960 15106 3998
rect 14928 3926 14935 3960
rect 14969 3926 15003 3960
rect 15037 3926 15071 3960
rect 15105 3926 15106 3960
rect 14928 3888 15106 3926
rect 14928 3854 14935 3888
rect 14969 3854 15003 3888
rect 15037 3854 15071 3888
rect 15105 3854 15106 3888
rect 14928 3816 15106 3854
rect 14928 3782 14935 3816
rect 14969 3782 15003 3816
rect 15037 3782 15071 3816
rect 15105 3782 15106 3816
rect 14928 3744 15106 3782
rect 14928 3710 14935 3744
rect 14969 3710 15003 3744
rect 15037 3710 15071 3744
rect 15105 3710 15106 3744
rect 14928 3672 15106 3710
rect 14928 3638 14935 3672
rect 14969 3638 15003 3672
rect 15037 3638 15071 3672
rect 15105 3638 15106 3672
rect 14928 3600 15106 3638
rect 14928 3566 14935 3600
rect 14969 3566 15003 3600
rect 15037 3566 15071 3600
rect 15105 3566 15106 3600
rect 14928 3528 15106 3566
rect 14928 3494 14935 3528
rect 14969 3494 15003 3528
rect 15037 3494 15071 3528
rect 15105 3494 15106 3528
rect 14928 3456 15106 3494
rect 14928 3422 14935 3456
rect 14969 3422 15003 3456
rect 15037 3422 15071 3456
rect 15105 3422 15106 3456
rect 14928 3384 15106 3422
rect 14928 3350 14935 3384
rect 14969 3350 15003 3384
rect 15037 3350 15071 3384
rect 15105 3350 15106 3384
rect 14928 3312 15106 3350
rect 14928 3278 14935 3312
rect 14969 3278 15003 3312
rect 15037 3278 15071 3312
rect 15105 3278 15106 3312
rect 14928 3240 15106 3278
rect 14928 3206 14935 3240
rect 14969 3206 15003 3240
rect 15037 3206 15071 3240
rect 15105 3206 15106 3240
rect 14928 3168 15106 3206
rect 14928 3134 14935 3168
rect 14969 3134 15003 3168
rect 15037 3134 15071 3168
rect 15105 3134 15106 3168
rect 14928 3096 15106 3134
rect 14928 3062 14935 3096
rect 14969 3062 15003 3096
rect 15037 3062 15071 3096
rect 15105 3062 15106 3096
rect 14928 3024 15106 3062
rect 14928 2990 14935 3024
rect 14969 2990 15003 3024
rect 15037 2990 15071 3024
rect 15105 2990 15106 3024
rect 14928 2952 15106 2990
rect 14928 2918 14935 2952
rect 14969 2918 15003 2952
rect 15037 2918 15071 2952
rect 15105 2918 15106 2952
rect 14928 2880 15106 2918
rect 14928 2846 14935 2880
rect 14969 2846 15003 2880
rect 15037 2846 15071 2880
rect 15105 2846 15106 2880
rect 14928 2808 15106 2846
rect 14928 2774 14935 2808
rect 14969 2774 15003 2808
rect 15037 2774 15071 2808
rect 15105 2774 15106 2808
rect 14928 2736 15106 2774
rect 14928 2702 14935 2736
rect 14969 2702 15003 2736
rect 15037 2702 15071 2736
rect 15105 2702 15106 2736
rect 14928 2664 15106 2702
rect 14928 2630 14935 2664
rect 14969 2630 15003 2664
rect 15037 2630 15071 2664
rect 15105 2630 15106 2664
rect 14928 2592 15106 2630
rect 14928 2558 14935 2592
rect 14969 2558 15003 2592
rect 15037 2558 15071 2592
rect 15105 2558 15106 2592
rect 14928 2520 15106 2558
rect 14928 2486 14935 2520
rect 14969 2486 15003 2520
rect 15037 2486 15071 2520
rect 15105 2486 15106 2520
rect 14928 2448 15106 2486
rect 14928 2414 14935 2448
rect 14969 2414 15003 2448
rect 15037 2414 15071 2448
rect 15105 2414 15106 2448
rect 14928 2376 15106 2414
rect 14928 2342 14935 2376
rect 14969 2342 15003 2376
rect 15037 2342 15071 2376
rect 15105 2342 15106 2376
rect 14928 2304 15106 2342
rect 14928 2270 14935 2304
rect 14969 2270 15003 2304
rect 15037 2270 15071 2304
rect 15105 2270 15106 2304
rect 14928 2232 15106 2270
rect 14928 2198 14935 2232
rect 14969 2198 15003 2232
rect 15037 2198 15071 2232
rect 15105 2198 15106 2232
rect 14928 2160 15106 2198
rect 14928 2126 14935 2160
rect 14969 2126 15003 2160
rect 15037 2126 15071 2160
rect 15105 2126 15106 2160
rect 14928 2088 15106 2126
rect 14928 2054 14935 2088
rect 14969 2054 15003 2088
rect 15037 2054 15071 2088
rect 15105 2054 15106 2088
rect 14928 2016 15106 2054
rect 14928 1982 14935 2016
rect 14969 1982 15003 2016
rect 15037 1982 15071 2016
rect 15105 1982 15106 2016
rect 14928 1944 15106 1982
rect 14928 1910 14935 1944
rect 14969 1910 15003 1944
rect 15037 1910 15071 1944
rect 15105 1910 15106 1944
rect 14928 1872 15106 1910
rect 14928 1838 14935 1872
rect 14969 1838 15003 1872
rect 15037 1838 15071 1872
rect 15105 1838 15106 1872
rect 14928 1800 15106 1838
rect 14928 1766 14935 1800
rect 14969 1766 15003 1800
rect 15037 1766 15071 1800
rect 15105 1766 15106 1800
rect 14928 1728 15106 1766
rect 14928 1694 14935 1728
rect 14969 1694 15003 1728
rect 15037 1694 15071 1728
rect 15105 1694 15106 1728
rect 14928 1656 15106 1694
rect 14928 1622 14935 1656
rect 14969 1622 15003 1656
rect 15037 1622 15071 1656
rect 15105 1622 15106 1656
rect 14928 1584 15106 1622
rect 14928 1550 14935 1584
rect 14969 1550 15003 1584
rect 15037 1550 15071 1584
rect 15105 1550 15106 1584
rect 14928 1512 15106 1550
rect 14928 1478 14935 1512
rect 14969 1478 15003 1512
rect 15037 1478 15071 1512
rect 15105 1478 15106 1512
rect 14928 1440 15106 1478
rect 14928 1406 14935 1440
rect 14969 1406 15003 1440
rect 15037 1406 15071 1440
rect 15105 1406 15106 1440
rect 14928 1368 15106 1406
rect 14928 1334 14935 1368
rect 14969 1334 15003 1368
rect 15037 1334 15071 1368
rect 15105 1334 15106 1368
rect 14928 1296 15106 1334
rect 14928 1262 14935 1296
rect 14969 1262 15003 1296
rect 15037 1262 15071 1296
rect 15105 1262 15106 1296
rect 14928 1224 15106 1262
rect 14928 1190 14935 1224
rect 14969 1190 15003 1224
rect 15037 1190 15071 1224
rect 15105 1190 15106 1224
rect 14928 1152 15106 1190
rect 14928 1118 14935 1152
rect 14969 1118 15003 1152
rect 15037 1118 15071 1152
rect 15105 1118 15106 1152
rect 14928 1080 15106 1118
rect 14928 1046 14935 1080
rect 14969 1046 15003 1080
rect 15037 1046 15071 1080
rect 15105 1046 15106 1080
rect 14928 1008 15106 1046
rect 14928 974 14935 1008
rect 14969 974 15003 1008
rect 15037 974 15071 1008
rect 15105 974 15106 1008
rect 14928 936 15106 974
rect 14928 902 14935 936
rect 14969 902 15003 936
rect 15037 902 15071 936
rect 15105 902 15106 936
rect 14928 864 15106 902
rect 14928 830 14935 864
rect 14969 830 15003 864
rect 15037 830 15071 864
rect 15105 830 15106 864
rect 14928 792 15106 830
rect 14928 758 14935 792
rect 14969 758 15003 792
rect 15037 758 15071 792
rect 15105 758 15106 792
rect 14928 720 15106 758
rect 14928 686 14935 720
rect 14969 686 15003 720
rect 15037 686 15071 720
rect 15105 686 15106 720
rect 14928 668 15106 686
rect 241 664 15106 668
rect 241 630 294 664
rect 328 630 363 664
rect 397 630 432 664
rect 466 630 501 664
rect 535 630 570 664
rect 604 630 639 664
rect 673 630 708 664
rect 742 630 777 664
rect 811 630 846 664
rect 880 630 915 664
rect 949 630 984 664
rect 1018 630 1053 664
rect 1087 630 1122 664
rect 1156 630 1191 664
rect 1225 630 1260 664
rect 1294 630 1329 664
rect 1363 630 1398 664
rect 1432 630 1467 664
rect 1501 630 1536 664
rect 1570 630 1605 664
rect 1639 630 1674 664
rect 1708 630 1743 664
rect 1777 630 1812 664
rect 1846 630 1881 664
rect 1915 630 1950 664
rect 1984 630 2019 664
rect 2053 630 2088 664
rect 2122 630 2157 664
rect 2191 630 2226 664
rect 2260 630 2295 664
rect 2329 630 2364 664
rect 2398 630 2433 664
rect 2467 630 2502 664
rect 2536 630 2571 664
rect 2605 630 2640 664
rect 2674 630 2709 664
rect 2743 630 2778 664
rect 2812 630 2847 664
rect 2881 630 2916 664
rect 2950 630 2985 664
rect 3019 630 3054 664
rect 3088 630 3123 664
rect 3157 630 3192 664
rect 3226 630 3261 664
rect 3295 630 3330 664
rect 3364 630 3399 664
rect 3433 630 3468 664
rect 3502 630 3537 664
rect 3571 630 3606 664
rect 3640 630 3675 664
rect 3709 630 3744 664
rect 3778 630 3813 664
rect 3847 630 3882 664
rect 3916 630 3951 664
rect 3985 630 4020 664
rect 4054 630 4089 664
rect 4123 630 4158 664
rect 4192 630 4227 664
rect 4261 630 4296 664
rect 4330 630 4365 664
rect 4399 630 4434 664
rect 4468 630 4503 664
rect 4537 630 4572 664
rect 4606 630 4641 664
rect 4675 630 4710 664
rect 241 596 4710 630
rect 241 562 294 596
rect 328 562 363 596
rect 397 562 432 596
rect 466 562 501 596
rect 535 562 570 596
rect 604 562 639 596
rect 673 562 708 596
rect 742 562 777 596
rect 811 562 846 596
rect 880 562 915 596
rect 949 562 984 596
rect 1018 562 1053 596
rect 1087 562 1122 596
rect 1156 562 1191 596
rect 1225 562 1260 596
rect 1294 562 1329 596
rect 1363 562 1398 596
rect 1432 562 1467 596
rect 1501 562 1536 596
rect 1570 562 1605 596
rect 1639 562 1674 596
rect 1708 562 1743 596
rect 1777 562 1812 596
rect 1846 562 1881 596
rect 1915 562 1950 596
rect 1984 562 2019 596
rect 2053 562 2088 596
rect 2122 562 2157 596
rect 2191 562 2226 596
rect 2260 562 2295 596
rect 2329 562 2364 596
rect 2398 562 2433 596
rect 2467 562 2502 596
rect 2536 562 2571 596
rect 2605 562 2640 596
rect 2674 562 2709 596
rect 2743 562 2778 596
rect 2812 562 2847 596
rect 2881 562 2916 596
rect 2950 562 2985 596
rect 3019 562 3054 596
rect 3088 562 3123 596
rect 3157 562 3192 596
rect 3226 562 3261 596
rect 3295 562 3330 596
rect 3364 562 3399 596
rect 3433 562 3468 596
rect 3502 562 3537 596
rect 3571 562 3606 596
rect 3640 562 3675 596
rect 3709 562 3744 596
rect 3778 562 3813 596
rect 3847 562 3882 596
rect 3916 562 3951 596
rect 3985 562 4020 596
rect 4054 562 4089 596
rect 4123 562 4158 596
rect 4192 562 4227 596
rect 4261 562 4296 596
rect 4330 562 4365 596
rect 4399 562 4434 596
rect 4468 562 4503 596
rect 4537 562 4572 596
rect 4606 562 4641 596
rect 4675 562 4710 596
rect 241 545 4710 562
rect 67 528 4710 545
rect 67 494 294 528
rect 328 494 363 528
rect 397 494 432 528
rect 466 494 501 528
rect 535 494 570 528
rect 604 494 639 528
rect 673 494 708 528
rect 742 494 777 528
rect 811 494 846 528
rect 880 494 915 528
rect 949 494 984 528
rect 1018 494 1053 528
rect 1087 494 1122 528
rect 1156 494 1191 528
rect 1225 494 1260 528
rect 1294 494 1329 528
rect 1363 494 1398 528
rect 1432 494 1467 528
rect 1501 494 1536 528
rect 1570 494 1605 528
rect 1639 494 1674 528
rect 1708 494 1743 528
rect 1777 494 1812 528
rect 1846 494 1881 528
rect 1915 494 1950 528
rect 1984 494 2019 528
rect 2053 494 2088 528
rect 2122 494 2157 528
rect 2191 494 2226 528
rect 2260 494 2295 528
rect 2329 494 2364 528
rect 2398 494 2433 528
rect 2467 494 2502 528
rect 2536 494 2571 528
rect 2605 494 2640 528
rect 2674 494 2709 528
rect 2743 494 2778 528
rect 2812 494 2847 528
rect 2881 494 2916 528
rect 2950 494 2985 528
rect 3019 494 3054 528
rect 3088 494 3123 528
rect 3157 494 3192 528
rect 3226 494 3261 528
rect 3295 494 3330 528
rect 3364 494 3399 528
rect 3433 494 3468 528
rect 3502 494 3537 528
rect 3571 494 3606 528
rect 3640 494 3675 528
rect 3709 494 3744 528
rect 3778 494 3813 528
rect 3847 494 3882 528
rect 3916 494 3951 528
rect 3985 494 4020 528
rect 4054 494 4089 528
rect 4123 494 4158 528
rect 4192 494 4227 528
rect 4261 494 4296 528
rect 4330 494 4365 528
rect 4399 494 4434 528
rect 4468 494 4503 528
rect 4537 494 4572 528
rect 4606 494 4641 528
rect 4675 494 4710 528
rect 14876 648 15106 664
rect 14876 614 14935 648
rect 14969 614 15003 648
rect 15037 614 15071 648
rect 15105 614 15106 648
rect 14876 576 15106 614
rect 14876 542 14935 576
rect 14969 542 15003 576
rect 15037 542 15071 576
rect 15105 542 15106 576
rect 14876 494 15106 542
rect 67 490 15106 494
<< mvpsubdiffcont >>
rect 657 4922 14495 4956
rect 14530 4922 14564 4956
rect 14599 4922 14633 4956
rect 555 4888 589 4922
rect 657 4888 14461 4922
rect 623 4854 14461 4888
rect 14496 4854 14530 4888
rect 14565 4854 14599 4888
rect 555 4816 589 4850
rect 623 4785 657 4819
rect 691 4786 14393 4854
rect 14428 4786 14462 4820
rect 14497 4786 14531 4820
rect 555 4744 589 4778
rect 623 4716 657 4750
rect 691 4717 725 4751
rect 555 4672 589 4706
rect 623 4647 657 4681
rect 691 4648 725 4682
rect 555 4600 589 4634
rect 555 4529 589 4563
rect 555 4458 589 4492
rect 555 4387 589 4421
rect 555 4316 589 4350
rect 555 4245 589 4279
rect 555 4174 589 4208
rect 555 4103 589 4137
rect 623 4103 725 4613
rect 14565 4784 14599 4818
rect 14633 4810 14667 4844
rect 14497 4716 14531 4750
rect 14565 4714 14599 4748
rect 14633 4737 14667 4771
rect 14497 4646 14531 4680
rect 14565 4644 14599 4678
rect 14633 4664 14667 4698
rect 14497 4576 14531 4610
rect 14565 4574 14599 4608
rect 14633 4591 14667 4625
rect 14497 4506 14531 4540
rect 14565 4504 14599 4538
rect 14633 4518 14667 4552
rect 14497 4436 14531 4470
rect 14565 4434 14599 4468
rect 14633 4445 14667 4479
rect 14497 4365 14531 4399
rect 14565 4364 14599 4398
rect 14633 4372 14667 4406
rect 14497 4294 14531 4328
rect 14565 4294 14599 4328
rect 14633 4299 14667 4333
rect 14497 4223 14531 4257
rect 14565 4223 14599 4257
rect 14633 4226 14667 4260
rect 14497 4152 14531 4186
rect 14565 4152 14599 4186
rect 14633 4152 14667 4186
rect 14565 4081 14599 4115
rect 14633 4081 14667 4115
rect 555 4007 589 4041
rect 623 4007 657 4041
rect 734 4000 768 4034
rect 555 3936 589 3970
rect 623 3936 657 3970
rect 734 3932 768 3966
rect 555 3862 589 3896
rect 623 3862 657 3896
rect 734 3864 768 3898
rect 555 3791 589 3825
rect 623 3791 657 3825
rect 734 3796 768 3830
rect 555 3717 589 3751
rect 623 3717 657 3751
rect 734 3728 768 3762
rect 555 3646 589 3680
rect 623 3646 657 3680
rect 734 3660 768 3694
rect 555 3572 589 3606
rect 623 3572 657 3606
rect 734 3592 768 3626
rect 555 3501 589 3535
rect 623 3501 657 3535
rect 734 3524 768 3558
rect 555 3427 589 3461
rect 623 3427 657 3461
rect 734 3456 768 3490
rect 555 3356 589 3390
rect 623 3356 657 3390
rect 734 3388 768 3422
rect 734 3320 768 3354
rect 555 3282 589 3316
rect 623 3282 657 3316
rect 734 3252 768 3286
rect 555 3211 589 3245
rect 623 3211 657 3245
rect 734 3184 768 3218
rect 555 3117 589 3151
rect 623 3117 657 3151
rect 734 3116 768 3150
rect 555 3013 657 3081
rect 1678 4012 1712 4046
rect 1678 3944 1712 3978
rect 1678 3876 1712 3910
rect 1678 3808 1712 3842
rect 1678 3740 1712 3774
rect 1678 3672 1712 3706
rect 1678 3604 1712 3638
rect 1678 3536 1712 3570
rect 1678 3468 1712 3502
rect 1678 3400 1712 3434
rect 1678 3332 1712 3366
rect 1678 3264 1712 3298
rect 1678 3196 1712 3230
rect 1678 3128 1712 3162
rect 2670 4012 2704 4046
rect 2670 3944 2704 3978
rect 2670 3876 2704 3910
rect 2670 3808 2704 3842
rect 2670 3740 2704 3774
rect 2670 3672 2704 3706
rect 2670 3604 2704 3638
rect 2670 3536 2704 3570
rect 2670 3468 2704 3502
rect 2670 3400 2704 3434
rect 2670 3332 2704 3366
rect 2670 3264 2704 3298
rect 2670 3196 2704 3230
rect 2670 3128 2704 3162
rect 3662 4012 3696 4046
rect 3662 3944 3696 3978
rect 3662 3876 3696 3910
rect 3662 3808 3696 3842
rect 3662 3740 3696 3774
rect 3662 3672 3696 3706
rect 3662 3604 3696 3638
rect 3662 3536 3696 3570
rect 3662 3468 3696 3502
rect 3662 3400 3696 3434
rect 3662 3332 3696 3366
rect 3662 3264 3696 3298
rect 3662 3196 3696 3230
rect 3662 3128 3696 3162
rect 4654 4012 4688 4046
rect 4654 3944 4688 3978
rect 4654 3876 4688 3910
rect 4654 3808 4688 3842
rect 4654 3740 4688 3774
rect 4654 3672 4688 3706
rect 4654 3604 4688 3638
rect 4654 3536 4688 3570
rect 4654 3468 4688 3502
rect 4654 3400 4688 3434
rect 4654 3332 4688 3366
rect 4654 3264 4688 3298
rect 4654 3196 4688 3230
rect 4654 3128 4688 3162
rect 5646 4012 5680 4046
rect 5646 3944 5680 3978
rect 5646 3876 5680 3910
rect 5646 3808 5680 3842
rect 5646 3740 5680 3774
rect 5646 3672 5680 3706
rect 5646 3604 5680 3638
rect 5646 3536 5680 3570
rect 5646 3468 5680 3502
rect 5646 3400 5680 3434
rect 5646 3332 5680 3366
rect 5646 3264 5680 3298
rect 5646 3196 5680 3230
rect 5646 3128 5680 3162
rect 6638 4012 6672 4046
rect 6638 3944 6672 3978
rect 6638 3876 6672 3910
rect 6638 3808 6672 3842
rect 6638 3740 6672 3774
rect 6638 3672 6672 3706
rect 6638 3604 6672 3638
rect 6638 3536 6672 3570
rect 6638 3468 6672 3502
rect 6638 3400 6672 3434
rect 6638 3332 6672 3366
rect 6638 3264 6672 3298
rect 6638 3196 6672 3230
rect 6638 3128 6672 3162
rect 7630 4012 7664 4046
rect 7630 3944 7664 3978
rect 7630 3876 7664 3910
rect 7630 3808 7664 3842
rect 7630 3740 7664 3774
rect 7630 3672 7664 3706
rect 7630 3604 7664 3638
rect 7630 3536 7664 3570
rect 7630 3468 7664 3502
rect 7630 3400 7664 3434
rect 7630 3332 7664 3366
rect 7630 3264 7664 3298
rect 7630 3196 7664 3230
rect 7630 3128 7664 3162
rect 8622 4012 8656 4046
rect 8622 3944 8656 3978
rect 8622 3876 8656 3910
rect 8622 3808 8656 3842
rect 8622 3740 8656 3774
rect 8622 3672 8656 3706
rect 8622 3604 8656 3638
rect 8622 3536 8656 3570
rect 8622 3468 8656 3502
rect 8622 3400 8656 3434
rect 8622 3332 8656 3366
rect 8622 3264 8656 3298
rect 8622 3196 8656 3230
rect 8622 3128 8656 3162
rect 9614 4012 9648 4046
rect 9614 3944 9648 3978
rect 9614 3876 9648 3910
rect 9614 3808 9648 3842
rect 9614 3740 9648 3774
rect 9614 3672 9648 3706
rect 9614 3604 9648 3638
rect 9614 3536 9648 3570
rect 9614 3468 9648 3502
rect 9614 3400 9648 3434
rect 9614 3332 9648 3366
rect 9614 3264 9648 3298
rect 9614 3196 9648 3230
rect 9614 3128 9648 3162
rect 10606 4012 10640 4046
rect 10606 3944 10640 3978
rect 10606 3876 10640 3910
rect 10606 3808 10640 3842
rect 10606 3740 10640 3774
rect 10606 3672 10640 3706
rect 10606 3604 10640 3638
rect 10606 3536 10640 3570
rect 10606 3468 10640 3502
rect 10606 3400 10640 3434
rect 10606 3332 10640 3366
rect 10606 3264 10640 3298
rect 10606 3196 10640 3230
rect 10606 3128 10640 3162
rect 11598 4012 11632 4046
rect 11598 3944 11632 3978
rect 11598 3876 11632 3910
rect 11598 3808 11632 3842
rect 11598 3740 11632 3774
rect 11598 3672 11632 3706
rect 11598 3604 11632 3638
rect 11598 3536 11632 3570
rect 11598 3468 11632 3502
rect 11598 3400 11632 3434
rect 11598 3332 11632 3366
rect 11598 3264 11632 3298
rect 11598 3196 11632 3230
rect 11598 3128 11632 3162
rect 12590 4012 12624 4046
rect 12590 3944 12624 3978
rect 12590 3876 12624 3910
rect 12590 3808 12624 3842
rect 12590 3740 12624 3774
rect 12590 3672 12624 3706
rect 12590 3604 12624 3638
rect 12590 3536 12624 3570
rect 12590 3468 12624 3502
rect 12590 3400 12624 3434
rect 12590 3332 12624 3366
rect 12590 3264 12624 3298
rect 12590 3196 12624 3230
rect 12590 3128 12624 3162
rect 13582 4012 13616 4046
rect 13582 3944 13616 3978
rect 13582 3876 13616 3910
rect 13582 3808 13616 3842
rect 13582 3740 13616 3774
rect 13582 3672 13616 3706
rect 13582 3604 13616 3638
rect 13582 3536 13616 3570
rect 13582 3468 13616 3502
rect 13582 3400 13616 3434
rect 13582 3332 13616 3366
rect 13582 3264 13616 3298
rect 13582 3196 13616 3230
rect 13582 3128 13616 3162
rect 14454 4000 14488 4034
rect 14565 4007 14599 4041
rect 14633 4007 14667 4041
rect 14454 3932 14488 3966
rect 14565 3936 14599 3970
rect 14633 3936 14667 3970
rect 14454 3864 14488 3898
rect 14565 3862 14599 3896
rect 14633 3862 14667 3896
rect 14454 3796 14488 3830
rect 14565 3791 14599 3825
rect 14633 3791 14667 3825
rect 14454 3728 14488 3762
rect 14565 3717 14599 3751
rect 14633 3717 14667 3751
rect 14454 3660 14488 3694
rect 14565 3646 14599 3680
rect 14633 3646 14667 3680
rect 14454 3592 14488 3626
rect 14565 3572 14599 3606
rect 14633 3572 14667 3606
rect 14454 3524 14488 3558
rect 14565 3501 14599 3535
rect 14633 3501 14667 3535
rect 14454 3456 14488 3490
rect 14565 3427 14599 3461
rect 14633 3427 14667 3461
rect 14454 3388 14488 3422
rect 14565 3356 14599 3390
rect 14633 3356 14667 3390
rect 14454 3320 14488 3354
rect 14454 3252 14488 3286
rect 14565 3282 14599 3316
rect 14633 3282 14667 3316
rect 14454 3184 14488 3218
rect 14565 3211 14599 3245
rect 14633 3211 14667 3245
rect 14454 3116 14488 3150
rect 14565 3117 14599 3151
rect 14633 3117 14667 3151
rect 555 2503 725 3013
rect 555 2367 657 2503
rect 1645 2901 1679 2935
rect 1713 2901 1747 2935
rect 1645 2821 1679 2855
rect 1713 2821 1747 2855
rect 1645 2741 1679 2775
rect 1713 2741 1747 2775
rect 1645 2661 1679 2695
rect 1713 2661 1747 2695
rect 1645 2580 1679 2614
rect 1713 2580 1747 2614
rect 2637 2901 2671 2935
rect 2705 2901 2739 2935
rect 2637 2821 2671 2855
rect 2705 2821 2739 2855
rect 2637 2741 2671 2775
rect 2705 2741 2739 2775
rect 2637 2661 2671 2695
rect 2705 2661 2739 2695
rect 2637 2580 2671 2614
rect 2705 2580 2739 2614
rect 3629 2901 3663 2935
rect 3697 2901 3731 2935
rect 3629 2821 3663 2855
rect 3697 2821 3731 2855
rect 3629 2741 3663 2775
rect 3697 2741 3731 2775
rect 3629 2661 3663 2695
rect 3697 2661 3731 2695
rect 3629 2580 3663 2614
rect 3697 2580 3731 2614
rect 4621 2901 4655 2935
rect 4689 2901 4723 2935
rect 4621 2821 4655 2855
rect 4689 2821 4723 2855
rect 4621 2741 4655 2775
rect 4689 2741 4723 2775
rect 4621 2661 4655 2695
rect 4689 2661 4723 2695
rect 4621 2580 4655 2614
rect 4689 2580 4723 2614
rect 5613 2901 5647 2935
rect 5681 2901 5715 2935
rect 5613 2821 5647 2855
rect 5681 2821 5715 2855
rect 5613 2741 5647 2775
rect 5681 2741 5715 2775
rect 5613 2661 5647 2695
rect 5681 2661 5715 2695
rect 5613 2580 5647 2614
rect 5681 2580 5715 2614
rect 6605 2901 6639 2935
rect 6673 2901 6707 2935
rect 6605 2821 6639 2855
rect 6673 2821 6707 2855
rect 6605 2741 6639 2775
rect 6673 2741 6707 2775
rect 6605 2661 6639 2695
rect 6673 2661 6707 2695
rect 6605 2580 6639 2614
rect 6673 2580 6707 2614
rect 7597 2901 7631 2935
rect 7665 2901 7699 2935
rect 7597 2821 7631 2855
rect 7665 2821 7699 2855
rect 7597 2741 7631 2775
rect 7665 2741 7699 2775
rect 7597 2661 7631 2695
rect 7665 2661 7699 2695
rect 7597 2580 7631 2614
rect 7665 2580 7699 2614
rect 8589 2901 8623 2935
rect 8657 2901 8691 2935
rect 8589 2821 8623 2855
rect 8657 2821 8691 2855
rect 8589 2741 8623 2775
rect 8657 2741 8691 2775
rect 8589 2661 8623 2695
rect 8657 2661 8691 2695
rect 8589 2580 8623 2614
rect 8657 2580 8691 2614
rect 9581 2901 9615 2935
rect 9649 2901 9683 2935
rect 9581 2821 9615 2855
rect 9649 2821 9683 2855
rect 9581 2741 9615 2775
rect 9649 2741 9683 2775
rect 9581 2661 9615 2695
rect 9649 2661 9683 2695
rect 9581 2580 9615 2614
rect 9649 2580 9683 2614
rect 10573 2901 10607 2935
rect 10641 2901 10675 2935
rect 10573 2821 10607 2855
rect 10641 2821 10675 2855
rect 10573 2741 10607 2775
rect 10641 2741 10675 2775
rect 10573 2661 10607 2695
rect 10641 2661 10675 2695
rect 10573 2580 10607 2614
rect 10641 2580 10675 2614
rect 11565 2901 11599 2935
rect 11633 2901 11667 2935
rect 11565 2821 11599 2855
rect 11633 2821 11667 2855
rect 11565 2741 11599 2775
rect 11633 2741 11667 2775
rect 11565 2661 11599 2695
rect 11633 2661 11667 2695
rect 11565 2580 11599 2614
rect 11633 2580 11667 2614
rect 12557 2901 12591 2935
rect 12625 2901 12659 2935
rect 12557 2821 12591 2855
rect 12625 2821 12659 2855
rect 12557 2741 12591 2775
rect 12625 2741 12659 2775
rect 12557 2661 12591 2695
rect 12625 2661 12659 2695
rect 12557 2580 12591 2614
rect 12625 2580 12659 2614
rect 13549 2901 13583 2935
rect 13617 2901 13651 2935
rect 13549 2821 13583 2855
rect 13617 2821 13651 2855
rect 13549 2741 13583 2775
rect 13617 2741 13651 2775
rect 13549 2661 13583 2695
rect 13617 2661 13651 2695
rect 13549 2580 13583 2614
rect 13617 2580 13651 2614
rect 14565 3032 14599 3066
rect 14633 3032 14667 3066
rect 14497 2530 14667 2972
rect 734 2399 768 2433
rect 734 2331 768 2365
rect 555 2293 589 2327
rect 623 2293 657 2327
rect 734 2263 768 2297
rect 555 2216 589 2250
rect 623 2216 657 2250
rect 734 2195 768 2229
rect 555 2122 589 2156
rect 623 2122 657 2156
rect 734 2127 768 2161
rect 555 2051 589 2085
rect 623 2051 657 2085
rect 734 2059 768 2093
rect 555 1977 589 2011
rect 623 1977 657 2011
rect 734 1991 768 2025
rect 555 1906 589 1940
rect 623 1906 657 1940
rect 734 1923 768 1957
rect 555 1832 589 1866
rect 623 1832 657 1866
rect 734 1855 768 1889
rect 555 1761 589 1795
rect 623 1761 657 1795
rect 734 1787 768 1821
rect 555 1687 589 1721
rect 623 1687 657 1721
rect 734 1719 768 1753
rect 734 1651 768 1685
rect 555 1616 589 1650
rect 623 1616 657 1650
rect 734 1583 768 1617
rect 555 1542 589 1576
rect 623 1542 657 1576
rect 734 1515 768 1549
rect 555 1471 589 1505
rect 623 1471 657 1505
rect 1678 2411 1712 2445
rect 1678 2343 1712 2377
rect 1678 2275 1712 2309
rect 1678 2207 1712 2241
rect 1678 2139 1712 2173
rect 1678 2071 1712 2105
rect 1678 2003 1712 2037
rect 1678 1935 1712 1969
rect 1678 1867 1712 1901
rect 1678 1799 1712 1833
rect 1678 1731 1712 1765
rect 1678 1663 1712 1697
rect 1678 1595 1712 1629
rect 1678 1527 1712 1561
rect 2670 2411 2704 2445
rect 2670 2343 2704 2377
rect 2670 2275 2704 2309
rect 2670 2207 2704 2241
rect 2670 2139 2704 2173
rect 2670 2071 2704 2105
rect 2670 2003 2704 2037
rect 2670 1935 2704 1969
rect 2670 1867 2704 1901
rect 2670 1799 2704 1833
rect 2670 1731 2704 1765
rect 2670 1663 2704 1697
rect 2670 1595 2704 1629
rect 2670 1527 2704 1561
rect 3662 2411 3696 2445
rect 3662 2343 3696 2377
rect 3662 2275 3696 2309
rect 3662 2207 3696 2241
rect 3662 2139 3696 2173
rect 3662 2071 3696 2105
rect 3662 2003 3696 2037
rect 3662 1935 3696 1969
rect 3662 1867 3696 1901
rect 3662 1799 3696 1833
rect 3662 1731 3696 1765
rect 3662 1663 3696 1697
rect 3662 1595 3696 1629
rect 3662 1527 3696 1561
rect 4654 2411 4688 2445
rect 4654 2343 4688 2377
rect 4654 2275 4688 2309
rect 4654 2207 4688 2241
rect 4654 2139 4688 2173
rect 4654 2071 4688 2105
rect 4654 2003 4688 2037
rect 4654 1935 4688 1969
rect 4654 1867 4688 1901
rect 4654 1799 4688 1833
rect 4654 1731 4688 1765
rect 4654 1663 4688 1697
rect 4654 1595 4688 1629
rect 4654 1527 4688 1561
rect 5646 2411 5680 2445
rect 5646 2343 5680 2377
rect 5646 2275 5680 2309
rect 5646 2207 5680 2241
rect 5646 2139 5680 2173
rect 5646 2071 5680 2105
rect 5646 2003 5680 2037
rect 5646 1935 5680 1969
rect 5646 1867 5680 1901
rect 5646 1799 5680 1833
rect 5646 1731 5680 1765
rect 5646 1663 5680 1697
rect 5646 1595 5680 1629
rect 5646 1527 5680 1561
rect 6638 2411 6672 2445
rect 6638 2343 6672 2377
rect 6638 2275 6672 2309
rect 6638 2207 6672 2241
rect 6638 2139 6672 2173
rect 6638 2071 6672 2105
rect 6638 2003 6672 2037
rect 6638 1935 6672 1969
rect 6638 1867 6672 1901
rect 6638 1799 6672 1833
rect 6638 1731 6672 1765
rect 6638 1663 6672 1697
rect 6638 1595 6672 1629
rect 6638 1527 6672 1561
rect 7630 2411 7664 2445
rect 7630 2343 7664 2377
rect 7630 2275 7664 2309
rect 7630 2207 7664 2241
rect 7630 2139 7664 2173
rect 7630 2071 7664 2105
rect 7630 2003 7664 2037
rect 7630 1935 7664 1969
rect 7630 1867 7664 1901
rect 7630 1799 7664 1833
rect 7630 1731 7664 1765
rect 7630 1663 7664 1697
rect 7630 1595 7664 1629
rect 7630 1527 7664 1561
rect 8622 2411 8656 2445
rect 8622 2343 8656 2377
rect 8622 2275 8656 2309
rect 8622 2207 8656 2241
rect 8622 2139 8656 2173
rect 8622 2071 8656 2105
rect 8622 2003 8656 2037
rect 8622 1935 8656 1969
rect 8622 1867 8656 1901
rect 8622 1799 8656 1833
rect 8622 1731 8656 1765
rect 8622 1663 8656 1697
rect 8622 1595 8656 1629
rect 8622 1527 8656 1561
rect 9614 2411 9648 2445
rect 9614 2343 9648 2377
rect 9614 2275 9648 2309
rect 9614 2207 9648 2241
rect 9614 2139 9648 2173
rect 9614 2071 9648 2105
rect 9614 2003 9648 2037
rect 9614 1935 9648 1969
rect 9614 1867 9648 1901
rect 9614 1799 9648 1833
rect 9614 1731 9648 1765
rect 9614 1663 9648 1697
rect 9614 1595 9648 1629
rect 9614 1527 9648 1561
rect 10606 2411 10640 2445
rect 10606 2343 10640 2377
rect 10606 2275 10640 2309
rect 10606 2207 10640 2241
rect 10606 2139 10640 2173
rect 10606 2071 10640 2105
rect 10606 2003 10640 2037
rect 10606 1935 10640 1969
rect 10606 1867 10640 1901
rect 10606 1799 10640 1833
rect 10606 1731 10640 1765
rect 10606 1663 10640 1697
rect 10606 1595 10640 1629
rect 10606 1527 10640 1561
rect 11598 2411 11632 2445
rect 11598 2343 11632 2377
rect 11598 2275 11632 2309
rect 11598 2207 11632 2241
rect 11598 2139 11632 2173
rect 11598 2071 11632 2105
rect 11598 2003 11632 2037
rect 11598 1935 11632 1969
rect 11598 1867 11632 1901
rect 11598 1799 11632 1833
rect 11598 1731 11632 1765
rect 11598 1663 11632 1697
rect 11598 1595 11632 1629
rect 11598 1527 11632 1561
rect 12590 2411 12624 2445
rect 12590 2343 12624 2377
rect 12590 2275 12624 2309
rect 12590 2207 12624 2241
rect 12590 2139 12624 2173
rect 12590 2071 12624 2105
rect 12590 2003 12624 2037
rect 12590 1935 12624 1969
rect 12590 1867 12624 1901
rect 12590 1799 12624 1833
rect 12590 1731 12624 1765
rect 12590 1663 12624 1697
rect 12590 1595 12624 1629
rect 12590 1527 12624 1561
rect 13582 2411 13616 2445
rect 13582 2343 13616 2377
rect 13582 2275 13616 2309
rect 13582 2207 13616 2241
rect 13582 2139 13616 2173
rect 13582 2071 13616 2105
rect 13582 2003 13616 2037
rect 13582 1935 13616 1969
rect 13582 1867 13616 1901
rect 13582 1799 13616 1833
rect 13582 1731 13616 1765
rect 13582 1663 13616 1697
rect 13582 1595 13616 1629
rect 13582 1527 13616 1561
rect 14565 2451 14599 2485
rect 14633 2451 14667 2485
rect 14454 2399 14488 2433
rect 14565 2369 14599 2403
rect 14633 2369 14667 2403
rect 14454 2331 14488 2365
rect 14454 2263 14488 2297
rect 14565 2293 14599 2327
rect 14633 2293 14667 2327
rect 14454 2195 14488 2229
rect 14565 2216 14599 2250
rect 14633 2216 14667 2250
rect 14454 2127 14488 2161
rect 14565 2122 14599 2156
rect 14633 2122 14667 2156
rect 14454 2059 14488 2093
rect 14565 2051 14599 2085
rect 14633 2051 14667 2085
rect 14454 1991 14488 2025
rect 14565 1977 14599 2011
rect 14633 1977 14667 2011
rect 14454 1923 14488 1957
rect 14565 1906 14599 1940
rect 14633 1906 14667 1940
rect 14454 1855 14488 1889
rect 14565 1832 14599 1866
rect 14633 1832 14667 1866
rect 14454 1787 14488 1821
rect 14565 1761 14599 1795
rect 14633 1761 14667 1795
rect 14454 1719 14488 1753
rect 14565 1687 14599 1721
rect 14633 1687 14667 1721
rect 14454 1651 14488 1685
rect 14454 1583 14488 1617
rect 14565 1616 14599 1650
rect 14633 1616 14667 1650
rect 14454 1515 14488 1549
rect 14565 1542 14599 1576
rect 14633 1542 14667 1576
rect 14565 1471 14599 1505
rect 14633 1471 14667 1505
rect 555 1341 589 1375
rect 623 1341 657 1375
rect 691 1341 725 1375
rect 14497 1353 14531 1387
rect 14565 1353 14599 1387
rect 14633 1353 14667 1387
rect 555 1187 589 1221
rect 623 1187 657 1221
rect 691 1185 725 1219
rect 555 1106 589 1140
rect 623 1116 657 1150
rect 14497 1274 14531 1308
rect 14565 1277 14599 1311
rect 14633 1285 14667 1319
rect 14497 1194 14531 1228
rect 14565 1200 14599 1234
rect 14633 1217 14667 1251
rect 691 1114 725 1148
rect 760 1114 794 1148
rect 829 1080 14531 1148
rect 14565 1123 14599 1157
rect 14633 1149 14667 1183
rect 14633 1081 14667 1115
rect 623 1046 657 1080
rect 692 1046 726 1080
rect 761 1046 14599 1080
rect 761 1012 14565 1046
rect 14633 1012 14667 1046
rect 589 978 623 1012
rect 658 978 692 1012
rect 727 978 14565 1012
<< mvnsubdiffcont >>
rect 71 5269 105 5303
rect 139 5269 173 5303
rect 207 5269 241 5303
rect 294 5252 10868 5422
rect 10903 5388 10937 5422
rect 10972 5388 11006 5422
rect 11041 5388 11075 5422
rect 11110 5388 11144 5422
rect 11179 5388 11213 5422
rect 11248 5388 11282 5422
rect 11317 5388 11351 5422
rect 11386 5388 11420 5422
rect 11455 5388 11489 5422
rect 11524 5388 11558 5422
rect 11593 5388 11627 5422
rect 11662 5388 11696 5422
rect 11731 5388 11765 5422
rect 11800 5388 11834 5422
rect 11869 5388 11903 5422
rect 11938 5388 11972 5422
rect 12007 5388 12041 5422
rect 12076 5388 12110 5422
rect 12145 5388 12179 5422
rect 12214 5388 12248 5422
rect 12283 5388 12317 5422
rect 12352 5388 12386 5422
rect 12421 5388 12455 5422
rect 12490 5388 12524 5422
rect 12559 5388 12593 5422
rect 12628 5388 12662 5422
rect 12697 5388 12731 5422
rect 12766 5388 12800 5422
rect 12835 5388 12869 5422
rect 12904 5388 12938 5422
rect 12973 5388 13007 5422
rect 13042 5388 13076 5422
rect 13111 5388 13145 5422
rect 13180 5388 13214 5422
rect 13249 5388 13283 5422
rect 13318 5388 13352 5422
rect 13387 5388 13421 5422
rect 13456 5388 13490 5422
rect 13525 5388 13559 5422
rect 13594 5388 13628 5422
rect 13663 5388 13697 5422
rect 13732 5388 13766 5422
rect 13801 5388 13835 5422
rect 13870 5388 13904 5422
rect 13939 5388 13973 5422
rect 14008 5388 14042 5422
rect 14077 5388 14111 5422
rect 14146 5388 14180 5422
rect 14215 5388 14249 5422
rect 14284 5388 14318 5422
rect 14353 5388 14387 5422
rect 14422 5388 14456 5422
rect 14491 5388 14525 5422
rect 14560 5388 14594 5422
rect 14629 5388 14663 5422
rect 14698 5388 14732 5422
rect 14767 5388 14801 5422
rect 14836 5388 14870 5422
rect 10903 5320 10937 5354
rect 10972 5320 11006 5354
rect 11041 5320 11075 5354
rect 11110 5320 11144 5354
rect 11179 5320 11213 5354
rect 11248 5320 11282 5354
rect 11317 5320 11351 5354
rect 11386 5320 11420 5354
rect 11455 5320 11489 5354
rect 11524 5320 11558 5354
rect 11593 5320 11627 5354
rect 11662 5320 11696 5354
rect 11731 5320 11765 5354
rect 11800 5320 11834 5354
rect 11869 5320 11903 5354
rect 11938 5320 11972 5354
rect 12007 5320 12041 5354
rect 12076 5320 12110 5354
rect 12145 5320 12179 5354
rect 12214 5320 12248 5354
rect 12283 5320 12317 5354
rect 12352 5320 12386 5354
rect 12421 5320 12455 5354
rect 12490 5320 12524 5354
rect 12559 5320 12593 5354
rect 12628 5320 12662 5354
rect 12697 5320 12731 5354
rect 12766 5320 12800 5354
rect 12835 5320 12869 5354
rect 12904 5320 12938 5354
rect 12973 5320 13007 5354
rect 13042 5320 13076 5354
rect 13111 5320 13145 5354
rect 13180 5320 13214 5354
rect 13249 5320 13283 5354
rect 13318 5320 13352 5354
rect 13387 5320 13421 5354
rect 13456 5320 13490 5354
rect 13525 5320 13559 5354
rect 13594 5320 13628 5354
rect 13663 5320 13697 5354
rect 13732 5320 13766 5354
rect 13801 5320 13835 5354
rect 13870 5320 13904 5354
rect 13939 5320 13973 5354
rect 14008 5320 14042 5354
rect 14077 5320 14111 5354
rect 14146 5320 14180 5354
rect 14215 5320 14249 5354
rect 14284 5320 14318 5354
rect 14353 5320 14387 5354
rect 14422 5320 14456 5354
rect 14491 5320 14525 5354
rect 14560 5320 14594 5354
rect 14629 5320 14663 5354
rect 14698 5320 14732 5354
rect 14767 5320 14801 5354
rect 14836 5320 14870 5354
rect 14935 5294 14969 5328
rect 15003 5294 15037 5328
rect 15071 5294 15105 5328
rect 10903 5252 10937 5286
rect 10972 5252 11006 5286
rect 11041 5252 11075 5286
rect 11110 5252 11144 5286
rect 11179 5252 11213 5286
rect 11248 5252 11282 5286
rect 11317 5252 11351 5286
rect 11386 5252 11420 5286
rect 11455 5252 11489 5286
rect 11524 5252 11558 5286
rect 11593 5252 11627 5286
rect 11662 5252 11696 5286
rect 11731 5252 11765 5286
rect 11800 5252 11834 5286
rect 11869 5252 11903 5286
rect 11938 5252 11972 5286
rect 12007 5252 12041 5286
rect 12076 5252 12110 5286
rect 12145 5252 12179 5286
rect 12214 5252 12248 5286
rect 12283 5252 12317 5286
rect 12352 5252 12386 5286
rect 12421 5252 12455 5286
rect 12490 5252 12524 5286
rect 12559 5252 12593 5286
rect 12628 5252 12662 5286
rect 12697 5252 12731 5286
rect 12766 5252 12800 5286
rect 12835 5252 12869 5286
rect 12904 5252 12938 5286
rect 12973 5252 13007 5286
rect 13042 5252 13076 5286
rect 13111 5252 13145 5286
rect 13180 5252 13214 5286
rect 13249 5252 13283 5286
rect 13318 5252 13352 5286
rect 13387 5252 13421 5286
rect 13456 5252 13490 5286
rect 13525 5252 13559 5286
rect 13594 5252 13628 5286
rect 13663 5252 13697 5286
rect 13732 5252 13766 5286
rect 13801 5252 13835 5286
rect 13870 5252 13904 5286
rect 13939 5252 13973 5286
rect 14008 5252 14042 5286
rect 14077 5252 14111 5286
rect 14146 5252 14180 5286
rect 14215 5252 14249 5286
rect 14284 5252 14318 5286
rect 14353 5252 14387 5286
rect 14422 5252 14456 5286
rect 14491 5252 14525 5286
rect 14560 5252 14594 5286
rect 14629 5252 14663 5286
rect 14698 5252 14732 5286
rect 14767 5252 14801 5286
rect 14836 5252 14870 5286
rect 71 5198 105 5232
rect 139 5198 173 5232
rect 207 5198 241 5232
rect 71 5127 105 5161
rect 139 5127 173 5161
rect 207 5127 241 5161
rect 71 5056 105 5090
rect 139 5056 173 5090
rect 207 5056 241 5090
rect 71 4986 105 5020
rect 139 4986 173 5020
rect 207 4986 241 5020
rect 14935 5222 14969 5256
rect 15003 5222 15037 5256
rect 15071 5222 15105 5256
rect 14935 5150 14969 5184
rect 15003 5150 15037 5184
rect 15071 5150 15105 5184
rect 14935 5078 14969 5112
rect 15003 5078 15037 5112
rect 15071 5078 15105 5112
rect 14935 5006 14969 5040
rect 15003 5006 15037 5040
rect 15071 5006 15105 5040
rect 71 4884 105 4918
rect 139 4884 173 4918
rect 207 4884 241 4918
rect 71 4815 105 4849
rect 139 4815 173 4849
rect 207 4815 241 4849
rect 71 4746 105 4780
rect 139 4746 173 4780
rect 207 4746 241 4780
rect 71 4677 105 4711
rect 139 4677 173 4711
rect 207 4677 241 4711
rect 71 4608 105 4642
rect 139 4608 173 4642
rect 207 4608 241 4642
rect 71 4539 105 4573
rect 139 4539 173 4573
rect 207 4539 241 4573
rect 71 4470 105 4504
rect 139 4470 173 4504
rect 207 4470 241 4504
rect 71 4401 105 4435
rect 139 4401 173 4435
rect 207 4401 241 4435
rect 71 4332 105 4366
rect 139 4332 173 4366
rect 207 4332 241 4366
rect 71 4263 105 4297
rect 139 4263 173 4297
rect 207 4263 241 4297
rect 71 4194 105 4228
rect 139 4194 173 4228
rect 207 4194 241 4228
rect 71 4125 105 4159
rect 139 4125 173 4159
rect 207 4125 241 4159
rect 71 4056 105 4090
rect 139 4056 173 4090
rect 207 4056 241 4090
rect 71 3987 105 4021
rect 139 3987 173 4021
rect 207 3987 241 4021
rect 71 3918 105 3952
rect 139 3918 173 3952
rect 207 3918 241 3952
rect 71 3849 105 3883
rect 139 3849 173 3883
rect 207 3849 241 3883
rect 71 3780 105 3814
rect 139 3780 173 3814
rect 207 3780 241 3814
rect 71 3711 105 3745
rect 139 3711 173 3745
rect 207 3711 241 3745
rect 71 3642 105 3676
rect 139 3642 173 3676
rect 207 3642 241 3676
rect 71 3573 105 3607
rect 139 3573 173 3607
rect 207 3573 241 3607
rect 71 3504 105 3538
rect 139 3504 173 3538
rect 207 3504 241 3538
rect 71 3435 105 3469
rect 139 3435 173 3469
rect 207 3435 241 3469
rect 71 3366 105 3400
rect 139 3366 173 3400
rect 207 3366 241 3400
rect 71 3297 105 3331
rect 139 3297 173 3331
rect 207 3297 241 3331
rect 71 3228 105 3262
rect 139 3228 173 3262
rect 207 3228 241 3262
rect 71 3159 105 3193
rect 139 3159 173 3193
rect 207 3159 241 3193
rect 71 3090 105 3124
rect 139 3090 173 3124
rect 207 3090 241 3124
rect 71 3021 105 3055
rect 139 3021 173 3055
rect 207 3021 241 3055
rect 71 2952 105 2986
rect 139 2952 173 2986
rect 207 2952 241 2986
rect 71 2883 105 2917
rect 139 2883 173 2917
rect 207 2883 241 2917
rect 71 2814 105 2848
rect 139 2814 173 2848
rect 207 2814 241 2848
rect 71 2745 105 2779
rect 139 2745 173 2779
rect 207 2745 241 2779
rect 71 2676 105 2710
rect 139 2676 173 2710
rect 207 2676 241 2710
rect 71 2607 105 2641
rect 139 2607 173 2641
rect 207 2607 241 2641
rect 71 2538 105 2572
rect 139 2538 173 2572
rect 207 2538 241 2572
rect 71 2469 105 2503
rect 139 2469 173 2503
rect 207 2469 241 2503
rect 71 2400 105 2434
rect 139 2400 173 2434
rect 207 2400 241 2434
rect 71 2331 105 2365
rect 139 2331 173 2365
rect 207 2331 241 2365
rect 71 2262 105 2296
rect 139 2262 173 2296
rect 207 2262 241 2296
rect 71 2193 105 2227
rect 139 2193 173 2227
rect 207 2193 241 2227
rect 71 2124 105 2158
rect 139 2124 173 2158
rect 207 2124 241 2158
rect 71 2055 105 2089
rect 139 2055 173 2089
rect 207 2055 241 2089
rect 71 1986 105 2020
rect 139 1986 173 2020
rect 207 1986 241 2020
rect 71 1917 105 1951
rect 139 1917 173 1951
rect 207 1917 241 1951
rect 71 1848 105 1882
rect 139 1848 173 1882
rect 207 1848 241 1882
rect 71 1779 105 1813
rect 139 1779 173 1813
rect 207 1779 241 1813
rect 71 1710 105 1744
rect 139 1710 173 1744
rect 207 1710 241 1744
rect 71 1641 105 1675
rect 139 1641 173 1675
rect 207 1641 241 1675
rect 71 1572 105 1606
rect 139 1572 173 1606
rect 207 1572 241 1606
rect 71 1503 105 1537
rect 139 1503 173 1537
rect 207 1503 241 1537
rect 71 1434 105 1468
rect 139 1434 173 1468
rect 207 1434 241 1468
rect 71 1365 105 1399
rect 139 1365 173 1399
rect 207 1365 241 1399
rect 71 1296 105 1330
rect 139 1296 173 1330
rect 207 1296 241 1330
rect 71 1227 105 1261
rect 139 1227 173 1261
rect 207 1227 241 1261
rect 71 1158 105 1192
rect 139 1158 173 1192
rect 207 1158 241 1192
rect 71 545 241 1123
rect 14935 4934 14969 4968
rect 15003 4934 15037 4968
rect 15071 4934 15105 4968
rect 14935 4862 14969 4896
rect 15003 4862 15037 4896
rect 15071 4862 15105 4896
rect 14935 4790 14969 4824
rect 15003 4790 15037 4824
rect 15071 4790 15105 4824
rect 14935 4718 14969 4752
rect 15003 4718 15037 4752
rect 15071 4718 15105 4752
rect 14935 4646 14969 4680
rect 15003 4646 15037 4680
rect 15071 4646 15105 4680
rect 14935 4574 14969 4608
rect 15003 4574 15037 4608
rect 15071 4574 15105 4608
rect 14935 4502 14969 4536
rect 15003 4502 15037 4536
rect 15071 4502 15105 4536
rect 14935 4430 14969 4464
rect 15003 4430 15037 4464
rect 15071 4430 15105 4464
rect 14935 4358 14969 4392
rect 15003 4358 15037 4392
rect 15071 4358 15105 4392
rect 14935 4286 14969 4320
rect 15003 4286 15037 4320
rect 15071 4286 15105 4320
rect 14935 4214 14969 4248
rect 15003 4214 15037 4248
rect 15071 4214 15105 4248
rect 14935 4142 14969 4176
rect 15003 4142 15037 4176
rect 15071 4142 15105 4176
rect 14935 4070 14969 4104
rect 15003 4070 15037 4104
rect 15071 4070 15105 4104
rect 14935 3998 14969 4032
rect 15003 3998 15037 4032
rect 15071 3998 15105 4032
rect 14935 3926 14969 3960
rect 15003 3926 15037 3960
rect 15071 3926 15105 3960
rect 14935 3854 14969 3888
rect 15003 3854 15037 3888
rect 15071 3854 15105 3888
rect 14935 3782 14969 3816
rect 15003 3782 15037 3816
rect 15071 3782 15105 3816
rect 14935 3710 14969 3744
rect 15003 3710 15037 3744
rect 15071 3710 15105 3744
rect 14935 3638 14969 3672
rect 15003 3638 15037 3672
rect 15071 3638 15105 3672
rect 14935 3566 14969 3600
rect 15003 3566 15037 3600
rect 15071 3566 15105 3600
rect 14935 3494 14969 3528
rect 15003 3494 15037 3528
rect 15071 3494 15105 3528
rect 14935 3422 14969 3456
rect 15003 3422 15037 3456
rect 15071 3422 15105 3456
rect 14935 3350 14969 3384
rect 15003 3350 15037 3384
rect 15071 3350 15105 3384
rect 14935 3278 14969 3312
rect 15003 3278 15037 3312
rect 15071 3278 15105 3312
rect 14935 3206 14969 3240
rect 15003 3206 15037 3240
rect 15071 3206 15105 3240
rect 14935 3134 14969 3168
rect 15003 3134 15037 3168
rect 15071 3134 15105 3168
rect 14935 3062 14969 3096
rect 15003 3062 15037 3096
rect 15071 3062 15105 3096
rect 14935 2990 14969 3024
rect 15003 2990 15037 3024
rect 15071 2990 15105 3024
rect 14935 2918 14969 2952
rect 15003 2918 15037 2952
rect 15071 2918 15105 2952
rect 14935 2846 14969 2880
rect 15003 2846 15037 2880
rect 15071 2846 15105 2880
rect 14935 2774 14969 2808
rect 15003 2774 15037 2808
rect 15071 2774 15105 2808
rect 14935 2702 14969 2736
rect 15003 2702 15037 2736
rect 15071 2702 15105 2736
rect 14935 2630 14969 2664
rect 15003 2630 15037 2664
rect 15071 2630 15105 2664
rect 14935 2558 14969 2592
rect 15003 2558 15037 2592
rect 15071 2558 15105 2592
rect 14935 2486 14969 2520
rect 15003 2486 15037 2520
rect 15071 2486 15105 2520
rect 14935 2414 14969 2448
rect 15003 2414 15037 2448
rect 15071 2414 15105 2448
rect 14935 2342 14969 2376
rect 15003 2342 15037 2376
rect 15071 2342 15105 2376
rect 14935 2270 14969 2304
rect 15003 2270 15037 2304
rect 15071 2270 15105 2304
rect 14935 2198 14969 2232
rect 15003 2198 15037 2232
rect 15071 2198 15105 2232
rect 14935 2126 14969 2160
rect 15003 2126 15037 2160
rect 15071 2126 15105 2160
rect 14935 2054 14969 2088
rect 15003 2054 15037 2088
rect 15071 2054 15105 2088
rect 14935 1982 14969 2016
rect 15003 1982 15037 2016
rect 15071 1982 15105 2016
rect 14935 1910 14969 1944
rect 15003 1910 15037 1944
rect 15071 1910 15105 1944
rect 14935 1838 14969 1872
rect 15003 1838 15037 1872
rect 15071 1838 15105 1872
rect 14935 1766 14969 1800
rect 15003 1766 15037 1800
rect 15071 1766 15105 1800
rect 14935 1694 14969 1728
rect 15003 1694 15037 1728
rect 15071 1694 15105 1728
rect 14935 1622 14969 1656
rect 15003 1622 15037 1656
rect 15071 1622 15105 1656
rect 14935 1550 14969 1584
rect 15003 1550 15037 1584
rect 15071 1550 15105 1584
rect 14935 1478 14969 1512
rect 15003 1478 15037 1512
rect 15071 1478 15105 1512
rect 14935 1406 14969 1440
rect 15003 1406 15037 1440
rect 15071 1406 15105 1440
rect 14935 1334 14969 1368
rect 15003 1334 15037 1368
rect 15071 1334 15105 1368
rect 14935 1262 14969 1296
rect 15003 1262 15037 1296
rect 15071 1262 15105 1296
rect 14935 1190 14969 1224
rect 15003 1190 15037 1224
rect 15071 1190 15105 1224
rect 14935 1118 14969 1152
rect 15003 1118 15037 1152
rect 15071 1118 15105 1152
rect 14935 1046 14969 1080
rect 15003 1046 15037 1080
rect 15071 1046 15105 1080
rect 14935 974 14969 1008
rect 15003 974 15037 1008
rect 15071 974 15105 1008
rect 14935 902 14969 936
rect 15003 902 15037 936
rect 15071 902 15105 936
rect 14935 830 14969 864
rect 15003 830 15037 864
rect 15071 830 15105 864
rect 14935 758 14969 792
rect 15003 758 15037 792
rect 15071 758 15105 792
rect 14935 686 14969 720
rect 15003 686 15037 720
rect 15071 686 15105 720
rect 294 630 328 664
rect 363 630 397 664
rect 432 630 466 664
rect 501 630 535 664
rect 570 630 604 664
rect 639 630 673 664
rect 708 630 742 664
rect 777 630 811 664
rect 846 630 880 664
rect 915 630 949 664
rect 984 630 1018 664
rect 1053 630 1087 664
rect 1122 630 1156 664
rect 1191 630 1225 664
rect 1260 630 1294 664
rect 1329 630 1363 664
rect 1398 630 1432 664
rect 1467 630 1501 664
rect 1536 630 1570 664
rect 1605 630 1639 664
rect 1674 630 1708 664
rect 1743 630 1777 664
rect 1812 630 1846 664
rect 1881 630 1915 664
rect 1950 630 1984 664
rect 2019 630 2053 664
rect 2088 630 2122 664
rect 2157 630 2191 664
rect 2226 630 2260 664
rect 2295 630 2329 664
rect 2364 630 2398 664
rect 2433 630 2467 664
rect 2502 630 2536 664
rect 2571 630 2605 664
rect 2640 630 2674 664
rect 2709 630 2743 664
rect 2778 630 2812 664
rect 2847 630 2881 664
rect 2916 630 2950 664
rect 2985 630 3019 664
rect 3054 630 3088 664
rect 3123 630 3157 664
rect 3192 630 3226 664
rect 3261 630 3295 664
rect 3330 630 3364 664
rect 3399 630 3433 664
rect 3468 630 3502 664
rect 3537 630 3571 664
rect 3606 630 3640 664
rect 3675 630 3709 664
rect 3744 630 3778 664
rect 3813 630 3847 664
rect 3882 630 3916 664
rect 3951 630 3985 664
rect 4020 630 4054 664
rect 4089 630 4123 664
rect 4158 630 4192 664
rect 4227 630 4261 664
rect 4296 630 4330 664
rect 4365 630 4399 664
rect 4434 630 4468 664
rect 4503 630 4537 664
rect 4572 630 4606 664
rect 4641 630 4675 664
rect 294 562 328 596
rect 363 562 397 596
rect 432 562 466 596
rect 501 562 535 596
rect 570 562 604 596
rect 639 562 673 596
rect 708 562 742 596
rect 777 562 811 596
rect 846 562 880 596
rect 915 562 949 596
rect 984 562 1018 596
rect 1053 562 1087 596
rect 1122 562 1156 596
rect 1191 562 1225 596
rect 1260 562 1294 596
rect 1329 562 1363 596
rect 1398 562 1432 596
rect 1467 562 1501 596
rect 1536 562 1570 596
rect 1605 562 1639 596
rect 1674 562 1708 596
rect 1743 562 1777 596
rect 1812 562 1846 596
rect 1881 562 1915 596
rect 1950 562 1984 596
rect 2019 562 2053 596
rect 2088 562 2122 596
rect 2157 562 2191 596
rect 2226 562 2260 596
rect 2295 562 2329 596
rect 2364 562 2398 596
rect 2433 562 2467 596
rect 2502 562 2536 596
rect 2571 562 2605 596
rect 2640 562 2674 596
rect 2709 562 2743 596
rect 2778 562 2812 596
rect 2847 562 2881 596
rect 2916 562 2950 596
rect 2985 562 3019 596
rect 3054 562 3088 596
rect 3123 562 3157 596
rect 3192 562 3226 596
rect 3261 562 3295 596
rect 3330 562 3364 596
rect 3399 562 3433 596
rect 3468 562 3502 596
rect 3537 562 3571 596
rect 3606 562 3640 596
rect 3675 562 3709 596
rect 3744 562 3778 596
rect 3813 562 3847 596
rect 3882 562 3916 596
rect 3951 562 3985 596
rect 4020 562 4054 596
rect 4089 562 4123 596
rect 4158 562 4192 596
rect 4227 562 4261 596
rect 4296 562 4330 596
rect 4365 562 4399 596
rect 4434 562 4468 596
rect 4503 562 4537 596
rect 4572 562 4606 596
rect 4641 562 4675 596
rect 294 494 328 528
rect 363 494 397 528
rect 432 494 466 528
rect 501 494 535 528
rect 570 494 604 528
rect 639 494 673 528
rect 708 494 742 528
rect 777 494 811 528
rect 846 494 880 528
rect 915 494 949 528
rect 984 494 1018 528
rect 1053 494 1087 528
rect 1122 494 1156 528
rect 1191 494 1225 528
rect 1260 494 1294 528
rect 1329 494 1363 528
rect 1398 494 1432 528
rect 1467 494 1501 528
rect 1536 494 1570 528
rect 1605 494 1639 528
rect 1674 494 1708 528
rect 1743 494 1777 528
rect 1812 494 1846 528
rect 1881 494 1915 528
rect 1950 494 1984 528
rect 2019 494 2053 528
rect 2088 494 2122 528
rect 2157 494 2191 528
rect 2226 494 2260 528
rect 2295 494 2329 528
rect 2364 494 2398 528
rect 2433 494 2467 528
rect 2502 494 2536 528
rect 2571 494 2605 528
rect 2640 494 2674 528
rect 2709 494 2743 528
rect 2778 494 2812 528
rect 2847 494 2881 528
rect 2916 494 2950 528
rect 2985 494 3019 528
rect 3054 494 3088 528
rect 3123 494 3157 528
rect 3192 494 3226 528
rect 3261 494 3295 528
rect 3330 494 3364 528
rect 3399 494 3433 528
rect 3468 494 3502 528
rect 3537 494 3571 528
rect 3606 494 3640 528
rect 3675 494 3709 528
rect 3744 494 3778 528
rect 3813 494 3847 528
rect 3882 494 3916 528
rect 3951 494 3985 528
rect 4020 494 4054 528
rect 4089 494 4123 528
rect 4158 494 4192 528
rect 4227 494 4261 528
rect 4296 494 4330 528
rect 4365 494 4399 528
rect 4434 494 4468 528
rect 4503 494 4537 528
rect 4572 494 4606 528
rect 4641 494 4675 528
rect 4710 494 14876 664
rect 14935 614 14969 648
rect 15003 614 15037 648
rect 15071 614 15105 648
rect 14935 542 14969 576
rect 15003 542 15037 576
rect 15071 542 15105 576
<< poly >>
rect 924 4214 1044 4230
rect 924 4180 967 4214
rect 1001 4180 1044 4214
rect 924 4140 1044 4180
rect 924 4106 967 4140
rect 1001 4106 1044 4140
rect 924 4058 1044 4106
rect 1354 4214 1474 4230
rect 1354 4180 1397 4214
rect 1431 4180 1474 4214
rect 1354 4140 1474 4180
rect 1354 4106 1397 4140
rect 1431 4106 1474 4140
rect 1354 4058 1474 4106
rect 1916 4214 2036 4230
rect 1916 4180 1959 4214
rect 1993 4180 2036 4214
rect 1916 4140 2036 4180
rect 1916 4106 1959 4140
rect 1993 4106 2036 4140
rect 1916 4058 2036 4106
rect 2346 4214 2466 4230
rect 2346 4180 2389 4214
rect 2423 4180 2466 4214
rect 2346 4140 2466 4180
rect 2346 4106 2389 4140
rect 2423 4106 2466 4140
rect 2346 4058 2466 4106
rect 2908 4214 3028 4230
rect 2908 4180 2951 4214
rect 2985 4180 3028 4214
rect 2908 4140 3028 4180
rect 2908 4106 2951 4140
rect 2985 4106 3028 4140
rect 2908 4058 3028 4106
rect 3338 4214 3458 4230
rect 3338 4180 3381 4214
rect 3415 4180 3458 4214
rect 3338 4140 3458 4180
rect 3338 4106 3381 4140
rect 3415 4106 3458 4140
rect 3338 4058 3458 4106
rect 3900 4214 4020 4230
rect 3900 4180 3943 4214
rect 3977 4180 4020 4214
rect 3900 4140 4020 4180
rect 3900 4106 3943 4140
rect 3977 4106 4020 4140
rect 3900 4058 4020 4106
rect 4330 4214 4450 4230
rect 4330 4180 4373 4214
rect 4407 4180 4450 4214
rect 4330 4140 4450 4180
rect 4330 4106 4373 4140
rect 4407 4106 4450 4140
rect 4330 4058 4450 4106
rect 4892 4214 5012 4230
rect 4892 4180 4935 4214
rect 4969 4180 5012 4214
rect 4892 4140 5012 4180
rect 4892 4106 4935 4140
rect 4969 4106 5012 4140
rect 4892 4058 5012 4106
rect 5322 4214 5442 4230
rect 5322 4180 5365 4214
rect 5399 4180 5442 4214
rect 5322 4140 5442 4180
rect 5322 4106 5365 4140
rect 5399 4106 5442 4140
rect 5322 4058 5442 4106
rect 5884 4214 6004 4230
rect 5884 4180 5927 4214
rect 5961 4180 6004 4214
rect 5884 4140 6004 4180
rect 5884 4106 5927 4140
rect 5961 4106 6004 4140
rect 5884 4058 6004 4106
rect 6314 4214 6434 4230
rect 6314 4180 6357 4214
rect 6391 4180 6434 4214
rect 6314 4140 6434 4180
rect 6314 4106 6357 4140
rect 6391 4106 6434 4140
rect 6314 4058 6434 4106
rect 6876 4214 6996 4230
rect 6876 4180 6919 4214
rect 6953 4180 6996 4214
rect 6876 4140 6996 4180
rect 6876 4106 6919 4140
rect 6953 4106 6996 4140
rect 6876 4058 6996 4106
rect 7306 4214 7426 4230
rect 7306 4180 7349 4214
rect 7383 4180 7426 4214
rect 7306 4140 7426 4180
rect 7306 4106 7349 4140
rect 7383 4106 7426 4140
rect 7306 4058 7426 4106
rect 7868 4214 7988 4230
rect 7868 4180 7911 4214
rect 7945 4180 7988 4214
rect 7868 4140 7988 4180
rect 7868 4106 7911 4140
rect 7945 4106 7988 4140
rect 7868 4058 7988 4106
rect 8298 4214 8418 4230
rect 8298 4180 8341 4214
rect 8375 4180 8418 4214
rect 8298 4140 8418 4180
rect 8298 4106 8341 4140
rect 8375 4106 8418 4140
rect 8298 4058 8418 4106
rect 8860 4214 8980 4230
rect 8860 4180 8903 4214
rect 8937 4180 8980 4214
rect 8860 4140 8980 4180
rect 8860 4106 8903 4140
rect 8937 4106 8980 4140
rect 8860 4058 8980 4106
rect 9290 4214 9410 4230
rect 9290 4180 9333 4214
rect 9367 4180 9410 4214
rect 9290 4140 9410 4180
rect 9290 4106 9333 4140
rect 9367 4106 9410 4140
rect 9290 4058 9410 4106
rect 9852 4214 9972 4230
rect 9852 4180 9895 4214
rect 9929 4180 9972 4214
rect 9852 4140 9972 4180
rect 9852 4106 9895 4140
rect 9929 4106 9972 4140
rect 9852 4058 9972 4106
rect 10282 4214 10402 4230
rect 10282 4180 10325 4214
rect 10359 4180 10402 4214
rect 10282 4140 10402 4180
rect 10282 4106 10325 4140
rect 10359 4106 10402 4140
rect 10282 4058 10402 4106
rect 10844 4214 10964 4230
rect 10844 4180 10887 4214
rect 10921 4180 10964 4214
rect 10844 4140 10964 4180
rect 10844 4106 10887 4140
rect 10921 4106 10964 4140
rect 10844 4058 10964 4106
rect 11274 4214 11394 4230
rect 11274 4180 11317 4214
rect 11351 4180 11394 4214
rect 11274 4140 11394 4180
rect 11274 4106 11317 4140
rect 11351 4106 11394 4140
rect 11274 4058 11394 4106
rect 11836 4214 11956 4230
rect 11836 4180 11879 4214
rect 11913 4180 11956 4214
rect 11836 4140 11956 4180
rect 11836 4106 11879 4140
rect 11913 4106 11956 4140
rect 11836 4058 11956 4106
rect 12266 4214 12386 4230
rect 12266 4180 12309 4214
rect 12343 4180 12386 4214
rect 12266 4140 12386 4180
rect 12266 4106 12309 4140
rect 12343 4106 12386 4140
rect 12266 4058 12386 4106
rect 12828 4214 12948 4230
rect 12828 4180 12871 4214
rect 12905 4180 12948 4214
rect 12828 4140 12948 4180
rect 12828 4106 12871 4140
rect 12905 4106 12948 4140
rect 12828 4058 12948 4106
rect 13258 4214 13378 4230
rect 13258 4180 13301 4214
rect 13335 4180 13378 4214
rect 13258 4140 13378 4180
rect 13258 4106 13301 4140
rect 13335 4106 13378 4140
rect 13258 4058 13378 4106
rect 13820 4214 13940 4230
rect 13820 4180 13863 4214
rect 13897 4180 13940 4214
rect 13820 4140 13940 4180
rect 13820 4106 13863 4140
rect 13897 4106 13940 4140
rect 13820 4058 13940 4106
rect 14178 4214 14298 4230
rect 14178 4180 14221 4214
rect 14255 4180 14298 4214
rect 14178 4140 14298 4180
rect 14178 4106 14221 4140
rect 14255 4106 14298 4140
rect 14178 4058 14298 4106
rect 924 3010 1044 3058
rect 924 2976 967 3010
rect 1001 2976 1044 3010
rect 924 2932 1044 2976
rect 924 2898 967 2932
rect 1001 2898 1044 2932
rect 924 2854 1044 2898
rect 924 2820 967 2854
rect 1001 2820 1044 2854
rect 924 2776 1044 2820
rect 924 2742 967 2776
rect 1001 2742 1044 2776
rect 924 2697 1044 2742
rect 924 2663 967 2697
rect 1001 2663 1044 2697
rect 924 2618 1044 2663
rect 924 2584 967 2618
rect 1001 2584 1044 2618
rect 924 2539 1044 2584
rect 924 2505 967 2539
rect 1001 2505 1044 2539
rect 924 2457 1044 2505
rect 1354 3010 1474 3058
rect 1354 2976 1397 3010
rect 1431 2976 1474 3010
rect 1354 2932 1474 2976
rect 1916 3010 2036 3058
rect 1916 2976 1959 3010
rect 1993 2976 2036 3010
rect 1354 2898 1397 2932
rect 1431 2898 1474 2932
rect 1354 2854 1474 2898
rect 1354 2820 1397 2854
rect 1431 2820 1474 2854
rect 1354 2776 1474 2820
rect 1354 2742 1397 2776
rect 1431 2742 1474 2776
rect 1354 2697 1474 2742
rect 1354 2663 1397 2697
rect 1431 2663 1474 2697
rect 1354 2618 1474 2663
rect 1354 2584 1397 2618
rect 1431 2584 1474 2618
rect 1354 2539 1474 2584
rect 1916 2932 2036 2976
rect 1916 2898 1959 2932
rect 1993 2898 2036 2932
rect 1916 2854 2036 2898
rect 1916 2820 1959 2854
rect 1993 2820 2036 2854
rect 1916 2776 2036 2820
rect 1916 2742 1959 2776
rect 1993 2742 2036 2776
rect 1916 2697 2036 2742
rect 1916 2663 1959 2697
rect 1993 2663 2036 2697
rect 1916 2618 2036 2663
rect 1916 2584 1959 2618
rect 1993 2584 2036 2618
rect 1354 2505 1397 2539
rect 1431 2505 1474 2539
rect 1354 2457 1474 2505
rect 1916 2539 2036 2584
rect 1916 2505 1959 2539
rect 1993 2505 2036 2539
rect 1916 2457 2036 2505
rect 2346 3010 2466 3058
rect 2346 2976 2389 3010
rect 2423 2976 2466 3010
rect 2346 2932 2466 2976
rect 2908 3010 3028 3058
rect 2908 2976 2951 3010
rect 2985 2976 3028 3010
rect 2346 2898 2389 2932
rect 2423 2898 2466 2932
rect 2346 2854 2466 2898
rect 2346 2820 2389 2854
rect 2423 2820 2466 2854
rect 2346 2776 2466 2820
rect 2346 2742 2389 2776
rect 2423 2742 2466 2776
rect 2346 2697 2466 2742
rect 2346 2663 2389 2697
rect 2423 2663 2466 2697
rect 2346 2618 2466 2663
rect 2346 2584 2389 2618
rect 2423 2584 2466 2618
rect 2346 2539 2466 2584
rect 2908 2932 3028 2976
rect 2908 2898 2951 2932
rect 2985 2898 3028 2932
rect 2908 2854 3028 2898
rect 2908 2820 2951 2854
rect 2985 2820 3028 2854
rect 2908 2776 3028 2820
rect 2908 2742 2951 2776
rect 2985 2742 3028 2776
rect 2908 2697 3028 2742
rect 2908 2663 2951 2697
rect 2985 2663 3028 2697
rect 2908 2618 3028 2663
rect 2908 2584 2951 2618
rect 2985 2584 3028 2618
rect 2346 2505 2389 2539
rect 2423 2505 2466 2539
rect 2346 2457 2466 2505
rect 2908 2539 3028 2584
rect 2908 2505 2951 2539
rect 2985 2505 3028 2539
rect 2908 2457 3028 2505
rect 3338 3010 3458 3058
rect 3338 2976 3381 3010
rect 3415 2976 3458 3010
rect 3338 2932 3458 2976
rect 3900 3010 4020 3058
rect 3900 2976 3943 3010
rect 3977 2976 4020 3010
rect 3338 2898 3381 2932
rect 3415 2898 3458 2932
rect 3338 2854 3458 2898
rect 3338 2820 3381 2854
rect 3415 2820 3458 2854
rect 3338 2776 3458 2820
rect 3338 2742 3381 2776
rect 3415 2742 3458 2776
rect 3338 2697 3458 2742
rect 3338 2663 3381 2697
rect 3415 2663 3458 2697
rect 3338 2618 3458 2663
rect 3338 2584 3381 2618
rect 3415 2584 3458 2618
rect 3338 2539 3458 2584
rect 3900 2932 4020 2976
rect 3900 2898 3943 2932
rect 3977 2898 4020 2932
rect 3900 2854 4020 2898
rect 3900 2820 3943 2854
rect 3977 2820 4020 2854
rect 3900 2776 4020 2820
rect 3900 2742 3943 2776
rect 3977 2742 4020 2776
rect 3900 2697 4020 2742
rect 3900 2663 3943 2697
rect 3977 2663 4020 2697
rect 3900 2618 4020 2663
rect 3900 2584 3943 2618
rect 3977 2584 4020 2618
rect 3338 2505 3381 2539
rect 3415 2505 3458 2539
rect 3338 2457 3458 2505
rect 3900 2539 4020 2584
rect 3900 2505 3943 2539
rect 3977 2505 4020 2539
rect 3900 2457 4020 2505
rect 4330 3010 4450 3058
rect 4330 2976 4373 3010
rect 4407 2976 4450 3010
rect 4330 2932 4450 2976
rect 4892 3010 5012 3058
rect 4892 2976 4935 3010
rect 4969 2976 5012 3010
rect 4330 2898 4373 2932
rect 4407 2898 4450 2932
rect 4330 2854 4450 2898
rect 4330 2820 4373 2854
rect 4407 2820 4450 2854
rect 4330 2776 4450 2820
rect 4330 2742 4373 2776
rect 4407 2742 4450 2776
rect 4330 2697 4450 2742
rect 4330 2663 4373 2697
rect 4407 2663 4450 2697
rect 4330 2618 4450 2663
rect 4330 2584 4373 2618
rect 4407 2584 4450 2618
rect 4330 2539 4450 2584
rect 4892 2932 5012 2976
rect 4892 2898 4935 2932
rect 4969 2898 5012 2932
rect 4892 2854 5012 2898
rect 4892 2820 4935 2854
rect 4969 2820 5012 2854
rect 4892 2776 5012 2820
rect 4892 2742 4935 2776
rect 4969 2742 5012 2776
rect 4892 2697 5012 2742
rect 4892 2663 4935 2697
rect 4969 2663 5012 2697
rect 4892 2618 5012 2663
rect 4892 2584 4935 2618
rect 4969 2584 5012 2618
rect 4330 2505 4373 2539
rect 4407 2505 4450 2539
rect 4330 2457 4450 2505
rect 4892 2539 5012 2584
rect 4892 2505 4935 2539
rect 4969 2505 5012 2539
rect 4892 2457 5012 2505
rect 5322 3010 5442 3058
rect 5322 2976 5365 3010
rect 5399 2976 5442 3010
rect 5322 2932 5442 2976
rect 5884 3010 6004 3058
rect 5884 2976 5927 3010
rect 5961 2976 6004 3010
rect 5322 2898 5365 2932
rect 5399 2898 5442 2932
rect 5322 2854 5442 2898
rect 5322 2820 5365 2854
rect 5399 2820 5442 2854
rect 5322 2776 5442 2820
rect 5322 2742 5365 2776
rect 5399 2742 5442 2776
rect 5322 2697 5442 2742
rect 5322 2663 5365 2697
rect 5399 2663 5442 2697
rect 5322 2618 5442 2663
rect 5322 2584 5365 2618
rect 5399 2584 5442 2618
rect 5322 2539 5442 2584
rect 5884 2932 6004 2976
rect 5884 2898 5927 2932
rect 5961 2898 6004 2932
rect 5884 2854 6004 2898
rect 5884 2820 5927 2854
rect 5961 2820 6004 2854
rect 5884 2776 6004 2820
rect 5884 2742 5927 2776
rect 5961 2742 6004 2776
rect 5884 2697 6004 2742
rect 5884 2663 5927 2697
rect 5961 2663 6004 2697
rect 5884 2618 6004 2663
rect 5884 2584 5927 2618
rect 5961 2584 6004 2618
rect 5322 2505 5365 2539
rect 5399 2505 5442 2539
rect 5322 2457 5442 2505
rect 5884 2539 6004 2584
rect 5884 2505 5927 2539
rect 5961 2505 6004 2539
rect 5884 2457 6004 2505
rect 6314 3010 6434 3058
rect 6314 2976 6357 3010
rect 6391 2976 6434 3010
rect 6314 2932 6434 2976
rect 6876 3010 6996 3058
rect 6876 2976 6919 3010
rect 6953 2976 6996 3010
rect 6314 2898 6357 2932
rect 6391 2898 6434 2932
rect 6314 2854 6434 2898
rect 6314 2820 6357 2854
rect 6391 2820 6434 2854
rect 6314 2776 6434 2820
rect 6314 2742 6357 2776
rect 6391 2742 6434 2776
rect 6314 2697 6434 2742
rect 6314 2663 6357 2697
rect 6391 2663 6434 2697
rect 6314 2618 6434 2663
rect 6314 2584 6357 2618
rect 6391 2584 6434 2618
rect 6314 2539 6434 2584
rect 6876 2932 6996 2976
rect 6876 2898 6919 2932
rect 6953 2898 6996 2932
rect 6876 2854 6996 2898
rect 6876 2820 6919 2854
rect 6953 2820 6996 2854
rect 6876 2776 6996 2820
rect 6876 2742 6919 2776
rect 6953 2742 6996 2776
rect 6876 2697 6996 2742
rect 6876 2663 6919 2697
rect 6953 2663 6996 2697
rect 6876 2618 6996 2663
rect 6876 2584 6919 2618
rect 6953 2584 6996 2618
rect 6314 2505 6357 2539
rect 6391 2505 6434 2539
rect 6314 2457 6434 2505
rect 6876 2539 6996 2584
rect 6876 2505 6919 2539
rect 6953 2505 6996 2539
rect 6876 2457 6996 2505
rect 7306 3010 7426 3058
rect 7306 2976 7349 3010
rect 7383 2976 7426 3010
rect 7306 2932 7426 2976
rect 7868 3010 7988 3058
rect 7868 2976 7911 3010
rect 7945 2976 7988 3010
rect 7306 2898 7349 2932
rect 7383 2898 7426 2932
rect 7306 2854 7426 2898
rect 7306 2820 7349 2854
rect 7383 2820 7426 2854
rect 7306 2776 7426 2820
rect 7306 2742 7349 2776
rect 7383 2742 7426 2776
rect 7306 2697 7426 2742
rect 7306 2663 7349 2697
rect 7383 2663 7426 2697
rect 7306 2618 7426 2663
rect 7306 2584 7349 2618
rect 7383 2584 7426 2618
rect 7306 2539 7426 2584
rect 7868 2932 7988 2976
rect 7868 2898 7911 2932
rect 7945 2898 7988 2932
rect 7868 2854 7988 2898
rect 7868 2820 7911 2854
rect 7945 2820 7988 2854
rect 7868 2776 7988 2820
rect 7868 2742 7911 2776
rect 7945 2742 7988 2776
rect 7868 2697 7988 2742
rect 7868 2663 7911 2697
rect 7945 2663 7988 2697
rect 7868 2618 7988 2663
rect 7868 2584 7911 2618
rect 7945 2584 7988 2618
rect 7306 2505 7349 2539
rect 7383 2505 7426 2539
rect 7306 2457 7426 2505
rect 7868 2539 7988 2584
rect 7868 2505 7911 2539
rect 7945 2505 7988 2539
rect 7868 2457 7988 2505
rect 8298 3010 8418 3058
rect 8298 2976 8341 3010
rect 8375 2976 8418 3010
rect 8298 2932 8418 2976
rect 8860 3010 8980 3058
rect 8860 2976 8903 3010
rect 8937 2976 8980 3010
rect 8298 2898 8341 2932
rect 8375 2898 8418 2932
rect 8298 2854 8418 2898
rect 8298 2820 8341 2854
rect 8375 2820 8418 2854
rect 8298 2776 8418 2820
rect 8298 2742 8341 2776
rect 8375 2742 8418 2776
rect 8298 2697 8418 2742
rect 8298 2663 8341 2697
rect 8375 2663 8418 2697
rect 8298 2618 8418 2663
rect 8298 2584 8341 2618
rect 8375 2584 8418 2618
rect 8298 2539 8418 2584
rect 8860 2932 8980 2976
rect 8860 2898 8903 2932
rect 8937 2898 8980 2932
rect 8860 2854 8980 2898
rect 8860 2820 8903 2854
rect 8937 2820 8980 2854
rect 8860 2776 8980 2820
rect 8860 2742 8903 2776
rect 8937 2742 8980 2776
rect 8860 2697 8980 2742
rect 8860 2663 8903 2697
rect 8937 2663 8980 2697
rect 8860 2618 8980 2663
rect 8860 2584 8903 2618
rect 8937 2584 8980 2618
rect 8298 2505 8341 2539
rect 8375 2505 8418 2539
rect 8298 2457 8418 2505
rect 8860 2539 8980 2584
rect 8860 2505 8903 2539
rect 8937 2505 8980 2539
rect 8860 2457 8980 2505
rect 9290 3010 9410 3058
rect 9290 2976 9333 3010
rect 9367 2976 9410 3010
rect 9290 2932 9410 2976
rect 9852 3010 9972 3058
rect 9852 2976 9895 3010
rect 9929 2976 9972 3010
rect 9290 2898 9333 2932
rect 9367 2898 9410 2932
rect 9290 2854 9410 2898
rect 9290 2820 9333 2854
rect 9367 2820 9410 2854
rect 9290 2776 9410 2820
rect 9290 2742 9333 2776
rect 9367 2742 9410 2776
rect 9290 2697 9410 2742
rect 9290 2663 9333 2697
rect 9367 2663 9410 2697
rect 9290 2618 9410 2663
rect 9290 2584 9333 2618
rect 9367 2584 9410 2618
rect 9290 2539 9410 2584
rect 9852 2932 9972 2976
rect 9852 2898 9895 2932
rect 9929 2898 9972 2932
rect 9852 2854 9972 2898
rect 9852 2820 9895 2854
rect 9929 2820 9972 2854
rect 9852 2776 9972 2820
rect 9852 2742 9895 2776
rect 9929 2742 9972 2776
rect 9852 2697 9972 2742
rect 9852 2663 9895 2697
rect 9929 2663 9972 2697
rect 9852 2618 9972 2663
rect 9852 2584 9895 2618
rect 9929 2584 9972 2618
rect 9290 2505 9333 2539
rect 9367 2505 9410 2539
rect 9290 2457 9410 2505
rect 9852 2539 9972 2584
rect 9852 2505 9895 2539
rect 9929 2505 9972 2539
rect 9852 2457 9972 2505
rect 10282 3010 10402 3058
rect 10282 2976 10325 3010
rect 10359 2976 10402 3010
rect 10282 2932 10402 2976
rect 10844 3010 10964 3058
rect 10844 2976 10887 3010
rect 10921 2976 10964 3010
rect 10282 2898 10325 2932
rect 10359 2898 10402 2932
rect 10282 2854 10402 2898
rect 10282 2820 10325 2854
rect 10359 2820 10402 2854
rect 10282 2776 10402 2820
rect 10282 2742 10325 2776
rect 10359 2742 10402 2776
rect 10282 2697 10402 2742
rect 10282 2663 10325 2697
rect 10359 2663 10402 2697
rect 10282 2618 10402 2663
rect 10282 2584 10325 2618
rect 10359 2584 10402 2618
rect 10282 2539 10402 2584
rect 10844 2932 10964 2976
rect 10844 2898 10887 2932
rect 10921 2898 10964 2932
rect 10844 2854 10964 2898
rect 10844 2820 10887 2854
rect 10921 2820 10964 2854
rect 10844 2776 10964 2820
rect 10844 2742 10887 2776
rect 10921 2742 10964 2776
rect 10844 2697 10964 2742
rect 10844 2663 10887 2697
rect 10921 2663 10964 2697
rect 10844 2618 10964 2663
rect 10844 2584 10887 2618
rect 10921 2584 10964 2618
rect 10282 2505 10325 2539
rect 10359 2505 10402 2539
rect 10282 2457 10402 2505
rect 10844 2539 10964 2584
rect 10844 2505 10887 2539
rect 10921 2505 10964 2539
rect 10844 2457 10964 2505
rect 11274 3010 11394 3058
rect 11274 2976 11317 3010
rect 11351 2976 11394 3010
rect 11274 2932 11394 2976
rect 11836 3010 11956 3058
rect 11836 2976 11879 3010
rect 11913 2976 11956 3010
rect 11274 2898 11317 2932
rect 11351 2898 11394 2932
rect 11274 2854 11394 2898
rect 11274 2820 11317 2854
rect 11351 2820 11394 2854
rect 11274 2776 11394 2820
rect 11274 2742 11317 2776
rect 11351 2742 11394 2776
rect 11274 2697 11394 2742
rect 11274 2663 11317 2697
rect 11351 2663 11394 2697
rect 11274 2618 11394 2663
rect 11274 2584 11317 2618
rect 11351 2584 11394 2618
rect 11274 2539 11394 2584
rect 11836 2932 11956 2976
rect 11836 2898 11879 2932
rect 11913 2898 11956 2932
rect 11836 2854 11956 2898
rect 11836 2820 11879 2854
rect 11913 2820 11956 2854
rect 11836 2776 11956 2820
rect 11836 2742 11879 2776
rect 11913 2742 11956 2776
rect 11836 2697 11956 2742
rect 11836 2663 11879 2697
rect 11913 2663 11956 2697
rect 11836 2618 11956 2663
rect 11836 2584 11879 2618
rect 11913 2584 11956 2618
rect 11274 2505 11317 2539
rect 11351 2505 11394 2539
rect 11274 2457 11394 2505
rect 11836 2539 11956 2584
rect 11836 2505 11879 2539
rect 11913 2505 11956 2539
rect 11836 2457 11956 2505
rect 12266 3010 12386 3058
rect 12266 2976 12309 3010
rect 12343 2976 12386 3010
rect 12266 2932 12386 2976
rect 12828 3010 12948 3058
rect 12828 2976 12871 3010
rect 12905 2976 12948 3010
rect 12266 2898 12309 2932
rect 12343 2898 12386 2932
rect 12266 2854 12386 2898
rect 12266 2820 12309 2854
rect 12343 2820 12386 2854
rect 12266 2776 12386 2820
rect 12266 2742 12309 2776
rect 12343 2742 12386 2776
rect 12266 2697 12386 2742
rect 12266 2663 12309 2697
rect 12343 2663 12386 2697
rect 12266 2618 12386 2663
rect 12266 2584 12309 2618
rect 12343 2584 12386 2618
rect 12266 2539 12386 2584
rect 12828 2932 12948 2976
rect 12828 2898 12871 2932
rect 12905 2898 12948 2932
rect 12828 2854 12948 2898
rect 12828 2820 12871 2854
rect 12905 2820 12948 2854
rect 12828 2776 12948 2820
rect 12828 2742 12871 2776
rect 12905 2742 12948 2776
rect 12828 2697 12948 2742
rect 12828 2663 12871 2697
rect 12905 2663 12948 2697
rect 12828 2618 12948 2663
rect 12828 2584 12871 2618
rect 12905 2584 12948 2618
rect 12266 2505 12309 2539
rect 12343 2505 12386 2539
rect 12266 2457 12386 2505
rect 12828 2539 12948 2584
rect 12828 2505 12871 2539
rect 12905 2505 12948 2539
rect 12828 2457 12948 2505
rect 13258 3010 13378 3058
rect 13258 2976 13301 3010
rect 13335 2976 13378 3010
rect 13258 2932 13378 2976
rect 13820 3010 13940 3058
rect 13820 2976 13863 3010
rect 13897 2976 13940 3010
rect 13258 2898 13301 2932
rect 13335 2898 13378 2932
rect 13258 2854 13378 2898
rect 13258 2820 13301 2854
rect 13335 2820 13378 2854
rect 13258 2776 13378 2820
rect 13258 2742 13301 2776
rect 13335 2742 13378 2776
rect 13258 2697 13378 2742
rect 13258 2663 13301 2697
rect 13335 2663 13378 2697
rect 13258 2618 13378 2663
rect 13258 2584 13301 2618
rect 13335 2584 13378 2618
rect 13258 2539 13378 2584
rect 13820 2932 13940 2976
rect 13820 2898 13863 2932
rect 13897 2898 13940 2932
rect 13820 2854 13940 2898
rect 13820 2820 13863 2854
rect 13897 2820 13940 2854
rect 13820 2776 13940 2820
rect 13820 2742 13863 2776
rect 13897 2742 13940 2776
rect 13820 2697 13940 2742
rect 13820 2663 13863 2697
rect 13897 2663 13940 2697
rect 13820 2618 13940 2663
rect 13820 2584 13863 2618
rect 13897 2584 13940 2618
rect 13258 2505 13301 2539
rect 13335 2505 13378 2539
rect 13258 2457 13378 2505
rect 13820 2539 13940 2584
rect 13820 2505 13863 2539
rect 13897 2505 13940 2539
rect 13820 2457 13940 2505
rect 14178 3010 14298 3058
rect 14178 2976 14221 3010
rect 14255 2976 14298 3010
rect 14178 2932 14298 2976
rect 14178 2898 14221 2932
rect 14255 2898 14298 2932
rect 14178 2854 14298 2898
rect 14178 2820 14221 2854
rect 14255 2820 14298 2854
rect 14178 2776 14298 2820
rect 14178 2742 14221 2776
rect 14255 2742 14298 2776
rect 14178 2697 14298 2742
rect 14178 2663 14221 2697
rect 14255 2663 14298 2697
rect 14178 2618 14298 2663
rect 14178 2584 14221 2618
rect 14255 2584 14298 2618
rect 14178 2539 14298 2584
rect 14178 2505 14221 2539
rect 14255 2505 14298 2539
rect 14178 2457 14298 2505
rect 924 1409 1044 1457
rect 924 1375 967 1409
rect 1001 1375 1044 1409
rect 924 1335 1044 1375
rect 924 1301 967 1335
rect 1001 1301 1044 1335
rect 924 1285 1044 1301
rect 1354 1409 1474 1457
rect 1354 1375 1397 1409
rect 1431 1375 1474 1409
rect 1354 1335 1474 1375
rect 1354 1301 1397 1335
rect 1431 1301 1474 1335
rect 1354 1285 1474 1301
rect 1916 1409 2036 1457
rect 1916 1375 1959 1409
rect 1993 1375 2036 1409
rect 1916 1335 2036 1375
rect 1916 1301 1959 1335
rect 1993 1301 2036 1335
rect 1916 1285 2036 1301
rect 2346 1409 2466 1457
rect 2346 1375 2389 1409
rect 2423 1375 2466 1409
rect 2346 1335 2466 1375
rect 2346 1301 2389 1335
rect 2423 1301 2466 1335
rect 2346 1285 2466 1301
rect 2908 1409 3028 1457
rect 2908 1375 2951 1409
rect 2985 1375 3028 1409
rect 2908 1335 3028 1375
rect 2908 1301 2951 1335
rect 2985 1301 3028 1335
rect 2908 1285 3028 1301
rect 3338 1409 3458 1457
rect 3338 1375 3381 1409
rect 3415 1375 3458 1409
rect 3338 1335 3458 1375
rect 3338 1301 3381 1335
rect 3415 1301 3458 1335
rect 3338 1285 3458 1301
rect 3900 1409 4020 1457
rect 3900 1375 3943 1409
rect 3977 1375 4020 1409
rect 3900 1335 4020 1375
rect 3900 1301 3943 1335
rect 3977 1301 4020 1335
rect 3900 1285 4020 1301
rect 4330 1409 4450 1457
rect 4330 1375 4373 1409
rect 4407 1375 4450 1409
rect 4330 1335 4450 1375
rect 4330 1301 4373 1335
rect 4407 1301 4450 1335
rect 4330 1285 4450 1301
rect 4892 1409 5012 1457
rect 4892 1375 4935 1409
rect 4969 1375 5012 1409
rect 4892 1335 5012 1375
rect 4892 1301 4935 1335
rect 4969 1301 5012 1335
rect 4892 1285 5012 1301
rect 5322 1409 5442 1457
rect 5322 1375 5365 1409
rect 5399 1375 5442 1409
rect 5322 1335 5442 1375
rect 5322 1301 5365 1335
rect 5399 1301 5442 1335
rect 5322 1285 5442 1301
rect 5884 1409 6004 1457
rect 5884 1375 5927 1409
rect 5961 1375 6004 1409
rect 5884 1335 6004 1375
rect 5884 1301 5927 1335
rect 5961 1301 6004 1335
rect 5884 1285 6004 1301
rect 6314 1409 6434 1457
rect 6314 1375 6357 1409
rect 6391 1375 6434 1409
rect 6314 1335 6434 1375
rect 6314 1301 6357 1335
rect 6391 1301 6434 1335
rect 6314 1285 6434 1301
rect 6876 1409 6996 1457
rect 6876 1375 6919 1409
rect 6953 1375 6996 1409
rect 6876 1335 6996 1375
rect 6876 1301 6919 1335
rect 6953 1301 6996 1335
rect 6876 1285 6996 1301
rect 7306 1409 7426 1457
rect 7306 1375 7349 1409
rect 7383 1375 7426 1409
rect 7306 1335 7426 1375
rect 7306 1301 7349 1335
rect 7383 1301 7426 1335
rect 7306 1285 7426 1301
rect 7868 1409 7988 1457
rect 7868 1375 7911 1409
rect 7945 1375 7988 1409
rect 7868 1335 7988 1375
rect 7868 1301 7911 1335
rect 7945 1301 7988 1335
rect 7868 1285 7988 1301
rect 8298 1409 8418 1457
rect 8298 1375 8341 1409
rect 8375 1375 8418 1409
rect 8298 1335 8418 1375
rect 8298 1301 8341 1335
rect 8375 1301 8418 1335
rect 8298 1285 8418 1301
rect 8860 1409 8980 1457
rect 8860 1375 8903 1409
rect 8937 1375 8980 1409
rect 8860 1335 8980 1375
rect 8860 1301 8903 1335
rect 8937 1301 8980 1335
rect 8860 1285 8980 1301
rect 9290 1409 9410 1457
rect 9290 1375 9333 1409
rect 9367 1375 9410 1409
rect 9290 1335 9410 1375
rect 9290 1301 9333 1335
rect 9367 1301 9410 1335
rect 9290 1285 9410 1301
rect 9852 1409 9972 1457
rect 9852 1375 9895 1409
rect 9929 1375 9972 1409
rect 9852 1335 9972 1375
rect 9852 1301 9895 1335
rect 9929 1301 9972 1335
rect 9852 1285 9972 1301
rect 10282 1409 10402 1457
rect 10282 1375 10325 1409
rect 10359 1375 10402 1409
rect 10282 1335 10402 1375
rect 10282 1301 10325 1335
rect 10359 1301 10402 1335
rect 10282 1285 10402 1301
rect 10844 1409 10964 1457
rect 10844 1375 10887 1409
rect 10921 1375 10964 1409
rect 10844 1335 10964 1375
rect 10844 1301 10887 1335
rect 10921 1301 10964 1335
rect 10844 1285 10964 1301
rect 11274 1409 11394 1457
rect 11274 1375 11317 1409
rect 11351 1375 11394 1409
rect 11274 1335 11394 1375
rect 11274 1301 11317 1335
rect 11351 1301 11394 1335
rect 11274 1285 11394 1301
rect 11836 1409 11956 1457
rect 11836 1375 11879 1409
rect 11913 1375 11956 1409
rect 11836 1335 11956 1375
rect 11836 1301 11879 1335
rect 11913 1301 11956 1335
rect 11836 1285 11956 1301
rect 12266 1409 12386 1457
rect 12266 1375 12309 1409
rect 12343 1375 12386 1409
rect 12266 1335 12386 1375
rect 12266 1301 12309 1335
rect 12343 1301 12386 1335
rect 12266 1285 12386 1301
rect 12828 1409 12948 1457
rect 12828 1375 12871 1409
rect 12905 1375 12948 1409
rect 12828 1335 12948 1375
rect 12828 1301 12871 1335
rect 12905 1301 12948 1335
rect 12828 1285 12948 1301
rect 13258 1409 13378 1457
rect 13258 1375 13301 1409
rect 13335 1375 13378 1409
rect 13258 1335 13378 1375
rect 13258 1301 13301 1335
rect 13335 1301 13378 1335
rect 13258 1285 13378 1301
rect 13820 1409 13940 1457
rect 13820 1375 13863 1409
rect 13897 1375 13940 1409
rect 13820 1335 13940 1375
rect 13820 1301 13863 1335
rect 13897 1301 13940 1335
rect 13820 1285 13940 1301
rect 14178 1409 14298 1457
rect 14178 1375 14221 1409
rect 14255 1375 14298 1409
rect 14178 1335 14298 1375
rect 14178 1301 14221 1335
rect 14255 1301 14298 1335
rect 14178 1285 14298 1301
<< polycont >>
rect 967 4180 1001 4214
rect 967 4106 1001 4140
rect 1397 4180 1431 4214
rect 1397 4106 1431 4140
rect 1959 4180 1993 4214
rect 1959 4106 1993 4140
rect 2389 4180 2423 4214
rect 2389 4106 2423 4140
rect 2951 4180 2985 4214
rect 2951 4106 2985 4140
rect 3381 4180 3415 4214
rect 3381 4106 3415 4140
rect 3943 4180 3977 4214
rect 3943 4106 3977 4140
rect 4373 4180 4407 4214
rect 4373 4106 4407 4140
rect 4935 4180 4969 4214
rect 4935 4106 4969 4140
rect 5365 4180 5399 4214
rect 5365 4106 5399 4140
rect 5927 4180 5961 4214
rect 5927 4106 5961 4140
rect 6357 4180 6391 4214
rect 6357 4106 6391 4140
rect 6919 4180 6953 4214
rect 6919 4106 6953 4140
rect 7349 4180 7383 4214
rect 7349 4106 7383 4140
rect 7911 4180 7945 4214
rect 7911 4106 7945 4140
rect 8341 4180 8375 4214
rect 8341 4106 8375 4140
rect 8903 4180 8937 4214
rect 8903 4106 8937 4140
rect 9333 4180 9367 4214
rect 9333 4106 9367 4140
rect 9895 4180 9929 4214
rect 9895 4106 9929 4140
rect 10325 4180 10359 4214
rect 10325 4106 10359 4140
rect 10887 4180 10921 4214
rect 10887 4106 10921 4140
rect 11317 4180 11351 4214
rect 11317 4106 11351 4140
rect 11879 4180 11913 4214
rect 11879 4106 11913 4140
rect 12309 4180 12343 4214
rect 12309 4106 12343 4140
rect 12871 4180 12905 4214
rect 12871 4106 12905 4140
rect 13301 4180 13335 4214
rect 13301 4106 13335 4140
rect 13863 4180 13897 4214
rect 13863 4106 13897 4140
rect 14221 4180 14255 4214
rect 14221 4106 14255 4140
rect 967 2976 1001 3010
rect 967 2898 1001 2932
rect 967 2820 1001 2854
rect 967 2742 1001 2776
rect 967 2663 1001 2697
rect 967 2584 1001 2618
rect 967 2505 1001 2539
rect 1397 2976 1431 3010
rect 1959 2976 1993 3010
rect 1397 2898 1431 2932
rect 1397 2820 1431 2854
rect 1397 2742 1431 2776
rect 1397 2663 1431 2697
rect 1397 2584 1431 2618
rect 1959 2898 1993 2932
rect 1959 2820 1993 2854
rect 1959 2742 1993 2776
rect 1959 2663 1993 2697
rect 1959 2584 1993 2618
rect 1397 2505 1431 2539
rect 1959 2505 1993 2539
rect 2389 2976 2423 3010
rect 2951 2976 2985 3010
rect 2389 2898 2423 2932
rect 2389 2820 2423 2854
rect 2389 2742 2423 2776
rect 2389 2663 2423 2697
rect 2389 2584 2423 2618
rect 2951 2898 2985 2932
rect 2951 2820 2985 2854
rect 2951 2742 2985 2776
rect 2951 2663 2985 2697
rect 2951 2584 2985 2618
rect 2389 2505 2423 2539
rect 2951 2505 2985 2539
rect 3381 2976 3415 3010
rect 3943 2976 3977 3010
rect 3381 2898 3415 2932
rect 3381 2820 3415 2854
rect 3381 2742 3415 2776
rect 3381 2663 3415 2697
rect 3381 2584 3415 2618
rect 3943 2898 3977 2932
rect 3943 2820 3977 2854
rect 3943 2742 3977 2776
rect 3943 2663 3977 2697
rect 3943 2584 3977 2618
rect 3381 2505 3415 2539
rect 3943 2505 3977 2539
rect 4373 2976 4407 3010
rect 4935 2976 4969 3010
rect 4373 2898 4407 2932
rect 4373 2820 4407 2854
rect 4373 2742 4407 2776
rect 4373 2663 4407 2697
rect 4373 2584 4407 2618
rect 4935 2898 4969 2932
rect 4935 2820 4969 2854
rect 4935 2742 4969 2776
rect 4935 2663 4969 2697
rect 4935 2584 4969 2618
rect 4373 2505 4407 2539
rect 4935 2505 4969 2539
rect 5365 2976 5399 3010
rect 5927 2976 5961 3010
rect 5365 2898 5399 2932
rect 5365 2820 5399 2854
rect 5365 2742 5399 2776
rect 5365 2663 5399 2697
rect 5365 2584 5399 2618
rect 5927 2898 5961 2932
rect 5927 2820 5961 2854
rect 5927 2742 5961 2776
rect 5927 2663 5961 2697
rect 5927 2584 5961 2618
rect 5365 2505 5399 2539
rect 5927 2505 5961 2539
rect 6357 2976 6391 3010
rect 6919 2976 6953 3010
rect 6357 2898 6391 2932
rect 6357 2820 6391 2854
rect 6357 2742 6391 2776
rect 6357 2663 6391 2697
rect 6357 2584 6391 2618
rect 6919 2898 6953 2932
rect 6919 2820 6953 2854
rect 6919 2742 6953 2776
rect 6919 2663 6953 2697
rect 6919 2584 6953 2618
rect 6357 2505 6391 2539
rect 6919 2505 6953 2539
rect 7349 2976 7383 3010
rect 7911 2976 7945 3010
rect 7349 2898 7383 2932
rect 7349 2820 7383 2854
rect 7349 2742 7383 2776
rect 7349 2663 7383 2697
rect 7349 2584 7383 2618
rect 7911 2898 7945 2932
rect 7911 2820 7945 2854
rect 7911 2742 7945 2776
rect 7911 2663 7945 2697
rect 7911 2584 7945 2618
rect 7349 2505 7383 2539
rect 7911 2505 7945 2539
rect 8341 2976 8375 3010
rect 8903 2976 8937 3010
rect 8341 2898 8375 2932
rect 8341 2820 8375 2854
rect 8341 2742 8375 2776
rect 8341 2663 8375 2697
rect 8341 2584 8375 2618
rect 8903 2898 8937 2932
rect 8903 2820 8937 2854
rect 8903 2742 8937 2776
rect 8903 2663 8937 2697
rect 8903 2584 8937 2618
rect 8341 2505 8375 2539
rect 8903 2505 8937 2539
rect 9333 2976 9367 3010
rect 9895 2976 9929 3010
rect 9333 2898 9367 2932
rect 9333 2820 9367 2854
rect 9333 2742 9367 2776
rect 9333 2663 9367 2697
rect 9333 2584 9367 2618
rect 9895 2898 9929 2932
rect 9895 2820 9929 2854
rect 9895 2742 9929 2776
rect 9895 2663 9929 2697
rect 9895 2584 9929 2618
rect 9333 2505 9367 2539
rect 9895 2505 9929 2539
rect 10325 2976 10359 3010
rect 10887 2976 10921 3010
rect 10325 2898 10359 2932
rect 10325 2820 10359 2854
rect 10325 2742 10359 2776
rect 10325 2663 10359 2697
rect 10325 2584 10359 2618
rect 10887 2898 10921 2932
rect 10887 2820 10921 2854
rect 10887 2742 10921 2776
rect 10887 2663 10921 2697
rect 10887 2584 10921 2618
rect 10325 2505 10359 2539
rect 10887 2505 10921 2539
rect 11317 2976 11351 3010
rect 11879 2976 11913 3010
rect 11317 2898 11351 2932
rect 11317 2820 11351 2854
rect 11317 2742 11351 2776
rect 11317 2663 11351 2697
rect 11317 2584 11351 2618
rect 11879 2898 11913 2932
rect 11879 2820 11913 2854
rect 11879 2742 11913 2776
rect 11879 2663 11913 2697
rect 11879 2584 11913 2618
rect 11317 2505 11351 2539
rect 11879 2505 11913 2539
rect 12309 2976 12343 3010
rect 12871 2976 12905 3010
rect 12309 2898 12343 2932
rect 12309 2820 12343 2854
rect 12309 2742 12343 2776
rect 12309 2663 12343 2697
rect 12309 2584 12343 2618
rect 12871 2898 12905 2932
rect 12871 2820 12905 2854
rect 12871 2742 12905 2776
rect 12871 2663 12905 2697
rect 12871 2584 12905 2618
rect 12309 2505 12343 2539
rect 12871 2505 12905 2539
rect 13301 2976 13335 3010
rect 13863 2976 13897 3010
rect 13301 2898 13335 2932
rect 13301 2820 13335 2854
rect 13301 2742 13335 2776
rect 13301 2663 13335 2697
rect 13301 2584 13335 2618
rect 13863 2898 13897 2932
rect 13863 2820 13897 2854
rect 13863 2742 13897 2776
rect 13863 2663 13897 2697
rect 13863 2584 13897 2618
rect 13301 2505 13335 2539
rect 13863 2505 13897 2539
rect 14221 2976 14255 3010
rect 14221 2898 14255 2932
rect 14221 2820 14255 2854
rect 14221 2742 14255 2776
rect 14221 2663 14255 2697
rect 14221 2584 14255 2618
rect 14221 2505 14255 2539
rect 967 1375 1001 1409
rect 967 1301 1001 1335
rect 1397 1375 1431 1409
rect 1397 1301 1431 1335
rect 1959 1375 1993 1409
rect 1959 1301 1993 1335
rect 2389 1375 2423 1409
rect 2389 1301 2423 1335
rect 2951 1375 2985 1409
rect 2951 1301 2985 1335
rect 3381 1375 3415 1409
rect 3381 1301 3415 1335
rect 3943 1375 3977 1409
rect 3943 1301 3977 1335
rect 4373 1375 4407 1409
rect 4373 1301 4407 1335
rect 4935 1375 4969 1409
rect 4935 1301 4969 1335
rect 5365 1375 5399 1409
rect 5365 1301 5399 1335
rect 5927 1375 5961 1409
rect 5927 1301 5961 1335
rect 6357 1375 6391 1409
rect 6357 1301 6391 1335
rect 6919 1375 6953 1409
rect 6919 1301 6953 1335
rect 7349 1375 7383 1409
rect 7349 1301 7383 1335
rect 7911 1375 7945 1409
rect 7911 1301 7945 1335
rect 8341 1375 8375 1409
rect 8341 1301 8375 1335
rect 8903 1375 8937 1409
rect 8903 1301 8937 1335
rect 9333 1375 9367 1409
rect 9333 1301 9367 1335
rect 9895 1375 9929 1409
rect 9895 1301 9929 1335
rect 10325 1375 10359 1409
rect 10325 1301 10359 1335
rect 10887 1375 10921 1409
rect 10887 1301 10921 1335
rect 11317 1375 11351 1409
rect 11317 1301 11351 1335
rect 11879 1375 11913 1409
rect 11879 1301 11913 1335
rect 12309 1375 12343 1409
rect 12309 1301 12343 1335
rect 12871 1375 12905 1409
rect 12871 1301 12905 1335
rect 13301 1375 13335 1409
rect 13301 1301 13335 1335
rect 13863 1375 13897 1409
rect 13863 1301 13897 1335
rect 14221 1375 14255 1409
rect 14221 1301 14255 1335
<< locali >>
rect 67 496 71 5426
rect 249 5422 308 5426
rect 249 5252 294 5422
rect 14886 5420 15106 5426
rect 249 5248 308 5252
rect 14886 5248 14927 5420
rect 555 4922 657 4956
rect 589 4888 657 4922
rect 555 4854 623 4888
rect 555 4850 691 4854
rect 589 4819 691 4850
rect 589 4816 623 4819
rect 555 4785 623 4816
rect 657 4786 691 4819
rect 14495 4922 14530 4956
rect 14564 4922 14599 4956
rect 14633 4922 14667 4956
rect 14461 4888 14667 4922
rect 14461 4854 14496 4888
rect 14530 4854 14565 4888
rect 14599 4854 14667 4888
rect 14393 4852 14667 4854
rect 14393 4818 14402 4852
rect 14436 4844 14667 4852
rect 14436 4820 14633 4844
rect 14393 4786 14428 4818
rect 14462 4786 14497 4820
rect 14531 4818 14633 4820
rect 14531 4786 14565 4818
rect 657 4785 822 4786
rect 555 4778 822 4785
rect 589 4774 822 4778
rect 589 4751 733 4774
rect 589 4750 691 4751
rect 589 4744 623 4750
rect 555 4710 587 4744
rect 621 4716 623 4744
rect 657 4744 691 4750
rect 657 4716 659 4744
rect 725 4740 733 4751
rect 767 4740 822 4774
rect 725 4717 822 4740
rect 621 4710 659 4716
rect 693 4710 822 4717
rect 555 4706 822 4710
rect 589 4701 822 4706
rect 589 4682 733 4701
rect 589 4681 691 4682
rect 589 4672 623 4681
rect 555 4670 623 4672
rect 555 4636 587 4670
rect 621 4647 623 4670
rect 657 4670 691 4681
rect 657 4647 659 4670
rect 725 4667 733 4682
rect 767 4667 822 4701
rect 725 4648 822 4667
rect 621 4636 659 4647
rect 693 4636 822 4648
rect 555 4634 822 4636
rect 589 4628 822 4634
rect 589 4613 733 4628
rect 589 4600 623 4613
rect 555 4596 623 4600
rect 555 4563 587 4596
rect 621 4562 623 4596
rect 725 4594 733 4613
rect 767 4594 822 4628
rect 589 4529 623 4562
rect 555 4522 623 4529
rect 725 4555 822 4594
rect 555 4492 587 4522
rect 621 4488 623 4522
rect 725 4521 733 4555
rect 767 4521 822 4555
rect 589 4458 623 4488
rect 555 4449 623 4458
rect 725 4482 822 4521
rect 14400 4784 14565 4786
rect 14599 4810 14633 4818
rect 14599 4784 14667 4810
rect 14400 4774 14667 4784
rect 14400 4740 14431 4774
rect 14465 4771 14667 4774
rect 14465 4750 14633 4771
rect 14465 4740 14497 4750
rect 14531 4748 14633 4750
rect 14531 4743 14565 4748
rect 14599 4743 14633 4748
rect 14400 4716 14497 4740
rect 14400 4709 14510 4716
rect 14544 4714 14565 4743
rect 14616 4737 14633 4743
rect 14544 4709 14582 4714
rect 14616 4709 14667 4737
rect 14400 4701 14667 4709
rect 14400 4667 14431 4701
rect 14465 4698 14667 4701
rect 14465 4680 14633 4698
rect 14465 4667 14497 4680
rect 14531 4678 14633 4680
rect 14531 4670 14565 4678
rect 14599 4670 14633 4678
rect 14400 4646 14497 4667
rect 14400 4636 14510 4646
rect 14544 4644 14565 4670
rect 14616 4664 14633 4670
rect 14544 4636 14582 4644
rect 14616 4636 14667 4664
rect 14400 4628 14667 4636
rect 14400 4594 14431 4628
rect 14465 4625 14667 4628
rect 14465 4610 14633 4625
rect 14465 4594 14497 4610
rect 14531 4608 14633 4610
rect 14531 4597 14565 4608
rect 14599 4597 14633 4608
rect 14400 4576 14497 4594
rect 14400 4563 14510 4576
rect 14544 4574 14565 4597
rect 14616 4591 14633 4597
rect 14544 4563 14582 4574
rect 14616 4563 14667 4591
rect 14400 4555 14667 4563
rect 14400 4521 14431 4555
rect 14465 4552 14667 4555
rect 14465 4540 14633 4552
rect 14465 4521 14497 4540
rect 14531 4538 14633 4540
rect 14531 4524 14565 4538
rect 14599 4524 14633 4538
rect 14400 4506 14497 4521
rect 555 4421 587 4449
rect 621 4415 623 4449
rect 725 4448 733 4482
rect 767 4448 822 4482
rect 589 4387 623 4415
rect 555 4376 623 4387
rect 725 4409 822 4448
rect 555 4350 587 4376
rect 621 4342 623 4376
rect 725 4375 733 4409
rect 767 4375 822 4409
rect 589 4316 623 4342
rect 555 4303 623 4316
rect 725 4336 822 4375
rect 555 4279 587 4303
rect 621 4269 623 4303
rect 725 4302 733 4336
rect 767 4302 822 4336
rect 589 4245 623 4269
rect 555 4230 623 4245
rect 725 4263 822 4302
rect 555 4208 587 4230
rect 621 4196 623 4230
rect 725 4229 733 4263
rect 767 4229 822 4263
rect 589 4174 623 4196
rect 555 4157 623 4174
rect 725 4190 822 4229
rect 555 4137 587 4157
rect 621 4123 623 4157
rect 725 4156 733 4190
rect 767 4156 822 4190
rect 589 4103 623 4123
rect 725 4117 822 4156
rect 725 4103 733 4117
rect 555 4084 733 4103
rect 555 4050 587 4084
rect 621 4050 659 4084
rect 693 4083 733 4084
rect 767 4083 822 4117
rect 693 4062 822 4083
rect 924 4388 931 4494
rect 1037 4388 1044 4494
rect 924 4214 1044 4388
rect 924 4180 967 4214
rect 1001 4180 1044 4214
rect 924 4140 1044 4180
rect 924 4106 967 4140
rect 1001 4106 1044 4140
rect 693 4050 836 4062
rect 555 4046 836 4050
rect 555 4044 802 4046
rect 555 4041 733 4044
rect 589 4011 623 4041
rect 621 4007 623 4011
rect 657 4011 733 4041
rect 767 4034 802 4044
rect 657 4007 659 4011
rect 555 3977 587 4007
rect 621 3977 659 4007
rect 693 4010 733 4011
rect 768 4012 802 4034
rect 693 4000 734 4010
rect 768 4000 836 4012
rect 693 3978 836 4000
rect 693 3977 802 3978
rect 555 3971 802 3977
rect 555 3970 733 3971
rect 589 3938 623 3970
rect 621 3936 623 3938
rect 657 3938 733 3970
rect 767 3966 802 3971
rect 657 3936 659 3938
rect 555 3904 587 3936
rect 621 3904 659 3936
rect 693 3937 733 3938
rect 768 3944 802 3966
rect 693 3932 734 3937
rect 768 3932 836 3944
rect 693 3910 836 3932
rect 693 3904 802 3910
rect 555 3898 802 3904
rect 555 3896 733 3898
rect 589 3865 623 3896
rect 621 3862 623 3865
rect 657 3865 733 3896
rect 657 3862 659 3865
rect 555 3831 587 3862
rect 621 3831 659 3862
rect 693 3864 733 3865
rect 768 3876 802 3898
rect 768 3864 836 3876
rect 693 3842 836 3864
rect 693 3831 802 3842
rect 555 3830 802 3831
rect 555 3825 734 3830
rect 589 3792 623 3825
rect 621 3791 623 3792
rect 657 3792 733 3825
rect 768 3808 802 3830
rect 768 3796 836 3808
rect 657 3791 659 3792
rect 555 3758 587 3791
rect 621 3758 659 3791
rect 693 3791 733 3792
rect 767 3791 836 3796
rect 693 3774 836 3791
rect 693 3762 802 3774
rect 693 3758 734 3762
rect 555 3752 734 3758
rect 555 3751 733 3752
rect 589 3719 623 3751
rect 621 3717 623 3719
rect 657 3719 733 3751
rect 768 3740 802 3762
rect 768 3728 836 3740
rect 657 3717 659 3719
rect 555 3685 587 3717
rect 621 3685 659 3717
rect 693 3718 733 3719
rect 767 3718 836 3728
rect 693 3706 836 3718
rect 693 3694 802 3706
rect 693 3685 734 3694
rect 555 3680 734 3685
rect 589 3646 623 3680
rect 657 3679 734 3680
rect 657 3646 733 3679
rect 768 3672 802 3694
rect 768 3660 836 3672
rect 555 3612 587 3646
rect 621 3612 659 3646
rect 693 3645 733 3646
rect 767 3645 836 3660
rect 693 3638 836 3645
rect 693 3626 802 3638
rect 693 3612 734 3626
rect 555 3606 734 3612
rect 589 3573 623 3606
rect 621 3572 623 3573
rect 657 3573 733 3606
rect 768 3604 802 3626
rect 768 3592 836 3604
rect 657 3572 659 3573
rect 555 3539 587 3572
rect 621 3539 659 3572
rect 693 3572 733 3573
rect 767 3572 836 3592
rect 693 3570 836 3572
rect 693 3558 802 3570
rect 693 3539 734 3558
rect 555 3535 734 3539
rect 589 3501 623 3535
rect 657 3533 734 3535
rect 768 3536 802 3558
rect 657 3501 733 3533
rect 768 3524 836 3536
rect 555 3500 733 3501
rect 555 3466 587 3500
rect 621 3466 659 3500
rect 693 3499 733 3500
rect 767 3502 836 3524
rect 767 3499 802 3502
rect 693 3490 802 3499
rect 693 3466 734 3490
rect 555 3461 734 3466
rect 589 3427 623 3461
rect 657 3460 734 3461
rect 768 3468 802 3490
rect 657 3427 733 3460
rect 768 3456 836 3468
rect 555 3393 587 3427
rect 621 3393 659 3427
rect 693 3426 733 3427
rect 767 3434 836 3456
rect 767 3426 802 3434
rect 693 3422 802 3426
rect 693 3393 734 3422
rect 555 3390 734 3393
rect 589 3356 623 3390
rect 657 3388 734 3390
rect 768 3400 802 3422
rect 768 3388 836 3400
rect 657 3387 836 3388
rect 657 3356 733 3387
rect 555 3354 733 3356
rect 767 3366 836 3387
rect 767 3354 802 3366
rect 555 3320 587 3354
rect 621 3320 659 3354
rect 693 3353 733 3354
rect 693 3320 734 3353
rect 768 3332 802 3354
rect 768 3320 836 3332
rect 555 3316 836 3320
rect 589 3282 623 3316
rect 657 3314 836 3316
rect 657 3282 733 3314
rect 767 3298 836 3314
rect 767 3286 802 3298
rect 555 3281 733 3282
rect 555 3247 587 3281
rect 621 3247 659 3281
rect 693 3280 733 3281
rect 693 3252 734 3280
rect 768 3264 802 3286
rect 768 3252 836 3264
rect 693 3247 836 3252
rect 555 3245 836 3247
rect 589 3211 623 3245
rect 657 3241 836 3245
rect 657 3211 733 3241
rect 767 3230 836 3241
rect 767 3218 802 3230
rect 555 3208 733 3211
rect 555 3174 587 3208
rect 621 3174 659 3208
rect 693 3207 733 3208
rect 693 3184 734 3207
rect 768 3196 802 3218
rect 768 3184 836 3196
rect 693 3174 836 3184
rect 555 3168 836 3174
rect 555 3151 733 3168
rect 589 3135 623 3151
rect 621 3117 623 3135
rect 657 3135 733 3151
rect 767 3162 836 3168
rect 767 3150 802 3162
rect 657 3117 659 3135
rect 555 3101 587 3117
rect 621 3101 659 3117
rect 693 3134 733 3135
rect 693 3116 734 3134
rect 768 3128 802 3150
rect 768 3116 836 3128
rect 693 3101 836 3116
rect 555 3100 836 3101
rect 555 3095 822 3100
rect 555 3081 733 3095
rect 657 3062 733 3081
rect 657 3028 659 3062
rect 693 3061 733 3062
rect 767 3061 822 3095
rect 693 3028 822 3061
rect 657 3022 822 3028
rect 657 3013 733 3022
rect 725 2988 733 3013
rect 767 2988 822 3022
rect 725 2949 822 2988
rect 725 2915 733 2949
rect 767 2915 822 2949
rect 725 2876 822 2915
rect 725 2842 733 2876
rect 767 2842 822 2876
rect 725 2803 822 2842
rect 725 2769 733 2803
rect 767 2769 822 2803
rect 725 2730 822 2769
rect 725 2696 733 2730
rect 767 2696 822 2730
rect 725 2657 822 2696
rect 725 2623 733 2657
rect 767 2623 822 2657
rect 725 2584 822 2623
rect 725 2550 733 2584
rect 767 2550 822 2584
rect 725 2511 822 2550
rect 725 2503 733 2511
rect 657 2478 733 2503
rect 657 2444 659 2478
rect 693 2477 733 2478
rect 767 2477 822 2511
rect 693 2461 822 2477
rect 924 3010 1044 4106
rect 1354 4388 1361 4494
rect 1467 4388 1474 4494
rect 1354 4214 1474 4388
rect 1354 4180 1397 4214
rect 1431 4180 1474 4214
rect 1354 4140 1474 4180
rect 1354 4106 1397 4140
rect 1431 4106 1474 4140
rect 924 2976 967 3010
rect 1001 2976 1044 3010
rect 924 2932 1044 2976
rect 924 2898 967 2932
rect 1001 2898 1044 2932
rect 924 2854 1044 2898
rect 924 2820 967 2854
rect 1001 2820 1044 2854
rect 924 2776 1044 2820
rect 924 2742 967 2776
rect 1001 2742 1044 2776
rect 924 2697 1044 2742
rect 924 2663 967 2697
rect 1001 2663 1044 2697
rect 924 2618 1044 2663
rect 924 2584 967 2618
rect 1001 2584 1044 2618
rect 924 2539 1044 2584
rect 924 2505 967 2539
rect 1001 2505 1044 2539
rect 693 2445 836 2461
rect 693 2444 802 2445
rect 657 2438 802 2444
rect 657 2405 733 2438
rect 767 2433 802 2438
rect 657 2371 659 2405
rect 693 2404 733 2405
rect 768 2411 802 2433
rect 693 2399 734 2404
rect 768 2399 836 2411
rect 693 2377 836 2399
rect 693 2371 802 2377
rect 657 2367 802 2371
rect 555 2365 802 2367
rect 555 2332 733 2365
rect 555 2327 587 2332
rect 621 2327 659 2332
rect 621 2298 623 2327
rect 589 2293 623 2298
rect 657 2298 659 2327
rect 693 2331 733 2332
rect 768 2343 802 2365
rect 768 2331 836 2343
rect 693 2309 836 2331
rect 693 2298 802 2309
rect 657 2297 802 2298
rect 657 2293 734 2297
rect 555 2292 734 2293
rect 555 2259 733 2292
rect 768 2275 802 2297
rect 768 2263 836 2275
rect 555 2250 587 2259
rect 621 2250 659 2259
rect 621 2225 623 2250
rect 589 2216 623 2225
rect 657 2225 659 2250
rect 693 2258 733 2259
rect 767 2258 836 2263
rect 693 2241 836 2258
rect 693 2229 802 2241
rect 693 2225 734 2229
rect 657 2219 734 2225
rect 657 2216 733 2219
rect 555 2186 733 2216
rect 768 2207 802 2229
rect 768 2195 836 2207
rect 555 2156 587 2186
rect 621 2156 659 2186
rect 621 2152 623 2156
rect 589 2122 623 2152
rect 657 2152 659 2156
rect 693 2185 733 2186
rect 767 2185 836 2195
rect 693 2173 836 2185
rect 693 2161 802 2173
rect 693 2152 734 2161
rect 657 2146 734 2152
rect 657 2122 733 2146
rect 768 2139 802 2161
rect 768 2127 836 2139
rect 555 2113 733 2122
rect 555 2085 587 2113
rect 621 2085 659 2113
rect 621 2079 623 2085
rect 589 2051 623 2079
rect 657 2079 659 2085
rect 693 2112 733 2113
rect 767 2112 836 2127
rect 693 2105 836 2112
rect 693 2093 802 2105
rect 693 2079 734 2093
rect 657 2073 734 2079
rect 657 2051 733 2073
rect 768 2071 802 2093
rect 768 2059 836 2071
rect 555 2040 733 2051
rect 555 2011 587 2040
rect 621 2011 659 2040
rect 621 2006 623 2011
rect 589 1977 623 2006
rect 657 2006 659 2011
rect 693 2039 733 2040
rect 767 2039 836 2059
rect 693 2037 836 2039
rect 693 2025 802 2037
rect 693 2006 734 2025
rect 657 2000 734 2006
rect 768 2003 802 2025
rect 657 1977 733 2000
rect 768 1991 836 2003
rect 555 1967 733 1977
rect 555 1940 587 1967
rect 621 1940 659 1967
rect 621 1933 623 1940
rect 589 1906 623 1933
rect 657 1933 659 1940
rect 693 1966 733 1967
rect 767 1969 836 1991
rect 767 1966 802 1969
rect 693 1957 802 1966
rect 693 1933 734 1957
rect 657 1927 734 1933
rect 768 1935 802 1957
rect 657 1906 733 1927
rect 768 1923 836 1935
rect 555 1894 733 1906
rect 555 1866 587 1894
rect 621 1866 659 1894
rect 621 1860 623 1866
rect 589 1832 623 1860
rect 657 1860 659 1866
rect 693 1893 733 1894
rect 767 1901 836 1923
rect 767 1893 802 1901
rect 693 1889 802 1893
rect 693 1860 734 1889
rect 657 1855 734 1860
rect 768 1867 802 1889
rect 768 1855 836 1867
rect 657 1854 836 1855
rect 657 1832 733 1854
rect 555 1821 733 1832
rect 767 1833 836 1854
rect 767 1821 802 1833
rect 555 1795 587 1821
rect 621 1795 659 1821
rect 621 1787 623 1795
rect 589 1761 623 1787
rect 657 1787 659 1795
rect 693 1820 733 1821
rect 693 1787 734 1820
rect 768 1799 802 1821
rect 768 1787 836 1799
rect 657 1781 836 1787
rect 657 1761 733 1781
rect 555 1748 733 1761
rect 767 1765 836 1781
rect 767 1753 802 1765
rect 555 1721 587 1748
rect 621 1721 659 1748
rect 621 1714 623 1721
rect 589 1687 623 1714
rect 657 1714 659 1721
rect 693 1747 733 1748
rect 693 1719 734 1747
rect 768 1731 802 1753
rect 768 1719 836 1731
rect 693 1714 836 1719
rect 657 1708 836 1714
rect 657 1687 733 1708
rect 555 1675 733 1687
rect 767 1697 836 1708
rect 767 1685 802 1697
rect 555 1650 587 1675
rect 621 1650 659 1675
rect 621 1641 623 1650
rect 589 1616 623 1641
rect 657 1641 659 1650
rect 693 1674 733 1675
rect 693 1651 734 1674
rect 768 1663 802 1685
rect 768 1651 836 1663
rect 693 1641 836 1651
rect 657 1635 836 1641
rect 657 1616 733 1635
rect 767 1629 836 1635
rect 767 1617 802 1629
rect 555 1602 733 1616
rect 555 1576 587 1602
rect 621 1576 659 1602
rect 621 1568 623 1576
rect 589 1542 623 1568
rect 657 1568 659 1576
rect 693 1601 733 1602
rect 693 1583 734 1601
rect 768 1595 802 1617
rect 768 1583 836 1595
rect 693 1568 836 1583
rect 657 1562 836 1568
rect 657 1542 733 1562
rect 767 1561 836 1562
rect 767 1549 802 1561
rect 555 1529 733 1542
rect 555 1505 587 1529
rect 621 1505 659 1529
rect 621 1495 623 1505
rect 589 1471 623 1495
rect 657 1495 659 1505
rect 693 1528 733 1529
rect 693 1515 734 1528
rect 768 1527 802 1549
rect 768 1515 836 1527
rect 693 1499 836 1515
rect 693 1495 822 1499
rect 657 1489 822 1495
rect 657 1471 733 1489
rect 555 1455 733 1471
rect 767 1455 822 1489
rect 555 1419 822 1455
rect 555 1385 587 1419
rect 621 1385 659 1419
rect 693 1416 822 1419
rect 693 1385 733 1416
rect 555 1382 733 1385
rect 767 1382 822 1416
rect 555 1375 822 1382
rect 589 1341 623 1375
rect 657 1341 691 1375
rect 725 1342 822 1375
rect 725 1341 733 1342
rect 555 1330 733 1341
rect 555 1296 587 1330
rect 621 1296 659 1330
rect 693 1308 733 1330
rect 767 1308 822 1342
rect 693 1296 822 1308
rect 555 1268 822 1296
rect 924 1409 1044 2505
rect 1109 4028 1110 4062
rect 1144 4046 1182 4062
rect 1144 4028 1146 4046
rect 1109 4012 1146 4028
rect 1180 4028 1182 4046
rect 1216 4046 1254 4062
rect 1216 4028 1218 4046
rect 1180 4012 1218 4028
rect 1252 4028 1254 4046
rect 1288 4028 1289 4062
rect 1252 4012 1289 4028
rect 1109 3988 1289 4012
rect 1109 3954 1110 3988
rect 1144 3978 1182 3988
rect 1144 3954 1146 3978
rect 1109 3944 1146 3954
rect 1180 3954 1182 3978
rect 1216 3978 1254 3988
rect 1216 3954 1218 3978
rect 1180 3944 1218 3954
rect 1252 3954 1254 3978
rect 1288 3954 1289 3988
rect 1252 3944 1289 3954
rect 1109 3914 1289 3944
rect 1109 3880 1110 3914
rect 1144 3910 1182 3914
rect 1144 3880 1146 3910
rect 1109 3876 1146 3880
rect 1180 3880 1182 3910
rect 1216 3910 1254 3914
rect 1216 3880 1218 3910
rect 1180 3876 1218 3880
rect 1252 3880 1254 3910
rect 1288 3880 1289 3914
rect 1252 3876 1289 3880
rect 1109 3842 1289 3876
rect 1109 3840 1146 3842
rect 1109 3806 1110 3840
rect 1144 3808 1146 3840
rect 1180 3840 1218 3842
rect 1180 3808 1182 3840
rect 1144 3806 1182 3808
rect 1216 3808 1218 3840
rect 1252 3840 1289 3842
rect 1252 3808 1254 3840
rect 1216 3806 1254 3808
rect 1288 3806 1289 3840
rect 1109 3774 1289 3806
rect 1109 3766 1146 3774
rect 1109 3732 1110 3766
rect 1144 3740 1146 3766
rect 1180 3766 1218 3774
rect 1180 3740 1182 3766
rect 1144 3732 1182 3740
rect 1216 3740 1218 3766
rect 1252 3766 1289 3774
rect 1252 3740 1254 3766
rect 1216 3732 1254 3740
rect 1288 3732 1289 3766
rect 1109 3706 1289 3732
rect 1109 3692 1146 3706
rect 1109 3658 1110 3692
rect 1144 3672 1146 3692
rect 1180 3692 1218 3706
rect 1180 3672 1182 3692
rect 1144 3658 1182 3672
rect 1216 3672 1218 3692
rect 1252 3692 1289 3706
rect 1252 3672 1254 3692
rect 1216 3658 1254 3672
rect 1288 3658 1289 3692
rect 1109 3638 1289 3658
rect 1109 3618 1146 3638
rect 1109 3584 1110 3618
rect 1144 3604 1146 3618
rect 1180 3618 1218 3638
rect 1180 3604 1182 3618
rect 1144 3584 1182 3604
rect 1216 3604 1218 3618
rect 1252 3618 1289 3638
rect 1252 3604 1254 3618
rect 1216 3584 1254 3604
rect 1288 3584 1289 3618
rect 1109 3570 1289 3584
rect 1109 3544 1146 3570
rect 1109 3510 1110 3544
rect 1144 3536 1146 3544
rect 1180 3544 1218 3570
rect 1180 3536 1182 3544
rect 1144 3510 1182 3536
rect 1216 3536 1218 3544
rect 1252 3544 1289 3570
rect 1252 3536 1254 3544
rect 1216 3510 1254 3536
rect 1288 3510 1289 3544
rect 1109 3502 1289 3510
rect 1109 3470 1146 3502
rect 1109 3436 1110 3470
rect 1144 3468 1146 3470
rect 1180 3470 1218 3502
rect 1180 3468 1182 3470
rect 1144 3436 1182 3468
rect 1216 3468 1218 3470
rect 1252 3470 1289 3502
rect 1252 3468 1254 3470
rect 1216 3436 1254 3468
rect 1288 3436 1289 3470
rect 1109 3434 1289 3436
rect 1109 3400 1146 3434
rect 1180 3400 1218 3434
rect 1252 3400 1289 3434
rect 1109 3396 1289 3400
rect 1109 3362 1110 3396
rect 1144 3366 1182 3396
rect 1144 3362 1146 3366
rect 1109 3332 1146 3362
rect 1180 3362 1182 3366
rect 1216 3366 1254 3396
rect 1216 3362 1218 3366
rect 1180 3332 1218 3362
rect 1252 3362 1254 3366
rect 1288 3362 1289 3396
rect 1252 3332 1289 3362
rect 1109 3322 1289 3332
rect 1109 3288 1110 3322
rect 1144 3298 1182 3322
rect 1144 3288 1146 3298
rect 1109 3264 1146 3288
rect 1180 3288 1182 3298
rect 1216 3298 1254 3322
rect 1216 3288 1218 3298
rect 1180 3264 1218 3288
rect 1252 3288 1254 3298
rect 1288 3288 1289 3322
rect 1252 3264 1289 3288
rect 1109 3248 1289 3264
rect 1109 3214 1110 3248
rect 1144 3230 1182 3248
rect 1144 3214 1146 3230
rect 1109 3196 1146 3214
rect 1180 3214 1182 3230
rect 1216 3230 1254 3248
rect 1216 3214 1218 3230
rect 1180 3196 1218 3214
rect 1252 3214 1254 3230
rect 1288 3214 1289 3248
rect 1252 3196 1289 3214
rect 1109 3174 1289 3196
rect 1109 3140 1110 3174
rect 1144 3162 1182 3174
rect 1144 3140 1146 3162
rect 1109 3128 1146 3140
rect 1180 3140 1182 3162
rect 1216 3162 1254 3174
rect 1216 3140 1218 3162
rect 1180 3128 1218 3140
rect 1252 3140 1254 3162
rect 1288 3140 1289 3174
rect 1252 3128 1289 3140
rect 1109 3100 1289 3128
rect 1109 3066 1110 3100
rect 1144 3066 1182 3100
rect 1216 3066 1254 3100
rect 1288 3066 1289 3100
rect 1109 3026 1289 3066
rect 1109 2992 1110 3026
rect 1144 2992 1182 3026
rect 1216 2992 1254 3026
rect 1288 2992 1289 3026
rect 1109 2952 1289 2992
rect 1109 2918 1110 2952
rect 1144 2918 1182 2952
rect 1216 2918 1254 2952
rect 1288 2918 1289 2952
rect 1109 2878 1289 2918
rect 1109 2844 1110 2878
rect 1144 2844 1182 2878
rect 1216 2844 1254 2878
rect 1288 2844 1289 2878
rect 1109 2804 1289 2844
rect 1109 2770 1110 2804
rect 1144 2770 1182 2804
rect 1216 2770 1254 2804
rect 1288 2770 1289 2804
rect 1109 2730 1289 2770
rect 1109 2696 1110 2730
rect 1144 2696 1182 2730
rect 1216 2696 1254 2730
rect 1288 2696 1289 2730
rect 1109 2656 1289 2696
rect 1109 2622 1110 2656
rect 1144 2622 1182 2656
rect 1216 2622 1254 2656
rect 1288 2622 1289 2656
rect 1109 2582 1289 2622
rect 1109 2548 1110 2582
rect 1144 2548 1182 2582
rect 1216 2548 1254 2582
rect 1288 2548 1289 2582
rect 1109 2508 1289 2548
rect 1109 2474 1110 2508
rect 1144 2474 1182 2508
rect 1216 2474 1254 2508
rect 1288 2474 1289 2508
rect 1109 2445 1289 2474
rect 1109 2434 1146 2445
rect 1109 2400 1110 2434
rect 1144 2411 1146 2434
rect 1180 2434 1218 2445
rect 1180 2411 1182 2434
rect 1144 2400 1182 2411
rect 1216 2411 1218 2434
rect 1252 2434 1289 2445
rect 1252 2411 1254 2434
rect 1216 2400 1254 2411
rect 1288 2400 1289 2434
rect 1109 2377 1289 2400
rect 1109 2360 1146 2377
rect 1109 2326 1110 2360
rect 1144 2343 1146 2360
rect 1180 2360 1218 2377
rect 1180 2343 1182 2360
rect 1144 2326 1182 2343
rect 1216 2343 1218 2360
rect 1252 2360 1289 2377
rect 1252 2343 1254 2360
rect 1216 2326 1254 2343
rect 1288 2326 1289 2360
rect 1109 2309 1289 2326
rect 1109 2286 1146 2309
rect 1109 2252 1110 2286
rect 1144 2275 1146 2286
rect 1180 2286 1218 2309
rect 1180 2275 1182 2286
rect 1144 2252 1182 2275
rect 1216 2275 1218 2286
rect 1252 2286 1289 2309
rect 1252 2275 1254 2286
rect 1216 2252 1254 2275
rect 1288 2252 1289 2286
rect 1109 2241 1289 2252
rect 1109 2212 1146 2241
rect 1109 2178 1110 2212
rect 1144 2207 1146 2212
rect 1180 2212 1218 2241
rect 1180 2207 1182 2212
rect 1144 2178 1182 2207
rect 1216 2207 1218 2212
rect 1252 2212 1289 2241
rect 1252 2207 1254 2212
rect 1216 2178 1254 2207
rect 1288 2178 1289 2212
rect 1109 2173 1289 2178
rect 1109 2139 1146 2173
rect 1180 2139 1218 2173
rect 1252 2139 1289 2173
rect 1109 2138 1289 2139
rect 1109 2104 1110 2138
rect 1144 2105 1182 2138
rect 1144 2104 1146 2105
rect 1109 2071 1146 2104
rect 1180 2104 1182 2105
rect 1216 2105 1254 2138
rect 1216 2104 1218 2105
rect 1180 2071 1218 2104
rect 1252 2104 1254 2105
rect 1288 2104 1289 2138
rect 1252 2071 1289 2104
rect 1109 2064 1289 2071
rect 1109 2030 1110 2064
rect 1144 2037 1182 2064
rect 1144 2030 1146 2037
rect 1109 2003 1146 2030
rect 1180 2030 1182 2037
rect 1216 2037 1254 2064
rect 1216 2030 1218 2037
rect 1180 2003 1218 2030
rect 1252 2030 1254 2037
rect 1288 2030 1289 2064
rect 1252 2003 1289 2030
rect 1109 1990 1289 2003
rect 1109 1956 1110 1990
rect 1144 1969 1182 1990
rect 1144 1956 1146 1969
rect 1109 1935 1146 1956
rect 1180 1956 1182 1969
rect 1216 1969 1254 1990
rect 1216 1956 1218 1969
rect 1180 1935 1218 1956
rect 1252 1956 1254 1969
rect 1288 1956 1289 1990
rect 1252 1935 1289 1956
rect 1109 1916 1289 1935
rect 1109 1882 1110 1916
rect 1144 1901 1182 1916
rect 1144 1882 1146 1901
rect 1109 1867 1146 1882
rect 1180 1882 1182 1901
rect 1216 1901 1254 1916
rect 1216 1882 1218 1901
rect 1180 1867 1218 1882
rect 1252 1882 1254 1901
rect 1288 1882 1289 1916
rect 1252 1867 1289 1882
rect 1109 1842 1289 1867
rect 1109 1808 1110 1842
rect 1144 1833 1182 1842
rect 1144 1808 1146 1833
rect 1109 1799 1146 1808
rect 1180 1808 1182 1833
rect 1216 1833 1254 1842
rect 1216 1808 1218 1833
rect 1180 1799 1218 1808
rect 1252 1808 1254 1833
rect 1288 1808 1289 1842
rect 1252 1799 1289 1808
rect 1109 1768 1289 1799
rect 1109 1734 1110 1768
rect 1144 1765 1182 1768
rect 1144 1734 1146 1765
rect 1109 1731 1146 1734
rect 1180 1734 1182 1765
rect 1216 1765 1254 1768
rect 1216 1734 1218 1765
rect 1180 1731 1218 1734
rect 1252 1734 1254 1765
rect 1288 1734 1289 1768
rect 1252 1731 1289 1734
rect 1109 1697 1289 1731
rect 1109 1694 1146 1697
rect 1109 1660 1110 1694
rect 1144 1663 1146 1694
rect 1180 1694 1218 1697
rect 1180 1663 1182 1694
rect 1144 1660 1182 1663
rect 1216 1663 1218 1694
rect 1252 1694 1289 1697
rect 1252 1663 1254 1694
rect 1216 1660 1254 1663
rect 1288 1660 1289 1694
rect 1109 1629 1289 1660
rect 1109 1620 1146 1629
rect 1109 1586 1110 1620
rect 1144 1595 1146 1620
rect 1180 1620 1218 1629
rect 1180 1595 1182 1620
rect 1144 1586 1182 1595
rect 1216 1595 1218 1620
rect 1252 1620 1289 1629
rect 1252 1595 1254 1620
rect 1216 1586 1254 1595
rect 1288 1586 1289 1620
rect 1109 1561 1289 1586
rect 1109 1545 1146 1561
rect 1109 1511 1110 1545
rect 1144 1527 1146 1545
rect 1180 1545 1218 1561
rect 1180 1527 1182 1545
rect 1144 1511 1182 1527
rect 1216 1527 1218 1545
rect 1252 1545 1289 1561
rect 1252 1527 1254 1545
rect 1216 1511 1254 1527
rect 1288 1511 1289 1545
rect 1354 3010 1474 4106
rect 1916 4388 1923 4494
rect 2029 4388 2036 4494
rect 1916 4214 2036 4388
rect 1916 4180 1959 4214
rect 1993 4180 2036 4214
rect 1916 4140 2036 4180
rect 1916 4106 1959 4140
rect 1993 4106 2036 4140
rect 1354 2976 1397 3010
rect 1431 2976 1474 3010
rect 1354 2932 1474 2976
rect 1354 2898 1397 2932
rect 1431 2898 1474 2932
rect 1354 2854 1474 2898
rect 1354 2820 1397 2854
rect 1431 2820 1474 2854
rect 1354 2776 1474 2820
rect 1354 2742 1397 2776
rect 1431 2742 1474 2776
rect 1354 2697 1474 2742
rect 1354 2663 1397 2697
rect 1431 2663 1474 2697
rect 1354 2618 1474 2663
rect 1354 2584 1397 2618
rect 1431 2584 1474 2618
rect 1354 2539 1474 2584
rect 1354 2505 1397 2539
rect 1431 2505 1474 2539
rect 1146 1491 1252 1511
rect 924 1375 967 1409
rect 1001 1375 1044 1409
rect 924 1335 1044 1375
rect 924 1301 967 1335
rect 1001 1301 1044 1335
rect 924 1285 1044 1301
rect 1354 1409 1474 2505
rect 1576 4050 1678 4062
rect 1712 4050 1814 4062
rect 1576 4046 1606 4050
rect 1784 4046 1814 4050
rect 1576 3978 1606 4012
rect 1784 3978 1814 4012
rect 1576 3910 1606 3944
rect 1784 3910 1814 3944
rect 1576 3842 1606 3876
rect 1784 3842 1814 3876
rect 1576 3774 1606 3808
rect 1784 3774 1814 3808
rect 1576 3706 1606 3740
rect 1784 3706 1814 3740
rect 1576 3638 1606 3672
rect 1784 3638 1814 3672
rect 1576 3570 1606 3604
rect 1784 3570 1814 3604
rect 1576 3502 1606 3536
rect 1784 3502 1814 3536
rect 1576 3434 1606 3468
rect 1784 3434 1814 3468
rect 1576 3366 1606 3400
rect 1784 3366 1814 3400
rect 1576 3298 1606 3332
rect 1784 3298 1814 3332
rect 1576 3230 1606 3264
rect 1784 3230 1814 3264
rect 1576 3162 1606 3196
rect 1784 3162 1814 3196
rect 1576 3080 1606 3128
rect 1640 3080 1750 3092
rect 1784 3080 1814 3128
rect 1576 3040 1814 3080
rect 1576 2574 1606 3040
rect 1784 2574 1814 3040
rect 1576 2535 1814 2574
rect 1576 2501 1606 2535
rect 1640 2501 1678 2535
rect 1712 2501 1750 2535
rect 1784 2501 1814 2535
rect 1576 2461 1814 2501
rect 1576 2449 1678 2461
rect 1712 2449 1814 2461
rect 1576 2445 1606 2449
rect 1784 2445 1814 2449
rect 1576 2377 1606 2411
rect 1784 2377 1814 2411
rect 1576 2309 1606 2343
rect 1784 2309 1814 2343
rect 1576 2241 1606 2275
rect 1784 2241 1814 2275
rect 1576 2173 1606 2207
rect 1784 2173 1814 2207
rect 1576 2105 1606 2139
rect 1784 2105 1814 2139
rect 1576 2037 1606 2071
rect 1784 2037 1814 2071
rect 1576 1969 1606 2003
rect 1784 1969 1814 2003
rect 1576 1901 1606 1935
rect 1784 1901 1814 1935
rect 1576 1833 1606 1867
rect 1784 1833 1814 1867
rect 1576 1765 1606 1799
rect 1784 1765 1814 1799
rect 1576 1697 1606 1731
rect 1784 1697 1814 1731
rect 1576 1629 1606 1663
rect 1784 1629 1814 1663
rect 1576 1561 1606 1595
rect 1784 1561 1814 1595
rect 1576 1479 1606 1527
rect 1640 1479 1750 1491
rect 1784 1479 1814 1527
rect 1576 1464 1814 1479
rect 1916 3010 2036 4106
rect 2346 4388 2353 4494
rect 2459 4388 2466 4494
rect 2346 4214 2466 4388
rect 2346 4180 2389 4214
rect 2423 4180 2466 4214
rect 2346 4140 2466 4180
rect 2346 4106 2389 4140
rect 2423 4106 2466 4140
rect 1916 2976 1959 3010
rect 1993 2976 2036 3010
rect 1916 2932 2036 2976
rect 1916 2898 1959 2932
rect 1993 2898 2036 2932
rect 1916 2854 2036 2898
rect 1916 2820 1959 2854
rect 1993 2820 2036 2854
rect 1916 2776 2036 2820
rect 1916 2742 1959 2776
rect 1993 2742 2036 2776
rect 1916 2697 2036 2742
rect 1916 2663 1959 2697
rect 1993 2663 2036 2697
rect 1916 2618 2036 2663
rect 1916 2584 1959 2618
rect 1993 2584 2036 2618
rect 1916 2539 2036 2584
rect 1916 2505 1959 2539
rect 1993 2505 2036 2539
rect 1354 1375 1397 1409
rect 1431 1375 1474 1409
rect 1354 1335 1474 1375
rect 1354 1301 1397 1335
rect 1431 1301 1474 1335
rect 1354 1285 1474 1301
rect 1916 1409 2036 2505
rect 2101 4028 2102 4062
rect 2136 4046 2174 4062
rect 2136 4028 2138 4046
rect 2101 4012 2138 4028
rect 2172 4028 2174 4046
rect 2208 4046 2246 4062
rect 2208 4028 2210 4046
rect 2172 4012 2210 4028
rect 2244 4028 2246 4046
rect 2280 4028 2281 4062
rect 2244 4012 2281 4028
rect 2101 3988 2281 4012
rect 2101 3954 2102 3988
rect 2136 3978 2174 3988
rect 2136 3954 2138 3978
rect 2101 3944 2138 3954
rect 2172 3954 2174 3978
rect 2208 3978 2246 3988
rect 2208 3954 2210 3978
rect 2172 3944 2210 3954
rect 2244 3954 2246 3978
rect 2280 3954 2281 3988
rect 2244 3944 2281 3954
rect 2101 3914 2281 3944
rect 2101 3880 2102 3914
rect 2136 3910 2174 3914
rect 2136 3880 2138 3910
rect 2101 3876 2138 3880
rect 2172 3880 2174 3910
rect 2208 3910 2246 3914
rect 2208 3880 2210 3910
rect 2172 3876 2210 3880
rect 2244 3880 2246 3910
rect 2280 3880 2281 3914
rect 2244 3876 2281 3880
rect 2101 3842 2281 3876
rect 2101 3840 2138 3842
rect 2101 3806 2102 3840
rect 2136 3808 2138 3840
rect 2172 3840 2210 3842
rect 2172 3808 2174 3840
rect 2136 3806 2174 3808
rect 2208 3808 2210 3840
rect 2244 3840 2281 3842
rect 2244 3808 2246 3840
rect 2208 3806 2246 3808
rect 2280 3806 2281 3840
rect 2101 3774 2281 3806
rect 2101 3766 2138 3774
rect 2101 3732 2102 3766
rect 2136 3740 2138 3766
rect 2172 3766 2210 3774
rect 2172 3740 2174 3766
rect 2136 3732 2174 3740
rect 2208 3740 2210 3766
rect 2244 3766 2281 3774
rect 2244 3740 2246 3766
rect 2208 3732 2246 3740
rect 2280 3732 2281 3766
rect 2101 3706 2281 3732
rect 2101 3692 2138 3706
rect 2101 3658 2102 3692
rect 2136 3672 2138 3692
rect 2172 3692 2210 3706
rect 2172 3672 2174 3692
rect 2136 3658 2174 3672
rect 2208 3672 2210 3692
rect 2244 3692 2281 3706
rect 2244 3672 2246 3692
rect 2208 3658 2246 3672
rect 2280 3658 2281 3692
rect 2101 3638 2281 3658
rect 2101 3618 2138 3638
rect 2101 3584 2102 3618
rect 2136 3604 2138 3618
rect 2172 3618 2210 3638
rect 2172 3604 2174 3618
rect 2136 3584 2174 3604
rect 2208 3604 2210 3618
rect 2244 3618 2281 3638
rect 2244 3604 2246 3618
rect 2208 3584 2246 3604
rect 2280 3584 2281 3618
rect 2101 3570 2281 3584
rect 2101 3544 2138 3570
rect 2101 3510 2102 3544
rect 2136 3536 2138 3544
rect 2172 3544 2210 3570
rect 2172 3536 2174 3544
rect 2136 3510 2174 3536
rect 2208 3536 2210 3544
rect 2244 3544 2281 3570
rect 2244 3536 2246 3544
rect 2208 3510 2246 3536
rect 2280 3510 2281 3544
rect 2101 3502 2281 3510
rect 2101 3470 2138 3502
rect 2101 3436 2102 3470
rect 2136 3468 2138 3470
rect 2172 3470 2210 3502
rect 2172 3468 2174 3470
rect 2136 3436 2174 3468
rect 2208 3468 2210 3470
rect 2244 3470 2281 3502
rect 2244 3468 2246 3470
rect 2208 3436 2246 3468
rect 2280 3436 2281 3470
rect 2101 3434 2281 3436
rect 2101 3400 2138 3434
rect 2172 3400 2210 3434
rect 2244 3400 2281 3434
rect 2101 3396 2281 3400
rect 2101 3362 2102 3396
rect 2136 3366 2174 3396
rect 2136 3362 2138 3366
rect 2101 3332 2138 3362
rect 2172 3362 2174 3366
rect 2208 3366 2246 3396
rect 2208 3362 2210 3366
rect 2172 3332 2210 3362
rect 2244 3362 2246 3366
rect 2280 3362 2281 3396
rect 2244 3332 2281 3362
rect 2101 3322 2281 3332
rect 2101 3288 2102 3322
rect 2136 3298 2174 3322
rect 2136 3288 2138 3298
rect 2101 3264 2138 3288
rect 2172 3288 2174 3298
rect 2208 3298 2246 3322
rect 2208 3288 2210 3298
rect 2172 3264 2210 3288
rect 2244 3288 2246 3298
rect 2280 3288 2281 3322
rect 2244 3264 2281 3288
rect 2101 3248 2281 3264
rect 2101 3214 2102 3248
rect 2136 3230 2174 3248
rect 2136 3214 2138 3230
rect 2101 3196 2138 3214
rect 2172 3214 2174 3230
rect 2208 3230 2246 3248
rect 2208 3214 2210 3230
rect 2172 3196 2210 3214
rect 2244 3214 2246 3230
rect 2280 3214 2281 3248
rect 2244 3196 2281 3214
rect 2101 3174 2281 3196
rect 2101 3140 2102 3174
rect 2136 3162 2174 3174
rect 2136 3140 2138 3162
rect 2101 3128 2138 3140
rect 2172 3140 2174 3162
rect 2208 3162 2246 3174
rect 2208 3140 2210 3162
rect 2172 3128 2210 3140
rect 2244 3140 2246 3162
rect 2280 3140 2281 3174
rect 2244 3128 2281 3140
rect 2101 3100 2281 3128
rect 2101 3066 2102 3100
rect 2136 3066 2174 3100
rect 2208 3066 2246 3100
rect 2280 3066 2281 3100
rect 2101 3026 2281 3066
rect 2101 2992 2102 3026
rect 2136 2992 2174 3026
rect 2208 2992 2246 3026
rect 2280 2992 2281 3026
rect 2101 2952 2281 2992
rect 2101 2918 2102 2952
rect 2136 2918 2174 2952
rect 2208 2918 2246 2952
rect 2280 2918 2281 2952
rect 2101 2878 2281 2918
rect 2101 2844 2102 2878
rect 2136 2844 2174 2878
rect 2208 2844 2246 2878
rect 2280 2844 2281 2878
rect 2101 2804 2281 2844
rect 2101 2770 2102 2804
rect 2136 2770 2174 2804
rect 2208 2770 2246 2804
rect 2280 2770 2281 2804
rect 2101 2730 2281 2770
rect 2101 2696 2102 2730
rect 2136 2696 2174 2730
rect 2208 2696 2246 2730
rect 2280 2696 2281 2730
rect 2101 2656 2281 2696
rect 2101 2622 2102 2656
rect 2136 2622 2174 2656
rect 2208 2622 2246 2656
rect 2280 2622 2281 2656
rect 2101 2582 2281 2622
rect 2101 2548 2102 2582
rect 2136 2548 2174 2582
rect 2208 2548 2246 2582
rect 2280 2548 2281 2582
rect 2101 2508 2281 2548
rect 2101 2474 2102 2508
rect 2136 2474 2174 2508
rect 2208 2474 2246 2508
rect 2280 2474 2281 2508
rect 2101 2445 2281 2474
rect 2101 2434 2138 2445
rect 2101 2400 2102 2434
rect 2136 2411 2138 2434
rect 2172 2434 2210 2445
rect 2172 2411 2174 2434
rect 2136 2400 2174 2411
rect 2208 2411 2210 2434
rect 2244 2434 2281 2445
rect 2244 2411 2246 2434
rect 2208 2400 2246 2411
rect 2280 2400 2281 2434
rect 2101 2377 2281 2400
rect 2101 2360 2138 2377
rect 2101 2326 2102 2360
rect 2136 2343 2138 2360
rect 2172 2360 2210 2377
rect 2172 2343 2174 2360
rect 2136 2326 2174 2343
rect 2208 2343 2210 2360
rect 2244 2360 2281 2377
rect 2244 2343 2246 2360
rect 2208 2326 2246 2343
rect 2280 2326 2281 2360
rect 2101 2309 2281 2326
rect 2101 2286 2138 2309
rect 2101 2252 2102 2286
rect 2136 2275 2138 2286
rect 2172 2286 2210 2309
rect 2172 2275 2174 2286
rect 2136 2252 2174 2275
rect 2208 2275 2210 2286
rect 2244 2286 2281 2309
rect 2244 2275 2246 2286
rect 2208 2252 2246 2275
rect 2280 2252 2281 2286
rect 2101 2241 2281 2252
rect 2101 2212 2138 2241
rect 2101 2178 2102 2212
rect 2136 2207 2138 2212
rect 2172 2212 2210 2241
rect 2172 2207 2174 2212
rect 2136 2178 2174 2207
rect 2208 2207 2210 2212
rect 2244 2212 2281 2241
rect 2244 2207 2246 2212
rect 2208 2178 2246 2207
rect 2280 2178 2281 2212
rect 2101 2173 2281 2178
rect 2101 2139 2138 2173
rect 2172 2139 2210 2173
rect 2244 2139 2281 2173
rect 2101 2138 2281 2139
rect 2101 2104 2102 2138
rect 2136 2105 2174 2138
rect 2136 2104 2138 2105
rect 2101 2071 2138 2104
rect 2172 2104 2174 2105
rect 2208 2105 2246 2138
rect 2208 2104 2210 2105
rect 2172 2071 2210 2104
rect 2244 2104 2246 2105
rect 2280 2104 2281 2138
rect 2244 2071 2281 2104
rect 2101 2064 2281 2071
rect 2101 2030 2102 2064
rect 2136 2037 2174 2064
rect 2136 2030 2138 2037
rect 2101 2003 2138 2030
rect 2172 2030 2174 2037
rect 2208 2037 2246 2064
rect 2208 2030 2210 2037
rect 2172 2003 2210 2030
rect 2244 2030 2246 2037
rect 2280 2030 2281 2064
rect 2244 2003 2281 2030
rect 2101 1990 2281 2003
rect 2101 1956 2102 1990
rect 2136 1969 2174 1990
rect 2136 1956 2138 1969
rect 2101 1935 2138 1956
rect 2172 1956 2174 1969
rect 2208 1969 2246 1990
rect 2208 1956 2210 1969
rect 2172 1935 2210 1956
rect 2244 1956 2246 1969
rect 2280 1956 2281 1990
rect 2244 1935 2281 1956
rect 2101 1916 2281 1935
rect 2101 1882 2102 1916
rect 2136 1901 2174 1916
rect 2136 1882 2138 1901
rect 2101 1867 2138 1882
rect 2172 1882 2174 1901
rect 2208 1901 2246 1916
rect 2208 1882 2210 1901
rect 2172 1867 2210 1882
rect 2244 1882 2246 1901
rect 2280 1882 2281 1916
rect 2244 1867 2281 1882
rect 2101 1842 2281 1867
rect 2101 1808 2102 1842
rect 2136 1833 2174 1842
rect 2136 1808 2138 1833
rect 2101 1799 2138 1808
rect 2172 1808 2174 1833
rect 2208 1833 2246 1842
rect 2208 1808 2210 1833
rect 2172 1799 2210 1808
rect 2244 1808 2246 1833
rect 2280 1808 2281 1842
rect 2244 1799 2281 1808
rect 2101 1768 2281 1799
rect 2101 1734 2102 1768
rect 2136 1765 2174 1768
rect 2136 1734 2138 1765
rect 2101 1731 2138 1734
rect 2172 1734 2174 1765
rect 2208 1765 2246 1768
rect 2208 1734 2210 1765
rect 2172 1731 2210 1734
rect 2244 1734 2246 1765
rect 2280 1734 2281 1768
rect 2244 1731 2281 1734
rect 2101 1697 2281 1731
rect 2101 1694 2138 1697
rect 2101 1660 2102 1694
rect 2136 1663 2138 1694
rect 2172 1694 2210 1697
rect 2172 1663 2174 1694
rect 2136 1660 2174 1663
rect 2208 1663 2210 1694
rect 2244 1694 2281 1697
rect 2244 1663 2246 1694
rect 2208 1660 2246 1663
rect 2280 1660 2281 1694
rect 2101 1629 2281 1660
rect 2101 1620 2138 1629
rect 2101 1586 2102 1620
rect 2136 1595 2138 1620
rect 2172 1620 2210 1629
rect 2172 1595 2174 1620
rect 2136 1586 2174 1595
rect 2208 1595 2210 1620
rect 2244 1620 2281 1629
rect 2244 1595 2246 1620
rect 2208 1586 2246 1595
rect 2280 1586 2281 1620
rect 2101 1561 2281 1586
rect 2101 1545 2138 1561
rect 2101 1511 2102 1545
rect 2136 1527 2138 1545
rect 2172 1545 2210 1561
rect 2172 1527 2174 1545
rect 2136 1511 2174 1527
rect 2208 1527 2210 1545
rect 2244 1545 2281 1561
rect 2244 1527 2246 1545
rect 2208 1511 2246 1527
rect 2280 1511 2281 1545
rect 2346 3010 2466 4106
rect 2908 4388 2915 4494
rect 3021 4388 3028 4494
rect 2908 4214 3028 4388
rect 2908 4180 2951 4214
rect 2985 4180 3028 4214
rect 2908 4140 3028 4180
rect 2908 4106 2951 4140
rect 2985 4106 3028 4140
rect 2346 2976 2389 3010
rect 2423 2976 2466 3010
rect 2346 2932 2466 2976
rect 2346 2898 2389 2932
rect 2423 2898 2466 2932
rect 2346 2854 2466 2898
rect 2346 2820 2389 2854
rect 2423 2820 2466 2854
rect 2346 2776 2466 2820
rect 2346 2742 2389 2776
rect 2423 2742 2466 2776
rect 2346 2697 2466 2742
rect 2346 2663 2389 2697
rect 2423 2663 2466 2697
rect 2346 2618 2466 2663
rect 2346 2584 2389 2618
rect 2423 2584 2466 2618
rect 2346 2539 2466 2584
rect 2346 2505 2389 2539
rect 2423 2505 2466 2539
rect 2138 1491 2244 1511
rect 1916 1375 1959 1409
rect 1993 1375 2036 1409
rect 1916 1335 2036 1375
rect 1916 1301 1959 1335
rect 1993 1301 2036 1335
rect 1916 1285 2036 1301
rect 2346 1409 2466 2505
rect 2568 4050 2670 4062
rect 2704 4050 2806 4062
rect 2568 4046 2598 4050
rect 2776 4046 2806 4050
rect 2568 3978 2598 4012
rect 2776 3978 2806 4012
rect 2568 3910 2598 3944
rect 2776 3910 2806 3944
rect 2568 3842 2598 3876
rect 2776 3842 2806 3876
rect 2568 3774 2598 3808
rect 2776 3774 2806 3808
rect 2568 3706 2598 3740
rect 2776 3706 2806 3740
rect 2568 3638 2598 3672
rect 2776 3638 2806 3672
rect 2568 3570 2598 3604
rect 2776 3570 2806 3604
rect 2568 3502 2598 3536
rect 2776 3502 2806 3536
rect 2568 3434 2598 3468
rect 2776 3434 2806 3468
rect 2568 3366 2598 3400
rect 2776 3366 2806 3400
rect 2568 3298 2598 3332
rect 2776 3298 2806 3332
rect 2568 3230 2598 3264
rect 2776 3230 2806 3264
rect 2568 3162 2598 3196
rect 2776 3162 2806 3196
rect 2568 3080 2598 3128
rect 2632 3080 2742 3092
rect 2776 3080 2806 3128
rect 2568 3040 2806 3080
rect 2568 2574 2598 3040
rect 2776 2574 2806 3040
rect 2568 2535 2806 2574
rect 2568 2501 2598 2535
rect 2632 2501 2670 2535
rect 2704 2501 2742 2535
rect 2776 2501 2806 2535
rect 2568 2461 2806 2501
rect 2568 2449 2670 2461
rect 2704 2449 2806 2461
rect 2568 2445 2598 2449
rect 2776 2445 2806 2449
rect 2568 2377 2598 2411
rect 2776 2377 2806 2411
rect 2568 2309 2598 2343
rect 2776 2309 2806 2343
rect 2568 2241 2598 2275
rect 2776 2241 2806 2275
rect 2568 2173 2598 2207
rect 2776 2173 2806 2207
rect 2568 2105 2598 2139
rect 2776 2105 2806 2139
rect 2568 2037 2598 2071
rect 2776 2037 2806 2071
rect 2568 1969 2598 2003
rect 2776 1969 2806 2003
rect 2568 1901 2598 1935
rect 2776 1901 2806 1935
rect 2568 1833 2598 1867
rect 2776 1833 2806 1867
rect 2568 1765 2598 1799
rect 2776 1765 2806 1799
rect 2568 1697 2598 1731
rect 2776 1697 2806 1731
rect 2568 1629 2598 1663
rect 2776 1629 2806 1663
rect 2568 1561 2598 1595
rect 2776 1561 2806 1595
rect 2568 1479 2598 1527
rect 2632 1479 2742 1491
rect 2776 1479 2806 1527
rect 2568 1464 2806 1479
rect 2908 3010 3028 4106
rect 3338 4388 3345 4494
rect 3451 4388 3458 4494
rect 3338 4214 3458 4388
rect 3338 4180 3381 4214
rect 3415 4180 3458 4214
rect 3338 4140 3458 4180
rect 3338 4106 3381 4140
rect 3415 4106 3458 4140
rect 2908 2976 2951 3010
rect 2985 2976 3028 3010
rect 2908 2932 3028 2976
rect 2908 2898 2951 2932
rect 2985 2898 3028 2932
rect 2908 2854 3028 2898
rect 2908 2820 2951 2854
rect 2985 2820 3028 2854
rect 2908 2776 3028 2820
rect 2908 2742 2951 2776
rect 2985 2742 3028 2776
rect 2908 2697 3028 2742
rect 2908 2663 2951 2697
rect 2985 2663 3028 2697
rect 2908 2618 3028 2663
rect 2908 2584 2951 2618
rect 2985 2584 3028 2618
rect 2908 2539 3028 2584
rect 2908 2505 2951 2539
rect 2985 2505 3028 2539
rect 2346 1375 2389 1409
rect 2423 1375 2466 1409
rect 2346 1335 2466 1375
rect 2346 1301 2389 1335
rect 2423 1301 2466 1335
rect 2346 1285 2466 1301
rect 2908 1409 3028 2505
rect 3093 4028 3094 4062
rect 3128 4046 3166 4062
rect 3128 4028 3130 4046
rect 3093 4012 3130 4028
rect 3164 4028 3166 4046
rect 3200 4046 3238 4062
rect 3200 4028 3202 4046
rect 3164 4012 3202 4028
rect 3236 4028 3238 4046
rect 3272 4028 3273 4062
rect 3236 4012 3273 4028
rect 3093 3988 3273 4012
rect 3093 3954 3094 3988
rect 3128 3978 3166 3988
rect 3128 3954 3130 3978
rect 3093 3944 3130 3954
rect 3164 3954 3166 3978
rect 3200 3978 3238 3988
rect 3200 3954 3202 3978
rect 3164 3944 3202 3954
rect 3236 3954 3238 3978
rect 3272 3954 3273 3988
rect 3236 3944 3273 3954
rect 3093 3914 3273 3944
rect 3093 3880 3094 3914
rect 3128 3910 3166 3914
rect 3128 3880 3130 3910
rect 3093 3876 3130 3880
rect 3164 3880 3166 3910
rect 3200 3910 3238 3914
rect 3200 3880 3202 3910
rect 3164 3876 3202 3880
rect 3236 3880 3238 3910
rect 3272 3880 3273 3914
rect 3236 3876 3273 3880
rect 3093 3842 3273 3876
rect 3093 3840 3130 3842
rect 3093 3806 3094 3840
rect 3128 3808 3130 3840
rect 3164 3840 3202 3842
rect 3164 3808 3166 3840
rect 3128 3806 3166 3808
rect 3200 3808 3202 3840
rect 3236 3840 3273 3842
rect 3236 3808 3238 3840
rect 3200 3806 3238 3808
rect 3272 3806 3273 3840
rect 3093 3774 3273 3806
rect 3093 3766 3130 3774
rect 3093 3732 3094 3766
rect 3128 3740 3130 3766
rect 3164 3766 3202 3774
rect 3164 3740 3166 3766
rect 3128 3732 3166 3740
rect 3200 3740 3202 3766
rect 3236 3766 3273 3774
rect 3236 3740 3238 3766
rect 3200 3732 3238 3740
rect 3272 3732 3273 3766
rect 3093 3706 3273 3732
rect 3093 3692 3130 3706
rect 3093 3658 3094 3692
rect 3128 3672 3130 3692
rect 3164 3692 3202 3706
rect 3164 3672 3166 3692
rect 3128 3658 3166 3672
rect 3200 3672 3202 3692
rect 3236 3692 3273 3706
rect 3236 3672 3238 3692
rect 3200 3658 3238 3672
rect 3272 3658 3273 3692
rect 3093 3638 3273 3658
rect 3093 3618 3130 3638
rect 3093 3584 3094 3618
rect 3128 3604 3130 3618
rect 3164 3618 3202 3638
rect 3164 3604 3166 3618
rect 3128 3584 3166 3604
rect 3200 3604 3202 3618
rect 3236 3618 3273 3638
rect 3236 3604 3238 3618
rect 3200 3584 3238 3604
rect 3272 3584 3273 3618
rect 3093 3570 3273 3584
rect 3093 3544 3130 3570
rect 3093 3510 3094 3544
rect 3128 3536 3130 3544
rect 3164 3544 3202 3570
rect 3164 3536 3166 3544
rect 3128 3510 3166 3536
rect 3200 3536 3202 3544
rect 3236 3544 3273 3570
rect 3236 3536 3238 3544
rect 3200 3510 3238 3536
rect 3272 3510 3273 3544
rect 3093 3502 3273 3510
rect 3093 3470 3130 3502
rect 3093 3436 3094 3470
rect 3128 3468 3130 3470
rect 3164 3470 3202 3502
rect 3164 3468 3166 3470
rect 3128 3436 3166 3468
rect 3200 3468 3202 3470
rect 3236 3470 3273 3502
rect 3236 3468 3238 3470
rect 3200 3436 3238 3468
rect 3272 3436 3273 3470
rect 3093 3434 3273 3436
rect 3093 3400 3130 3434
rect 3164 3400 3202 3434
rect 3236 3400 3273 3434
rect 3093 3396 3273 3400
rect 3093 3362 3094 3396
rect 3128 3366 3166 3396
rect 3128 3362 3130 3366
rect 3093 3332 3130 3362
rect 3164 3362 3166 3366
rect 3200 3366 3238 3396
rect 3200 3362 3202 3366
rect 3164 3332 3202 3362
rect 3236 3362 3238 3366
rect 3272 3362 3273 3396
rect 3236 3332 3273 3362
rect 3093 3322 3273 3332
rect 3093 3288 3094 3322
rect 3128 3298 3166 3322
rect 3128 3288 3130 3298
rect 3093 3264 3130 3288
rect 3164 3288 3166 3298
rect 3200 3298 3238 3322
rect 3200 3288 3202 3298
rect 3164 3264 3202 3288
rect 3236 3288 3238 3298
rect 3272 3288 3273 3322
rect 3236 3264 3273 3288
rect 3093 3248 3273 3264
rect 3093 3214 3094 3248
rect 3128 3230 3166 3248
rect 3128 3214 3130 3230
rect 3093 3196 3130 3214
rect 3164 3214 3166 3230
rect 3200 3230 3238 3248
rect 3200 3214 3202 3230
rect 3164 3196 3202 3214
rect 3236 3214 3238 3230
rect 3272 3214 3273 3248
rect 3236 3196 3273 3214
rect 3093 3174 3273 3196
rect 3093 3140 3094 3174
rect 3128 3162 3166 3174
rect 3128 3140 3130 3162
rect 3093 3128 3130 3140
rect 3164 3140 3166 3162
rect 3200 3162 3238 3174
rect 3200 3140 3202 3162
rect 3164 3128 3202 3140
rect 3236 3140 3238 3162
rect 3272 3140 3273 3174
rect 3236 3128 3273 3140
rect 3093 3100 3273 3128
rect 3093 3066 3094 3100
rect 3128 3066 3166 3100
rect 3200 3066 3238 3100
rect 3272 3066 3273 3100
rect 3093 3026 3273 3066
rect 3093 2992 3094 3026
rect 3128 2992 3166 3026
rect 3200 2992 3238 3026
rect 3272 2992 3273 3026
rect 3093 2952 3273 2992
rect 3093 2918 3094 2952
rect 3128 2918 3166 2952
rect 3200 2918 3238 2952
rect 3272 2918 3273 2952
rect 3093 2878 3273 2918
rect 3093 2844 3094 2878
rect 3128 2844 3166 2878
rect 3200 2844 3238 2878
rect 3272 2844 3273 2878
rect 3093 2804 3273 2844
rect 3093 2770 3094 2804
rect 3128 2770 3166 2804
rect 3200 2770 3238 2804
rect 3272 2770 3273 2804
rect 3093 2730 3273 2770
rect 3093 2696 3094 2730
rect 3128 2696 3166 2730
rect 3200 2696 3238 2730
rect 3272 2696 3273 2730
rect 3093 2656 3273 2696
rect 3093 2622 3094 2656
rect 3128 2622 3166 2656
rect 3200 2622 3238 2656
rect 3272 2622 3273 2656
rect 3093 2582 3273 2622
rect 3093 2548 3094 2582
rect 3128 2548 3166 2582
rect 3200 2548 3238 2582
rect 3272 2548 3273 2582
rect 3093 2508 3273 2548
rect 3093 2474 3094 2508
rect 3128 2474 3166 2508
rect 3200 2474 3238 2508
rect 3272 2474 3273 2508
rect 3093 2445 3273 2474
rect 3093 2434 3130 2445
rect 3093 2400 3094 2434
rect 3128 2411 3130 2434
rect 3164 2434 3202 2445
rect 3164 2411 3166 2434
rect 3128 2400 3166 2411
rect 3200 2411 3202 2434
rect 3236 2434 3273 2445
rect 3236 2411 3238 2434
rect 3200 2400 3238 2411
rect 3272 2400 3273 2434
rect 3093 2377 3273 2400
rect 3093 2360 3130 2377
rect 3093 2326 3094 2360
rect 3128 2343 3130 2360
rect 3164 2360 3202 2377
rect 3164 2343 3166 2360
rect 3128 2326 3166 2343
rect 3200 2343 3202 2360
rect 3236 2360 3273 2377
rect 3236 2343 3238 2360
rect 3200 2326 3238 2343
rect 3272 2326 3273 2360
rect 3093 2309 3273 2326
rect 3093 2286 3130 2309
rect 3093 2252 3094 2286
rect 3128 2275 3130 2286
rect 3164 2286 3202 2309
rect 3164 2275 3166 2286
rect 3128 2252 3166 2275
rect 3200 2275 3202 2286
rect 3236 2286 3273 2309
rect 3236 2275 3238 2286
rect 3200 2252 3238 2275
rect 3272 2252 3273 2286
rect 3093 2241 3273 2252
rect 3093 2212 3130 2241
rect 3093 2178 3094 2212
rect 3128 2207 3130 2212
rect 3164 2212 3202 2241
rect 3164 2207 3166 2212
rect 3128 2178 3166 2207
rect 3200 2207 3202 2212
rect 3236 2212 3273 2241
rect 3236 2207 3238 2212
rect 3200 2178 3238 2207
rect 3272 2178 3273 2212
rect 3093 2173 3273 2178
rect 3093 2139 3130 2173
rect 3164 2139 3202 2173
rect 3236 2139 3273 2173
rect 3093 2138 3273 2139
rect 3093 2104 3094 2138
rect 3128 2105 3166 2138
rect 3128 2104 3130 2105
rect 3093 2071 3130 2104
rect 3164 2104 3166 2105
rect 3200 2105 3238 2138
rect 3200 2104 3202 2105
rect 3164 2071 3202 2104
rect 3236 2104 3238 2105
rect 3272 2104 3273 2138
rect 3236 2071 3273 2104
rect 3093 2064 3273 2071
rect 3093 2030 3094 2064
rect 3128 2037 3166 2064
rect 3128 2030 3130 2037
rect 3093 2003 3130 2030
rect 3164 2030 3166 2037
rect 3200 2037 3238 2064
rect 3200 2030 3202 2037
rect 3164 2003 3202 2030
rect 3236 2030 3238 2037
rect 3272 2030 3273 2064
rect 3236 2003 3273 2030
rect 3093 1990 3273 2003
rect 3093 1956 3094 1990
rect 3128 1969 3166 1990
rect 3128 1956 3130 1969
rect 3093 1935 3130 1956
rect 3164 1956 3166 1969
rect 3200 1969 3238 1990
rect 3200 1956 3202 1969
rect 3164 1935 3202 1956
rect 3236 1956 3238 1969
rect 3272 1956 3273 1990
rect 3236 1935 3273 1956
rect 3093 1916 3273 1935
rect 3093 1882 3094 1916
rect 3128 1901 3166 1916
rect 3128 1882 3130 1901
rect 3093 1867 3130 1882
rect 3164 1882 3166 1901
rect 3200 1901 3238 1916
rect 3200 1882 3202 1901
rect 3164 1867 3202 1882
rect 3236 1882 3238 1901
rect 3272 1882 3273 1916
rect 3236 1867 3273 1882
rect 3093 1842 3273 1867
rect 3093 1808 3094 1842
rect 3128 1833 3166 1842
rect 3128 1808 3130 1833
rect 3093 1799 3130 1808
rect 3164 1808 3166 1833
rect 3200 1833 3238 1842
rect 3200 1808 3202 1833
rect 3164 1799 3202 1808
rect 3236 1808 3238 1833
rect 3272 1808 3273 1842
rect 3236 1799 3273 1808
rect 3093 1768 3273 1799
rect 3093 1734 3094 1768
rect 3128 1765 3166 1768
rect 3128 1734 3130 1765
rect 3093 1731 3130 1734
rect 3164 1734 3166 1765
rect 3200 1765 3238 1768
rect 3200 1734 3202 1765
rect 3164 1731 3202 1734
rect 3236 1734 3238 1765
rect 3272 1734 3273 1768
rect 3236 1731 3273 1734
rect 3093 1697 3273 1731
rect 3093 1694 3130 1697
rect 3093 1660 3094 1694
rect 3128 1663 3130 1694
rect 3164 1694 3202 1697
rect 3164 1663 3166 1694
rect 3128 1660 3166 1663
rect 3200 1663 3202 1694
rect 3236 1694 3273 1697
rect 3236 1663 3238 1694
rect 3200 1660 3238 1663
rect 3272 1660 3273 1694
rect 3093 1629 3273 1660
rect 3093 1620 3130 1629
rect 3093 1586 3094 1620
rect 3128 1595 3130 1620
rect 3164 1620 3202 1629
rect 3164 1595 3166 1620
rect 3128 1586 3166 1595
rect 3200 1595 3202 1620
rect 3236 1620 3273 1629
rect 3236 1595 3238 1620
rect 3200 1586 3238 1595
rect 3272 1586 3273 1620
rect 3093 1561 3273 1586
rect 3093 1545 3130 1561
rect 3093 1511 3094 1545
rect 3128 1527 3130 1545
rect 3164 1545 3202 1561
rect 3164 1527 3166 1545
rect 3128 1511 3166 1527
rect 3200 1527 3202 1545
rect 3236 1545 3273 1561
rect 3236 1527 3238 1545
rect 3200 1511 3238 1527
rect 3272 1511 3273 1545
rect 3338 3010 3458 4106
rect 3900 4388 3907 4494
rect 4013 4388 4020 4494
rect 3900 4214 4020 4388
rect 3900 4180 3943 4214
rect 3977 4180 4020 4214
rect 3900 4140 4020 4180
rect 3900 4106 3943 4140
rect 3977 4106 4020 4140
rect 3338 2976 3381 3010
rect 3415 2976 3458 3010
rect 3338 2932 3458 2976
rect 3338 2898 3381 2932
rect 3415 2898 3458 2932
rect 3338 2854 3458 2898
rect 3338 2820 3381 2854
rect 3415 2820 3458 2854
rect 3338 2776 3458 2820
rect 3338 2742 3381 2776
rect 3415 2742 3458 2776
rect 3338 2697 3458 2742
rect 3338 2663 3381 2697
rect 3415 2663 3458 2697
rect 3338 2618 3458 2663
rect 3338 2584 3381 2618
rect 3415 2584 3458 2618
rect 3338 2539 3458 2584
rect 3338 2505 3381 2539
rect 3415 2505 3458 2539
rect 3130 1491 3236 1511
rect 2908 1375 2951 1409
rect 2985 1375 3028 1409
rect 2908 1335 3028 1375
rect 2908 1301 2951 1335
rect 2985 1301 3028 1335
rect 2908 1285 3028 1301
rect 3338 1409 3458 2505
rect 3560 4050 3662 4062
rect 3696 4050 3798 4062
rect 3560 4046 3590 4050
rect 3768 4046 3798 4050
rect 3560 3978 3590 4012
rect 3768 3978 3798 4012
rect 3560 3910 3590 3944
rect 3768 3910 3798 3944
rect 3560 3842 3590 3876
rect 3768 3842 3798 3876
rect 3560 3774 3590 3808
rect 3768 3774 3798 3808
rect 3560 3706 3590 3740
rect 3768 3706 3798 3740
rect 3560 3638 3590 3672
rect 3768 3638 3798 3672
rect 3560 3570 3590 3604
rect 3768 3570 3798 3604
rect 3560 3502 3590 3536
rect 3768 3502 3798 3536
rect 3560 3434 3590 3468
rect 3768 3434 3798 3468
rect 3560 3366 3590 3400
rect 3768 3366 3798 3400
rect 3560 3298 3590 3332
rect 3768 3298 3798 3332
rect 3560 3230 3590 3264
rect 3768 3230 3798 3264
rect 3560 3162 3590 3196
rect 3768 3162 3798 3196
rect 3560 3080 3590 3128
rect 3624 3080 3734 3092
rect 3768 3080 3798 3128
rect 3560 3040 3798 3080
rect 3560 2574 3590 3040
rect 3768 2574 3798 3040
rect 3560 2535 3798 2574
rect 3560 2501 3590 2535
rect 3624 2501 3662 2535
rect 3696 2501 3734 2535
rect 3768 2501 3798 2535
rect 3560 2461 3798 2501
rect 3560 2449 3662 2461
rect 3696 2449 3798 2461
rect 3560 2445 3590 2449
rect 3768 2445 3798 2449
rect 3560 2377 3590 2411
rect 3768 2377 3798 2411
rect 3560 2309 3590 2343
rect 3768 2309 3798 2343
rect 3560 2241 3590 2275
rect 3768 2241 3798 2275
rect 3560 2173 3590 2207
rect 3768 2173 3798 2207
rect 3560 2105 3590 2139
rect 3768 2105 3798 2139
rect 3560 2037 3590 2071
rect 3768 2037 3798 2071
rect 3560 1969 3590 2003
rect 3768 1969 3798 2003
rect 3560 1901 3590 1935
rect 3768 1901 3798 1935
rect 3560 1833 3590 1867
rect 3768 1833 3798 1867
rect 3560 1765 3590 1799
rect 3768 1765 3798 1799
rect 3560 1697 3590 1731
rect 3768 1697 3798 1731
rect 3560 1629 3590 1663
rect 3768 1629 3798 1663
rect 3560 1561 3590 1595
rect 3768 1561 3798 1595
rect 3560 1479 3590 1527
rect 3624 1479 3734 1491
rect 3768 1479 3798 1527
rect 3560 1464 3798 1479
rect 3900 3010 4020 4106
rect 4330 4388 4337 4494
rect 4443 4388 4450 4494
rect 4330 4214 4450 4388
rect 4330 4180 4373 4214
rect 4407 4180 4450 4214
rect 4330 4140 4450 4180
rect 4330 4106 4373 4140
rect 4407 4106 4450 4140
rect 3900 2976 3943 3010
rect 3977 2976 4020 3010
rect 3900 2932 4020 2976
rect 3900 2898 3943 2932
rect 3977 2898 4020 2932
rect 3900 2854 4020 2898
rect 3900 2820 3943 2854
rect 3977 2820 4020 2854
rect 3900 2776 4020 2820
rect 3900 2742 3943 2776
rect 3977 2742 4020 2776
rect 3900 2697 4020 2742
rect 3900 2663 3943 2697
rect 3977 2663 4020 2697
rect 3900 2618 4020 2663
rect 3900 2584 3943 2618
rect 3977 2584 4020 2618
rect 3900 2539 4020 2584
rect 3900 2505 3943 2539
rect 3977 2505 4020 2539
rect 3338 1375 3381 1409
rect 3415 1375 3458 1409
rect 3338 1335 3458 1375
rect 3338 1301 3381 1335
rect 3415 1301 3458 1335
rect 3338 1285 3458 1301
rect 3900 1409 4020 2505
rect 4085 4028 4086 4062
rect 4120 4046 4158 4062
rect 4120 4028 4122 4046
rect 4085 4012 4122 4028
rect 4156 4028 4158 4046
rect 4192 4046 4230 4062
rect 4192 4028 4194 4046
rect 4156 4012 4194 4028
rect 4228 4028 4230 4046
rect 4264 4028 4265 4062
rect 4228 4012 4265 4028
rect 4085 3988 4265 4012
rect 4085 3954 4086 3988
rect 4120 3978 4158 3988
rect 4120 3954 4122 3978
rect 4085 3944 4122 3954
rect 4156 3954 4158 3978
rect 4192 3978 4230 3988
rect 4192 3954 4194 3978
rect 4156 3944 4194 3954
rect 4228 3954 4230 3978
rect 4264 3954 4265 3988
rect 4228 3944 4265 3954
rect 4085 3914 4265 3944
rect 4085 3880 4086 3914
rect 4120 3910 4158 3914
rect 4120 3880 4122 3910
rect 4085 3876 4122 3880
rect 4156 3880 4158 3910
rect 4192 3910 4230 3914
rect 4192 3880 4194 3910
rect 4156 3876 4194 3880
rect 4228 3880 4230 3910
rect 4264 3880 4265 3914
rect 4228 3876 4265 3880
rect 4085 3842 4265 3876
rect 4085 3840 4122 3842
rect 4085 3806 4086 3840
rect 4120 3808 4122 3840
rect 4156 3840 4194 3842
rect 4156 3808 4158 3840
rect 4120 3806 4158 3808
rect 4192 3808 4194 3840
rect 4228 3840 4265 3842
rect 4228 3808 4230 3840
rect 4192 3806 4230 3808
rect 4264 3806 4265 3840
rect 4085 3774 4265 3806
rect 4085 3766 4122 3774
rect 4085 3732 4086 3766
rect 4120 3740 4122 3766
rect 4156 3766 4194 3774
rect 4156 3740 4158 3766
rect 4120 3732 4158 3740
rect 4192 3740 4194 3766
rect 4228 3766 4265 3774
rect 4228 3740 4230 3766
rect 4192 3732 4230 3740
rect 4264 3732 4265 3766
rect 4085 3706 4265 3732
rect 4085 3692 4122 3706
rect 4085 3658 4086 3692
rect 4120 3672 4122 3692
rect 4156 3692 4194 3706
rect 4156 3672 4158 3692
rect 4120 3658 4158 3672
rect 4192 3672 4194 3692
rect 4228 3692 4265 3706
rect 4228 3672 4230 3692
rect 4192 3658 4230 3672
rect 4264 3658 4265 3692
rect 4085 3638 4265 3658
rect 4085 3618 4122 3638
rect 4085 3584 4086 3618
rect 4120 3604 4122 3618
rect 4156 3618 4194 3638
rect 4156 3604 4158 3618
rect 4120 3584 4158 3604
rect 4192 3604 4194 3618
rect 4228 3618 4265 3638
rect 4228 3604 4230 3618
rect 4192 3584 4230 3604
rect 4264 3584 4265 3618
rect 4085 3570 4265 3584
rect 4085 3544 4122 3570
rect 4085 3510 4086 3544
rect 4120 3536 4122 3544
rect 4156 3544 4194 3570
rect 4156 3536 4158 3544
rect 4120 3510 4158 3536
rect 4192 3536 4194 3544
rect 4228 3544 4265 3570
rect 4228 3536 4230 3544
rect 4192 3510 4230 3536
rect 4264 3510 4265 3544
rect 4085 3502 4265 3510
rect 4085 3470 4122 3502
rect 4085 3436 4086 3470
rect 4120 3468 4122 3470
rect 4156 3470 4194 3502
rect 4156 3468 4158 3470
rect 4120 3436 4158 3468
rect 4192 3468 4194 3470
rect 4228 3470 4265 3502
rect 4228 3468 4230 3470
rect 4192 3436 4230 3468
rect 4264 3436 4265 3470
rect 4085 3434 4265 3436
rect 4085 3400 4122 3434
rect 4156 3400 4194 3434
rect 4228 3400 4265 3434
rect 4085 3396 4265 3400
rect 4085 3362 4086 3396
rect 4120 3366 4158 3396
rect 4120 3362 4122 3366
rect 4085 3332 4122 3362
rect 4156 3362 4158 3366
rect 4192 3366 4230 3396
rect 4192 3362 4194 3366
rect 4156 3332 4194 3362
rect 4228 3362 4230 3366
rect 4264 3362 4265 3396
rect 4228 3332 4265 3362
rect 4085 3322 4265 3332
rect 4085 3288 4086 3322
rect 4120 3298 4158 3322
rect 4120 3288 4122 3298
rect 4085 3264 4122 3288
rect 4156 3288 4158 3298
rect 4192 3298 4230 3322
rect 4192 3288 4194 3298
rect 4156 3264 4194 3288
rect 4228 3288 4230 3298
rect 4264 3288 4265 3322
rect 4228 3264 4265 3288
rect 4085 3248 4265 3264
rect 4085 3214 4086 3248
rect 4120 3230 4158 3248
rect 4120 3214 4122 3230
rect 4085 3196 4122 3214
rect 4156 3214 4158 3230
rect 4192 3230 4230 3248
rect 4192 3214 4194 3230
rect 4156 3196 4194 3214
rect 4228 3214 4230 3230
rect 4264 3214 4265 3248
rect 4228 3196 4265 3214
rect 4085 3174 4265 3196
rect 4085 3140 4086 3174
rect 4120 3162 4158 3174
rect 4120 3140 4122 3162
rect 4085 3128 4122 3140
rect 4156 3140 4158 3162
rect 4192 3162 4230 3174
rect 4192 3140 4194 3162
rect 4156 3128 4194 3140
rect 4228 3140 4230 3162
rect 4264 3140 4265 3174
rect 4228 3128 4265 3140
rect 4085 3100 4265 3128
rect 4085 3066 4086 3100
rect 4120 3066 4158 3100
rect 4192 3066 4230 3100
rect 4264 3066 4265 3100
rect 4085 3026 4265 3066
rect 4085 2992 4086 3026
rect 4120 2992 4158 3026
rect 4192 2992 4230 3026
rect 4264 2992 4265 3026
rect 4085 2952 4265 2992
rect 4085 2918 4086 2952
rect 4120 2918 4158 2952
rect 4192 2918 4230 2952
rect 4264 2918 4265 2952
rect 4085 2878 4265 2918
rect 4085 2844 4086 2878
rect 4120 2844 4158 2878
rect 4192 2844 4230 2878
rect 4264 2844 4265 2878
rect 4085 2804 4265 2844
rect 4085 2770 4086 2804
rect 4120 2770 4158 2804
rect 4192 2770 4230 2804
rect 4264 2770 4265 2804
rect 4085 2730 4265 2770
rect 4085 2696 4086 2730
rect 4120 2696 4158 2730
rect 4192 2696 4230 2730
rect 4264 2696 4265 2730
rect 4085 2656 4265 2696
rect 4085 2622 4086 2656
rect 4120 2622 4158 2656
rect 4192 2622 4230 2656
rect 4264 2622 4265 2656
rect 4085 2582 4265 2622
rect 4085 2548 4086 2582
rect 4120 2548 4158 2582
rect 4192 2548 4230 2582
rect 4264 2548 4265 2582
rect 4085 2508 4265 2548
rect 4085 2474 4086 2508
rect 4120 2474 4158 2508
rect 4192 2474 4230 2508
rect 4264 2474 4265 2508
rect 4085 2445 4265 2474
rect 4085 2434 4122 2445
rect 4085 2400 4086 2434
rect 4120 2411 4122 2434
rect 4156 2434 4194 2445
rect 4156 2411 4158 2434
rect 4120 2400 4158 2411
rect 4192 2411 4194 2434
rect 4228 2434 4265 2445
rect 4228 2411 4230 2434
rect 4192 2400 4230 2411
rect 4264 2400 4265 2434
rect 4085 2377 4265 2400
rect 4085 2360 4122 2377
rect 4085 2326 4086 2360
rect 4120 2343 4122 2360
rect 4156 2360 4194 2377
rect 4156 2343 4158 2360
rect 4120 2326 4158 2343
rect 4192 2343 4194 2360
rect 4228 2360 4265 2377
rect 4228 2343 4230 2360
rect 4192 2326 4230 2343
rect 4264 2326 4265 2360
rect 4085 2309 4265 2326
rect 4085 2286 4122 2309
rect 4085 2252 4086 2286
rect 4120 2275 4122 2286
rect 4156 2286 4194 2309
rect 4156 2275 4158 2286
rect 4120 2252 4158 2275
rect 4192 2275 4194 2286
rect 4228 2286 4265 2309
rect 4228 2275 4230 2286
rect 4192 2252 4230 2275
rect 4264 2252 4265 2286
rect 4085 2241 4265 2252
rect 4085 2212 4122 2241
rect 4085 2178 4086 2212
rect 4120 2207 4122 2212
rect 4156 2212 4194 2241
rect 4156 2207 4158 2212
rect 4120 2178 4158 2207
rect 4192 2207 4194 2212
rect 4228 2212 4265 2241
rect 4228 2207 4230 2212
rect 4192 2178 4230 2207
rect 4264 2178 4265 2212
rect 4085 2173 4265 2178
rect 4085 2139 4122 2173
rect 4156 2139 4194 2173
rect 4228 2139 4265 2173
rect 4085 2138 4265 2139
rect 4085 2104 4086 2138
rect 4120 2105 4158 2138
rect 4120 2104 4122 2105
rect 4085 2071 4122 2104
rect 4156 2104 4158 2105
rect 4192 2105 4230 2138
rect 4192 2104 4194 2105
rect 4156 2071 4194 2104
rect 4228 2104 4230 2105
rect 4264 2104 4265 2138
rect 4228 2071 4265 2104
rect 4085 2064 4265 2071
rect 4085 2030 4086 2064
rect 4120 2037 4158 2064
rect 4120 2030 4122 2037
rect 4085 2003 4122 2030
rect 4156 2030 4158 2037
rect 4192 2037 4230 2064
rect 4192 2030 4194 2037
rect 4156 2003 4194 2030
rect 4228 2030 4230 2037
rect 4264 2030 4265 2064
rect 4228 2003 4265 2030
rect 4085 1990 4265 2003
rect 4085 1956 4086 1990
rect 4120 1969 4158 1990
rect 4120 1956 4122 1969
rect 4085 1935 4122 1956
rect 4156 1956 4158 1969
rect 4192 1969 4230 1990
rect 4192 1956 4194 1969
rect 4156 1935 4194 1956
rect 4228 1956 4230 1969
rect 4264 1956 4265 1990
rect 4228 1935 4265 1956
rect 4085 1916 4265 1935
rect 4085 1882 4086 1916
rect 4120 1901 4158 1916
rect 4120 1882 4122 1901
rect 4085 1867 4122 1882
rect 4156 1882 4158 1901
rect 4192 1901 4230 1916
rect 4192 1882 4194 1901
rect 4156 1867 4194 1882
rect 4228 1882 4230 1901
rect 4264 1882 4265 1916
rect 4228 1867 4265 1882
rect 4085 1842 4265 1867
rect 4085 1808 4086 1842
rect 4120 1833 4158 1842
rect 4120 1808 4122 1833
rect 4085 1799 4122 1808
rect 4156 1808 4158 1833
rect 4192 1833 4230 1842
rect 4192 1808 4194 1833
rect 4156 1799 4194 1808
rect 4228 1808 4230 1833
rect 4264 1808 4265 1842
rect 4228 1799 4265 1808
rect 4085 1768 4265 1799
rect 4085 1734 4086 1768
rect 4120 1765 4158 1768
rect 4120 1734 4122 1765
rect 4085 1731 4122 1734
rect 4156 1734 4158 1765
rect 4192 1765 4230 1768
rect 4192 1734 4194 1765
rect 4156 1731 4194 1734
rect 4228 1734 4230 1765
rect 4264 1734 4265 1768
rect 4228 1731 4265 1734
rect 4085 1697 4265 1731
rect 4085 1694 4122 1697
rect 4085 1660 4086 1694
rect 4120 1663 4122 1694
rect 4156 1694 4194 1697
rect 4156 1663 4158 1694
rect 4120 1660 4158 1663
rect 4192 1663 4194 1694
rect 4228 1694 4265 1697
rect 4228 1663 4230 1694
rect 4192 1660 4230 1663
rect 4264 1660 4265 1694
rect 4085 1629 4265 1660
rect 4085 1620 4122 1629
rect 4085 1586 4086 1620
rect 4120 1595 4122 1620
rect 4156 1620 4194 1629
rect 4156 1595 4158 1620
rect 4120 1586 4158 1595
rect 4192 1595 4194 1620
rect 4228 1620 4265 1629
rect 4228 1595 4230 1620
rect 4192 1586 4230 1595
rect 4264 1586 4265 1620
rect 4085 1561 4265 1586
rect 4085 1545 4122 1561
rect 4085 1511 4086 1545
rect 4120 1527 4122 1545
rect 4156 1545 4194 1561
rect 4156 1527 4158 1545
rect 4120 1511 4158 1527
rect 4192 1527 4194 1545
rect 4228 1545 4265 1561
rect 4228 1527 4230 1545
rect 4192 1511 4230 1527
rect 4264 1511 4265 1545
rect 4330 3010 4450 4106
rect 4892 4388 4899 4494
rect 5005 4388 5012 4494
rect 4892 4214 5012 4388
rect 4892 4180 4935 4214
rect 4969 4180 5012 4214
rect 4892 4140 5012 4180
rect 4892 4106 4935 4140
rect 4969 4106 5012 4140
rect 4330 2976 4373 3010
rect 4407 2976 4450 3010
rect 4330 2932 4450 2976
rect 4330 2898 4373 2932
rect 4407 2898 4450 2932
rect 4330 2854 4450 2898
rect 4330 2820 4373 2854
rect 4407 2820 4450 2854
rect 4330 2776 4450 2820
rect 4330 2742 4373 2776
rect 4407 2742 4450 2776
rect 4330 2697 4450 2742
rect 4330 2663 4373 2697
rect 4407 2663 4450 2697
rect 4330 2618 4450 2663
rect 4330 2584 4373 2618
rect 4407 2584 4450 2618
rect 4330 2539 4450 2584
rect 4330 2505 4373 2539
rect 4407 2505 4450 2539
rect 4122 1491 4228 1511
rect 3900 1375 3943 1409
rect 3977 1375 4020 1409
rect 3900 1335 4020 1375
rect 3900 1301 3943 1335
rect 3977 1301 4020 1335
rect 3900 1285 4020 1301
rect 4330 1409 4450 2505
rect 4552 4050 4654 4062
rect 4688 4050 4790 4062
rect 4552 4046 4582 4050
rect 4760 4046 4790 4050
rect 4552 3978 4582 4012
rect 4760 3978 4790 4012
rect 4552 3910 4582 3944
rect 4760 3910 4790 3944
rect 4552 3842 4582 3876
rect 4760 3842 4790 3876
rect 4552 3774 4582 3808
rect 4760 3774 4790 3808
rect 4552 3706 4582 3740
rect 4760 3706 4790 3740
rect 4552 3638 4582 3672
rect 4760 3638 4790 3672
rect 4552 3570 4582 3604
rect 4760 3570 4790 3604
rect 4552 3502 4582 3536
rect 4760 3502 4790 3536
rect 4552 3434 4582 3468
rect 4760 3434 4790 3468
rect 4552 3366 4582 3400
rect 4760 3366 4790 3400
rect 4552 3298 4582 3332
rect 4760 3298 4790 3332
rect 4552 3230 4582 3264
rect 4760 3230 4790 3264
rect 4552 3162 4582 3196
rect 4760 3162 4790 3196
rect 4552 3080 4582 3128
rect 4616 3080 4726 3092
rect 4760 3080 4790 3128
rect 4552 3040 4790 3080
rect 4552 2574 4582 3040
rect 4760 2574 4790 3040
rect 4552 2535 4790 2574
rect 4552 2501 4582 2535
rect 4616 2501 4654 2535
rect 4688 2501 4726 2535
rect 4760 2501 4790 2535
rect 4552 2461 4790 2501
rect 4552 2449 4654 2461
rect 4688 2449 4790 2461
rect 4552 2445 4582 2449
rect 4760 2445 4790 2449
rect 4552 2377 4582 2411
rect 4760 2377 4790 2411
rect 4552 2309 4582 2343
rect 4760 2309 4790 2343
rect 4552 2241 4582 2275
rect 4760 2241 4790 2275
rect 4552 2173 4582 2207
rect 4760 2173 4790 2207
rect 4552 2105 4582 2139
rect 4760 2105 4790 2139
rect 4552 2037 4582 2071
rect 4760 2037 4790 2071
rect 4552 1969 4582 2003
rect 4760 1969 4790 2003
rect 4552 1901 4582 1935
rect 4760 1901 4790 1935
rect 4552 1833 4582 1867
rect 4760 1833 4790 1867
rect 4552 1765 4582 1799
rect 4760 1765 4790 1799
rect 4552 1697 4582 1731
rect 4760 1697 4790 1731
rect 4552 1629 4582 1663
rect 4760 1629 4790 1663
rect 4552 1561 4582 1595
rect 4760 1561 4790 1595
rect 4552 1479 4582 1527
rect 4616 1479 4726 1491
rect 4760 1479 4790 1527
rect 4552 1464 4790 1479
rect 4892 3010 5012 4106
rect 5322 4388 5329 4494
rect 5435 4388 5442 4494
rect 5322 4214 5442 4388
rect 5322 4180 5365 4214
rect 5399 4180 5442 4214
rect 5322 4140 5442 4180
rect 5322 4106 5365 4140
rect 5399 4106 5442 4140
rect 4892 2976 4935 3010
rect 4969 2976 5012 3010
rect 4892 2932 5012 2976
rect 4892 2898 4935 2932
rect 4969 2898 5012 2932
rect 4892 2854 5012 2898
rect 4892 2820 4935 2854
rect 4969 2820 5012 2854
rect 4892 2776 5012 2820
rect 4892 2742 4935 2776
rect 4969 2742 5012 2776
rect 4892 2697 5012 2742
rect 4892 2663 4935 2697
rect 4969 2663 5012 2697
rect 4892 2618 5012 2663
rect 4892 2584 4935 2618
rect 4969 2584 5012 2618
rect 4892 2539 5012 2584
rect 4892 2505 4935 2539
rect 4969 2505 5012 2539
rect 4330 1375 4373 1409
rect 4407 1375 4450 1409
rect 4330 1335 4450 1375
rect 4330 1301 4373 1335
rect 4407 1301 4450 1335
rect 4330 1285 4450 1301
rect 4892 1409 5012 2505
rect 5077 4028 5078 4062
rect 5112 4046 5150 4062
rect 5112 4028 5114 4046
rect 5077 4012 5114 4028
rect 5148 4028 5150 4046
rect 5184 4046 5222 4062
rect 5184 4028 5186 4046
rect 5148 4012 5186 4028
rect 5220 4028 5222 4046
rect 5256 4028 5257 4062
rect 5220 4012 5257 4028
rect 5077 3988 5257 4012
rect 5077 3954 5078 3988
rect 5112 3978 5150 3988
rect 5112 3954 5114 3978
rect 5077 3944 5114 3954
rect 5148 3954 5150 3978
rect 5184 3978 5222 3988
rect 5184 3954 5186 3978
rect 5148 3944 5186 3954
rect 5220 3954 5222 3978
rect 5256 3954 5257 3988
rect 5220 3944 5257 3954
rect 5077 3914 5257 3944
rect 5077 3880 5078 3914
rect 5112 3910 5150 3914
rect 5112 3880 5114 3910
rect 5077 3876 5114 3880
rect 5148 3880 5150 3910
rect 5184 3910 5222 3914
rect 5184 3880 5186 3910
rect 5148 3876 5186 3880
rect 5220 3880 5222 3910
rect 5256 3880 5257 3914
rect 5220 3876 5257 3880
rect 5077 3842 5257 3876
rect 5077 3840 5114 3842
rect 5077 3806 5078 3840
rect 5112 3808 5114 3840
rect 5148 3840 5186 3842
rect 5148 3808 5150 3840
rect 5112 3806 5150 3808
rect 5184 3808 5186 3840
rect 5220 3840 5257 3842
rect 5220 3808 5222 3840
rect 5184 3806 5222 3808
rect 5256 3806 5257 3840
rect 5077 3774 5257 3806
rect 5077 3766 5114 3774
rect 5077 3732 5078 3766
rect 5112 3740 5114 3766
rect 5148 3766 5186 3774
rect 5148 3740 5150 3766
rect 5112 3732 5150 3740
rect 5184 3740 5186 3766
rect 5220 3766 5257 3774
rect 5220 3740 5222 3766
rect 5184 3732 5222 3740
rect 5256 3732 5257 3766
rect 5077 3706 5257 3732
rect 5077 3692 5114 3706
rect 5077 3658 5078 3692
rect 5112 3672 5114 3692
rect 5148 3692 5186 3706
rect 5148 3672 5150 3692
rect 5112 3658 5150 3672
rect 5184 3672 5186 3692
rect 5220 3692 5257 3706
rect 5220 3672 5222 3692
rect 5184 3658 5222 3672
rect 5256 3658 5257 3692
rect 5077 3638 5257 3658
rect 5077 3618 5114 3638
rect 5077 3584 5078 3618
rect 5112 3604 5114 3618
rect 5148 3618 5186 3638
rect 5148 3604 5150 3618
rect 5112 3584 5150 3604
rect 5184 3604 5186 3618
rect 5220 3618 5257 3638
rect 5220 3604 5222 3618
rect 5184 3584 5222 3604
rect 5256 3584 5257 3618
rect 5077 3570 5257 3584
rect 5077 3544 5114 3570
rect 5077 3510 5078 3544
rect 5112 3536 5114 3544
rect 5148 3544 5186 3570
rect 5148 3536 5150 3544
rect 5112 3510 5150 3536
rect 5184 3536 5186 3544
rect 5220 3544 5257 3570
rect 5220 3536 5222 3544
rect 5184 3510 5222 3536
rect 5256 3510 5257 3544
rect 5077 3502 5257 3510
rect 5077 3470 5114 3502
rect 5077 3436 5078 3470
rect 5112 3468 5114 3470
rect 5148 3470 5186 3502
rect 5148 3468 5150 3470
rect 5112 3436 5150 3468
rect 5184 3468 5186 3470
rect 5220 3470 5257 3502
rect 5220 3468 5222 3470
rect 5184 3436 5222 3468
rect 5256 3436 5257 3470
rect 5077 3434 5257 3436
rect 5077 3400 5114 3434
rect 5148 3400 5186 3434
rect 5220 3400 5257 3434
rect 5077 3396 5257 3400
rect 5077 3362 5078 3396
rect 5112 3366 5150 3396
rect 5112 3362 5114 3366
rect 5077 3332 5114 3362
rect 5148 3362 5150 3366
rect 5184 3366 5222 3396
rect 5184 3362 5186 3366
rect 5148 3332 5186 3362
rect 5220 3362 5222 3366
rect 5256 3362 5257 3396
rect 5220 3332 5257 3362
rect 5077 3322 5257 3332
rect 5077 3288 5078 3322
rect 5112 3298 5150 3322
rect 5112 3288 5114 3298
rect 5077 3264 5114 3288
rect 5148 3288 5150 3298
rect 5184 3298 5222 3322
rect 5184 3288 5186 3298
rect 5148 3264 5186 3288
rect 5220 3288 5222 3298
rect 5256 3288 5257 3322
rect 5220 3264 5257 3288
rect 5077 3248 5257 3264
rect 5077 3214 5078 3248
rect 5112 3230 5150 3248
rect 5112 3214 5114 3230
rect 5077 3196 5114 3214
rect 5148 3214 5150 3230
rect 5184 3230 5222 3248
rect 5184 3214 5186 3230
rect 5148 3196 5186 3214
rect 5220 3214 5222 3230
rect 5256 3214 5257 3248
rect 5220 3196 5257 3214
rect 5077 3174 5257 3196
rect 5077 3140 5078 3174
rect 5112 3162 5150 3174
rect 5112 3140 5114 3162
rect 5077 3128 5114 3140
rect 5148 3140 5150 3162
rect 5184 3162 5222 3174
rect 5184 3140 5186 3162
rect 5148 3128 5186 3140
rect 5220 3140 5222 3162
rect 5256 3140 5257 3174
rect 5220 3128 5257 3140
rect 5077 3100 5257 3128
rect 5077 3066 5078 3100
rect 5112 3066 5150 3100
rect 5184 3066 5222 3100
rect 5256 3066 5257 3100
rect 5077 3026 5257 3066
rect 5077 2992 5078 3026
rect 5112 2992 5150 3026
rect 5184 2992 5222 3026
rect 5256 2992 5257 3026
rect 5077 2952 5257 2992
rect 5077 2918 5078 2952
rect 5112 2918 5150 2952
rect 5184 2918 5222 2952
rect 5256 2918 5257 2952
rect 5077 2878 5257 2918
rect 5077 2844 5078 2878
rect 5112 2844 5150 2878
rect 5184 2844 5222 2878
rect 5256 2844 5257 2878
rect 5077 2804 5257 2844
rect 5077 2770 5078 2804
rect 5112 2770 5150 2804
rect 5184 2770 5222 2804
rect 5256 2770 5257 2804
rect 5077 2730 5257 2770
rect 5077 2696 5078 2730
rect 5112 2696 5150 2730
rect 5184 2696 5222 2730
rect 5256 2696 5257 2730
rect 5077 2656 5257 2696
rect 5077 2622 5078 2656
rect 5112 2622 5150 2656
rect 5184 2622 5222 2656
rect 5256 2622 5257 2656
rect 5077 2582 5257 2622
rect 5077 2548 5078 2582
rect 5112 2548 5150 2582
rect 5184 2548 5222 2582
rect 5256 2548 5257 2582
rect 5077 2508 5257 2548
rect 5077 2474 5078 2508
rect 5112 2474 5150 2508
rect 5184 2474 5222 2508
rect 5256 2474 5257 2508
rect 5077 2445 5257 2474
rect 5077 2434 5114 2445
rect 5077 2400 5078 2434
rect 5112 2411 5114 2434
rect 5148 2434 5186 2445
rect 5148 2411 5150 2434
rect 5112 2400 5150 2411
rect 5184 2411 5186 2434
rect 5220 2434 5257 2445
rect 5220 2411 5222 2434
rect 5184 2400 5222 2411
rect 5256 2400 5257 2434
rect 5077 2377 5257 2400
rect 5077 2360 5114 2377
rect 5077 2326 5078 2360
rect 5112 2343 5114 2360
rect 5148 2360 5186 2377
rect 5148 2343 5150 2360
rect 5112 2326 5150 2343
rect 5184 2343 5186 2360
rect 5220 2360 5257 2377
rect 5220 2343 5222 2360
rect 5184 2326 5222 2343
rect 5256 2326 5257 2360
rect 5077 2309 5257 2326
rect 5077 2286 5114 2309
rect 5077 2252 5078 2286
rect 5112 2275 5114 2286
rect 5148 2286 5186 2309
rect 5148 2275 5150 2286
rect 5112 2252 5150 2275
rect 5184 2275 5186 2286
rect 5220 2286 5257 2309
rect 5220 2275 5222 2286
rect 5184 2252 5222 2275
rect 5256 2252 5257 2286
rect 5077 2241 5257 2252
rect 5077 2212 5114 2241
rect 5077 2178 5078 2212
rect 5112 2207 5114 2212
rect 5148 2212 5186 2241
rect 5148 2207 5150 2212
rect 5112 2178 5150 2207
rect 5184 2207 5186 2212
rect 5220 2212 5257 2241
rect 5220 2207 5222 2212
rect 5184 2178 5222 2207
rect 5256 2178 5257 2212
rect 5077 2173 5257 2178
rect 5077 2139 5114 2173
rect 5148 2139 5186 2173
rect 5220 2139 5257 2173
rect 5077 2138 5257 2139
rect 5077 2104 5078 2138
rect 5112 2105 5150 2138
rect 5112 2104 5114 2105
rect 5077 2071 5114 2104
rect 5148 2104 5150 2105
rect 5184 2105 5222 2138
rect 5184 2104 5186 2105
rect 5148 2071 5186 2104
rect 5220 2104 5222 2105
rect 5256 2104 5257 2138
rect 5220 2071 5257 2104
rect 5077 2064 5257 2071
rect 5077 2030 5078 2064
rect 5112 2037 5150 2064
rect 5112 2030 5114 2037
rect 5077 2003 5114 2030
rect 5148 2030 5150 2037
rect 5184 2037 5222 2064
rect 5184 2030 5186 2037
rect 5148 2003 5186 2030
rect 5220 2030 5222 2037
rect 5256 2030 5257 2064
rect 5220 2003 5257 2030
rect 5077 1990 5257 2003
rect 5077 1956 5078 1990
rect 5112 1969 5150 1990
rect 5112 1956 5114 1969
rect 5077 1935 5114 1956
rect 5148 1956 5150 1969
rect 5184 1969 5222 1990
rect 5184 1956 5186 1969
rect 5148 1935 5186 1956
rect 5220 1956 5222 1969
rect 5256 1956 5257 1990
rect 5220 1935 5257 1956
rect 5077 1916 5257 1935
rect 5077 1882 5078 1916
rect 5112 1901 5150 1916
rect 5112 1882 5114 1901
rect 5077 1867 5114 1882
rect 5148 1882 5150 1901
rect 5184 1901 5222 1916
rect 5184 1882 5186 1901
rect 5148 1867 5186 1882
rect 5220 1882 5222 1901
rect 5256 1882 5257 1916
rect 5220 1867 5257 1882
rect 5077 1842 5257 1867
rect 5077 1808 5078 1842
rect 5112 1833 5150 1842
rect 5112 1808 5114 1833
rect 5077 1799 5114 1808
rect 5148 1808 5150 1833
rect 5184 1833 5222 1842
rect 5184 1808 5186 1833
rect 5148 1799 5186 1808
rect 5220 1808 5222 1833
rect 5256 1808 5257 1842
rect 5220 1799 5257 1808
rect 5077 1768 5257 1799
rect 5077 1734 5078 1768
rect 5112 1765 5150 1768
rect 5112 1734 5114 1765
rect 5077 1731 5114 1734
rect 5148 1734 5150 1765
rect 5184 1765 5222 1768
rect 5184 1734 5186 1765
rect 5148 1731 5186 1734
rect 5220 1734 5222 1765
rect 5256 1734 5257 1768
rect 5220 1731 5257 1734
rect 5077 1697 5257 1731
rect 5077 1694 5114 1697
rect 5077 1660 5078 1694
rect 5112 1663 5114 1694
rect 5148 1694 5186 1697
rect 5148 1663 5150 1694
rect 5112 1660 5150 1663
rect 5184 1663 5186 1694
rect 5220 1694 5257 1697
rect 5220 1663 5222 1694
rect 5184 1660 5222 1663
rect 5256 1660 5257 1694
rect 5077 1629 5257 1660
rect 5077 1620 5114 1629
rect 5077 1586 5078 1620
rect 5112 1595 5114 1620
rect 5148 1620 5186 1629
rect 5148 1595 5150 1620
rect 5112 1586 5150 1595
rect 5184 1595 5186 1620
rect 5220 1620 5257 1629
rect 5220 1595 5222 1620
rect 5184 1586 5222 1595
rect 5256 1586 5257 1620
rect 5077 1561 5257 1586
rect 5077 1545 5114 1561
rect 5077 1511 5078 1545
rect 5112 1527 5114 1545
rect 5148 1545 5186 1561
rect 5148 1527 5150 1545
rect 5112 1511 5150 1527
rect 5184 1527 5186 1545
rect 5220 1545 5257 1561
rect 5220 1527 5222 1545
rect 5184 1511 5222 1527
rect 5256 1511 5257 1545
rect 5322 3010 5442 4106
rect 5884 4388 5891 4494
rect 5997 4388 6004 4494
rect 5884 4214 6004 4388
rect 5884 4180 5927 4214
rect 5961 4180 6004 4214
rect 5884 4140 6004 4180
rect 5884 4106 5927 4140
rect 5961 4106 6004 4140
rect 5322 2976 5365 3010
rect 5399 2976 5442 3010
rect 5322 2932 5442 2976
rect 5322 2898 5365 2932
rect 5399 2898 5442 2932
rect 5322 2854 5442 2898
rect 5322 2820 5365 2854
rect 5399 2820 5442 2854
rect 5322 2776 5442 2820
rect 5322 2742 5365 2776
rect 5399 2742 5442 2776
rect 5322 2697 5442 2742
rect 5322 2663 5365 2697
rect 5399 2663 5442 2697
rect 5322 2618 5442 2663
rect 5322 2584 5365 2618
rect 5399 2584 5442 2618
rect 5322 2539 5442 2584
rect 5322 2505 5365 2539
rect 5399 2505 5442 2539
rect 5114 1491 5220 1511
rect 4892 1375 4935 1409
rect 4969 1375 5012 1409
rect 4892 1335 5012 1375
rect 4892 1301 4935 1335
rect 4969 1301 5012 1335
rect 4892 1285 5012 1301
rect 5322 1409 5442 2505
rect 5544 4050 5646 4062
rect 5680 4050 5782 4062
rect 5544 4046 5574 4050
rect 5752 4046 5782 4050
rect 5544 3978 5574 4012
rect 5752 3978 5782 4012
rect 5544 3910 5574 3944
rect 5752 3910 5782 3944
rect 5544 3842 5574 3876
rect 5752 3842 5782 3876
rect 5544 3774 5574 3808
rect 5752 3774 5782 3808
rect 5544 3706 5574 3740
rect 5752 3706 5782 3740
rect 5544 3638 5574 3672
rect 5752 3638 5782 3672
rect 5544 3570 5574 3604
rect 5752 3570 5782 3604
rect 5544 3502 5574 3536
rect 5752 3502 5782 3536
rect 5544 3434 5574 3468
rect 5752 3434 5782 3468
rect 5544 3366 5574 3400
rect 5752 3366 5782 3400
rect 5544 3298 5574 3332
rect 5752 3298 5782 3332
rect 5544 3230 5574 3264
rect 5752 3230 5782 3264
rect 5544 3162 5574 3196
rect 5752 3162 5782 3196
rect 5544 3080 5574 3128
rect 5608 3080 5718 3092
rect 5752 3080 5782 3128
rect 5544 3040 5782 3080
rect 5544 2574 5574 3040
rect 5752 2574 5782 3040
rect 5544 2535 5782 2574
rect 5544 2501 5574 2535
rect 5608 2501 5646 2535
rect 5680 2501 5718 2535
rect 5752 2501 5782 2535
rect 5544 2461 5782 2501
rect 5544 2449 5646 2461
rect 5680 2449 5782 2461
rect 5544 2445 5574 2449
rect 5752 2445 5782 2449
rect 5544 2377 5574 2411
rect 5752 2377 5782 2411
rect 5544 2309 5574 2343
rect 5752 2309 5782 2343
rect 5544 2241 5574 2275
rect 5752 2241 5782 2275
rect 5544 2173 5574 2207
rect 5752 2173 5782 2207
rect 5544 2105 5574 2139
rect 5752 2105 5782 2139
rect 5544 2037 5574 2071
rect 5752 2037 5782 2071
rect 5544 1969 5574 2003
rect 5752 1969 5782 2003
rect 5544 1901 5574 1935
rect 5752 1901 5782 1935
rect 5544 1833 5574 1867
rect 5752 1833 5782 1867
rect 5544 1765 5574 1799
rect 5752 1765 5782 1799
rect 5544 1697 5574 1731
rect 5752 1697 5782 1731
rect 5544 1629 5574 1663
rect 5752 1629 5782 1663
rect 5544 1561 5574 1595
rect 5752 1561 5782 1595
rect 5544 1479 5574 1527
rect 5608 1479 5718 1491
rect 5752 1479 5782 1527
rect 5544 1464 5782 1479
rect 5884 3010 6004 4106
rect 6314 4388 6321 4494
rect 6427 4388 6434 4494
rect 6974 4388 6996 4494
rect 6314 4214 6434 4388
rect 6314 4180 6357 4214
rect 6391 4180 6434 4214
rect 6314 4140 6434 4180
rect 6314 4106 6357 4140
rect 6391 4106 6434 4140
rect 5884 2976 5927 3010
rect 5961 2976 6004 3010
rect 5884 2932 6004 2976
rect 5884 2898 5927 2932
rect 5961 2898 6004 2932
rect 5884 2854 6004 2898
rect 5884 2820 5927 2854
rect 5961 2820 6004 2854
rect 5884 2776 6004 2820
rect 5884 2742 5927 2776
rect 5961 2742 6004 2776
rect 5884 2697 6004 2742
rect 5884 2663 5927 2697
rect 5961 2663 6004 2697
rect 5884 2618 6004 2663
rect 5884 2584 5927 2618
rect 5961 2584 6004 2618
rect 5884 2539 6004 2584
rect 5884 2505 5927 2539
rect 5961 2505 6004 2539
rect 5322 1375 5365 1409
rect 5399 1375 5442 1409
rect 5322 1335 5442 1375
rect 5322 1301 5365 1335
rect 5399 1301 5442 1335
rect 5322 1285 5442 1301
rect 5884 1409 6004 2505
rect 6069 4028 6070 4062
rect 6104 4046 6142 4062
rect 6104 4028 6106 4046
rect 6069 4012 6106 4028
rect 6140 4028 6142 4046
rect 6176 4046 6214 4062
rect 6176 4028 6178 4046
rect 6140 4012 6178 4028
rect 6212 4028 6214 4046
rect 6248 4028 6249 4062
rect 6212 4012 6249 4028
rect 6069 3988 6249 4012
rect 6069 3954 6070 3988
rect 6104 3978 6142 3988
rect 6104 3954 6106 3978
rect 6069 3944 6106 3954
rect 6140 3954 6142 3978
rect 6176 3978 6214 3988
rect 6176 3954 6178 3978
rect 6140 3944 6178 3954
rect 6212 3954 6214 3978
rect 6248 3954 6249 3988
rect 6212 3944 6249 3954
rect 6069 3914 6249 3944
rect 6069 3880 6070 3914
rect 6104 3910 6142 3914
rect 6104 3880 6106 3910
rect 6069 3876 6106 3880
rect 6140 3880 6142 3910
rect 6176 3910 6214 3914
rect 6176 3880 6178 3910
rect 6140 3876 6178 3880
rect 6212 3880 6214 3910
rect 6248 3880 6249 3914
rect 6212 3876 6249 3880
rect 6069 3842 6249 3876
rect 6069 3840 6106 3842
rect 6069 3806 6070 3840
rect 6104 3808 6106 3840
rect 6140 3840 6178 3842
rect 6140 3808 6142 3840
rect 6104 3806 6142 3808
rect 6176 3808 6178 3840
rect 6212 3840 6249 3842
rect 6212 3808 6214 3840
rect 6176 3806 6214 3808
rect 6248 3806 6249 3840
rect 6069 3774 6249 3806
rect 6069 3766 6106 3774
rect 6069 3732 6070 3766
rect 6104 3740 6106 3766
rect 6140 3766 6178 3774
rect 6140 3740 6142 3766
rect 6104 3732 6142 3740
rect 6176 3740 6178 3766
rect 6212 3766 6249 3774
rect 6212 3740 6214 3766
rect 6176 3732 6214 3740
rect 6248 3732 6249 3766
rect 6069 3706 6249 3732
rect 6069 3692 6106 3706
rect 6069 3658 6070 3692
rect 6104 3672 6106 3692
rect 6140 3692 6178 3706
rect 6140 3672 6142 3692
rect 6104 3658 6142 3672
rect 6176 3672 6178 3692
rect 6212 3692 6249 3706
rect 6212 3672 6214 3692
rect 6176 3658 6214 3672
rect 6248 3658 6249 3692
rect 6069 3638 6249 3658
rect 6069 3618 6106 3638
rect 6069 3584 6070 3618
rect 6104 3604 6106 3618
rect 6140 3618 6178 3638
rect 6140 3604 6142 3618
rect 6104 3584 6142 3604
rect 6176 3604 6178 3618
rect 6212 3618 6249 3638
rect 6212 3604 6214 3618
rect 6176 3584 6214 3604
rect 6248 3584 6249 3618
rect 6069 3570 6249 3584
rect 6069 3544 6106 3570
rect 6069 3510 6070 3544
rect 6104 3536 6106 3544
rect 6140 3544 6178 3570
rect 6140 3536 6142 3544
rect 6104 3510 6142 3536
rect 6176 3536 6178 3544
rect 6212 3544 6249 3570
rect 6212 3536 6214 3544
rect 6176 3510 6214 3536
rect 6248 3510 6249 3544
rect 6069 3502 6249 3510
rect 6069 3470 6106 3502
rect 6069 3436 6070 3470
rect 6104 3468 6106 3470
rect 6140 3470 6178 3502
rect 6140 3468 6142 3470
rect 6104 3436 6142 3468
rect 6176 3468 6178 3470
rect 6212 3470 6249 3502
rect 6212 3468 6214 3470
rect 6176 3436 6214 3468
rect 6248 3436 6249 3470
rect 6069 3434 6249 3436
rect 6069 3400 6106 3434
rect 6140 3400 6178 3434
rect 6212 3400 6249 3434
rect 6069 3396 6249 3400
rect 6069 3362 6070 3396
rect 6104 3366 6142 3396
rect 6104 3362 6106 3366
rect 6069 3332 6106 3362
rect 6140 3362 6142 3366
rect 6176 3366 6214 3396
rect 6176 3362 6178 3366
rect 6140 3332 6178 3362
rect 6212 3362 6214 3366
rect 6248 3362 6249 3396
rect 6212 3332 6249 3362
rect 6069 3322 6249 3332
rect 6069 3288 6070 3322
rect 6104 3298 6142 3322
rect 6104 3288 6106 3298
rect 6069 3264 6106 3288
rect 6140 3288 6142 3298
rect 6176 3298 6214 3322
rect 6176 3288 6178 3298
rect 6140 3264 6178 3288
rect 6212 3288 6214 3298
rect 6248 3288 6249 3322
rect 6212 3264 6249 3288
rect 6069 3248 6249 3264
rect 6069 3214 6070 3248
rect 6104 3230 6142 3248
rect 6104 3214 6106 3230
rect 6069 3196 6106 3214
rect 6140 3214 6142 3230
rect 6176 3230 6214 3248
rect 6176 3214 6178 3230
rect 6140 3196 6178 3214
rect 6212 3214 6214 3230
rect 6248 3214 6249 3248
rect 6212 3196 6249 3214
rect 6069 3174 6249 3196
rect 6069 3140 6070 3174
rect 6104 3162 6142 3174
rect 6104 3140 6106 3162
rect 6069 3128 6106 3140
rect 6140 3140 6142 3162
rect 6176 3162 6214 3174
rect 6176 3140 6178 3162
rect 6140 3128 6178 3140
rect 6212 3140 6214 3162
rect 6248 3140 6249 3174
rect 6212 3128 6249 3140
rect 6069 3100 6249 3128
rect 6069 3066 6070 3100
rect 6104 3066 6142 3100
rect 6176 3066 6214 3100
rect 6248 3066 6249 3100
rect 6069 3026 6249 3066
rect 6069 2992 6070 3026
rect 6104 2992 6142 3026
rect 6176 2992 6214 3026
rect 6248 2992 6249 3026
rect 6069 2952 6249 2992
rect 6069 2918 6070 2952
rect 6104 2918 6142 2952
rect 6176 2918 6214 2952
rect 6248 2918 6249 2952
rect 6069 2878 6249 2918
rect 6069 2844 6070 2878
rect 6104 2844 6142 2878
rect 6176 2844 6214 2878
rect 6248 2844 6249 2878
rect 6069 2804 6249 2844
rect 6069 2770 6070 2804
rect 6104 2770 6142 2804
rect 6176 2770 6214 2804
rect 6248 2770 6249 2804
rect 6069 2730 6249 2770
rect 6069 2696 6070 2730
rect 6104 2696 6142 2730
rect 6176 2696 6214 2730
rect 6248 2696 6249 2730
rect 6069 2656 6249 2696
rect 6069 2622 6070 2656
rect 6104 2622 6142 2656
rect 6176 2622 6214 2656
rect 6248 2622 6249 2656
rect 6069 2582 6249 2622
rect 6069 2548 6070 2582
rect 6104 2548 6142 2582
rect 6176 2548 6214 2582
rect 6248 2548 6249 2582
rect 6069 2508 6249 2548
rect 6069 2474 6070 2508
rect 6104 2474 6142 2508
rect 6176 2474 6214 2508
rect 6248 2474 6249 2508
rect 6069 2445 6249 2474
rect 6069 2434 6106 2445
rect 6069 2400 6070 2434
rect 6104 2411 6106 2434
rect 6140 2434 6178 2445
rect 6140 2411 6142 2434
rect 6104 2400 6142 2411
rect 6176 2411 6178 2434
rect 6212 2434 6249 2445
rect 6212 2411 6214 2434
rect 6176 2400 6214 2411
rect 6248 2400 6249 2434
rect 6069 2377 6249 2400
rect 6069 2360 6106 2377
rect 6069 2326 6070 2360
rect 6104 2343 6106 2360
rect 6140 2360 6178 2377
rect 6140 2343 6142 2360
rect 6104 2326 6142 2343
rect 6176 2343 6178 2360
rect 6212 2360 6249 2377
rect 6212 2343 6214 2360
rect 6176 2326 6214 2343
rect 6248 2326 6249 2360
rect 6069 2309 6249 2326
rect 6069 2286 6106 2309
rect 6069 2252 6070 2286
rect 6104 2275 6106 2286
rect 6140 2286 6178 2309
rect 6140 2275 6142 2286
rect 6104 2252 6142 2275
rect 6176 2275 6178 2286
rect 6212 2286 6249 2309
rect 6212 2275 6214 2286
rect 6176 2252 6214 2275
rect 6248 2252 6249 2286
rect 6069 2241 6249 2252
rect 6069 2212 6106 2241
rect 6069 2178 6070 2212
rect 6104 2207 6106 2212
rect 6140 2212 6178 2241
rect 6140 2207 6142 2212
rect 6104 2178 6142 2207
rect 6176 2207 6178 2212
rect 6212 2212 6249 2241
rect 6212 2207 6214 2212
rect 6176 2178 6214 2207
rect 6248 2178 6249 2212
rect 6069 2173 6249 2178
rect 6069 2139 6106 2173
rect 6140 2139 6178 2173
rect 6212 2139 6249 2173
rect 6069 2138 6249 2139
rect 6069 2104 6070 2138
rect 6104 2105 6142 2138
rect 6104 2104 6106 2105
rect 6069 2071 6106 2104
rect 6140 2104 6142 2105
rect 6176 2105 6214 2138
rect 6176 2104 6178 2105
rect 6140 2071 6178 2104
rect 6212 2104 6214 2105
rect 6248 2104 6249 2138
rect 6212 2071 6249 2104
rect 6069 2064 6249 2071
rect 6069 2030 6070 2064
rect 6104 2037 6142 2064
rect 6104 2030 6106 2037
rect 6069 2003 6106 2030
rect 6140 2030 6142 2037
rect 6176 2037 6214 2064
rect 6176 2030 6178 2037
rect 6140 2003 6178 2030
rect 6212 2030 6214 2037
rect 6248 2030 6249 2064
rect 6212 2003 6249 2030
rect 6069 1990 6249 2003
rect 6069 1956 6070 1990
rect 6104 1969 6142 1990
rect 6104 1956 6106 1969
rect 6069 1935 6106 1956
rect 6140 1956 6142 1969
rect 6176 1969 6214 1990
rect 6176 1956 6178 1969
rect 6140 1935 6178 1956
rect 6212 1956 6214 1969
rect 6248 1956 6249 1990
rect 6212 1935 6249 1956
rect 6069 1916 6249 1935
rect 6069 1882 6070 1916
rect 6104 1901 6142 1916
rect 6104 1882 6106 1901
rect 6069 1867 6106 1882
rect 6140 1882 6142 1901
rect 6176 1901 6214 1916
rect 6176 1882 6178 1901
rect 6140 1867 6178 1882
rect 6212 1882 6214 1901
rect 6248 1882 6249 1916
rect 6212 1867 6249 1882
rect 6069 1842 6249 1867
rect 6069 1808 6070 1842
rect 6104 1833 6142 1842
rect 6104 1808 6106 1833
rect 6069 1799 6106 1808
rect 6140 1808 6142 1833
rect 6176 1833 6214 1842
rect 6176 1808 6178 1833
rect 6140 1799 6178 1808
rect 6212 1808 6214 1833
rect 6248 1808 6249 1842
rect 6212 1799 6249 1808
rect 6069 1768 6249 1799
rect 6069 1734 6070 1768
rect 6104 1765 6142 1768
rect 6104 1734 6106 1765
rect 6069 1731 6106 1734
rect 6140 1734 6142 1765
rect 6176 1765 6214 1768
rect 6176 1734 6178 1765
rect 6140 1731 6178 1734
rect 6212 1734 6214 1765
rect 6248 1734 6249 1768
rect 6212 1731 6249 1734
rect 6069 1697 6249 1731
rect 6069 1694 6106 1697
rect 6069 1660 6070 1694
rect 6104 1663 6106 1694
rect 6140 1694 6178 1697
rect 6140 1663 6142 1694
rect 6104 1660 6142 1663
rect 6176 1663 6178 1694
rect 6212 1694 6249 1697
rect 6212 1663 6214 1694
rect 6176 1660 6214 1663
rect 6248 1660 6249 1694
rect 6069 1629 6249 1660
rect 6069 1620 6106 1629
rect 6069 1586 6070 1620
rect 6104 1595 6106 1620
rect 6140 1620 6178 1629
rect 6140 1595 6142 1620
rect 6104 1586 6142 1595
rect 6176 1595 6178 1620
rect 6212 1620 6249 1629
rect 6212 1595 6214 1620
rect 6176 1586 6214 1595
rect 6248 1586 6249 1620
rect 6069 1561 6249 1586
rect 6069 1545 6106 1561
rect 6069 1511 6070 1545
rect 6104 1527 6106 1545
rect 6140 1545 6178 1561
rect 6140 1527 6142 1545
rect 6104 1511 6142 1527
rect 6176 1527 6178 1545
rect 6212 1545 6249 1561
rect 6212 1527 6214 1545
rect 6176 1511 6214 1527
rect 6248 1511 6249 1545
rect 6314 3010 6434 4106
rect 6876 4214 6996 4388
rect 6876 4180 6919 4214
rect 6953 4180 6996 4214
rect 6876 4140 6996 4180
rect 6876 4106 6919 4140
rect 6953 4106 6996 4140
rect 6314 2976 6357 3010
rect 6391 2976 6434 3010
rect 6314 2932 6434 2976
rect 6314 2898 6357 2932
rect 6391 2898 6434 2932
rect 6314 2854 6434 2898
rect 6314 2820 6357 2854
rect 6391 2820 6434 2854
rect 6314 2776 6434 2820
rect 6314 2742 6357 2776
rect 6391 2742 6434 2776
rect 6314 2697 6434 2742
rect 6314 2663 6357 2697
rect 6391 2663 6434 2697
rect 6314 2618 6434 2663
rect 6314 2584 6357 2618
rect 6391 2584 6434 2618
rect 6314 2539 6434 2584
rect 6314 2505 6357 2539
rect 6391 2505 6434 2539
rect 6106 1491 6212 1511
rect 5884 1375 5927 1409
rect 5961 1375 6004 1409
rect 5884 1335 6004 1375
rect 5884 1301 5927 1335
rect 5961 1301 6004 1335
rect 5884 1285 6004 1301
rect 6314 1409 6434 2505
rect 6536 4050 6638 4062
rect 6672 4050 6774 4062
rect 6536 4046 6566 4050
rect 6744 4046 6774 4050
rect 6536 3978 6566 4012
rect 6744 3978 6774 4012
rect 6536 3910 6566 3944
rect 6744 3910 6774 3944
rect 6536 3842 6566 3876
rect 6744 3842 6774 3876
rect 6536 3774 6566 3808
rect 6744 3774 6774 3808
rect 6536 3706 6566 3740
rect 6744 3706 6774 3740
rect 6536 3638 6566 3672
rect 6744 3638 6774 3672
rect 6536 3570 6566 3604
rect 6744 3570 6774 3604
rect 6536 3502 6566 3536
rect 6744 3502 6774 3536
rect 6536 3434 6566 3468
rect 6744 3434 6774 3468
rect 6536 3366 6566 3400
rect 6744 3366 6774 3400
rect 6536 3298 6566 3332
rect 6744 3298 6774 3332
rect 6536 3230 6566 3264
rect 6744 3230 6774 3264
rect 6536 3162 6566 3196
rect 6744 3162 6774 3196
rect 6536 3080 6566 3128
rect 6600 3080 6710 3092
rect 6744 3080 6774 3128
rect 6536 3040 6774 3080
rect 6536 2574 6566 3040
rect 6744 2574 6774 3040
rect 6536 2535 6774 2574
rect 6536 2501 6566 2535
rect 6600 2501 6638 2535
rect 6672 2501 6710 2535
rect 6744 2501 6774 2535
rect 6536 2461 6774 2501
rect 6536 2449 6638 2461
rect 6672 2449 6774 2461
rect 6536 2445 6566 2449
rect 6744 2445 6774 2449
rect 6536 2377 6566 2411
rect 6744 2377 6774 2411
rect 6536 2309 6566 2343
rect 6744 2309 6774 2343
rect 6536 2241 6566 2275
rect 6744 2241 6774 2275
rect 6536 2173 6566 2207
rect 6744 2173 6774 2207
rect 6536 2105 6566 2139
rect 6744 2105 6774 2139
rect 6536 2037 6566 2071
rect 6744 2037 6774 2071
rect 6536 1969 6566 2003
rect 6744 1969 6774 2003
rect 6536 1901 6566 1935
rect 6744 1901 6774 1935
rect 6536 1833 6566 1867
rect 6744 1833 6774 1867
rect 6536 1765 6566 1799
rect 6744 1765 6774 1799
rect 6536 1697 6566 1731
rect 6744 1697 6774 1731
rect 6536 1629 6566 1663
rect 6744 1629 6774 1663
rect 6536 1561 6566 1595
rect 6744 1561 6774 1595
rect 6536 1479 6566 1527
rect 6600 1479 6710 1491
rect 6744 1479 6774 1527
rect 6536 1464 6774 1479
rect 6876 3010 6996 4106
rect 7306 4388 7313 4494
rect 7419 4388 7426 4494
rect 7306 4214 7426 4388
rect 7306 4180 7349 4214
rect 7383 4180 7426 4214
rect 7306 4140 7426 4180
rect 7306 4106 7349 4140
rect 7383 4106 7426 4140
rect 6876 2976 6919 3010
rect 6953 2976 6996 3010
rect 6876 2932 6996 2976
rect 6876 2898 6919 2932
rect 6953 2898 6996 2932
rect 6876 2854 6996 2898
rect 6876 2820 6919 2854
rect 6953 2820 6996 2854
rect 6876 2776 6996 2820
rect 6876 2742 6919 2776
rect 6953 2742 6996 2776
rect 6876 2697 6996 2742
rect 6876 2663 6919 2697
rect 6953 2663 6996 2697
rect 6876 2618 6996 2663
rect 6876 2584 6919 2618
rect 6953 2584 6996 2618
rect 6876 2539 6996 2584
rect 6876 2505 6919 2539
rect 6953 2505 6996 2539
rect 6314 1375 6357 1409
rect 6391 1375 6434 1409
rect 6314 1335 6434 1375
rect 6314 1301 6357 1335
rect 6391 1301 6434 1335
rect 6314 1285 6434 1301
rect 6876 1409 6996 2505
rect 7061 4028 7062 4062
rect 7096 4046 7134 4062
rect 7096 4028 7098 4046
rect 7061 4012 7098 4028
rect 7132 4028 7134 4046
rect 7168 4046 7206 4062
rect 7168 4028 7170 4046
rect 7132 4012 7170 4028
rect 7204 4028 7206 4046
rect 7240 4028 7241 4062
rect 7204 4012 7241 4028
rect 7061 3988 7241 4012
rect 7061 3954 7062 3988
rect 7096 3978 7134 3988
rect 7096 3954 7098 3978
rect 7061 3944 7098 3954
rect 7132 3954 7134 3978
rect 7168 3978 7206 3988
rect 7168 3954 7170 3978
rect 7132 3944 7170 3954
rect 7204 3954 7206 3978
rect 7240 3954 7241 3988
rect 7204 3944 7241 3954
rect 7061 3914 7241 3944
rect 7061 3880 7062 3914
rect 7096 3910 7134 3914
rect 7096 3880 7098 3910
rect 7061 3876 7098 3880
rect 7132 3880 7134 3910
rect 7168 3910 7206 3914
rect 7168 3880 7170 3910
rect 7132 3876 7170 3880
rect 7204 3880 7206 3910
rect 7240 3880 7241 3914
rect 7204 3876 7241 3880
rect 7061 3842 7241 3876
rect 7061 3840 7098 3842
rect 7061 3806 7062 3840
rect 7096 3808 7098 3840
rect 7132 3840 7170 3842
rect 7132 3808 7134 3840
rect 7096 3806 7134 3808
rect 7168 3808 7170 3840
rect 7204 3840 7241 3842
rect 7204 3808 7206 3840
rect 7168 3806 7206 3808
rect 7240 3806 7241 3840
rect 7061 3774 7241 3806
rect 7061 3766 7098 3774
rect 7061 3732 7062 3766
rect 7096 3740 7098 3766
rect 7132 3766 7170 3774
rect 7132 3740 7134 3766
rect 7096 3732 7134 3740
rect 7168 3740 7170 3766
rect 7204 3766 7241 3774
rect 7204 3740 7206 3766
rect 7168 3732 7206 3740
rect 7240 3732 7241 3766
rect 7061 3706 7241 3732
rect 7061 3692 7098 3706
rect 7061 3658 7062 3692
rect 7096 3672 7098 3692
rect 7132 3692 7170 3706
rect 7132 3672 7134 3692
rect 7096 3658 7134 3672
rect 7168 3672 7170 3692
rect 7204 3692 7241 3706
rect 7204 3672 7206 3692
rect 7168 3658 7206 3672
rect 7240 3658 7241 3692
rect 7061 3638 7241 3658
rect 7061 3618 7098 3638
rect 7061 3584 7062 3618
rect 7096 3604 7098 3618
rect 7132 3618 7170 3638
rect 7132 3604 7134 3618
rect 7096 3584 7134 3604
rect 7168 3604 7170 3618
rect 7204 3618 7241 3638
rect 7204 3604 7206 3618
rect 7168 3584 7206 3604
rect 7240 3584 7241 3618
rect 7061 3570 7241 3584
rect 7061 3544 7098 3570
rect 7061 3510 7062 3544
rect 7096 3536 7098 3544
rect 7132 3544 7170 3570
rect 7132 3536 7134 3544
rect 7096 3510 7134 3536
rect 7168 3536 7170 3544
rect 7204 3544 7241 3570
rect 7204 3536 7206 3544
rect 7168 3510 7206 3536
rect 7240 3510 7241 3544
rect 7061 3502 7241 3510
rect 7061 3470 7098 3502
rect 7061 3436 7062 3470
rect 7096 3468 7098 3470
rect 7132 3470 7170 3502
rect 7132 3468 7134 3470
rect 7096 3436 7134 3468
rect 7168 3468 7170 3470
rect 7204 3470 7241 3502
rect 7204 3468 7206 3470
rect 7168 3436 7206 3468
rect 7240 3436 7241 3470
rect 7061 3434 7241 3436
rect 7061 3400 7098 3434
rect 7132 3400 7170 3434
rect 7204 3400 7241 3434
rect 7061 3396 7241 3400
rect 7061 3362 7062 3396
rect 7096 3366 7134 3396
rect 7096 3362 7098 3366
rect 7061 3332 7098 3362
rect 7132 3362 7134 3366
rect 7168 3366 7206 3396
rect 7168 3362 7170 3366
rect 7132 3332 7170 3362
rect 7204 3362 7206 3366
rect 7240 3362 7241 3396
rect 7204 3332 7241 3362
rect 7061 3322 7241 3332
rect 7061 3288 7062 3322
rect 7096 3298 7134 3322
rect 7096 3288 7098 3298
rect 7061 3264 7098 3288
rect 7132 3288 7134 3298
rect 7168 3298 7206 3322
rect 7168 3288 7170 3298
rect 7132 3264 7170 3288
rect 7204 3288 7206 3298
rect 7240 3288 7241 3322
rect 7204 3264 7241 3288
rect 7061 3248 7241 3264
rect 7061 3214 7062 3248
rect 7096 3230 7134 3248
rect 7096 3214 7098 3230
rect 7061 3196 7098 3214
rect 7132 3214 7134 3230
rect 7168 3230 7206 3248
rect 7168 3214 7170 3230
rect 7132 3196 7170 3214
rect 7204 3214 7206 3230
rect 7240 3214 7241 3248
rect 7204 3196 7241 3214
rect 7061 3174 7241 3196
rect 7061 3140 7062 3174
rect 7096 3162 7134 3174
rect 7096 3140 7098 3162
rect 7061 3128 7098 3140
rect 7132 3140 7134 3162
rect 7168 3162 7206 3174
rect 7168 3140 7170 3162
rect 7132 3128 7170 3140
rect 7204 3140 7206 3162
rect 7240 3140 7241 3174
rect 7204 3128 7241 3140
rect 7061 3100 7241 3128
rect 7061 3066 7062 3100
rect 7096 3066 7134 3100
rect 7168 3066 7206 3100
rect 7240 3066 7241 3100
rect 7061 3026 7241 3066
rect 7061 2992 7062 3026
rect 7096 2992 7134 3026
rect 7168 2992 7206 3026
rect 7240 2992 7241 3026
rect 7061 2952 7241 2992
rect 7061 2918 7062 2952
rect 7096 2918 7134 2952
rect 7168 2918 7206 2952
rect 7240 2918 7241 2952
rect 7061 2878 7241 2918
rect 7061 2844 7062 2878
rect 7096 2844 7134 2878
rect 7168 2844 7206 2878
rect 7240 2844 7241 2878
rect 7061 2804 7241 2844
rect 7061 2770 7062 2804
rect 7096 2770 7134 2804
rect 7168 2770 7206 2804
rect 7240 2770 7241 2804
rect 7061 2730 7241 2770
rect 7061 2696 7062 2730
rect 7096 2696 7134 2730
rect 7168 2696 7206 2730
rect 7240 2696 7241 2730
rect 7061 2656 7241 2696
rect 7061 2622 7062 2656
rect 7096 2622 7134 2656
rect 7168 2622 7206 2656
rect 7240 2622 7241 2656
rect 7061 2582 7241 2622
rect 7061 2548 7062 2582
rect 7096 2548 7134 2582
rect 7168 2548 7206 2582
rect 7240 2548 7241 2582
rect 7061 2508 7241 2548
rect 7061 2474 7062 2508
rect 7096 2474 7134 2508
rect 7168 2474 7206 2508
rect 7240 2474 7241 2508
rect 7061 2445 7241 2474
rect 7061 2434 7098 2445
rect 7061 2400 7062 2434
rect 7096 2411 7098 2434
rect 7132 2434 7170 2445
rect 7132 2411 7134 2434
rect 7096 2400 7134 2411
rect 7168 2411 7170 2434
rect 7204 2434 7241 2445
rect 7204 2411 7206 2434
rect 7168 2400 7206 2411
rect 7240 2400 7241 2434
rect 7061 2377 7241 2400
rect 7061 2360 7098 2377
rect 7061 2326 7062 2360
rect 7096 2343 7098 2360
rect 7132 2360 7170 2377
rect 7132 2343 7134 2360
rect 7096 2326 7134 2343
rect 7168 2343 7170 2360
rect 7204 2360 7241 2377
rect 7204 2343 7206 2360
rect 7168 2326 7206 2343
rect 7240 2326 7241 2360
rect 7061 2309 7241 2326
rect 7061 2286 7098 2309
rect 7061 2252 7062 2286
rect 7096 2275 7098 2286
rect 7132 2286 7170 2309
rect 7132 2275 7134 2286
rect 7096 2252 7134 2275
rect 7168 2275 7170 2286
rect 7204 2286 7241 2309
rect 7204 2275 7206 2286
rect 7168 2252 7206 2275
rect 7240 2252 7241 2286
rect 7061 2241 7241 2252
rect 7061 2212 7098 2241
rect 7061 2178 7062 2212
rect 7096 2207 7098 2212
rect 7132 2212 7170 2241
rect 7132 2207 7134 2212
rect 7096 2178 7134 2207
rect 7168 2207 7170 2212
rect 7204 2212 7241 2241
rect 7204 2207 7206 2212
rect 7168 2178 7206 2207
rect 7240 2178 7241 2212
rect 7061 2173 7241 2178
rect 7061 2139 7098 2173
rect 7132 2139 7170 2173
rect 7204 2139 7241 2173
rect 7061 2138 7241 2139
rect 7061 2104 7062 2138
rect 7096 2105 7134 2138
rect 7096 2104 7098 2105
rect 7061 2071 7098 2104
rect 7132 2104 7134 2105
rect 7168 2105 7206 2138
rect 7168 2104 7170 2105
rect 7132 2071 7170 2104
rect 7204 2104 7206 2105
rect 7240 2104 7241 2138
rect 7204 2071 7241 2104
rect 7061 2064 7241 2071
rect 7061 2030 7062 2064
rect 7096 2037 7134 2064
rect 7096 2030 7098 2037
rect 7061 2003 7098 2030
rect 7132 2030 7134 2037
rect 7168 2037 7206 2064
rect 7168 2030 7170 2037
rect 7132 2003 7170 2030
rect 7204 2030 7206 2037
rect 7240 2030 7241 2064
rect 7204 2003 7241 2030
rect 7061 1990 7241 2003
rect 7061 1956 7062 1990
rect 7096 1969 7134 1990
rect 7096 1956 7098 1969
rect 7061 1935 7098 1956
rect 7132 1956 7134 1969
rect 7168 1969 7206 1990
rect 7168 1956 7170 1969
rect 7132 1935 7170 1956
rect 7204 1956 7206 1969
rect 7240 1956 7241 1990
rect 7204 1935 7241 1956
rect 7061 1916 7241 1935
rect 7061 1882 7062 1916
rect 7096 1901 7134 1916
rect 7096 1882 7098 1901
rect 7061 1867 7098 1882
rect 7132 1882 7134 1901
rect 7168 1901 7206 1916
rect 7168 1882 7170 1901
rect 7132 1867 7170 1882
rect 7204 1882 7206 1901
rect 7240 1882 7241 1916
rect 7204 1867 7241 1882
rect 7061 1842 7241 1867
rect 7061 1808 7062 1842
rect 7096 1833 7134 1842
rect 7096 1808 7098 1833
rect 7061 1799 7098 1808
rect 7132 1808 7134 1833
rect 7168 1833 7206 1842
rect 7168 1808 7170 1833
rect 7132 1799 7170 1808
rect 7204 1808 7206 1833
rect 7240 1808 7241 1842
rect 7204 1799 7241 1808
rect 7061 1768 7241 1799
rect 7061 1734 7062 1768
rect 7096 1765 7134 1768
rect 7096 1734 7098 1765
rect 7061 1731 7098 1734
rect 7132 1734 7134 1765
rect 7168 1765 7206 1768
rect 7168 1734 7170 1765
rect 7132 1731 7170 1734
rect 7204 1734 7206 1765
rect 7240 1734 7241 1768
rect 7204 1731 7241 1734
rect 7061 1697 7241 1731
rect 7061 1694 7098 1697
rect 7061 1660 7062 1694
rect 7096 1663 7098 1694
rect 7132 1694 7170 1697
rect 7132 1663 7134 1694
rect 7096 1660 7134 1663
rect 7168 1663 7170 1694
rect 7204 1694 7241 1697
rect 7204 1663 7206 1694
rect 7168 1660 7206 1663
rect 7240 1660 7241 1694
rect 7061 1629 7241 1660
rect 7061 1620 7098 1629
rect 7061 1586 7062 1620
rect 7096 1595 7098 1620
rect 7132 1620 7170 1629
rect 7132 1595 7134 1620
rect 7096 1586 7134 1595
rect 7168 1595 7170 1620
rect 7204 1620 7241 1629
rect 7204 1595 7206 1620
rect 7168 1586 7206 1595
rect 7240 1586 7241 1620
rect 7061 1561 7241 1586
rect 7061 1545 7098 1561
rect 7061 1511 7062 1545
rect 7096 1527 7098 1545
rect 7132 1545 7170 1561
rect 7132 1527 7134 1545
rect 7096 1511 7134 1527
rect 7168 1527 7170 1545
rect 7204 1545 7241 1561
rect 7204 1527 7206 1545
rect 7168 1511 7206 1527
rect 7240 1511 7241 1545
rect 7306 3010 7426 4106
rect 7868 4388 7875 4494
rect 7981 4388 7988 4494
rect 7868 4214 7988 4388
rect 7868 4180 7911 4214
rect 7945 4180 7988 4214
rect 7868 4140 7988 4180
rect 7868 4106 7911 4140
rect 7945 4106 7988 4140
rect 7306 2976 7349 3010
rect 7383 2976 7426 3010
rect 7306 2932 7426 2976
rect 7306 2898 7349 2932
rect 7383 2898 7426 2932
rect 7306 2854 7426 2898
rect 7306 2820 7349 2854
rect 7383 2820 7426 2854
rect 7306 2776 7426 2820
rect 7306 2742 7349 2776
rect 7383 2742 7426 2776
rect 7306 2697 7426 2742
rect 7306 2663 7349 2697
rect 7383 2663 7426 2697
rect 7306 2618 7426 2663
rect 7306 2584 7349 2618
rect 7383 2584 7426 2618
rect 7306 2539 7426 2584
rect 7306 2505 7349 2539
rect 7383 2505 7426 2539
rect 7098 1491 7204 1511
rect 6876 1375 6919 1409
rect 6953 1375 6996 1409
rect 6876 1335 6996 1375
rect 6876 1301 6919 1335
rect 6953 1301 6996 1335
rect 6876 1285 6996 1301
rect 7306 1409 7426 2505
rect 7528 4050 7630 4062
rect 7664 4050 7766 4062
rect 7528 4046 7558 4050
rect 7736 4046 7766 4050
rect 7528 3978 7558 4012
rect 7736 3978 7766 4012
rect 7528 3910 7558 3944
rect 7736 3910 7766 3944
rect 7528 3842 7558 3876
rect 7736 3842 7766 3876
rect 7528 3774 7558 3808
rect 7736 3774 7766 3808
rect 7528 3706 7558 3740
rect 7736 3706 7766 3740
rect 7528 3638 7558 3672
rect 7736 3638 7766 3672
rect 7528 3570 7558 3604
rect 7736 3570 7766 3604
rect 7528 3502 7558 3536
rect 7736 3502 7766 3536
rect 7528 3434 7558 3468
rect 7736 3434 7766 3468
rect 7528 3366 7558 3400
rect 7736 3366 7766 3400
rect 7528 3298 7558 3332
rect 7736 3298 7766 3332
rect 7528 3230 7558 3264
rect 7736 3230 7766 3264
rect 7528 3162 7558 3196
rect 7736 3162 7766 3196
rect 7528 3080 7558 3128
rect 7592 3080 7702 3092
rect 7736 3080 7766 3128
rect 7528 3040 7766 3080
rect 7528 2574 7558 3040
rect 7736 2574 7766 3040
rect 7528 2535 7766 2574
rect 7528 2501 7558 2535
rect 7592 2501 7630 2535
rect 7664 2501 7702 2535
rect 7736 2501 7766 2535
rect 7528 2461 7766 2501
rect 7528 2449 7630 2461
rect 7664 2449 7766 2461
rect 7528 2445 7558 2449
rect 7736 2445 7766 2449
rect 7528 2377 7558 2411
rect 7736 2377 7766 2411
rect 7528 2309 7558 2343
rect 7736 2309 7766 2343
rect 7528 2241 7558 2275
rect 7736 2241 7766 2275
rect 7528 2173 7558 2207
rect 7736 2173 7766 2207
rect 7528 2105 7558 2139
rect 7736 2105 7766 2139
rect 7528 2037 7558 2071
rect 7736 2037 7766 2071
rect 7528 1969 7558 2003
rect 7736 1969 7766 2003
rect 7528 1901 7558 1935
rect 7736 1901 7766 1935
rect 7528 1833 7558 1867
rect 7736 1833 7766 1867
rect 7528 1765 7558 1799
rect 7736 1765 7766 1799
rect 7528 1697 7558 1731
rect 7736 1697 7766 1731
rect 7528 1629 7558 1663
rect 7736 1629 7766 1663
rect 7528 1561 7558 1595
rect 7736 1561 7766 1595
rect 7528 1479 7558 1527
rect 7592 1479 7702 1491
rect 7736 1479 7766 1527
rect 7528 1464 7766 1479
rect 7868 3010 7988 4106
rect 8298 4388 8305 4494
rect 8411 4388 8418 4494
rect 8298 4214 8418 4388
rect 8298 4180 8341 4214
rect 8375 4180 8418 4214
rect 8298 4140 8418 4180
rect 8298 4106 8341 4140
rect 8375 4106 8418 4140
rect 7868 2976 7911 3010
rect 7945 2976 7988 3010
rect 7868 2932 7988 2976
rect 7868 2898 7911 2932
rect 7945 2898 7988 2932
rect 7868 2854 7988 2898
rect 7868 2820 7911 2854
rect 7945 2820 7988 2854
rect 7868 2776 7988 2820
rect 7868 2742 7911 2776
rect 7945 2742 7988 2776
rect 7868 2697 7988 2742
rect 7868 2663 7911 2697
rect 7945 2663 7988 2697
rect 7868 2618 7988 2663
rect 7868 2584 7911 2618
rect 7945 2584 7988 2618
rect 7868 2539 7988 2584
rect 7868 2505 7911 2539
rect 7945 2505 7988 2539
rect 7306 1375 7349 1409
rect 7383 1375 7426 1409
rect 7306 1335 7426 1375
rect 7306 1301 7349 1335
rect 7383 1301 7426 1335
rect 7306 1285 7426 1301
rect 7868 1409 7988 2505
rect 8053 4028 8054 4062
rect 8088 4046 8126 4062
rect 8088 4028 8090 4046
rect 8053 4012 8090 4028
rect 8124 4028 8126 4046
rect 8160 4046 8198 4062
rect 8160 4028 8162 4046
rect 8124 4012 8162 4028
rect 8196 4028 8198 4046
rect 8232 4028 8233 4062
rect 8196 4012 8233 4028
rect 8053 3988 8233 4012
rect 8053 3954 8054 3988
rect 8088 3978 8126 3988
rect 8088 3954 8090 3978
rect 8053 3944 8090 3954
rect 8124 3954 8126 3978
rect 8160 3978 8198 3988
rect 8160 3954 8162 3978
rect 8124 3944 8162 3954
rect 8196 3954 8198 3978
rect 8232 3954 8233 3988
rect 8196 3944 8233 3954
rect 8053 3914 8233 3944
rect 8053 3880 8054 3914
rect 8088 3910 8126 3914
rect 8088 3880 8090 3910
rect 8053 3876 8090 3880
rect 8124 3880 8126 3910
rect 8160 3910 8198 3914
rect 8160 3880 8162 3910
rect 8124 3876 8162 3880
rect 8196 3880 8198 3910
rect 8232 3880 8233 3914
rect 8196 3876 8233 3880
rect 8053 3842 8233 3876
rect 8053 3840 8090 3842
rect 8053 3806 8054 3840
rect 8088 3808 8090 3840
rect 8124 3840 8162 3842
rect 8124 3808 8126 3840
rect 8088 3806 8126 3808
rect 8160 3808 8162 3840
rect 8196 3840 8233 3842
rect 8196 3808 8198 3840
rect 8160 3806 8198 3808
rect 8232 3806 8233 3840
rect 8053 3774 8233 3806
rect 8053 3766 8090 3774
rect 8053 3732 8054 3766
rect 8088 3740 8090 3766
rect 8124 3766 8162 3774
rect 8124 3740 8126 3766
rect 8088 3732 8126 3740
rect 8160 3740 8162 3766
rect 8196 3766 8233 3774
rect 8196 3740 8198 3766
rect 8160 3732 8198 3740
rect 8232 3732 8233 3766
rect 8053 3706 8233 3732
rect 8053 3692 8090 3706
rect 8053 3658 8054 3692
rect 8088 3672 8090 3692
rect 8124 3692 8162 3706
rect 8124 3672 8126 3692
rect 8088 3658 8126 3672
rect 8160 3672 8162 3692
rect 8196 3692 8233 3706
rect 8196 3672 8198 3692
rect 8160 3658 8198 3672
rect 8232 3658 8233 3692
rect 8053 3638 8233 3658
rect 8053 3618 8090 3638
rect 8053 3584 8054 3618
rect 8088 3604 8090 3618
rect 8124 3618 8162 3638
rect 8124 3604 8126 3618
rect 8088 3584 8126 3604
rect 8160 3604 8162 3618
rect 8196 3618 8233 3638
rect 8196 3604 8198 3618
rect 8160 3584 8198 3604
rect 8232 3584 8233 3618
rect 8053 3570 8233 3584
rect 8053 3544 8090 3570
rect 8053 3510 8054 3544
rect 8088 3536 8090 3544
rect 8124 3544 8162 3570
rect 8124 3536 8126 3544
rect 8088 3510 8126 3536
rect 8160 3536 8162 3544
rect 8196 3544 8233 3570
rect 8196 3536 8198 3544
rect 8160 3510 8198 3536
rect 8232 3510 8233 3544
rect 8053 3502 8233 3510
rect 8053 3470 8090 3502
rect 8053 3436 8054 3470
rect 8088 3468 8090 3470
rect 8124 3470 8162 3502
rect 8124 3468 8126 3470
rect 8088 3436 8126 3468
rect 8160 3468 8162 3470
rect 8196 3470 8233 3502
rect 8196 3468 8198 3470
rect 8160 3436 8198 3468
rect 8232 3436 8233 3470
rect 8053 3434 8233 3436
rect 8053 3400 8090 3434
rect 8124 3400 8162 3434
rect 8196 3400 8233 3434
rect 8053 3396 8233 3400
rect 8053 3362 8054 3396
rect 8088 3366 8126 3396
rect 8088 3362 8090 3366
rect 8053 3332 8090 3362
rect 8124 3362 8126 3366
rect 8160 3366 8198 3396
rect 8160 3362 8162 3366
rect 8124 3332 8162 3362
rect 8196 3362 8198 3366
rect 8232 3362 8233 3396
rect 8196 3332 8233 3362
rect 8053 3322 8233 3332
rect 8053 3288 8054 3322
rect 8088 3298 8126 3322
rect 8088 3288 8090 3298
rect 8053 3264 8090 3288
rect 8124 3288 8126 3298
rect 8160 3298 8198 3322
rect 8160 3288 8162 3298
rect 8124 3264 8162 3288
rect 8196 3288 8198 3298
rect 8232 3288 8233 3322
rect 8196 3264 8233 3288
rect 8053 3248 8233 3264
rect 8053 3214 8054 3248
rect 8088 3230 8126 3248
rect 8088 3214 8090 3230
rect 8053 3196 8090 3214
rect 8124 3214 8126 3230
rect 8160 3230 8198 3248
rect 8160 3214 8162 3230
rect 8124 3196 8162 3214
rect 8196 3214 8198 3230
rect 8232 3214 8233 3248
rect 8196 3196 8233 3214
rect 8053 3174 8233 3196
rect 8053 3140 8054 3174
rect 8088 3162 8126 3174
rect 8088 3140 8090 3162
rect 8053 3128 8090 3140
rect 8124 3140 8126 3162
rect 8160 3162 8198 3174
rect 8160 3140 8162 3162
rect 8124 3128 8162 3140
rect 8196 3140 8198 3162
rect 8232 3140 8233 3174
rect 8196 3128 8233 3140
rect 8053 3100 8233 3128
rect 8053 3066 8054 3100
rect 8088 3066 8126 3100
rect 8160 3066 8198 3100
rect 8232 3066 8233 3100
rect 8053 3026 8233 3066
rect 8053 2992 8054 3026
rect 8088 2992 8126 3026
rect 8160 2992 8198 3026
rect 8232 2992 8233 3026
rect 8053 2952 8233 2992
rect 8053 2918 8054 2952
rect 8088 2918 8126 2952
rect 8160 2918 8198 2952
rect 8232 2918 8233 2952
rect 8053 2878 8233 2918
rect 8053 2844 8054 2878
rect 8088 2844 8126 2878
rect 8160 2844 8198 2878
rect 8232 2844 8233 2878
rect 8053 2804 8233 2844
rect 8053 2770 8054 2804
rect 8088 2770 8126 2804
rect 8160 2770 8198 2804
rect 8232 2770 8233 2804
rect 8053 2730 8233 2770
rect 8053 2696 8054 2730
rect 8088 2696 8126 2730
rect 8160 2696 8198 2730
rect 8232 2696 8233 2730
rect 8053 2656 8233 2696
rect 8053 2622 8054 2656
rect 8088 2622 8126 2656
rect 8160 2622 8198 2656
rect 8232 2622 8233 2656
rect 8053 2582 8233 2622
rect 8053 2548 8054 2582
rect 8088 2548 8126 2582
rect 8160 2548 8198 2582
rect 8232 2548 8233 2582
rect 8053 2508 8233 2548
rect 8053 2474 8054 2508
rect 8088 2474 8126 2508
rect 8160 2474 8198 2508
rect 8232 2474 8233 2508
rect 8053 2445 8233 2474
rect 8053 2434 8090 2445
rect 8053 2400 8054 2434
rect 8088 2411 8090 2434
rect 8124 2434 8162 2445
rect 8124 2411 8126 2434
rect 8088 2400 8126 2411
rect 8160 2411 8162 2434
rect 8196 2434 8233 2445
rect 8196 2411 8198 2434
rect 8160 2400 8198 2411
rect 8232 2400 8233 2434
rect 8053 2377 8233 2400
rect 8053 2360 8090 2377
rect 8053 2326 8054 2360
rect 8088 2343 8090 2360
rect 8124 2360 8162 2377
rect 8124 2343 8126 2360
rect 8088 2326 8126 2343
rect 8160 2343 8162 2360
rect 8196 2360 8233 2377
rect 8196 2343 8198 2360
rect 8160 2326 8198 2343
rect 8232 2326 8233 2360
rect 8053 2309 8233 2326
rect 8053 2286 8090 2309
rect 8053 2252 8054 2286
rect 8088 2275 8090 2286
rect 8124 2286 8162 2309
rect 8124 2275 8126 2286
rect 8088 2252 8126 2275
rect 8160 2275 8162 2286
rect 8196 2286 8233 2309
rect 8196 2275 8198 2286
rect 8160 2252 8198 2275
rect 8232 2252 8233 2286
rect 8053 2241 8233 2252
rect 8053 2212 8090 2241
rect 8053 2178 8054 2212
rect 8088 2207 8090 2212
rect 8124 2212 8162 2241
rect 8124 2207 8126 2212
rect 8088 2178 8126 2207
rect 8160 2207 8162 2212
rect 8196 2212 8233 2241
rect 8196 2207 8198 2212
rect 8160 2178 8198 2207
rect 8232 2178 8233 2212
rect 8053 2173 8233 2178
rect 8053 2139 8090 2173
rect 8124 2139 8162 2173
rect 8196 2139 8233 2173
rect 8053 2138 8233 2139
rect 8053 2104 8054 2138
rect 8088 2105 8126 2138
rect 8088 2104 8090 2105
rect 8053 2071 8090 2104
rect 8124 2104 8126 2105
rect 8160 2105 8198 2138
rect 8160 2104 8162 2105
rect 8124 2071 8162 2104
rect 8196 2104 8198 2105
rect 8232 2104 8233 2138
rect 8196 2071 8233 2104
rect 8053 2064 8233 2071
rect 8053 2030 8054 2064
rect 8088 2037 8126 2064
rect 8088 2030 8090 2037
rect 8053 2003 8090 2030
rect 8124 2030 8126 2037
rect 8160 2037 8198 2064
rect 8160 2030 8162 2037
rect 8124 2003 8162 2030
rect 8196 2030 8198 2037
rect 8232 2030 8233 2064
rect 8196 2003 8233 2030
rect 8053 1990 8233 2003
rect 8053 1956 8054 1990
rect 8088 1969 8126 1990
rect 8088 1956 8090 1969
rect 8053 1935 8090 1956
rect 8124 1956 8126 1969
rect 8160 1969 8198 1990
rect 8160 1956 8162 1969
rect 8124 1935 8162 1956
rect 8196 1956 8198 1969
rect 8232 1956 8233 1990
rect 8196 1935 8233 1956
rect 8053 1916 8233 1935
rect 8053 1882 8054 1916
rect 8088 1901 8126 1916
rect 8088 1882 8090 1901
rect 8053 1867 8090 1882
rect 8124 1882 8126 1901
rect 8160 1901 8198 1916
rect 8160 1882 8162 1901
rect 8124 1867 8162 1882
rect 8196 1882 8198 1901
rect 8232 1882 8233 1916
rect 8196 1867 8233 1882
rect 8053 1842 8233 1867
rect 8053 1808 8054 1842
rect 8088 1833 8126 1842
rect 8088 1808 8090 1833
rect 8053 1799 8090 1808
rect 8124 1808 8126 1833
rect 8160 1833 8198 1842
rect 8160 1808 8162 1833
rect 8124 1799 8162 1808
rect 8196 1808 8198 1833
rect 8232 1808 8233 1842
rect 8196 1799 8233 1808
rect 8053 1768 8233 1799
rect 8053 1734 8054 1768
rect 8088 1765 8126 1768
rect 8088 1734 8090 1765
rect 8053 1731 8090 1734
rect 8124 1734 8126 1765
rect 8160 1765 8198 1768
rect 8160 1734 8162 1765
rect 8124 1731 8162 1734
rect 8196 1734 8198 1765
rect 8232 1734 8233 1768
rect 8196 1731 8233 1734
rect 8053 1697 8233 1731
rect 8053 1694 8090 1697
rect 8053 1660 8054 1694
rect 8088 1663 8090 1694
rect 8124 1694 8162 1697
rect 8124 1663 8126 1694
rect 8088 1660 8126 1663
rect 8160 1663 8162 1694
rect 8196 1694 8233 1697
rect 8196 1663 8198 1694
rect 8160 1660 8198 1663
rect 8232 1660 8233 1694
rect 8053 1629 8233 1660
rect 8053 1620 8090 1629
rect 8053 1586 8054 1620
rect 8088 1595 8090 1620
rect 8124 1620 8162 1629
rect 8124 1595 8126 1620
rect 8088 1586 8126 1595
rect 8160 1595 8162 1620
rect 8196 1620 8233 1629
rect 8196 1595 8198 1620
rect 8160 1586 8198 1595
rect 8232 1586 8233 1620
rect 8053 1561 8233 1586
rect 8053 1545 8090 1561
rect 8053 1511 8054 1545
rect 8088 1527 8090 1545
rect 8124 1545 8162 1561
rect 8124 1527 8126 1545
rect 8088 1511 8126 1527
rect 8160 1527 8162 1545
rect 8196 1545 8233 1561
rect 8196 1527 8198 1545
rect 8160 1511 8198 1527
rect 8232 1511 8233 1545
rect 8298 3010 8418 4106
rect 8860 4388 8867 4494
rect 8973 4388 8980 4494
rect 8860 4214 8980 4388
rect 8860 4180 8903 4214
rect 8937 4180 8980 4214
rect 8860 4140 8980 4180
rect 8860 4106 8903 4140
rect 8937 4106 8980 4140
rect 8298 2976 8341 3010
rect 8375 2976 8418 3010
rect 8298 2932 8418 2976
rect 8298 2898 8341 2932
rect 8375 2898 8418 2932
rect 8298 2854 8418 2898
rect 8298 2820 8341 2854
rect 8375 2820 8418 2854
rect 8298 2776 8418 2820
rect 8298 2742 8341 2776
rect 8375 2742 8418 2776
rect 8298 2697 8418 2742
rect 8298 2663 8341 2697
rect 8375 2663 8418 2697
rect 8298 2618 8418 2663
rect 8298 2584 8341 2618
rect 8375 2584 8418 2618
rect 8298 2539 8418 2584
rect 8298 2505 8341 2539
rect 8375 2505 8418 2539
rect 8090 1491 8196 1511
rect 7868 1375 7911 1409
rect 7945 1375 7988 1409
rect 7868 1335 7988 1375
rect 7868 1301 7911 1335
rect 7945 1301 7988 1335
rect 7868 1285 7988 1301
rect 8298 1409 8418 2505
rect 8520 4050 8622 4062
rect 8656 4050 8758 4062
rect 8520 4046 8550 4050
rect 8728 4046 8758 4050
rect 8520 3978 8550 4012
rect 8728 3978 8758 4012
rect 8520 3910 8550 3944
rect 8728 3910 8758 3944
rect 8520 3842 8550 3876
rect 8728 3842 8758 3876
rect 8520 3774 8550 3808
rect 8728 3774 8758 3808
rect 8520 3706 8550 3740
rect 8728 3706 8758 3740
rect 8520 3638 8550 3672
rect 8728 3638 8758 3672
rect 8520 3570 8550 3604
rect 8728 3570 8758 3604
rect 8520 3502 8550 3536
rect 8728 3502 8758 3536
rect 8520 3434 8550 3468
rect 8728 3434 8758 3468
rect 8520 3366 8550 3400
rect 8728 3366 8758 3400
rect 8520 3298 8550 3332
rect 8728 3298 8758 3332
rect 8520 3230 8550 3264
rect 8728 3230 8758 3264
rect 8520 3162 8550 3196
rect 8728 3162 8758 3196
rect 8520 3080 8550 3128
rect 8584 3080 8694 3092
rect 8728 3080 8758 3128
rect 8520 3040 8758 3080
rect 8520 2574 8550 3040
rect 8728 2574 8758 3040
rect 8520 2535 8758 2574
rect 8520 2501 8550 2535
rect 8584 2501 8622 2535
rect 8656 2501 8694 2535
rect 8728 2501 8758 2535
rect 8520 2461 8758 2501
rect 8520 2449 8622 2461
rect 8656 2449 8758 2461
rect 8520 2445 8550 2449
rect 8728 2445 8758 2449
rect 8520 2377 8550 2411
rect 8728 2377 8758 2411
rect 8520 2309 8550 2343
rect 8728 2309 8758 2343
rect 8520 2241 8550 2275
rect 8728 2241 8758 2275
rect 8520 2173 8550 2207
rect 8728 2173 8758 2207
rect 8520 2105 8550 2139
rect 8728 2105 8758 2139
rect 8520 2037 8550 2071
rect 8728 2037 8758 2071
rect 8520 1969 8550 2003
rect 8728 1969 8758 2003
rect 8520 1901 8550 1935
rect 8728 1901 8758 1935
rect 8520 1833 8550 1867
rect 8728 1833 8758 1867
rect 8520 1765 8550 1799
rect 8728 1765 8758 1799
rect 8520 1697 8550 1731
rect 8728 1697 8758 1731
rect 8520 1629 8550 1663
rect 8728 1629 8758 1663
rect 8520 1561 8550 1595
rect 8728 1561 8758 1595
rect 8520 1479 8550 1527
rect 8584 1479 8694 1491
rect 8728 1479 8758 1527
rect 8520 1464 8758 1479
rect 8860 3010 8980 4106
rect 9290 4388 9297 4494
rect 9403 4388 9410 4494
rect 9290 4214 9410 4388
rect 9290 4180 9333 4214
rect 9367 4180 9410 4214
rect 9290 4140 9410 4180
rect 9290 4106 9333 4140
rect 9367 4106 9410 4140
rect 8860 2976 8903 3010
rect 8937 2976 8980 3010
rect 8860 2932 8980 2976
rect 8860 2898 8903 2932
rect 8937 2898 8980 2932
rect 8860 2854 8980 2898
rect 8860 2820 8903 2854
rect 8937 2820 8980 2854
rect 8860 2776 8980 2820
rect 8860 2742 8903 2776
rect 8937 2742 8980 2776
rect 8860 2697 8980 2742
rect 8860 2663 8903 2697
rect 8937 2663 8980 2697
rect 8860 2618 8980 2663
rect 8860 2584 8903 2618
rect 8937 2584 8980 2618
rect 8860 2539 8980 2584
rect 8860 2505 8903 2539
rect 8937 2505 8980 2539
rect 8298 1375 8341 1409
rect 8375 1375 8418 1409
rect 8298 1335 8418 1375
rect 8298 1301 8341 1335
rect 8375 1301 8418 1335
rect 8298 1285 8418 1301
rect 8860 1409 8980 2505
rect 9045 4028 9046 4062
rect 9080 4046 9118 4062
rect 9080 4028 9082 4046
rect 9045 4012 9082 4028
rect 9116 4028 9118 4046
rect 9152 4046 9190 4062
rect 9152 4028 9154 4046
rect 9116 4012 9154 4028
rect 9188 4028 9190 4046
rect 9224 4028 9225 4062
rect 9188 4012 9225 4028
rect 9045 3988 9225 4012
rect 9045 3954 9046 3988
rect 9080 3978 9118 3988
rect 9080 3954 9082 3978
rect 9045 3944 9082 3954
rect 9116 3954 9118 3978
rect 9152 3978 9190 3988
rect 9152 3954 9154 3978
rect 9116 3944 9154 3954
rect 9188 3954 9190 3978
rect 9224 3954 9225 3988
rect 9188 3944 9225 3954
rect 9045 3914 9225 3944
rect 9045 3880 9046 3914
rect 9080 3910 9118 3914
rect 9080 3880 9082 3910
rect 9045 3876 9082 3880
rect 9116 3880 9118 3910
rect 9152 3910 9190 3914
rect 9152 3880 9154 3910
rect 9116 3876 9154 3880
rect 9188 3880 9190 3910
rect 9224 3880 9225 3914
rect 9188 3876 9225 3880
rect 9045 3842 9225 3876
rect 9045 3840 9082 3842
rect 9045 3806 9046 3840
rect 9080 3808 9082 3840
rect 9116 3840 9154 3842
rect 9116 3808 9118 3840
rect 9080 3806 9118 3808
rect 9152 3808 9154 3840
rect 9188 3840 9225 3842
rect 9188 3808 9190 3840
rect 9152 3806 9190 3808
rect 9224 3806 9225 3840
rect 9045 3774 9225 3806
rect 9045 3766 9082 3774
rect 9045 3732 9046 3766
rect 9080 3740 9082 3766
rect 9116 3766 9154 3774
rect 9116 3740 9118 3766
rect 9080 3732 9118 3740
rect 9152 3740 9154 3766
rect 9188 3766 9225 3774
rect 9188 3740 9190 3766
rect 9152 3732 9190 3740
rect 9224 3732 9225 3766
rect 9045 3706 9225 3732
rect 9045 3692 9082 3706
rect 9045 3658 9046 3692
rect 9080 3672 9082 3692
rect 9116 3692 9154 3706
rect 9116 3672 9118 3692
rect 9080 3658 9118 3672
rect 9152 3672 9154 3692
rect 9188 3692 9225 3706
rect 9188 3672 9190 3692
rect 9152 3658 9190 3672
rect 9224 3658 9225 3692
rect 9045 3638 9225 3658
rect 9045 3618 9082 3638
rect 9045 3584 9046 3618
rect 9080 3604 9082 3618
rect 9116 3618 9154 3638
rect 9116 3604 9118 3618
rect 9080 3584 9118 3604
rect 9152 3604 9154 3618
rect 9188 3618 9225 3638
rect 9188 3604 9190 3618
rect 9152 3584 9190 3604
rect 9224 3584 9225 3618
rect 9045 3570 9225 3584
rect 9045 3544 9082 3570
rect 9045 3510 9046 3544
rect 9080 3536 9082 3544
rect 9116 3544 9154 3570
rect 9116 3536 9118 3544
rect 9080 3510 9118 3536
rect 9152 3536 9154 3544
rect 9188 3544 9225 3570
rect 9188 3536 9190 3544
rect 9152 3510 9190 3536
rect 9224 3510 9225 3544
rect 9045 3502 9225 3510
rect 9045 3470 9082 3502
rect 9045 3436 9046 3470
rect 9080 3468 9082 3470
rect 9116 3470 9154 3502
rect 9116 3468 9118 3470
rect 9080 3436 9118 3468
rect 9152 3468 9154 3470
rect 9188 3470 9225 3502
rect 9188 3468 9190 3470
rect 9152 3436 9190 3468
rect 9224 3436 9225 3470
rect 9045 3434 9225 3436
rect 9045 3400 9082 3434
rect 9116 3400 9154 3434
rect 9188 3400 9225 3434
rect 9045 3396 9225 3400
rect 9045 3362 9046 3396
rect 9080 3366 9118 3396
rect 9080 3362 9082 3366
rect 9045 3332 9082 3362
rect 9116 3362 9118 3366
rect 9152 3366 9190 3396
rect 9152 3362 9154 3366
rect 9116 3332 9154 3362
rect 9188 3362 9190 3366
rect 9224 3362 9225 3396
rect 9188 3332 9225 3362
rect 9045 3322 9225 3332
rect 9045 3288 9046 3322
rect 9080 3298 9118 3322
rect 9080 3288 9082 3298
rect 9045 3264 9082 3288
rect 9116 3288 9118 3298
rect 9152 3298 9190 3322
rect 9152 3288 9154 3298
rect 9116 3264 9154 3288
rect 9188 3288 9190 3298
rect 9224 3288 9225 3322
rect 9188 3264 9225 3288
rect 9045 3248 9225 3264
rect 9045 3214 9046 3248
rect 9080 3230 9118 3248
rect 9080 3214 9082 3230
rect 9045 3196 9082 3214
rect 9116 3214 9118 3230
rect 9152 3230 9190 3248
rect 9152 3214 9154 3230
rect 9116 3196 9154 3214
rect 9188 3214 9190 3230
rect 9224 3214 9225 3248
rect 9188 3196 9225 3214
rect 9045 3174 9225 3196
rect 9045 3140 9046 3174
rect 9080 3162 9118 3174
rect 9080 3140 9082 3162
rect 9045 3128 9082 3140
rect 9116 3140 9118 3162
rect 9152 3162 9190 3174
rect 9152 3140 9154 3162
rect 9116 3128 9154 3140
rect 9188 3140 9190 3162
rect 9224 3140 9225 3174
rect 9188 3128 9225 3140
rect 9045 3100 9225 3128
rect 9045 3066 9046 3100
rect 9080 3066 9118 3100
rect 9152 3066 9190 3100
rect 9224 3066 9225 3100
rect 9045 3026 9225 3066
rect 9045 2992 9046 3026
rect 9080 2992 9118 3026
rect 9152 2992 9190 3026
rect 9224 2992 9225 3026
rect 9045 2952 9225 2992
rect 9045 2918 9046 2952
rect 9080 2918 9118 2952
rect 9152 2918 9190 2952
rect 9224 2918 9225 2952
rect 9045 2878 9225 2918
rect 9045 2844 9046 2878
rect 9080 2844 9118 2878
rect 9152 2844 9190 2878
rect 9224 2844 9225 2878
rect 9045 2804 9225 2844
rect 9045 2770 9046 2804
rect 9080 2770 9118 2804
rect 9152 2770 9190 2804
rect 9224 2770 9225 2804
rect 9045 2730 9225 2770
rect 9045 2696 9046 2730
rect 9080 2696 9118 2730
rect 9152 2696 9190 2730
rect 9224 2696 9225 2730
rect 9045 2656 9225 2696
rect 9045 2622 9046 2656
rect 9080 2622 9118 2656
rect 9152 2622 9190 2656
rect 9224 2622 9225 2656
rect 9045 2582 9225 2622
rect 9045 2548 9046 2582
rect 9080 2548 9118 2582
rect 9152 2548 9190 2582
rect 9224 2548 9225 2582
rect 9045 2508 9225 2548
rect 9045 2474 9046 2508
rect 9080 2474 9118 2508
rect 9152 2474 9190 2508
rect 9224 2474 9225 2508
rect 9045 2445 9225 2474
rect 9045 2434 9082 2445
rect 9045 2400 9046 2434
rect 9080 2411 9082 2434
rect 9116 2434 9154 2445
rect 9116 2411 9118 2434
rect 9080 2400 9118 2411
rect 9152 2411 9154 2434
rect 9188 2434 9225 2445
rect 9188 2411 9190 2434
rect 9152 2400 9190 2411
rect 9224 2400 9225 2434
rect 9045 2377 9225 2400
rect 9045 2360 9082 2377
rect 9045 2326 9046 2360
rect 9080 2343 9082 2360
rect 9116 2360 9154 2377
rect 9116 2343 9118 2360
rect 9080 2326 9118 2343
rect 9152 2343 9154 2360
rect 9188 2360 9225 2377
rect 9188 2343 9190 2360
rect 9152 2326 9190 2343
rect 9224 2326 9225 2360
rect 9045 2309 9225 2326
rect 9045 2286 9082 2309
rect 9045 2252 9046 2286
rect 9080 2275 9082 2286
rect 9116 2286 9154 2309
rect 9116 2275 9118 2286
rect 9080 2252 9118 2275
rect 9152 2275 9154 2286
rect 9188 2286 9225 2309
rect 9188 2275 9190 2286
rect 9152 2252 9190 2275
rect 9224 2252 9225 2286
rect 9045 2241 9225 2252
rect 9045 2212 9082 2241
rect 9045 2178 9046 2212
rect 9080 2207 9082 2212
rect 9116 2212 9154 2241
rect 9116 2207 9118 2212
rect 9080 2178 9118 2207
rect 9152 2207 9154 2212
rect 9188 2212 9225 2241
rect 9188 2207 9190 2212
rect 9152 2178 9190 2207
rect 9224 2178 9225 2212
rect 9045 2173 9225 2178
rect 9045 2139 9082 2173
rect 9116 2139 9154 2173
rect 9188 2139 9225 2173
rect 9045 2138 9225 2139
rect 9045 2104 9046 2138
rect 9080 2105 9118 2138
rect 9080 2104 9082 2105
rect 9045 2071 9082 2104
rect 9116 2104 9118 2105
rect 9152 2105 9190 2138
rect 9152 2104 9154 2105
rect 9116 2071 9154 2104
rect 9188 2104 9190 2105
rect 9224 2104 9225 2138
rect 9188 2071 9225 2104
rect 9045 2064 9225 2071
rect 9045 2030 9046 2064
rect 9080 2037 9118 2064
rect 9080 2030 9082 2037
rect 9045 2003 9082 2030
rect 9116 2030 9118 2037
rect 9152 2037 9190 2064
rect 9152 2030 9154 2037
rect 9116 2003 9154 2030
rect 9188 2030 9190 2037
rect 9224 2030 9225 2064
rect 9188 2003 9225 2030
rect 9045 1990 9225 2003
rect 9045 1956 9046 1990
rect 9080 1969 9118 1990
rect 9080 1956 9082 1969
rect 9045 1935 9082 1956
rect 9116 1956 9118 1969
rect 9152 1969 9190 1990
rect 9152 1956 9154 1969
rect 9116 1935 9154 1956
rect 9188 1956 9190 1969
rect 9224 1956 9225 1990
rect 9188 1935 9225 1956
rect 9045 1916 9225 1935
rect 9045 1882 9046 1916
rect 9080 1901 9118 1916
rect 9080 1882 9082 1901
rect 9045 1867 9082 1882
rect 9116 1882 9118 1901
rect 9152 1901 9190 1916
rect 9152 1882 9154 1901
rect 9116 1867 9154 1882
rect 9188 1882 9190 1901
rect 9224 1882 9225 1916
rect 9188 1867 9225 1882
rect 9045 1842 9225 1867
rect 9045 1808 9046 1842
rect 9080 1833 9118 1842
rect 9080 1808 9082 1833
rect 9045 1799 9082 1808
rect 9116 1808 9118 1833
rect 9152 1833 9190 1842
rect 9152 1808 9154 1833
rect 9116 1799 9154 1808
rect 9188 1808 9190 1833
rect 9224 1808 9225 1842
rect 9188 1799 9225 1808
rect 9045 1768 9225 1799
rect 9045 1734 9046 1768
rect 9080 1765 9118 1768
rect 9080 1734 9082 1765
rect 9045 1731 9082 1734
rect 9116 1734 9118 1765
rect 9152 1765 9190 1768
rect 9152 1734 9154 1765
rect 9116 1731 9154 1734
rect 9188 1734 9190 1765
rect 9224 1734 9225 1768
rect 9188 1731 9225 1734
rect 9045 1697 9225 1731
rect 9045 1694 9082 1697
rect 9045 1660 9046 1694
rect 9080 1663 9082 1694
rect 9116 1694 9154 1697
rect 9116 1663 9118 1694
rect 9080 1660 9118 1663
rect 9152 1663 9154 1694
rect 9188 1694 9225 1697
rect 9188 1663 9190 1694
rect 9152 1660 9190 1663
rect 9224 1660 9225 1694
rect 9045 1629 9225 1660
rect 9045 1620 9082 1629
rect 9045 1586 9046 1620
rect 9080 1595 9082 1620
rect 9116 1620 9154 1629
rect 9116 1595 9118 1620
rect 9080 1586 9118 1595
rect 9152 1595 9154 1620
rect 9188 1620 9225 1629
rect 9188 1595 9190 1620
rect 9152 1586 9190 1595
rect 9224 1586 9225 1620
rect 9045 1561 9225 1586
rect 9045 1545 9082 1561
rect 9045 1511 9046 1545
rect 9080 1527 9082 1545
rect 9116 1545 9154 1561
rect 9116 1527 9118 1545
rect 9080 1511 9118 1527
rect 9152 1527 9154 1545
rect 9188 1545 9225 1561
rect 9188 1527 9190 1545
rect 9152 1511 9190 1527
rect 9224 1511 9225 1545
rect 9290 3010 9410 4106
rect 9852 4388 9859 4494
rect 9965 4388 9972 4494
rect 9852 4214 9972 4388
rect 9852 4180 9895 4214
rect 9929 4180 9972 4214
rect 9852 4140 9972 4180
rect 9852 4106 9895 4140
rect 9929 4106 9972 4140
rect 9290 2976 9333 3010
rect 9367 2976 9410 3010
rect 9290 2932 9410 2976
rect 9290 2898 9333 2932
rect 9367 2898 9410 2932
rect 9290 2854 9410 2898
rect 9290 2820 9333 2854
rect 9367 2820 9410 2854
rect 9290 2776 9410 2820
rect 9290 2742 9333 2776
rect 9367 2742 9410 2776
rect 9290 2697 9410 2742
rect 9290 2663 9333 2697
rect 9367 2663 9410 2697
rect 9290 2618 9410 2663
rect 9290 2584 9333 2618
rect 9367 2584 9410 2618
rect 9290 2539 9410 2584
rect 9290 2505 9333 2539
rect 9367 2505 9410 2539
rect 9082 1491 9188 1511
rect 8860 1375 8903 1409
rect 8937 1375 8980 1409
rect 8860 1335 8980 1375
rect 8860 1301 8903 1335
rect 8937 1301 8980 1335
rect 8860 1285 8980 1301
rect 9290 1409 9410 2505
rect 9512 4050 9614 4062
rect 9648 4050 9750 4062
rect 9512 4046 9542 4050
rect 9720 4046 9750 4050
rect 9512 3978 9542 4012
rect 9720 3978 9750 4012
rect 9512 3910 9542 3944
rect 9720 3910 9750 3944
rect 9512 3842 9542 3876
rect 9720 3842 9750 3876
rect 9512 3774 9542 3808
rect 9720 3774 9750 3808
rect 9512 3706 9542 3740
rect 9720 3706 9750 3740
rect 9512 3638 9542 3672
rect 9720 3638 9750 3672
rect 9512 3570 9542 3604
rect 9720 3570 9750 3604
rect 9512 3502 9542 3536
rect 9720 3502 9750 3536
rect 9512 3434 9542 3468
rect 9720 3434 9750 3468
rect 9512 3366 9542 3400
rect 9720 3366 9750 3400
rect 9512 3298 9542 3332
rect 9720 3298 9750 3332
rect 9512 3230 9542 3264
rect 9720 3230 9750 3264
rect 9512 3162 9542 3196
rect 9720 3162 9750 3196
rect 9512 3080 9542 3128
rect 9576 3080 9686 3092
rect 9720 3080 9750 3128
rect 9512 3040 9750 3080
rect 9512 2574 9542 3040
rect 9720 2574 9750 3040
rect 9512 2535 9750 2574
rect 9512 2501 9542 2535
rect 9576 2501 9614 2535
rect 9648 2501 9686 2535
rect 9720 2501 9750 2535
rect 9512 2461 9750 2501
rect 9512 2449 9614 2461
rect 9648 2449 9750 2461
rect 9512 2445 9542 2449
rect 9720 2445 9750 2449
rect 9512 2377 9542 2411
rect 9720 2377 9750 2411
rect 9512 2309 9542 2343
rect 9720 2309 9750 2343
rect 9512 2241 9542 2275
rect 9720 2241 9750 2275
rect 9512 2173 9542 2207
rect 9720 2173 9750 2207
rect 9512 2105 9542 2139
rect 9720 2105 9750 2139
rect 9512 2037 9542 2071
rect 9720 2037 9750 2071
rect 9512 1969 9542 2003
rect 9720 1969 9750 2003
rect 9512 1901 9542 1935
rect 9720 1901 9750 1935
rect 9512 1833 9542 1867
rect 9720 1833 9750 1867
rect 9512 1765 9542 1799
rect 9720 1765 9750 1799
rect 9512 1697 9542 1731
rect 9720 1697 9750 1731
rect 9512 1629 9542 1663
rect 9720 1629 9750 1663
rect 9512 1561 9542 1595
rect 9720 1561 9750 1595
rect 9512 1479 9542 1527
rect 9576 1479 9686 1491
rect 9720 1479 9750 1527
rect 9512 1464 9750 1479
rect 9852 3010 9972 4106
rect 10282 4388 10289 4494
rect 10395 4388 10402 4494
rect 10282 4214 10402 4388
rect 10282 4180 10325 4214
rect 10359 4180 10402 4214
rect 10282 4140 10402 4180
rect 10282 4106 10325 4140
rect 10359 4106 10402 4140
rect 9852 2976 9895 3010
rect 9929 2976 9972 3010
rect 9852 2932 9972 2976
rect 9852 2898 9895 2932
rect 9929 2898 9972 2932
rect 9852 2854 9972 2898
rect 9852 2820 9895 2854
rect 9929 2820 9972 2854
rect 9852 2776 9972 2820
rect 9852 2742 9895 2776
rect 9929 2742 9972 2776
rect 9852 2697 9972 2742
rect 9852 2663 9895 2697
rect 9929 2663 9972 2697
rect 9852 2618 9972 2663
rect 9852 2584 9895 2618
rect 9929 2584 9972 2618
rect 9852 2539 9972 2584
rect 9852 2505 9895 2539
rect 9929 2505 9972 2539
rect 9290 1375 9333 1409
rect 9367 1375 9410 1409
rect 9290 1335 9410 1375
rect 9290 1301 9333 1335
rect 9367 1301 9410 1335
rect 9290 1285 9410 1301
rect 9852 1409 9972 2505
rect 10037 4028 10038 4062
rect 10072 4046 10110 4062
rect 10072 4028 10074 4046
rect 10037 4012 10074 4028
rect 10108 4028 10110 4046
rect 10144 4046 10182 4062
rect 10144 4028 10146 4046
rect 10108 4012 10146 4028
rect 10180 4028 10182 4046
rect 10216 4028 10217 4062
rect 10180 4012 10217 4028
rect 10037 3988 10217 4012
rect 10037 3954 10038 3988
rect 10072 3978 10110 3988
rect 10072 3954 10074 3978
rect 10037 3944 10074 3954
rect 10108 3954 10110 3978
rect 10144 3978 10182 3988
rect 10144 3954 10146 3978
rect 10108 3944 10146 3954
rect 10180 3954 10182 3978
rect 10216 3954 10217 3988
rect 10180 3944 10217 3954
rect 10037 3914 10217 3944
rect 10037 3880 10038 3914
rect 10072 3910 10110 3914
rect 10072 3880 10074 3910
rect 10037 3876 10074 3880
rect 10108 3880 10110 3910
rect 10144 3910 10182 3914
rect 10144 3880 10146 3910
rect 10108 3876 10146 3880
rect 10180 3880 10182 3910
rect 10216 3880 10217 3914
rect 10180 3876 10217 3880
rect 10037 3842 10217 3876
rect 10037 3840 10074 3842
rect 10037 3806 10038 3840
rect 10072 3808 10074 3840
rect 10108 3840 10146 3842
rect 10108 3808 10110 3840
rect 10072 3806 10110 3808
rect 10144 3808 10146 3840
rect 10180 3840 10217 3842
rect 10180 3808 10182 3840
rect 10144 3806 10182 3808
rect 10216 3806 10217 3840
rect 10037 3774 10217 3806
rect 10037 3766 10074 3774
rect 10037 3732 10038 3766
rect 10072 3740 10074 3766
rect 10108 3766 10146 3774
rect 10108 3740 10110 3766
rect 10072 3732 10110 3740
rect 10144 3740 10146 3766
rect 10180 3766 10217 3774
rect 10180 3740 10182 3766
rect 10144 3732 10182 3740
rect 10216 3732 10217 3766
rect 10037 3706 10217 3732
rect 10037 3692 10074 3706
rect 10037 3658 10038 3692
rect 10072 3672 10074 3692
rect 10108 3692 10146 3706
rect 10108 3672 10110 3692
rect 10072 3658 10110 3672
rect 10144 3672 10146 3692
rect 10180 3692 10217 3706
rect 10180 3672 10182 3692
rect 10144 3658 10182 3672
rect 10216 3658 10217 3692
rect 10037 3638 10217 3658
rect 10037 3618 10074 3638
rect 10037 3584 10038 3618
rect 10072 3604 10074 3618
rect 10108 3618 10146 3638
rect 10108 3604 10110 3618
rect 10072 3584 10110 3604
rect 10144 3604 10146 3618
rect 10180 3618 10217 3638
rect 10180 3604 10182 3618
rect 10144 3584 10182 3604
rect 10216 3584 10217 3618
rect 10037 3570 10217 3584
rect 10037 3544 10074 3570
rect 10037 3510 10038 3544
rect 10072 3536 10074 3544
rect 10108 3544 10146 3570
rect 10108 3536 10110 3544
rect 10072 3510 10110 3536
rect 10144 3536 10146 3544
rect 10180 3544 10217 3570
rect 10180 3536 10182 3544
rect 10144 3510 10182 3536
rect 10216 3510 10217 3544
rect 10037 3502 10217 3510
rect 10037 3470 10074 3502
rect 10037 3436 10038 3470
rect 10072 3468 10074 3470
rect 10108 3470 10146 3502
rect 10108 3468 10110 3470
rect 10072 3436 10110 3468
rect 10144 3468 10146 3470
rect 10180 3470 10217 3502
rect 10180 3468 10182 3470
rect 10144 3436 10182 3468
rect 10216 3436 10217 3470
rect 10037 3434 10217 3436
rect 10037 3400 10074 3434
rect 10108 3400 10146 3434
rect 10180 3400 10217 3434
rect 10037 3396 10217 3400
rect 10037 3362 10038 3396
rect 10072 3366 10110 3396
rect 10072 3362 10074 3366
rect 10037 3332 10074 3362
rect 10108 3362 10110 3366
rect 10144 3366 10182 3396
rect 10144 3362 10146 3366
rect 10108 3332 10146 3362
rect 10180 3362 10182 3366
rect 10216 3362 10217 3396
rect 10180 3332 10217 3362
rect 10037 3322 10217 3332
rect 10037 3288 10038 3322
rect 10072 3298 10110 3322
rect 10072 3288 10074 3298
rect 10037 3264 10074 3288
rect 10108 3288 10110 3298
rect 10144 3298 10182 3322
rect 10144 3288 10146 3298
rect 10108 3264 10146 3288
rect 10180 3288 10182 3298
rect 10216 3288 10217 3322
rect 10180 3264 10217 3288
rect 10037 3248 10217 3264
rect 10037 3214 10038 3248
rect 10072 3230 10110 3248
rect 10072 3214 10074 3230
rect 10037 3196 10074 3214
rect 10108 3214 10110 3230
rect 10144 3230 10182 3248
rect 10144 3214 10146 3230
rect 10108 3196 10146 3214
rect 10180 3214 10182 3230
rect 10216 3214 10217 3248
rect 10180 3196 10217 3214
rect 10037 3174 10217 3196
rect 10037 3140 10038 3174
rect 10072 3162 10110 3174
rect 10072 3140 10074 3162
rect 10037 3128 10074 3140
rect 10108 3140 10110 3162
rect 10144 3162 10182 3174
rect 10144 3140 10146 3162
rect 10108 3128 10146 3140
rect 10180 3140 10182 3162
rect 10216 3140 10217 3174
rect 10180 3128 10217 3140
rect 10037 3100 10217 3128
rect 10037 3066 10038 3100
rect 10072 3066 10110 3100
rect 10144 3066 10182 3100
rect 10216 3066 10217 3100
rect 10037 3026 10217 3066
rect 10037 2992 10038 3026
rect 10072 2992 10110 3026
rect 10144 2992 10182 3026
rect 10216 2992 10217 3026
rect 10037 2952 10217 2992
rect 10037 2918 10038 2952
rect 10072 2918 10110 2952
rect 10144 2918 10182 2952
rect 10216 2918 10217 2952
rect 10037 2878 10217 2918
rect 10037 2844 10038 2878
rect 10072 2844 10110 2878
rect 10144 2844 10182 2878
rect 10216 2844 10217 2878
rect 10037 2804 10217 2844
rect 10037 2770 10038 2804
rect 10072 2770 10110 2804
rect 10144 2770 10182 2804
rect 10216 2770 10217 2804
rect 10037 2730 10217 2770
rect 10037 2696 10038 2730
rect 10072 2696 10110 2730
rect 10144 2696 10182 2730
rect 10216 2696 10217 2730
rect 10037 2656 10217 2696
rect 10037 2622 10038 2656
rect 10072 2622 10110 2656
rect 10144 2622 10182 2656
rect 10216 2622 10217 2656
rect 10037 2582 10217 2622
rect 10037 2548 10038 2582
rect 10072 2548 10110 2582
rect 10144 2548 10182 2582
rect 10216 2548 10217 2582
rect 10037 2508 10217 2548
rect 10037 2474 10038 2508
rect 10072 2474 10110 2508
rect 10144 2474 10182 2508
rect 10216 2474 10217 2508
rect 10037 2445 10217 2474
rect 10037 2434 10074 2445
rect 10037 2400 10038 2434
rect 10072 2411 10074 2434
rect 10108 2434 10146 2445
rect 10108 2411 10110 2434
rect 10072 2400 10110 2411
rect 10144 2411 10146 2434
rect 10180 2434 10217 2445
rect 10180 2411 10182 2434
rect 10144 2400 10182 2411
rect 10216 2400 10217 2434
rect 10037 2377 10217 2400
rect 10037 2360 10074 2377
rect 10037 2326 10038 2360
rect 10072 2343 10074 2360
rect 10108 2360 10146 2377
rect 10108 2343 10110 2360
rect 10072 2326 10110 2343
rect 10144 2343 10146 2360
rect 10180 2360 10217 2377
rect 10180 2343 10182 2360
rect 10144 2326 10182 2343
rect 10216 2326 10217 2360
rect 10037 2309 10217 2326
rect 10037 2286 10074 2309
rect 10037 2252 10038 2286
rect 10072 2275 10074 2286
rect 10108 2286 10146 2309
rect 10108 2275 10110 2286
rect 10072 2252 10110 2275
rect 10144 2275 10146 2286
rect 10180 2286 10217 2309
rect 10180 2275 10182 2286
rect 10144 2252 10182 2275
rect 10216 2252 10217 2286
rect 10037 2241 10217 2252
rect 10037 2212 10074 2241
rect 10037 2178 10038 2212
rect 10072 2207 10074 2212
rect 10108 2212 10146 2241
rect 10108 2207 10110 2212
rect 10072 2178 10110 2207
rect 10144 2207 10146 2212
rect 10180 2212 10217 2241
rect 10180 2207 10182 2212
rect 10144 2178 10182 2207
rect 10216 2178 10217 2212
rect 10037 2173 10217 2178
rect 10037 2139 10074 2173
rect 10108 2139 10146 2173
rect 10180 2139 10217 2173
rect 10037 2138 10217 2139
rect 10037 2104 10038 2138
rect 10072 2105 10110 2138
rect 10072 2104 10074 2105
rect 10037 2071 10074 2104
rect 10108 2104 10110 2105
rect 10144 2105 10182 2138
rect 10144 2104 10146 2105
rect 10108 2071 10146 2104
rect 10180 2104 10182 2105
rect 10216 2104 10217 2138
rect 10180 2071 10217 2104
rect 10037 2064 10217 2071
rect 10037 2030 10038 2064
rect 10072 2037 10110 2064
rect 10072 2030 10074 2037
rect 10037 2003 10074 2030
rect 10108 2030 10110 2037
rect 10144 2037 10182 2064
rect 10144 2030 10146 2037
rect 10108 2003 10146 2030
rect 10180 2030 10182 2037
rect 10216 2030 10217 2064
rect 10180 2003 10217 2030
rect 10037 1990 10217 2003
rect 10037 1956 10038 1990
rect 10072 1969 10110 1990
rect 10072 1956 10074 1969
rect 10037 1935 10074 1956
rect 10108 1956 10110 1969
rect 10144 1969 10182 1990
rect 10144 1956 10146 1969
rect 10108 1935 10146 1956
rect 10180 1956 10182 1969
rect 10216 1956 10217 1990
rect 10180 1935 10217 1956
rect 10037 1916 10217 1935
rect 10037 1882 10038 1916
rect 10072 1901 10110 1916
rect 10072 1882 10074 1901
rect 10037 1867 10074 1882
rect 10108 1882 10110 1901
rect 10144 1901 10182 1916
rect 10144 1882 10146 1901
rect 10108 1867 10146 1882
rect 10180 1882 10182 1901
rect 10216 1882 10217 1916
rect 10180 1867 10217 1882
rect 10037 1842 10217 1867
rect 10037 1808 10038 1842
rect 10072 1833 10110 1842
rect 10072 1808 10074 1833
rect 10037 1799 10074 1808
rect 10108 1808 10110 1833
rect 10144 1833 10182 1842
rect 10144 1808 10146 1833
rect 10108 1799 10146 1808
rect 10180 1808 10182 1833
rect 10216 1808 10217 1842
rect 10180 1799 10217 1808
rect 10037 1768 10217 1799
rect 10037 1734 10038 1768
rect 10072 1765 10110 1768
rect 10072 1734 10074 1765
rect 10037 1731 10074 1734
rect 10108 1734 10110 1765
rect 10144 1765 10182 1768
rect 10144 1734 10146 1765
rect 10108 1731 10146 1734
rect 10180 1734 10182 1765
rect 10216 1734 10217 1768
rect 10180 1731 10217 1734
rect 10037 1697 10217 1731
rect 10037 1694 10074 1697
rect 10037 1660 10038 1694
rect 10072 1663 10074 1694
rect 10108 1694 10146 1697
rect 10108 1663 10110 1694
rect 10072 1660 10110 1663
rect 10144 1663 10146 1694
rect 10180 1694 10217 1697
rect 10180 1663 10182 1694
rect 10144 1660 10182 1663
rect 10216 1660 10217 1694
rect 10037 1629 10217 1660
rect 10037 1620 10074 1629
rect 10037 1586 10038 1620
rect 10072 1595 10074 1620
rect 10108 1620 10146 1629
rect 10108 1595 10110 1620
rect 10072 1586 10110 1595
rect 10144 1595 10146 1620
rect 10180 1620 10217 1629
rect 10180 1595 10182 1620
rect 10144 1586 10182 1595
rect 10216 1586 10217 1620
rect 10037 1561 10217 1586
rect 10037 1545 10074 1561
rect 10037 1511 10038 1545
rect 10072 1527 10074 1545
rect 10108 1545 10146 1561
rect 10108 1527 10110 1545
rect 10072 1511 10110 1527
rect 10144 1527 10146 1545
rect 10180 1545 10217 1561
rect 10180 1527 10182 1545
rect 10144 1511 10182 1527
rect 10216 1511 10217 1545
rect 10282 3010 10402 4106
rect 10844 4388 10851 4494
rect 10957 4388 10964 4494
rect 10844 4214 10964 4388
rect 10844 4180 10887 4214
rect 10921 4180 10964 4214
rect 10844 4140 10964 4180
rect 10844 4106 10887 4140
rect 10921 4106 10964 4140
rect 10282 2976 10325 3010
rect 10359 2976 10402 3010
rect 10282 2932 10402 2976
rect 10282 2898 10325 2932
rect 10359 2898 10402 2932
rect 10282 2854 10402 2898
rect 10282 2820 10325 2854
rect 10359 2820 10402 2854
rect 10282 2776 10402 2820
rect 10282 2742 10325 2776
rect 10359 2742 10402 2776
rect 10282 2697 10402 2742
rect 10282 2663 10325 2697
rect 10359 2663 10402 2697
rect 10282 2618 10402 2663
rect 10282 2584 10325 2618
rect 10359 2584 10402 2618
rect 10282 2539 10402 2584
rect 10282 2505 10325 2539
rect 10359 2505 10402 2539
rect 10074 1491 10180 1511
rect 9852 1375 9895 1409
rect 9929 1375 9972 1409
rect 9852 1335 9972 1375
rect 9852 1301 9895 1335
rect 9929 1301 9972 1335
rect 9852 1285 9972 1301
rect 10282 1409 10402 2505
rect 10504 4050 10606 4062
rect 10640 4050 10742 4062
rect 10504 4046 10534 4050
rect 10712 4046 10742 4050
rect 10504 3978 10534 4012
rect 10712 3978 10742 4012
rect 10504 3910 10534 3944
rect 10712 3910 10742 3944
rect 10504 3842 10534 3876
rect 10712 3842 10742 3876
rect 10504 3774 10534 3808
rect 10712 3774 10742 3808
rect 10504 3706 10534 3740
rect 10712 3706 10742 3740
rect 10504 3638 10534 3672
rect 10712 3638 10742 3672
rect 10504 3570 10534 3604
rect 10712 3570 10742 3604
rect 10504 3502 10534 3536
rect 10712 3502 10742 3536
rect 10504 3434 10534 3468
rect 10712 3434 10742 3468
rect 10504 3366 10534 3400
rect 10712 3366 10742 3400
rect 10504 3298 10534 3332
rect 10712 3298 10742 3332
rect 10504 3230 10534 3264
rect 10712 3230 10742 3264
rect 10504 3162 10534 3196
rect 10712 3162 10742 3196
rect 10504 3080 10534 3128
rect 10568 3080 10678 3092
rect 10712 3080 10742 3128
rect 10504 3037 10742 3080
rect 10504 3003 10534 3037
rect 10568 3003 10606 3037
rect 10640 3003 10678 3037
rect 10712 3003 10742 3037
rect 10504 2954 10742 3003
rect 10504 2920 10534 2954
rect 10568 2935 10606 2954
rect 10640 2935 10678 2954
rect 10568 2920 10573 2935
rect 10640 2920 10641 2935
rect 10504 2901 10573 2920
rect 10607 2901 10641 2920
rect 10675 2920 10678 2935
rect 10712 2920 10742 2954
rect 10675 2901 10742 2920
rect 10504 2871 10742 2901
rect 10504 2837 10534 2871
rect 10568 2855 10606 2871
rect 10640 2855 10678 2871
rect 10568 2837 10573 2855
rect 10640 2837 10641 2855
rect 10504 2821 10573 2837
rect 10607 2821 10641 2837
rect 10675 2837 10678 2855
rect 10712 2837 10742 2871
rect 10675 2821 10742 2837
rect 10504 2787 10742 2821
rect 10504 2753 10534 2787
rect 10568 2775 10606 2787
rect 10640 2775 10678 2787
rect 10568 2753 10573 2775
rect 10640 2753 10641 2775
rect 10504 2741 10573 2753
rect 10607 2741 10641 2753
rect 10675 2753 10678 2775
rect 10712 2753 10742 2787
rect 10675 2741 10742 2753
rect 10504 2703 10742 2741
rect 10504 2669 10534 2703
rect 10568 2695 10606 2703
rect 10640 2695 10678 2703
rect 10568 2669 10573 2695
rect 10640 2669 10641 2695
rect 10504 2661 10573 2669
rect 10607 2661 10641 2669
rect 10675 2669 10678 2695
rect 10712 2669 10742 2703
rect 10675 2661 10742 2669
rect 10504 2619 10742 2661
rect 10504 2585 10534 2619
rect 10568 2614 10606 2619
rect 10640 2614 10678 2619
rect 10568 2585 10573 2614
rect 10640 2585 10641 2614
rect 10504 2580 10573 2585
rect 10607 2580 10641 2585
rect 10675 2585 10678 2614
rect 10712 2585 10742 2619
rect 10675 2580 10742 2585
rect 10504 2535 10742 2580
rect 10504 2501 10534 2535
rect 10568 2501 10606 2535
rect 10640 2501 10678 2535
rect 10712 2501 10742 2535
rect 10504 2461 10742 2501
rect 10504 2449 10606 2461
rect 10640 2449 10742 2461
rect 10504 2445 10534 2449
rect 10712 2445 10742 2449
rect 10504 2377 10534 2411
rect 10712 2377 10742 2411
rect 10504 2309 10534 2343
rect 10712 2309 10742 2343
rect 10504 2241 10534 2275
rect 10712 2241 10742 2275
rect 10504 2173 10534 2207
rect 10712 2173 10742 2207
rect 10504 2105 10534 2139
rect 10712 2105 10742 2139
rect 10504 2037 10534 2071
rect 10712 2037 10742 2071
rect 10504 1969 10534 2003
rect 10712 1969 10742 2003
rect 10504 1901 10534 1935
rect 10712 1901 10742 1935
rect 10504 1833 10534 1867
rect 10712 1833 10742 1867
rect 10504 1765 10534 1799
rect 10712 1765 10742 1799
rect 10504 1697 10534 1731
rect 10712 1697 10742 1731
rect 10504 1629 10534 1663
rect 10712 1629 10742 1663
rect 10504 1561 10534 1595
rect 10712 1561 10742 1595
rect 10504 1479 10534 1527
rect 10568 1479 10678 1491
rect 10712 1479 10742 1527
rect 10504 1464 10742 1479
rect 10844 3010 10964 4106
rect 11274 4388 11281 4494
rect 11387 4388 11394 4494
rect 11274 4214 11394 4388
rect 11274 4180 11317 4214
rect 11351 4180 11394 4214
rect 11274 4140 11394 4180
rect 11274 4106 11317 4140
rect 11351 4106 11394 4140
rect 10844 2976 10887 3010
rect 10921 2976 10964 3010
rect 10844 2932 10964 2976
rect 10844 2898 10887 2932
rect 10921 2898 10964 2932
rect 10844 2854 10964 2898
rect 10844 2820 10887 2854
rect 10921 2820 10964 2854
rect 10844 2776 10964 2820
rect 10844 2742 10887 2776
rect 10921 2742 10964 2776
rect 10844 2697 10964 2742
rect 10844 2663 10887 2697
rect 10921 2663 10964 2697
rect 10844 2618 10964 2663
rect 10844 2584 10887 2618
rect 10921 2584 10964 2618
rect 10844 2539 10964 2584
rect 10844 2505 10887 2539
rect 10921 2505 10964 2539
rect 10282 1375 10325 1409
rect 10359 1375 10402 1409
rect 10282 1335 10402 1375
rect 10282 1301 10325 1335
rect 10359 1301 10402 1335
rect 10282 1285 10402 1301
rect 10844 1409 10964 2505
rect 11029 4028 11030 4062
rect 11064 4046 11102 4062
rect 11064 4028 11066 4046
rect 11029 4012 11066 4028
rect 11100 4028 11102 4046
rect 11136 4046 11174 4062
rect 11136 4028 11138 4046
rect 11100 4012 11138 4028
rect 11172 4028 11174 4046
rect 11208 4028 11209 4062
rect 11172 4012 11209 4028
rect 11029 3988 11209 4012
rect 11029 3954 11030 3988
rect 11064 3978 11102 3988
rect 11064 3954 11066 3978
rect 11029 3944 11066 3954
rect 11100 3954 11102 3978
rect 11136 3978 11174 3988
rect 11136 3954 11138 3978
rect 11100 3944 11138 3954
rect 11172 3954 11174 3978
rect 11208 3954 11209 3988
rect 11172 3944 11209 3954
rect 11029 3914 11209 3944
rect 11029 3880 11030 3914
rect 11064 3910 11102 3914
rect 11064 3880 11066 3910
rect 11029 3876 11066 3880
rect 11100 3880 11102 3910
rect 11136 3910 11174 3914
rect 11136 3880 11138 3910
rect 11100 3876 11138 3880
rect 11172 3880 11174 3910
rect 11208 3880 11209 3914
rect 11172 3876 11209 3880
rect 11029 3842 11209 3876
rect 11029 3840 11066 3842
rect 11029 3806 11030 3840
rect 11064 3808 11066 3840
rect 11100 3840 11138 3842
rect 11100 3808 11102 3840
rect 11064 3806 11102 3808
rect 11136 3808 11138 3840
rect 11172 3840 11209 3842
rect 11172 3808 11174 3840
rect 11136 3806 11174 3808
rect 11208 3806 11209 3840
rect 11029 3774 11209 3806
rect 11029 3766 11066 3774
rect 11029 3732 11030 3766
rect 11064 3740 11066 3766
rect 11100 3766 11138 3774
rect 11100 3740 11102 3766
rect 11064 3732 11102 3740
rect 11136 3740 11138 3766
rect 11172 3766 11209 3774
rect 11172 3740 11174 3766
rect 11136 3732 11174 3740
rect 11208 3732 11209 3766
rect 11029 3706 11209 3732
rect 11029 3692 11066 3706
rect 11029 3658 11030 3692
rect 11064 3672 11066 3692
rect 11100 3692 11138 3706
rect 11100 3672 11102 3692
rect 11064 3658 11102 3672
rect 11136 3672 11138 3692
rect 11172 3692 11209 3706
rect 11172 3672 11174 3692
rect 11136 3658 11174 3672
rect 11208 3658 11209 3692
rect 11029 3638 11209 3658
rect 11029 3618 11066 3638
rect 11029 3584 11030 3618
rect 11064 3604 11066 3618
rect 11100 3618 11138 3638
rect 11100 3604 11102 3618
rect 11064 3584 11102 3604
rect 11136 3604 11138 3618
rect 11172 3618 11209 3638
rect 11172 3604 11174 3618
rect 11136 3584 11174 3604
rect 11208 3584 11209 3618
rect 11029 3570 11209 3584
rect 11029 3544 11066 3570
rect 11029 3510 11030 3544
rect 11064 3536 11066 3544
rect 11100 3544 11138 3570
rect 11100 3536 11102 3544
rect 11064 3510 11102 3536
rect 11136 3536 11138 3544
rect 11172 3544 11209 3570
rect 11172 3536 11174 3544
rect 11136 3510 11174 3536
rect 11208 3510 11209 3544
rect 11029 3502 11209 3510
rect 11029 3470 11066 3502
rect 11029 3436 11030 3470
rect 11064 3468 11066 3470
rect 11100 3470 11138 3502
rect 11100 3468 11102 3470
rect 11064 3436 11102 3468
rect 11136 3468 11138 3470
rect 11172 3470 11209 3502
rect 11172 3468 11174 3470
rect 11136 3436 11174 3468
rect 11208 3436 11209 3470
rect 11029 3434 11209 3436
rect 11029 3400 11066 3434
rect 11100 3400 11138 3434
rect 11172 3400 11209 3434
rect 11029 3396 11209 3400
rect 11029 3362 11030 3396
rect 11064 3366 11102 3396
rect 11064 3362 11066 3366
rect 11029 3332 11066 3362
rect 11100 3362 11102 3366
rect 11136 3366 11174 3396
rect 11136 3362 11138 3366
rect 11100 3332 11138 3362
rect 11172 3362 11174 3366
rect 11208 3362 11209 3396
rect 11172 3332 11209 3362
rect 11029 3322 11209 3332
rect 11029 3288 11030 3322
rect 11064 3298 11102 3322
rect 11064 3288 11066 3298
rect 11029 3264 11066 3288
rect 11100 3288 11102 3298
rect 11136 3298 11174 3322
rect 11136 3288 11138 3298
rect 11100 3264 11138 3288
rect 11172 3288 11174 3298
rect 11208 3288 11209 3322
rect 11172 3264 11209 3288
rect 11029 3248 11209 3264
rect 11029 3214 11030 3248
rect 11064 3230 11102 3248
rect 11064 3214 11066 3230
rect 11029 3196 11066 3214
rect 11100 3214 11102 3230
rect 11136 3230 11174 3248
rect 11136 3214 11138 3230
rect 11100 3196 11138 3214
rect 11172 3214 11174 3230
rect 11208 3214 11209 3248
rect 11172 3196 11209 3214
rect 11029 3174 11209 3196
rect 11029 3140 11030 3174
rect 11064 3162 11102 3174
rect 11064 3140 11066 3162
rect 11029 3128 11066 3140
rect 11100 3140 11102 3162
rect 11136 3162 11174 3174
rect 11136 3140 11138 3162
rect 11100 3128 11138 3140
rect 11172 3140 11174 3162
rect 11208 3140 11209 3174
rect 11172 3128 11209 3140
rect 11029 3100 11209 3128
rect 11029 3066 11030 3100
rect 11064 3066 11102 3100
rect 11136 3066 11174 3100
rect 11208 3066 11209 3100
rect 11029 3026 11209 3066
rect 11029 2992 11030 3026
rect 11064 2992 11102 3026
rect 11136 2992 11174 3026
rect 11208 2992 11209 3026
rect 11029 2952 11209 2992
rect 11029 2918 11030 2952
rect 11064 2918 11102 2952
rect 11136 2918 11174 2952
rect 11208 2918 11209 2952
rect 11029 2878 11209 2918
rect 11029 2844 11030 2878
rect 11064 2844 11102 2878
rect 11136 2844 11174 2878
rect 11208 2844 11209 2878
rect 11029 2804 11209 2844
rect 11029 2770 11030 2804
rect 11064 2770 11102 2804
rect 11136 2770 11174 2804
rect 11208 2770 11209 2804
rect 11029 2730 11209 2770
rect 11029 2696 11030 2730
rect 11064 2696 11102 2730
rect 11136 2696 11174 2730
rect 11208 2696 11209 2730
rect 11029 2656 11209 2696
rect 11029 2622 11030 2656
rect 11064 2622 11102 2656
rect 11136 2622 11174 2656
rect 11208 2622 11209 2656
rect 11029 2582 11209 2622
rect 11029 2548 11030 2582
rect 11064 2548 11102 2582
rect 11136 2548 11174 2582
rect 11208 2548 11209 2582
rect 11029 2508 11209 2548
rect 11029 2474 11030 2508
rect 11064 2474 11102 2508
rect 11136 2474 11174 2508
rect 11208 2474 11209 2508
rect 11029 2445 11209 2474
rect 11029 2434 11066 2445
rect 11029 2400 11030 2434
rect 11064 2411 11066 2434
rect 11100 2434 11138 2445
rect 11100 2411 11102 2434
rect 11064 2400 11102 2411
rect 11136 2411 11138 2434
rect 11172 2434 11209 2445
rect 11172 2411 11174 2434
rect 11136 2400 11174 2411
rect 11208 2400 11209 2434
rect 11029 2377 11209 2400
rect 11029 2360 11066 2377
rect 11029 2326 11030 2360
rect 11064 2343 11066 2360
rect 11100 2360 11138 2377
rect 11100 2343 11102 2360
rect 11064 2326 11102 2343
rect 11136 2343 11138 2360
rect 11172 2360 11209 2377
rect 11172 2343 11174 2360
rect 11136 2326 11174 2343
rect 11208 2326 11209 2360
rect 11029 2309 11209 2326
rect 11029 2286 11066 2309
rect 11029 2252 11030 2286
rect 11064 2275 11066 2286
rect 11100 2286 11138 2309
rect 11100 2275 11102 2286
rect 11064 2252 11102 2275
rect 11136 2275 11138 2286
rect 11172 2286 11209 2309
rect 11172 2275 11174 2286
rect 11136 2252 11174 2275
rect 11208 2252 11209 2286
rect 11029 2241 11209 2252
rect 11029 2212 11066 2241
rect 11029 2178 11030 2212
rect 11064 2207 11066 2212
rect 11100 2212 11138 2241
rect 11100 2207 11102 2212
rect 11064 2178 11102 2207
rect 11136 2207 11138 2212
rect 11172 2212 11209 2241
rect 11172 2207 11174 2212
rect 11136 2178 11174 2207
rect 11208 2178 11209 2212
rect 11029 2173 11209 2178
rect 11029 2139 11066 2173
rect 11100 2139 11138 2173
rect 11172 2139 11209 2173
rect 11029 2138 11209 2139
rect 11029 2104 11030 2138
rect 11064 2105 11102 2138
rect 11064 2104 11066 2105
rect 11029 2071 11066 2104
rect 11100 2104 11102 2105
rect 11136 2105 11174 2138
rect 11136 2104 11138 2105
rect 11100 2071 11138 2104
rect 11172 2104 11174 2105
rect 11208 2104 11209 2138
rect 11172 2071 11209 2104
rect 11029 2064 11209 2071
rect 11029 2030 11030 2064
rect 11064 2037 11102 2064
rect 11064 2030 11066 2037
rect 11029 2003 11066 2030
rect 11100 2030 11102 2037
rect 11136 2037 11174 2064
rect 11136 2030 11138 2037
rect 11100 2003 11138 2030
rect 11172 2030 11174 2037
rect 11208 2030 11209 2064
rect 11172 2003 11209 2030
rect 11029 1990 11209 2003
rect 11029 1956 11030 1990
rect 11064 1969 11102 1990
rect 11064 1956 11066 1969
rect 11029 1935 11066 1956
rect 11100 1956 11102 1969
rect 11136 1969 11174 1990
rect 11136 1956 11138 1969
rect 11100 1935 11138 1956
rect 11172 1956 11174 1969
rect 11208 1956 11209 1990
rect 11172 1935 11209 1956
rect 11029 1916 11209 1935
rect 11029 1882 11030 1916
rect 11064 1901 11102 1916
rect 11064 1882 11066 1901
rect 11029 1867 11066 1882
rect 11100 1882 11102 1901
rect 11136 1901 11174 1916
rect 11136 1882 11138 1901
rect 11100 1867 11138 1882
rect 11172 1882 11174 1901
rect 11208 1882 11209 1916
rect 11172 1867 11209 1882
rect 11029 1842 11209 1867
rect 11029 1808 11030 1842
rect 11064 1833 11102 1842
rect 11064 1808 11066 1833
rect 11029 1799 11066 1808
rect 11100 1808 11102 1833
rect 11136 1833 11174 1842
rect 11136 1808 11138 1833
rect 11100 1799 11138 1808
rect 11172 1808 11174 1833
rect 11208 1808 11209 1842
rect 11172 1799 11209 1808
rect 11029 1768 11209 1799
rect 11029 1734 11030 1768
rect 11064 1765 11102 1768
rect 11064 1734 11066 1765
rect 11029 1731 11066 1734
rect 11100 1734 11102 1765
rect 11136 1765 11174 1768
rect 11136 1734 11138 1765
rect 11100 1731 11138 1734
rect 11172 1734 11174 1765
rect 11208 1734 11209 1768
rect 11172 1731 11209 1734
rect 11029 1697 11209 1731
rect 11029 1694 11066 1697
rect 11029 1660 11030 1694
rect 11064 1663 11066 1694
rect 11100 1694 11138 1697
rect 11100 1663 11102 1694
rect 11064 1660 11102 1663
rect 11136 1663 11138 1694
rect 11172 1694 11209 1697
rect 11172 1663 11174 1694
rect 11136 1660 11174 1663
rect 11208 1660 11209 1694
rect 11029 1629 11209 1660
rect 11029 1620 11066 1629
rect 11029 1586 11030 1620
rect 11064 1595 11066 1620
rect 11100 1620 11138 1629
rect 11100 1595 11102 1620
rect 11064 1586 11102 1595
rect 11136 1595 11138 1620
rect 11172 1620 11209 1629
rect 11172 1595 11174 1620
rect 11136 1586 11174 1595
rect 11208 1586 11209 1620
rect 11029 1561 11209 1586
rect 11029 1545 11066 1561
rect 11029 1511 11030 1545
rect 11064 1527 11066 1545
rect 11100 1545 11138 1561
rect 11100 1527 11102 1545
rect 11064 1511 11102 1527
rect 11136 1527 11138 1545
rect 11172 1545 11209 1561
rect 11172 1527 11174 1545
rect 11136 1511 11174 1527
rect 11208 1511 11209 1545
rect 11274 3010 11394 4106
rect 11836 4388 11843 4494
rect 11949 4388 11956 4494
rect 11836 4214 11956 4388
rect 11836 4180 11879 4214
rect 11913 4180 11956 4214
rect 11836 4140 11956 4180
rect 11836 4106 11879 4140
rect 11913 4106 11956 4140
rect 11274 2976 11317 3010
rect 11351 2976 11394 3010
rect 11274 2932 11394 2976
rect 11274 2898 11317 2932
rect 11351 2898 11394 2932
rect 11274 2854 11394 2898
rect 11274 2820 11317 2854
rect 11351 2820 11394 2854
rect 11274 2776 11394 2820
rect 11274 2742 11317 2776
rect 11351 2742 11394 2776
rect 11274 2697 11394 2742
rect 11274 2663 11317 2697
rect 11351 2663 11394 2697
rect 11274 2618 11394 2663
rect 11274 2584 11317 2618
rect 11351 2584 11394 2618
rect 11274 2539 11394 2584
rect 11274 2505 11317 2539
rect 11351 2505 11394 2539
rect 11066 1491 11172 1511
rect 10844 1375 10887 1409
rect 10921 1375 10964 1409
rect 10844 1335 10964 1375
rect 10844 1301 10887 1335
rect 10921 1301 10964 1335
rect 10844 1285 10964 1301
rect 11274 1409 11394 2505
rect 11496 4050 11598 4062
rect 11632 4050 11734 4062
rect 11496 4046 11526 4050
rect 11704 4046 11734 4050
rect 11496 3978 11526 4012
rect 11704 3978 11734 4012
rect 11496 3910 11526 3944
rect 11704 3910 11734 3944
rect 11496 3842 11526 3876
rect 11704 3842 11734 3876
rect 11496 3774 11526 3808
rect 11704 3774 11734 3808
rect 11496 3706 11526 3740
rect 11704 3706 11734 3740
rect 11496 3638 11526 3672
rect 11704 3638 11734 3672
rect 11496 3570 11526 3604
rect 11704 3570 11734 3604
rect 11496 3502 11526 3536
rect 11704 3502 11734 3536
rect 11496 3434 11526 3468
rect 11704 3434 11734 3468
rect 11496 3366 11526 3400
rect 11704 3366 11734 3400
rect 11496 3298 11526 3332
rect 11704 3298 11734 3332
rect 11496 3230 11526 3264
rect 11704 3230 11734 3264
rect 11496 3162 11526 3196
rect 11704 3162 11734 3196
rect 11496 3080 11526 3128
rect 11560 3080 11670 3092
rect 11704 3080 11734 3128
rect 11496 3037 11734 3080
rect 11496 3003 11526 3037
rect 11560 3003 11598 3037
rect 11632 3003 11670 3037
rect 11704 3003 11734 3037
rect 11496 2954 11734 3003
rect 11496 2920 11526 2954
rect 11560 2935 11598 2954
rect 11632 2935 11670 2954
rect 11560 2920 11565 2935
rect 11632 2920 11633 2935
rect 11496 2901 11565 2920
rect 11599 2901 11633 2920
rect 11667 2920 11670 2935
rect 11704 2920 11734 2954
rect 11667 2901 11734 2920
rect 11496 2871 11734 2901
rect 11496 2837 11526 2871
rect 11560 2855 11598 2871
rect 11632 2855 11670 2871
rect 11560 2837 11565 2855
rect 11632 2837 11633 2855
rect 11496 2821 11565 2837
rect 11599 2821 11633 2837
rect 11667 2837 11670 2855
rect 11704 2837 11734 2871
rect 11667 2821 11734 2837
rect 11496 2787 11734 2821
rect 11496 2753 11526 2787
rect 11560 2775 11598 2787
rect 11632 2775 11670 2787
rect 11560 2753 11565 2775
rect 11632 2753 11633 2775
rect 11496 2741 11565 2753
rect 11599 2741 11633 2753
rect 11667 2753 11670 2775
rect 11704 2753 11734 2787
rect 11667 2741 11734 2753
rect 11496 2703 11734 2741
rect 11496 2669 11526 2703
rect 11560 2695 11598 2703
rect 11632 2695 11670 2703
rect 11560 2669 11565 2695
rect 11632 2669 11633 2695
rect 11496 2661 11565 2669
rect 11599 2661 11633 2669
rect 11667 2669 11670 2695
rect 11704 2669 11734 2703
rect 11667 2661 11734 2669
rect 11496 2619 11734 2661
rect 11496 2585 11526 2619
rect 11560 2614 11598 2619
rect 11632 2614 11670 2619
rect 11560 2585 11565 2614
rect 11632 2585 11633 2614
rect 11496 2580 11565 2585
rect 11599 2580 11633 2585
rect 11667 2585 11670 2614
rect 11704 2585 11734 2619
rect 11667 2580 11734 2585
rect 11496 2535 11734 2580
rect 11496 2501 11526 2535
rect 11560 2501 11598 2535
rect 11632 2501 11670 2535
rect 11704 2501 11734 2535
rect 11496 2461 11734 2501
rect 11496 2449 11598 2461
rect 11632 2449 11734 2461
rect 11496 2445 11526 2449
rect 11704 2445 11734 2449
rect 11496 2377 11526 2411
rect 11704 2377 11734 2411
rect 11496 2309 11526 2343
rect 11704 2309 11734 2343
rect 11496 2241 11526 2275
rect 11704 2241 11734 2275
rect 11496 2173 11526 2207
rect 11704 2173 11734 2207
rect 11496 2105 11526 2139
rect 11704 2105 11734 2139
rect 11496 2037 11526 2071
rect 11704 2037 11734 2071
rect 11496 1969 11526 2003
rect 11704 1969 11734 2003
rect 11496 1901 11526 1935
rect 11704 1901 11734 1935
rect 11496 1833 11526 1867
rect 11704 1833 11734 1867
rect 11496 1765 11526 1799
rect 11704 1765 11734 1799
rect 11496 1697 11526 1731
rect 11704 1697 11734 1731
rect 11496 1629 11526 1663
rect 11704 1629 11734 1663
rect 11496 1561 11526 1595
rect 11704 1561 11734 1595
rect 11496 1479 11526 1527
rect 11560 1479 11670 1491
rect 11704 1479 11734 1527
rect 11496 1464 11734 1479
rect 11836 3010 11956 4106
rect 12266 4388 12273 4494
rect 12379 4388 12386 4494
rect 12266 4214 12386 4388
rect 12266 4180 12309 4214
rect 12343 4180 12386 4214
rect 12266 4140 12386 4180
rect 12266 4106 12309 4140
rect 12343 4106 12386 4140
rect 11836 2976 11879 3010
rect 11913 2976 11956 3010
rect 11836 2932 11956 2976
rect 11836 2898 11879 2932
rect 11913 2898 11956 2932
rect 11836 2854 11956 2898
rect 11836 2820 11879 2854
rect 11913 2820 11956 2854
rect 11836 2776 11956 2820
rect 11836 2742 11879 2776
rect 11913 2742 11956 2776
rect 11836 2697 11956 2742
rect 11836 2663 11879 2697
rect 11913 2663 11956 2697
rect 11836 2618 11956 2663
rect 11836 2584 11879 2618
rect 11913 2584 11956 2618
rect 11836 2539 11956 2584
rect 11836 2505 11879 2539
rect 11913 2505 11956 2539
rect 11274 1375 11317 1409
rect 11351 1375 11394 1409
rect 11274 1335 11394 1375
rect 11274 1301 11317 1335
rect 11351 1301 11394 1335
rect 11274 1285 11394 1301
rect 11836 1409 11956 2505
rect 12021 4028 12022 4062
rect 12056 4046 12094 4062
rect 12056 4028 12058 4046
rect 12021 4012 12058 4028
rect 12092 4028 12094 4046
rect 12128 4046 12166 4062
rect 12128 4028 12130 4046
rect 12092 4012 12130 4028
rect 12164 4028 12166 4046
rect 12200 4028 12201 4062
rect 12164 4012 12201 4028
rect 12021 3988 12201 4012
rect 12021 3954 12022 3988
rect 12056 3978 12094 3988
rect 12056 3954 12058 3978
rect 12021 3944 12058 3954
rect 12092 3954 12094 3978
rect 12128 3978 12166 3988
rect 12128 3954 12130 3978
rect 12092 3944 12130 3954
rect 12164 3954 12166 3978
rect 12200 3954 12201 3988
rect 12164 3944 12201 3954
rect 12021 3914 12201 3944
rect 12021 3880 12022 3914
rect 12056 3910 12094 3914
rect 12056 3880 12058 3910
rect 12021 3876 12058 3880
rect 12092 3880 12094 3910
rect 12128 3910 12166 3914
rect 12128 3880 12130 3910
rect 12092 3876 12130 3880
rect 12164 3880 12166 3910
rect 12200 3880 12201 3914
rect 12164 3876 12201 3880
rect 12021 3842 12201 3876
rect 12021 3840 12058 3842
rect 12021 3806 12022 3840
rect 12056 3808 12058 3840
rect 12092 3840 12130 3842
rect 12092 3808 12094 3840
rect 12056 3806 12094 3808
rect 12128 3808 12130 3840
rect 12164 3840 12201 3842
rect 12164 3808 12166 3840
rect 12128 3806 12166 3808
rect 12200 3806 12201 3840
rect 12021 3774 12201 3806
rect 12021 3766 12058 3774
rect 12021 3732 12022 3766
rect 12056 3740 12058 3766
rect 12092 3766 12130 3774
rect 12092 3740 12094 3766
rect 12056 3732 12094 3740
rect 12128 3740 12130 3766
rect 12164 3766 12201 3774
rect 12164 3740 12166 3766
rect 12128 3732 12166 3740
rect 12200 3732 12201 3766
rect 12021 3706 12201 3732
rect 12021 3692 12058 3706
rect 12021 3658 12022 3692
rect 12056 3672 12058 3692
rect 12092 3692 12130 3706
rect 12092 3672 12094 3692
rect 12056 3658 12094 3672
rect 12128 3672 12130 3692
rect 12164 3692 12201 3706
rect 12164 3672 12166 3692
rect 12128 3658 12166 3672
rect 12200 3658 12201 3692
rect 12021 3638 12201 3658
rect 12021 3618 12058 3638
rect 12021 3584 12022 3618
rect 12056 3604 12058 3618
rect 12092 3618 12130 3638
rect 12092 3604 12094 3618
rect 12056 3584 12094 3604
rect 12128 3604 12130 3618
rect 12164 3618 12201 3638
rect 12164 3604 12166 3618
rect 12128 3584 12166 3604
rect 12200 3584 12201 3618
rect 12021 3570 12201 3584
rect 12021 3544 12058 3570
rect 12021 3510 12022 3544
rect 12056 3536 12058 3544
rect 12092 3544 12130 3570
rect 12092 3536 12094 3544
rect 12056 3510 12094 3536
rect 12128 3536 12130 3544
rect 12164 3544 12201 3570
rect 12164 3536 12166 3544
rect 12128 3510 12166 3536
rect 12200 3510 12201 3544
rect 12021 3502 12201 3510
rect 12021 3470 12058 3502
rect 12021 3436 12022 3470
rect 12056 3468 12058 3470
rect 12092 3470 12130 3502
rect 12092 3468 12094 3470
rect 12056 3436 12094 3468
rect 12128 3468 12130 3470
rect 12164 3470 12201 3502
rect 12164 3468 12166 3470
rect 12128 3436 12166 3468
rect 12200 3436 12201 3470
rect 12021 3434 12201 3436
rect 12021 3400 12058 3434
rect 12092 3400 12130 3434
rect 12164 3400 12201 3434
rect 12021 3396 12201 3400
rect 12021 3362 12022 3396
rect 12056 3366 12094 3396
rect 12056 3362 12058 3366
rect 12021 3332 12058 3362
rect 12092 3362 12094 3366
rect 12128 3366 12166 3396
rect 12128 3362 12130 3366
rect 12092 3332 12130 3362
rect 12164 3362 12166 3366
rect 12200 3362 12201 3396
rect 12164 3332 12201 3362
rect 12021 3322 12201 3332
rect 12021 3288 12022 3322
rect 12056 3298 12094 3322
rect 12056 3288 12058 3298
rect 12021 3264 12058 3288
rect 12092 3288 12094 3298
rect 12128 3298 12166 3322
rect 12128 3288 12130 3298
rect 12092 3264 12130 3288
rect 12164 3288 12166 3298
rect 12200 3288 12201 3322
rect 12164 3264 12201 3288
rect 12021 3248 12201 3264
rect 12021 3214 12022 3248
rect 12056 3230 12094 3248
rect 12056 3214 12058 3230
rect 12021 3196 12058 3214
rect 12092 3214 12094 3230
rect 12128 3230 12166 3248
rect 12128 3214 12130 3230
rect 12092 3196 12130 3214
rect 12164 3214 12166 3230
rect 12200 3214 12201 3248
rect 12164 3196 12201 3214
rect 12021 3174 12201 3196
rect 12021 3140 12022 3174
rect 12056 3162 12094 3174
rect 12056 3140 12058 3162
rect 12021 3128 12058 3140
rect 12092 3140 12094 3162
rect 12128 3162 12166 3174
rect 12128 3140 12130 3162
rect 12092 3128 12130 3140
rect 12164 3140 12166 3162
rect 12200 3140 12201 3174
rect 12164 3128 12201 3140
rect 12021 3100 12201 3128
rect 12021 3066 12022 3100
rect 12056 3066 12094 3100
rect 12128 3066 12166 3100
rect 12200 3066 12201 3100
rect 12021 3026 12201 3066
rect 12021 2992 12022 3026
rect 12056 2992 12094 3026
rect 12128 2992 12166 3026
rect 12200 2992 12201 3026
rect 12021 2952 12201 2992
rect 12021 2918 12022 2952
rect 12056 2918 12094 2952
rect 12128 2918 12166 2952
rect 12200 2918 12201 2952
rect 12021 2878 12201 2918
rect 12021 2844 12022 2878
rect 12056 2844 12094 2878
rect 12128 2844 12166 2878
rect 12200 2844 12201 2878
rect 12021 2804 12201 2844
rect 12021 2770 12022 2804
rect 12056 2770 12094 2804
rect 12128 2770 12166 2804
rect 12200 2770 12201 2804
rect 12021 2730 12201 2770
rect 12021 2696 12022 2730
rect 12056 2696 12094 2730
rect 12128 2696 12166 2730
rect 12200 2696 12201 2730
rect 12021 2656 12201 2696
rect 12021 2622 12022 2656
rect 12056 2622 12094 2656
rect 12128 2622 12166 2656
rect 12200 2622 12201 2656
rect 12021 2582 12201 2622
rect 12021 2548 12022 2582
rect 12056 2548 12094 2582
rect 12128 2548 12166 2582
rect 12200 2548 12201 2582
rect 12021 2508 12201 2548
rect 12021 2474 12022 2508
rect 12056 2474 12094 2508
rect 12128 2474 12166 2508
rect 12200 2474 12201 2508
rect 12021 2445 12201 2474
rect 12021 2434 12058 2445
rect 12021 2400 12022 2434
rect 12056 2411 12058 2434
rect 12092 2434 12130 2445
rect 12092 2411 12094 2434
rect 12056 2400 12094 2411
rect 12128 2411 12130 2434
rect 12164 2434 12201 2445
rect 12164 2411 12166 2434
rect 12128 2400 12166 2411
rect 12200 2400 12201 2434
rect 12021 2377 12201 2400
rect 12021 2360 12058 2377
rect 12021 2326 12022 2360
rect 12056 2343 12058 2360
rect 12092 2360 12130 2377
rect 12092 2343 12094 2360
rect 12056 2326 12094 2343
rect 12128 2343 12130 2360
rect 12164 2360 12201 2377
rect 12164 2343 12166 2360
rect 12128 2326 12166 2343
rect 12200 2326 12201 2360
rect 12021 2309 12201 2326
rect 12021 2286 12058 2309
rect 12021 2252 12022 2286
rect 12056 2275 12058 2286
rect 12092 2286 12130 2309
rect 12092 2275 12094 2286
rect 12056 2252 12094 2275
rect 12128 2275 12130 2286
rect 12164 2286 12201 2309
rect 12164 2275 12166 2286
rect 12128 2252 12166 2275
rect 12200 2252 12201 2286
rect 12021 2241 12201 2252
rect 12021 2212 12058 2241
rect 12021 2178 12022 2212
rect 12056 2207 12058 2212
rect 12092 2212 12130 2241
rect 12092 2207 12094 2212
rect 12056 2178 12094 2207
rect 12128 2207 12130 2212
rect 12164 2212 12201 2241
rect 12164 2207 12166 2212
rect 12128 2178 12166 2207
rect 12200 2178 12201 2212
rect 12021 2173 12201 2178
rect 12021 2139 12058 2173
rect 12092 2139 12130 2173
rect 12164 2139 12201 2173
rect 12021 2138 12201 2139
rect 12021 2104 12022 2138
rect 12056 2105 12094 2138
rect 12056 2104 12058 2105
rect 12021 2071 12058 2104
rect 12092 2104 12094 2105
rect 12128 2105 12166 2138
rect 12128 2104 12130 2105
rect 12092 2071 12130 2104
rect 12164 2104 12166 2105
rect 12200 2104 12201 2138
rect 12164 2071 12201 2104
rect 12021 2064 12201 2071
rect 12021 2030 12022 2064
rect 12056 2037 12094 2064
rect 12056 2030 12058 2037
rect 12021 2003 12058 2030
rect 12092 2030 12094 2037
rect 12128 2037 12166 2064
rect 12128 2030 12130 2037
rect 12092 2003 12130 2030
rect 12164 2030 12166 2037
rect 12200 2030 12201 2064
rect 12164 2003 12201 2030
rect 12021 1990 12201 2003
rect 12021 1956 12022 1990
rect 12056 1969 12094 1990
rect 12056 1956 12058 1969
rect 12021 1935 12058 1956
rect 12092 1956 12094 1969
rect 12128 1969 12166 1990
rect 12128 1956 12130 1969
rect 12092 1935 12130 1956
rect 12164 1956 12166 1969
rect 12200 1956 12201 1990
rect 12164 1935 12201 1956
rect 12021 1916 12201 1935
rect 12021 1882 12022 1916
rect 12056 1901 12094 1916
rect 12056 1882 12058 1901
rect 12021 1867 12058 1882
rect 12092 1882 12094 1901
rect 12128 1901 12166 1916
rect 12128 1882 12130 1901
rect 12092 1867 12130 1882
rect 12164 1882 12166 1901
rect 12200 1882 12201 1916
rect 12164 1867 12201 1882
rect 12021 1842 12201 1867
rect 12021 1808 12022 1842
rect 12056 1833 12094 1842
rect 12056 1808 12058 1833
rect 12021 1799 12058 1808
rect 12092 1808 12094 1833
rect 12128 1833 12166 1842
rect 12128 1808 12130 1833
rect 12092 1799 12130 1808
rect 12164 1808 12166 1833
rect 12200 1808 12201 1842
rect 12164 1799 12201 1808
rect 12021 1768 12201 1799
rect 12021 1734 12022 1768
rect 12056 1765 12094 1768
rect 12056 1734 12058 1765
rect 12021 1731 12058 1734
rect 12092 1734 12094 1765
rect 12128 1765 12166 1768
rect 12128 1734 12130 1765
rect 12092 1731 12130 1734
rect 12164 1734 12166 1765
rect 12200 1734 12201 1768
rect 12164 1731 12201 1734
rect 12021 1697 12201 1731
rect 12021 1694 12058 1697
rect 12021 1660 12022 1694
rect 12056 1663 12058 1694
rect 12092 1694 12130 1697
rect 12092 1663 12094 1694
rect 12056 1660 12094 1663
rect 12128 1663 12130 1694
rect 12164 1694 12201 1697
rect 12164 1663 12166 1694
rect 12128 1660 12166 1663
rect 12200 1660 12201 1694
rect 12021 1629 12201 1660
rect 12021 1620 12058 1629
rect 12021 1586 12022 1620
rect 12056 1595 12058 1620
rect 12092 1620 12130 1629
rect 12092 1595 12094 1620
rect 12056 1586 12094 1595
rect 12128 1595 12130 1620
rect 12164 1620 12201 1629
rect 12164 1595 12166 1620
rect 12128 1586 12166 1595
rect 12200 1586 12201 1620
rect 12021 1561 12201 1586
rect 12021 1545 12058 1561
rect 12021 1511 12022 1545
rect 12056 1527 12058 1545
rect 12092 1545 12130 1561
rect 12092 1527 12094 1545
rect 12056 1511 12094 1527
rect 12128 1527 12130 1545
rect 12164 1545 12201 1561
rect 12164 1527 12166 1545
rect 12128 1511 12166 1527
rect 12200 1511 12201 1545
rect 12266 3010 12386 4106
rect 12828 4388 12835 4494
rect 12941 4388 12948 4494
rect 12828 4214 12948 4388
rect 12828 4180 12871 4214
rect 12905 4180 12948 4214
rect 12828 4140 12948 4180
rect 12828 4106 12871 4140
rect 12905 4106 12948 4140
rect 12266 2976 12309 3010
rect 12343 2976 12386 3010
rect 12266 2932 12386 2976
rect 12266 2898 12309 2932
rect 12343 2898 12386 2932
rect 12266 2854 12386 2898
rect 12266 2820 12309 2854
rect 12343 2820 12386 2854
rect 12266 2776 12386 2820
rect 12266 2742 12309 2776
rect 12343 2742 12386 2776
rect 12266 2697 12386 2742
rect 12266 2663 12309 2697
rect 12343 2663 12386 2697
rect 12266 2618 12386 2663
rect 12266 2584 12309 2618
rect 12343 2584 12386 2618
rect 12266 2539 12386 2584
rect 12266 2505 12309 2539
rect 12343 2505 12386 2539
rect 12058 1491 12164 1511
rect 11836 1375 11879 1409
rect 11913 1375 11956 1409
rect 11836 1335 11956 1375
rect 11836 1301 11879 1335
rect 11913 1301 11956 1335
rect 11836 1285 11956 1301
rect 12266 1409 12386 2505
rect 12488 4050 12590 4062
rect 12624 4050 12726 4062
rect 12488 4046 12518 4050
rect 12696 4046 12726 4050
rect 12488 3978 12518 4012
rect 12696 3978 12726 4012
rect 12488 3910 12518 3944
rect 12696 3910 12726 3944
rect 12488 3842 12518 3876
rect 12696 3842 12726 3876
rect 12488 3774 12518 3808
rect 12696 3774 12726 3808
rect 12488 3706 12518 3740
rect 12696 3706 12726 3740
rect 12488 3638 12518 3672
rect 12696 3638 12726 3672
rect 12488 3570 12518 3604
rect 12696 3570 12726 3604
rect 12488 3502 12518 3536
rect 12696 3502 12726 3536
rect 12488 3434 12518 3468
rect 12696 3434 12726 3468
rect 12488 3366 12518 3400
rect 12696 3366 12726 3400
rect 12488 3298 12518 3332
rect 12696 3298 12726 3332
rect 12488 3230 12518 3264
rect 12696 3230 12726 3264
rect 12488 3162 12518 3196
rect 12696 3162 12726 3196
rect 12488 3080 12518 3128
rect 12552 3080 12662 3092
rect 12696 3080 12726 3128
rect 12488 3038 12726 3080
rect 12488 3004 12518 3038
rect 12552 3004 12590 3038
rect 12624 3004 12662 3038
rect 12696 3004 12726 3038
rect 12488 2955 12726 3004
rect 12488 2921 12518 2955
rect 12552 2935 12590 2955
rect 12624 2935 12662 2955
rect 12552 2921 12557 2935
rect 12624 2921 12625 2935
rect 12488 2901 12557 2921
rect 12591 2901 12625 2921
rect 12659 2921 12662 2935
rect 12696 2921 12726 2955
rect 12659 2901 12726 2921
rect 12488 2871 12726 2901
rect 12488 2837 12518 2871
rect 12552 2855 12590 2871
rect 12624 2855 12662 2871
rect 12552 2837 12557 2855
rect 12624 2837 12625 2855
rect 12488 2821 12557 2837
rect 12591 2821 12625 2837
rect 12659 2837 12662 2855
rect 12696 2837 12726 2871
rect 12659 2821 12726 2837
rect 12488 2787 12726 2821
rect 12488 2753 12518 2787
rect 12552 2775 12590 2787
rect 12624 2775 12662 2787
rect 12552 2753 12557 2775
rect 12624 2753 12625 2775
rect 12488 2741 12557 2753
rect 12591 2741 12625 2753
rect 12659 2753 12662 2775
rect 12696 2753 12726 2787
rect 12659 2741 12726 2753
rect 12488 2703 12726 2741
rect 12488 2669 12518 2703
rect 12552 2695 12590 2703
rect 12624 2695 12662 2703
rect 12552 2669 12557 2695
rect 12624 2669 12625 2695
rect 12488 2661 12557 2669
rect 12591 2661 12625 2669
rect 12659 2669 12662 2695
rect 12696 2669 12726 2703
rect 12659 2661 12726 2669
rect 12488 2619 12726 2661
rect 12488 2585 12518 2619
rect 12552 2614 12590 2619
rect 12624 2614 12662 2619
rect 12552 2585 12557 2614
rect 12624 2585 12625 2614
rect 12488 2580 12557 2585
rect 12591 2580 12625 2585
rect 12659 2585 12662 2614
rect 12696 2585 12726 2619
rect 12659 2580 12726 2585
rect 12488 2535 12726 2580
rect 12488 2501 12518 2535
rect 12552 2501 12590 2535
rect 12624 2501 12662 2535
rect 12696 2501 12726 2535
rect 12488 2461 12726 2501
rect 12488 2449 12590 2461
rect 12624 2449 12726 2461
rect 12488 2445 12518 2449
rect 12696 2445 12726 2449
rect 12488 2377 12518 2411
rect 12696 2377 12726 2411
rect 12488 2309 12518 2343
rect 12696 2309 12726 2343
rect 12488 2241 12518 2275
rect 12696 2241 12726 2275
rect 12488 2173 12518 2207
rect 12696 2173 12726 2207
rect 12488 2105 12518 2139
rect 12696 2105 12726 2139
rect 12488 2037 12518 2071
rect 12696 2037 12726 2071
rect 12488 1969 12518 2003
rect 12696 1969 12726 2003
rect 12488 1901 12518 1935
rect 12696 1901 12726 1935
rect 12488 1833 12518 1867
rect 12696 1833 12726 1867
rect 12488 1765 12518 1799
rect 12696 1765 12726 1799
rect 12488 1697 12518 1731
rect 12696 1697 12726 1731
rect 12488 1629 12518 1663
rect 12696 1629 12726 1663
rect 12488 1561 12518 1595
rect 12696 1561 12726 1595
rect 12488 1479 12518 1527
rect 12552 1479 12662 1491
rect 12696 1479 12726 1527
rect 12488 1464 12726 1479
rect 12828 3010 12948 4106
rect 13258 4388 13265 4494
rect 13371 4388 13378 4494
rect 13258 4214 13378 4388
rect 13258 4180 13301 4214
rect 13335 4180 13378 4214
rect 13258 4140 13378 4180
rect 13258 4106 13301 4140
rect 13335 4106 13378 4140
rect 12828 2976 12871 3010
rect 12905 2976 12948 3010
rect 12828 2932 12948 2976
rect 12828 2898 12871 2932
rect 12905 2898 12948 2932
rect 12828 2854 12948 2898
rect 12828 2820 12871 2854
rect 12905 2820 12948 2854
rect 12828 2776 12948 2820
rect 12828 2742 12871 2776
rect 12905 2742 12948 2776
rect 12828 2697 12948 2742
rect 12828 2663 12871 2697
rect 12905 2663 12948 2697
rect 12828 2618 12948 2663
rect 12828 2584 12871 2618
rect 12905 2584 12948 2618
rect 12828 2539 12948 2584
rect 12828 2505 12871 2539
rect 12905 2505 12948 2539
rect 12266 1375 12309 1409
rect 12343 1375 12386 1409
rect 12266 1335 12386 1375
rect 12266 1301 12309 1335
rect 12343 1301 12386 1335
rect 12266 1285 12386 1301
rect 12828 1409 12948 2505
rect 13013 4028 13014 4062
rect 13048 4046 13086 4062
rect 13048 4028 13050 4046
rect 13013 4012 13050 4028
rect 13084 4028 13086 4046
rect 13120 4046 13158 4062
rect 13120 4028 13122 4046
rect 13084 4012 13122 4028
rect 13156 4028 13158 4046
rect 13192 4028 13193 4062
rect 13156 4012 13193 4028
rect 13013 3988 13193 4012
rect 13013 3954 13014 3988
rect 13048 3978 13086 3988
rect 13048 3954 13050 3978
rect 13013 3944 13050 3954
rect 13084 3954 13086 3978
rect 13120 3978 13158 3988
rect 13120 3954 13122 3978
rect 13084 3944 13122 3954
rect 13156 3954 13158 3978
rect 13192 3954 13193 3988
rect 13156 3944 13193 3954
rect 13013 3914 13193 3944
rect 13013 3880 13014 3914
rect 13048 3910 13086 3914
rect 13048 3880 13050 3910
rect 13013 3876 13050 3880
rect 13084 3880 13086 3910
rect 13120 3910 13158 3914
rect 13120 3880 13122 3910
rect 13084 3876 13122 3880
rect 13156 3880 13158 3910
rect 13192 3880 13193 3914
rect 13156 3876 13193 3880
rect 13013 3842 13193 3876
rect 13013 3840 13050 3842
rect 13013 3806 13014 3840
rect 13048 3808 13050 3840
rect 13084 3840 13122 3842
rect 13084 3808 13086 3840
rect 13048 3806 13086 3808
rect 13120 3808 13122 3840
rect 13156 3840 13193 3842
rect 13156 3808 13158 3840
rect 13120 3806 13158 3808
rect 13192 3806 13193 3840
rect 13013 3774 13193 3806
rect 13013 3766 13050 3774
rect 13013 3732 13014 3766
rect 13048 3740 13050 3766
rect 13084 3766 13122 3774
rect 13084 3740 13086 3766
rect 13048 3732 13086 3740
rect 13120 3740 13122 3766
rect 13156 3766 13193 3774
rect 13156 3740 13158 3766
rect 13120 3732 13158 3740
rect 13192 3732 13193 3766
rect 13013 3706 13193 3732
rect 13013 3692 13050 3706
rect 13013 3658 13014 3692
rect 13048 3672 13050 3692
rect 13084 3692 13122 3706
rect 13084 3672 13086 3692
rect 13048 3658 13086 3672
rect 13120 3672 13122 3692
rect 13156 3692 13193 3706
rect 13156 3672 13158 3692
rect 13120 3658 13158 3672
rect 13192 3658 13193 3692
rect 13013 3638 13193 3658
rect 13013 3618 13050 3638
rect 13013 3584 13014 3618
rect 13048 3604 13050 3618
rect 13084 3618 13122 3638
rect 13084 3604 13086 3618
rect 13048 3584 13086 3604
rect 13120 3604 13122 3618
rect 13156 3618 13193 3638
rect 13156 3604 13158 3618
rect 13120 3584 13158 3604
rect 13192 3584 13193 3618
rect 13013 3570 13193 3584
rect 13013 3544 13050 3570
rect 13013 3510 13014 3544
rect 13048 3536 13050 3544
rect 13084 3544 13122 3570
rect 13084 3536 13086 3544
rect 13048 3510 13086 3536
rect 13120 3536 13122 3544
rect 13156 3544 13193 3570
rect 13156 3536 13158 3544
rect 13120 3510 13158 3536
rect 13192 3510 13193 3544
rect 13013 3502 13193 3510
rect 13013 3470 13050 3502
rect 13013 3436 13014 3470
rect 13048 3468 13050 3470
rect 13084 3470 13122 3502
rect 13084 3468 13086 3470
rect 13048 3436 13086 3468
rect 13120 3468 13122 3470
rect 13156 3470 13193 3502
rect 13156 3468 13158 3470
rect 13120 3436 13158 3468
rect 13192 3436 13193 3470
rect 13013 3434 13193 3436
rect 13013 3400 13050 3434
rect 13084 3400 13122 3434
rect 13156 3400 13193 3434
rect 13013 3396 13193 3400
rect 13013 3362 13014 3396
rect 13048 3366 13086 3396
rect 13048 3362 13050 3366
rect 13013 3332 13050 3362
rect 13084 3362 13086 3366
rect 13120 3366 13158 3396
rect 13120 3362 13122 3366
rect 13084 3332 13122 3362
rect 13156 3362 13158 3366
rect 13192 3362 13193 3396
rect 13156 3332 13193 3362
rect 13013 3322 13193 3332
rect 13013 3288 13014 3322
rect 13048 3298 13086 3322
rect 13048 3288 13050 3298
rect 13013 3264 13050 3288
rect 13084 3288 13086 3298
rect 13120 3298 13158 3322
rect 13120 3288 13122 3298
rect 13084 3264 13122 3288
rect 13156 3288 13158 3298
rect 13192 3288 13193 3322
rect 13156 3264 13193 3288
rect 13013 3248 13193 3264
rect 13013 3214 13014 3248
rect 13048 3230 13086 3248
rect 13048 3214 13050 3230
rect 13013 3196 13050 3214
rect 13084 3214 13086 3230
rect 13120 3230 13158 3248
rect 13120 3214 13122 3230
rect 13084 3196 13122 3214
rect 13156 3214 13158 3230
rect 13192 3214 13193 3248
rect 13156 3196 13193 3214
rect 13013 3174 13193 3196
rect 13013 3140 13014 3174
rect 13048 3162 13086 3174
rect 13048 3140 13050 3162
rect 13013 3128 13050 3140
rect 13084 3140 13086 3162
rect 13120 3162 13158 3174
rect 13120 3140 13122 3162
rect 13084 3128 13122 3140
rect 13156 3140 13158 3162
rect 13192 3140 13193 3174
rect 13156 3128 13193 3140
rect 13013 3100 13193 3128
rect 13013 3066 13014 3100
rect 13048 3066 13086 3100
rect 13120 3066 13158 3100
rect 13192 3066 13193 3100
rect 13013 3026 13193 3066
rect 13013 2992 13014 3026
rect 13048 2992 13086 3026
rect 13120 2992 13158 3026
rect 13192 2992 13193 3026
rect 13013 2952 13193 2992
rect 13013 2918 13014 2952
rect 13048 2918 13086 2952
rect 13120 2918 13158 2952
rect 13192 2918 13193 2952
rect 13013 2878 13193 2918
rect 13013 2844 13014 2878
rect 13048 2844 13086 2878
rect 13120 2844 13158 2878
rect 13192 2844 13193 2878
rect 13013 2804 13193 2844
rect 13013 2770 13014 2804
rect 13048 2770 13086 2804
rect 13120 2770 13158 2804
rect 13192 2770 13193 2804
rect 13013 2730 13193 2770
rect 13013 2696 13014 2730
rect 13048 2696 13086 2730
rect 13120 2696 13158 2730
rect 13192 2696 13193 2730
rect 13013 2656 13193 2696
rect 13013 2622 13014 2656
rect 13048 2622 13086 2656
rect 13120 2622 13158 2656
rect 13192 2622 13193 2656
rect 13013 2582 13193 2622
rect 13013 2548 13014 2582
rect 13048 2548 13086 2582
rect 13120 2548 13158 2582
rect 13192 2548 13193 2582
rect 13013 2508 13193 2548
rect 13013 2474 13014 2508
rect 13048 2474 13086 2508
rect 13120 2474 13158 2508
rect 13192 2474 13193 2508
rect 13013 2445 13193 2474
rect 13013 2434 13050 2445
rect 13013 2400 13014 2434
rect 13048 2411 13050 2434
rect 13084 2434 13122 2445
rect 13084 2411 13086 2434
rect 13048 2400 13086 2411
rect 13120 2411 13122 2434
rect 13156 2434 13193 2445
rect 13156 2411 13158 2434
rect 13120 2400 13158 2411
rect 13192 2400 13193 2434
rect 13013 2377 13193 2400
rect 13013 2360 13050 2377
rect 13013 2326 13014 2360
rect 13048 2343 13050 2360
rect 13084 2360 13122 2377
rect 13084 2343 13086 2360
rect 13048 2326 13086 2343
rect 13120 2343 13122 2360
rect 13156 2360 13193 2377
rect 13156 2343 13158 2360
rect 13120 2326 13158 2343
rect 13192 2326 13193 2360
rect 13013 2309 13193 2326
rect 13013 2286 13050 2309
rect 13013 2252 13014 2286
rect 13048 2275 13050 2286
rect 13084 2286 13122 2309
rect 13084 2275 13086 2286
rect 13048 2252 13086 2275
rect 13120 2275 13122 2286
rect 13156 2286 13193 2309
rect 13156 2275 13158 2286
rect 13120 2252 13158 2275
rect 13192 2252 13193 2286
rect 13013 2241 13193 2252
rect 13013 2212 13050 2241
rect 13013 2178 13014 2212
rect 13048 2207 13050 2212
rect 13084 2212 13122 2241
rect 13084 2207 13086 2212
rect 13048 2178 13086 2207
rect 13120 2207 13122 2212
rect 13156 2212 13193 2241
rect 13156 2207 13158 2212
rect 13120 2178 13158 2207
rect 13192 2178 13193 2212
rect 13013 2173 13193 2178
rect 13013 2139 13050 2173
rect 13084 2139 13122 2173
rect 13156 2139 13193 2173
rect 13013 2138 13193 2139
rect 13013 2104 13014 2138
rect 13048 2105 13086 2138
rect 13048 2104 13050 2105
rect 13013 2071 13050 2104
rect 13084 2104 13086 2105
rect 13120 2105 13158 2138
rect 13120 2104 13122 2105
rect 13084 2071 13122 2104
rect 13156 2104 13158 2105
rect 13192 2104 13193 2138
rect 13156 2071 13193 2104
rect 13013 2064 13193 2071
rect 13013 2030 13014 2064
rect 13048 2037 13086 2064
rect 13048 2030 13050 2037
rect 13013 2003 13050 2030
rect 13084 2030 13086 2037
rect 13120 2037 13158 2064
rect 13120 2030 13122 2037
rect 13084 2003 13122 2030
rect 13156 2030 13158 2037
rect 13192 2030 13193 2064
rect 13156 2003 13193 2030
rect 13013 1990 13193 2003
rect 13013 1956 13014 1990
rect 13048 1969 13086 1990
rect 13048 1956 13050 1969
rect 13013 1935 13050 1956
rect 13084 1956 13086 1969
rect 13120 1969 13158 1990
rect 13120 1956 13122 1969
rect 13084 1935 13122 1956
rect 13156 1956 13158 1969
rect 13192 1956 13193 1990
rect 13156 1935 13193 1956
rect 13013 1916 13193 1935
rect 13013 1882 13014 1916
rect 13048 1901 13086 1916
rect 13048 1882 13050 1901
rect 13013 1867 13050 1882
rect 13084 1882 13086 1901
rect 13120 1901 13158 1916
rect 13120 1882 13122 1901
rect 13084 1867 13122 1882
rect 13156 1882 13158 1901
rect 13192 1882 13193 1916
rect 13156 1867 13193 1882
rect 13013 1842 13193 1867
rect 13013 1808 13014 1842
rect 13048 1833 13086 1842
rect 13048 1808 13050 1833
rect 13013 1799 13050 1808
rect 13084 1808 13086 1833
rect 13120 1833 13158 1842
rect 13120 1808 13122 1833
rect 13084 1799 13122 1808
rect 13156 1808 13158 1833
rect 13192 1808 13193 1842
rect 13156 1799 13193 1808
rect 13013 1768 13193 1799
rect 13013 1734 13014 1768
rect 13048 1765 13086 1768
rect 13048 1734 13050 1765
rect 13013 1731 13050 1734
rect 13084 1734 13086 1765
rect 13120 1765 13158 1768
rect 13120 1734 13122 1765
rect 13084 1731 13122 1734
rect 13156 1734 13158 1765
rect 13192 1734 13193 1768
rect 13156 1731 13193 1734
rect 13013 1697 13193 1731
rect 13013 1694 13050 1697
rect 13013 1660 13014 1694
rect 13048 1663 13050 1694
rect 13084 1694 13122 1697
rect 13084 1663 13086 1694
rect 13048 1660 13086 1663
rect 13120 1663 13122 1694
rect 13156 1694 13193 1697
rect 13156 1663 13158 1694
rect 13120 1660 13158 1663
rect 13192 1660 13193 1694
rect 13013 1629 13193 1660
rect 13013 1620 13050 1629
rect 13013 1586 13014 1620
rect 13048 1595 13050 1620
rect 13084 1620 13122 1629
rect 13084 1595 13086 1620
rect 13048 1586 13086 1595
rect 13120 1595 13122 1620
rect 13156 1620 13193 1629
rect 13156 1595 13158 1620
rect 13120 1586 13158 1595
rect 13192 1586 13193 1620
rect 13013 1561 13193 1586
rect 13013 1545 13050 1561
rect 13013 1511 13014 1545
rect 13048 1527 13050 1545
rect 13084 1545 13122 1561
rect 13084 1527 13086 1545
rect 13048 1511 13086 1527
rect 13120 1527 13122 1545
rect 13156 1545 13193 1561
rect 13156 1527 13158 1545
rect 13120 1511 13158 1527
rect 13192 1511 13193 1545
rect 13258 3010 13378 4106
rect 13820 4388 13827 4494
rect 13933 4388 13940 4494
rect 13820 4214 13940 4388
rect 13820 4180 13863 4214
rect 13897 4180 13940 4214
rect 13820 4140 13940 4180
rect 13820 4106 13863 4140
rect 13897 4106 13940 4140
rect 13258 2976 13301 3010
rect 13335 2976 13378 3010
rect 13258 2932 13378 2976
rect 13258 2898 13301 2932
rect 13335 2898 13378 2932
rect 13258 2854 13378 2898
rect 13258 2820 13301 2854
rect 13335 2820 13378 2854
rect 13258 2776 13378 2820
rect 13258 2742 13301 2776
rect 13335 2742 13378 2776
rect 13258 2697 13378 2742
rect 13258 2663 13301 2697
rect 13335 2663 13378 2697
rect 13258 2618 13378 2663
rect 13258 2584 13301 2618
rect 13335 2584 13378 2618
rect 13258 2539 13378 2584
rect 13258 2505 13301 2539
rect 13335 2505 13378 2539
rect 12828 1375 12871 1409
rect 12905 1375 12948 1409
rect 12828 1335 12948 1375
rect 12828 1301 12871 1335
rect 12905 1301 12948 1335
rect 12828 1285 12948 1301
rect 13258 1409 13378 2505
rect 13480 4050 13582 4062
rect 13616 4050 13718 4062
rect 13480 4046 13510 4050
rect 13688 4046 13718 4050
rect 13480 3978 13510 4012
rect 13688 3978 13718 4012
rect 13480 3910 13510 3944
rect 13688 3910 13718 3944
rect 13480 3842 13510 3876
rect 13688 3842 13718 3876
rect 13480 3774 13510 3808
rect 13688 3774 13718 3808
rect 13480 3706 13510 3740
rect 13688 3706 13718 3740
rect 13480 3638 13510 3672
rect 13688 3638 13718 3672
rect 13480 3570 13510 3604
rect 13688 3570 13718 3604
rect 13480 3502 13510 3536
rect 13688 3502 13718 3536
rect 13480 3434 13510 3468
rect 13688 3434 13718 3468
rect 13480 3366 13510 3400
rect 13688 3366 13718 3400
rect 13480 3298 13510 3332
rect 13688 3298 13718 3332
rect 13480 3230 13510 3264
rect 13688 3230 13718 3264
rect 13480 3162 13510 3196
rect 13688 3162 13718 3196
rect 13480 3080 13510 3128
rect 13544 3080 13654 3092
rect 13688 3080 13718 3128
rect 13480 3040 13718 3080
rect 13480 2574 13510 3040
rect 13688 2574 13718 3040
rect 13480 2535 13718 2574
rect 13480 2501 13510 2535
rect 13544 2501 13582 2535
rect 13616 2501 13654 2535
rect 13688 2501 13718 2535
rect 13480 2461 13718 2501
rect 13480 2449 13582 2461
rect 13616 2449 13718 2461
rect 13480 2445 13510 2449
rect 13688 2445 13718 2449
rect 13480 2377 13510 2411
rect 13688 2377 13718 2411
rect 13480 2309 13510 2343
rect 13688 2309 13718 2343
rect 13480 2241 13510 2275
rect 13688 2241 13718 2275
rect 13480 2173 13510 2207
rect 13688 2173 13718 2207
rect 13480 2105 13510 2139
rect 13688 2105 13718 2139
rect 13480 2037 13510 2071
rect 13688 2037 13718 2071
rect 13480 1969 13510 2003
rect 13688 1969 13718 2003
rect 13480 1901 13510 1935
rect 13688 1901 13718 1935
rect 13480 1833 13510 1867
rect 13688 1833 13718 1867
rect 13480 1765 13510 1799
rect 13688 1765 13718 1799
rect 13480 1697 13510 1731
rect 13688 1697 13718 1731
rect 13480 1629 13510 1663
rect 13688 1629 13718 1663
rect 13480 1561 13510 1595
rect 13688 1561 13718 1595
rect 13480 1479 13510 1527
rect 13544 1479 13654 1491
rect 13688 1479 13718 1527
rect 13480 1464 13718 1479
rect 13820 3010 13940 4106
rect 14178 4388 14185 4494
rect 14291 4388 14298 4494
rect 14178 4214 14298 4388
rect 14178 4180 14221 4214
rect 14255 4180 14298 4214
rect 14178 4140 14298 4180
rect 14178 4106 14221 4140
rect 14255 4106 14298 4140
rect 13820 2976 13863 3010
rect 13897 2976 13940 3010
rect 13820 2932 13940 2976
rect 13820 2898 13863 2932
rect 13897 2898 13940 2932
rect 13820 2854 13940 2898
rect 13820 2820 13863 2854
rect 13897 2820 13940 2854
rect 13820 2776 13940 2820
rect 13820 2742 13863 2776
rect 13897 2742 13940 2776
rect 13820 2697 13940 2742
rect 13820 2663 13863 2697
rect 13897 2663 13940 2697
rect 13820 2618 13940 2663
rect 13820 2584 13863 2618
rect 13897 2584 13940 2618
rect 13820 2539 13940 2584
rect 13820 2505 13863 2539
rect 13897 2505 13940 2539
rect 13258 1375 13301 1409
rect 13335 1375 13378 1409
rect 13258 1335 13378 1375
rect 13258 1301 13301 1335
rect 13335 1301 13378 1335
rect 13258 1285 13378 1301
rect 13820 1409 13940 2505
rect 14042 3990 14076 4012
rect 14042 3918 14076 3944
rect 14042 3846 14076 3876
rect 14042 3774 14076 3808
rect 14042 3706 14076 3740
rect 14042 3638 14076 3668
rect 14042 3570 14076 3596
rect 14042 3502 14076 3524
rect 14042 3434 14076 3452
rect 14042 3366 14076 3380
rect 14042 3298 14076 3308
rect 14042 3230 14076 3236
rect 14042 3162 14076 3164
rect 14042 3126 14076 3128
rect 14042 3054 14076 3092
rect 14042 2982 14076 3020
rect 14042 2910 14076 2948
rect 14042 2838 14076 2876
rect 14042 2766 14076 2804
rect 14042 2693 14076 2732
rect 14042 2620 14076 2659
rect 14042 2547 14076 2586
rect 14042 2474 14076 2513
rect 14042 2401 14076 2411
rect 14042 2328 14076 2343
rect 14042 2255 14076 2275
rect 14042 2182 14076 2207
rect 14042 2109 14076 2139
rect 14042 2037 14076 2071
rect 14042 1969 14076 2002
rect 14042 1901 14076 1929
rect 14042 1833 14076 1856
rect 14042 1765 14076 1783
rect 14042 1697 14076 1710
rect 14042 1629 14076 1637
rect 14042 1561 14076 1564
rect 14042 1525 14076 1527
rect 14178 3010 14298 4106
rect 14400 4490 14510 4506
rect 14544 4504 14565 4524
rect 14616 4518 14633 4524
rect 14544 4490 14582 4504
rect 14616 4490 14667 4518
rect 14400 4482 14667 4490
rect 14400 4448 14431 4482
rect 14465 4479 14667 4482
rect 14465 4470 14633 4479
rect 14465 4448 14497 4470
rect 14531 4468 14633 4470
rect 14531 4451 14565 4468
rect 14599 4451 14633 4468
rect 14400 4436 14497 4448
rect 14400 4417 14510 4436
rect 14544 4434 14565 4451
rect 14616 4445 14633 4451
rect 14544 4417 14582 4434
rect 14616 4417 14667 4445
rect 14400 4409 14667 4417
rect 14400 4375 14431 4409
rect 14465 4406 14667 4409
rect 14465 4399 14633 4406
rect 14465 4375 14497 4399
rect 14531 4398 14633 4399
rect 14531 4378 14565 4398
rect 14599 4378 14633 4398
rect 14400 4365 14497 4375
rect 14400 4344 14510 4365
rect 14544 4364 14565 4378
rect 14616 4372 14633 4378
rect 14544 4344 14582 4364
rect 14616 4344 14667 4372
rect 14400 4336 14667 4344
rect 14400 4302 14431 4336
rect 14465 4333 14667 4336
rect 14465 4328 14633 4333
rect 14465 4302 14497 4328
rect 14531 4305 14565 4328
rect 14599 4305 14633 4328
rect 14400 4294 14497 4302
rect 14544 4294 14565 4305
rect 14616 4299 14633 4305
rect 14400 4271 14510 4294
rect 14544 4271 14582 4294
rect 14616 4271 14667 4299
rect 14400 4263 14667 4271
rect 14400 4229 14431 4263
rect 14465 4260 14667 4263
rect 14465 4257 14633 4260
rect 14465 4229 14497 4257
rect 14531 4232 14565 4257
rect 14599 4232 14633 4257
rect 14400 4223 14497 4229
rect 14544 4223 14565 4232
rect 14616 4226 14633 4232
rect 14400 4198 14510 4223
rect 14544 4198 14582 4223
rect 14616 4198 14667 4226
rect 14400 4190 14667 4198
rect 14400 4156 14431 4190
rect 14465 4186 14667 4190
rect 14465 4156 14497 4186
rect 14531 4159 14565 4186
rect 14599 4159 14633 4186
rect 14400 4152 14497 4156
rect 14544 4152 14565 4159
rect 14616 4152 14633 4159
rect 14400 4125 14510 4152
rect 14544 4125 14582 4152
rect 14616 4125 14667 4152
rect 14400 4117 14667 4125
rect 14400 4083 14431 4117
rect 14465 4115 14667 4117
rect 14465 4086 14565 4115
rect 14599 4086 14633 4115
rect 14465 4083 14510 4086
rect 14400 4062 14510 4083
rect 14386 4052 14510 4062
rect 14544 4081 14565 4086
rect 14616 4081 14633 4086
rect 14544 4052 14582 4081
rect 14616 4052 14667 4081
rect 14386 4046 14667 4052
rect 14420 4044 14667 4046
rect 14420 4012 14431 4044
rect 14465 4041 14667 4044
rect 14465 4034 14565 4041
rect 14386 4010 14431 4012
rect 14488 4013 14565 4034
rect 14599 4013 14633 4041
rect 14386 4000 14454 4010
rect 14488 4000 14510 4013
rect 14386 3979 14510 4000
rect 14544 4007 14565 4013
rect 14616 4007 14633 4013
rect 14544 3979 14582 4007
rect 14616 3979 14667 4007
rect 14386 3978 14667 3979
rect 14420 3971 14667 3978
rect 14420 3944 14431 3971
rect 14465 3970 14667 3971
rect 14465 3966 14565 3970
rect 14386 3937 14431 3944
rect 14488 3940 14565 3966
rect 14599 3940 14633 3970
rect 14386 3932 14454 3937
rect 14488 3932 14510 3940
rect 14386 3910 14510 3932
rect 14420 3906 14510 3910
rect 14544 3936 14565 3940
rect 14616 3936 14633 3940
rect 14544 3906 14582 3936
rect 14616 3906 14667 3936
rect 14420 3898 14667 3906
rect 14420 3876 14431 3898
rect 14386 3864 14431 3876
rect 14488 3896 14667 3898
rect 14488 3867 14565 3896
rect 14599 3867 14633 3896
rect 14488 3864 14510 3867
rect 14386 3842 14510 3864
rect 14420 3833 14510 3842
rect 14544 3862 14565 3867
rect 14616 3862 14633 3867
rect 14544 3833 14582 3862
rect 14616 3833 14667 3862
rect 14420 3830 14667 3833
rect 14420 3825 14454 3830
rect 14488 3825 14667 3830
rect 14420 3808 14431 3825
rect 14386 3791 14431 3808
rect 14488 3796 14565 3825
rect 14465 3794 14565 3796
rect 14599 3794 14633 3825
rect 14465 3791 14510 3794
rect 14386 3774 14510 3791
rect 14420 3762 14510 3774
rect 14420 3752 14454 3762
rect 14488 3760 14510 3762
rect 14544 3791 14565 3794
rect 14616 3791 14633 3794
rect 14544 3760 14582 3791
rect 14616 3760 14667 3791
rect 14420 3740 14431 3752
rect 14386 3718 14431 3740
rect 14488 3751 14667 3760
rect 14488 3728 14565 3751
rect 14465 3721 14565 3728
rect 14599 3721 14633 3751
rect 14465 3718 14510 3721
rect 14386 3706 14510 3718
rect 14420 3694 14510 3706
rect 14420 3679 14454 3694
rect 14488 3687 14510 3694
rect 14544 3717 14565 3721
rect 14616 3717 14633 3721
rect 14544 3687 14582 3717
rect 14616 3687 14667 3717
rect 14488 3680 14667 3687
rect 14420 3672 14431 3679
rect 14386 3645 14431 3672
rect 14488 3660 14565 3680
rect 14465 3648 14565 3660
rect 14599 3648 14633 3680
rect 14465 3645 14510 3648
rect 14386 3638 14510 3645
rect 14420 3626 14510 3638
rect 14420 3606 14454 3626
rect 14488 3614 14510 3626
rect 14544 3646 14565 3648
rect 14616 3646 14633 3648
rect 14544 3614 14582 3646
rect 14616 3614 14667 3646
rect 14488 3606 14667 3614
rect 14420 3604 14431 3606
rect 14386 3572 14431 3604
rect 14488 3592 14565 3606
rect 14465 3575 14565 3592
rect 14599 3575 14633 3606
rect 14465 3572 14510 3575
rect 14386 3570 14510 3572
rect 14420 3558 14510 3570
rect 14420 3536 14454 3558
rect 14386 3533 14454 3536
rect 14488 3541 14510 3558
rect 14544 3572 14565 3575
rect 14616 3572 14633 3575
rect 14544 3541 14582 3572
rect 14616 3541 14667 3572
rect 14488 3535 14667 3541
rect 14386 3502 14431 3533
rect 14488 3524 14565 3535
rect 14420 3499 14431 3502
rect 14465 3502 14565 3524
rect 14599 3502 14633 3535
rect 14465 3499 14510 3502
rect 14420 3490 14510 3499
rect 14420 3468 14454 3490
rect 14386 3460 14454 3468
rect 14488 3468 14510 3490
rect 14544 3501 14565 3502
rect 14616 3501 14633 3502
rect 14544 3468 14582 3501
rect 14616 3468 14667 3501
rect 14488 3461 14667 3468
rect 14386 3434 14431 3460
rect 14488 3456 14565 3461
rect 14420 3426 14431 3434
rect 14465 3429 14565 3456
rect 14599 3429 14633 3461
rect 14465 3426 14510 3429
rect 14420 3422 14510 3426
rect 14420 3400 14454 3422
rect 14386 3388 14454 3400
rect 14488 3395 14510 3422
rect 14544 3427 14565 3429
rect 14616 3427 14633 3429
rect 14544 3395 14582 3427
rect 14616 3395 14667 3427
rect 14488 3390 14667 3395
rect 14488 3388 14565 3390
rect 14386 3387 14565 3388
rect 14386 3366 14431 3387
rect 14420 3353 14431 3366
rect 14465 3356 14565 3387
rect 14599 3356 14633 3390
rect 14465 3354 14510 3356
rect 14420 3332 14454 3353
rect 14386 3320 14454 3332
rect 14488 3322 14510 3354
rect 14544 3322 14582 3356
rect 14616 3322 14667 3356
rect 14488 3320 14667 3322
rect 14386 3316 14667 3320
rect 14386 3314 14565 3316
rect 14386 3298 14431 3314
rect 14420 3280 14431 3298
rect 14465 3286 14565 3314
rect 14488 3283 14565 3286
rect 14599 3283 14633 3316
rect 14420 3264 14454 3280
rect 14386 3252 14454 3264
rect 14488 3252 14510 3283
rect 14386 3249 14510 3252
rect 14544 3282 14565 3283
rect 14616 3282 14633 3283
rect 14544 3249 14582 3282
rect 14616 3249 14667 3282
rect 14386 3245 14667 3249
rect 14386 3241 14565 3245
rect 14386 3230 14431 3241
rect 14420 3207 14431 3230
rect 14465 3218 14565 3241
rect 14488 3211 14565 3218
rect 14599 3211 14633 3245
rect 14488 3210 14667 3211
rect 14420 3196 14454 3207
rect 14386 3184 14454 3196
rect 14488 3184 14510 3210
rect 14386 3176 14510 3184
rect 14544 3176 14582 3210
rect 14616 3176 14667 3210
rect 14386 3168 14667 3176
rect 14386 3162 14431 3168
rect 14420 3134 14431 3162
rect 14465 3151 14667 3168
rect 14465 3150 14565 3151
rect 14488 3137 14565 3150
rect 14599 3137 14633 3151
rect 14420 3128 14454 3134
rect 14386 3116 14454 3128
rect 14488 3116 14510 3137
rect 14386 3103 14510 3116
rect 14544 3117 14565 3137
rect 14616 3117 14633 3137
rect 14544 3103 14582 3117
rect 14616 3103 14667 3117
rect 14386 3100 14667 3103
rect 14178 2976 14221 3010
rect 14255 2976 14298 3010
rect 14178 2932 14298 2976
rect 14178 2898 14221 2932
rect 14255 2898 14298 2932
rect 14178 2854 14298 2898
rect 14178 2820 14221 2854
rect 14255 2820 14298 2854
rect 14178 2776 14298 2820
rect 14178 2742 14221 2776
rect 14255 2742 14298 2776
rect 14178 2697 14298 2742
rect 14178 2663 14221 2697
rect 14255 2663 14298 2697
rect 14178 2618 14298 2663
rect 14178 2584 14221 2618
rect 14255 2584 14298 2618
rect 14178 2539 14298 2584
rect 14178 2505 14221 2539
rect 14255 2505 14298 2539
rect 13820 1375 13863 1409
rect 13897 1375 13940 1409
rect 13820 1335 13940 1375
rect 13820 1301 13863 1335
rect 13897 1301 13940 1335
rect 13820 1285 13940 1301
rect 14178 1409 14298 2505
rect 14400 3095 14667 3100
rect 14400 3061 14431 3095
rect 14465 3066 14667 3095
rect 14465 3064 14565 3066
rect 14599 3064 14633 3066
rect 14465 3061 14510 3064
rect 14400 3030 14510 3061
rect 14544 3032 14565 3064
rect 14616 3032 14633 3064
rect 14544 3030 14582 3032
rect 14616 3030 14667 3032
rect 14400 3022 14667 3030
rect 14400 2988 14431 3022
rect 14465 2991 14667 3022
rect 14465 2988 14510 2991
rect 14400 2972 14510 2988
rect 14544 2972 14582 2991
rect 14616 2972 14667 2991
rect 14400 2949 14497 2972
rect 14400 2915 14431 2949
rect 14465 2915 14497 2949
rect 14400 2876 14497 2915
rect 14400 2842 14431 2876
rect 14465 2842 14497 2876
rect 14400 2803 14497 2842
rect 14400 2769 14431 2803
rect 14465 2769 14497 2803
rect 14400 2730 14497 2769
rect 14400 2696 14431 2730
rect 14465 2696 14497 2730
rect 14400 2657 14497 2696
rect 14400 2623 14431 2657
rect 14465 2623 14497 2657
rect 14400 2584 14497 2623
rect 14400 2550 14431 2584
rect 14465 2550 14497 2584
rect 14400 2530 14497 2550
rect 14400 2519 14510 2530
rect 14544 2519 14582 2530
rect 14616 2519 14667 2530
rect 14400 2511 14667 2519
rect 14400 2477 14431 2511
rect 14465 2485 14667 2511
rect 14465 2480 14565 2485
rect 14599 2480 14633 2485
rect 14465 2477 14510 2480
rect 14400 2461 14510 2477
rect 14386 2446 14510 2461
rect 14544 2451 14565 2480
rect 14616 2451 14633 2480
rect 14544 2446 14582 2451
rect 14616 2446 14667 2451
rect 14386 2445 14667 2446
rect 14420 2438 14667 2445
rect 14420 2411 14431 2438
rect 14465 2433 14667 2438
rect 14386 2404 14431 2411
rect 14488 2407 14667 2433
rect 14386 2399 14454 2404
rect 14488 2399 14510 2407
rect 14386 2377 14510 2399
rect 14420 2373 14510 2377
rect 14544 2403 14582 2407
rect 14616 2403 14667 2407
rect 14544 2373 14565 2403
rect 14616 2373 14633 2403
rect 14420 2369 14565 2373
rect 14599 2369 14633 2373
rect 14420 2365 14667 2369
rect 14420 2343 14431 2365
rect 14386 2331 14431 2343
rect 14488 2334 14667 2365
rect 14488 2331 14510 2334
rect 14386 2309 14510 2331
rect 14420 2300 14510 2309
rect 14544 2327 14582 2334
rect 14616 2327 14667 2334
rect 14544 2300 14565 2327
rect 14616 2300 14633 2327
rect 14420 2297 14565 2300
rect 14420 2292 14454 2297
rect 14488 2293 14565 2297
rect 14599 2293 14633 2300
rect 14420 2275 14431 2292
rect 14386 2258 14431 2275
rect 14488 2263 14667 2293
rect 14465 2260 14667 2263
rect 14465 2258 14510 2260
rect 14386 2241 14510 2258
rect 14420 2229 14510 2241
rect 14420 2219 14454 2229
rect 14488 2226 14510 2229
rect 14544 2250 14582 2260
rect 14616 2250 14667 2260
rect 14544 2226 14565 2250
rect 14616 2226 14633 2250
rect 14420 2207 14431 2219
rect 14386 2185 14431 2207
rect 14488 2216 14565 2226
rect 14599 2216 14633 2226
rect 14488 2195 14667 2216
rect 14465 2186 14667 2195
rect 14465 2185 14510 2186
rect 14386 2173 14510 2185
rect 14420 2161 14510 2173
rect 14420 2146 14454 2161
rect 14488 2152 14510 2161
rect 14544 2156 14582 2186
rect 14616 2156 14667 2186
rect 14544 2152 14565 2156
rect 14616 2152 14633 2156
rect 14420 2139 14431 2146
rect 14386 2112 14431 2139
rect 14488 2127 14565 2152
rect 14465 2122 14565 2127
rect 14599 2122 14633 2152
rect 14465 2112 14667 2122
rect 14386 2105 14510 2112
rect 14420 2093 14510 2105
rect 14420 2073 14454 2093
rect 14488 2078 14510 2093
rect 14544 2085 14582 2112
rect 14616 2085 14667 2112
rect 14544 2078 14565 2085
rect 14616 2078 14633 2085
rect 14420 2071 14431 2073
rect 14386 2039 14431 2071
rect 14488 2059 14565 2078
rect 14465 2051 14565 2059
rect 14599 2051 14633 2078
rect 14465 2039 14667 2051
rect 14386 2038 14667 2039
rect 14386 2037 14510 2038
rect 14420 2025 14510 2037
rect 14420 2003 14454 2025
rect 14386 2000 14454 2003
rect 14488 2004 14510 2025
rect 14544 2011 14582 2038
rect 14616 2011 14667 2038
rect 14544 2004 14565 2011
rect 14616 2004 14633 2011
rect 14386 1969 14431 2000
rect 14488 1991 14565 2004
rect 14420 1966 14431 1969
rect 14465 1977 14565 1991
rect 14599 1977 14633 2004
rect 14465 1966 14667 1977
rect 14420 1964 14667 1966
rect 14420 1957 14510 1964
rect 14420 1935 14454 1957
rect 14386 1927 14454 1935
rect 14488 1930 14510 1957
rect 14544 1940 14582 1964
rect 14616 1940 14667 1964
rect 14544 1930 14565 1940
rect 14616 1930 14633 1940
rect 14386 1901 14431 1927
rect 14488 1923 14565 1930
rect 14420 1893 14431 1901
rect 14465 1906 14565 1923
rect 14599 1906 14633 1930
rect 14465 1893 14667 1906
rect 14420 1890 14667 1893
rect 14420 1889 14510 1890
rect 14420 1867 14454 1889
rect 14386 1855 14454 1867
rect 14488 1856 14510 1889
rect 14544 1866 14582 1890
rect 14616 1866 14667 1890
rect 14544 1856 14565 1866
rect 14616 1856 14633 1866
rect 14488 1855 14565 1856
rect 14386 1854 14565 1855
rect 14386 1833 14431 1854
rect 14420 1820 14431 1833
rect 14465 1832 14565 1854
rect 14599 1832 14633 1856
rect 14465 1821 14667 1832
rect 14420 1799 14454 1820
rect 14386 1787 14454 1799
rect 14488 1816 14667 1821
rect 14488 1787 14510 1816
rect 14386 1782 14510 1787
rect 14544 1795 14582 1816
rect 14616 1795 14667 1816
rect 14544 1782 14565 1795
rect 14616 1782 14633 1795
rect 14386 1781 14565 1782
rect 14386 1765 14431 1781
rect 14420 1747 14431 1765
rect 14465 1761 14565 1781
rect 14599 1761 14633 1782
rect 14465 1753 14667 1761
rect 14420 1731 14454 1747
rect 14386 1719 14454 1731
rect 14488 1742 14667 1753
rect 14488 1719 14510 1742
rect 14386 1708 14510 1719
rect 14544 1721 14582 1742
rect 14616 1721 14667 1742
rect 14544 1708 14565 1721
rect 14616 1708 14633 1721
rect 14386 1697 14431 1708
rect 14420 1674 14431 1697
rect 14465 1687 14565 1708
rect 14599 1687 14633 1708
rect 14465 1685 14667 1687
rect 14420 1663 14454 1674
rect 14386 1651 14454 1663
rect 14488 1668 14667 1685
rect 14488 1651 14510 1668
rect 14386 1635 14510 1651
rect 14386 1629 14431 1635
rect 14420 1601 14431 1629
rect 14465 1634 14510 1635
rect 14544 1650 14582 1668
rect 14616 1650 14667 1668
rect 14544 1634 14565 1650
rect 14616 1634 14633 1650
rect 14465 1617 14565 1634
rect 14488 1616 14565 1617
rect 14599 1616 14633 1634
rect 14420 1595 14454 1601
rect 14386 1583 14454 1595
rect 14488 1594 14667 1616
rect 14488 1583 14510 1594
rect 14386 1562 14510 1583
rect 14386 1561 14431 1562
rect 14420 1528 14431 1561
rect 14465 1560 14510 1562
rect 14544 1576 14582 1594
rect 14616 1576 14667 1594
rect 14544 1560 14565 1576
rect 14616 1560 14633 1576
rect 14465 1549 14565 1560
rect 14488 1542 14565 1549
rect 14599 1542 14633 1560
rect 14420 1527 14454 1528
rect 14386 1515 14454 1527
rect 14488 1520 14667 1542
rect 14488 1515 14510 1520
rect 14386 1499 14510 1515
rect 14178 1375 14221 1409
rect 14255 1375 14298 1409
rect 14178 1335 14298 1375
rect 14178 1301 14221 1335
rect 14255 1301 14298 1335
rect 14178 1285 14298 1301
rect 14400 1489 14510 1499
rect 14400 1455 14431 1489
rect 14465 1486 14510 1489
rect 14544 1505 14582 1520
rect 14616 1505 14667 1520
rect 14544 1486 14565 1505
rect 14616 1486 14633 1505
rect 14465 1471 14565 1486
rect 14599 1471 14633 1486
rect 14465 1455 14667 1471
rect 14400 1446 14667 1455
rect 14400 1416 14510 1446
rect 14400 1382 14431 1416
rect 14465 1412 14510 1416
rect 14544 1412 14582 1446
rect 14616 1412 14667 1446
rect 14465 1387 14667 1412
rect 14465 1382 14497 1387
rect 14400 1353 14497 1382
rect 14531 1372 14565 1387
rect 14599 1372 14633 1387
rect 14544 1353 14565 1372
rect 14616 1353 14633 1372
rect 14400 1342 14510 1353
rect 14400 1308 14431 1342
rect 14465 1338 14510 1342
rect 14544 1338 14582 1353
rect 14616 1338 14667 1353
rect 14465 1319 14667 1338
rect 14465 1311 14633 1319
rect 14465 1308 14565 1311
rect 555 1241 733 1268
rect 555 1221 587 1241
rect 621 1221 659 1241
rect 621 1207 623 1221
rect 589 1187 623 1207
rect 657 1207 659 1221
rect 693 1234 733 1241
rect 767 1234 822 1268
rect 693 1219 822 1234
rect 657 1187 691 1207
rect 555 1185 691 1187
rect 725 1194 822 1219
rect 725 1185 733 1194
rect 555 1160 733 1185
rect 767 1160 822 1194
rect 555 1150 822 1160
rect 555 1140 623 1150
rect 589 1116 623 1140
rect 657 1148 822 1150
rect 14400 1274 14497 1308
rect 14531 1298 14565 1308
rect 14599 1298 14633 1311
rect 14544 1277 14565 1298
rect 14616 1285 14633 1298
rect 14400 1268 14510 1274
rect 14400 1234 14431 1268
rect 14465 1264 14510 1268
rect 14544 1264 14582 1277
rect 14616 1264 14667 1285
rect 14465 1251 14667 1264
rect 14465 1234 14633 1251
rect 14400 1228 14565 1234
rect 14400 1194 14497 1228
rect 14531 1224 14565 1228
rect 14599 1224 14633 1234
rect 14544 1200 14565 1224
rect 14616 1217 14633 1224
rect 14400 1160 14431 1194
rect 14465 1190 14510 1194
rect 14544 1190 14582 1200
rect 14616 1190 14667 1217
rect 14465 1183 14667 1190
rect 14465 1160 14633 1183
rect 14400 1157 14633 1160
rect 14400 1148 14565 1157
rect 657 1116 691 1148
rect 589 1114 691 1116
rect 725 1114 760 1148
rect 794 1116 829 1148
rect 14531 1123 14565 1148
rect 14599 1149 14633 1157
rect 14599 1123 14667 1149
rect 589 1106 767 1114
rect 555 1082 767 1106
rect 801 1082 829 1116
rect 555 1080 829 1082
rect 555 1046 623 1080
rect 657 1046 692 1080
rect 726 1046 761 1080
rect 555 1012 761 1046
rect 555 978 589 1012
rect 623 978 658 1012
rect 692 978 727 1012
rect 14531 1115 14667 1123
rect 14531 1081 14633 1115
rect 14531 1080 14667 1081
rect 14599 1046 14667 1080
rect 14565 1012 14633 1046
rect 14565 978 14667 1012
rect 249 664 308 668
rect 249 630 294 664
rect 249 596 308 630
rect 249 562 294 596
rect 249 528 308 562
rect 249 496 294 528
rect 67 494 294 496
rect 67 490 308 494
rect 14886 490 14927 668
rect 15105 490 15106 5420
<< viali >>
rect 71 5303 249 5426
rect 308 5422 14886 5426
rect 71 5269 105 5303
rect 105 5269 139 5303
rect 139 5269 173 5303
rect 173 5269 207 5303
rect 207 5269 241 5303
rect 241 5269 249 5303
rect 71 5232 249 5269
rect 308 5252 10868 5422
rect 10868 5388 10903 5422
rect 10903 5388 10937 5422
rect 10937 5388 10972 5422
rect 10972 5388 11006 5422
rect 11006 5388 11041 5422
rect 11041 5388 11075 5422
rect 11075 5388 11110 5422
rect 11110 5388 11144 5422
rect 11144 5388 11179 5422
rect 11179 5388 11213 5422
rect 11213 5388 11248 5422
rect 11248 5388 11282 5422
rect 11282 5388 11317 5422
rect 11317 5388 11351 5422
rect 11351 5388 11386 5422
rect 11386 5388 11420 5422
rect 11420 5388 11455 5422
rect 11455 5388 11489 5422
rect 11489 5388 11524 5422
rect 11524 5388 11558 5422
rect 11558 5388 11593 5422
rect 11593 5388 11627 5422
rect 11627 5388 11662 5422
rect 11662 5388 11696 5422
rect 11696 5388 11731 5422
rect 11731 5388 11765 5422
rect 11765 5388 11800 5422
rect 11800 5388 11834 5422
rect 11834 5388 11869 5422
rect 11869 5388 11903 5422
rect 11903 5388 11938 5422
rect 11938 5388 11972 5422
rect 11972 5388 12007 5422
rect 12007 5388 12041 5422
rect 12041 5388 12076 5422
rect 12076 5388 12110 5422
rect 12110 5388 12145 5422
rect 12145 5388 12179 5422
rect 12179 5388 12214 5422
rect 12214 5388 12248 5422
rect 12248 5388 12283 5422
rect 12283 5388 12317 5422
rect 12317 5388 12352 5422
rect 12352 5388 12386 5422
rect 12386 5388 12421 5422
rect 12421 5388 12455 5422
rect 12455 5388 12490 5422
rect 12490 5388 12524 5422
rect 12524 5388 12559 5422
rect 12559 5388 12593 5422
rect 12593 5388 12628 5422
rect 12628 5388 12662 5422
rect 12662 5388 12697 5422
rect 12697 5388 12731 5422
rect 12731 5388 12766 5422
rect 12766 5388 12800 5422
rect 12800 5388 12835 5422
rect 12835 5388 12869 5422
rect 12869 5388 12904 5422
rect 12904 5388 12938 5422
rect 12938 5388 12973 5422
rect 12973 5388 13007 5422
rect 13007 5388 13042 5422
rect 13042 5388 13076 5422
rect 13076 5388 13111 5422
rect 13111 5388 13145 5422
rect 13145 5388 13180 5422
rect 13180 5388 13214 5422
rect 13214 5388 13249 5422
rect 13249 5388 13283 5422
rect 13283 5388 13318 5422
rect 13318 5388 13352 5422
rect 13352 5388 13387 5422
rect 13387 5388 13421 5422
rect 13421 5388 13456 5422
rect 13456 5388 13490 5422
rect 13490 5388 13525 5422
rect 13525 5388 13559 5422
rect 13559 5388 13594 5422
rect 13594 5388 13628 5422
rect 13628 5388 13663 5422
rect 13663 5388 13697 5422
rect 13697 5388 13732 5422
rect 13732 5388 13766 5422
rect 13766 5388 13801 5422
rect 13801 5388 13835 5422
rect 13835 5388 13870 5422
rect 13870 5388 13904 5422
rect 13904 5388 13939 5422
rect 13939 5388 13973 5422
rect 13973 5388 14008 5422
rect 14008 5388 14042 5422
rect 14042 5388 14077 5422
rect 14077 5388 14111 5422
rect 14111 5388 14146 5422
rect 14146 5388 14180 5422
rect 14180 5388 14215 5422
rect 14215 5388 14249 5422
rect 14249 5388 14284 5422
rect 14284 5388 14318 5422
rect 14318 5388 14353 5422
rect 14353 5388 14387 5422
rect 14387 5388 14422 5422
rect 14422 5388 14456 5422
rect 14456 5388 14491 5422
rect 14491 5388 14525 5422
rect 14525 5388 14560 5422
rect 14560 5388 14594 5422
rect 14594 5388 14629 5422
rect 14629 5388 14663 5422
rect 14663 5388 14698 5422
rect 14698 5388 14732 5422
rect 14732 5388 14767 5422
rect 14767 5388 14801 5422
rect 14801 5388 14836 5422
rect 14836 5388 14870 5422
rect 14870 5388 14886 5422
rect 10868 5354 14886 5388
rect 10868 5320 10903 5354
rect 10903 5320 10937 5354
rect 10937 5320 10972 5354
rect 10972 5320 11006 5354
rect 11006 5320 11041 5354
rect 11041 5320 11075 5354
rect 11075 5320 11110 5354
rect 11110 5320 11144 5354
rect 11144 5320 11179 5354
rect 11179 5320 11213 5354
rect 11213 5320 11248 5354
rect 11248 5320 11282 5354
rect 11282 5320 11317 5354
rect 11317 5320 11351 5354
rect 11351 5320 11386 5354
rect 11386 5320 11420 5354
rect 11420 5320 11455 5354
rect 11455 5320 11489 5354
rect 11489 5320 11524 5354
rect 11524 5320 11558 5354
rect 11558 5320 11593 5354
rect 11593 5320 11627 5354
rect 11627 5320 11662 5354
rect 11662 5320 11696 5354
rect 11696 5320 11731 5354
rect 11731 5320 11765 5354
rect 11765 5320 11800 5354
rect 11800 5320 11834 5354
rect 11834 5320 11869 5354
rect 11869 5320 11903 5354
rect 11903 5320 11938 5354
rect 11938 5320 11972 5354
rect 11972 5320 12007 5354
rect 12007 5320 12041 5354
rect 12041 5320 12076 5354
rect 12076 5320 12110 5354
rect 12110 5320 12145 5354
rect 12145 5320 12179 5354
rect 12179 5320 12214 5354
rect 12214 5320 12248 5354
rect 12248 5320 12283 5354
rect 12283 5320 12317 5354
rect 12317 5320 12352 5354
rect 12352 5320 12386 5354
rect 12386 5320 12421 5354
rect 12421 5320 12455 5354
rect 12455 5320 12490 5354
rect 12490 5320 12524 5354
rect 12524 5320 12559 5354
rect 12559 5320 12593 5354
rect 12593 5320 12628 5354
rect 12628 5320 12662 5354
rect 12662 5320 12697 5354
rect 12697 5320 12731 5354
rect 12731 5320 12766 5354
rect 12766 5320 12800 5354
rect 12800 5320 12835 5354
rect 12835 5320 12869 5354
rect 12869 5320 12904 5354
rect 12904 5320 12938 5354
rect 12938 5320 12973 5354
rect 12973 5320 13007 5354
rect 13007 5320 13042 5354
rect 13042 5320 13076 5354
rect 13076 5320 13111 5354
rect 13111 5320 13145 5354
rect 13145 5320 13180 5354
rect 13180 5320 13214 5354
rect 13214 5320 13249 5354
rect 13249 5320 13283 5354
rect 13283 5320 13318 5354
rect 13318 5320 13352 5354
rect 13352 5320 13387 5354
rect 13387 5320 13421 5354
rect 13421 5320 13456 5354
rect 13456 5320 13490 5354
rect 13490 5320 13525 5354
rect 13525 5320 13559 5354
rect 13559 5320 13594 5354
rect 13594 5320 13628 5354
rect 13628 5320 13663 5354
rect 13663 5320 13697 5354
rect 13697 5320 13732 5354
rect 13732 5320 13766 5354
rect 13766 5320 13801 5354
rect 13801 5320 13835 5354
rect 13835 5320 13870 5354
rect 13870 5320 13904 5354
rect 13904 5320 13939 5354
rect 13939 5320 13973 5354
rect 13973 5320 14008 5354
rect 14008 5320 14042 5354
rect 14042 5320 14077 5354
rect 14077 5320 14111 5354
rect 14111 5320 14146 5354
rect 14146 5320 14180 5354
rect 14180 5320 14215 5354
rect 14215 5320 14249 5354
rect 14249 5320 14284 5354
rect 14284 5320 14318 5354
rect 14318 5320 14353 5354
rect 14353 5320 14387 5354
rect 14387 5320 14422 5354
rect 14422 5320 14456 5354
rect 14456 5320 14491 5354
rect 14491 5320 14525 5354
rect 14525 5320 14560 5354
rect 14560 5320 14594 5354
rect 14594 5320 14629 5354
rect 14629 5320 14663 5354
rect 14663 5320 14698 5354
rect 14698 5320 14732 5354
rect 14732 5320 14767 5354
rect 14767 5320 14801 5354
rect 14801 5320 14836 5354
rect 14836 5320 14870 5354
rect 14870 5320 14886 5354
rect 10868 5286 14886 5320
rect 10868 5252 10903 5286
rect 10903 5252 10937 5286
rect 10937 5252 10972 5286
rect 10972 5252 11006 5286
rect 11006 5252 11041 5286
rect 11041 5252 11075 5286
rect 11075 5252 11110 5286
rect 11110 5252 11144 5286
rect 11144 5252 11179 5286
rect 11179 5252 11213 5286
rect 11213 5252 11248 5286
rect 11248 5252 11282 5286
rect 11282 5252 11317 5286
rect 11317 5252 11351 5286
rect 11351 5252 11386 5286
rect 11386 5252 11420 5286
rect 11420 5252 11455 5286
rect 11455 5252 11489 5286
rect 11489 5252 11524 5286
rect 11524 5252 11558 5286
rect 11558 5252 11593 5286
rect 11593 5252 11627 5286
rect 11627 5252 11662 5286
rect 11662 5252 11696 5286
rect 11696 5252 11731 5286
rect 11731 5252 11765 5286
rect 11765 5252 11800 5286
rect 11800 5252 11834 5286
rect 11834 5252 11869 5286
rect 11869 5252 11903 5286
rect 11903 5252 11938 5286
rect 11938 5252 11972 5286
rect 11972 5252 12007 5286
rect 12007 5252 12041 5286
rect 12041 5252 12076 5286
rect 12076 5252 12110 5286
rect 12110 5252 12145 5286
rect 12145 5252 12179 5286
rect 12179 5252 12214 5286
rect 12214 5252 12248 5286
rect 12248 5252 12283 5286
rect 12283 5252 12317 5286
rect 12317 5252 12352 5286
rect 12352 5252 12386 5286
rect 12386 5252 12421 5286
rect 12421 5252 12455 5286
rect 12455 5252 12490 5286
rect 12490 5252 12524 5286
rect 12524 5252 12559 5286
rect 12559 5252 12593 5286
rect 12593 5252 12628 5286
rect 12628 5252 12662 5286
rect 12662 5252 12697 5286
rect 12697 5252 12731 5286
rect 12731 5252 12766 5286
rect 12766 5252 12800 5286
rect 12800 5252 12835 5286
rect 12835 5252 12869 5286
rect 12869 5252 12904 5286
rect 12904 5252 12938 5286
rect 12938 5252 12973 5286
rect 12973 5252 13007 5286
rect 13007 5252 13042 5286
rect 13042 5252 13076 5286
rect 13076 5252 13111 5286
rect 13111 5252 13145 5286
rect 13145 5252 13180 5286
rect 13180 5252 13214 5286
rect 13214 5252 13249 5286
rect 13249 5252 13283 5286
rect 13283 5252 13318 5286
rect 13318 5252 13352 5286
rect 13352 5252 13387 5286
rect 13387 5252 13421 5286
rect 13421 5252 13456 5286
rect 13456 5252 13490 5286
rect 13490 5252 13525 5286
rect 13525 5252 13559 5286
rect 13559 5252 13594 5286
rect 13594 5252 13628 5286
rect 13628 5252 13663 5286
rect 13663 5252 13697 5286
rect 13697 5252 13732 5286
rect 13732 5252 13766 5286
rect 13766 5252 13801 5286
rect 13801 5252 13835 5286
rect 13835 5252 13870 5286
rect 13870 5252 13904 5286
rect 13904 5252 13939 5286
rect 13939 5252 13973 5286
rect 13973 5252 14008 5286
rect 14008 5252 14042 5286
rect 14042 5252 14077 5286
rect 14077 5252 14111 5286
rect 14111 5252 14146 5286
rect 14146 5252 14180 5286
rect 14180 5252 14215 5286
rect 14215 5252 14249 5286
rect 14249 5252 14284 5286
rect 14284 5252 14318 5286
rect 14318 5252 14353 5286
rect 14353 5252 14387 5286
rect 14387 5252 14422 5286
rect 14422 5252 14456 5286
rect 14456 5252 14491 5286
rect 14491 5252 14525 5286
rect 14525 5252 14560 5286
rect 14560 5252 14594 5286
rect 14594 5252 14629 5286
rect 14629 5252 14663 5286
rect 14663 5252 14698 5286
rect 14698 5252 14732 5286
rect 14732 5252 14767 5286
rect 14767 5252 14801 5286
rect 14801 5252 14836 5286
rect 14836 5252 14870 5286
rect 14870 5252 14886 5286
rect 308 5248 14886 5252
rect 14927 5328 15105 5420
rect 14927 5294 14935 5328
rect 14935 5294 14969 5328
rect 14969 5294 15003 5328
rect 15003 5294 15037 5328
rect 15037 5294 15071 5328
rect 15071 5294 15105 5328
rect 14927 5256 15105 5294
rect 71 5198 105 5232
rect 105 5198 139 5232
rect 139 5198 173 5232
rect 173 5198 207 5232
rect 207 5198 241 5232
rect 241 5198 249 5232
rect 71 5161 249 5198
rect 71 5127 105 5161
rect 105 5127 139 5161
rect 139 5127 173 5161
rect 173 5127 207 5161
rect 207 5127 241 5161
rect 241 5127 249 5161
rect 71 5090 249 5127
rect 71 5056 105 5090
rect 105 5056 139 5090
rect 139 5056 173 5090
rect 173 5056 207 5090
rect 207 5056 241 5090
rect 241 5056 249 5090
rect 71 5020 249 5056
rect 71 4986 105 5020
rect 105 4986 139 5020
rect 139 4986 173 5020
rect 173 4986 207 5020
rect 207 4986 241 5020
rect 241 4986 249 5020
rect 71 4918 249 4986
rect 14927 5222 14935 5256
rect 14935 5222 14969 5256
rect 14969 5222 15003 5256
rect 15003 5222 15037 5256
rect 15037 5222 15071 5256
rect 15071 5222 15105 5256
rect 14927 5184 15105 5222
rect 14927 5150 14935 5184
rect 14935 5150 14969 5184
rect 14969 5150 15003 5184
rect 15003 5150 15037 5184
rect 15037 5150 15071 5184
rect 15071 5150 15105 5184
rect 14927 5112 15105 5150
rect 14927 5078 14935 5112
rect 14935 5078 14969 5112
rect 14969 5078 15003 5112
rect 15003 5078 15037 5112
rect 15037 5078 15071 5112
rect 15071 5078 15105 5112
rect 14927 5040 15105 5078
rect 14927 5006 14935 5040
rect 14935 5006 14969 5040
rect 14969 5006 15003 5040
rect 15003 5006 15037 5040
rect 15037 5006 15071 5040
rect 15071 5006 15105 5040
rect 14927 4968 15105 5006
rect 71 4884 105 4918
rect 105 4884 139 4918
rect 139 4884 173 4918
rect 173 4884 207 4918
rect 207 4884 241 4918
rect 241 4884 249 4918
rect 71 4849 249 4884
rect 71 4815 105 4849
rect 105 4815 139 4849
rect 139 4815 173 4849
rect 173 4815 207 4849
rect 207 4815 241 4849
rect 241 4815 249 4849
rect 71 4780 249 4815
rect 71 4746 105 4780
rect 105 4746 139 4780
rect 139 4746 173 4780
rect 173 4746 207 4780
rect 207 4746 241 4780
rect 241 4746 249 4780
rect 71 4711 249 4746
rect 71 4677 105 4711
rect 105 4677 139 4711
rect 139 4677 173 4711
rect 173 4677 207 4711
rect 207 4677 241 4711
rect 241 4677 249 4711
rect 71 4642 249 4677
rect 71 4608 105 4642
rect 105 4608 139 4642
rect 139 4608 173 4642
rect 173 4608 207 4642
rect 207 4608 241 4642
rect 241 4608 249 4642
rect 71 4573 249 4608
rect 71 4539 105 4573
rect 105 4539 139 4573
rect 139 4539 173 4573
rect 173 4539 207 4573
rect 207 4539 241 4573
rect 241 4539 249 4573
rect 71 4504 249 4539
rect 71 4470 105 4504
rect 105 4470 139 4504
rect 139 4470 173 4504
rect 173 4470 207 4504
rect 207 4470 241 4504
rect 241 4470 249 4504
rect 71 4435 249 4470
rect 71 4401 105 4435
rect 105 4401 139 4435
rect 139 4401 173 4435
rect 173 4401 207 4435
rect 207 4401 241 4435
rect 241 4401 249 4435
rect 71 4366 249 4401
rect 71 4332 105 4366
rect 105 4332 139 4366
rect 139 4332 173 4366
rect 173 4332 207 4366
rect 207 4332 241 4366
rect 241 4332 249 4366
rect 71 4297 249 4332
rect 71 4263 105 4297
rect 105 4263 139 4297
rect 139 4263 173 4297
rect 173 4263 207 4297
rect 207 4263 241 4297
rect 241 4263 249 4297
rect 71 4228 249 4263
rect 71 4194 105 4228
rect 105 4194 139 4228
rect 139 4194 173 4228
rect 173 4194 207 4228
rect 207 4194 241 4228
rect 241 4194 249 4228
rect 71 4159 249 4194
rect 71 4125 105 4159
rect 105 4125 139 4159
rect 139 4125 173 4159
rect 173 4125 207 4159
rect 207 4125 241 4159
rect 241 4125 249 4159
rect 71 4090 249 4125
rect 71 4056 105 4090
rect 105 4056 139 4090
rect 139 4056 173 4090
rect 173 4056 207 4090
rect 207 4056 241 4090
rect 241 4056 249 4090
rect 71 4021 249 4056
rect 71 3987 105 4021
rect 105 3987 139 4021
rect 139 3987 173 4021
rect 173 3987 207 4021
rect 207 3987 241 4021
rect 241 3987 249 4021
rect 71 3952 249 3987
rect 71 3918 105 3952
rect 105 3918 139 3952
rect 139 3918 173 3952
rect 173 3918 207 3952
rect 207 3918 241 3952
rect 241 3918 249 3952
rect 71 3883 249 3918
rect 71 3849 105 3883
rect 105 3849 139 3883
rect 139 3849 173 3883
rect 173 3849 207 3883
rect 207 3849 241 3883
rect 241 3849 249 3883
rect 71 3814 249 3849
rect 71 3780 105 3814
rect 105 3780 139 3814
rect 139 3780 173 3814
rect 173 3780 207 3814
rect 207 3780 241 3814
rect 241 3780 249 3814
rect 71 3745 249 3780
rect 71 3711 105 3745
rect 105 3711 139 3745
rect 139 3711 173 3745
rect 173 3711 207 3745
rect 207 3711 241 3745
rect 241 3711 249 3745
rect 71 3676 249 3711
rect 71 3642 105 3676
rect 105 3642 139 3676
rect 139 3642 173 3676
rect 173 3642 207 3676
rect 207 3642 241 3676
rect 241 3642 249 3676
rect 71 3607 249 3642
rect 71 3573 105 3607
rect 105 3573 139 3607
rect 139 3573 173 3607
rect 173 3573 207 3607
rect 207 3573 241 3607
rect 241 3573 249 3607
rect 71 3538 249 3573
rect 71 3504 105 3538
rect 105 3504 139 3538
rect 139 3504 173 3538
rect 173 3504 207 3538
rect 207 3504 241 3538
rect 241 3504 249 3538
rect 71 3469 249 3504
rect 71 3435 105 3469
rect 105 3435 139 3469
rect 139 3435 173 3469
rect 173 3435 207 3469
rect 207 3435 241 3469
rect 241 3435 249 3469
rect 71 3400 249 3435
rect 71 3366 105 3400
rect 105 3366 139 3400
rect 139 3366 173 3400
rect 173 3366 207 3400
rect 207 3366 241 3400
rect 241 3366 249 3400
rect 71 3331 249 3366
rect 71 3297 105 3331
rect 105 3297 139 3331
rect 139 3297 173 3331
rect 173 3297 207 3331
rect 207 3297 241 3331
rect 241 3297 249 3331
rect 71 3262 249 3297
rect 71 3228 105 3262
rect 105 3228 139 3262
rect 139 3228 173 3262
rect 173 3228 207 3262
rect 207 3228 241 3262
rect 241 3228 249 3262
rect 71 3193 249 3228
rect 71 3159 105 3193
rect 105 3159 139 3193
rect 139 3159 173 3193
rect 173 3159 207 3193
rect 207 3159 241 3193
rect 241 3159 249 3193
rect 71 3124 249 3159
rect 71 3090 105 3124
rect 105 3090 139 3124
rect 139 3090 173 3124
rect 173 3090 207 3124
rect 207 3090 241 3124
rect 241 3090 249 3124
rect 71 3055 249 3090
rect 71 3021 105 3055
rect 105 3021 139 3055
rect 139 3021 173 3055
rect 173 3021 207 3055
rect 207 3021 241 3055
rect 241 3021 249 3055
rect 71 2986 249 3021
rect 71 2952 105 2986
rect 105 2952 139 2986
rect 139 2952 173 2986
rect 173 2952 207 2986
rect 207 2952 241 2986
rect 241 2952 249 2986
rect 71 2917 249 2952
rect 71 2883 105 2917
rect 105 2883 139 2917
rect 139 2883 173 2917
rect 173 2883 207 2917
rect 207 2883 241 2917
rect 241 2883 249 2917
rect 71 2848 249 2883
rect 71 2814 105 2848
rect 105 2814 139 2848
rect 139 2814 173 2848
rect 173 2814 207 2848
rect 207 2814 241 2848
rect 241 2814 249 2848
rect 71 2779 249 2814
rect 71 2745 105 2779
rect 105 2745 139 2779
rect 139 2745 173 2779
rect 173 2745 207 2779
rect 207 2745 241 2779
rect 241 2745 249 2779
rect 71 2710 249 2745
rect 71 2676 105 2710
rect 105 2676 139 2710
rect 139 2676 173 2710
rect 173 2676 207 2710
rect 207 2676 241 2710
rect 241 2676 249 2710
rect 71 2641 249 2676
rect 71 2607 105 2641
rect 105 2607 139 2641
rect 139 2607 173 2641
rect 173 2607 207 2641
rect 207 2607 241 2641
rect 241 2607 249 2641
rect 71 2572 249 2607
rect 71 2538 105 2572
rect 105 2538 139 2572
rect 139 2538 173 2572
rect 173 2538 207 2572
rect 207 2538 241 2572
rect 241 2538 249 2572
rect 71 2503 249 2538
rect 71 2469 105 2503
rect 105 2469 139 2503
rect 139 2469 173 2503
rect 173 2469 207 2503
rect 207 2469 241 2503
rect 241 2469 249 2503
rect 71 2434 249 2469
rect 71 2400 105 2434
rect 105 2400 139 2434
rect 139 2400 173 2434
rect 173 2400 207 2434
rect 207 2400 241 2434
rect 241 2400 249 2434
rect 71 2365 249 2400
rect 71 2331 105 2365
rect 105 2331 139 2365
rect 139 2331 173 2365
rect 173 2331 207 2365
rect 207 2331 241 2365
rect 241 2331 249 2365
rect 71 2296 249 2331
rect 71 2262 105 2296
rect 105 2262 139 2296
rect 139 2262 173 2296
rect 173 2262 207 2296
rect 207 2262 241 2296
rect 241 2262 249 2296
rect 71 2227 249 2262
rect 71 2193 105 2227
rect 105 2193 139 2227
rect 139 2193 173 2227
rect 173 2193 207 2227
rect 207 2193 241 2227
rect 241 2193 249 2227
rect 71 2158 249 2193
rect 71 2124 105 2158
rect 105 2124 139 2158
rect 139 2124 173 2158
rect 173 2124 207 2158
rect 207 2124 241 2158
rect 241 2124 249 2158
rect 71 2089 249 2124
rect 71 2055 105 2089
rect 105 2055 139 2089
rect 139 2055 173 2089
rect 173 2055 207 2089
rect 207 2055 241 2089
rect 241 2055 249 2089
rect 71 2020 249 2055
rect 71 1986 105 2020
rect 105 1986 139 2020
rect 139 1986 173 2020
rect 173 1986 207 2020
rect 207 1986 241 2020
rect 241 1986 249 2020
rect 71 1951 249 1986
rect 71 1917 105 1951
rect 105 1917 139 1951
rect 139 1917 173 1951
rect 173 1917 207 1951
rect 207 1917 241 1951
rect 241 1917 249 1951
rect 71 1882 249 1917
rect 71 1848 105 1882
rect 105 1848 139 1882
rect 139 1848 173 1882
rect 173 1848 207 1882
rect 207 1848 241 1882
rect 241 1848 249 1882
rect 71 1813 249 1848
rect 71 1779 105 1813
rect 105 1779 139 1813
rect 139 1779 173 1813
rect 173 1779 207 1813
rect 207 1779 241 1813
rect 241 1779 249 1813
rect 71 1744 249 1779
rect 71 1710 105 1744
rect 105 1710 139 1744
rect 139 1710 173 1744
rect 173 1710 207 1744
rect 207 1710 241 1744
rect 241 1710 249 1744
rect 71 1675 249 1710
rect 71 1641 105 1675
rect 105 1641 139 1675
rect 139 1641 173 1675
rect 173 1641 207 1675
rect 207 1641 241 1675
rect 241 1641 249 1675
rect 71 1606 249 1641
rect 71 1572 105 1606
rect 105 1572 139 1606
rect 139 1572 173 1606
rect 173 1572 207 1606
rect 207 1572 241 1606
rect 241 1572 249 1606
rect 71 1537 249 1572
rect 71 1503 105 1537
rect 105 1503 139 1537
rect 139 1503 173 1537
rect 173 1503 207 1537
rect 207 1503 241 1537
rect 241 1503 249 1537
rect 71 1468 249 1503
rect 71 1434 105 1468
rect 105 1434 139 1468
rect 139 1434 173 1468
rect 173 1434 207 1468
rect 207 1434 241 1468
rect 241 1434 249 1468
rect 71 1399 249 1434
rect 71 1365 105 1399
rect 105 1365 139 1399
rect 139 1365 173 1399
rect 173 1365 207 1399
rect 207 1365 241 1399
rect 241 1365 249 1399
rect 71 1330 249 1365
rect 71 1296 105 1330
rect 105 1296 139 1330
rect 139 1296 173 1330
rect 173 1296 207 1330
rect 207 1296 241 1330
rect 241 1296 249 1330
rect 71 1261 249 1296
rect 71 1227 105 1261
rect 105 1227 139 1261
rect 139 1227 173 1261
rect 173 1227 207 1261
rect 207 1227 241 1261
rect 241 1227 249 1261
rect 71 1192 249 1227
rect 71 1158 105 1192
rect 105 1158 139 1192
rect 139 1158 173 1192
rect 173 1158 207 1192
rect 207 1158 241 1192
rect 241 1158 249 1192
rect 71 1123 249 1158
rect 71 545 241 1123
rect 241 545 249 1123
rect 767 4818 12465 4924
rect 12504 4890 12538 4924
rect 12577 4890 12611 4924
rect 12650 4890 12684 4924
rect 12723 4890 12757 4924
rect 12796 4890 12830 4924
rect 12869 4890 12903 4924
rect 12942 4890 12976 4924
rect 13015 4890 13049 4924
rect 13088 4890 13122 4924
rect 13161 4890 13195 4924
rect 13234 4890 13268 4924
rect 13307 4890 13341 4924
rect 13380 4890 13414 4924
rect 13453 4890 13487 4924
rect 13526 4890 13560 4924
rect 13599 4890 13633 4924
rect 13672 4890 13706 4924
rect 13745 4890 13779 4924
rect 13818 4890 13852 4924
rect 13891 4890 13925 4924
rect 13964 4890 13998 4924
rect 14037 4890 14071 4924
rect 14110 4890 14144 4924
rect 14183 4890 14217 4924
rect 14256 4890 14290 4924
rect 14329 4890 14363 4924
rect 14402 4890 14436 4924
rect 12504 4818 12538 4852
rect 12577 4818 12611 4852
rect 12650 4818 12684 4852
rect 12723 4818 12757 4852
rect 12796 4818 12830 4852
rect 12869 4818 12903 4852
rect 12942 4818 12976 4852
rect 13015 4818 13049 4852
rect 13088 4818 13122 4852
rect 13161 4818 13195 4852
rect 13234 4818 13268 4852
rect 13307 4818 13341 4852
rect 13380 4818 13414 4852
rect 13453 4818 13487 4852
rect 13526 4818 13560 4852
rect 13599 4818 13633 4852
rect 13672 4818 13706 4852
rect 13745 4818 13779 4852
rect 13818 4818 13852 4852
rect 13891 4818 13925 4852
rect 13964 4818 13998 4852
rect 14037 4818 14071 4852
rect 14110 4818 14144 4852
rect 14183 4818 14217 4852
rect 14256 4818 14290 4852
rect 14329 4818 14363 4852
rect 14402 4820 14436 4852
rect 14402 4818 14428 4820
rect 14428 4818 14436 4820
rect 587 4710 621 4744
rect 659 4717 691 4744
rect 691 4717 693 4744
rect 733 4740 767 4774
rect 659 4710 693 4717
rect 587 4636 621 4670
rect 659 4648 691 4670
rect 691 4648 693 4670
rect 733 4667 767 4701
rect 659 4636 693 4648
rect 587 4563 621 4596
rect 587 4562 589 4563
rect 589 4562 621 4563
rect 659 4562 693 4596
rect 733 4594 767 4628
rect 587 4492 621 4522
rect 587 4488 589 4492
rect 589 4488 621 4492
rect 659 4488 693 4522
rect 733 4521 767 4555
rect 14431 4740 14465 4774
rect 14510 4716 14531 4743
rect 14531 4716 14544 4743
rect 14510 4709 14544 4716
rect 14582 4714 14599 4743
rect 14599 4714 14616 4743
rect 14582 4709 14616 4714
rect 14431 4667 14465 4701
rect 14510 4646 14531 4670
rect 14531 4646 14544 4670
rect 14510 4636 14544 4646
rect 14582 4644 14599 4670
rect 14599 4644 14616 4670
rect 14582 4636 14616 4644
rect 14431 4594 14465 4628
rect 14510 4576 14531 4597
rect 14531 4576 14544 4597
rect 14510 4563 14544 4576
rect 14582 4574 14599 4597
rect 14599 4574 14616 4597
rect 14582 4563 14616 4574
rect 14431 4521 14465 4555
rect 14510 4506 14531 4524
rect 14531 4506 14544 4524
rect 587 4421 621 4449
rect 587 4415 589 4421
rect 589 4415 621 4421
rect 659 4415 693 4449
rect 733 4448 767 4482
rect 587 4350 621 4376
rect 587 4342 589 4350
rect 589 4342 621 4350
rect 659 4342 693 4376
rect 733 4375 767 4409
rect 587 4279 621 4303
rect 587 4269 589 4279
rect 589 4269 621 4279
rect 659 4269 693 4303
rect 733 4302 767 4336
rect 587 4208 621 4230
rect 587 4196 589 4208
rect 589 4196 621 4208
rect 659 4196 693 4230
rect 733 4229 767 4263
rect 587 4137 621 4157
rect 587 4123 589 4137
rect 589 4123 621 4137
rect 659 4123 693 4157
rect 733 4156 767 4190
rect 587 4050 621 4084
rect 659 4050 693 4084
rect 733 4083 767 4117
rect 931 4388 1037 4494
rect 587 4007 589 4011
rect 589 4007 621 4011
rect 733 4034 767 4044
rect 587 3977 621 4007
rect 659 3977 693 4011
rect 733 4010 734 4034
rect 734 4010 767 4034
rect 587 3936 589 3938
rect 589 3936 621 3938
rect 733 3966 767 3971
rect 587 3904 621 3936
rect 659 3904 693 3938
rect 733 3937 734 3966
rect 734 3937 767 3966
rect 587 3862 589 3865
rect 589 3862 621 3865
rect 587 3831 621 3862
rect 659 3831 693 3865
rect 733 3864 734 3898
rect 734 3864 767 3898
rect 587 3791 589 3792
rect 589 3791 621 3792
rect 733 3796 734 3825
rect 734 3796 767 3825
rect 587 3758 621 3791
rect 659 3758 693 3792
rect 733 3791 767 3796
rect 587 3717 589 3719
rect 589 3717 621 3719
rect 733 3728 734 3752
rect 734 3728 767 3752
rect 587 3685 621 3717
rect 659 3685 693 3719
rect 733 3718 767 3728
rect 733 3660 734 3679
rect 734 3660 767 3679
rect 587 3612 621 3646
rect 659 3612 693 3646
rect 733 3645 767 3660
rect 587 3572 589 3573
rect 589 3572 621 3573
rect 733 3592 734 3606
rect 734 3592 767 3606
rect 587 3539 621 3572
rect 659 3539 693 3573
rect 733 3572 767 3592
rect 733 3524 734 3533
rect 734 3524 767 3533
rect 587 3466 621 3500
rect 659 3466 693 3500
rect 733 3499 767 3524
rect 733 3456 734 3460
rect 734 3456 767 3460
rect 587 3393 621 3427
rect 659 3393 693 3427
rect 733 3426 767 3456
rect 733 3354 767 3387
rect 587 3320 621 3354
rect 659 3320 693 3354
rect 733 3353 734 3354
rect 734 3353 767 3354
rect 733 3286 767 3314
rect 587 3247 621 3281
rect 659 3247 693 3281
rect 733 3280 734 3286
rect 734 3280 767 3286
rect 733 3218 767 3241
rect 587 3174 621 3208
rect 659 3174 693 3208
rect 733 3207 734 3218
rect 734 3207 767 3218
rect 587 3117 589 3135
rect 589 3117 621 3135
rect 733 3150 767 3168
rect 587 3101 621 3117
rect 659 3101 693 3135
rect 733 3134 734 3150
rect 734 3134 767 3150
rect 587 3028 621 3062
rect 659 3028 693 3062
rect 733 3061 767 3095
rect 587 2955 621 2989
rect 659 2955 693 2989
rect 733 2988 767 3022
rect 587 2882 621 2916
rect 659 2882 693 2916
rect 733 2915 767 2949
rect 587 2809 621 2843
rect 659 2809 693 2843
rect 733 2842 767 2876
rect 587 2736 621 2770
rect 659 2736 693 2770
rect 733 2769 767 2803
rect 587 2663 621 2697
rect 659 2663 693 2697
rect 733 2696 767 2730
rect 587 2590 621 2624
rect 659 2590 693 2624
rect 733 2623 767 2657
rect 587 2517 621 2551
rect 659 2517 693 2551
rect 733 2550 767 2584
rect 587 2444 621 2478
rect 659 2444 693 2478
rect 733 2477 767 2511
rect 1361 4388 1467 4494
rect 733 2433 767 2438
rect 587 2371 621 2405
rect 659 2371 693 2405
rect 733 2404 734 2433
rect 734 2404 767 2433
rect 587 2327 621 2332
rect 587 2298 589 2327
rect 589 2298 621 2327
rect 659 2298 693 2332
rect 733 2331 734 2365
rect 734 2331 767 2365
rect 733 2263 734 2292
rect 734 2263 767 2292
rect 587 2250 621 2259
rect 587 2225 589 2250
rect 589 2225 621 2250
rect 659 2225 693 2259
rect 733 2258 767 2263
rect 733 2195 734 2219
rect 734 2195 767 2219
rect 587 2156 621 2186
rect 587 2152 589 2156
rect 589 2152 621 2156
rect 659 2152 693 2186
rect 733 2185 767 2195
rect 733 2127 734 2146
rect 734 2127 767 2146
rect 587 2085 621 2113
rect 587 2079 589 2085
rect 589 2079 621 2085
rect 659 2079 693 2113
rect 733 2112 767 2127
rect 733 2059 734 2073
rect 734 2059 767 2073
rect 587 2011 621 2040
rect 587 2006 589 2011
rect 589 2006 621 2011
rect 659 2006 693 2040
rect 733 2039 767 2059
rect 733 1991 734 2000
rect 734 1991 767 2000
rect 587 1940 621 1967
rect 587 1933 589 1940
rect 589 1933 621 1940
rect 659 1933 693 1967
rect 733 1966 767 1991
rect 733 1923 734 1927
rect 734 1923 767 1927
rect 587 1866 621 1894
rect 587 1860 589 1866
rect 589 1860 621 1866
rect 659 1860 693 1894
rect 733 1893 767 1923
rect 733 1821 767 1854
rect 587 1795 621 1821
rect 587 1787 589 1795
rect 589 1787 621 1795
rect 659 1787 693 1821
rect 733 1820 734 1821
rect 734 1820 767 1821
rect 733 1753 767 1781
rect 587 1721 621 1748
rect 587 1714 589 1721
rect 589 1714 621 1721
rect 659 1714 693 1748
rect 733 1747 734 1753
rect 734 1747 767 1753
rect 733 1685 767 1708
rect 587 1650 621 1675
rect 587 1641 589 1650
rect 589 1641 621 1650
rect 659 1641 693 1675
rect 733 1674 734 1685
rect 734 1674 767 1685
rect 733 1617 767 1635
rect 587 1576 621 1602
rect 587 1568 589 1576
rect 589 1568 621 1576
rect 659 1568 693 1602
rect 733 1601 734 1617
rect 734 1601 767 1617
rect 733 1549 767 1562
rect 587 1505 621 1529
rect 587 1495 589 1505
rect 589 1495 621 1505
rect 659 1495 693 1529
rect 733 1528 734 1549
rect 734 1528 767 1549
rect 733 1455 767 1489
rect 587 1385 621 1419
rect 659 1385 693 1419
rect 733 1382 767 1416
rect 587 1296 621 1330
rect 659 1296 693 1330
rect 733 1308 767 1342
rect 1110 4028 1144 4062
rect 1182 4028 1216 4062
rect 1254 4028 1288 4062
rect 1110 3954 1144 3988
rect 1182 3954 1216 3988
rect 1254 3954 1288 3988
rect 1110 3880 1144 3914
rect 1182 3880 1216 3914
rect 1254 3880 1288 3914
rect 1110 3806 1144 3840
rect 1182 3806 1216 3840
rect 1254 3806 1288 3840
rect 1110 3732 1144 3766
rect 1182 3732 1216 3766
rect 1254 3732 1288 3766
rect 1110 3658 1144 3692
rect 1182 3658 1216 3692
rect 1254 3658 1288 3692
rect 1110 3584 1144 3618
rect 1182 3584 1216 3618
rect 1254 3584 1288 3618
rect 1110 3510 1144 3544
rect 1182 3510 1216 3544
rect 1254 3510 1288 3544
rect 1110 3436 1144 3470
rect 1182 3436 1216 3470
rect 1254 3436 1288 3470
rect 1110 3362 1144 3396
rect 1182 3362 1216 3396
rect 1254 3362 1288 3396
rect 1110 3288 1144 3322
rect 1182 3288 1216 3322
rect 1254 3288 1288 3322
rect 1110 3214 1144 3248
rect 1182 3214 1216 3248
rect 1254 3214 1288 3248
rect 1110 3140 1144 3174
rect 1182 3140 1216 3174
rect 1254 3140 1288 3174
rect 1110 3066 1144 3100
rect 1182 3066 1216 3100
rect 1254 3066 1288 3100
rect 1110 2992 1144 3026
rect 1182 2992 1216 3026
rect 1254 2992 1288 3026
rect 1110 2918 1144 2952
rect 1182 2918 1216 2952
rect 1254 2918 1288 2952
rect 1110 2844 1144 2878
rect 1182 2844 1216 2878
rect 1254 2844 1288 2878
rect 1110 2770 1144 2804
rect 1182 2770 1216 2804
rect 1254 2770 1288 2804
rect 1110 2696 1144 2730
rect 1182 2696 1216 2730
rect 1254 2696 1288 2730
rect 1110 2622 1144 2656
rect 1182 2622 1216 2656
rect 1254 2622 1288 2656
rect 1110 2548 1144 2582
rect 1182 2548 1216 2582
rect 1254 2548 1288 2582
rect 1110 2474 1144 2508
rect 1182 2474 1216 2508
rect 1254 2474 1288 2508
rect 1110 2400 1144 2434
rect 1182 2400 1216 2434
rect 1254 2400 1288 2434
rect 1110 2326 1144 2360
rect 1182 2326 1216 2360
rect 1254 2326 1288 2360
rect 1110 2252 1144 2286
rect 1182 2252 1216 2286
rect 1254 2252 1288 2286
rect 1110 2178 1144 2212
rect 1182 2178 1216 2212
rect 1254 2178 1288 2212
rect 1110 2104 1144 2138
rect 1182 2104 1216 2138
rect 1254 2104 1288 2138
rect 1110 2030 1144 2064
rect 1182 2030 1216 2064
rect 1254 2030 1288 2064
rect 1110 1956 1144 1990
rect 1182 1956 1216 1990
rect 1254 1956 1288 1990
rect 1110 1882 1144 1916
rect 1182 1882 1216 1916
rect 1254 1882 1288 1916
rect 1110 1808 1144 1842
rect 1182 1808 1216 1842
rect 1254 1808 1288 1842
rect 1110 1734 1144 1768
rect 1182 1734 1216 1768
rect 1254 1734 1288 1768
rect 1110 1660 1144 1694
rect 1182 1660 1216 1694
rect 1254 1660 1288 1694
rect 1110 1586 1144 1620
rect 1182 1586 1216 1620
rect 1254 1586 1288 1620
rect 1110 1511 1144 1545
rect 1182 1511 1216 1545
rect 1254 1511 1288 1545
rect 1923 4388 2029 4494
rect 1678 4050 1712 4062
rect 1606 4046 1784 4050
rect 1606 4012 1610 4046
rect 1610 4012 1678 4046
rect 1678 4012 1712 4046
rect 1712 4012 1780 4046
rect 1780 4012 1784 4046
rect 1606 3978 1784 4012
rect 1606 3944 1610 3978
rect 1610 3944 1678 3978
rect 1678 3944 1712 3978
rect 1712 3944 1780 3978
rect 1780 3944 1784 3978
rect 1606 3910 1784 3944
rect 1606 3876 1610 3910
rect 1610 3876 1678 3910
rect 1678 3876 1712 3910
rect 1712 3876 1780 3910
rect 1780 3876 1784 3910
rect 1606 3842 1784 3876
rect 1606 3808 1610 3842
rect 1610 3808 1678 3842
rect 1678 3808 1712 3842
rect 1712 3808 1780 3842
rect 1780 3808 1784 3842
rect 1606 3774 1784 3808
rect 1606 3740 1610 3774
rect 1610 3740 1678 3774
rect 1678 3740 1712 3774
rect 1712 3740 1780 3774
rect 1780 3740 1784 3774
rect 1606 3706 1784 3740
rect 1606 3672 1610 3706
rect 1610 3672 1678 3706
rect 1678 3672 1712 3706
rect 1712 3672 1780 3706
rect 1780 3672 1784 3706
rect 1606 3638 1784 3672
rect 1606 3604 1610 3638
rect 1610 3604 1678 3638
rect 1678 3604 1712 3638
rect 1712 3604 1780 3638
rect 1780 3604 1784 3638
rect 1606 3570 1784 3604
rect 1606 3536 1610 3570
rect 1610 3536 1678 3570
rect 1678 3536 1712 3570
rect 1712 3536 1780 3570
rect 1780 3536 1784 3570
rect 1606 3502 1784 3536
rect 1606 3468 1610 3502
rect 1610 3468 1678 3502
rect 1678 3468 1712 3502
rect 1712 3468 1780 3502
rect 1780 3468 1784 3502
rect 1606 3434 1784 3468
rect 1606 3400 1610 3434
rect 1610 3400 1678 3434
rect 1678 3400 1712 3434
rect 1712 3400 1780 3434
rect 1780 3400 1784 3434
rect 1606 3366 1784 3400
rect 1606 3332 1610 3366
rect 1610 3332 1678 3366
rect 1678 3332 1712 3366
rect 1712 3332 1780 3366
rect 1780 3332 1784 3366
rect 1606 3298 1784 3332
rect 1606 3264 1610 3298
rect 1610 3264 1678 3298
rect 1678 3264 1712 3298
rect 1712 3264 1780 3298
rect 1780 3264 1784 3298
rect 1606 3230 1784 3264
rect 1606 3196 1610 3230
rect 1610 3196 1678 3230
rect 1678 3196 1712 3230
rect 1712 3196 1780 3230
rect 1780 3196 1784 3230
rect 1606 3162 1784 3196
rect 1606 3128 1610 3162
rect 1610 3128 1678 3162
rect 1678 3128 1712 3162
rect 1712 3128 1780 3162
rect 1780 3128 1784 3162
rect 1606 3092 1784 3128
rect 1606 3080 1640 3092
rect 1750 3080 1784 3092
rect 1606 2935 1784 3040
rect 1606 2901 1645 2935
rect 1645 2901 1679 2935
rect 1679 2901 1713 2935
rect 1713 2901 1747 2935
rect 1747 2901 1784 2935
rect 1606 2855 1784 2901
rect 1606 2821 1645 2855
rect 1645 2821 1679 2855
rect 1679 2821 1713 2855
rect 1713 2821 1747 2855
rect 1747 2821 1784 2855
rect 1606 2775 1784 2821
rect 1606 2741 1645 2775
rect 1645 2741 1679 2775
rect 1679 2741 1713 2775
rect 1713 2741 1747 2775
rect 1747 2741 1784 2775
rect 1606 2695 1784 2741
rect 1606 2661 1645 2695
rect 1645 2661 1679 2695
rect 1679 2661 1713 2695
rect 1713 2661 1747 2695
rect 1747 2661 1784 2695
rect 1606 2614 1784 2661
rect 1606 2580 1645 2614
rect 1645 2580 1679 2614
rect 1679 2580 1713 2614
rect 1713 2580 1747 2614
rect 1747 2580 1784 2614
rect 1606 2574 1784 2580
rect 1606 2501 1640 2535
rect 1678 2501 1712 2535
rect 1750 2501 1784 2535
rect 1678 2449 1712 2461
rect 1606 2445 1784 2449
rect 1606 2411 1610 2445
rect 1610 2411 1678 2445
rect 1678 2411 1712 2445
rect 1712 2411 1780 2445
rect 1780 2411 1784 2445
rect 1606 2377 1784 2411
rect 1606 2343 1610 2377
rect 1610 2343 1678 2377
rect 1678 2343 1712 2377
rect 1712 2343 1780 2377
rect 1780 2343 1784 2377
rect 1606 2309 1784 2343
rect 1606 2275 1610 2309
rect 1610 2275 1678 2309
rect 1678 2275 1712 2309
rect 1712 2275 1780 2309
rect 1780 2275 1784 2309
rect 1606 2241 1784 2275
rect 1606 2207 1610 2241
rect 1610 2207 1678 2241
rect 1678 2207 1712 2241
rect 1712 2207 1780 2241
rect 1780 2207 1784 2241
rect 1606 2173 1784 2207
rect 1606 2139 1610 2173
rect 1610 2139 1678 2173
rect 1678 2139 1712 2173
rect 1712 2139 1780 2173
rect 1780 2139 1784 2173
rect 1606 2105 1784 2139
rect 1606 2071 1610 2105
rect 1610 2071 1678 2105
rect 1678 2071 1712 2105
rect 1712 2071 1780 2105
rect 1780 2071 1784 2105
rect 1606 2037 1784 2071
rect 1606 2003 1610 2037
rect 1610 2003 1678 2037
rect 1678 2003 1712 2037
rect 1712 2003 1780 2037
rect 1780 2003 1784 2037
rect 1606 1969 1784 2003
rect 1606 1935 1610 1969
rect 1610 1935 1678 1969
rect 1678 1935 1712 1969
rect 1712 1935 1780 1969
rect 1780 1935 1784 1969
rect 1606 1901 1784 1935
rect 1606 1867 1610 1901
rect 1610 1867 1678 1901
rect 1678 1867 1712 1901
rect 1712 1867 1780 1901
rect 1780 1867 1784 1901
rect 1606 1833 1784 1867
rect 1606 1799 1610 1833
rect 1610 1799 1678 1833
rect 1678 1799 1712 1833
rect 1712 1799 1780 1833
rect 1780 1799 1784 1833
rect 1606 1765 1784 1799
rect 1606 1731 1610 1765
rect 1610 1731 1678 1765
rect 1678 1731 1712 1765
rect 1712 1731 1780 1765
rect 1780 1731 1784 1765
rect 1606 1697 1784 1731
rect 1606 1663 1610 1697
rect 1610 1663 1678 1697
rect 1678 1663 1712 1697
rect 1712 1663 1780 1697
rect 1780 1663 1784 1697
rect 1606 1629 1784 1663
rect 1606 1595 1610 1629
rect 1610 1595 1678 1629
rect 1678 1595 1712 1629
rect 1712 1595 1780 1629
rect 1780 1595 1784 1629
rect 1606 1561 1784 1595
rect 1606 1527 1610 1561
rect 1610 1527 1678 1561
rect 1678 1527 1712 1561
rect 1712 1527 1780 1561
rect 1780 1527 1784 1561
rect 1606 1491 1784 1527
rect 1606 1479 1640 1491
rect 1750 1479 1784 1491
rect 2353 4388 2459 4494
rect 2102 4028 2136 4062
rect 2174 4028 2208 4062
rect 2246 4028 2280 4062
rect 2102 3954 2136 3988
rect 2174 3954 2208 3988
rect 2246 3954 2280 3988
rect 2102 3880 2136 3914
rect 2174 3880 2208 3914
rect 2246 3880 2280 3914
rect 2102 3806 2136 3840
rect 2174 3806 2208 3840
rect 2246 3806 2280 3840
rect 2102 3732 2136 3766
rect 2174 3732 2208 3766
rect 2246 3732 2280 3766
rect 2102 3658 2136 3692
rect 2174 3658 2208 3692
rect 2246 3658 2280 3692
rect 2102 3584 2136 3618
rect 2174 3584 2208 3618
rect 2246 3584 2280 3618
rect 2102 3510 2136 3544
rect 2174 3510 2208 3544
rect 2246 3510 2280 3544
rect 2102 3436 2136 3470
rect 2174 3436 2208 3470
rect 2246 3436 2280 3470
rect 2102 3362 2136 3396
rect 2174 3362 2208 3396
rect 2246 3362 2280 3396
rect 2102 3288 2136 3322
rect 2174 3288 2208 3322
rect 2246 3288 2280 3322
rect 2102 3214 2136 3248
rect 2174 3214 2208 3248
rect 2246 3214 2280 3248
rect 2102 3140 2136 3174
rect 2174 3140 2208 3174
rect 2246 3140 2280 3174
rect 2102 3066 2136 3100
rect 2174 3066 2208 3100
rect 2246 3066 2280 3100
rect 2102 2992 2136 3026
rect 2174 2992 2208 3026
rect 2246 2992 2280 3026
rect 2102 2918 2136 2952
rect 2174 2918 2208 2952
rect 2246 2918 2280 2952
rect 2102 2844 2136 2878
rect 2174 2844 2208 2878
rect 2246 2844 2280 2878
rect 2102 2770 2136 2804
rect 2174 2770 2208 2804
rect 2246 2770 2280 2804
rect 2102 2696 2136 2730
rect 2174 2696 2208 2730
rect 2246 2696 2280 2730
rect 2102 2622 2136 2656
rect 2174 2622 2208 2656
rect 2246 2622 2280 2656
rect 2102 2548 2136 2582
rect 2174 2548 2208 2582
rect 2246 2548 2280 2582
rect 2102 2474 2136 2508
rect 2174 2474 2208 2508
rect 2246 2474 2280 2508
rect 2102 2400 2136 2434
rect 2174 2400 2208 2434
rect 2246 2400 2280 2434
rect 2102 2326 2136 2360
rect 2174 2326 2208 2360
rect 2246 2326 2280 2360
rect 2102 2252 2136 2286
rect 2174 2252 2208 2286
rect 2246 2252 2280 2286
rect 2102 2178 2136 2212
rect 2174 2178 2208 2212
rect 2246 2178 2280 2212
rect 2102 2104 2136 2138
rect 2174 2104 2208 2138
rect 2246 2104 2280 2138
rect 2102 2030 2136 2064
rect 2174 2030 2208 2064
rect 2246 2030 2280 2064
rect 2102 1956 2136 1990
rect 2174 1956 2208 1990
rect 2246 1956 2280 1990
rect 2102 1882 2136 1916
rect 2174 1882 2208 1916
rect 2246 1882 2280 1916
rect 2102 1808 2136 1842
rect 2174 1808 2208 1842
rect 2246 1808 2280 1842
rect 2102 1734 2136 1768
rect 2174 1734 2208 1768
rect 2246 1734 2280 1768
rect 2102 1660 2136 1694
rect 2174 1660 2208 1694
rect 2246 1660 2280 1694
rect 2102 1586 2136 1620
rect 2174 1586 2208 1620
rect 2246 1586 2280 1620
rect 2102 1511 2136 1545
rect 2174 1511 2208 1545
rect 2246 1511 2280 1545
rect 2915 4388 3021 4494
rect 2670 4050 2704 4062
rect 2598 4046 2776 4050
rect 2598 4012 2602 4046
rect 2602 4012 2670 4046
rect 2670 4012 2704 4046
rect 2704 4012 2772 4046
rect 2772 4012 2776 4046
rect 2598 3978 2776 4012
rect 2598 3944 2602 3978
rect 2602 3944 2670 3978
rect 2670 3944 2704 3978
rect 2704 3944 2772 3978
rect 2772 3944 2776 3978
rect 2598 3910 2776 3944
rect 2598 3876 2602 3910
rect 2602 3876 2670 3910
rect 2670 3876 2704 3910
rect 2704 3876 2772 3910
rect 2772 3876 2776 3910
rect 2598 3842 2776 3876
rect 2598 3808 2602 3842
rect 2602 3808 2670 3842
rect 2670 3808 2704 3842
rect 2704 3808 2772 3842
rect 2772 3808 2776 3842
rect 2598 3774 2776 3808
rect 2598 3740 2602 3774
rect 2602 3740 2670 3774
rect 2670 3740 2704 3774
rect 2704 3740 2772 3774
rect 2772 3740 2776 3774
rect 2598 3706 2776 3740
rect 2598 3672 2602 3706
rect 2602 3672 2670 3706
rect 2670 3672 2704 3706
rect 2704 3672 2772 3706
rect 2772 3672 2776 3706
rect 2598 3638 2776 3672
rect 2598 3604 2602 3638
rect 2602 3604 2670 3638
rect 2670 3604 2704 3638
rect 2704 3604 2772 3638
rect 2772 3604 2776 3638
rect 2598 3570 2776 3604
rect 2598 3536 2602 3570
rect 2602 3536 2670 3570
rect 2670 3536 2704 3570
rect 2704 3536 2772 3570
rect 2772 3536 2776 3570
rect 2598 3502 2776 3536
rect 2598 3468 2602 3502
rect 2602 3468 2670 3502
rect 2670 3468 2704 3502
rect 2704 3468 2772 3502
rect 2772 3468 2776 3502
rect 2598 3434 2776 3468
rect 2598 3400 2602 3434
rect 2602 3400 2670 3434
rect 2670 3400 2704 3434
rect 2704 3400 2772 3434
rect 2772 3400 2776 3434
rect 2598 3366 2776 3400
rect 2598 3332 2602 3366
rect 2602 3332 2670 3366
rect 2670 3332 2704 3366
rect 2704 3332 2772 3366
rect 2772 3332 2776 3366
rect 2598 3298 2776 3332
rect 2598 3264 2602 3298
rect 2602 3264 2670 3298
rect 2670 3264 2704 3298
rect 2704 3264 2772 3298
rect 2772 3264 2776 3298
rect 2598 3230 2776 3264
rect 2598 3196 2602 3230
rect 2602 3196 2670 3230
rect 2670 3196 2704 3230
rect 2704 3196 2772 3230
rect 2772 3196 2776 3230
rect 2598 3162 2776 3196
rect 2598 3128 2602 3162
rect 2602 3128 2670 3162
rect 2670 3128 2704 3162
rect 2704 3128 2772 3162
rect 2772 3128 2776 3162
rect 2598 3092 2776 3128
rect 2598 3080 2632 3092
rect 2742 3080 2776 3092
rect 2598 2935 2776 3040
rect 2598 2901 2637 2935
rect 2637 2901 2671 2935
rect 2671 2901 2705 2935
rect 2705 2901 2739 2935
rect 2739 2901 2776 2935
rect 2598 2855 2776 2901
rect 2598 2821 2637 2855
rect 2637 2821 2671 2855
rect 2671 2821 2705 2855
rect 2705 2821 2739 2855
rect 2739 2821 2776 2855
rect 2598 2775 2776 2821
rect 2598 2741 2637 2775
rect 2637 2741 2671 2775
rect 2671 2741 2705 2775
rect 2705 2741 2739 2775
rect 2739 2741 2776 2775
rect 2598 2695 2776 2741
rect 2598 2661 2637 2695
rect 2637 2661 2671 2695
rect 2671 2661 2705 2695
rect 2705 2661 2739 2695
rect 2739 2661 2776 2695
rect 2598 2614 2776 2661
rect 2598 2580 2637 2614
rect 2637 2580 2671 2614
rect 2671 2580 2705 2614
rect 2705 2580 2739 2614
rect 2739 2580 2776 2614
rect 2598 2574 2776 2580
rect 2598 2501 2632 2535
rect 2670 2501 2704 2535
rect 2742 2501 2776 2535
rect 2670 2449 2704 2461
rect 2598 2445 2776 2449
rect 2598 2411 2602 2445
rect 2602 2411 2670 2445
rect 2670 2411 2704 2445
rect 2704 2411 2772 2445
rect 2772 2411 2776 2445
rect 2598 2377 2776 2411
rect 2598 2343 2602 2377
rect 2602 2343 2670 2377
rect 2670 2343 2704 2377
rect 2704 2343 2772 2377
rect 2772 2343 2776 2377
rect 2598 2309 2776 2343
rect 2598 2275 2602 2309
rect 2602 2275 2670 2309
rect 2670 2275 2704 2309
rect 2704 2275 2772 2309
rect 2772 2275 2776 2309
rect 2598 2241 2776 2275
rect 2598 2207 2602 2241
rect 2602 2207 2670 2241
rect 2670 2207 2704 2241
rect 2704 2207 2772 2241
rect 2772 2207 2776 2241
rect 2598 2173 2776 2207
rect 2598 2139 2602 2173
rect 2602 2139 2670 2173
rect 2670 2139 2704 2173
rect 2704 2139 2772 2173
rect 2772 2139 2776 2173
rect 2598 2105 2776 2139
rect 2598 2071 2602 2105
rect 2602 2071 2670 2105
rect 2670 2071 2704 2105
rect 2704 2071 2772 2105
rect 2772 2071 2776 2105
rect 2598 2037 2776 2071
rect 2598 2003 2602 2037
rect 2602 2003 2670 2037
rect 2670 2003 2704 2037
rect 2704 2003 2772 2037
rect 2772 2003 2776 2037
rect 2598 1969 2776 2003
rect 2598 1935 2602 1969
rect 2602 1935 2670 1969
rect 2670 1935 2704 1969
rect 2704 1935 2772 1969
rect 2772 1935 2776 1969
rect 2598 1901 2776 1935
rect 2598 1867 2602 1901
rect 2602 1867 2670 1901
rect 2670 1867 2704 1901
rect 2704 1867 2772 1901
rect 2772 1867 2776 1901
rect 2598 1833 2776 1867
rect 2598 1799 2602 1833
rect 2602 1799 2670 1833
rect 2670 1799 2704 1833
rect 2704 1799 2772 1833
rect 2772 1799 2776 1833
rect 2598 1765 2776 1799
rect 2598 1731 2602 1765
rect 2602 1731 2670 1765
rect 2670 1731 2704 1765
rect 2704 1731 2772 1765
rect 2772 1731 2776 1765
rect 2598 1697 2776 1731
rect 2598 1663 2602 1697
rect 2602 1663 2670 1697
rect 2670 1663 2704 1697
rect 2704 1663 2772 1697
rect 2772 1663 2776 1697
rect 2598 1629 2776 1663
rect 2598 1595 2602 1629
rect 2602 1595 2670 1629
rect 2670 1595 2704 1629
rect 2704 1595 2772 1629
rect 2772 1595 2776 1629
rect 2598 1561 2776 1595
rect 2598 1527 2602 1561
rect 2602 1527 2670 1561
rect 2670 1527 2704 1561
rect 2704 1527 2772 1561
rect 2772 1527 2776 1561
rect 2598 1491 2776 1527
rect 2598 1479 2632 1491
rect 2742 1479 2776 1491
rect 3345 4388 3451 4494
rect 3094 4028 3128 4062
rect 3166 4028 3200 4062
rect 3238 4028 3272 4062
rect 3094 3954 3128 3988
rect 3166 3954 3200 3988
rect 3238 3954 3272 3988
rect 3094 3880 3128 3914
rect 3166 3880 3200 3914
rect 3238 3880 3272 3914
rect 3094 3806 3128 3840
rect 3166 3806 3200 3840
rect 3238 3806 3272 3840
rect 3094 3732 3128 3766
rect 3166 3732 3200 3766
rect 3238 3732 3272 3766
rect 3094 3658 3128 3692
rect 3166 3658 3200 3692
rect 3238 3658 3272 3692
rect 3094 3584 3128 3618
rect 3166 3584 3200 3618
rect 3238 3584 3272 3618
rect 3094 3510 3128 3544
rect 3166 3510 3200 3544
rect 3238 3510 3272 3544
rect 3094 3436 3128 3470
rect 3166 3436 3200 3470
rect 3238 3436 3272 3470
rect 3094 3362 3128 3396
rect 3166 3362 3200 3396
rect 3238 3362 3272 3396
rect 3094 3288 3128 3322
rect 3166 3288 3200 3322
rect 3238 3288 3272 3322
rect 3094 3214 3128 3248
rect 3166 3214 3200 3248
rect 3238 3214 3272 3248
rect 3094 3140 3128 3174
rect 3166 3140 3200 3174
rect 3238 3140 3272 3174
rect 3094 3066 3128 3100
rect 3166 3066 3200 3100
rect 3238 3066 3272 3100
rect 3094 2992 3128 3026
rect 3166 2992 3200 3026
rect 3238 2992 3272 3026
rect 3094 2918 3128 2952
rect 3166 2918 3200 2952
rect 3238 2918 3272 2952
rect 3094 2844 3128 2878
rect 3166 2844 3200 2878
rect 3238 2844 3272 2878
rect 3094 2770 3128 2804
rect 3166 2770 3200 2804
rect 3238 2770 3272 2804
rect 3094 2696 3128 2730
rect 3166 2696 3200 2730
rect 3238 2696 3272 2730
rect 3094 2622 3128 2656
rect 3166 2622 3200 2656
rect 3238 2622 3272 2656
rect 3094 2548 3128 2582
rect 3166 2548 3200 2582
rect 3238 2548 3272 2582
rect 3094 2474 3128 2508
rect 3166 2474 3200 2508
rect 3238 2474 3272 2508
rect 3094 2400 3128 2434
rect 3166 2400 3200 2434
rect 3238 2400 3272 2434
rect 3094 2326 3128 2360
rect 3166 2326 3200 2360
rect 3238 2326 3272 2360
rect 3094 2252 3128 2286
rect 3166 2252 3200 2286
rect 3238 2252 3272 2286
rect 3094 2178 3128 2212
rect 3166 2178 3200 2212
rect 3238 2178 3272 2212
rect 3094 2104 3128 2138
rect 3166 2104 3200 2138
rect 3238 2104 3272 2138
rect 3094 2030 3128 2064
rect 3166 2030 3200 2064
rect 3238 2030 3272 2064
rect 3094 1956 3128 1990
rect 3166 1956 3200 1990
rect 3238 1956 3272 1990
rect 3094 1882 3128 1916
rect 3166 1882 3200 1916
rect 3238 1882 3272 1916
rect 3094 1808 3128 1842
rect 3166 1808 3200 1842
rect 3238 1808 3272 1842
rect 3094 1734 3128 1768
rect 3166 1734 3200 1768
rect 3238 1734 3272 1768
rect 3094 1660 3128 1694
rect 3166 1660 3200 1694
rect 3238 1660 3272 1694
rect 3094 1586 3128 1620
rect 3166 1586 3200 1620
rect 3238 1586 3272 1620
rect 3094 1511 3128 1545
rect 3166 1511 3200 1545
rect 3238 1511 3272 1545
rect 3907 4388 4013 4494
rect 3662 4050 3696 4062
rect 3590 4046 3768 4050
rect 3590 4012 3594 4046
rect 3594 4012 3662 4046
rect 3662 4012 3696 4046
rect 3696 4012 3764 4046
rect 3764 4012 3768 4046
rect 3590 3978 3768 4012
rect 3590 3944 3594 3978
rect 3594 3944 3662 3978
rect 3662 3944 3696 3978
rect 3696 3944 3764 3978
rect 3764 3944 3768 3978
rect 3590 3910 3768 3944
rect 3590 3876 3594 3910
rect 3594 3876 3662 3910
rect 3662 3876 3696 3910
rect 3696 3876 3764 3910
rect 3764 3876 3768 3910
rect 3590 3842 3768 3876
rect 3590 3808 3594 3842
rect 3594 3808 3662 3842
rect 3662 3808 3696 3842
rect 3696 3808 3764 3842
rect 3764 3808 3768 3842
rect 3590 3774 3768 3808
rect 3590 3740 3594 3774
rect 3594 3740 3662 3774
rect 3662 3740 3696 3774
rect 3696 3740 3764 3774
rect 3764 3740 3768 3774
rect 3590 3706 3768 3740
rect 3590 3672 3594 3706
rect 3594 3672 3662 3706
rect 3662 3672 3696 3706
rect 3696 3672 3764 3706
rect 3764 3672 3768 3706
rect 3590 3638 3768 3672
rect 3590 3604 3594 3638
rect 3594 3604 3662 3638
rect 3662 3604 3696 3638
rect 3696 3604 3764 3638
rect 3764 3604 3768 3638
rect 3590 3570 3768 3604
rect 3590 3536 3594 3570
rect 3594 3536 3662 3570
rect 3662 3536 3696 3570
rect 3696 3536 3764 3570
rect 3764 3536 3768 3570
rect 3590 3502 3768 3536
rect 3590 3468 3594 3502
rect 3594 3468 3662 3502
rect 3662 3468 3696 3502
rect 3696 3468 3764 3502
rect 3764 3468 3768 3502
rect 3590 3434 3768 3468
rect 3590 3400 3594 3434
rect 3594 3400 3662 3434
rect 3662 3400 3696 3434
rect 3696 3400 3764 3434
rect 3764 3400 3768 3434
rect 3590 3366 3768 3400
rect 3590 3332 3594 3366
rect 3594 3332 3662 3366
rect 3662 3332 3696 3366
rect 3696 3332 3764 3366
rect 3764 3332 3768 3366
rect 3590 3298 3768 3332
rect 3590 3264 3594 3298
rect 3594 3264 3662 3298
rect 3662 3264 3696 3298
rect 3696 3264 3764 3298
rect 3764 3264 3768 3298
rect 3590 3230 3768 3264
rect 3590 3196 3594 3230
rect 3594 3196 3662 3230
rect 3662 3196 3696 3230
rect 3696 3196 3764 3230
rect 3764 3196 3768 3230
rect 3590 3162 3768 3196
rect 3590 3128 3594 3162
rect 3594 3128 3662 3162
rect 3662 3128 3696 3162
rect 3696 3128 3764 3162
rect 3764 3128 3768 3162
rect 3590 3092 3768 3128
rect 3590 3080 3624 3092
rect 3734 3080 3768 3092
rect 3590 2935 3768 3040
rect 3590 2901 3629 2935
rect 3629 2901 3663 2935
rect 3663 2901 3697 2935
rect 3697 2901 3731 2935
rect 3731 2901 3768 2935
rect 3590 2855 3768 2901
rect 3590 2821 3629 2855
rect 3629 2821 3663 2855
rect 3663 2821 3697 2855
rect 3697 2821 3731 2855
rect 3731 2821 3768 2855
rect 3590 2775 3768 2821
rect 3590 2741 3629 2775
rect 3629 2741 3663 2775
rect 3663 2741 3697 2775
rect 3697 2741 3731 2775
rect 3731 2741 3768 2775
rect 3590 2695 3768 2741
rect 3590 2661 3629 2695
rect 3629 2661 3663 2695
rect 3663 2661 3697 2695
rect 3697 2661 3731 2695
rect 3731 2661 3768 2695
rect 3590 2614 3768 2661
rect 3590 2580 3629 2614
rect 3629 2580 3663 2614
rect 3663 2580 3697 2614
rect 3697 2580 3731 2614
rect 3731 2580 3768 2614
rect 3590 2574 3768 2580
rect 3590 2501 3624 2535
rect 3662 2501 3696 2535
rect 3734 2501 3768 2535
rect 3662 2449 3696 2461
rect 3590 2445 3768 2449
rect 3590 2411 3594 2445
rect 3594 2411 3662 2445
rect 3662 2411 3696 2445
rect 3696 2411 3764 2445
rect 3764 2411 3768 2445
rect 3590 2377 3768 2411
rect 3590 2343 3594 2377
rect 3594 2343 3662 2377
rect 3662 2343 3696 2377
rect 3696 2343 3764 2377
rect 3764 2343 3768 2377
rect 3590 2309 3768 2343
rect 3590 2275 3594 2309
rect 3594 2275 3662 2309
rect 3662 2275 3696 2309
rect 3696 2275 3764 2309
rect 3764 2275 3768 2309
rect 3590 2241 3768 2275
rect 3590 2207 3594 2241
rect 3594 2207 3662 2241
rect 3662 2207 3696 2241
rect 3696 2207 3764 2241
rect 3764 2207 3768 2241
rect 3590 2173 3768 2207
rect 3590 2139 3594 2173
rect 3594 2139 3662 2173
rect 3662 2139 3696 2173
rect 3696 2139 3764 2173
rect 3764 2139 3768 2173
rect 3590 2105 3768 2139
rect 3590 2071 3594 2105
rect 3594 2071 3662 2105
rect 3662 2071 3696 2105
rect 3696 2071 3764 2105
rect 3764 2071 3768 2105
rect 3590 2037 3768 2071
rect 3590 2003 3594 2037
rect 3594 2003 3662 2037
rect 3662 2003 3696 2037
rect 3696 2003 3764 2037
rect 3764 2003 3768 2037
rect 3590 1969 3768 2003
rect 3590 1935 3594 1969
rect 3594 1935 3662 1969
rect 3662 1935 3696 1969
rect 3696 1935 3764 1969
rect 3764 1935 3768 1969
rect 3590 1901 3768 1935
rect 3590 1867 3594 1901
rect 3594 1867 3662 1901
rect 3662 1867 3696 1901
rect 3696 1867 3764 1901
rect 3764 1867 3768 1901
rect 3590 1833 3768 1867
rect 3590 1799 3594 1833
rect 3594 1799 3662 1833
rect 3662 1799 3696 1833
rect 3696 1799 3764 1833
rect 3764 1799 3768 1833
rect 3590 1765 3768 1799
rect 3590 1731 3594 1765
rect 3594 1731 3662 1765
rect 3662 1731 3696 1765
rect 3696 1731 3764 1765
rect 3764 1731 3768 1765
rect 3590 1697 3768 1731
rect 3590 1663 3594 1697
rect 3594 1663 3662 1697
rect 3662 1663 3696 1697
rect 3696 1663 3764 1697
rect 3764 1663 3768 1697
rect 3590 1629 3768 1663
rect 3590 1595 3594 1629
rect 3594 1595 3662 1629
rect 3662 1595 3696 1629
rect 3696 1595 3764 1629
rect 3764 1595 3768 1629
rect 3590 1561 3768 1595
rect 3590 1527 3594 1561
rect 3594 1527 3662 1561
rect 3662 1527 3696 1561
rect 3696 1527 3764 1561
rect 3764 1527 3768 1561
rect 3590 1491 3768 1527
rect 3590 1479 3624 1491
rect 3734 1479 3768 1491
rect 4337 4388 4443 4494
rect 4086 4028 4120 4062
rect 4158 4028 4192 4062
rect 4230 4028 4264 4062
rect 4086 3954 4120 3988
rect 4158 3954 4192 3988
rect 4230 3954 4264 3988
rect 4086 3880 4120 3914
rect 4158 3880 4192 3914
rect 4230 3880 4264 3914
rect 4086 3806 4120 3840
rect 4158 3806 4192 3840
rect 4230 3806 4264 3840
rect 4086 3732 4120 3766
rect 4158 3732 4192 3766
rect 4230 3732 4264 3766
rect 4086 3658 4120 3692
rect 4158 3658 4192 3692
rect 4230 3658 4264 3692
rect 4086 3584 4120 3618
rect 4158 3584 4192 3618
rect 4230 3584 4264 3618
rect 4086 3510 4120 3544
rect 4158 3510 4192 3544
rect 4230 3510 4264 3544
rect 4086 3436 4120 3470
rect 4158 3436 4192 3470
rect 4230 3436 4264 3470
rect 4086 3362 4120 3396
rect 4158 3362 4192 3396
rect 4230 3362 4264 3396
rect 4086 3288 4120 3322
rect 4158 3288 4192 3322
rect 4230 3288 4264 3322
rect 4086 3214 4120 3248
rect 4158 3214 4192 3248
rect 4230 3214 4264 3248
rect 4086 3140 4120 3174
rect 4158 3140 4192 3174
rect 4230 3140 4264 3174
rect 4086 3066 4120 3100
rect 4158 3066 4192 3100
rect 4230 3066 4264 3100
rect 4086 2992 4120 3026
rect 4158 2992 4192 3026
rect 4230 2992 4264 3026
rect 4086 2918 4120 2952
rect 4158 2918 4192 2952
rect 4230 2918 4264 2952
rect 4086 2844 4120 2878
rect 4158 2844 4192 2878
rect 4230 2844 4264 2878
rect 4086 2770 4120 2804
rect 4158 2770 4192 2804
rect 4230 2770 4264 2804
rect 4086 2696 4120 2730
rect 4158 2696 4192 2730
rect 4230 2696 4264 2730
rect 4086 2622 4120 2656
rect 4158 2622 4192 2656
rect 4230 2622 4264 2656
rect 4086 2548 4120 2582
rect 4158 2548 4192 2582
rect 4230 2548 4264 2582
rect 4086 2474 4120 2508
rect 4158 2474 4192 2508
rect 4230 2474 4264 2508
rect 4086 2400 4120 2434
rect 4158 2400 4192 2434
rect 4230 2400 4264 2434
rect 4086 2326 4120 2360
rect 4158 2326 4192 2360
rect 4230 2326 4264 2360
rect 4086 2252 4120 2286
rect 4158 2252 4192 2286
rect 4230 2252 4264 2286
rect 4086 2178 4120 2212
rect 4158 2178 4192 2212
rect 4230 2178 4264 2212
rect 4086 2104 4120 2138
rect 4158 2104 4192 2138
rect 4230 2104 4264 2138
rect 4086 2030 4120 2064
rect 4158 2030 4192 2064
rect 4230 2030 4264 2064
rect 4086 1956 4120 1990
rect 4158 1956 4192 1990
rect 4230 1956 4264 1990
rect 4086 1882 4120 1916
rect 4158 1882 4192 1916
rect 4230 1882 4264 1916
rect 4086 1808 4120 1842
rect 4158 1808 4192 1842
rect 4230 1808 4264 1842
rect 4086 1734 4120 1768
rect 4158 1734 4192 1768
rect 4230 1734 4264 1768
rect 4086 1660 4120 1694
rect 4158 1660 4192 1694
rect 4230 1660 4264 1694
rect 4086 1586 4120 1620
rect 4158 1586 4192 1620
rect 4230 1586 4264 1620
rect 4086 1511 4120 1545
rect 4158 1511 4192 1545
rect 4230 1511 4264 1545
rect 4899 4388 5005 4494
rect 4654 4050 4688 4062
rect 4582 4046 4760 4050
rect 4582 4012 4586 4046
rect 4586 4012 4654 4046
rect 4654 4012 4688 4046
rect 4688 4012 4756 4046
rect 4756 4012 4760 4046
rect 4582 3978 4760 4012
rect 4582 3944 4586 3978
rect 4586 3944 4654 3978
rect 4654 3944 4688 3978
rect 4688 3944 4756 3978
rect 4756 3944 4760 3978
rect 4582 3910 4760 3944
rect 4582 3876 4586 3910
rect 4586 3876 4654 3910
rect 4654 3876 4688 3910
rect 4688 3876 4756 3910
rect 4756 3876 4760 3910
rect 4582 3842 4760 3876
rect 4582 3808 4586 3842
rect 4586 3808 4654 3842
rect 4654 3808 4688 3842
rect 4688 3808 4756 3842
rect 4756 3808 4760 3842
rect 4582 3774 4760 3808
rect 4582 3740 4586 3774
rect 4586 3740 4654 3774
rect 4654 3740 4688 3774
rect 4688 3740 4756 3774
rect 4756 3740 4760 3774
rect 4582 3706 4760 3740
rect 4582 3672 4586 3706
rect 4586 3672 4654 3706
rect 4654 3672 4688 3706
rect 4688 3672 4756 3706
rect 4756 3672 4760 3706
rect 4582 3638 4760 3672
rect 4582 3604 4586 3638
rect 4586 3604 4654 3638
rect 4654 3604 4688 3638
rect 4688 3604 4756 3638
rect 4756 3604 4760 3638
rect 4582 3570 4760 3604
rect 4582 3536 4586 3570
rect 4586 3536 4654 3570
rect 4654 3536 4688 3570
rect 4688 3536 4756 3570
rect 4756 3536 4760 3570
rect 4582 3502 4760 3536
rect 4582 3468 4586 3502
rect 4586 3468 4654 3502
rect 4654 3468 4688 3502
rect 4688 3468 4756 3502
rect 4756 3468 4760 3502
rect 4582 3434 4760 3468
rect 4582 3400 4586 3434
rect 4586 3400 4654 3434
rect 4654 3400 4688 3434
rect 4688 3400 4756 3434
rect 4756 3400 4760 3434
rect 4582 3366 4760 3400
rect 4582 3332 4586 3366
rect 4586 3332 4654 3366
rect 4654 3332 4688 3366
rect 4688 3332 4756 3366
rect 4756 3332 4760 3366
rect 4582 3298 4760 3332
rect 4582 3264 4586 3298
rect 4586 3264 4654 3298
rect 4654 3264 4688 3298
rect 4688 3264 4756 3298
rect 4756 3264 4760 3298
rect 4582 3230 4760 3264
rect 4582 3196 4586 3230
rect 4586 3196 4654 3230
rect 4654 3196 4688 3230
rect 4688 3196 4756 3230
rect 4756 3196 4760 3230
rect 4582 3162 4760 3196
rect 4582 3128 4586 3162
rect 4586 3128 4654 3162
rect 4654 3128 4688 3162
rect 4688 3128 4756 3162
rect 4756 3128 4760 3162
rect 4582 3092 4760 3128
rect 4582 3080 4616 3092
rect 4726 3080 4760 3092
rect 4582 2935 4760 3040
rect 4582 2901 4621 2935
rect 4621 2901 4655 2935
rect 4655 2901 4689 2935
rect 4689 2901 4723 2935
rect 4723 2901 4760 2935
rect 4582 2855 4760 2901
rect 4582 2821 4621 2855
rect 4621 2821 4655 2855
rect 4655 2821 4689 2855
rect 4689 2821 4723 2855
rect 4723 2821 4760 2855
rect 4582 2775 4760 2821
rect 4582 2741 4621 2775
rect 4621 2741 4655 2775
rect 4655 2741 4689 2775
rect 4689 2741 4723 2775
rect 4723 2741 4760 2775
rect 4582 2695 4760 2741
rect 4582 2661 4621 2695
rect 4621 2661 4655 2695
rect 4655 2661 4689 2695
rect 4689 2661 4723 2695
rect 4723 2661 4760 2695
rect 4582 2614 4760 2661
rect 4582 2580 4621 2614
rect 4621 2580 4655 2614
rect 4655 2580 4689 2614
rect 4689 2580 4723 2614
rect 4723 2580 4760 2614
rect 4582 2574 4760 2580
rect 4582 2501 4616 2535
rect 4654 2501 4688 2535
rect 4726 2501 4760 2535
rect 4654 2449 4688 2461
rect 4582 2445 4760 2449
rect 4582 2411 4586 2445
rect 4586 2411 4654 2445
rect 4654 2411 4688 2445
rect 4688 2411 4756 2445
rect 4756 2411 4760 2445
rect 4582 2377 4760 2411
rect 4582 2343 4586 2377
rect 4586 2343 4654 2377
rect 4654 2343 4688 2377
rect 4688 2343 4756 2377
rect 4756 2343 4760 2377
rect 4582 2309 4760 2343
rect 4582 2275 4586 2309
rect 4586 2275 4654 2309
rect 4654 2275 4688 2309
rect 4688 2275 4756 2309
rect 4756 2275 4760 2309
rect 4582 2241 4760 2275
rect 4582 2207 4586 2241
rect 4586 2207 4654 2241
rect 4654 2207 4688 2241
rect 4688 2207 4756 2241
rect 4756 2207 4760 2241
rect 4582 2173 4760 2207
rect 4582 2139 4586 2173
rect 4586 2139 4654 2173
rect 4654 2139 4688 2173
rect 4688 2139 4756 2173
rect 4756 2139 4760 2173
rect 4582 2105 4760 2139
rect 4582 2071 4586 2105
rect 4586 2071 4654 2105
rect 4654 2071 4688 2105
rect 4688 2071 4756 2105
rect 4756 2071 4760 2105
rect 4582 2037 4760 2071
rect 4582 2003 4586 2037
rect 4586 2003 4654 2037
rect 4654 2003 4688 2037
rect 4688 2003 4756 2037
rect 4756 2003 4760 2037
rect 4582 1969 4760 2003
rect 4582 1935 4586 1969
rect 4586 1935 4654 1969
rect 4654 1935 4688 1969
rect 4688 1935 4756 1969
rect 4756 1935 4760 1969
rect 4582 1901 4760 1935
rect 4582 1867 4586 1901
rect 4586 1867 4654 1901
rect 4654 1867 4688 1901
rect 4688 1867 4756 1901
rect 4756 1867 4760 1901
rect 4582 1833 4760 1867
rect 4582 1799 4586 1833
rect 4586 1799 4654 1833
rect 4654 1799 4688 1833
rect 4688 1799 4756 1833
rect 4756 1799 4760 1833
rect 4582 1765 4760 1799
rect 4582 1731 4586 1765
rect 4586 1731 4654 1765
rect 4654 1731 4688 1765
rect 4688 1731 4756 1765
rect 4756 1731 4760 1765
rect 4582 1697 4760 1731
rect 4582 1663 4586 1697
rect 4586 1663 4654 1697
rect 4654 1663 4688 1697
rect 4688 1663 4756 1697
rect 4756 1663 4760 1697
rect 4582 1629 4760 1663
rect 4582 1595 4586 1629
rect 4586 1595 4654 1629
rect 4654 1595 4688 1629
rect 4688 1595 4756 1629
rect 4756 1595 4760 1629
rect 4582 1561 4760 1595
rect 4582 1527 4586 1561
rect 4586 1527 4654 1561
rect 4654 1527 4688 1561
rect 4688 1527 4756 1561
rect 4756 1527 4760 1561
rect 4582 1491 4760 1527
rect 4582 1479 4616 1491
rect 4726 1479 4760 1491
rect 5329 4388 5435 4494
rect 5078 4028 5112 4062
rect 5150 4028 5184 4062
rect 5222 4028 5256 4062
rect 5078 3954 5112 3988
rect 5150 3954 5184 3988
rect 5222 3954 5256 3988
rect 5078 3880 5112 3914
rect 5150 3880 5184 3914
rect 5222 3880 5256 3914
rect 5078 3806 5112 3840
rect 5150 3806 5184 3840
rect 5222 3806 5256 3840
rect 5078 3732 5112 3766
rect 5150 3732 5184 3766
rect 5222 3732 5256 3766
rect 5078 3658 5112 3692
rect 5150 3658 5184 3692
rect 5222 3658 5256 3692
rect 5078 3584 5112 3618
rect 5150 3584 5184 3618
rect 5222 3584 5256 3618
rect 5078 3510 5112 3544
rect 5150 3510 5184 3544
rect 5222 3510 5256 3544
rect 5078 3436 5112 3470
rect 5150 3436 5184 3470
rect 5222 3436 5256 3470
rect 5078 3362 5112 3396
rect 5150 3362 5184 3396
rect 5222 3362 5256 3396
rect 5078 3288 5112 3322
rect 5150 3288 5184 3322
rect 5222 3288 5256 3322
rect 5078 3214 5112 3248
rect 5150 3214 5184 3248
rect 5222 3214 5256 3248
rect 5078 3140 5112 3174
rect 5150 3140 5184 3174
rect 5222 3140 5256 3174
rect 5078 3066 5112 3100
rect 5150 3066 5184 3100
rect 5222 3066 5256 3100
rect 5078 2992 5112 3026
rect 5150 2992 5184 3026
rect 5222 2992 5256 3026
rect 5078 2918 5112 2952
rect 5150 2918 5184 2952
rect 5222 2918 5256 2952
rect 5078 2844 5112 2878
rect 5150 2844 5184 2878
rect 5222 2844 5256 2878
rect 5078 2770 5112 2804
rect 5150 2770 5184 2804
rect 5222 2770 5256 2804
rect 5078 2696 5112 2730
rect 5150 2696 5184 2730
rect 5222 2696 5256 2730
rect 5078 2622 5112 2656
rect 5150 2622 5184 2656
rect 5222 2622 5256 2656
rect 5078 2548 5112 2582
rect 5150 2548 5184 2582
rect 5222 2548 5256 2582
rect 5078 2474 5112 2508
rect 5150 2474 5184 2508
rect 5222 2474 5256 2508
rect 5078 2400 5112 2434
rect 5150 2400 5184 2434
rect 5222 2400 5256 2434
rect 5078 2326 5112 2360
rect 5150 2326 5184 2360
rect 5222 2326 5256 2360
rect 5078 2252 5112 2286
rect 5150 2252 5184 2286
rect 5222 2252 5256 2286
rect 5078 2178 5112 2212
rect 5150 2178 5184 2212
rect 5222 2178 5256 2212
rect 5078 2104 5112 2138
rect 5150 2104 5184 2138
rect 5222 2104 5256 2138
rect 5078 2030 5112 2064
rect 5150 2030 5184 2064
rect 5222 2030 5256 2064
rect 5078 1956 5112 1990
rect 5150 1956 5184 1990
rect 5222 1956 5256 1990
rect 5078 1882 5112 1916
rect 5150 1882 5184 1916
rect 5222 1882 5256 1916
rect 5078 1808 5112 1842
rect 5150 1808 5184 1842
rect 5222 1808 5256 1842
rect 5078 1734 5112 1768
rect 5150 1734 5184 1768
rect 5222 1734 5256 1768
rect 5078 1660 5112 1694
rect 5150 1660 5184 1694
rect 5222 1660 5256 1694
rect 5078 1586 5112 1620
rect 5150 1586 5184 1620
rect 5222 1586 5256 1620
rect 5078 1511 5112 1545
rect 5150 1511 5184 1545
rect 5222 1511 5256 1545
rect 5891 4388 5997 4494
rect 5646 4050 5680 4062
rect 5574 4046 5752 4050
rect 5574 4012 5578 4046
rect 5578 4012 5646 4046
rect 5646 4012 5680 4046
rect 5680 4012 5748 4046
rect 5748 4012 5752 4046
rect 5574 3978 5752 4012
rect 5574 3944 5578 3978
rect 5578 3944 5646 3978
rect 5646 3944 5680 3978
rect 5680 3944 5748 3978
rect 5748 3944 5752 3978
rect 5574 3910 5752 3944
rect 5574 3876 5578 3910
rect 5578 3876 5646 3910
rect 5646 3876 5680 3910
rect 5680 3876 5748 3910
rect 5748 3876 5752 3910
rect 5574 3842 5752 3876
rect 5574 3808 5578 3842
rect 5578 3808 5646 3842
rect 5646 3808 5680 3842
rect 5680 3808 5748 3842
rect 5748 3808 5752 3842
rect 5574 3774 5752 3808
rect 5574 3740 5578 3774
rect 5578 3740 5646 3774
rect 5646 3740 5680 3774
rect 5680 3740 5748 3774
rect 5748 3740 5752 3774
rect 5574 3706 5752 3740
rect 5574 3672 5578 3706
rect 5578 3672 5646 3706
rect 5646 3672 5680 3706
rect 5680 3672 5748 3706
rect 5748 3672 5752 3706
rect 5574 3638 5752 3672
rect 5574 3604 5578 3638
rect 5578 3604 5646 3638
rect 5646 3604 5680 3638
rect 5680 3604 5748 3638
rect 5748 3604 5752 3638
rect 5574 3570 5752 3604
rect 5574 3536 5578 3570
rect 5578 3536 5646 3570
rect 5646 3536 5680 3570
rect 5680 3536 5748 3570
rect 5748 3536 5752 3570
rect 5574 3502 5752 3536
rect 5574 3468 5578 3502
rect 5578 3468 5646 3502
rect 5646 3468 5680 3502
rect 5680 3468 5748 3502
rect 5748 3468 5752 3502
rect 5574 3434 5752 3468
rect 5574 3400 5578 3434
rect 5578 3400 5646 3434
rect 5646 3400 5680 3434
rect 5680 3400 5748 3434
rect 5748 3400 5752 3434
rect 5574 3366 5752 3400
rect 5574 3332 5578 3366
rect 5578 3332 5646 3366
rect 5646 3332 5680 3366
rect 5680 3332 5748 3366
rect 5748 3332 5752 3366
rect 5574 3298 5752 3332
rect 5574 3264 5578 3298
rect 5578 3264 5646 3298
rect 5646 3264 5680 3298
rect 5680 3264 5748 3298
rect 5748 3264 5752 3298
rect 5574 3230 5752 3264
rect 5574 3196 5578 3230
rect 5578 3196 5646 3230
rect 5646 3196 5680 3230
rect 5680 3196 5748 3230
rect 5748 3196 5752 3230
rect 5574 3162 5752 3196
rect 5574 3128 5578 3162
rect 5578 3128 5646 3162
rect 5646 3128 5680 3162
rect 5680 3128 5748 3162
rect 5748 3128 5752 3162
rect 5574 3092 5752 3128
rect 5574 3080 5608 3092
rect 5718 3080 5752 3092
rect 5574 2935 5752 3040
rect 5574 2901 5613 2935
rect 5613 2901 5647 2935
rect 5647 2901 5681 2935
rect 5681 2901 5715 2935
rect 5715 2901 5752 2935
rect 5574 2855 5752 2901
rect 5574 2821 5613 2855
rect 5613 2821 5647 2855
rect 5647 2821 5681 2855
rect 5681 2821 5715 2855
rect 5715 2821 5752 2855
rect 5574 2775 5752 2821
rect 5574 2741 5613 2775
rect 5613 2741 5647 2775
rect 5647 2741 5681 2775
rect 5681 2741 5715 2775
rect 5715 2741 5752 2775
rect 5574 2695 5752 2741
rect 5574 2661 5613 2695
rect 5613 2661 5647 2695
rect 5647 2661 5681 2695
rect 5681 2661 5715 2695
rect 5715 2661 5752 2695
rect 5574 2614 5752 2661
rect 5574 2580 5613 2614
rect 5613 2580 5647 2614
rect 5647 2580 5681 2614
rect 5681 2580 5715 2614
rect 5715 2580 5752 2614
rect 5574 2574 5752 2580
rect 5574 2501 5608 2535
rect 5646 2501 5680 2535
rect 5718 2501 5752 2535
rect 5646 2449 5680 2461
rect 5574 2445 5752 2449
rect 5574 2411 5578 2445
rect 5578 2411 5646 2445
rect 5646 2411 5680 2445
rect 5680 2411 5748 2445
rect 5748 2411 5752 2445
rect 5574 2377 5752 2411
rect 5574 2343 5578 2377
rect 5578 2343 5646 2377
rect 5646 2343 5680 2377
rect 5680 2343 5748 2377
rect 5748 2343 5752 2377
rect 5574 2309 5752 2343
rect 5574 2275 5578 2309
rect 5578 2275 5646 2309
rect 5646 2275 5680 2309
rect 5680 2275 5748 2309
rect 5748 2275 5752 2309
rect 5574 2241 5752 2275
rect 5574 2207 5578 2241
rect 5578 2207 5646 2241
rect 5646 2207 5680 2241
rect 5680 2207 5748 2241
rect 5748 2207 5752 2241
rect 5574 2173 5752 2207
rect 5574 2139 5578 2173
rect 5578 2139 5646 2173
rect 5646 2139 5680 2173
rect 5680 2139 5748 2173
rect 5748 2139 5752 2173
rect 5574 2105 5752 2139
rect 5574 2071 5578 2105
rect 5578 2071 5646 2105
rect 5646 2071 5680 2105
rect 5680 2071 5748 2105
rect 5748 2071 5752 2105
rect 5574 2037 5752 2071
rect 5574 2003 5578 2037
rect 5578 2003 5646 2037
rect 5646 2003 5680 2037
rect 5680 2003 5748 2037
rect 5748 2003 5752 2037
rect 5574 1969 5752 2003
rect 5574 1935 5578 1969
rect 5578 1935 5646 1969
rect 5646 1935 5680 1969
rect 5680 1935 5748 1969
rect 5748 1935 5752 1969
rect 5574 1901 5752 1935
rect 5574 1867 5578 1901
rect 5578 1867 5646 1901
rect 5646 1867 5680 1901
rect 5680 1867 5748 1901
rect 5748 1867 5752 1901
rect 5574 1833 5752 1867
rect 5574 1799 5578 1833
rect 5578 1799 5646 1833
rect 5646 1799 5680 1833
rect 5680 1799 5748 1833
rect 5748 1799 5752 1833
rect 5574 1765 5752 1799
rect 5574 1731 5578 1765
rect 5578 1731 5646 1765
rect 5646 1731 5680 1765
rect 5680 1731 5748 1765
rect 5748 1731 5752 1765
rect 5574 1697 5752 1731
rect 5574 1663 5578 1697
rect 5578 1663 5646 1697
rect 5646 1663 5680 1697
rect 5680 1663 5748 1697
rect 5748 1663 5752 1697
rect 5574 1629 5752 1663
rect 5574 1595 5578 1629
rect 5578 1595 5646 1629
rect 5646 1595 5680 1629
rect 5680 1595 5748 1629
rect 5748 1595 5752 1629
rect 5574 1561 5752 1595
rect 5574 1527 5578 1561
rect 5578 1527 5646 1561
rect 5646 1527 5680 1561
rect 5680 1527 5748 1561
rect 5748 1527 5752 1561
rect 5574 1491 5752 1527
rect 5574 1479 5608 1491
rect 5718 1479 5752 1491
rect 6321 4388 6427 4494
rect 6868 4388 6974 4494
rect 6070 4028 6104 4062
rect 6142 4028 6176 4062
rect 6214 4028 6248 4062
rect 6070 3954 6104 3988
rect 6142 3954 6176 3988
rect 6214 3954 6248 3988
rect 6070 3880 6104 3914
rect 6142 3880 6176 3914
rect 6214 3880 6248 3914
rect 6070 3806 6104 3840
rect 6142 3806 6176 3840
rect 6214 3806 6248 3840
rect 6070 3732 6104 3766
rect 6142 3732 6176 3766
rect 6214 3732 6248 3766
rect 6070 3658 6104 3692
rect 6142 3658 6176 3692
rect 6214 3658 6248 3692
rect 6070 3584 6104 3618
rect 6142 3584 6176 3618
rect 6214 3584 6248 3618
rect 6070 3510 6104 3544
rect 6142 3510 6176 3544
rect 6214 3510 6248 3544
rect 6070 3436 6104 3470
rect 6142 3436 6176 3470
rect 6214 3436 6248 3470
rect 6070 3362 6104 3396
rect 6142 3362 6176 3396
rect 6214 3362 6248 3396
rect 6070 3288 6104 3322
rect 6142 3288 6176 3322
rect 6214 3288 6248 3322
rect 6070 3214 6104 3248
rect 6142 3214 6176 3248
rect 6214 3214 6248 3248
rect 6070 3140 6104 3174
rect 6142 3140 6176 3174
rect 6214 3140 6248 3174
rect 6070 3066 6104 3100
rect 6142 3066 6176 3100
rect 6214 3066 6248 3100
rect 6070 2992 6104 3026
rect 6142 2992 6176 3026
rect 6214 2992 6248 3026
rect 6070 2918 6104 2952
rect 6142 2918 6176 2952
rect 6214 2918 6248 2952
rect 6070 2844 6104 2878
rect 6142 2844 6176 2878
rect 6214 2844 6248 2878
rect 6070 2770 6104 2804
rect 6142 2770 6176 2804
rect 6214 2770 6248 2804
rect 6070 2696 6104 2730
rect 6142 2696 6176 2730
rect 6214 2696 6248 2730
rect 6070 2622 6104 2656
rect 6142 2622 6176 2656
rect 6214 2622 6248 2656
rect 6070 2548 6104 2582
rect 6142 2548 6176 2582
rect 6214 2548 6248 2582
rect 6070 2474 6104 2508
rect 6142 2474 6176 2508
rect 6214 2474 6248 2508
rect 6070 2400 6104 2434
rect 6142 2400 6176 2434
rect 6214 2400 6248 2434
rect 6070 2326 6104 2360
rect 6142 2326 6176 2360
rect 6214 2326 6248 2360
rect 6070 2252 6104 2286
rect 6142 2252 6176 2286
rect 6214 2252 6248 2286
rect 6070 2178 6104 2212
rect 6142 2178 6176 2212
rect 6214 2178 6248 2212
rect 6070 2104 6104 2138
rect 6142 2104 6176 2138
rect 6214 2104 6248 2138
rect 6070 2030 6104 2064
rect 6142 2030 6176 2064
rect 6214 2030 6248 2064
rect 6070 1956 6104 1990
rect 6142 1956 6176 1990
rect 6214 1956 6248 1990
rect 6070 1882 6104 1916
rect 6142 1882 6176 1916
rect 6214 1882 6248 1916
rect 6070 1808 6104 1842
rect 6142 1808 6176 1842
rect 6214 1808 6248 1842
rect 6070 1734 6104 1768
rect 6142 1734 6176 1768
rect 6214 1734 6248 1768
rect 6070 1660 6104 1694
rect 6142 1660 6176 1694
rect 6214 1660 6248 1694
rect 6070 1586 6104 1620
rect 6142 1586 6176 1620
rect 6214 1586 6248 1620
rect 6070 1511 6104 1545
rect 6142 1511 6176 1545
rect 6214 1511 6248 1545
rect 6638 4050 6672 4062
rect 6566 4046 6744 4050
rect 6566 4012 6570 4046
rect 6570 4012 6638 4046
rect 6638 4012 6672 4046
rect 6672 4012 6740 4046
rect 6740 4012 6744 4046
rect 6566 3978 6744 4012
rect 6566 3944 6570 3978
rect 6570 3944 6638 3978
rect 6638 3944 6672 3978
rect 6672 3944 6740 3978
rect 6740 3944 6744 3978
rect 6566 3910 6744 3944
rect 6566 3876 6570 3910
rect 6570 3876 6638 3910
rect 6638 3876 6672 3910
rect 6672 3876 6740 3910
rect 6740 3876 6744 3910
rect 6566 3842 6744 3876
rect 6566 3808 6570 3842
rect 6570 3808 6638 3842
rect 6638 3808 6672 3842
rect 6672 3808 6740 3842
rect 6740 3808 6744 3842
rect 6566 3774 6744 3808
rect 6566 3740 6570 3774
rect 6570 3740 6638 3774
rect 6638 3740 6672 3774
rect 6672 3740 6740 3774
rect 6740 3740 6744 3774
rect 6566 3706 6744 3740
rect 6566 3672 6570 3706
rect 6570 3672 6638 3706
rect 6638 3672 6672 3706
rect 6672 3672 6740 3706
rect 6740 3672 6744 3706
rect 6566 3638 6744 3672
rect 6566 3604 6570 3638
rect 6570 3604 6638 3638
rect 6638 3604 6672 3638
rect 6672 3604 6740 3638
rect 6740 3604 6744 3638
rect 6566 3570 6744 3604
rect 6566 3536 6570 3570
rect 6570 3536 6638 3570
rect 6638 3536 6672 3570
rect 6672 3536 6740 3570
rect 6740 3536 6744 3570
rect 6566 3502 6744 3536
rect 6566 3468 6570 3502
rect 6570 3468 6638 3502
rect 6638 3468 6672 3502
rect 6672 3468 6740 3502
rect 6740 3468 6744 3502
rect 6566 3434 6744 3468
rect 6566 3400 6570 3434
rect 6570 3400 6638 3434
rect 6638 3400 6672 3434
rect 6672 3400 6740 3434
rect 6740 3400 6744 3434
rect 6566 3366 6744 3400
rect 6566 3332 6570 3366
rect 6570 3332 6638 3366
rect 6638 3332 6672 3366
rect 6672 3332 6740 3366
rect 6740 3332 6744 3366
rect 6566 3298 6744 3332
rect 6566 3264 6570 3298
rect 6570 3264 6638 3298
rect 6638 3264 6672 3298
rect 6672 3264 6740 3298
rect 6740 3264 6744 3298
rect 6566 3230 6744 3264
rect 6566 3196 6570 3230
rect 6570 3196 6638 3230
rect 6638 3196 6672 3230
rect 6672 3196 6740 3230
rect 6740 3196 6744 3230
rect 6566 3162 6744 3196
rect 6566 3128 6570 3162
rect 6570 3128 6638 3162
rect 6638 3128 6672 3162
rect 6672 3128 6740 3162
rect 6740 3128 6744 3162
rect 6566 3092 6744 3128
rect 6566 3080 6600 3092
rect 6710 3080 6744 3092
rect 6566 2935 6744 3040
rect 6566 2901 6605 2935
rect 6605 2901 6639 2935
rect 6639 2901 6673 2935
rect 6673 2901 6707 2935
rect 6707 2901 6744 2935
rect 6566 2855 6744 2901
rect 6566 2821 6605 2855
rect 6605 2821 6639 2855
rect 6639 2821 6673 2855
rect 6673 2821 6707 2855
rect 6707 2821 6744 2855
rect 6566 2775 6744 2821
rect 6566 2741 6605 2775
rect 6605 2741 6639 2775
rect 6639 2741 6673 2775
rect 6673 2741 6707 2775
rect 6707 2741 6744 2775
rect 6566 2695 6744 2741
rect 6566 2661 6605 2695
rect 6605 2661 6639 2695
rect 6639 2661 6673 2695
rect 6673 2661 6707 2695
rect 6707 2661 6744 2695
rect 6566 2614 6744 2661
rect 6566 2580 6605 2614
rect 6605 2580 6639 2614
rect 6639 2580 6673 2614
rect 6673 2580 6707 2614
rect 6707 2580 6744 2614
rect 6566 2574 6744 2580
rect 6566 2501 6600 2535
rect 6638 2501 6672 2535
rect 6710 2501 6744 2535
rect 6638 2449 6672 2461
rect 6566 2445 6744 2449
rect 6566 2411 6570 2445
rect 6570 2411 6638 2445
rect 6638 2411 6672 2445
rect 6672 2411 6740 2445
rect 6740 2411 6744 2445
rect 6566 2377 6744 2411
rect 6566 2343 6570 2377
rect 6570 2343 6638 2377
rect 6638 2343 6672 2377
rect 6672 2343 6740 2377
rect 6740 2343 6744 2377
rect 6566 2309 6744 2343
rect 6566 2275 6570 2309
rect 6570 2275 6638 2309
rect 6638 2275 6672 2309
rect 6672 2275 6740 2309
rect 6740 2275 6744 2309
rect 6566 2241 6744 2275
rect 6566 2207 6570 2241
rect 6570 2207 6638 2241
rect 6638 2207 6672 2241
rect 6672 2207 6740 2241
rect 6740 2207 6744 2241
rect 6566 2173 6744 2207
rect 6566 2139 6570 2173
rect 6570 2139 6638 2173
rect 6638 2139 6672 2173
rect 6672 2139 6740 2173
rect 6740 2139 6744 2173
rect 6566 2105 6744 2139
rect 6566 2071 6570 2105
rect 6570 2071 6638 2105
rect 6638 2071 6672 2105
rect 6672 2071 6740 2105
rect 6740 2071 6744 2105
rect 6566 2037 6744 2071
rect 6566 2003 6570 2037
rect 6570 2003 6638 2037
rect 6638 2003 6672 2037
rect 6672 2003 6740 2037
rect 6740 2003 6744 2037
rect 6566 1969 6744 2003
rect 6566 1935 6570 1969
rect 6570 1935 6638 1969
rect 6638 1935 6672 1969
rect 6672 1935 6740 1969
rect 6740 1935 6744 1969
rect 6566 1901 6744 1935
rect 6566 1867 6570 1901
rect 6570 1867 6638 1901
rect 6638 1867 6672 1901
rect 6672 1867 6740 1901
rect 6740 1867 6744 1901
rect 6566 1833 6744 1867
rect 6566 1799 6570 1833
rect 6570 1799 6638 1833
rect 6638 1799 6672 1833
rect 6672 1799 6740 1833
rect 6740 1799 6744 1833
rect 6566 1765 6744 1799
rect 6566 1731 6570 1765
rect 6570 1731 6638 1765
rect 6638 1731 6672 1765
rect 6672 1731 6740 1765
rect 6740 1731 6744 1765
rect 6566 1697 6744 1731
rect 6566 1663 6570 1697
rect 6570 1663 6638 1697
rect 6638 1663 6672 1697
rect 6672 1663 6740 1697
rect 6740 1663 6744 1697
rect 6566 1629 6744 1663
rect 6566 1595 6570 1629
rect 6570 1595 6638 1629
rect 6638 1595 6672 1629
rect 6672 1595 6740 1629
rect 6740 1595 6744 1629
rect 6566 1561 6744 1595
rect 6566 1527 6570 1561
rect 6570 1527 6638 1561
rect 6638 1527 6672 1561
rect 6672 1527 6740 1561
rect 6740 1527 6744 1561
rect 6566 1491 6744 1527
rect 6566 1479 6600 1491
rect 6710 1479 6744 1491
rect 7313 4388 7419 4494
rect 7062 4028 7096 4062
rect 7134 4028 7168 4062
rect 7206 4028 7240 4062
rect 7062 3954 7096 3988
rect 7134 3954 7168 3988
rect 7206 3954 7240 3988
rect 7062 3880 7096 3914
rect 7134 3880 7168 3914
rect 7206 3880 7240 3914
rect 7062 3806 7096 3840
rect 7134 3806 7168 3840
rect 7206 3806 7240 3840
rect 7062 3732 7096 3766
rect 7134 3732 7168 3766
rect 7206 3732 7240 3766
rect 7062 3658 7096 3692
rect 7134 3658 7168 3692
rect 7206 3658 7240 3692
rect 7062 3584 7096 3618
rect 7134 3584 7168 3618
rect 7206 3584 7240 3618
rect 7062 3510 7096 3544
rect 7134 3510 7168 3544
rect 7206 3510 7240 3544
rect 7062 3436 7096 3470
rect 7134 3436 7168 3470
rect 7206 3436 7240 3470
rect 7062 3362 7096 3396
rect 7134 3362 7168 3396
rect 7206 3362 7240 3396
rect 7062 3288 7096 3322
rect 7134 3288 7168 3322
rect 7206 3288 7240 3322
rect 7062 3214 7096 3248
rect 7134 3214 7168 3248
rect 7206 3214 7240 3248
rect 7062 3140 7096 3174
rect 7134 3140 7168 3174
rect 7206 3140 7240 3174
rect 7062 3066 7096 3100
rect 7134 3066 7168 3100
rect 7206 3066 7240 3100
rect 7062 2992 7096 3026
rect 7134 2992 7168 3026
rect 7206 2992 7240 3026
rect 7062 2918 7096 2952
rect 7134 2918 7168 2952
rect 7206 2918 7240 2952
rect 7062 2844 7096 2878
rect 7134 2844 7168 2878
rect 7206 2844 7240 2878
rect 7062 2770 7096 2804
rect 7134 2770 7168 2804
rect 7206 2770 7240 2804
rect 7062 2696 7096 2730
rect 7134 2696 7168 2730
rect 7206 2696 7240 2730
rect 7062 2622 7096 2656
rect 7134 2622 7168 2656
rect 7206 2622 7240 2656
rect 7062 2548 7096 2582
rect 7134 2548 7168 2582
rect 7206 2548 7240 2582
rect 7062 2474 7096 2508
rect 7134 2474 7168 2508
rect 7206 2474 7240 2508
rect 7062 2400 7096 2434
rect 7134 2400 7168 2434
rect 7206 2400 7240 2434
rect 7062 2326 7096 2360
rect 7134 2326 7168 2360
rect 7206 2326 7240 2360
rect 7062 2252 7096 2286
rect 7134 2252 7168 2286
rect 7206 2252 7240 2286
rect 7062 2178 7096 2212
rect 7134 2178 7168 2212
rect 7206 2178 7240 2212
rect 7062 2104 7096 2138
rect 7134 2104 7168 2138
rect 7206 2104 7240 2138
rect 7062 2030 7096 2064
rect 7134 2030 7168 2064
rect 7206 2030 7240 2064
rect 7062 1956 7096 1990
rect 7134 1956 7168 1990
rect 7206 1956 7240 1990
rect 7062 1882 7096 1916
rect 7134 1882 7168 1916
rect 7206 1882 7240 1916
rect 7062 1808 7096 1842
rect 7134 1808 7168 1842
rect 7206 1808 7240 1842
rect 7062 1734 7096 1768
rect 7134 1734 7168 1768
rect 7206 1734 7240 1768
rect 7062 1660 7096 1694
rect 7134 1660 7168 1694
rect 7206 1660 7240 1694
rect 7062 1586 7096 1620
rect 7134 1586 7168 1620
rect 7206 1586 7240 1620
rect 7062 1511 7096 1545
rect 7134 1511 7168 1545
rect 7206 1511 7240 1545
rect 7875 4388 7981 4494
rect 7630 4050 7664 4062
rect 7558 4046 7736 4050
rect 7558 4012 7562 4046
rect 7562 4012 7630 4046
rect 7630 4012 7664 4046
rect 7664 4012 7732 4046
rect 7732 4012 7736 4046
rect 7558 3978 7736 4012
rect 7558 3944 7562 3978
rect 7562 3944 7630 3978
rect 7630 3944 7664 3978
rect 7664 3944 7732 3978
rect 7732 3944 7736 3978
rect 7558 3910 7736 3944
rect 7558 3876 7562 3910
rect 7562 3876 7630 3910
rect 7630 3876 7664 3910
rect 7664 3876 7732 3910
rect 7732 3876 7736 3910
rect 7558 3842 7736 3876
rect 7558 3808 7562 3842
rect 7562 3808 7630 3842
rect 7630 3808 7664 3842
rect 7664 3808 7732 3842
rect 7732 3808 7736 3842
rect 7558 3774 7736 3808
rect 7558 3740 7562 3774
rect 7562 3740 7630 3774
rect 7630 3740 7664 3774
rect 7664 3740 7732 3774
rect 7732 3740 7736 3774
rect 7558 3706 7736 3740
rect 7558 3672 7562 3706
rect 7562 3672 7630 3706
rect 7630 3672 7664 3706
rect 7664 3672 7732 3706
rect 7732 3672 7736 3706
rect 7558 3638 7736 3672
rect 7558 3604 7562 3638
rect 7562 3604 7630 3638
rect 7630 3604 7664 3638
rect 7664 3604 7732 3638
rect 7732 3604 7736 3638
rect 7558 3570 7736 3604
rect 7558 3536 7562 3570
rect 7562 3536 7630 3570
rect 7630 3536 7664 3570
rect 7664 3536 7732 3570
rect 7732 3536 7736 3570
rect 7558 3502 7736 3536
rect 7558 3468 7562 3502
rect 7562 3468 7630 3502
rect 7630 3468 7664 3502
rect 7664 3468 7732 3502
rect 7732 3468 7736 3502
rect 7558 3434 7736 3468
rect 7558 3400 7562 3434
rect 7562 3400 7630 3434
rect 7630 3400 7664 3434
rect 7664 3400 7732 3434
rect 7732 3400 7736 3434
rect 7558 3366 7736 3400
rect 7558 3332 7562 3366
rect 7562 3332 7630 3366
rect 7630 3332 7664 3366
rect 7664 3332 7732 3366
rect 7732 3332 7736 3366
rect 7558 3298 7736 3332
rect 7558 3264 7562 3298
rect 7562 3264 7630 3298
rect 7630 3264 7664 3298
rect 7664 3264 7732 3298
rect 7732 3264 7736 3298
rect 7558 3230 7736 3264
rect 7558 3196 7562 3230
rect 7562 3196 7630 3230
rect 7630 3196 7664 3230
rect 7664 3196 7732 3230
rect 7732 3196 7736 3230
rect 7558 3162 7736 3196
rect 7558 3128 7562 3162
rect 7562 3128 7630 3162
rect 7630 3128 7664 3162
rect 7664 3128 7732 3162
rect 7732 3128 7736 3162
rect 7558 3092 7736 3128
rect 7558 3080 7592 3092
rect 7702 3080 7736 3092
rect 7558 2935 7736 3040
rect 7558 2901 7597 2935
rect 7597 2901 7631 2935
rect 7631 2901 7665 2935
rect 7665 2901 7699 2935
rect 7699 2901 7736 2935
rect 7558 2855 7736 2901
rect 7558 2821 7597 2855
rect 7597 2821 7631 2855
rect 7631 2821 7665 2855
rect 7665 2821 7699 2855
rect 7699 2821 7736 2855
rect 7558 2775 7736 2821
rect 7558 2741 7597 2775
rect 7597 2741 7631 2775
rect 7631 2741 7665 2775
rect 7665 2741 7699 2775
rect 7699 2741 7736 2775
rect 7558 2695 7736 2741
rect 7558 2661 7597 2695
rect 7597 2661 7631 2695
rect 7631 2661 7665 2695
rect 7665 2661 7699 2695
rect 7699 2661 7736 2695
rect 7558 2614 7736 2661
rect 7558 2580 7597 2614
rect 7597 2580 7631 2614
rect 7631 2580 7665 2614
rect 7665 2580 7699 2614
rect 7699 2580 7736 2614
rect 7558 2574 7736 2580
rect 7558 2501 7592 2535
rect 7630 2501 7664 2535
rect 7702 2501 7736 2535
rect 7630 2449 7664 2461
rect 7558 2445 7736 2449
rect 7558 2411 7562 2445
rect 7562 2411 7630 2445
rect 7630 2411 7664 2445
rect 7664 2411 7732 2445
rect 7732 2411 7736 2445
rect 7558 2377 7736 2411
rect 7558 2343 7562 2377
rect 7562 2343 7630 2377
rect 7630 2343 7664 2377
rect 7664 2343 7732 2377
rect 7732 2343 7736 2377
rect 7558 2309 7736 2343
rect 7558 2275 7562 2309
rect 7562 2275 7630 2309
rect 7630 2275 7664 2309
rect 7664 2275 7732 2309
rect 7732 2275 7736 2309
rect 7558 2241 7736 2275
rect 7558 2207 7562 2241
rect 7562 2207 7630 2241
rect 7630 2207 7664 2241
rect 7664 2207 7732 2241
rect 7732 2207 7736 2241
rect 7558 2173 7736 2207
rect 7558 2139 7562 2173
rect 7562 2139 7630 2173
rect 7630 2139 7664 2173
rect 7664 2139 7732 2173
rect 7732 2139 7736 2173
rect 7558 2105 7736 2139
rect 7558 2071 7562 2105
rect 7562 2071 7630 2105
rect 7630 2071 7664 2105
rect 7664 2071 7732 2105
rect 7732 2071 7736 2105
rect 7558 2037 7736 2071
rect 7558 2003 7562 2037
rect 7562 2003 7630 2037
rect 7630 2003 7664 2037
rect 7664 2003 7732 2037
rect 7732 2003 7736 2037
rect 7558 1969 7736 2003
rect 7558 1935 7562 1969
rect 7562 1935 7630 1969
rect 7630 1935 7664 1969
rect 7664 1935 7732 1969
rect 7732 1935 7736 1969
rect 7558 1901 7736 1935
rect 7558 1867 7562 1901
rect 7562 1867 7630 1901
rect 7630 1867 7664 1901
rect 7664 1867 7732 1901
rect 7732 1867 7736 1901
rect 7558 1833 7736 1867
rect 7558 1799 7562 1833
rect 7562 1799 7630 1833
rect 7630 1799 7664 1833
rect 7664 1799 7732 1833
rect 7732 1799 7736 1833
rect 7558 1765 7736 1799
rect 7558 1731 7562 1765
rect 7562 1731 7630 1765
rect 7630 1731 7664 1765
rect 7664 1731 7732 1765
rect 7732 1731 7736 1765
rect 7558 1697 7736 1731
rect 7558 1663 7562 1697
rect 7562 1663 7630 1697
rect 7630 1663 7664 1697
rect 7664 1663 7732 1697
rect 7732 1663 7736 1697
rect 7558 1629 7736 1663
rect 7558 1595 7562 1629
rect 7562 1595 7630 1629
rect 7630 1595 7664 1629
rect 7664 1595 7732 1629
rect 7732 1595 7736 1629
rect 7558 1561 7736 1595
rect 7558 1527 7562 1561
rect 7562 1527 7630 1561
rect 7630 1527 7664 1561
rect 7664 1527 7732 1561
rect 7732 1527 7736 1561
rect 7558 1491 7736 1527
rect 7558 1479 7592 1491
rect 7702 1479 7736 1491
rect 8305 4388 8411 4494
rect 8054 4028 8088 4062
rect 8126 4028 8160 4062
rect 8198 4028 8232 4062
rect 8054 3954 8088 3988
rect 8126 3954 8160 3988
rect 8198 3954 8232 3988
rect 8054 3880 8088 3914
rect 8126 3880 8160 3914
rect 8198 3880 8232 3914
rect 8054 3806 8088 3840
rect 8126 3806 8160 3840
rect 8198 3806 8232 3840
rect 8054 3732 8088 3766
rect 8126 3732 8160 3766
rect 8198 3732 8232 3766
rect 8054 3658 8088 3692
rect 8126 3658 8160 3692
rect 8198 3658 8232 3692
rect 8054 3584 8088 3618
rect 8126 3584 8160 3618
rect 8198 3584 8232 3618
rect 8054 3510 8088 3544
rect 8126 3510 8160 3544
rect 8198 3510 8232 3544
rect 8054 3436 8088 3470
rect 8126 3436 8160 3470
rect 8198 3436 8232 3470
rect 8054 3362 8088 3396
rect 8126 3362 8160 3396
rect 8198 3362 8232 3396
rect 8054 3288 8088 3322
rect 8126 3288 8160 3322
rect 8198 3288 8232 3322
rect 8054 3214 8088 3248
rect 8126 3214 8160 3248
rect 8198 3214 8232 3248
rect 8054 3140 8088 3174
rect 8126 3140 8160 3174
rect 8198 3140 8232 3174
rect 8054 3066 8088 3100
rect 8126 3066 8160 3100
rect 8198 3066 8232 3100
rect 8054 2992 8088 3026
rect 8126 2992 8160 3026
rect 8198 2992 8232 3026
rect 8054 2918 8088 2952
rect 8126 2918 8160 2952
rect 8198 2918 8232 2952
rect 8054 2844 8088 2878
rect 8126 2844 8160 2878
rect 8198 2844 8232 2878
rect 8054 2770 8088 2804
rect 8126 2770 8160 2804
rect 8198 2770 8232 2804
rect 8054 2696 8088 2730
rect 8126 2696 8160 2730
rect 8198 2696 8232 2730
rect 8054 2622 8088 2656
rect 8126 2622 8160 2656
rect 8198 2622 8232 2656
rect 8054 2548 8088 2582
rect 8126 2548 8160 2582
rect 8198 2548 8232 2582
rect 8054 2474 8088 2508
rect 8126 2474 8160 2508
rect 8198 2474 8232 2508
rect 8054 2400 8088 2434
rect 8126 2400 8160 2434
rect 8198 2400 8232 2434
rect 8054 2326 8088 2360
rect 8126 2326 8160 2360
rect 8198 2326 8232 2360
rect 8054 2252 8088 2286
rect 8126 2252 8160 2286
rect 8198 2252 8232 2286
rect 8054 2178 8088 2212
rect 8126 2178 8160 2212
rect 8198 2178 8232 2212
rect 8054 2104 8088 2138
rect 8126 2104 8160 2138
rect 8198 2104 8232 2138
rect 8054 2030 8088 2064
rect 8126 2030 8160 2064
rect 8198 2030 8232 2064
rect 8054 1956 8088 1990
rect 8126 1956 8160 1990
rect 8198 1956 8232 1990
rect 8054 1882 8088 1916
rect 8126 1882 8160 1916
rect 8198 1882 8232 1916
rect 8054 1808 8088 1842
rect 8126 1808 8160 1842
rect 8198 1808 8232 1842
rect 8054 1734 8088 1768
rect 8126 1734 8160 1768
rect 8198 1734 8232 1768
rect 8054 1660 8088 1694
rect 8126 1660 8160 1694
rect 8198 1660 8232 1694
rect 8054 1586 8088 1620
rect 8126 1586 8160 1620
rect 8198 1586 8232 1620
rect 8054 1511 8088 1545
rect 8126 1511 8160 1545
rect 8198 1511 8232 1545
rect 8867 4388 8973 4494
rect 8622 4050 8656 4062
rect 8550 4046 8728 4050
rect 8550 4012 8554 4046
rect 8554 4012 8622 4046
rect 8622 4012 8656 4046
rect 8656 4012 8724 4046
rect 8724 4012 8728 4046
rect 8550 3978 8728 4012
rect 8550 3944 8554 3978
rect 8554 3944 8622 3978
rect 8622 3944 8656 3978
rect 8656 3944 8724 3978
rect 8724 3944 8728 3978
rect 8550 3910 8728 3944
rect 8550 3876 8554 3910
rect 8554 3876 8622 3910
rect 8622 3876 8656 3910
rect 8656 3876 8724 3910
rect 8724 3876 8728 3910
rect 8550 3842 8728 3876
rect 8550 3808 8554 3842
rect 8554 3808 8622 3842
rect 8622 3808 8656 3842
rect 8656 3808 8724 3842
rect 8724 3808 8728 3842
rect 8550 3774 8728 3808
rect 8550 3740 8554 3774
rect 8554 3740 8622 3774
rect 8622 3740 8656 3774
rect 8656 3740 8724 3774
rect 8724 3740 8728 3774
rect 8550 3706 8728 3740
rect 8550 3672 8554 3706
rect 8554 3672 8622 3706
rect 8622 3672 8656 3706
rect 8656 3672 8724 3706
rect 8724 3672 8728 3706
rect 8550 3638 8728 3672
rect 8550 3604 8554 3638
rect 8554 3604 8622 3638
rect 8622 3604 8656 3638
rect 8656 3604 8724 3638
rect 8724 3604 8728 3638
rect 8550 3570 8728 3604
rect 8550 3536 8554 3570
rect 8554 3536 8622 3570
rect 8622 3536 8656 3570
rect 8656 3536 8724 3570
rect 8724 3536 8728 3570
rect 8550 3502 8728 3536
rect 8550 3468 8554 3502
rect 8554 3468 8622 3502
rect 8622 3468 8656 3502
rect 8656 3468 8724 3502
rect 8724 3468 8728 3502
rect 8550 3434 8728 3468
rect 8550 3400 8554 3434
rect 8554 3400 8622 3434
rect 8622 3400 8656 3434
rect 8656 3400 8724 3434
rect 8724 3400 8728 3434
rect 8550 3366 8728 3400
rect 8550 3332 8554 3366
rect 8554 3332 8622 3366
rect 8622 3332 8656 3366
rect 8656 3332 8724 3366
rect 8724 3332 8728 3366
rect 8550 3298 8728 3332
rect 8550 3264 8554 3298
rect 8554 3264 8622 3298
rect 8622 3264 8656 3298
rect 8656 3264 8724 3298
rect 8724 3264 8728 3298
rect 8550 3230 8728 3264
rect 8550 3196 8554 3230
rect 8554 3196 8622 3230
rect 8622 3196 8656 3230
rect 8656 3196 8724 3230
rect 8724 3196 8728 3230
rect 8550 3162 8728 3196
rect 8550 3128 8554 3162
rect 8554 3128 8622 3162
rect 8622 3128 8656 3162
rect 8656 3128 8724 3162
rect 8724 3128 8728 3162
rect 8550 3092 8728 3128
rect 8550 3080 8584 3092
rect 8694 3080 8728 3092
rect 8550 2935 8728 3040
rect 8550 2901 8589 2935
rect 8589 2901 8623 2935
rect 8623 2901 8657 2935
rect 8657 2901 8691 2935
rect 8691 2901 8728 2935
rect 8550 2855 8728 2901
rect 8550 2821 8589 2855
rect 8589 2821 8623 2855
rect 8623 2821 8657 2855
rect 8657 2821 8691 2855
rect 8691 2821 8728 2855
rect 8550 2775 8728 2821
rect 8550 2741 8589 2775
rect 8589 2741 8623 2775
rect 8623 2741 8657 2775
rect 8657 2741 8691 2775
rect 8691 2741 8728 2775
rect 8550 2695 8728 2741
rect 8550 2661 8589 2695
rect 8589 2661 8623 2695
rect 8623 2661 8657 2695
rect 8657 2661 8691 2695
rect 8691 2661 8728 2695
rect 8550 2614 8728 2661
rect 8550 2580 8589 2614
rect 8589 2580 8623 2614
rect 8623 2580 8657 2614
rect 8657 2580 8691 2614
rect 8691 2580 8728 2614
rect 8550 2574 8728 2580
rect 8550 2501 8584 2535
rect 8622 2501 8656 2535
rect 8694 2501 8728 2535
rect 8622 2449 8656 2461
rect 8550 2445 8728 2449
rect 8550 2411 8554 2445
rect 8554 2411 8622 2445
rect 8622 2411 8656 2445
rect 8656 2411 8724 2445
rect 8724 2411 8728 2445
rect 8550 2377 8728 2411
rect 8550 2343 8554 2377
rect 8554 2343 8622 2377
rect 8622 2343 8656 2377
rect 8656 2343 8724 2377
rect 8724 2343 8728 2377
rect 8550 2309 8728 2343
rect 8550 2275 8554 2309
rect 8554 2275 8622 2309
rect 8622 2275 8656 2309
rect 8656 2275 8724 2309
rect 8724 2275 8728 2309
rect 8550 2241 8728 2275
rect 8550 2207 8554 2241
rect 8554 2207 8622 2241
rect 8622 2207 8656 2241
rect 8656 2207 8724 2241
rect 8724 2207 8728 2241
rect 8550 2173 8728 2207
rect 8550 2139 8554 2173
rect 8554 2139 8622 2173
rect 8622 2139 8656 2173
rect 8656 2139 8724 2173
rect 8724 2139 8728 2173
rect 8550 2105 8728 2139
rect 8550 2071 8554 2105
rect 8554 2071 8622 2105
rect 8622 2071 8656 2105
rect 8656 2071 8724 2105
rect 8724 2071 8728 2105
rect 8550 2037 8728 2071
rect 8550 2003 8554 2037
rect 8554 2003 8622 2037
rect 8622 2003 8656 2037
rect 8656 2003 8724 2037
rect 8724 2003 8728 2037
rect 8550 1969 8728 2003
rect 8550 1935 8554 1969
rect 8554 1935 8622 1969
rect 8622 1935 8656 1969
rect 8656 1935 8724 1969
rect 8724 1935 8728 1969
rect 8550 1901 8728 1935
rect 8550 1867 8554 1901
rect 8554 1867 8622 1901
rect 8622 1867 8656 1901
rect 8656 1867 8724 1901
rect 8724 1867 8728 1901
rect 8550 1833 8728 1867
rect 8550 1799 8554 1833
rect 8554 1799 8622 1833
rect 8622 1799 8656 1833
rect 8656 1799 8724 1833
rect 8724 1799 8728 1833
rect 8550 1765 8728 1799
rect 8550 1731 8554 1765
rect 8554 1731 8622 1765
rect 8622 1731 8656 1765
rect 8656 1731 8724 1765
rect 8724 1731 8728 1765
rect 8550 1697 8728 1731
rect 8550 1663 8554 1697
rect 8554 1663 8622 1697
rect 8622 1663 8656 1697
rect 8656 1663 8724 1697
rect 8724 1663 8728 1697
rect 8550 1629 8728 1663
rect 8550 1595 8554 1629
rect 8554 1595 8622 1629
rect 8622 1595 8656 1629
rect 8656 1595 8724 1629
rect 8724 1595 8728 1629
rect 8550 1561 8728 1595
rect 8550 1527 8554 1561
rect 8554 1527 8622 1561
rect 8622 1527 8656 1561
rect 8656 1527 8724 1561
rect 8724 1527 8728 1561
rect 8550 1491 8728 1527
rect 8550 1479 8584 1491
rect 8694 1479 8728 1491
rect 9297 4388 9403 4494
rect 9046 4028 9080 4062
rect 9118 4028 9152 4062
rect 9190 4028 9224 4062
rect 9046 3954 9080 3988
rect 9118 3954 9152 3988
rect 9190 3954 9224 3988
rect 9046 3880 9080 3914
rect 9118 3880 9152 3914
rect 9190 3880 9224 3914
rect 9046 3806 9080 3840
rect 9118 3806 9152 3840
rect 9190 3806 9224 3840
rect 9046 3732 9080 3766
rect 9118 3732 9152 3766
rect 9190 3732 9224 3766
rect 9046 3658 9080 3692
rect 9118 3658 9152 3692
rect 9190 3658 9224 3692
rect 9046 3584 9080 3618
rect 9118 3584 9152 3618
rect 9190 3584 9224 3618
rect 9046 3510 9080 3544
rect 9118 3510 9152 3544
rect 9190 3510 9224 3544
rect 9046 3436 9080 3470
rect 9118 3436 9152 3470
rect 9190 3436 9224 3470
rect 9046 3362 9080 3396
rect 9118 3362 9152 3396
rect 9190 3362 9224 3396
rect 9046 3288 9080 3322
rect 9118 3288 9152 3322
rect 9190 3288 9224 3322
rect 9046 3214 9080 3248
rect 9118 3214 9152 3248
rect 9190 3214 9224 3248
rect 9046 3140 9080 3174
rect 9118 3140 9152 3174
rect 9190 3140 9224 3174
rect 9046 3066 9080 3100
rect 9118 3066 9152 3100
rect 9190 3066 9224 3100
rect 9046 2992 9080 3026
rect 9118 2992 9152 3026
rect 9190 2992 9224 3026
rect 9046 2918 9080 2952
rect 9118 2918 9152 2952
rect 9190 2918 9224 2952
rect 9046 2844 9080 2878
rect 9118 2844 9152 2878
rect 9190 2844 9224 2878
rect 9046 2770 9080 2804
rect 9118 2770 9152 2804
rect 9190 2770 9224 2804
rect 9046 2696 9080 2730
rect 9118 2696 9152 2730
rect 9190 2696 9224 2730
rect 9046 2622 9080 2656
rect 9118 2622 9152 2656
rect 9190 2622 9224 2656
rect 9046 2548 9080 2582
rect 9118 2548 9152 2582
rect 9190 2548 9224 2582
rect 9046 2474 9080 2508
rect 9118 2474 9152 2508
rect 9190 2474 9224 2508
rect 9046 2400 9080 2434
rect 9118 2400 9152 2434
rect 9190 2400 9224 2434
rect 9046 2326 9080 2360
rect 9118 2326 9152 2360
rect 9190 2326 9224 2360
rect 9046 2252 9080 2286
rect 9118 2252 9152 2286
rect 9190 2252 9224 2286
rect 9046 2178 9080 2212
rect 9118 2178 9152 2212
rect 9190 2178 9224 2212
rect 9046 2104 9080 2138
rect 9118 2104 9152 2138
rect 9190 2104 9224 2138
rect 9046 2030 9080 2064
rect 9118 2030 9152 2064
rect 9190 2030 9224 2064
rect 9046 1956 9080 1990
rect 9118 1956 9152 1990
rect 9190 1956 9224 1990
rect 9046 1882 9080 1916
rect 9118 1882 9152 1916
rect 9190 1882 9224 1916
rect 9046 1808 9080 1842
rect 9118 1808 9152 1842
rect 9190 1808 9224 1842
rect 9046 1734 9080 1768
rect 9118 1734 9152 1768
rect 9190 1734 9224 1768
rect 9046 1660 9080 1694
rect 9118 1660 9152 1694
rect 9190 1660 9224 1694
rect 9046 1586 9080 1620
rect 9118 1586 9152 1620
rect 9190 1586 9224 1620
rect 9046 1511 9080 1545
rect 9118 1511 9152 1545
rect 9190 1511 9224 1545
rect 9859 4388 9965 4494
rect 9614 4050 9648 4062
rect 9542 4046 9720 4050
rect 9542 4012 9546 4046
rect 9546 4012 9614 4046
rect 9614 4012 9648 4046
rect 9648 4012 9716 4046
rect 9716 4012 9720 4046
rect 9542 3978 9720 4012
rect 9542 3944 9546 3978
rect 9546 3944 9614 3978
rect 9614 3944 9648 3978
rect 9648 3944 9716 3978
rect 9716 3944 9720 3978
rect 9542 3910 9720 3944
rect 9542 3876 9546 3910
rect 9546 3876 9614 3910
rect 9614 3876 9648 3910
rect 9648 3876 9716 3910
rect 9716 3876 9720 3910
rect 9542 3842 9720 3876
rect 9542 3808 9546 3842
rect 9546 3808 9614 3842
rect 9614 3808 9648 3842
rect 9648 3808 9716 3842
rect 9716 3808 9720 3842
rect 9542 3774 9720 3808
rect 9542 3740 9546 3774
rect 9546 3740 9614 3774
rect 9614 3740 9648 3774
rect 9648 3740 9716 3774
rect 9716 3740 9720 3774
rect 9542 3706 9720 3740
rect 9542 3672 9546 3706
rect 9546 3672 9614 3706
rect 9614 3672 9648 3706
rect 9648 3672 9716 3706
rect 9716 3672 9720 3706
rect 9542 3638 9720 3672
rect 9542 3604 9546 3638
rect 9546 3604 9614 3638
rect 9614 3604 9648 3638
rect 9648 3604 9716 3638
rect 9716 3604 9720 3638
rect 9542 3570 9720 3604
rect 9542 3536 9546 3570
rect 9546 3536 9614 3570
rect 9614 3536 9648 3570
rect 9648 3536 9716 3570
rect 9716 3536 9720 3570
rect 9542 3502 9720 3536
rect 9542 3468 9546 3502
rect 9546 3468 9614 3502
rect 9614 3468 9648 3502
rect 9648 3468 9716 3502
rect 9716 3468 9720 3502
rect 9542 3434 9720 3468
rect 9542 3400 9546 3434
rect 9546 3400 9614 3434
rect 9614 3400 9648 3434
rect 9648 3400 9716 3434
rect 9716 3400 9720 3434
rect 9542 3366 9720 3400
rect 9542 3332 9546 3366
rect 9546 3332 9614 3366
rect 9614 3332 9648 3366
rect 9648 3332 9716 3366
rect 9716 3332 9720 3366
rect 9542 3298 9720 3332
rect 9542 3264 9546 3298
rect 9546 3264 9614 3298
rect 9614 3264 9648 3298
rect 9648 3264 9716 3298
rect 9716 3264 9720 3298
rect 9542 3230 9720 3264
rect 9542 3196 9546 3230
rect 9546 3196 9614 3230
rect 9614 3196 9648 3230
rect 9648 3196 9716 3230
rect 9716 3196 9720 3230
rect 9542 3162 9720 3196
rect 9542 3128 9546 3162
rect 9546 3128 9614 3162
rect 9614 3128 9648 3162
rect 9648 3128 9716 3162
rect 9716 3128 9720 3162
rect 9542 3092 9720 3128
rect 9542 3080 9576 3092
rect 9686 3080 9720 3092
rect 9542 2935 9720 3040
rect 9542 2901 9581 2935
rect 9581 2901 9615 2935
rect 9615 2901 9649 2935
rect 9649 2901 9683 2935
rect 9683 2901 9720 2935
rect 9542 2855 9720 2901
rect 9542 2821 9581 2855
rect 9581 2821 9615 2855
rect 9615 2821 9649 2855
rect 9649 2821 9683 2855
rect 9683 2821 9720 2855
rect 9542 2775 9720 2821
rect 9542 2741 9581 2775
rect 9581 2741 9615 2775
rect 9615 2741 9649 2775
rect 9649 2741 9683 2775
rect 9683 2741 9720 2775
rect 9542 2695 9720 2741
rect 9542 2661 9581 2695
rect 9581 2661 9615 2695
rect 9615 2661 9649 2695
rect 9649 2661 9683 2695
rect 9683 2661 9720 2695
rect 9542 2614 9720 2661
rect 9542 2580 9581 2614
rect 9581 2580 9615 2614
rect 9615 2580 9649 2614
rect 9649 2580 9683 2614
rect 9683 2580 9720 2614
rect 9542 2574 9720 2580
rect 9542 2501 9576 2535
rect 9614 2501 9648 2535
rect 9686 2501 9720 2535
rect 9614 2449 9648 2461
rect 9542 2445 9720 2449
rect 9542 2411 9546 2445
rect 9546 2411 9614 2445
rect 9614 2411 9648 2445
rect 9648 2411 9716 2445
rect 9716 2411 9720 2445
rect 9542 2377 9720 2411
rect 9542 2343 9546 2377
rect 9546 2343 9614 2377
rect 9614 2343 9648 2377
rect 9648 2343 9716 2377
rect 9716 2343 9720 2377
rect 9542 2309 9720 2343
rect 9542 2275 9546 2309
rect 9546 2275 9614 2309
rect 9614 2275 9648 2309
rect 9648 2275 9716 2309
rect 9716 2275 9720 2309
rect 9542 2241 9720 2275
rect 9542 2207 9546 2241
rect 9546 2207 9614 2241
rect 9614 2207 9648 2241
rect 9648 2207 9716 2241
rect 9716 2207 9720 2241
rect 9542 2173 9720 2207
rect 9542 2139 9546 2173
rect 9546 2139 9614 2173
rect 9614 2139 9648 2173
rect 9648 2139 9716 2173
rect 9716 2139 9720 2173
rect 9542 2105 9720 2139
rect 9542 2071 9546 2105
rect 9546 2071 9614 2105
rect 9614 2071 9648 2105
rect 9648 2071 9716 2105
rect 9716 2071 9720 2105
rect 9542 2037 9720 2071
rect 9542 2003 9546 2037
rect 9546 2003 9614 2037
rect 9614 2003 9648 2037
rect 9648 2003 9716 2037
rect 9716 2003 9720 2037
rect 9542 1969 9720 2003
rect 9542 1935 9546 1969
rect 9546 1935 9614 1969
rect 9614 1935 9648 1969
rect 9648 1935 9716 1969
rect 9716 1935 9720 1969
rect 9542 1901 9720 1935
rect 9542 1867 9546 1901
rect 9546 1867 9614 1901
rect 9614 1867 9648 1901
rect 9648 1867 9716 1901
rect 9716 1867 9720 1901
rect 9542 1833 9720 1867
rect 9542 1799 9546 1833
rect 9546 1799 9614 1833
rect 9614 1799 9648 1833
rect 9648 1799 9716 1833
rect 9716 1799 9720 1833
rect 9542 1765 9720 1799
rect 9542 1731 9546 1765
rect 9546 1731 9614 1765
rect 9614 1731 9648 1765
rect 9648 1731 9716 1765
rect 9716 1731 9720 1765
rect 9542 1697 9720 1731
rect 9542 1663 9546 1697
rect 9546 1663 9614 1697
rect 9614 1663 9648 1697
rect 9648 1663 9716 1697
rect 9716 1663 9720 1697
rect 9542 1629 9720 1663
rect 9542 1595 9546 1629
rect 9546 1595 9614 1629
rect 9614 1595 9648 1629
rect 9648 1595 9716 1629
rect 9716 1595 9720 1629
rect 9542 1561 9720 1595
rect 9542 1527 9546 1561
rect 9546 1527 9614 1561
rect 9614 1527 9648 1561
rect 9648 1527 9716 1561
rect 9716 1527 9720 1561
rect 9542 1491 9720 1527
rect 9542 1479 9576 1491
rect 9686 1479 9720 1491
rect 10289 4388 10395 4494
rect 10038 4028 10072 4062
rect 10110 4028 10144 4062
rect 10182 4028 10216 4062
rect 10038 3954 10072 3988
rect 10110 3954 10144 3988
rect 10182 3954 10216 3988
rect 10038 3880 10072 3914
rect 10110 3880 10144 3914
rect 10182 3880 10216 3914
rect 10038 3806 10072 3840
rect 10110 3806 10144 3840
rect 10182 3806 10216 3840
rect 10038 3732 10072 3766
rect 10110 3732 10144 3766
rect 10182 3732 10216 3766
rect 10038 3658 10072 3692
rect 10110 3658 10144 3692
rect 10182 3658 10216 3692
rect 10038 3584 10072 3618
rect 10110 3584 10144 3618
rect 10182 3584 10216 3618
rect 10038 3510 10072 3544
rect 10110 3510 10144 3544
rect 10182 3510 10216 3544
rect 10038 3436 10072 3470
rect 10110 3436 10144 3470
rect 10182 3436 10216 3470
rect 10038 3362 10072 3396
rect 10110 3362 10144 3396
rect 10182 3362 10216 3396
rect 10038 3288 10072 3322
rect 10110 3288 10144 3322
rect 10182 3288 10216 3322
rect 10038 3214 10072 3248
rect 10110 3214 10144 3248
rect 10182 3214 10216 3248
rect 10038 3140 10072 3174
rect 10110 3140 10144 3174
rect 10182 3140 10216 3174
rect 10038 3066 10072 3100
rect 10110 3066 10144 3100
rect 10182 3066 10216 3100
rect 10038 2992 10072 3026
rect 10110 2992 10144 3026
rect 10182 2992 10216 3026
rect 10038 2918 10072 2952
rect 10110 2918 10144 2952
rect 10182 2918 10216 2952
rect 10038 2844 10072 2878
rect 10110 2844 10144 2878
rect 10182 2844 10216 2878
rect 10038 2770 10072 2804
rect 10110 2770 10144 2804
rect 10182 2770 10216 2804
rect 10038 2696 10072 2730
rect 10110 2696 10144 2730
rect 10182 2696 10216 2730
rect 10038 2622 10072 2656
rect 10110 2622 10144 2656
rect 10182 2622 10216 2656
rect 10038 2548 10072 2582
rect 10110 2548 10144 2582
rect 10182 2548 10216 2582
rect 10038 2474 10072 2508
rect 10110 2474 10144 2508
rect 10182 2474 10216 2508
rect 10038 2400 10072 2434
rect 10110 2400 10144 2434
rect 10182 2400 10216 2434
rect 10038 2326 10072 2360
rect 10110 2326 10144 2360
rect 10182 2326 10216 2360
rect 10038 2252 10072 2286
rect 10110 2252 10144 2286
rect 10182 2252 10216 2286
rect 10038 2178 10072 2212
rect 10110 2178 10144 2212
rect 10182 2178 10216 2212
rect 10038 2104 10072 2138
rect 10110 2104 10144 2138
rect 10182 2104 10216 2138
rect 10038 2030 10072 2064
rect 10110 2030 10144 2064
rect 10182 2030 10216 2064
rect 10038 1956 10072 1990
rect 10110 1956 10144 1990
rect 10182 1956 10216 1990
rect 10038 1882 10072 1916
rect 10110 1882 10144 1916
rect 10182 1882 10216 1916
rect 10038 1808 10072 1842
rect 10110 1808 10144 1842
rect 10182 1808 10216 1842
rect 10038 1734 10072 1768
rect 10110 1734 10144 1768
rect 10182 1734 10216 1768
rect 10038 1660 10072 1694
rect 10110 1660 10144 1694
rect 10182 1660 10216 1694
rect 10038 1586 10072 1620
rect 10110 1586 10144 1620
rect 10182 1586 10216 1620
rect 10038 1511 10072 1545
rect 10110 1511 10144 1545
rect 10182 1511 10216 1545
rect 10851 4388 10957 4494
rect 10606 4050 10640 4062
rect 10534 4046 10712 4050
rect 10534 4012 10538 4046
rect 10538 4012 10606 4046
rect 10606 4012 10640 4046
rect 10640 4012 10708 4046
rect 10708 4012 10712 4046
rect 10534 3978 10712 4012
rect 10534 3944 10538 3978
rect 10538 3944 10606 3978
rect 10606 3944 10640 3978
rect 10640 3944 10708 3978
rect 10708 3944 10712 3978
rect 10534 3910 10712 3944
rect 10534 3876 10538 3910
rect 10538 3876 10606 3910
rect 10606 3876 10640 3910
rect 10640 3876 10708 3910
rect 10708 3876 10712 3910
rect 10534 3842 10712 3876
rect 10534 3808 10538 3842
rect 10538 3808 10606 3842
rect 10606 3808 10640 3842
rect 10640 3808 10708 3842
rect 10708 3808 10712 3842
rect 10534 3774 10712 3808
rect 10534 3740 10538 3774
rect 10538 3740 10606 3774
rect 10606 3740 10640 3774
rect 10640 3740 10708 3774
rect 10708 3740 10712 3774
rect 10534 3706 10712 3740
rect 10534 3672 10538 3706
rect 10538 3672 10606 3706
rect 10606 3672 10640 3706
rect 10640 3672 10708 3706
rect 10708 3672 10712 3706
rect 10534 3638 10712 3672
rect 10534 3604 10538 3638
rect 10538 3604 10606 3638
rect 10606 3604 10640 3638
rect 10640 3604 10708 3638
rect 10708 3604 10712 3638
rect 10534 3570 10712 3604
rect 10534 3536 10538 3570
rect 10538 3536 10606 3570
rect 10606 3536 10640 3570
rect 10640 3536 10708 3570
rect 10708 3536 10712 3570
rect 10534 3502 10712 3536
rect 10534 3468 10538 3502
rect 10538 3468 10606 3502
rect 10606 3468 10640 3502
rect 10640 3468 10708 3502
rect 10708 3468 10712 3502
rect 10534 3434 10712 3468
rect 10534 3400 10538 3434
rect 10538 3400 10606 3434
rect 10606 3400 10640 3434
rect 10640 3400 10708 3434
rect 10708 3400 10712 3434
rect 10534 3366 10712 3400
rect 10534 3332 10538 3366
rect 10538 3332 10606 3366
rect 10606 3332 10640 3366
rect 10640 3332 10708 3366
rect 10708 3332 10712 3366
rect 10534 3298 10712 3332
rect 10534 3264 10538 3298
rect 10538 3264 10606 3298
rect 10606 3264 10640 3298
rect 10640 3264 10708 3298
rect 10708 3264 10712 3298
rect 10534 3230 10712 3264
rect 10534 3196 10538 3230
rect 10538 3196 10606 3230
rect 10606 3196 10640 3230
rect 10640 3196 10708 3230
rect 10708 3196 10712 3230
rect 10534 3162 10712 3196
rect 10534 3128 10538 3162
rect 10538 3128 10606 3162
rect 10606 3128 10640 3162
rect 10640 3128 10708 3162
rect 10708 3128 10712 3162
rect 10534 3092 10712 3128
rect 10534 3080 10568 3092
rect 10678 3080 10712 3092
rect 10534 3003 10568 3037
rect 10606 3003 10640 3037
rect 10678 3003 10712 3037
rect 10534 2920 10568 2954
rect 10606 2935 10640 2954
rect 10606 2920 10607 2935
rect 10607 2920 10640 2935
rect 10678 2920 10712 2954
rect 10534 2837 10568 2871
rect 10606 2855 10640 2871
rect 10606 2837 10607 2855
rect 10607 2837 10640 2855
rect 10678 2837 10712 2871
rect 10534 2753 10568 2787
rect 10606 2775 10640 2787
rect 10606 2753 10607 2775
rect 10607 2753 10640 2775
rect 10678 2753 10712 2787
rect 10534 2669 10568 2703
rect 10606 2695 10640 2703
rect 10606 2669 10607 2695
rect 10607 2669 10640 2695
rect 10678 2669 10712 2703
rect 10534 2585 10568 2619
rect 10606 2614 10640 2619
rect 10606 2585 10607 2614
rect 10607 2585 10640 2614
rect 10678 2585 10712 2619
rect 10534 2501 10568 2535
rect 10606 2501 10640 2535
rect 10678 2501 10712 2535
rect 10606 2449 10640 2461
rect 10534 2445 10712 2449
rect 10534 2411 10538 2445
rect 10538 2411 10606 2445
rect 10606 2411 10640 2445
rect 10640 2411 10708 2445
rect 10708 2411 10712 2445
rect 10534 2377 10712 2411
rect 10534 2343 10538 2377
rect 10538 2343 10606 2377
rect 10606 2343 10640 2377
rect 10640 2343 10708 2377
rect 10708 2343 10712 2377
rect 10534 2309 10712 2343
rect 10534 2275 10538 2309
rect 10538 2275 10606 2309
rect 10606 2275 10640 2309
rect 10640 2275 10708 2309
rect 10708 2275 10712 2309
rect 10534 2241 10712 2275
rect 10534 2207 10538 2241
rect 10538 2207 10606 2241
rect 10606 2207 10640 2241
rect 10640 2207 10708 2241
rect 10708 2207 10712 2241
rect 10534 2173 10712 2207
rect 10534 2139 10538 2173
rect 10538 2139 10606 2173
rect 10606 2139 10640 2173
rect 10640 2139 10708 2173
rect 10708 2139 10712 2173
rect 10534 2105 10712 2139
rect 10534 2071 10538 2105
rect 10538 2071 10606 2105
rect 10606 2071 10640 2105
rect 10640 2071 10708 2105
rect 10708 2071 10712 2105
rect 10534 2037 10712 2071
rect 10534 2003 10538 2037
rect 10538 2003 10606 2037
rect 10606 2003 10640 2037
rect 10640 2003 10708 2037
rect 10708 2003 10712 2037
rect 10534 1969 10712 2003
rect 10534 1935 10538 1969
rect 10538 1935 10606 1969
rect 10606 1935 10640 1969
rect 10640 1935 10708 1969
rect 10708 1935 10712 1969
rect 10534 1901 10712 1935
rect 10534 1867 10538 1901
rect 10538 1867 10606 1901
rect 10606 1867 10640 1901
rect 10640 1867 10708 1901
rect 10708 1867 10712 1901
rect 10534 1833 10712 1867
rect 10534 1799 10538 1833
rect 10538 1799 10606 1833
rect 10606 1799 10640 1833
rect 10640 1799 10708 1833
rect 10708 1799 10712 1833
rect 10534 1765 10712 1799
rect 10534 1731 10538 1765
rect 10538 1731 10606 1765
rect 10606 1731 10640 1765
rect 10640 1731 10708 1765
rect 10708 1731 10712 1765
rect 10534 1697 10712 1731
rect 10534 1663 10538 1697
rect 10538 1663 10606 1697
rect 10606 1663 10640 1697
rect 10640 1663 10708 1697
rect 10708 1663 10712 1697
rect 10534 1629 10712 1663
rect 10534 1595 10538 1629
rect 10538 1595 10606 1629
rect 10606 1595 10640 1629
rect 10640 1595 10708 1629
rect 10708 1595 10712 1629
rect 10534 1561 10712 1595
rect 10534 1527 10538 1561
rect 10538 1527 10606 1561
rect 10606 1527 10640 1561
rect 10640 1527 10708 1561
rect 10708 1527 10712 1561
rect 10534 1491 10712 1527
rect 10534 1479 10568 1491
rect 10678 1479 10712 1491
rect 11281 4388 11387 4494
rect 11030 4028 11064 4062
rect 11102 4028 11136 4062
rect 11174 4028 11208 4062
rect 11030 3954 11064 3988
rect 11102 3954 11136 3988
rect 11174 3954 11208 3988
rect 11030 3880 11064 3914
rect 11102 3880 11136 3914
rect 11174 3880 11208 3914
rect 11030 3806 11064 3840
rect 11102 3806 11136 3840
rect 11174 3806 11208 3840
rect 11030 3732 11064 3766
rect 11102 3732 11136 3766
rect 11174 3732 11208 3766
rect 11030 3658 11064 3692
rect 11102 3658 11136 3692
rect 11174 3658 11208 3692
rect 11030 3584 11064 3618
rect 11102 3584 11136 3618
rect 11174 3584 11208 3618
rect 11030 3510 11064 3544
rect 11102 3510 11136 3544
rect 11174 3510 11208 3544
rect 11030 3436 11064 3470
rect 11102 3436 11136 3470
rect 11174 3436 11208 3470
rect 11030 3362 11064 3396
rect 11102 3362 11136 3396
rect 11174 3362 11208 3396
rect 11030 3288 11064 3322
rect 11102 3288 11136 3322
rect 11174 3288 11208 3322
rect 11030 3214 11064 3248
rect 11102 3214 11136 3248
rect 11174 3214 11208 3248
rect 11030 3140 11064 3174
rect 11102 3140 11136 3174
rect 11174 3140 11208 3174
rect 11030 3066 11064 3100
rect 11102 3066 11136 3100
rect 11174 3066 11208 3100
rect 11030 2992 11064 3026
rect 11102 2992 11136 3026
rect 11174 2992 11208 3026
rect 11030 2918 11064 2952
rect 11102 2918 11136 2952
rect 11174 2918 11208 2952
rect 11030 2844 11064 2878
rect 11102 2844 11136 2878
rect 11174 2844 11208 2878
rect 11030 2770 11064 2804
rect 11102 2770 11136 2804
rect 11174 2770 11208 2804
rect 11030 2696 11064 2730
rect 11102 2696 11136 2730
rect 11174 2696 11208 2730
rect 11030 2622 11064 2656
rect 11102 2622 11136 2656
rect 11174 2622 11208 2656
rect 11030 2548 11064 2582
rect 11102 2548 11136 2582
rect 11174 2548 11208 2582
rect 11030 2474 11064 2508
rect 11102 2474 11136 2508
rect 11174 2474 11208 2508
rect 11030 2400 11064 2434
rect 11102 2400 11136 2434
rect 11174 2400 11208 2434
rect 11030 2326 11064 2360
rect 11102 2326 11136 2360
rect 11174 2326 11208 2360
rect 11030 2252 11064 2286
rect 11102 2252 11136 2286
rect 11174 2252 11208 2286
rect 11030 2178 11064 2212
rect 11102 2178 11136 2212
rect 11174 2178 11208 2212
rect 11030 2104 11064 2138
rect 11102 2104 11136 2138
rect 11174 2104 11208 2138
rect 11030 2030 11064 2064
rect 11102 2030 11136 2064
rect 11174 2030 11208 2064
rect 11030 1956 11064 1990
rect 11102 1956 11136 1990
rect 11174 1956 11208 1990
rect 11030 1882 11064 1916
rect 11102 1882 11136 1916
rect 11174 1882 11208 1916
rect 11030 1808 11064 1842
rect 11102 1808 11136 1842
rect 11174 1808 11208 1842
rect 11030 1734 11064 1768
rect 11102 1734 11136 1768
rect 11174 1734 11208 1768
rect 11030 1660 11064 1694
rect 11102 1660 11136 1694
rect 11174 1660 11208 1694
rect 11030 1586 11064 1620
rect 11102 1586 11136 1620
rect 11174 1586 11208 1620
rect 11030 1511 11064 1545
rect 11102 1511 11136 1545
rect 11174 1511 11208 1545
rect 11843 4388 11949 4494
rect 11598 4050 11632 4062
rect 11526 4046 11704 4050
rect 11526 4012 11530 4046
rect 11530 4012 11598 4046
rect 11598 4012 11632 4046
rect 11632 4012 11700 4046
rect 11700 4012 11704 4046
rect 11526 3978 11704 4012
rect 11526 3944 11530 3978
rect 11530 3944 11598 3978
rect 11598 3944 11632 3978
rect 11632 3944 11700 3978
rect 11700 3944 11704 3978
rect 11526 3910 11704 3944
rect 11526 3876 11530 3910
rect 11530 3876 11598 3910
rect 11598 3876 11632 3910
rect 11632 3876 11700 3910
rect 11700 3876 11704 3910
rect 11526 3842 11704 3876
rect 11526 3808 11530 3842
rect 11530 3808 11598 3842
rect 11598 3808 11632 3842
rect 11632 3808 11700 3842
rect 11700 3808 11704 3842
rect 11526 3774 11704 3808
rect 11526 3740 11530 3774
rect 11530 3740 11598 3774
rect 11598 3740 11632 3774
rect 11632 3740 11700 3774
rect 11700 3740 11704 3774
rect 11526 3706 11704 3740
rect 11526 3672 11530 3706
rect 11530 3672 11598 3706
rect 11598 3672 11632 3706
rect 11632 3672 11700 3706
rect 11700 3672 11704 3706
rect 11526 3638 11704 3672
rect 11526 3604 11530 3638
rect 11530 3604 11598 3638
rect 11598 3604 11632 3638
rect 11632 3604 11700 3638
rect 11700 3604 11704 3638
rect 11526 3570 11704 3604
rect 11526 3536 11530 3570
rect 11530 3536 11598 3570
rect 11598 3536 11632 3570
rect 11632 3536 11700 3570
rect 11700 3536 11704 3570
rect 11526 3502 11704 3536
rect 11526 3468 11530 3502
rect 11530 3468 11598 3502
rect 11598 3468 11632 3502
rect 11632 3468 11700 3502
rect 11700 3468 11704 3502
rect 11526 3434 11704 3468
rect 11526 3400 11530 3434
rect 11530 3400 11598 3434
rect 11598 3400 11632 3434
rect 11632 3400 11700 3434
rect 11700 3400 11704 3434
rect 11526 3366 11704 3400
rect 11526 3332 11530 3366
rect 11530 3332 11598 3366
rect 11598 3332 11632 3366
rect 11632 3332 11700 3366
rect 11700 3332 11704 3366
rect 11526 3298 11704 3332
rect 11526 3264 11530 3298
rect 11530 3264 11598 3298
rect 11598 3264 11632 3298
rect 11632 3264 11700 3298
rect 11700 3264 11704 3298
rect 11526 3230 11704 3264
rect 11526 3196 11530 3230
rect 11530 3196 11598 3230
rect 11598 3196 11632 3230
rect 11632 3196 11700 3230
rect 11700 3196 11704 3230
rect 11526 3162 11704 3196
rect 11526 3128 11530 3162
rect 11530 3128 11598 3162
rect 11598 3128 11632 3162
rect 11632 3128 11700 3162
rect 11700 3128 11704 3162
rect 11526 3092 11704 3128
rect 11526 3080 11560 3092
rect 11670 3080 11704 3092
rect 11526 3003 11560 3037
rect 11598 3003 11632 3037
rect 11670 3003 11704 3037
rect 11526 2920 11560 2954
rect 11598 2935 11632 2954
rect 11598 2920 11599 2935
rect 11599 2920 11632 2935
rect 11670 2920 11704 2954
rect 11526 2837 11560 2871
rect 11598 2855 11632 2871
rect 11598 2837 11599 2855
rect 11599 2837 11632 2855
rect 11670 2837 11704 2871
rect 11526 2753 11560 2787
rect 11598 2775 11632 2787
rect 11598 2753 11599 2775
rect 11599 2753 11632 2775
rect 11670 2753 11704 2787
rect 11526 2669 11560 2703
rect 11598 2695 11632 2703
rect 11598 2669 11599 2695
rect 11599 2669 11632 2695
rect 11670 2669 11704 2703
rect 11526 2585 11560 2619
rect 11598 2614 11632 2619
rect 11598 2585 11599 2614
rect 11599 2585 11632 2614
rect 11670 2585 11704 2619
rect 11526 2501 11560 2535
rect 11598 2501 11632 2535
rect 11670 2501 11704 2535
rect 11598 2449 11632 2461
rect 11526 2445 11704 2449
rect 11526 2411 11530 2445
rect 11530 2411 11598 2445
rect 11598 2411 11632 2445
rect 11632 2411 11700 2445
rect 11700 2411 11704 2445
rect 11526 2377 11704 2411
rect 11526 2343 11530 2377
rect 11530 2343 11598 2377
rect 11598 2343 11632 2377
rect 11632 2343 11700 2377
rect 11700 2343 11704 2377
rect 11526 2309 11704 2343
rect 11526 2275 11530 2309
rect 11530 2275 11598 2309
rect 11598 2275 11632 2309
rect 11632 2275 11700 2309
rect 11700 2275 11704 2309
rect 11526 2241 11704 2275
rect 11526 2207 11530 2241
rect 11530 2207 11598 2241
rect 11598 2207 11632 2241
rect 11632 2207 11700 2241
rect 11700 2207 11704 2241
rect 11526 2173 11704 2207
rect 11526 2139 11530 2173
rect 11530 2139 11598 2173
rect 11598 2139 11632 2173
rect 11632 2139 11700 2173
rect 11700 2139 11704 2173
rect 11526 2105 11704 2139
rect 11526 2071 11530 2105
rect 11530 2071 11598 2105
rect 11598 2071 11632 2105
rect 11632 2071 11700 2105
rect 11700 2071 11704 2105
rect 11526 2037 11704 2071
rect 11526 2003 11530 2037
rect 11530 2003 11598 2037
rect 11598 2003 11632 2037
rect 11632 2003 11700 2037
rect 11700 2003 11704 2037
rect 11526 1969 11704 2003
rect 11526 1935 11530 1969
rect 11530 1935 11598 1969
rect 11598 1935 11632 1969
rect 11632 1935 11700 1969
rect 11700 1935 11704 1969
rect 11526 1901 11704 1935
rect 11526 1867 11530 1901
rect 11530 1867 11598 1901
rect 11598 1867 11632 1901
rect 11632 1867 11700 1901
rect 11700 1867 11704 1901
rect 11526 1833 11704 1867
rect 11526 1799 11530 1833
rect 11530 1799 11598 1833
rect 11598 1799 11632 1833
rect 11632 1799 11700 1833
rect 11700 1799 11704 1833
rect 11526 1765 11704 1799
rect 11526 1731 11530 1765
rect 11530 1731 11598 1765
rect 11598 1731 11632 1765
rect 11632 1731 11700 1765
rect 11700 1731 11704 1765
rect 11526 1697 11704 1731
rect 11526 1663 11530 1697
rect 11530 1663 11598 1697
rect 11598 1663 11632 1697
rect 11632 1663 11700 1697
rect 11700 1663 11704 1697
rect 11526 1629 11704 1663
rect 11526 1595 11530 1629
rect 11530 1595 11598 1629
rect 11598 1595 11632 1629
rect 11632 1595 11700 1629
rect 11700 1595 11704 1629
rect 11526 1561 11704 1595
rect 11526 1527 11530 1561
rect 11530 1527 11598 1561
rect 11598 1527 11632 1561
rect 11632 1527 11700 1561
rect 11700 1527 11704 1561
rect 11526 1491 11704 1527
rect 11526 1479 11560 1491
rect 11670 1479 11704 1491
rect 12273 4388 12379 4494
rect 12022 4028 12056 4062
rect 12094 4028 12128 4062
rect 12166 4028 12200 4062
rect 12022 3954 12056 3988
rect 12094 3954 12128 3988
rect 12166 3954 12200 3988
rect 12022 3880 12056 3914
rect 12094 3880 12128 3914
rect 12166 3880 12200 3914
rect 12022 3806 12056 3840
rect 12094 3806 12128 3840
rect 12166 3806 12200 3840
rect 12022 3732 12056 3766
rect 12094 3732 12128 3766
rect 12166 3732 12200 3766
rect 12022 3658 12056 3692
rect 12094 3658 12128 3692
rect 12166 3658 12200 3692
rect 12022 3584 12056 3618
rect 12094 3584 12128 3618
rect 12166 3584 12200 3618
rect 12022 3510 12056 3544
rect 12094 3510 12128 3544
rect 12166 3510 12200 3544
rect 12022 3436 12056 3470
rect 12094 3436 12128 3470
rect 12166 3436 12200 3470
rect 12022 3362 12056 3396
rect 12094 3362 12128 3396
rect 12166 3362 12200 3396
rect 12022 3288 12056 3322
rect 12094 3288 12128 3322
rect 12166 3288 12200 3322
rect 12022 3214 12056 3248
rect 12094 3214 12128 3248
rect 12166 3214 12200 3248
rect 12022 3140 12056 3174
rect 12094 3140 12128 3174
rect 12166 3140 12200 3174
rect 12022 3066 12056 3100
rect 12094 3066 12128 3100
rect 12166 3066 12200 3100
rect 12022 2992 12056 3026
rect 12094 2992 12128 3026
rect 12166 2992 12200 3026
rect 12022 2918 12056 2952
rect 12094 2918 12128 2952
rect 12166 2918 12200 2952
rect 12022 2844 12056 2878
rect 12094 2844 12128 2878
rect 12166 2844 12200 2878
rect 12022 2770 12056 2804
rect 12094 2770 12128 2804
rect 12166 2770 12200 2804
rect 12022 2696 12056 2730
rect 12094 2696 12128 2730
rect 12166 2696 12200 2730
rect 12022 2622 12056 2656
rect 12094 2622 12128 2656
rect 12166 2622 12200 2656
rect 12022 2548 12056 2582
rect 12094 2548 12128 2582
rect 12166 2548 12200 2582
rect 12022 2474 12056 2508
rect 12094 2474 12128 2508
rect 12166 2474 12200 2508
rect 12022 2400 12056 2434
rect 12094 2400 12128 2434
rect 12166 2400 12200 2434
rect 12022 2326 12056 2360
rect 12094 2326 12128 2360
rect 12166 2326 12200 2360
rect 12022 2252 12056 2286
rect 12094 2252 12128 2286
rect 12166 2252 12200 2286
rect 12022 2178 12056 2212
rect 12094 2178 12128 2212
rect 12166 2178 12200 2212
rect 12022 2104 12056 2138
rect 12094 2104 12128 2138
rect 12166 2104 12200 2138
rect 12022 2030 12056 2064
rect 12094 2030 12128 2064
rect 12166 2030 12200 2064
rect 12022 1956 12056 1990
rect 12094 1956 12128 1990
rect 12166 1956 12200 1990
rect 12022 1882 12056 1916
rect 12094 1882 12128 1916
rect 12166 1882 12200 1916
rect 12022 1808 12056 1842
rect 12094 1808 12128 1842
rect 12166 1808 12200 1842
rect 12022 1734 12056 1768
rect 12094 1734 12128 1768
rect 12166 1734 12200 1768
rect 12022 1660 12056 1694
rect 12094 1660 12128 1694
rect 12166 1660 12200 1694
rect 12022 1586 12056 1620
rect 12094 1586 12128 1620
rect 12166 1586 12200 1620
rect 12022 1511 12056 1545
rect 12094 1511 12128 1545
rect 12166 1511 12200 1545
rect 12835 4388 12941 4494
rect 12590 4050 12624 4062
rect 12518 4046 12696 4050
rect 12518 4012 12522 4046
rect 12522 4012 12590 4046
rect 12590 4012 12624 4046
rect 12624 4012 12692 4046
rect 12692 4012 12696 4046
rect 12518 3978 12696 4012
rect 12518 3944 12522 3978
rect 12522 3944 12590 3978
rect 12590 3944 12624 3978
rect 12624 3944 12692 3978
rect 12692 3944 12696 3978
rect 12518 3910 12696 3944
rect 12518 3876 12522 3910
rect 12522 3876 12590 3910
rect 12590 3876 12624 3910
rect 12624 3876 12692 3910
rect 12692 3876 12696 3910
rect 12518 3842 12696 3876
rect 12518 3808 12522 3842
rect 12522 3808 12590 3842
rect 12590 3808 12624 3842
rect 12624 3808 12692 3842
rect 12692 3808 12696 3842
rect 12518 3774 12696 3808
rect 12518 3740 12522 3774
rect 12522 3740 12590 3774
rect 12590 3740 12624 3774
rect 12624 3740 12692 3774
rect 12692 3740 12696 3774
rect 12518 3706 12696 3740
rect 12518 3672 12522 3706
rect 12522 3672 12590 3706
rect 12590 3672 12624 3706
rect 12624 3672 12692 3706
rect 12692 3672 12696 3706
rect 12518 3638 12696 3672
rect 12518 3604 12522 3638
rect 12522 3604 12590 3638
rect 12590 3604 12624 3638
rect 12624 3604 12692 3638
rect 12692 3604 12696 3638
rect 12518 3570 12696 3604
rect 12518 3536 12522 3570
rect 12522 3536 12590 3570
rect 12590 3536 12624 3570
rect 12624 3536 12692 3570
rect 12692 3536 12696 3570
rect 12518 3502 12696 3536
rect 12518 3468 12522 3502
rect 12522 3468 12590 3502
rect 12590 3468 12624 3502
rect 12624 3468 12692 3502
rect 12692 3468 12696 3502
rect 12518 3434 12696 3468
rect 12518 3400 12522 3434
rect 12522 3400 12590 3434
rect 12590 3400 12624 3434
rect 12624 3400 12692 3434
rect 12692 3400 12696 3434
rect 12518 3366 12696 3400
rect 12518 3332 12522 3366
rect 12522 3332 12590 3366
rect 12590 3332 12624 3366
rect 12624 3332 12692 3366
rect 12692 3332 12696 3366
rect 12518 3298 12696 3332
rect 12518 3264 12522 3298
rect 12522 3264 12590 3298
rect 12590 3264 12624 3298
rect 12624 3264 12692 3298
rect 12692 3264 12696 3298
rect 12518 3230 12696 3264
rect 12518 3196 12522 3230
rect 12522 3196 12590 3230
rect 12590 3196 12624 3230
rect 12624 3196 12692 3230
rect 12692 3196 12696 3230
rect 12518 3162 12696 3196
rect 12518 3128 12522 3162
rect 12522 3128 12590 3162
rect 12590 3128 12624 3162
rect 12624 3128 12692 3162
rect 12692 3128 12696 3162
rect 12518 3092 12696 3128
rect 12518 3080 12552 3092
rect 12662 3080 12696 3092
rect 12518 3004 12552 3038
rect 12590 3004 12624 3038
rect 12662 3004 12696 3038
rect 12518 2921 12552 2955
rect 12590 2935 12624 2955
rect 12590 2921 12591 2935
rect 12591 2921 12624 2935
rect 12662 2921 12696 2955
rect 12518 2837 12552 2871
rect 12590 2855 12624 2871
rect 12590 2837 12591 2855
rect 12591 2837 12624 2855
rect 12662 2837 12696 2871
rect 12518 2753 12552 2787
rect 12590 2775 12624 2787
rect 12590 2753 12591 2775
rect 12591 2753 12624 2775
rect 12662 2753 12696 2787
rect 12518 2669 12552 2703
rect 12590 2695 12624 2703
rect 12590 2669 12591 2695
rect 12591 2669 12624 2695
rect 12662 2669 12696 2703
rect 12518 2585 12552 2619
rect 12590 2614 12624 2619
rect 12590 2585 12591 2614
rect 12591 2585 12624 2614
rect 12662 2585 12696 2619
rect 12518 2501 12552 2535
rect 12590 2501 12624 2535
rect 12662 2501 12696 2535
rect 12590 2449 12624 2461
rect 12518 2445 12696 2449
rect 12518 2411 12522 2445
rect 12522 2411 12590 2445
rect 12590 2411 12624 2445
rect 12624 2411 12692 2445
rect 12692 2411 12696 2445
rect 12518 2377 12696 2411
rect 12518 2343 12522 2377
rect 12522 2343 12590 2377
rect 12590 2343 12624 2377
rect 12624 2343 12692 2377
rect 12692 2343 12696 2377
rect 12518 2309 12696 2343
rect 12518 2275 12522 2309
rect 12522 2275 12590 2309
rect 12590 2275 12624 2309
rect 12624 2275 12692 2309
rect 12692 2275 12696 2309
rect 12518 2241 12696 2275
rect 12518 2207 12522 2241
rect 12522 2207 12590 2241
rect 12590 2207 12624 2241
rect 12624 2207 12692 2241
rect 12692 2207 12696 2241
rect 12518 2173 12696 2207
rect 12518 2139 12522 2173
rect 12522 2139 12590 2173
rect 12590 2139 12624 2173
rect 12624 2139 12692 2173
rect 12692 2139 12696 2173
rect 12518 2105 12696 2139
rect 12518 2071 12522 2105
rect 12522 2071 12590 2105
rect 12590 2071 12624 2105
rect 12624 2071 12692 2105
rect 12692 2071 12696 2105
rect 12518 2037 12696 2071
rect 12518 2003 12522 2037
rect 12522 2003 12590 2037
rect 12590 2003 12624 2037
rect 12624 2003 12692 2037
rect 12692 2003 12696 2037
rect 12518 1969 12696 2003
rect 12518 1935 12522 1969
rect 12522 1935 12590 1969
rect 12590 1935 12624 1969
rect 12624 1935 12692 1969
rect 12692 1935 12696 1969
rect 12518 1901 12696 1935
rect 12518 1867 12522 1901
rect 12522 1867 12590 1901
rect 12590 1867 12624 1901
rect 12624 1867 12692 1901
rect 12692 1867 12696 1901
rect 12518 1833 12696 1867
rect 12518 1799 12522 1833
rect 12522 1799 12590 1833
rect 12590 1799 12624 1833
rect 12624 1799 12692 1833
rect 12692 1799 12696 1833
rect 12518 1765 12696 1799
rect 12518 1731 12522 1765
rect 12522 1731 12590 1765
rect 12590 1731 12624 1765
rect 12624 1731 12692 1765
rect 12692 1731 12696 1765
rect 12518 1697 12696 1731
rect 12518 1663 12522 1697
rect 12522 1663 12590 1697
rect 12590 1663 12624 1697
rect 12624 1663 12692 1697
rect 12692 1663 12696 1697
rect 12518 1629 12696 1663
rect 12518 1595 12522 1629
rect 12522 1595 12590 1629
rect 12590 1595 12624 1629
rect 12624 1595 12692 1629
rect 12692 1595 12696 1629
rect 12518 1561 12696 1595
rect 12518 1527 12522 1561
rect 12522 1527 12590 1561
rect 12590 1527 12624 1561
rect 12624 1527 12692 1561
rect 12692 1527 12696 1561
rect 12518 1491 12696 1527
rect 12518 1479 12552 1491
rect 12662 1479 12696 1491
rect 13265 4388 13371 4494
rect 13014 4028 13048 4062
rect 13086 4028 13120 4062
rect 13158 4028 13192 4062
rect 13014 3954 13048 3988
rect 13086 3954 13120 3988
rect 13158 3954 13192 3988
rect 13014 3880 13048 3914
rect 13086 3880 13120 3914
rect 13158 3880 13192 3914
rect 13014 3806 13048 3840
rect 13086 3806 13120 3840
rect 13158 3806 13192 3840
rect 13014 3732 13048 3766
rect 13086 3732 13120 3766
rect 13158 3732 13192 3766
rect 13014 3658 13048 3692
rect 13086 3658 13120 3692
rect 13158 3658 13192 3692
rect 13014 3584 13048 3618
rect 13086 3584 13120 3618
rect 13158 3584 13192 3618
rect 13014 3510 13048 3544
rect 13086 3510 13120 3544
rect 13158 3510 13192 3544
rect 13014 3436 13048 3470
rect 13086 3436 13120 3470
rect 13158 3436 13192 3470
rect 13014 3362 13048 3396
rect 13086 3362 13120 3396
rect 13158 3362 13192 3396
rect 13014 3288 13048 3322
rect 13086 3288 13120 3322
rect 13158 3288 13192 3322
rect 13014 3214 13048 3248
rect 13086 3214 13120 3248
rect 13158 3214 13192 3248
rect 13014 3140 13048 3174
rect 13086 3140 13120 3174
rect 13158 3140 13192 3174
rect 13014 3066 13048 3100
rect 13086 3066 13120 3100
rect 13158 3066 13192 3100
rect 13014 2992 13048 3026
rect 13086 2992 13120 3026
rect 13158 2992 13192 3026
rect 13014 2918 13048 2952
rect 13086 2918 13120 2952
rect 13158 2918 13192 2952
rect 13014 2844 13048 2878
rect 13086 2844 13120 2878
rect 13158 2844 13192 2878
rect 13014 2770 13048 2804
rect 13086 2770 13120 2804
rect 13158 2770 13192 2804
rect 13014 2696 13048 2730
rect 13086 2696 13120 2730
rect 13158 2696 13192 2730
rect 13014 2622 13048 2656
rect 13086 2622 13120 2656
rect 13158 2622 13192 2656
rect 13014 2548 13048 2582
rect 13086 2548 13120 2582
rect 13158 2548 13192 2582
rect 13014 2474 13048 2508
rect 13086 2474 13120 2508
rect 13158 2474 13192 2508
rect 13014 2400 13048 2434
rect 13086 2400 13120 2434
rect 13158 2400 13192 2434
rect 13014 2326 13048 2360
rect 13086 2326 13120 2360
rect 13158 2326 13192 2360
rect 13014 2252 13048 2286
rect 13086 2252 13120 2286
rect 13158 2252 13192 2286
rect 13014 2178 13048 2212
rect 13086 2178 13120 2212
rect 13158 2178 13192 2212
rect 13014 2104 13048 2138
rect 13086 2104 13120 2138
rect 13158 2104 13192 2138
rect 13014 2030 13048 2064
rect 13086 2030 13120 2064
rect 13158 2030 13192 2064
rect 13014 1956 13048 1990
rect 13086 1956 13120 1990
rect 13158 1956 13192 1990
rect 13014 1882 13048 1916
rect 13086 1882 13120 1916
rect 13158 1882 13192 1916
rect 13014 1808 13048 1842
rect 13086 1808 13120 1842
rect 13158 1808 13192 1842
rect 13014 1734 13048 1768
rect 13086 1734 13120 1768
rect 13158 1734 13192 1768
rect 13014 1660 13048 1694
rect 13086 1660 13120 1694
rect 13158 1660 13192 1694
rect 13014 1586 13048 1620
rect 13086 1586 13120 1620
rect 13158 1586 13192 1620
rect 13014 1511 13048 1545
rect 13086 1511 13120 1545
rect 13158 1511 13192 1545
rect 13827 4388 13933 4494
rect 13582 4050 13616 4062
rect 13510 4046 13688 4050
rect 13510 4012 13514 4046
rect 13514 4012 13582 4046
rect 13582 4012 13616 4046
rect 13616 4012 13684 4046
rect 13684 4012 13688 4046
rect 13510 3978 13688 4012
rect 13510 3944 13514 3978
rect 13514 3944 13582 3978
rect 13582 3944 13616 3978
rect 13616 3944 13684 3978
rect 13684 3944 13688 3978
rect 13510 3910 13688 3944
rect 13510 3876 13514 3910
rect 13514 3876 13582 3910
rect 13582 3876 13616 3910
rect 13616 3876 13684 3910
rect 13684 3876 13688 3910
rect 13510 3842 13688 3876
rect 13510 3808 13514 3842
rect 13514 3808 13582 3842
rect 13582 3808 13616 3842
rect 13616 3808 13684 3842
rect 13684 3808 13688 3842
rect 13510 3774 13688 3808
rect 13510 3740 13514 3774
rect 13514 3740 13582 3774
rect 13582 3740 13616 3774
rect 13616 3740 13684 3774
rect 13684 3740 13688 3774
rect 13510 3706 13688 3740
rect 13510 3672 13514 3706
rect 13514 3672 13582 3706
rect 13582 3672 13616 3706
rect 13616 3672 13684 3706
rect 13684 3672 13688 3706
rect 13510 3638 13688 3672
rect 13510 3604 13514 3638
rect 13514 3604 13582 3638
rect 13582 3604 13616 3638
rect 13616 3604 13684 3638
rect 13684 3604 13688 3638
rect 13510 3570 13688 3604
rect 13510 3536 13514 3570
rect 13514 3536 13582 3570
rect 13582 3536 13616 3570
rect 13616 3536 13684 3570
rect 13684 3536 13688 3570
rect 13510 3502 13688 3536
rect 13510 3468 13514 3502
rect 13514 3468 13582 3502
rect 13582 3468 13616 3502
rect 13616 3468 13684 3502
rect 13684 3468 13688 3502
rect 13510 3434 13688 3468
rect 13510 3400 13514 3434
rect 13514 3400 13582 3434
rect 13582 3400 13616 3434
rect 13616 3400 13684 3434
rect 13684 3400 13688 3434
rect 13510 3366 13688 3400
rect 13510 3332 13514 3366
rect 13514 3332 13582 3366
rect 13582 3332 13616 3366
rect 13616 3332 13684 3366
rect 13684 3332 13688 3366
rect 13510 3298 13688 3332
rect 13510 3264 13514 3298
rect 13514 3264 13582 3298
rect 13582 3264 13616 3298
rect 13616 3264 13684 3298
rect 13684 3264 13688 3298
rect 13510 3230 13688 3264
rect 13510 3196 13514 3230
rect 13514 3196 13582 3230
rect 13582 3196 13616 3230
rect 13616 3196 13684 3230
rect 13684 3196 13688 3230
rect 13510 3162 13688 3196
rect 13510 3128 13514 3162
rect 13514 3128 13582 3162
rect 13582 3128 13616 3162
rect 13616 3128 13684 3162
rect 13684 3128 13688 3162
rect 13510 3092 13688 3128
rect 13510 3080 13544 3092
rect 13654 3080 13688 3092
rect 13510 2935 13688 3040
rect 13510 2901 13549 2935
rect 13549 2901 13583 2935
rect 13583 2901 13617 2935
rect 13617 2901 13651 2935
rect 13651 2901 13688 2935
rect 13510 2855 13688 2901
rect 13510 2821 13549 2855
rect 13549 2821 13583 2855
rect 13583 2821 13617 2855
rect 13617 2821 13651 2855
rect 13651 2821 13688 2855
rect 13510 2775 13688 2821
rect 13510 2741 13549 2775
rect 13549 2741 13583 2775
rect 13583 2741 13617 2775
rect 13617 2741 13651 2775
rect 13651 2741 13688 2775
rect 13510 2695 13688 2741
rect 13510 2661 13549 2695
rect 13549 2661 13583 2695
rect 13583 2661 13617 2695
rect 13617 2661 13651 2695
rect 13651 2661 13688 2695
rect 13510 2614 13688 2661
rect 13510 2580 13549 2614
rect 13549 2580 13583 2614
rect 13583 2580 13617 2614
rect 13617 2580 13651 2614
rect 13651 2580 13688 2614
rect 13510 2574 13688 2580
rect 13510 2501 13544 2535
rect 13582 2501 13616 2535
rect 13654 2501 13688 2535
rect 13582 2449 13616 2461
rect 13510 2445 13688 2449
rect 13510 2411 13514 2445
rect 13514 2411 13582 2445
rect 13582 2411 13616 2445
rect 13616 2411 13684 2445
rect 13684 2411 13688 2445
rect 13510 2377 13688 2411
rect 13510 2343 13514 2377
rect 13514 2343 13582 2377
rect 13582 2343 13616 2377
rect 13616 2343 13684 2377
rect 13684 2343 13688 2377
rect 13510 2309 13688 2343
rect 13510 2275 13514 2309
rect 13514 2275 13582 2309
rect 13582 2275 13616 2309
rect 13616 2275 13684 2309
rect 13684 2275 13688 2309
rect 13510 2241 13688 2275
rect 13510 2207 13514 2241
rect 13514 2207 13582 2241
rect 13582 2207 13616 2241
rect 13616 2207 13684 2241
rect 13684 2207 13688 2241
rect 13510 2173 13688 2207
rect 13510 2139 13514 2173
rect 13514 2139 13582 2173
rect 13582 2139 13616 2173
rect 13616 2139 13684 2173
rect 13684 2139 13688 2173
rect 13510 2105 13688 2139
rect 13510 2071 13514 2105
rect 13514 2071 13582 2105
rect 13582 2071 13616 2105
rect 13616 2071 13684 2105
rect 13684 2071 13688 2105
rect 13510 2037 13688 2071
rect 13510 2003 13514 2037
rect 13514 2003 13582 2037
rect 13582 2003 13616 2037
rect 13616 2003 13684 2037
rect 13684 2003 13688 2037
rect 13510 1969 13688 2003
rect 13510 1935 13514 1969
rect 13514 1935 13582 1969
rect 13582 1935 13616 1969
rect 13616 1935 13684 1969
rect 13684 1935 13688 1969
rect 13510 1901 13688 1935
rect 13510 1867 13514 1901
rect 13514 1867 13582 1901
rect 13582 1867 13616 1901
rect 13616 1867 13684 1901
rect 13684 1867 13688 1901
rect 13510 1833 13688 1867
rect 13510 1799 13514 1833
rect 13514 1799 13582 1833
rect 13582 1799 13616 1833
rect 13616 1799 13684 1833
rect 13684 1799 13688 1833
rect 13510 1765 13688 1799
rect 13510 1731 13514 1765
rect 13514 1731 13582 1765
rect 13582 1731 13616 1765
rect 13616 1731 13684 1765
rect 13684 1731 13688 1765
rect 13510 1697 13688 1731
rect 13510 1663 13514 1697
rect 13514 1663 13582 1697
rect 13582 1663 13616 1697
rect 13616 1663 13684 1697
rect 13684 1663 13688 1697
rect 13510 1629 13688 1663
rect 13510 1595 13514 1629
rect 13514 1595 13582 1629
rect 13582 1595 13616 1629
rect 13616 1595 13684 1629
rect 13684 1595 13688 1629
rect 13510 1561 13688 1595
rect 13510 1527 13514 1561
rect 13514 1527 13582 1561
rect 13582 1527 13616 1561
rect 13616 1527 13684 1561
rect 13684 1527 13688 1561
rect 13510 1491 13688 1527
rect 13510 1479 13544 1491
rect 13654 1479 13688 1491
rect 14185 4388 14291 4494
rect 14042 4046 14076 4062
rect 14042 4028 14076 4046
rect 14042 3978 14076 3990
rect 14042 3956 14076 3978
rect 14042 3910 14076 3918
rect 14042 3884 14076 3910
rect 14042 3842 14076 3846
rect 14042 3812 14076 3842
rect 14042 3740 14076 3774
rect 14042 3672 14076 3702
rect 14042 3668 14076 3672
rect 14042 3604 14076 3630
rect 14042 3596 14076 3604
rect 14042 3536 14076 3558
rect 14042 3524 14076 3536
rect 14042 3468 14076 3486
rect 14042 3452 14076 3468
rect 14042 3400 14076 3414
rect 14042 3380 14076 3400
rect 14042 3332 14076 3342
rect 14042 3308 14076 3332
rect 14042 3264 14076 3270
rect 14042 3236 14076 3264
rect 14042 3196 14076 3198
rect 14042 3164 14076 3196
rect 14042 3092 14076 3126
rect 14042 3020 14076 3054
rect 14042 2948 14076 2982
rect 14042 2876 14076 2910
rect 14042 2804 14076 2838
rect 14042 2732 14076 2766
rect 14042 2659 14076 2693
rect 14042 2586 14076 2620
rect 14042 2513 14076 2547
rect 14042 2445 14076 2474
rect 14042 2440 14076 2445
rect 14042 2377 14076 2401
rect 14042 2367 14076 2377
rect 14042 2309 14076 2328
rect 14042 2294 14076 2309
rect 14042 2241 14076 2255
rect 14042 2221 14076 2241
rect 14042 2173 14076 2182
rect 14042 2148 14076 2173
rect 14042 2105 14076 2109
rect 14042 2075 14076 2105
rect 14042 2003 14076 2036
rect 14042 2002 14076 2003
rect 14042 1935 14076 1963
rect 14042 1929 14076 1935
rect 14042 1867 14076 1890
rect 14042 1856 14076 1867
rect 14042 1799 14076 1817
rect 14042 1783 14076 1799
rect 14042 1731 14076 1744
rect 14042 1710 14076 1731
rect 14042 1663 14076 1671
rect 14042 1637 14076 1663
rect 14042 1595 14076 1598
rect 14042 1564 14076 1595
rect 14042 1491 14076 1525
rect 14510 4490 14544 4506
rect 14582 4504 14599 4524
rect 14599 4504 14616 4524
rect 14582 4490 14616 4504
rect 14431 4448 14465 4482
rect 14510 4436 14531 4451
rect 14531 4436 14544 4451
rect 14510 4417 14544 4436
rect 14582 4434 14599 4451
rect 14599 4434 14616 4451
rect 14582 4417 14616 4434
rect 14431 4375 14465 4409
rect 14510 4365 14531 4378
rect 14531 4365 14544 4378
rect 14510 4344 14544 4365
rect 14582 4364 14599 4378
rect 14599 4364 14616 4378
rect 14582 4344 14616 4364
rect 14431 4302 14465 4336
rect 14510 4294 14531 4305
rect 14531 4294 14544 4305
rect 14582 4294 14599 4305
rect 14599 4294 14616 4305
rect 14510 4271 14544 4294
rect 14582 4271 14616 4294
rect 14431 4229 14465 4263
rect 14510 4223 14531 4232
rect 14531 4223 14544 4232
rect 14582 4223 14599 4232
rect 14599 4223 14616 4232
rect 14510 4198 14544 4223
rect 14582 4198 14616 4223
rect 14431 4156 14465 4190
rect 14510 4152 14531 4159
rect 14531 4152 14544 4159
rect 14582 4152 14599 4159
rect 14599 4152 14616 4159
rect 14510 4125 14544 4152
rect 14582 4125 14616 4152
rect 14431 4083 14465 4117
rect 14510 4052 14544 4086
rect 14582 4081 14599 4086
rect 14599 4081 14616 4086
rect 14582 4052 14616 4081
rect 14431 4034 14465 4044
rect 14431 4010 14454 4034
rect 14454 4010 14465 4034
rect 14510 3979 14544 4013
rect 14582 4007 14599 4013
rect 14599 4007 14616 4013
rect 14582 3979 14616 4007
rect 14431 3966 14465 3971
rect 14431 3937 14454 3966
rect 14454 3937 14465 3966
rect 14510 3906 14544 3940
rect 14582 3936 14599 3940
rect 14599 3936 14616 3940
rect 14582 3906 14616 3936
rect 14431 3864 14454 3898
rect 14454 3864 14465 3898
rect 14510 3833 14544 3867
rect 14582 3862 14599 3867
rect 14599 3862 14616 3867
rect 14582 3833 14616 3862
rect 14431 3796 14454 3825
rect 14454 3796 14465 3825
rect 14431 3791 14465 3796
rect 14510 3760 14544 3794
rect 14582 3791 14599 3794
rect 14599 3791 14616 3794
rect 14582 3760 14616 3791
rect 14431 3728 14454 3752
rect 14454 3728 14465 3752
rect 14431 3718 14465 3728
rect 14510 3687 14544 3721
rect 14582 3717 14599 3721
rect 14599 3717 14616 3721
rect 14582 3687 14616 3717
rect 14431 3660 14454 3679
rect 14454 3660 14465 3679
rect 14431 3645 14465 3660
rect 14510 3614 14544 3648
rect 14582 3646 14599 3648
rect 14599 3646 14616 3648
rect 14582 3614 14616 3646
rect 14431 3592 14454 3606
rect 14454 3592 14465 3606
rect 14431 3572 14465 3592
rect 14510 3541 14544 3575
rect 14582 3572 14599 3575
rect 14599 3572 14616 3575
rect 14582 3541 14616 3572
rect 14431 3524 14454 3533
rect 14454 3524 14465 3533
rect 14431 3499 14465 3524
rect 14510 3468 14544 3502
rect 14582 3501 14599 3502
rect 14599 3501 14616 3502
rect 14582 3468 14616 3501
rect 14431 3456 14454 3460
rect 14454 3456 14465 3460
rect 14431 3426 14465 3456
rect 14510 3395 14544 3429
rect 14582 3427 14599 3429
rect 14599 3427 14616 3429
rect 14582 3395 14616 3427
rect 14431 3354 14465 3387
rect 14431 3353 14454 3354
rect 14454 3353 14465 3354
rect 14510 3322 14544 3356
rect 14582 3322 14616 3356
rect 14431 3286 14465 3314
rect 14431 3280 14454 3286
rect 14454 3280 14465 3286
rect 14510 3249 14544 3283
rect 14582 3282 14599 3283
rect 14599 3282 14616 3283
rect 14582 3249 14616 3282
rect 14431 3218 14465 3241
rect 14431 3207 14454 3218
rect 14454 3207 14465 3218
rect 14510 3176 14544 3210
rect 14582 3176 14616 3210
rect 14431 3150 14465 3168
rect 14431 3134 14454 3150
rect 14454 3134 14465 3150
rect 14510 3103 14544 3137
rect 14582 3117 14599 3137
rect 14599 3117 14616 3137
rect 14582 3103 14616 3117
rect 14431 3061 14465 3095
rect 14510 3030 14544 3064
rect 14582 3032 14599 3064
rect 14599 3032 14616 3064
rect 14582 3030 14616 3032
rect 14431 2988 14465 3022
rect 14510 2972 14544 2991
rect 14582 2972 14616 2991
rect 14510 2957 14544 2972
rect 14582 2957 14616 2972
rect 14431 2915 14465 2949
rect 14510 2884 14544 2918
rect 14582 2884 14616 2918
rect 14431 2842 14465 2876
rect 14510 2811 14544 2845
rect 14582 2811 14616 2845
rect 14431 2769 14465 2803
rect 14510 2738 14544 2772
rect 14582 2738 14616 2772
rect 14431 2696 14465 2730
rect 14510 2665 14544 2699
rect 14582 2665 14616 2699
rect 14431 2623 14465 2657
rect 14510 2592 14544 2626
rect 14582 2592 14616 2626
rect 14431 2550 14465 2584
rect 14510 2530 14544 2553
rect 14582 2530 14616 2553
rect 14510 2519 14544 2530
rect 14582 2519 14616 2530
rect 14431 2477 14465 2511
rect 14510 2446 14544 2480
rect 14582 2451 14599 2480
rect 14599 2451 14616 2480
rect 14582 2446 14616 2451
rect 14431 2433 14465 2438
rect 14431 2404 14454 2433
rect 14454 2404 14465 2433
rect 14510 2373 14544 2407
rect 14582 2403 14616 2407
rect 14582 2373 14599 2403
rect 14599 2373 14616 2403
rect 14431 2331 14454 2365
rect 14454 2331 14465 2365
rect 14510 2300 14544 2334
rect 14582 2327 14616 2334
rect 14582 2300 14599 2327
rect 14599 2300 14616 2327
rect 14431 2263 14454 2292
rect 14454 2263 14465 2292
rect 14431 2258 14465 2263
rect 14510 2226 14544 2260
rect 14582 2250 14616 2260
rect 14582 2226 14599 2250
rect 14599 2226 14616 2250
rect 14431 2195 14454 2219
rect 14454 2195 14465 2219
rect 14431 2185 14465 2195
rect 14510 2152 14544 2186
rect 14582 2156 14616 2186
rect 14582 2152 14599 2156
rect 14599 2152 14616 2156
rect 14431 2127 14454 2146
rect 14454 2127 14465 2146
rect 14431 2112 14465 2127
rect 14510 2078 14544 2112
rect 14582 2085 14616 2112
rect 14582 2078 14599 2085
rect 14599 2078 14616 2085
rect 14431 2059 14454 2073
rect 14454 2059 14465 2073
rect 14431 2039 14465 2059
rect 14510 2004 14544 2038
rect 14582 2011 14616 2038
rect 14582 2004 14599 2011
rect 14599 2004 14616 2011
rect 14431 1991 14454 2000
rect 14454 1991 14465 2000
rect 14431 1966 14465 1991
rect 14510 1930 14544 1964
rect 14582 1940 14616 1964
rect 14582 1930 14599 1940
rect 14599 1930 14616 1940
rect 14431 1923 14454 1927
rect 14454 1923 14465 1927
rect 14431 1893 14465 1923
rect 14510 1856 14544 1890
rect 14582 1866 14616 1890
rect 14582 1856 14599 1866
rect 14599 1856 14616 1866
rect 14431 1821 14465 1854
rect 14431 1820 14454 1821
rect 14454 1820 14465 1821
rect 14510 1782 14544 1816
rect 14582 1795 14616 1816
rect 14582 1782 14599 1795
rect 14599 1782 14616 1795
rect 14431 1753 14465 1781
rect 14431 1747 14454 1753
rect 14454 1747 14465 1753
rect 14510 1708 14544 1742
rect 14582 1721 14616 1742
rect 14582 1708 14599 1721
rect 14599 1708 14616 1721
rect 14431 1685 14465 1708
rect 14431 1674 14454 1685
rect 14454 1674 14465 1685
rect 14431 1617 14465 1635
rect 14510 1634 14544 1668
rect 14582 1650 14616 1668
rect 14582 1634 14599 1650
rect 14599 1634 14616 1650
rect 14431 1601 14454 1617
rect 14454 1601 14465 1617
rect 14431 1549 14465 1562
rect 14510 1560 14544 1594
rect 14582 1576 14616 1594
rect 14582 1560 14599 1576
rect 14599 1560 14616 1576
rect 14431 1528 14454 1549
rect 14454 1528 14465 1549
rect 14431 1455 14465 1489
rect 14510 1486 14544 1520
rect 14582 1505 14616 1520
rect 14582 1486 14599 1505
rect 14599 1486 14616 1505
rect 14431 1382 14465 1416
rect 14510 1412 14544 1446
rect 14582 1412 14616 1446
rect 14510 1353 14531 1372
rect 14531 1353 14544 1372
rect 14582 1353 14599 1372
rect 14599 1353 14616 1372
rect 14431 1308 14465 1342
rect 14510 1338 14544 1353
rect 14582 1338 14616 1353
rect 587 1221 621 1241
rect 587 1207 589 1221
rect 589 1207 621 1221
rect 659 1219 693 1241
rect 733 1234 767 1268
rect 659 1207 691 1219
rect 691 1207 693 1219
rect 733 1160 767 1194
rect 14510 1274 14531 1298
rect 14531 1274 14544 1298
rect 14582 1277 14599 1298
rect 14599 1277 14616 1298
rect 14431 1234 14465 1268
rect 14510 1264 14544 1274
rect 14582 1264 14616 1277
rect 14510 1194 14531 1224
rect 14531 1194 14544 1224
rect 14582 1200 14599 1224
rect 14599 1200 14616 1224
rect 14431 1160 14465 1194
rect 14510 1190 14544 1194
rect 14582 1190 14616 1200
rect 767 1114 794 1116
rect 794 1114 801 1116
rect 767 1082 801 1114
rect 840 1082 874 1116
rect 913 1082 947 1116
rect 986 1082 1020 1116
rect 1059 1082 1093 1116
rect 1132 1082 1166 1116
rect 1205 1082 1239 1116
rect 1278 1082 1312 1116
rect 1351 1082 1385 1116
rect 1424 1082 1458 1116
rect 1497 1082 1531 1116
rect 1570 1082 1604 1116
rect 1643 1082 1677 1116
rect 1716 1082 1750 1116
rect 1789 1082 1823 1116
rect 1862 1082 1896 1116
rect 1935 1082 1969 1116
rect 2008 1082 2042 1116
rect 2081 1082 2115 1116
rect 2154 1082 2188 1116
rect 2227 1082 2261 1116
rect 2300 1082 2334 1116
rect 2373 1082 2407 1116
rect 2446 1082 2480 1116
rect 2519 1082 2553 1116
rect 2592 1082 2626 1116
rect 2665 1082 2699 1116
rect 767 1010 801 1044
rect 840 1010 874 1044
rect 913 1010 947 1044
rect 986 1010 1020 1044
rect 1059 1010 1093 1044
rect 1132 1010 1166 1044
rect 1205 1010 1239 1044
rect 1278 1010 1312 1044
rect 1351 1010 1385 1044
rect 1424 1010 1458 1044
rect 1497 1010 1531 1044
rect 1570 1010 1604 1044
rect 1643 1010 1677 1044
rect 1716 1010 1750 1044
rect 1789 1010 1823 1044
rect 1862 1010 1896 1044
rect 1935 1010 1969 1044
rect 2008 1010 2042 1044
rect 2081 1010 2115 1044
rect 2154 1010 2188 1044
rect 2227 1010 2261 1044
rect 2300 1010 2334 1044
rect 2373 1010 2407 1044
rect 2446 1010 2480 1044
rect 2519 1010 2553 1044
rect 2592 1010 2626 1044
rect 2665 1010 2699 1044
rect 2738 1010 14436 1116
rect 14927 4934 14935 4968
rect 14935 4934 14969 4968
rect 14969 4934 15003 4968
rect 15003 4934 15037 4968
rect 15037 4934 15071 4968
rect 15071 4934 15105 4968
rect 14927 4896 15105 4934
rect 14927 4862 14935 4896
rect 14935 4862 14969 4896
rect 14969 4862 15003 4896
rect 15003 4862 15037 4896
rect 15037 4862 15071 4896
rect 15071 4862 15105 4896
rect 14927 4824 15105 4862
rect 14927 4790 14935 4824
rect 14935 4790 14969 4824
rect 14969 4790 15003 4824
rect 15003 4790 15037 4824
rect 15037 4790 15071 4824
rect 15071 4790 15105 4824
rect 14927 4752 15105 4790
rect 14927 4718 14935 4752
rect 14935 4718 14969 4752
rect 14969 4718 15003 4752
rect 15003 4718 15037 4752
rect 15037 4718 15071 4752
rect 15071 4718 15105 4752
rect 14927 4680 15105 4718
rect 14927 4646 14935 4680
rect 14935 4646 14969 4680
rect 14969 4646 15003 4680
rect 15003 4646 15037 4680
rect 15037 4646 15071 4680
rect 15071 4646 15105 4680
rect 14927 4608 15105 4646
rect 14927 4574 14935 4608
rect 14935 4574 14969 4608
rect 14969 4574 15003 4608
rect 15003 4574 15037 4608
rect 15037 4574 15071 4608
rect 15071 4574 15105 4608
rect 14927 4536 15105 4574
rect 14927 4502 14935 4536
rect 14935 4502 14969 4536
rect 14969 4502 15003 4536
rect 15003 4502 15037 4536
rect 15037 4502 15071 4536
rect 15071 4502 15105 4536
rect 14927 4464 15105 4502
rect 14927 4430 14935 4464
rect 14935 4430 14969 4464
rect 14969 4430 15003 4464
rect 15003 4430 15037 4464
rect 15037 4430 15071 4464
rect 15071 4430 15105 4464
rect 14927 4392 15105 4430
rect 14927 4358 14935 4392
rect 14935 4358 14969 4392
rect 14969 4358 15003 4392
rect 15003 4358 15037 4392
rect 15037 4358 15071 4392
rect 15071 4358 15105 4392
rect 14927 4320 15105 4358
rect 14927 4286 14935 4320
rect 14935 4286 14969 4320
rect 14969 4286 15003 4320
rect 15003 4286 15037 4320
rect 15037 4286 15071 4320
rect 15071 4286 15105 4320
rect 14927 4248 15105 4286
rect 14927 4214 14935 4248
rect 14935 4214 14969 4248
rect 14969 4214 15003 4248
rect 15003 4214 15037 4248
rect 15037 4214 15071 4248
rect 15071 4214 15105 4248
rect 14927 4176 15105 4214
rect 14927 4142 14935 4176
rect 14935 4142 14969 4176
rect 14969 4142 15003 4176
rect 15003 4142 15037 4176
rect 15037 4142 15071 4176
rect 15071 4142 15105 4176
rect 14927 4104 15105 4142
rect 14927 4070 14935 4104
rect 14935 4070 14969 4104
rect 14969 4070 15003 4104
rect 15003 4070 15037 4104
rect 15037 4070 15071 4104
rect 15071 4070 15105 4104
rect 14927 4032 15105 4070
rect 14927 3998 14935 4032
rect 14935 3998 14969 4032
rect 14969 3998 15003 4032
rect 15003 3998 15037 4032
rect 15037 3998 15071 4032
rect 15071 3998 15105 4032
rect 14927 3960 15105 3998
rect 14927 3926 14935 3960
rect 14935 3926 14969 3960
rect 14969 3926 15003 3960
rect 15003 3926 15037 3960
rect 15037 3926 15071 3960
rect 15071 3926 15105 3960
rect 14927 3888 15105 3926
rect 14927 3854 14935 3888
rect 14935 3854 14969 3888
rect 14969 3854 15003 3888
rect 15003 3854 15037 3888
rect 15037 3854 15071 3888
rect 15071 3854 15105 3888
rect 14927 3816 15105 3854
rect 14927 3782 14935 3816
rect 14935 3782 14969 3816
rect 14969 3782 15003 3816
rect 15003 3782 15037 3816
rect 15037 3782 15071 3816
rect 15071 3782 15105 3816
rect 14927 3744 15105 3782
rect 14927 3710 14935 3744
rect 14935 3710 14969 3744
rect 14969 3710 15003 3744
rect 15003 3710 15037 3744
rect 15037 3710 15071 3744
rect 15071 3710 15105 3744
rect 14927 3672 15105 3710
rect 14927 3638 14935 3672
rect 14935 3638 14969 3672
rect 14969 3638 15003 3672
rect 15003 3638 15037 3672
rect 15037 3638 15071 3672
rect 15071 3638 15105 3672
rect 14927 3600 15105 3638
rect 14927 3566 14935 3600
rect 14935 3566 14969 3600
rect 14969 3566 15003 3600
rect 15003 3566 15037 3600
rect 15037 3566 15071 3600
rect 15071 3566 15105 3600
rect 14927 3528 15105 3566
rect 14927 3494 14935 3528
rect 14935 3494 14969 3528
rect 14969 3494 15003 3528
rect 15003 3494 15037 3528
rect 15037 3494 15071 3528
rect 15071 3494 15105 3528
rect 14927 3456 15105 3494
rect 14927 3422 14935 3456
rect 14935 3422 14969 3456
rect 14969 3422 15003 3456
rect 15003 3422 15037 3456
rect 15037 3422 15071 3456
rect 15071 3422 15105 3456
rect 14927 3384 15105 3422
rect 14927 3350 14935 3384
rect 14935 3350 14969 3384
rect 14969 3350 15003 3384
rect 15003 3350 15037 3384
rect 15037 3350 15071 3384
rect 15071 3350 15105 3384
rect 14927 3312 15105 3350
rect 14927 3278 14935 3312
rect 14935 3278 14969 3312
rect 14969 3278 15003 3312
rect 15003 3278 15037 3312
rect 15037 3278 15071 3312
rect 15071 3278 15105 3312
rect 14927 3240 15105 3278
rect 14927 3206 14935 3240
rect 14935 3206 14969 3240
rect 14969 3206 15003 3240
rect 15003 3206 15037 3240
rect 15037 3206 15071 3240
rect 15071 3206 15105 3240
rect 14927 3168 15105 3206
rect 14927 3134 14935 3168
rect 14935 3134 14969 3168
rect 14969 3134 15003 3168
rect 15003 3134 15037 3168
rect 15037 3134 15071 3168
rect 15071 3134 15105 3168
rect 14927 3096 15105 3134
rect 14927 3062 14935 3096
rect 14935 3062 14969 3096
rect 14969 3062 15003 3096
rect 15003 3062 15037 3096
rect 15037 3062 15071 3096
rect 15071 3062 15105 3096
rect 14927 3024 15105 3062
rect 14927 2990 14935 3024
rect 14935 2990 14969 3024
rect 14969 2990 15003 3024
rect 15003 2990 15037 3024
rect 15037 2990 15071 3024
rect 15071 2990 15105 3024
rect 14927 2952 15105 2990
rect 14927 2918 14935 2952
rect 14935 2918 14969 2952
rect 14969 2918 15003 2952
rect 15003 2918 15037 2952
rect 15037 2918 15071 2952
rect 15071 2918 15105 2952
rect 14927 2880 15105 2918
rect 14927 2846 14935 2880
rect 14935 2846 14969 2880
rect 14969 2846 15003 2880
rect 15003 2846 15037 2880
rect 15037 2846 15071 2880
rect 15071 2846 15105 2880
rect 14927 2808 15105 2846
rect 14927 2774 14935 2808
rect 14935 2774 14969 2808
rect 14969 2774 15003 2808
rect 15003 2774 15037 2808
rect 15037 2774 15071 2808
rect 15071 2774 15105 2808
rect 14927 2736 15105 2774
rect 14927 2702 14935 2736
rect 14935 2702 14969 2736
rect 14969 2702 15003 2736
rect 15003 2702 15037 2736
rect 15037 2702 15071 2736
rect 15071 2702 15105 2736
rect 14927 2664 15105 2702
rect 14927 2630 14935 2664
rect 14935 2630 14969 2664
rect 14969 2630 15003 2664
rect 15003 2630 15037 2664
rect 15037 2630 15071 2664
rect 15071 2630 15105 2664
rect 14927 2592 15105 2630
rect 14927 2558 14935 2592
rect 14935 2558 14969 2592
rect 14969 2558 15003 2592
rect 15003 2558 15037 2592
rect 15037 2558 15071 2592
rect 15071 2558 15105 2592
rect 14927 2520 15105 2558
rect 14927 2486 14935 2520
rect 14935 2486 14969 2520
rect 14969 2486 15003 2520
rect 15003 2486 15037 2520
rect 15037 2486 15071 2520
rect 15071 2486 15105 2520
rect 14927 2448 15105 2486
rect 14927 2414 14935 2448
rect 14935 2414 14969 2448
rect 14969 2414 15003 2448
rect 15003 2414 15037 2448
rect 15037 2414 15071 2448
rect 15071 2414 15105 2448
rect 14927 2376 15105 2414
rect 14927 2342 14935 2376
rect 14935 2342 14969 2376
rect 14969 2342 15003 2376
rect 15003 2342 15037 2376
rect 15037 2342 15071 2376
rect 15071 2342 15105 2376
rect 14927 2304 15105 2342
rect 14927 2270 14935 2304
rect 14935 2270 14969 2304
rect 14969 2270 15003 2304
rect 15003 2270 15037 2304
rect 15037 2270 15071 2304
rect 15071 2270 15105 2304
rect 14927 2232 15105 2270
rect 14927 2198 14935 2232
rect 14935 2198 14969 2232
rect 14969 2198 15003 2232
rect 15003 2198 15037 2232
rect 15037 2198 15071 2232
rect 15071 2198 15105 2232
rect 14927 2160 15105 2198
rect 14927 2126 14935 2160
rect 14935 2126 14969 2160
rect 14969 2126 15003 2160
rect 15003 2126 15037 2160
rect 15037 2126 15071 2160
rect 15071 2126 15105 2160
rect 14927 2088 15105 2126
rect 14927 2054 14935 2088
rect 14935 2054 14969 2088
rect 14969 2054 15003 2088
rect 15003 2054 15037 2088
rect 15037 2054 15071 2088
rect 15071 2054 15105 2088
rect 14927 2016 15105 2054
rect 14927 1982 14935 2016
rect 14935 1982 14969 2016
rect 14969 1982 15003 2016
rect 15003 1982 15037 2016
rect 15037 1982 15071 2016
rect 15071 1982 15105 2016
rect 14927 1944 15105 1982
rect 14927 1910 14935 1944
rect 14935 1910 14969 1944
rect 14969 1910 15003 1944
rect 15003 1910 15037 1944
rect 15037 1910 15071 1944
rect 15071 1910 15105 1944
rect 14927 1872 15105 1910
rect 14927 1838 14935 1872
rect 14935 1838 14969 1872
rect 14969 1838 15003 1872
rect 15003 1838 15037 1872
rect 15037 1838 15071 1872
rect 15071 1838 15105 1872
rect 14927 1800 15105 1838
rect 14927 1766 14935 1800
rect 14935 1766 14969 1800
rect 14969 1766 15003 1800
rect 15003 1766 15037 1800
rect 15037 1766 15071 1800
rect 15071 1766 15105 1800
rect 14927 1728 15105 1766
rect 14927 1694 14935 1728
rect 14935 1694 14969 1728
rect 14969 1694 15003 1728
rect 15003 1694 15037 1728
rect 15037 1694 15071 1728
rect 15071 1694 15105 1728
rect 14927 1656 15105 1694
rect 14927 1622 14935 1656
rect 14935 1622 14969 1656
rect 14969 1622 15003 1656
rect 15003 1622 15037 1656
rect 15037 1622 15071 1656
rect 15071 1622 15105 1656
rect 14927 1584 15105 1622
rect 14927 1550 14935 1584
rect 14935 1550 14969 1584
rect 14969 1550 15003 1584
rect 15003 1550 15037 1584
rect 15037 1550 15071 1584
rect 15071 1550 15105 1584
rect 14927 1512 15105 1550
rect 14927 1478 14935 1512
rect 14935 1478 14969 1512
rect 14969 1478 15003 1512
rect 15003 1478 15037 1512
rect 15037 1478 15071 1512
rect 15071 1478 15105 1512
rect 14927 1440 15105 1478
rect 14927 1406 14935 1440
rect 14935 1406 14969 1440
rect 14969 1406 15003 1440
rect 15003 1406 15037 1440
rect 15037 1406 15071 1440
rect 15071 1406 15105 1440
rect 14927 1368 15105 1406
rect 14927 1334 14935 1368
rect 14935 1334 14969 1368
rect 14969 1334 15003 1368
rect 15003 1334 15037 1368
rect 15037 1334 15071 1368
rect 15071 1334 15105 1368
rect 14927 1296 15105 1334
rect 14927 1262 14935 1296
rect 14935 1262 14969 1296
rect 14969 1262 15003 1296
rect 15003 1262 15037 1296
rect 15037 1262 15071 1296
rect 15071 1262 15105 1296
rect 14927 1224 15105 1262
rect 14927 1190 14935 1224
rect 14935 1190 14969 1224
rect 14969 1190 15003 1224
rect 15003 1190 15037 1224
rect 15037 1190 15071 1224
rect 15071 1190 15105 1224
rect 14927 1152 15105 1190
rect 14927 1118 14935 1152
rect 14935 1118 14969 1152
rect 14969 1118 15003 1152
rect 15003 1118 15037 1152
rect 15037 1118 15071 1152
rect 15071 1118 15105 1152
rect 14927 1080 15105 1118
rect 14927 1046 14935 1080
rect 14935 1046 14969 1080
rect 14969 1046 15003 1080
rect 15003 1046 15037 1080
rect 15037 1046 15071 1080
rect 15071 1046 15105 1080
rect 14927 1008 15105 1046
rect 14927 974 14935 1008
rect 14935 974 14969 1008
rect 14969 974 15003 1008
rect 15003 974 15037 1008
rect 15037 974 15071 1008
rect 15071 974 15105 1008
rect 14927 936 15105 974
rect 14927 902 14935 936
rect 14935 902 14969 936
rect 14969 902 15003 936
rect 15003 902 15037 936
rect 15037 902 15071 936
rect 15071 902 15105 936
rect 14927 864 15105 902
rect 14927 830 14935 864
rect 14935 830 14969 864
rect 14969 830 15003 864
rect 15003 830 15037 864
rect 15037 830 15071 864
rect 15071 830 15105 864
rect 14927 792 15105 830
rect 14927 758 14935 792
rect 14935 758 14969 792
rect 14969 758 15003 792
rect 15003 758 15037 792
rect 15037 758 15071 792
rect 15071 758 15105 792
rect 14927 720 15105 758
rect 14927 686 14935 720
rect 14935 686 14969 720
rect 14969 686 15003 720
rect 15003 686 15037 720
rect 15037 686 15071 720
rect 15071 686 15105 720
rect 308 664 14886 668
rect 308 630 328 664
rect 328 630 363 664
rect 363 630 397 664
rect 397 630 432 664
rect 432 630 466 664
rect 466 630 501 664
rect 501 630 535 664
rect 535 630 570 664
rect 570 630 604 664
rect 604 630 639 664
rect 639 630 673 664
rect 673 630 708 664
rect 708 630 742 664
rect 742 630 777 664
rect 777 630 811 664
rect 811 630 846 664
rect 846 630 880 664
rect 880 630 915 664
rect 915 630 949 664
rect 949 630 984 664
rect 984 630 1018 664
rect 1018 630 1053 664
rect 1053 630 1087 664
rect 1087 630 1122 664
rect 1122 630 1156 664
rect 1156 630 1191 664
rect 1191 630 1225 664
rect 1225 630 1260 664
rect 1260 630 1294 664
rect 1294 630 1329 664
rect 1329 630 1363 664
rect 1363 630 1398 664
rect 1398 630 1432 664
rect 1432 630 1467 664
rect 1467 630 1501 664
rect 1501 630 1536 664
rect 1536 630 1570 664
rect 1570 630 1605 664
rect 1605 630 1639 664
rect 1639 630 1674 664
rect 1674 630 1708 664
rect 1708 630 1743 664
rect 1743 630 1777 664
rect 1777 630 1812 664
rect 1812 630 1846 664
rect 1846 630 1881 664
rect 1881 630 1915 664
rect 1915 630 1950 664
rect 1950 630 1984 664
rect 1984 630 2019 664
rect 2019 630 2053 664
rect 2053 630 2088 664
rect 2088 630 2122 664
rect 2122 630 2157 664
rect 2157 630 2191 664
rect 2191 630 2226 664
rect 2226 630 2260 664
rect 2260 630 2295 664
rect 2295 630 2329 664
rect 2329 630 2364 664
rect 2364 630 2398 664
rect 2398 630 2433 664
rect 2433 630 2467 664
rect 2467 630 2502 664
rect 2502 630 2536 664
rect 2536 630 2571 664
rect 2571 630 2605 664
rect 2605 630 2640 664
rect 2640 630 2674 664
rect 2674 630 2709 664
rect 2709 630 2743 664
rect 2743 630 2778 664
rect 2778 630 2812 664
rect 2812 630 2847 664
rect 2847 630 2881 664
rect 2881 630 2916 664
rect 2916 630 2950 664
rect 2950 630 2985 664
rect 2985 630 3019 664
rect 3019 630 3054 664
rect 3054 630 3088 664
rect 3088 630 3123 664
rect 3123 630 3157 664
rect 3157 630 3192 664
rect 3192 630 3226 664
rect 3226 630 3261 664
rect 3261 630 3295 664
rect 3295 630 3330 664
rect 3330 630 3364 664
rect 3364 630 3399 664
rect 3399 630 3433 664
rect 3433 630 3468 664
rect 3468 630 3502 664
rect 3502 630 3537 664
rect 3537 630 3571 664
rect 3571 630 3606 664
rect 3606 630 3640 664
rect 3640 630 3675 664
rect 3675 630 3709 664
rect 3709 630 3744 664
rect 3744 630 3778 664
rect 3778 630 3813 664
rect 3813 630 3847 664
rect 3847 630 3882 664
rect 3882 630 3916 664
rect 3916 630 3951 664
rect 3951 630 3985 664
rect 3985 630 4020 664
rect 4020 630 4054 664
rect 4054 630 4089 664
rect 4089 630 4123 664
rect 4123 630 4158 664
rect 4158 630 4192 664
rect 4192 630 4227 664
rect 4227 630 4261 664
rect 4261 630 4296 664
rect 4296 630 4330 664
rect 4330 630 4365 664
rect 4365 630 4399 664
rect 4399 630 4434 664
rect 4434 630 4468 664
rect 4468 630 4503 664
rect 4503 630 4537 664
rect 4537 630 4572 664
rect 4572 630 4606 664
rect 4606 630 4641 664
rect 4641 630 4675 664
rect 4675 630 4710 664
rect 308 596 4710 630
rect 308 562 328 596
rect 328 562 363 596
rect 363 562 397 596
rect 397 562 432 596
rect 432 562 466 596
rect 466 562 501 596
rect 501 562 535 596
rect 535 562 570 596
rect 570 562 604 596
rect 604 562 639 596
rect 639 562 673 596
rect 673 562 708 596
rect 708 562 742 596
rect 742 562 777 596
rect 777 562 811 596
rect 811 562 846 596
rect 846 562 880 596
rect 880 562 915 596
rect 915 562 949 596
rect 949 562 984 596
rect 984 562 1018 596
rect 1018 562 1053 596
rect 1053 562 1087 596
rect 1087 562 1122 596
rect 1122 562 1156 596
rect 1156 562 1191 596
rect 1191 562 1225 596
rect 1225 562 1260 596
rect 1260 562 1294 596
rect 1294 562 1329 596
rect 1329 562 1363 596
rect 1363 562 1398 596
rect 1398 562 1432 596
rect 1432 562 1467 596
rect 1467 562 1501 596
rect 1501 562 1536 596
rect 1536 562 1570 596
rect 1570 562 1605 596
rect 1605 562 1639 596
rect 1639 562 1674 596
rect 1674 562 1708 596
rect 1708 562 1743 596
rect 1743 562 1777 596
rect 1777 562 1812 596
rect 1812 562 1846 596
rect 1846 562 1881 596
rect 1881 562 1915 596
rect 1915 562 1950 596
rect 1950 562 1984 596
rect 1984 562 2019 596
rect 2019 562 2053 596
rect 2053 562 2088 596
rect 2088 562 2122 596
rect 2122 562 2157 596
rect 2157 562 2191 596
rect 2191 562 2226 596
rect 2226 562 2260 596
rect 2260 562 2295 596
rect 2295 562 2329 596
rect 2329 562 2364 596
rect 2364 562 2398 596
rect 2398 562 2433 596
rect 2433 562 2467 596
rect 2467 562 2502 596
rect 2502 562 2536 596
rect 2536 562 2571 596
rect 2571 562 2605 596
rect 2605 562 2640 596
rect 2640 562 2674 596
rect 2674 562 2709 596
rect 2709 562 2743 596
rect 2743 562 2778 596
rect 2778 562 2812 596
rect 2812 562 2847 596
rect 2847 562 2881 596
rect 2881 562 2916 596
rect 2916 562 2950 596
rect 2950 562 2985 596
rect 2985 562 3019 596
rect 3019 562 3054 596
rect 3054 562 3088 596
rect 3088 562 3123 596
rect 3123 562 3157 596
rect 3157 562 3192 596
rect 3192 562 3226 596
rect 3226 562 3261 596
rect 3261 562 3295 596
rect 3295 562 3330 596
rect 3330 562 3364 596
rect 3364 562 3399 596
rect 3399 562 3433 596
rect 3433 562 3468 596
rect 3468 562 3502 596
rect 3502 562 3537 596
rect 3537 562 3571 596
rect 3571 562 3606 596
rect 3606 562 3640 596
rect 3640 562 3675 596
rect 3675 562 3709 596
rect 3709 562 3744 596
rect 3744 562 3778 596
rect 3778 562 3813 596
rect 3813 562 3847 596
rect 3847 562 3882 596
rect 3882 562 3916 596
rect 3916 562 3951 596
rect 3951 562 3985 596
rect 3985 562 4020 596
rect 4020 562 4054 596
rect 4054 562 4089 596
rect 4089 562 4123 596
rect 4123 562 4158 596
rect 4158 562 4192 596
rect 4192 562 4227 596
rect 4227 562 4261 596
rect 4261 562 4296 596
rect 4296 562 4330 596
rect 4330 562 4365 596
rect 4365 562 4399 596
rect 4399 562 4434 596
rect 4434 562 4468 596
rect 4468 562 4503 596
rect 4503 562 4537 596
rect 4537 562 4572 596
rect 4572 562 4606 596
rect 4606 562 4641 596
rect 4641 562 4675 596
rect 4675 562 4710 596
rect 71 496 249 545
rect 308 528 4710 562
rect 308 494 328 528
rect 328 494 363 528
rect 363 494 397 528
rect 397 494 432 528
rect 432 494 466 528
rect 466 494 501 528
rect 501 494 535 528
rect 535 494 570 528
rect 570 494 604 528
rect 604 494 639 528
rect 639 494 673 528
rect 673 494 708 528
rect 708 494 742 528
rect 742 494 777 528
rect 777 494 811 528
rect 811 494 846 528
rect 846 494 880 528
rect 880 494 915 528
rect 915 494 949 528
rect 949 494 984 528
rect 984 494 1018 528
rect 1018 494 1053 528
rect 1053 494 1087 528
rect 1087 494 1122 528
rect 1122 494 1156 528
rect 1156 494 1191 528
rect 1191 494 1225 528
rect 1225 494 1260 528
rect 1260 494 1294 528
rect 1294 494 1329 528
rect 1329 494 1363 528
rect 1363 494 1398 528
rect 1398 494 1432 528
rect 1432 494 1467 528
rect 1467 494 1501 528
rect 1501 494 1536 528
rect 1536 494 1570 528
rect 1570 494 1605 528
rect 1605 494 1639 528
rect 1639 494 1674 528
rect 1674 494 1708 528
rect 1708 494 1743 528
rect 1743 494 1777 528
rect 1777 494 1812 528
rect 1812 494 1846 528
rect 1846 494 1881 528
rect 1881 494 1915 528
rect 1915 494 1950 528
rect 1950 494 1984 528
rect 1984 494 2019 528
rect 2019 494 2053 528
rect 2053 494 2088 528
rect 2088 494 2122 528
rect 2122 494 2157 528
rect 2157 494 2191 528
rect 2191 494 2226 528
rect 2226 494 2260 528
rect 2260 494 2295 528
rect 2295 494 2329 528
rect 2329 494 2364 528
rect 2364 494 2398 528
rect 2398 494 2433 528
rect 2433 494 2467 528
rect 2467 494 2502 528
rect 2502 494 2536 528
rect 2536 494 2571 528
rect 2571 494 2605 528
rect 2605 494 2640 528
rect 2640 494 2674 528
rect 2674 494 2709 528
rect 2709 494 2743 528
rect 2743 494 2778 528
rect 2778 494 2812 528
rect 2812 494 2847 528
rect 2847 494 2881 528
rect 2881 494 2916 528
rect 2916 494 2950 528
rect 2950 494 2985 528
rect 2985 494 3019 528
rect 3019 494 3054 528
rect 3054 494 3088 528
rect 3088 494 3123 528
rect 3123 494 3157 528
rect 3157 494 3192 528
rect 3192 494 3226 528
rect 3226 494 3261 528
rect 3261 494 3295 528
rect 3295 494 3330 528
rect 3330 494 3364 528
rect 3364 494 3399 528
rect 3399 494 3433 528
rect 3433 494 3468 528
rect 3468 494 3502 528
rect 3502 494 3537 528
rect 3537 494 3571 528
rect 3571 494 3606 528
rect 3606 494 3640 528
rect 3640 494 3675 528
rect 3675 494 3709 528
rect 3709 494 3744 528
rect 3744 494 3778 528
rect 3778 494 3813 528
rect 3813 494 3847 528
rect 3847 494 3882 528
rect 3882 494 3916 528
rect 3916 494 3951 528
rect 3951 494 3985 528
rect 3985 494 4020 528
rect 4020 494 4054 528
rect 4054 494 4089 528
rect 4089 494 4123 528
rect 4123 494 4158 528
rect 4158 494 4192 528
rect 4192 494 4227 528
rect 4227 494 4261 528
rect 4261 494 4296 528
rect 4296 494 4330 528
rect 4330 494 4365 528
rect 4365 494 4399 528
rect 4399 494 4434 528
rect 4434 494 4468 528
rect 4468 494 4503 528
rect 4503 494 4537 528
rect 4537 494 4572 528
rect 4572 494 4606 528
rect 4606 494 4641 528
rect 4641 494 4675 528
rect 4675 494 4710 528
rect 4710 494 14876 664
rect 14876 494 14886 664
rect 308 490 14886 494
rect 14927 648 15105 686
rect 14927 614 14935 648
rect 14935 614 14969 648
rect 14969 614 15003 648
rect 15003 614 15037 648
rect 15037 614 15071 648
rect 15071 614 15105 648
rect 14927 576 15105 614
rect 14927 542 14935 576
rect 14935 542 14969 576
rect 14969 542 15003 576
rect 15003 542 15037 576
rect 15037 542 15071 576
rect 15071 542 15105 576
rect 14927 490 15105 542
<< metal1 >>
rect 59 5426 15117 5438
rect 59 496 71 5426
rect 249 5248 308 5426
rect 14886 5420 15117 5426
rect 14886 5248 14927 5420
rect 249 5236 14927 5248
rect 249 680 261 5236
tri 261 4960 537 5236 nw
tri 14638 4960 14914 5236 ne
rect 14914 4960 14927 5236
tri 14914 4959 14915 4960 ne
tri 679 4924 691 4936 se
rect 691 4924 14512 4936
tri 575 4820 679 4924 se
rect 679 4820 767 4924
rect 575 4818 767 4820
rect 12465 4890 12504 4924
rect 12538 4890 12577 4924
rect 12611 4890 12650 4924
rect 12684 4890 12723 4924
rect 12757 4890 12796 4924
rect 12830 4890 12869 4924
rect 12903 4890 12942 4924
rect 12976 4890 13015 4924
rect 13049 4890 13088 4924
rect 13122 4890 13161 4924
rect 13195 4890 13234 4924
rect 13268 4890 13307 4924
rect 13341 4890 13380 4924
rect 13414 4890 13453 4924
rect 13487 4890 13526 4924
rect 13560 4890 13599 4924
rect 13633 4890 13672 4924
rect 13706 4890 13745 4924
rect 13779 4890 13818 4924
rect 13852 4890 13891 4924
rect 13925 4890 13964 4924
rect 13998 4890 14037 4924
rect 14071 4890 14110 4924
rect 14144 4890 14183 4924
rect 14217 4890 14256 4924
rect 14290 4890 14329 4924
rect 14363 4890 14402 4924
rect 14436 4890 14512 4924
rect 12465 4852 14512 4890
rect 12465 4818 12504 4852
rect 12538 4818 12577 4852
rect 12611 4818 12650 4852
rect 12684 4818 12723 4852
rect 12757 4818 12796 4852
rect 12830 4818 12869 4852
rect 12903 4818 12942 4852
rect 12976 4818 13015 4852
rect 13049 4818 13088 4852
rect 13122 4818 13161 4852
rect 13195 4818 13234 4852
rect 13268 4818 13307 4852
rect 13341 4818 13380 4852
rect 13414 4818 13453 4852
rect 13487 4818 13526 4852
rect 13560 4818 13599 4852
rect 13633 4818 13672 4852
rect 13706 4818 13745 4852
rect 13779 4818 13818 4852
rect 13852 4818 13891 4852
rect 13925 4818 13964 4852
rect 13998 4818 14037 4852
rect 14071 4818 14110 4852
rect 14144 4818 14183 4852
rect 14217 4818 14256 4852
rect 14290 4818 14329 4852
rect 14363 4818 14402 4852
rect 14436 4820 14512 4852
tri 14512 4820 14628 4936 sw
rect 14436 4818 14628 4820
rect 575 4806 14628 4818
rect 575 4774 980 4806
tri 980 4774 1012 4806 nw
tri 14210 4786 14230 4806 ne
rect 14230 4786 14628 4806
tri 14230 4774 14242 4786 ne
rect 14242 4774 14628 4786
rect 575 4744 733 4774
rect 575 4710 587 4744
rect 621 4710 659 4744
rect 693 4740 733 4744
rect 767 4740 946 4774
tri 946 4740 980 4774 nw
tri 14242 4740 14276 4774 ne
rect 14276 4740 14431 4774
rect 14465 4743 14628 4774
rect 14465 4740 14510 4743
rect 693 4710 915 4740
rect 575 4709 915 4710
tri 915 4709 946 4740 nw
tri 14276 4709 14307 4740 ne
rect 14307 4709 14510 4740
rect 14544 4709 14582 4743
rect 14616 4709 14628 4743
rect 575 4701 907 4709
tri 907 4701 915 4709 nw
tri 14307 4701 14315 4709 ne
rect 14315 4701 14628 4709
rect 575 4670 733 4701
rect 575 4636 587 4670
rect 621 4636 659 4670
rect 693 4667 733 4670
rect 767 4667 873 4701
tri 873 4667 907 4701 nw
tri 14315 4667 14349 4701 ne
rect 14349 4667 14431 4701
rect 14465 4670 14628 4701
rect 14465 4667 14510 4670
rect 693 4636 842 4667
tri 842 4636 873 4667 nw
tri 14349 4636 14380 4667 ne
rect 14380 4636 14510 4667
rect 14544 4636 14582 4670
rect 14616 4636 14628 4670
rect 575 4628 834 4636
tri 834 4628 842 4636 nw
tri 14380 4628 14388 4636 ne
rect 14388 4628 14628 4636
rect 575 4596 733 4628
rect 575 4562 587 4596
rect 621 4562 659 4596
rect 693 4594 733 4596
rect 767 4594 803 4628
tri 803 4597 834 4628 nw
tri 14388 4616 14400 4628 ne
rect 693 4562 803 4594
rect 575 4555 803 4562
rect 575 4522 733 4555
rect 575 4488 587 4522
rect 621 4488 659 4522
rect 693 4521 733 4522
rect 767 4521 803 4555
rect 693 4488 803 4521
rect 14400 4594 14431 4628
rect 14465 4597 14628 4628
rect 14465 4594 14510 4597
rect 14400 4563 14510 4594
rect 14544 4563 14582 4597
rect 14616 4563 14628 4597
rect 14400 4555 14628 4563
rect 14400 4521 14431 4555
rect 14465 4524 14628 4555
rect 14465 4521 14510 4524
rect 575 4482 803 4488
rect 575 4449 733 4482
rect 575 4415 587 4449
rect 621 4415 659 4449
rect 693 4448 733 4449
rect 767 4448 803 4482
rect 693 4415 803 4448
rect 575 4409 803 4415
rect 575 4376 733 4409
rect 575 4342 587 4376
rect 621 4342 659 4376
rect 693 4375 733 4376
rect 767 4375 803 4409
rect 919 4494 1049 4506
rect 919 4388 931 4494
rect 1037 4388 1049 4494
rect 919 4376 1049 4388
rect 1349 4494 1479 4506
rect 1349 4388 1361 4494
rect 1467 4388 1479 4494
rect 1349 4376 1479 4388
rect 1911 4494 2041 4506
rect 1911 4388 1923 4494
rect 2029 4388 2041 4494
rect 1911 4376 2041 4388
rect 2341 4494 2471 4506
rect 2341 4388 2353 4494
rect 2459 4388 2471 4494
rect 2341 4376 2471 4388
rect 2903 4494 3033 4506
rect 2903 4388 2915 4494
rect 3021 4388 3033 4494
rect 2903 4376 3033 4388
rect 3333 4494 3463 4506
rect 3333 4388 3345 4494
rect 3451 4388 3463 4494
rect 3333 4376 3463 4388
rect 3895 4494 4025 4506
rect 3895 4388 3907 4494
rect 4013 4388 4025 4494
rect 3895 4376 4025 4388
rect 4325 4494 4455 4506
rect 4325 4388 4337 4494
rect 4443 4388 4455 4494
rect 4325 4376 4455 4388
rect 4887 4494 5017 4506
rect 4887 4388 4899 4494
rect 5005 4388 5017 4494
rect 4887 4376 5017 4388
rect 5317 4494 5447 4506
rect 5317 4388 5329 4494
rect 5435 4388 5447 4494
rect 5317 4376 5447 4388
rect 5879 4494 6009 4506
rect 5879 4388 5891 4494
rect 5997 4388 6009 4494
rect 5879 4376 6009 4388
rect 6309 4494 6439 4506
rect 6309 4388 6321 4494
rect 6427 4388 6439 4494
rect 6309 4376 6439 4388
rect 6856 4494 6986 4506
rect 6856 4388 6868 4494
rect 6974 4388 6986 4494
rect 6856 4376 6986 4388
rect 7301 4494 7431 4506
rect 7301 4388 7313 4494
rect 7419 4388 7431 4494
rect 7301 4376 7431 4388
rect 7863 4494 7993 4506
rect 7863 4388 7875 4494
rect 7981 4388 7993 4494
rect 7863 4376 7993 4388
rect 8293 4494 8423 4506
rect 8293 4388 8305 4494
rect 8411 4388 8423 4494
rect 8293 4376 8423 4388
rect 8855 4494 8985 4506
rect 8855 4388 8867 4494
rect 8973 4388 8985 4494
rect 8855 4376 8985 4388
rect 9285 4494 9415 4506
rect 9285 4388 9297 4494
rect 9403 4388 9415 4494
rect 9285 4376 9415 4388
rect 9847 4494 9977 4506
rect 9847 4388 9859 4494
rect 9965 4388 9977 4494
rect 9847 4376 9977 4388
rect 10277 4494 10407 4506
rect 10277 4388 10289 4494
rect 10395 4388 10407 4494
rect 10277 4376 10407 4388
rect 10839 4494 10969 4506
rect 10839 4388 10851 4494
rect 10957 4388 10969 4494
rect 10839 4376 10969 4388
rect 11269 4494 11399 4506
rect 11269 4388 11281 4494
rect 11387 4388 11399 4494
rect 11269 4376 11399 4388
rect 11831 4494 11961 4506
rect 11831 4388 11843 4494
rect 11949 4388 11961 4494
rect 11831 4376 11961 4388
rect 12261 4494 12391 4506
rect 12261 4388 12273 4494
rect 12379 4388 12391 4494
rect 12261 4376 12391 4388
rect 12823 4494 12953 4506
rect 12823 4388 12835 4494
rect 12941 4388 12953 4494
rect 12823 4376 12953 4388
rect 13253 4494 13383 4506
rect 13253 4388 13265 4494
rect 13371 4388 13383 4494
rect 13253 4376 13383 4388
rect 13815 4494 13945 4506
rect 13815 4388 13827 4494
rect 13933 4388 13945 4494
rect 13815 4376 13945 4388
rect 14173 4494 14303 4506
rect 14173 4388 14185 4494
rect 14291 4388 14303 4494
rect 14173 4376 14303 4388
rect 14400 4490 14510 4521
rect 14544 4490 14582 4524
rect 14616 4490 14628 4524
rect 14400 4482 14628 4490
rect 14400 4448 14431 4482
rect 14465 4451 14628 4482
rect 14465 4448 14510 4451
rect 14400 4417 14510 4448
rect 14544 4417 14582 4451
rect 14616 4417 14628 4451
rect 14400 4409 14628 4417
rect 693 4342 803 4375
rect 575 4336 803 4342
rect 575 4303 733 4336
rect 575 4269 587 4303
rect 621 4269 659 4303
rect 693 4302 733 4303
rect 767 4302 803 4336
rect 693 4269 803 4302
rect 575 4263 803 4269
rect 575 4230 733 4263
rect 575 4196 587 4230
rect 621 4196 659 4230
rect 693 4229 733 4230
rect 767 4229 803 4263
rect 693 4196 803 4229
rect 575 4190 803 4196
rect 575 4157 733 4190
rect 575 4123 587 4157
rect 621 4123 659 4157
rect 693 4156 733 4157
rect 767 4156 803 4190
rect 693 4123 803 4156
rect 575 4117 803 4123
rect 575 4084 733 4117
rect 575 4068 587 4084
rect 621 4068 659 4084
rect 693 4083 733 4084
rect 767 4083 803 4117
rect 693 4068 803 4083
rect 14400 4375 14431 4409
rect 14465 4378 14628 4409
rect 14465 4375 14510 4378
rect 14400 4344 14510 4375
rect 14544 4344 14582 4378
rect 14616 4344 14628 4378
rect 14400 4336 14628 4344
rect 14400 4302 14431 4336
rect 14465 4305 14628 4336
rect 14465 4302 14510 4305
rect 14400 4271 14510 4302
rect 14544 4271 14582 4305
rect 14616 4271 14628 4305
rect 14400 4263 14628 4271
rect 14400 4229 14431 4263
rect 14465 4232 14628 4263
rect 14465 4229 14510 4232
rect 14400 4198 14510 4229
rect 14544 4198 14582 4232
rect 14616 4198 14628 4232
rect 14400 4190 14628 4198
rect 14400 4156 14431 4190
rect 14465 4159 14628 4190
rect 14465 4156 14510 4159
rect 14400 4125 14510 4156
rect 14544 4125 14582 4159
rect 14616 4125 14628 4159
rect 14400 4117 14628 4125
rect 14400 4083 14431 4117
rect 14465 4086 14628 4117
rect 14465 4083 14510 4086
rect 627 4050 659 4068
rect 627 4016 663 4050
rect 715 4044 751 4068
rect 715 4016 733 4044
rect 575 4011 733 4016
rect 575 4004 587 4011
rect 621 4004 659 4011
rect 693 4010 733 4011
rect 767 4010 803 4016
rect 693 4004 803 4010
rect 627 3977 659 4004
rect 627 3952 663 3977
rect 715 3971 751 4004
rect 715 3952 733 3971
rect 575 3940 733 3952
rect 767 3940 803 3952
rect 627 3938 663 3940
rect 627 3904 659 3938
rect 715 3937 733 3940
rect 627 3888 663 3904
rect 715 3898 751 3937
rect 715 3888 733 3898
rect 575 3876 733 3888
rect 767 3876 803 3888
rect 627 3865 663 3876
rect 627 3831 659 3865
rect 715 3864 733 3876
rect 627 3824 663 3831
rect 715 3825 751 3864
rect 715 3824 733 3825
rect 575 3812 733 3824
rect 767 3812 803 3824
rect 627 3792 663 3812
rect 627 3760 659 3792
rect 715 3791 733 3812
rect 715 3760 751 3791
rect 575 3758 587 3760
rect 621 3758 659 3760
rect 693 3758 803 3760
rect 575 3752 803 3758
rect 575 3748 733 3752
rect 767 3748 803 3752
rect 627 3719 663 3748
rect 627 3696 659 3719
rect 715 3718 733 3748
rect 715 3696 751 3718
rect 575 3685 587 3696
rect 621 3685 659 3696
rect 693 3685 803 3696
rect 575 3684 803 3685
rect 627 3646 663 3684
rect 715 3679 751 3684
rect 627 3632 659 3646
rect 715 3645 733 3679
rect 715 3632 751 3645
rect 575 3620 587 3632
rect 621 3620 659 3632
rect 693 3620 803 3632
rect 627 3612 659 3620
rect 627 3573 663 3612
rect 715 3606 751 3620
rect 627 3568 659 3573
rect 715 3572 733 3606
rect 715 3568 751 3572
rect 575 3556 587 3568
rect 621 3556 659 3568
rect 693 3556 803 3568
rect 627 3539 659 3556
rect 627 3504 663 3539
rect 715 3533 751 3556
rect 715 3504 733 3533
rect 575 3500 733 3504
rect 575 3492 587 3500
rect 621 3492 659 3500
rect 693 3499 733 3500
rect 767 3499 803 3504
rect 693 3492 803 3499
rect 627 3466 659 3492
rect 627 3440 663 3466
rect 715 3460 751 3492
rect 715 3440 733 3460
rect 575 3428 733 3440
rect 767 3428 803 3440
rect 627 3427 663 3428
rect 627 3393 659 3427
rect 715 3426 733 3428
rect 627 3376 663 3393
rect 715 3387 751 3426
rect 715 3376 733 3387
rect 575 3364 733 3376
rect 767 3364 803 3376
rect 627 3354 663 3364
rect 627 3320 659 3354
rect 715 3353 733 3364
rect 627 3312 663 3320
rect 715 3314 751 3353
rect 715 3312 733 3314
rect 575 3300 733 3312
rect 767 3300 803 3312
rect 627 3281 663 3300
rect 627 3248 659 3281
rect 715 3280 733 3300
rect 715 3248 751 3280
rect 575 3247 587 3248
rect 621 3247 659 3248
rect 693 3247 803 3248
rect 575 3241 803 3247
rect 575 3236 733 3241
rect 767 3236 803 3241
rect 627 3208 663 3236
rect 627 3184 659 3208
rect 715 3207 733 3236
rect 715 3184 751 3207
rect 575 3174 587 3184
rect 621 3174 659 3184
rect 693 3174 803 3184
rect 575 3172 803 3174
rect 627 3135 663 3172
rect 715 3168 751 3172
rect 627 3120 659 3135
rect 715 3134 733 3168
rect 715 3120 751 3134
rect 575 3108 587 3120
rect 621 3108 659 3120
rect 693 3108 803 3120
rect 627 3101 659 3108
rect 627 3062 663 3101
rect 715 3095 751 3108
rect 627 3056 659 3062
rect 715 3061 733 3095
rect 715 3056 751 3061
rect 575 3044 587 3056
rect 621 3044 659 3056
rect 693 3044 803 3056
rect 627 3028 659 3044
rect 627 2992 663 3028
rect 715 3022 751 3044
rect 715 2992 733 3022
rect 575 2989 733 2992
rect 575 2979 587 2989
rect 621 2979 659 2989
rect 693 2988 733 2989
rect 767 2988 803 2992
rect 693 2979 803 2988
rect 627 2955 659 2979
rect 627 2927 663 2955
rect 715 2949 751 2979
rect 715 2927 733 2949
rect 575 2916 733 2927
rect 575 2882 587 2916
rect 621 2882 659 2916
rect 693 2915 733 2916
rect 767 2915 803 2927
rect 693 2882 803 2915
rect 575 2876 803 2882
rect 575 2843 733 2876
rect 575 2809 587 2843
rect 621 2809 659 2843
rect 693 2842 733 2843
rect 767 2842 803 2876
rect 693 2809 803 2842
rect 575 2803 803 2809
rect 575 2770 733 2803
rect 575 2736 587 2770
rect 621 2736 659 2770
rect 693 2769 733 2770
rect 767 2769 803 2803
rect 693 2736 803 2769
rect 575 2730 803 2736
rect 575 2697 733 2730
rect 575 2663 587 2697
rect 621 2663 659 2697
rect 693 2696 733 2697
rect 767 2696 803 2730
rect 693 2663 803 2696
rect 575 2657 803 2663
rect 575 2624 733 2657
rect 575 2590 587 2624
rect 621 2590 659 2624
rect 693 2623 733 2624
rect 767 2623 803 2657
rect 693 2590 803 2623
rect 575 2584 803 2590
rect 575 2551 733 2584
rect 575 2517 587 2551
rect 621 2517 659 2551
rect 693 2550 733 2551
rect 767 2550 803 2584
rect 693 2517 803 2550
rect 575 2511 803 2517
rect 575 2478 733 2511
rect 575 2444 587 2478
rect 621 2444 659 2478
rect 693 2477 733 2478
rect 767 2477 803 2511
rect 693 2444 803 2477
rect 575 2438 803 2444
rect 575 2405 733 2438
rect 575 2371 587 2405
rect 621 2371 659 2405
rect 693 2404 733 2405
rect 767 2404 803 2438
rect 693 2371 803 2404
rect 575 2365 803 2371
rect 575 2332 733 2365
rect 575 2298 587 2332
rect 621 2298 659 2332
rect 693 2331 733 2332
rect 767 2331 803 2365
rect 693 2298 803 2331
rect 575 2292 803 2298
rect 575 2259 733 2292
rect 575 2225 587 2259
rect 621 2225 659 2259
rect 693 2258 733 2259
rect 767 2258 803 2292
rect 693 2225 803 2258
rect 575 2219 803 2225
rect 575 2186 733 2219
rect 575 2152 587 2186
rect 621 2152 659 2186
rect 693 2185 733 2186
rect 767 2185 803 2219
rect 693 2152 803 2185
rect 575 2146 803 2152
rect 575 2113 733 2146
rect 575 2079 587 2113
rect 621 2079 659 2113
rect 693 2112 733 2113
rect 767 2112 803 2146
rect 693 2079 803 2112
rect 575 2073 803 2079
rect 575 2040 733 2073
rect 575 2006 587 2040
rect 621 2006 659 2040
rect 693 2039 733 2040
rect 767 2039 803 2073
rect 693 2006 803 2039
rect 575 2000 803 2006
rect 575 1967 733 2000
rect 575 1933 587 1967
rect 621 1933 659 1967
rect 693 1966 733 1967
rect 767 1966 803 2000
rect 693 1933 803 1966
rect 575 1927 803 1933
rect 575 1894 733 1927
rect 575 1860 587 1894
rect 621 1860 659 1894
rect 693 1893 733 1894
rect 767 1893 803 1927
rect 693 1860 803 1893
rect 575 1854 803 1860
rect 575 1821 733 1854
rect 575 1787 587 1821
rect 621 1787 659 1821
rect 693 1820 733 1821
rect 767 1820 803 1854
rect 693 1787 803 1820
rect 575 1781 803 1787
rect 575 1748 733 1781
rect 575 1714 587 1748
rect 621 1714 659 1748
rect 693 1747 733 1748
rect 767 1747 803 1781
rect 693 1714 803 1747
rect 575 1708 803 1714
rect 575 1675 733 1708
rect 575 1641 587 1675
rect 621 1641 659 1675
rect 693 1674 733 1675
rect 767 1674 803 1708
rect 693 1641 803 1674
rect 575 1635 803 1641
rect 575 1602 733 1635
rect 575 1568 587 1602
rect 621 1568 659 1602
rect 693 1601 733 1602
rect 767 1601 803 1635
rect 693 1568 803 1601
rect 575 1562 803 1568
rect 575 1529 733 1562
rect 575 1495 587 1529
rect 621 1495 659 1529
rect 693 1528 733 1529
rect 767 1528 803 1562
rect 693 1495 803 1528
rect 575 1489 803 1495
rect 575 1455 733 1489
rect 767 1455 803 1489
rect 1103 4062 1295 4074
rect 1103 4028 1110 4062
rect 1144 4028 1182 4062
rect 1216 4028 1254 4062
rect 1288 4028 1295 4062
rect 1103 3988 1295 4028
rect 1103 3954 1110 3988
rect 1144 3954 1182 3988
rect 1216 3954 1254 3988
rect 1288 3954 1295 3988
rect 1103 3914 1295 3954
rect 1103 3880 1110 3914
rect 1144 3880 1182 3914
rect 1216 3880 1254 3914
rect 1288 3880 1295 3914
rect 1103 3840 1295 3880
rect 1103 3806 1110 3840
rect 1144 3806 1182 3840
rect 1216 3806 1254 3840
rect 1288 3806 1295 3840
rect 1103 3766 1295 3806
rect 1103 3732 1110 3766
rect 1144 3732 1182 3766
rect 1216 3732 1254 3766
rect 1288 3732 1295 3766
rect 1103 3692 1295 3732
rect 1103 3658 1110 3692
rect 1144 3658 1182 3692
rect 1216 3658 1254 3692
rect 1288 3658 1295 3692
rect 1103 3618 1295 3658
rect 1103 3584 1110 3618
rect 1144 3584 1182 3618
rect 1216 3584 1254 3618
rect 1288 3584 1295 3618
rect 1103 3544 1295 3584
rect 1103 3510 1110 3544
rect 1144 3510 1182 3544
rect 1216 3510 1254 3544
rect 1288 3510 1295 3544
rect 1103 3470 1295 3510
rect 1103 3436 1110 3470
rect 1144 3436 1182 3470
rect 1216 3436 1254 3470
rect 1288 3436 1295 3470
rect 1103 3396 1295 3436
rect 1103 3362 1110 3396
rect 1144 3362 1182 3396
rect 1216 3362 1254 3396
rect 1288 3362 1295 3396
rect 1103 3322 1295 3362
rect 1103 3288 1110 3322
rect 1144 3288 1182 3322
rect 1216 3288 1254 3322
rect 1288 3288 1295 3322
rect 1103 3248 1295 3288
rect 1103 3214 1110 3248
rect 1144 3214 1182 3248
rect 1216 3214 1254 3248
rect 1288 3214 1295 3248
rect 1103 3174 1295 3214
rect 1103 3140 1110 3174
rect 1144 3140 1182 3174
rect 1216 3140 1254 3174
rect 1288 3140 1295 3174
rect 1103 3100 1295 3140
rect 1103 3066 1110 3100
rect 1144 3066 1182 3100
rect 1216 3066 1254 3100
rect 1288 3066 1295 3100
rect 1103 3026 1295 3066
rect 1103 2992 1110 3026
rect 1144 2992 1182 3026
rect 1216 2992 1254 3026
rect 1288 2992 1295 3026
rect 1103 2952 1295 2992
rect 1103 2918 1110 2952
rect 1144 2918 1182 2952
rect 1216 2918 1254 2952
rect 1288 2918 1295 2952
rect 1103 2878 1295 2918
rect 1103 2844 1110 2878
rect 1144 2844 1182 2878
rect 1216 2844 1254 2878
rect 1288 2844 1295 2878
rect 1103 2804 1295 2844
rect 1103 2770 1110 2804
rect 1144 2770 1182 2804
rect 1216 2770 1254 2804
rect 1288 2770 1295 2804
rect 1103 2730 1295 2770
rect 1103 2696 1110 2730
rect 1144 2696 1182 2730
rect 1216 2696 1254 2730
rect 1288 2696 1295 2730
rect 1103 2656 1295 2696
rect 1103 2622 1110 2656
rect 1144 2622 1182 2656
rect 1216 2622 1254 2656
rect 1288 2622 1295 2656
rect 1103 2614 1295 2622
rect 1103 1538 1109 2614
rect 1289 1538 1295 2614
rect 1103 1525 1110 1538
rect 1144 1525 1182 1538
rect 1216 1525 1254 1538
rect 1288 1525 1295 1538
rect 1103 1473 1109 1525
rect 1161 1473 1173 1525
rect 1225 1473 1237 1525
rect 1289 1473 1295 1525
rect 1103 1467 1295 1473
rect 1599 4068 1791 4074
rect 1599 2992 1605 4068
rect 1785 2992 1791 4068
rect 1599 2979 1606 2992
rect 1784 2979 1791 2992
rect 1599 2927 1605 2979
rect 1785 2927 1791 2979
rect 1599 2574 1606 2927
rect 1784 2574 1791 2927
rect 1599 2535 1791 2574
rect 1599 2501 1606 2535
rect 1640 2501 1678 2535
rect 1712 2501 1750 2535
rect 1784 2501 1791 2535
rect 1599 2461 1791 2501
rect 1599 2449 1678 2461
rect 1712 2449 1791 2461
rect 1599 1479 1606 2449
rect 1640 1479 1750 1491
rect 1784 1479 1791 2449
rect 1599 1467 1791 1479
rect 2095 4062 2287 4074
rect 2095 4028 2102 4062
rect 2136 4028 2174 4062
rect 2208 4028 2246 4062
rect 2280 4028 2287 4062
rect 2095 3988 2287 4028
rect 2095 3954 2102 3988
rect 2136 3954 2174 3988
rect 2208 3954 2246 3988
rect 2280 3954 2287 3988
rect 2095 3914 2287 3954
rect 2095 3880 2102 3914
rect 2136 3880 2174 3914
rect 2208 3880 2246 3914
rect 2280 3880 2287 3914
rect 2095 3840 2287 3880
rect 2095 3806 2102 3840
rect 2136 3806 2174 3840
rect 2208 3806 2246 3840
rect 2280 3806 2287 3840
rect 2095 3766 2287 3806
rect 2095 3732 2102 3766
rect 2136 3732 2174 3766
rect 2208 3732 2246 3766
rect 2280 3732 2287 3766
rect 2095 3692 2287 3732
rect 2095 3658 2102 3692
rect 2136 3658 2174 3692
rect 2208 3658 2246 3692
rect 2280 3658 2287 3692
rect 2095 3618 2287 3658
rect 2095 3584 2102 3618
rect 2136 3584 2174 3618
rect 2208 3584 2246 3618
rect 2280 3584 2287 3618
rect 2095 3544 2287 3584
rect 2095 3510 2102 3544
rect 2136 3510 2174 3544
rect 2208 3510 2246 3544
rect 2280 3510 2287 3544
rect 2095 3470 2287 3510
rect 2095 3436 2102 3470
rect 2136 3436 2174 3470
rect 2208 3436 2246 3470
rect 2280 3436 2287 3470
rect 2095 3396 2287 3436
rect 2095 3362 2102 3396
rect 2136 3362 2174 3396
rect 2208 3362 2246 3396
rect 2280 3362 2287 3396
rect 2095 3322 2287 3362
rect 2095 3288 2102 3322
rect 2136 3288 2174 3322
rect 2208 3288 2246 3322
rect 2280 3288 2287 3322
rect 2095 3248 2287 3288
rect 2095 3214 2102 3248
rect 2136 3214 2174 3248
rect 2208 3214 2246 3248
rect 2280 3214 2287 3248
rect 2095 3174 2287 3214
rect 2095 3140 2102 3174
rect 2136 3140 2174 3174
rect 2208 3140 2246 3174
rect 2280 3140 2287 3174
rect 2095 3100 2287 3140
rect 2095 3066 2102 3100
rect 2136 3066 2174 3100
rect 2208 3066 2246 3100
rect 2280 3066 2287 3100
rect 2095 3026 2287 3066
rect 2095 2992 2102 3026
rect 2136 2992 2174 3026
rect 2208 2992 2246 3026
rect 2280 2992 2287 3026
rect 2095 2952 2287 2992
rect 2095 2918 2102 2952
rect 2136 2918 2174 2952
rect 2208 2918 2246 2952
rect 2280 2918 2287 2952
rect 2095 2878 2287 2918
rect 2095 2844 2102 2878
rect 2136 2844 2174 2878
rect 2208 2844 2246 2878
rect 2280 2844 2287 2878
rect 2095 2804 2287 2844
rect 2095 2770 2102 2804
rect 2136 2770 2174 2804
rect 2208 2770 2246 2804
rect 2280 2770 2287 2804
rect 2095 2730 2287 2770
rect 2095 2696 2102 2730
rect 2136 2696 2174 2730
rect 2208 2696 2246 2730
rect 2280 2696 2287 2730
rect 2095 2656 2287 2696
rect 2095 2622 2102 2656
rect 2136 2622 2174 2656
rect 2208 2622 2246 2656
rect 2280 2622 2287 2656
rect 2095 2614 2287 2622
rect 2095 1538 2101 2614
rect 2281 1538 2287 2614
rect 2095 1525 2102 1538
rect 2136 1525 2174 1538
rect 2208 1525 2246 1538
rect 2280 1525 2287 1538
rect 2095 1473 2101 1525
rect 2153 1473 2165 1525
rect 2217 1473 2229 1525
rect 2281 1473 2287 1525
rect 2095 1467 2287 1473
rect 2591 4068 2783 4074
rect 2591 2992 2597 4068
rect 2777 2992 2783 4068
rect 2591 2979 2598 2992
rect 2776 2979 2783 2992
rect 2591 2927 2597 2979
rect 2777 2927 2783 2979
rect 2591 2574 2598 2927
rect 2776 2574 2783 2927
rect 2591 2535 2783 2574
rect 2591 2501 2598 2535
rect 2632 2501 2670 2535
rect 2704 2501 2742 2535
rect 2776 2501 2783 2535
rect 2591 2461 2783 2501
rect 2591 2449 2670 2461
rect 2704 2449 2783 2461
rect 2591 1479 2598 2449
rect 2632 1479 2742 1491
rect 2776 1479 2783 2449
rect 2591 1467 2783 1479
rect 3087 4062 3279 4074
rect 3087 4028 3094 4062
rect 3128 4028 3166 4062
rect 3200 4028 3238 4062
rect 3272 4028 3279 4062
rect 3087 3988 3279 4028
rect 3087 3954 3094 3988
rect 3128 3954 3166 3988
rect 3200 3954 3238 3988
rect 3272 3954 3279 3988
rect 3087 3914 3279 3954
rect 3087 3880 3094 3914
rect 3128 3880 3166 3914
rect 3200 3880 3238 3914
rect 3272 3880 3279 3914
rect 3087 3840 3279 3880
rect 3087 3806 3094 3840
rect 3128 3806 3166 3840
rect 3200 3806 3238 3840
rect 3272 3806 3279 3840
rect 3087 3766 3279 3806
rect 3087 3732 3094 3766
rect 3128 3732 3166 3766
rect 3200 3732 3238 3766
rect 3272 3732 3279 3766
rect 3087 3692 3279 3732
rect 3087 3658 3094 3692
rect 3128 3658 3166 3692
rect 3200 3658 3238 3692
rect 3272 3658 3279 3692
rect 3087 3618 3279 3658
rect 3087 3584 3094 3618
rect 3128 3584 3166 3618
rect 3200 3584 3238 3618
rect 3272 3584 3279 3618
rect 3087 3544 3279 3584
rect 3087 3510 3094 3544
rect 3128 3510 3166 3544
rect 3200 3510 3238 3544
rect 3272 3510 3279 3544
rect 3087 3470 3279 3510
rect 3087 3436 3094 3470
rect 3128 3436 3166 3470
rect 3200 3436 3238 3470
rect 3272 3436 3279 3470
rect 3087 3396 3279 3436
rect 3087 3362 3094 3396
rect 3128 3362 3166 3396
rect 3200 3362 3238 3396
rect 3272 3362 3279 3396
rect 3087 3322 3279 3362
rect 3087 3288 3094 3322
rect 3128 3288 3166 3322
rect 3200 3288 3238 3322
rect 3272 3288 3279 3322
rect 3087 3248 3279 3288
rect 3087 3214 3094 3248
rect 3128 3214 3166 3248
rect 3200 3214 3238 3248
rect 3272 3214 3279 3248
rect 3087 3174 3279 3214
rect 3087 3140 3094 3174
rect 3128 3140 3166 3174
rect 3200 3140 3238 3174
rect 3272 3140 3279 3174
rect 3087 3100 3279 3140
rect 3087 3066 3094 3100
rect 3128 3066 3166 3100
rect 3200 3066 3238 3100
rect 3272 3066 3279 3100
rect 3087 3026 3279 3066
rect 3087 2992 3094 3026
rect 3128 2992 3166 3026
rect 3200 2992 3238 3026
rect 3272 2992 3279 3026
rect 3087 2952 3279 2992
rect 3087 2918 3094 2952
rect 3128 2918 3166 2952
rect 3200 2918 3238 2952
rect 3272 2918 3279 2952
rect 3087 2878 3279 2918
rect 3087 2844 3094 2878
rect 3128 2844 3166 2878
rect 3200 2844 3238 2878
rect 3272 2844 3279 2878
rect 3087 2804 3279 2844
rect 3087 2770 3094 2804
rect 3128 2770 3166 2804
rect 3200 2770 3238 2804
rect 3272 2770 3279 2804
rect 3087 2730 3279 2770
rect 3087 2696 3094 2730
rect 3128 2696 3166 2730
rect 3200 2696 3238 2730
rect 3272 2696 3279 2730
rect 3087 2656 3279 2696
rect 3087 2622 3094 2656
rect 3128 2622 3166 2656
rect 3200 2622 3238 2656
rect 3272 2622 3279 2656
rect 3087 2614 3279 2622
rect 3087 1538 3093 2614
rect 3273 1538 3279 2614
rect 3087 1525 3094 1538
rect 3128 1525 3166 1538
rect 3200 1525 3238 1538
rect 3272 1525 3279 1538
rect 3087 1473 3093 1525
rect 3145 1473 3157 1525
rect 3209 1473 3221 1525
rect 3273 1473 3279 1525
rect 3087 1467 3279 1473
rect 3583 4068 3775 4074
rect 3583 2992 3589 4068
rect 3769 2992 3775 4068
rect 3583 2979 3590 2992
rect 3768 2979 3775 2992
rect 3583 2927 3589 2979
rect 3769 2927 3775 2979
rect 3583 2574 3590 2927
rect 3768 2574 3775 2927
rect 3583 2535 3775 2574
rect 3583 2501 3590 2535
rect 3624 2501 3662 2535
rect 3696 2501 3734 2535
rect 3768 2501 3775 2535
rect 3583 2461 3775 2501
rect 3583 2449 3662 2461
rect 3696 2449 3775 2461
rect 3583 1479 3590 2449
rect 3624 1479 3734 1491
rect 3768 1479 3775 2449
rect 3583 1467 3775 1479
rect 4079 4062 4271 4074
rect 4079 4028 4086 4062
rect 4120 4028 4158 4062
rect 4192 4028 4230 4062
rect 4264 4028 4271 4062
rect 4079 3988 4271 4028
rect 4079 3954 4086 3988
rect 4120 3954 4158 3988
rect 4192 3954 4230 3988
rect 4264 3954 4271 3988
rect 4079 3914 4271 3954
rect 4079 3880 4086 3914
rect 4120 3880 4158 3914
rect 4192 3880 4230 3914
rect 4264 3880 4271 3914
rect 4079 3840 4271 3880
rect 4079 3806 4086 3840
rect 4120 3806 4158 3840
rect 4192 3806 4230 3840
rect 4264 3806 4271 3840
rect 4079 3766 4271 3806
rect 4079 3732 4086 3766
rect 4120 3732 4158 3766
rect 4192 3732 4230 3766
rect 4264 3732 4271 3766
rect 4079 3692 4271 3732
rect 4079 3658 4086 3692
rect 4120 3658 4158 3692
rect 4192 3658 4230 3692
rect 4264 3658 4271 3692
rect 4079 3618 4271 3658
rect 4079 3584 4086 3618
rect 4120 3584 4158 3618
rect 4192 3584 4230 3618
rect 4264 3584 4271 3618
rect 4079 3544 4271 3584
rect 4079 3510 4086 3544
rect 4120 3510 4158 3544
rect 4192 3510 4230 3544
rect 4264 3510 4271 3544
rect 4079 3470 4271 3510
rect 4079 3436 4086 3470
rect 4120 3436 4158 3470
rect 4192 3436 4230 3470
rect 4264 3436 4271 3470
rect 4079 3396 4271 3436
rect 4079 3362 4086 3396
rect 4120 3362 4158 3396
rect 4192 3362 4230 3396
rect 4264 3362 4271 3396
rect 4079 3322 4271 3362
rect 4079 3288 4086 3322
rect 4120 3288 4158 3322
rect 4192 3288 4230 3322
rect 4264 3288 4271 3322
rect 4079 3248 4271 3288
rect 4079 3214 4086 3248
rect 4120 3214 4158 3248
rect 4192 3214 4230 3248
rect 4264 3214 4271 3248
rect 4079 3174 4271 3214
rect 4079 3140 4086 3174
rect 4120 3140 4158 3174
rect 4192 3140 4230 3174
rect 4264 3140 4271 3174
rect 4079 3100 4271 3140
rect 4079 3066 4086 3100
rect 4120 3066 4158 3100
rect 4192 3066 4230 3100
rect 4264 3066 4271 3100
rect 4079 3026 4271 3066
rect 4079 2992 4086 3026
rect 4120 2992 4158 3026
rect 4192 2992 4230 3026
rect 4264 2992 4271 3026
rect 4079 2952 4271 2992
rect 4079 2918 4086 2952
rect 4120 2918 4158 2952
rect 4192 2918 4230 2952
rect 4264 2918 4271 2952
rect 4079 2878 4271 2918
rect 4079 2844 4086 2878
rect 4120 2844 4158 2878
rect 4192 2844 4230 2878
rect 4264 2844 4271 2878
rect 4079 2804 4271 2844
rect 4079 2770 4086 2804
rect 4120 2770 4158 2804
rect 4192 2770 4230 2804
rect 4264 2770 4271 2804
rect 4079 2730 4271 2770
rect 4079 2696 4086 2730
rect 4120 2696 4158 2730
rect 4192 2696 4230 2730
rect 4264 2696 4271 2730
rect 4079 2656 4271 2696
rect 4079 2622 4086 2656
rect 4120 2622 4158 2656
rect 4192 2622 4230 2656
rect 4264 2622 4271 2656
rect 4079 2614 4271 2622
rect 4079 1538 4085 2614
rect 4265 1538 4271 2614
rect 4079 1525 4086 1538
rect 4120 1525 4158 1538
rect 4192 1525 4230 1538
rect 4264 1525 4271 1538
rect 4079 1473 4085 1525
rect 4137 1473 4149 1525
rect 4201 1473 4213 1525
rect 4265 1473 4271 1525
rect 4079 1467 4271 1473
rect 4575 4068 4767 4074
rect 4575 2992 4581 4068
rect 4761 2992 4767 4068
rect 4575 2979 4582 2992
rect 4760 2979 4767 2992
rect 4575 2927 4581 2979
rect 4761 2927 4767 2979
rect 4575 2574 4582 2927
rect 4760 2574 4767 2927
rect 4575 2535 4767 2574
rect 4575 2501 4582 2535
rect 4616 2501 4654 2535
rect 4688 2501 4726 2535
rect 4760 2501 4767 2535
rect 4575 2461 4767 2501
rect 4575 2449 4654 2461
rect 4688 2449 4767 2461
rect 4575 1479 4582 2449
rect 4616 1479 4726 1491
rect 4760 1479 4767 2449
rect 4575 1467 4767 1479
rect 5071 4062 5263 4074
rect 5071 4028 5078 4062
rect 5112 4028 5150 4062
rect 5184 4028 5222 4062
rect 5256 4028 5263 4062
rect 5071 3988 5263 4028
rect 5071 3954 5078 3988
rect 5112 3954 5150 3988
rect 5184 3954 5222 3988
rect 5256 3954 5263 3988
rect 5071 3914 5263 3954
rect 5071 3880 5078 3914
rect 5112 3880 5150 3914
rect 5184 3880 5222 3914
rect 5256 3880 5263 3914
rect 5071 3840 5263 3880
rect 5071 3806 5078 3840
rect 5112 3806 5150 3840
rect 5184 3806 5222 3840
rect 5256 3806 5263 3840
rect 5071 3766 5263 3806
rect 5071 3732 5078 3766
rect 5112 3732 5150 3766
rect 5184 3732 5222 3766
rect 5256 3732 5263 3766
rect 5071 3692 5263 3732
rect 5071 3658 5078 3692
rect 5112 3658 5150 3692
rect 5184 3658 5222 3692
rect 5256 3658 5263 3692
rect 5071 3618 5263 3658
rect 5071 3584 5078 3618
rect 5112 3584 5150 3618
rect 5184 3584 5222 3618
rect 5256 3584 5263 3618
rect 5071 3544 5263 3584
rect 5071 3510 5078 3544
rect 5112 3510 5150 3544
rect 5184 3510 5222 3544
rect 5256 3510 5263 3544
rect 5071 3470 5263 3510
rect 5071 3436 5078 3470
rect 5112 3436 5150 3470
rect 5184 3436 5222 3470
rect 5256 3436 5263 3470
rect 5071 3396 5263 3436
rect 5071 3362 5078 3396
rect 5112 3362 5150 3396
rect 5184 3362 5222 3396
rect 5256 3362 5263 3396
rect 5071 3322 5263 3362
rect 5071 3288 5078 3322
rect 5112 3288 5150 3322
rect 5184 3288 5222 3322
rect 5256 3288 5263 3322
rect 5071 3248 5263 3288
rect 5071 3214 5078 3248
rect 5112 3214 5150 3248
rect 5184 3214 5222 3248
rect 5256 3214 5263 3248
rect 5071 3174 5263 3214
rect 5071 3140 5078 3174
rect 5112 3140 5150 3174
rect 5184 3140 5222 3174
rect 5256 3140 5263 3174
rect 5071 3100 5263 3140
rect 5071 3066 5078 3100
rect 5112 3066 5150 3100
rect 5184 3066 5222 3100
rect 5256 3066 5263 3100
rect 5071 3026 5263 3066
rect 5071 2992 5078 3026
rect 5112 2992 5150 3026
rect 5184 2992 5222 3026
rect 5256 2992 5263 3026
rect 5071 2952 5263 2992
rect 5071 2918 5078 2952
rect 5112 2918 5150 2952
rect 5184 2918 5222 2952
rect 5256 2918 5263 2952
rect 5071 2878 5263 2918
rect 5071 2844 5078 2878
rect 5112 2844 5150 2878
rect 5184 2844 5222 2878
rect 5256 2844 5263 2878
rect 5071 2804 5263 2844
rect 5071 2770 5078 2804
rect 5112 2770 5150 2804
rect 5184 2770 5222 2804
rect 5256 2770 5263 2804
rect 5071 2730 5263 2770
rect 5071 2696 5078 2730
rect 5112 2696 5150 2730
rect 5184 2696 5222 2730
rect 5256 2696 5263 2730
rect 5071 2656 5263 2696
rect 5071 2622 5078 2656
rect 5112 2622 5150 2656
rect 5184 2622 5222 2656
rect 5256 2622 5263 2656
rect 5071 2614 5263 2622
rect 5071 1538 5077 2614
rect 5257 1538 5263 2614
rect 5071 1525 5078 1538
rect 5112 1525 5150 1538
rect 5184 1525 5222 1538
rect 5256 1525 5263 1538
rect 5071 1473 5077 1525
rect 5129 1473 5141 1525
rect 5193 1473 5205 1525
rect 5257 1473 5263 1525
rect 5071 1467 5263 1473
rect 5567 4068 5759 4074
rect 5567 2992 5573 4068
rect 5753 2992 5759 4068
rect 5567 2979 5574 2992
rect 5752 2979 5759 2992
rect 5567 2927 5573 2979
rect 5753 2927 5759 2979
rect 5567 2574 5574 2927
rect 5752 2574 5759 2927
rect 5567 2535 5759 2574
rect 5567 2501 5574 2535
rect 5608 2501 5646 2535
rect 5680 2501 5718 2535
rect 5752 2501 5759 2535
rect 5567 2461 5759 2501
rect 5567 2449 5646 2461
rect 5680 2449 5759 2461
rect 5567 1479 5574 2449
rect 5608 1479 5718 1491
rect 5752 1479 5759 2449
rect 5567 1467 5759 1479
rect 6063 4062 6255 4074
rect 6063 4028 6070 4062
rect 6104 4028 6142 4062
rect 6176 4028 6214 4062
rect 6248 4028 6255 4062
rect 6063 3988 6255 4028
rect 6063 3954 6070 3988
rect 6104 3954 6142 3988
rect 6176 3954 6214 3988
rect 6248 3954 6255 3988
rect 6063 3914 6255 3954
rect 6063 3880 6070 3914
rect 6104 3880 6142 3914
rect 6176 3880 6214 3914
rect 6248 3880 6255 3914
rect 6063 3840 6255 3880
rect 6063 3806 6070 3840
rect 6104 3806 6142 3840
rect 6176 3806 6214 3840
rect 6248 3806 6255 3840
rect 6063 3766 6255 3806
rect 6063 3732 6070 3766
rect 6104 3732 6142 3766
rect 6176 3732 6214 3766
rect 6248 3732 6255 3766
rect 6063 3692 6255 3732
rect 6063 3658 6070 3692
rect 6104 3658 6142 3692
rect 6176 3658 6214 3692
rect 6248 3658 6255 3692
rect 6063 3618 6255 3658
rect 6063 3584 6070 3618
rect 6104 3584 6142 3618
rect 6176 3584 6214 3618
rect 6248 3584 6255 3618
rect 6063 3544 6255 3584
rect 6063 3510 6070 3544
rect 6104 3510 6142 3544
rect 6176 3510 6214 3544
rect 6248 3510 6255 3544
rect 6063 3470 6255 3510
rect 6063 3436 6070 3470
rect 6104 3436 6142 3470
rect 6176 3436 6214 3470
rect 6248 3436 6255 3470
rect 6063 3396 6255 3436
rect 6063 3362 6070 3396
rect 6104 3362 6142 3396
rect 6176 3362 6214 3396
rect 6248 3362 6255 3396
rect 6063 3322 6255 3362
rect 6063 3288 6070 3322
rect 6104 3288 6142 3322
rect 6176 3288 6214 3322
rect 6248 3288 6255 3322
rect 6063 3248 6255 3288
rect 6063 3214 6070 3248
rect 6104 3214 6142 3248
rect 6176 3214 6214 3248
rect 6248 3214 6255 3248
rect 6063 3174 6255 3214
rect 6063 3140 6070 3174
rect 6104 3140 6142 3174
rect 6176 3140 6214 3174
rect 6248 3140 6255 3174
rect 6063 3100 6255 3140
rect 6063 3066 6070 3100
rect 6104 3066 6142 3100
rect 6176 3066 6214 3100
rect 6248 3066 6255 3100
rect 6063 3026 6255 3066
rect 6063 2992 6070 3026
rect 6104 2992 6142 3026
rect 6176 2992 6214 3026
rect 6248 2992 6255 3026
rect 6063 2952 6255 2992
rect 6063 2918 6070 2952
rect 6104 2918 6142 2952
rect 6176 2918 6214 2952
rect 6248 2918 6255 2952
rect 6063 2878 6255 2918
rect 6063 2844 6070 2878
rect 6104 2844 6142 2878
rect 6176 2844 6214 2878
rect 6248 2844 6255 2878
rect 6063 2804 6255 2844
rect 6063 2770 6070 2804
rect 6104 2770 6142 2804
rect 6176 2770 6214 2804
rect 6248 2770 6255 2804
rect 6063 2730 6255 2770
rect 6063 2696 6070 2730
rect 6104 2696 6142 2730
rect 6176 2696 6214 2730
rect 6248 2696 6255 2730
rect 6063 2656 6255 2696
rect 6063 2622 6070 2656
rect 6104 2622 6142 2656
rect 6176 2622 6214 2656
rect 6248 2622 6255 2656
rect 6063 2614 6255 2622
rect 6063 1538 6069 2614
rect 6249 1538 6255 2614
rect 6063 1525 6070 1538
rect 6104 1525 6142 1538
rect 6176 1525 6214 1538
rect 6248 1525 6255 1538
rect 6063 1473 6069 1525
rect 6121 1473 6133 1525
rect 6185 1473 6197 1525
rect 6249 1473 6255 1525
rect 6063 1467 6255 1473
rect 6559 4068 6751 4074
rect 6559 2992 6565 4068
rect 6745 2992 6751 4068
rect 6559 2979 6566 2992
rect 6744 2979 6751 2992
rect 6559 2927 6565 2979
rect 6745 2927 6751 2979
rect 6559 2574 6566 2927
rect 6744 2574 6751 2927
rect 6559 2535 6751 2574
rect 6559 2501 6566 2535
rect 6600 2501 6638 2535
rect 6672 2501 6710 2535
rect 6744 2501 6751 2535
rect 6559 2461 6751 2501
rect 6559 2449 6638 2461
rect 6672 2449 6751 2461
rect 6559 1479 6566 2449
rect 6600 1479 6710 1491
rect 6744 1479 6751 2449
rect 6559 1467 6751 1479
rect 7055 4062 7247 4074
rect 7055 4028 7062 4062
rect 7096 4028 7134 4062
rect 7168 4028 7206 4062
rect 7240 4028 7247 4062
rect 7055 3988 7247 4028
rect 7055 3954 7062 3988
rect 7096 3954 7134 3988
rect 7168 3954 7206 3988
rect 7240 3954 7247 3988
rect 7055 3914 7247 3954
rect 7055 3880 7062 3914
rect 7096 3880 7134 3914
rect 7168 3880 7206 3914
rect 7240 3880 7247 3914
rect 7055 3840 7247 3880
rect 7055 3806 7062 3840
rect 7096 3806 7134 3840
rect 7168 3806 7206 3840
rect 7240 3806 7247 3840
rect 7055 3766 7247 3806
rect 7055 3732 7062 3766
rect 7096 3732 7134 3766
rect 7168 3732 7206 3766
rect 7240 3732 7247 3766
rect 7055 3692 7247 3732
rect 7055 3658 7062 3692
rect 7096 3658 7134 3692
rect 7168 3658 7206 3692
rect 7240 3658 7247 3692
rect 7055 3618 7247 3658
rect 7055 3584 7062 3618
rect 7096 3584 7134 3618
rect 7168 3584 7206 3618
rect 7240 3584 7247 3618
rect 7055 3544 7247 3584
rect 7055 3510 7062 3544
rect 7096 3510 7134 3544
rect 7168 3510 7206 3544
rect 7240 3510 7247 3544
rect 7055 3470 7247 3510
rect 7055 3436 7062 3470
rect 7096 3436 7134 3470
rect 7168 3436 7206 3470
rect 7240 3436 7247 3470
rect 7055 3396 7247 3436
rect 7055 3362 7062 3396
rect 7096 3362 7134 3396
rect 7168 3362 7206 3396
rect 7240 3362 7247 3396
rect 7055 3322 7247 3362
rect 7055 3288 7062 3322
rect 7096 3288 7134 3322
rect 7168 3288 7206 3322
rect 7240 3288 7247 3322
rect 7055 3248 7247 3288
rect 7055 3214 7062 3248
rect 7096 3214 7134 3248
rect 7168 3214 7206 3248
rect 7240 3214 7247 3248
rect 7055 3174 7247 3214
rect 7055 3140 7062 3174
rect 7096 3140 7134 3174
rect 7168 3140 7206 3174
rect 7240 3140 7247 3174
rect 7055 3100 7247 3140
rect 7055 3066 7062 3100
rect 7096 3066 7134 3100
rect 7168 3066 7206 3100
rect 7240 3066 7247 3100
rect 7055 3026 7247 3066
rect 7055 2992 7062 3026
rect 7096 2992 7134 3026
rect 7168 2992 7206 3026
rect 7240 2992 7247 3026
rect 7055 2952 7247 2992
rect 7055 2918 7062 2952
rect 7096 2918 7134 2952
rect 7168 2918 7206 2952
rect 7240 2918 7247 2952
rect 7055 2878 7247 2918
rect 7055 2844 7062 2878
rect 7096 2844 7134 2878
rect 7168 2844 7206 2878
rect 7240 2844 7247 2878
rect 7055 2804 7247 2844
rect 7055 2770 7062 2804
rect 7096 2770 7134 2804
rect 7168 2770 7206 2804
rect 7240 2770 7247 2804
rect 7055 2730 7247 2770
rect 7055 2696 7062 2730
rect 7096 2696 7134 2730
rect 7168 2696 7206 2730
rect 7240 2696 7247 2730
rect 7055 2656 7247 2696
rect 7055 2622 7062 2656
rect 7096 2622 7134 2656
rect 7168 2622 7206 2656
rect 7240 2622 7247 2656
rect 7055 2614 7247 2622
rect 7055 1538 7061 2614
rect 7241 1538 7247 2614
rect 7055 1525 7062 1538
rect 7096 1525 7134 1538
rect 7168 1525 7206 1538
rect 7240 1525 7247 1538
rect 7055 1473 7061 1525
rect 7113 1473 7125 1525
rect 7177 1473 7189 1525
rect 7241 1473 7247 1525
rect 7055 1467 7247 1473
rect 7551 4068 7743 4074
rect 7551 2992 7557 4068
rect 7737 2992 7743 4068
rect 7551 2979 7558 2992
rect 7736 2979 7743 2992
rect 7551 2927 7557 2979
rect 7737 2927 7743 2979
rect 7551 2574 7558 2927
rect 7736 2574 7743 2927
rect 7551 2535 7743 2574
rect 7551 2501 7558 2535
rect 7592 2501 7630 2535
rect 7664 2501 7702 2535
rect 7736 2501 7743 2535
rect 7551 2461 7743 2501
rect 7551 2449 7630 2461
rect 7664 2449 7743 2461
rect 7551 1479 7558 2449
rect 7592 1479 7702 1491
rect 7736 1479 7743 2449
rect 7551 1467 7743 1479
rect 8047 4062 8239 4074
rect 8047 4028 8054 4062
rect 8088 4028 8126 4062
rect 8160 4028 8198 4062
rect 8232 4028 8239 4062
rect 8047 3988 8239 4028
rect 8047 3954 8054 3988
rect 8088 3954 8126 3988
rect 8160 3954 8198 3988
rect 8232 3954 8239 3988
rect 8047 3914 8239 3954
rect 8047 3880 8054 3914
rect 8088 3880 8126 3914
rect 8160 3880 8198 3914
rect 8232 3880 8239 3914
rect 8047 3840 8239 3880
rect 8047 3806 8054 3840
rect 8088 3806 8126 3840
rect 8160 3806 8198 3840
rect 8232 3806 8239 3840
rect 8047 3766 8239 3806
rect 8047 3732 8054 3766
rect 8088 3732 8126 3766
rect 8160 3732 8198 3766
rect 8232 3732 8239 3766
rect 8047 3692 8239 3732
rect 8047 3658 8054 3692
rect 8088 3658 8126 3692
rect 8160 3658 8198 3692
rect 8232 3658 8239 3692
rect 8047 3618 8239 3658
rect 8047 3584 8054 3618
rect 8088 3584 8126 3618
rect 8160 3584 8198 3618
rect 8232 3584 8239 3618
rect 8047 3544 8239 3584
rect 8047 3510 8054 3544
rect 8088 3510 8126 3544
rect 8160 3510 8198 3544
rect 8232 3510 8239 3544
rect 8047 3470 8239 3510
rect 8047 3436 8054 3470
rect 8088 3436 8126 3470
rect 8160 3436 8198 3470
rect 8232 3436 8239 3470
rect 8047 3396 8239 3436
rect 8047 3362 8054 3396
rect 8088 3362 8126 3396
rect 8160 3362 8198 3396
rect 8232 3362 8239 3396
rect 8047 3322 8239 3362
rect 8047 3288 8054 3322
rect 8088 3288 8126 3322
rect 8160 3288 8198 3322
rect 8232 3288 8239 3322
rect 8047 3248 8239 3288
rect 8047 3214 8054 3248
rect 8088 3214 8126 3248
rect 8160 3214 8198 3248
rect 8232 3214 8239 3248
rect 8047 3174 8239 3214
rect 8047 3140 8054 3174
rect 8088 3140 8126 3174
rect 8160 3140 8198 3174
rect 8232 3140 8239 3174
rect 8047 3100 8239 3140
rect 8047 3066 8054 3100
rect 8088 3066 8126 3100
rect 8160 3066 8198 3100
rect 8232 3066 8239 3100
rect 8047 3026 8239 3066
rect 8047 2992 8054 3026
rect 8088 2992 8126 3026
rect 8160 2992 8198 3026
rect 8232 2992 8239 3026
rect 8047 2952 8239 2992
rect 8047 2918 8054 2952
rect 8088 2918 8126 2952
rect 8160 2918 8198 2952
rect 8232 2918 8239 2952
rect 8047 2878 8239 2918
rect 8047 2844 8054 2878
rect 8088 2844 8126 2878
rect 8160 2844 8198 2878
rect 8232 2844 8239 2878
rect 8047 2804 8239 2844
rect 8047 2770 8054 2804
rect 8088 2770 8126 2804
rect 8160 2770 8198 2804
rect 8232 2770 8239 2804
rect 8047 2730 8239 2770
rect 8047 2696 8054 2730
rect 8088 2696 8126 2730
rect 8160 2696 8198 2730
rect 8232 2696 8239 2730
rect 8047 2656 8239 2696
rect 8047 2622 8054 2656
rect 8088 2622 8126 2656
rect 8160 2622 8198 2656
rect 8232 2622 8239 2656
rect 8047 2614 8239 2622
rect 8047 1538 8053 2614
rect 8233 1538 8239 2614
rect 8047 1525 8054 1538
rect 8088 1525 8126 1538
rect 8160 1525 8198 1538
rect 8232 1525 8239 1538
rect 8047 1473 8053 1525
rect 8105 1473 8117 1525
rect 8169 1473 8181 1525
rect 8233 1473 8239 1525
rect 8047 1467 8239 1473
rect 8543 4068 8735 4074
rect 8543 2992 8549 4068
rect 8729 2992 8735 4068
rect 8543 2979 8550 2992
rect 8728 2979 8735 2992
rect 8543 2927 8549 2979
rect 8729 2927 8735 2979
rect 8543 2574 8550 2927
rect 8728 2574 8735 2927
rect 8543 2535 8735 2574
rect 8543 2501 8550 2535
rect 8584 2501 8622 2535
rect 8656 2501 8694 2535
rect 8728 2501 8735 2535
rect 8543 2461 8735 2501
rect 8543 2449 8622 2461
rect 8656 2449 8735 2461
rect 8543 1479 8550 2449
rect 8584 1479 8694 1491
rect 8728 1479 8735 2449
rect 8543 1467 8735 1479
rect 9039 4062 9231 4074
rect 9039 4028 9046 4062
rect 9080 4028 9118 4062
rect 9152 4028 9190 4062
rect 9224 4028 9231 4062
rect 9039 3988 9231 4028
rect 9039 3954 9046 3988
rect 9080 3954 9118 3988
rect 9152 3954 9190 3988
rect 9224 3954 9231 3988
rect 9039 3914 9231 3954
rect 9039 3880 9046 3914
rect 9080 3880 9118 3914
rect 9152 3880 9190 3914
rect 9224 3880 9231 3914
rect 9039 3840 9231 3880
rect 9039 3806 9046 3840
rect 9080 3806 9118 3840
rect 9152 3806 9190 3840
rect 9224 3806 9231 3840
rect 9039 3766 9231 3806
rect 9039 3732 9046 3766
rect 9080 3732 9118 3766
rect 9152 3732 9190 3766
rect 9224 3732 9231 3766
rect 9039 3692 9231 3732
rect 9039 3658 9046 3692
rect 9080 3658 9118 3692
rect 9152 3658 9190 3692
rect 9224 3658 9231 3692
rect 9039 3618 9231 3658
rect 9039 3584 9046 3618
rect 9080 3584 9118 3618
rect 9152 3584 9190 3618
rect 9224 3584 9231 3618
rect 9039 3544 9231 3584
rect 9039 3510 9046 3544
rect 9080 3510 9118 3544
rect 9152 3510 9190 3544
rect 9224 3510 9231 3544
rect 9039 3470 9231 3510
rect 9039 3436 9046 3470
rect 9080 3436 9118 3470
rect 9152 3436 9190 3470
rect 9224 3436 9231 3470
rect 9039 3396 9231 3436
rect 9039 3362 9046 3396
rect 9080 3362 9118 3396
rect 9152 3362 9190 3396
rect 9224 3362 9231 3396
rect 9039 3322 9231 3362
rect 9039 3288 9046 3322
rect 9080 3288 9118 3322
rect 9152 3288 9190 3322
rect 9224 3288 9231 3322
rect 9039 3248 9231 3288
rect 9039 3214 9046 3248
rect 9080 3214 9118 3248
rect 9152 3214 9190 3248
rect 9224 3214 9231 3248
rect 9039 3174 9231 3214
rect 9039 3140 9046 3174
rect 9080 3140 9118 3174
rect 9152 3140 9190 3174
rect 9224 3140 9231 3174
rect 9039 3100 9231 3140
rect 9039 3066 9046 3100
rect 9080 3066 9118 3100
rect 9152 3066 9190 3100
rect 9224 3066 9231 3100
rect 9039 3026 9231 3066
rect 9039 2992 9046 3026
rect 9080 2992 9118 3026
rect 9152 2992 9190 3026
rect 9224 2992 9231 3026
rect 9039 2952 9231 2992
rect 9039 2918 9046 2952
rect 9080 2918 9118 2952
rect 9152 2918 9190 2952
rect 9224 2918 9231 2952
rect 9039 2878 9231 2918
rect 9039 2844 9046 2878
rect 9080 2844 9118 2878
rect 9152 2844 9190 2878
rect 9224 2844 9231 2878
rect 9039 2804 9231 2844
rect 9039 2770 9046 2804
rect 9080 2770 9118 2804
rect 9152 2770 9190 2804
rect 9224 2770 9231 2804
rect 9039 2730 9231 2770
rect 9039 2696 9046 2730
rect 9080 2696 9118 2730
rect 9152 2696 9190 2730
rect 9224 2696 9231 2730
rect 9039 2656 9231 2696
rect 9039 2622 9046 2656
rect 9080 2622 9118 2656
rect 9152 2622 9190 2656
rect 9224 2622 9231 2656
rect 9039 2614 9231 2622
rect 9039 1538 9045 2614
rect 9225 1538 9231 2614
rect 9039 1525 9046 1538
rect 9080 1525 9118 1538
rect 9152 1525 9190 1538
rect 9224 1525 9231 1538
rect 9039 1473 9045 1525
rect 9097 1473 9109 1525
rect 9161 1473 9173 1525
rect 9225 1473 9231 1525
rect 9039 1467 9231 1473
rect 9535 4068 9727 4074
rect 9535 2992 9541 4068
rect 9721 2992 9727 4068
rect 9535 2979 9542 2992
rect 9720 2979 9727 2992
rect 9535 2927 9541 2979
rect 9721 2927 9727 2979
rect 9535 2574 9542 2927
rect 9720 2574 9727 2927
rect 9535 2535 9727 2574
rect 9535 2501 9542 2535
rect 9576 2501 9614 2535
rect 9648 2501 9686 2535
rect 9720 2501 9727 2535
rect 9535 2461 9727 2501
rect 9535 2449 9614 2461
rect 9648 2449 9727 2461
rect 9535 1479 9542 2449
rect 9576 1479 9686 1491
rect 9720 1479 9727 2449
rect 9535 1467 9727 1479
rect 10031 4062 10223 4074
rect 10031 4028 10038 4062
rect 10072 4028 10110 4062
rect 10144 4028 10182 4062
rect 10216 4028 10223 4062
rect 10031 3988 10223 4028
rect 10031 3954 10038 3988
rect 10072 3954 10110 3988
rect 10144 3954 10182 3988
rect 10216 3954 10223 3988
rect 10031 3914 10223 3954
rect 10031 3880 10038 3914
rect 10072 3880 10110 3914
rect 10144 3880 10182 3914
rect 10216 3880 10223 3914
rect 10031 3840 10223 3880
rect 10031 3806 10038 3840
rect 10072 3806 10110 3840
rect 10144 3806 10182 3840
rect 10216 3806 10223 3840
rect 10031 3766 10223 3806
rect 10031 3732 10038 3766
rect 10072 3732 10110 3766
rect 10144 3732 10182 3766
rect 10216 3732 10223 3766
rect 10031 3692 10223 3732
rect 10031 3658 10038 3692
rect 10072 3658 10110 3692
rect 10144 3658 10182 3692
rect 10216 3658 10223 3692
rect 10031 3618 10223 3658
rect 10031 3584 10038 3618
rect 10072 3584 10110 3618
rect 10144 3584 10182 3618
rect 10216 3584 10223 3618
rect 10031 3544 10223 3584
rect 10031 3510 10038 3544
rect 10072 3510 10110 3544
rect 10144 3510 10182 3544
rect 10216 3510 10223 3544
rect 10031 3470 10223 3510
rect 10031 3436 10038 3470
rect 10072 3436 10110 3470
rect 10144 3436 10182 3470
rect 10216 3436 10223 3470
rect 10031 3396 10223 3436
rect 10031 3362 10038 3396
rect 10072 3362 10110 3396
rect 10144 3362 10182 3396
rect 10216 3362 10223 3396
rect 10031 3322 10223 3362
rect 10031 3288 10038 3322
rect 10072 3288 10110 3322
rect 10144 3288 10182 3322
rect 10216 3288 10223 3322
rect 10031 3248 10223 3288
rect 10031 3214 10038 3248
rect 10072 3214 10110 3248
rect 10144 3214 10182 3248
rect 10216 3214 10223 3248
rect 10031 3174 10223 3214
rect 10031 3140 10038 3174
rect 10072 3140 10110 3174
rect 10144 3140 10182 3174
rect 10216 3140 10223 3174
rect 10031 3100 10223 3140
rect 10031 3066 10038 3100
rect 10072 3066 10110 3100
rect 10144 3066 10182 3100
rect 10216 3066 10223 3100
rect 10031 3026 10223 3066
rect 10031 2992 10038 3026
rect 10072 2992 10110 3026
rect 10144 2992 10182 3026
rect 10216 2992 10223 3026
rect 10031 2952 10223 2992
rect 10031 2918 10038 2952
rect 10072 2918 10110 2952
rect 10144 2918 10182 2952
rect 10216 2918 10223 2952
rect 10031 2878 10223 2918
rect 10031 2844 10038 2878
rect 10072 2844 10110 2878
rect 10144 2844 10182 2878
rect 10216 2844 10223 2878
rect 10031 2804 10223 2844
rect 10031 2770 10038 2804
rect 10072 2770 10110 2804
rect 10144 2770 10182 2804
rect 10216 2770 10223 2804
rect 10031 2730 10223 2770
rect 10031 2696 10038 2730
rect 10072 2696 10110 2730
rect 10144 2696 10182 2730
rect 10216 2696 10223 2730
rect 10031 2656 10223 2696
rect 10031 2622 10038 2656
rect 10072 2622 10110 2656
rect 10144 2622 10182 2656
rect 10216 2622 10223 2656
rect 10031 2614 10223 2622
rect 10031 1538 10037 2614
rect 10217 1538 10223 2614
rect 10031 1525 10038 1538
rect 10072 1525 10110 1538
rect 10144 1525 10182 1538
rect 10216 1525 10223 1538
rect 10031 1473 10037 1525
rect 10089 1473 10101 1525
rect 10153 1473 10165 1525
rect 10217 1473 10223 1525
rect 10031 1467 10223 1473
rect 10527 4068 10719 4074
rect 10527 2992 10533 4068
rect 10713 2992 10719 4068
rect 10527 2979 10719 2992
rect 10527 2927 10533 2979
rect 10585 2927 10597 2979
rect 10649 2927 10661 2979
rect 10713 2927 10719 2979
rect 10527 2920 10534 2927
rect 10568 2920 10606 2927
rect 10640 2920 10678 2927
rect 10712 2920 10719 2927
rect 10527 2871 10719 2920
rect 10527 2837 10534 2871
rect 10568 2837 10606 2871
rect 10640 2837 10678 2871
rect 10712 2837 10719 2871
rect 10527 2787 10719 2837
rect 10527 2753 10534 2787
rect 10568 2753 10606 2787
rect 10640 2753 10678 2787
rect 10712 2753 10719 2787
rect 10527 2703 10719 2753
rect 10527 2669 10534 2703
rect 10568 2669 10606 2703
rect 10640 2669 10678 2703
rect 10712 2669 10719 2703
rect 10527 2619 10719 2669
rect 10527 2585 10534 2619
rect 10568 2585 10606 2619
rect 10640 2585 10678 2619
rect 10712 2585 10719 2619
rect 10527 2535 10719 2585
rect 10527 2501 10534 2535
rect 10568 2501 10606 2535
rect 10640 2501 10678 2535
rect 10712 2501 10719 2535
rect 10527 2461 10719 2501
rect 10527 2449 10606 2461
rect 10640 2449 10719 2461
rect 10527 1479 10534 2449
rect 10568 1479 10678 1491
rect 10712 1479 10719 2449
rect 10527 1467 10719 1479
rect 11023 4062 11215 4074
rect 11023 4028 11030 4062
rect 11064 4028 11102 4062
rect 11136 4028 11174 4062
rect 11208 4028 11215 4062
rect 11023 3988 11215 4028
rect 11023 3954 11030 3988
rect 11064 3954 11102 3988
rect 11136 3954 11174 3988
rect 11208 3954 11215 3988
rect 11023 3914 11215 3954
rect 11023 3880 11030 3914
rect 11064 3880 11102 3914
rect 11136 3880 11174 3914
rect 11208 3880 11215 3914
rect 11023 3840 11215 3880
rect 11023 3806 11030 3840
rect 11064 3806 11102 3840
rect 11136 3806 11174 3840
rect 11208 3806 11215 3840
rect 11023 3766 11215 3806
rect 11023 3732 11030 3766
rect 11064 3732 11102 3766
rect 11136 3732 11174 3766
rect 11208 3732 11215 3766
rect 11023 3692 11215 3732
rect 11023 3658 11030 3692
rect 11064 3658 11102 3692
rect 11136 3658 11174 3692
rect 11208 3658 11215 3692
rect 11023 3618 11215 3658
rect 11023 3584 11030 3618
rect 11064 3584 11102 3618
rect 11136 3584 11174 3618
rect 11208 3584 11215 3618
rect 11023 3544 11215 3584
rect 11023 3510 11030 3544
rect 11064 3510 11102 3544
rect 11136 3510 11174 3544
rect 11208 3510 11215 3544
rect 11023 3470 11215 3510
rect 11023 3436 11030 3470
rect 11064 3436 11102 3470
rect 11136 3436 11174 3470
rect 11208 3436 11215 3470
rect 11023 3396 11215 3436
rect 11023 3362 11030 3396
rect 11064 3362 11102 3396
rect 11136 3362 11174 3396
rect 11208 3362 11215 3396
rect 11023 3322 11215 3362
rect 11023 3288 11030 3322
rect 11064 3288 11102 3322
rect 11136 3288 11174 3322
rect 11208 3288 11215 3322
rect 11023 3248 11215 3288
rect 11023 3214 11030 3248
rect 11064 3214 11102 3248
rect 11136 3214 11174 3248
rect 11208 3214 11215 3248
rect 11023 3174 11215 3214
rect 11023 3140 11030 3174
rect 11064 3140 11102 3174
rect 11136 3140 11174 3174
rect 11208 3140 11215 3174
rect 11023 3100 11215 3140
rect 11023 3066 11030 3100
rect 11064 3066 11102 3100
rect 11136 3066 11174 3100
rect 11208 3066 11215 3100
rect 11023 3026 11215 3066
rect 11023 2992 11030 3026
rect 11064 2992 11102 3026
rect 11136 2992 11174 3026
rect 11208 2992 11215 3026
rect 11023 2952 11215 2992
rect 11023 2918 11030 2952
rect 11064 2918 11102 2952
rect 11136 2918 11174 2952
rect 11208 2918 11215 2952
rect 11023 2878 11215 2918
rect 11023 2844 11030 2878
rect 11064 2844 11102 2878
rect 11136 2844 11174 2878
rect 11208 2844 11215 2878
rect 11023 2804 11215 2844
rect 11023 2770 11030 2804
rect 11064 2770 11102 2804
rect 11136 2770 11174 2804
rect 11208 2770 11215 2804
rect 11023 2730 11215 2770
rect 11023 2696 11030 2730
rect 11064 2696 11102 2730
rect 11136 2696 11174 2730
rect 11208 2696 11215 2730
rect 11023 2656 11215 2696
rect 11023 2622 11030 2656
rect 11064 2622 11102 2656
rect 11136 2622 11174 2656
rect 11208 2622 11215 2656
rect 11023 2614 11215 2622
rect 11023 1538 11029 2614
rect 11209 1538 11215 2614
rect 11023 1525 11030 1538
rect 11064 1525 11102 1538
rect 11136 1525 11174 1538
rect 11208 1525 11215 1538
rect 11023 1473 11029 1525
rect 11081 1473 11093 1525
rect 11145 1473 11157 1525
rect 11209 1473 11215 1525
rect 11023 1467 11215 1473
rect 11519 4068 11711 4074
rect 11519 2992 11525 4068
rect 11705 2992 11711 4068
rect 11519 2979 11711 2992
rect 11519 2927 11525 2979
rect 11577 2927 11589 2979
rect 11641 2927 11653 2979
rect 11705 2927 11711 2979
rect 11519 2920 11526 2927
rect 11560 2920 11598 2927
rect 11632 2920 11670 2927
rect 11704 2920 11711 2927
rect 11519 2871 11711 2920
rect 11519 2837 11526 2871
rect 11560 2837 11598 2871
rect 11632 2837 11670 2871
rect 11704 2837 11711 2871
rect 11519 2787 11711 2837
rect 11519 2753 11526 2787
rect 11560 2753 11598 2787
rect 11632 2753 11670 2787
rect 11704 2753 11711 2787
rect 11519 2703 11711 2753
rect 11519 2669 11526 2703
rect 11560 2669 11598 2703
rect 11632 2669 11670 2703
rect 11704 2669 11711 2703
rect 11519 2619 11711 2669
rect 11519 2585 11526 2619
rect 11560 2585 11598 2619
rect 11632 2585 11670 2619
rect 11704 2585 11711 2619
rect 11519 2535 11711 2585
rect 11519 2501 11526 2535
rect 11560 2501 11598 2535
rect 11632 2501 11670 2535
rect 11704 2501 11711 2535
rect 11519 2461 11711 2501
rect 11519 2449 11598 2461
rect 11632 2449 11711 2461
rect 11519 1479 11526 2449
rect 11560 1479 11670 1491
rect 11704 1479 11711 2449
rect 11519 1467 11711 1479
rect 12015 4062 12207 4074
rect 12015 4028 12022 4062
rect 12056 4028 12094 4062
rect 12128 4028 12166 4062
rect 12200 4028 12207 4062
rect 12015 3988 12207 4028
rect 12015 3954 12022 3988
rect 12056 3954 12094 3988
rect 12128 3954 12166 3988
rect 12200 3954 12207 3988
rect 12015 3914 12207 3954
rect 12015 3880 12022 3914
rect 12056 3880 12094 3914
rect 12128 3880 12166 3914
rect 12200 3880 12207 3914
rect 12015 3840 12207 3880
rect 12015 3806 12022 3840
rect 12056 3806 12094 3840
rect 12128 3806 12166 3840
rect 12200 3806 12207 3840
rect 12015 3766 12207 3806
rect 12015 3732 12022 3766
rect 12056 3732 12094 3766
rect 12128 3732 12166 3766
rect 12200 3732 12207 3766
rect 12015 3692 12207 3732
rect 12015 3658 12022 3692
rect 12056 3658 12094 3692
rect 12128 3658 12166 3692
rect 12200 3658 12207 3692
rect 12015 3618 12207 3658
rect 12015 3584 12022 3618
rect 12056 3584 12094 3618
rect 12128 3584 12166 3618
rect 12200 3584 12207 3618
rect 12015 3544 12207 3584
rect 12015 3510 12022 3544
rect 12056 3510 12094 3544
rect 12128 3510 12166 3544
rect 12200 3510 12207 3544
rect 12015 3470 12207 3510
rect 12015 3436 12022 3470
rect 12056 3436 12094 3470
rect 12128 3436 12166 3470
rect 12200 3436 12207 3470
rect 12015 3396 12207 3436
rect 12015 3362 12022 3396
rect 12056 3362 12094 3396
rect 12128 3362 12166 3396
rect 12200 3362 12207 3396
rect 12015 3322 12207 3362
rect 12015 3288 12022 3322
rect 12056 3288 12094 3322
rect 12128 3288 12166 3322
rect 12200 3288 12207 3322
rect 12015 3248 12207 3288
rect 12015 3214 12022 3248
rect 12056 3214 12094 3248
rect 12128 3214 12166 3248
rect 12200 3214 12207 3248
rect 12015 3174 12207 3214
rect 12015 3140 12022 3174
rect 12056 3140 12094 3174
rect 12128 3140 12166 3174
rect 12200 3140 12207 3174
rect 12015 3100 12207 3140
rect 12015 3066 12022 3100
rect 12056 3066 12094 3100
rect 12128 3066 12166 3100
rect 12200 3066 12207 3100
rect 12015 3026 12207 3066
rect 12015 2992 12022 3026
rect 12056 2992 12094 3026
rect 12128 2992 12166 3026
rect 12200 2992 12207 3026
rect 12015 2952 12207 2992
rect 12015 2918 12022 2952
rect 12056 2918 12094 2952
rect 12128 2918 12166 2952
rect 12200 2918 12207 2952
rect 12015 2878 12207 2918
rect 12015 2844 12022 2878
rect 12056 2844 12094 2878
rect 12128 2844 12166 2878
rect 12200 2844 12207 2878
rect 12015 2804 12207 2844
rect 12015 2770 12022 2804
rect 12056 2770 12094 2804
rect 12128 2770 12166 2804
rect 12200 2770 12207 2804
rect 12015 2730 12207 2770
rect 12015 2696 12022 2730
rect 12056 2696 12094 2730
rect 12128 2696 12166 2730
rect 12200 2696 12207 2730
rect 12015 2656 12207 2696
rect 12015 2622 12022 2656
rect 12056 2622 12094 2656
rect 12128 2622 12166 2656
rect 12200 2622 12207 2656
rect 12015 2614 12207 2622
rect 12015 1538 12021 2614
rect 12201 1538 12207 2614
rect 12015 1525 12022 1538
rect 12056 1525 12094 1538
rect 12128 1525 12166 1538
rect 12200 1525 12207 1538
rect 12015 1473 12021 1525
rect 12073 1473 12085 1525
rect 12137 1473 12149 1525
rect 12201 1473 12207 1525
rect 12015 1467 12207 1473
rect 12511 4068 12703 4074
rect 12511 2992 12517 4068
rect 12697 2992 12703 4068
rect 12511 2979 12703 2992
rect 12511 2927 12517 2979
rect 12569 2927 12581 2979
rect 12633 2927 12645 2979
rect 12697 2927 12703 2979
rect 12511 2921 12518 2927
rect 12552 2921 12590 2927
rect 12624 2921 12662 2927
rect 12696 2921 12703 2927
rect 12511 2871 12703 2921
rect 12511 2837 12518 2871
rect 12552 2837 12590 2871
rect 12624 2837 12662 2871
rect 12696 2837 12703 2871
rect 12511 2787 12703 2837
rect 12511 2753 12518 2787
rect 12552 2753 12590 2787
rect 12624 2753 12662 2787
rect 12696 2753 12703 2787
rect 12511 2703 12703 2753
rect 12511 2669 12518 2703
rect 12552 2669 12590 2703
rect 12624 2669 12662 2703
rect 12696 2669 12703 2703
rect 12511 2619 12703 2669
rect 12511 2585 12518 2619
rect 12552 2585 12590 2619
rect 12624 2585 12662 2619
rect 12696 2585 12703 2619
rect 12511 2535 12703 2585
rect 12511 2501 12518 2535
rect 12552 2501 12590 2535
rect 12624 2501 12662 2535
rect 12696 2501 12703 2535
rect 12511 2461 12703 2501
rect 12511 2449 12590 2461
rect 12624 2449 12703 2461
rect 12511 1479 12518 2449
rect 12552 1479 12662 1491
rect 12696 1479 12703 2449
rect 12511 1467 12703 1479
rect 13007 4062 13199 4074
rect 13007 4028 13014 4062
rect 13048 4028 13086 4062
rect 13120 4028 13158 4062
rect 13192 4028 13199 4062
rect 13007 3988 13199 4028
rect 13007 3954 13014 3988
rect 13048 3954 13086 3988
rect 13120 3954 13158 3988
rect 13192 3954 13199 3988
rect 13007 3914 13199 3954
rect 13007 3880 13014 3914
rect 13048 3880 13086 3914
rect 13120 3880 13158 3914
rect 13192 3880 13199 3914
rect 13007 3840 13199 3880
rect 13007 3806 13014 3840
rect 13048 3806 13086 3840
rect 13120 3806 13158 3840
rect 13192 3806 13199 3840
rect 13007 3766 13199 3806
rect 13007 3732 13014 3766
rect 13048 3732 13086 3766
rect 13120 3732 13158 3766
rect 13192 3732 13199 3766
rect 13007 3692 13199 3732
rect 13007 3658 13014 3692
rect 13048 3658 13086 3692
rect 13120 3658 13158 3692
rect 13192 3658 13199 3692
rect 13007 3618 13199 3658
rect 13007 3584 13014 3618
rect 13048 3584 13086 3618
rect 13120 3584 13158 3618
rect 13192 3584 13199 3618
rect 13007 3544 13199 3584
rect 13007 3510 13014 3544
rect 13048 3510 13086 3544
rect 13120 3510 13158 3544
rect 13192 3510 13199 3544
rect 13007 3470 13199 3510
rect 13007 3436 13014 3470
rect 13048 3436 13086 3470
rect 13120 3436 13158 3470
rect 13192 3436 13199 3470
rect 13007 3396 13199 3436
rect 13007 3362 13014 3396
rect 13048 3362 13086 3396
rect 13120 3362 13158 3396
rect 13192 3362 13199 3396
rect 13007 3322 13199 3362
rect 13007 3288 13014 3322
rect 13048 3288 13086 3322
rect 13120 3288 13158 3322
rect 13192 3288 13199 3322
rect 13007 3248 13199 3288
rect 13007 3214 13014 3248
rect 13048 3214 13086 3248
rect 13120 3214 13158 3248
rect 13192 3214 13199 3248
rect 13007 3174 13199 3214
rect 13007 3140 13014 3174
rect 13048 3140 13086 3174
rect 13120 3140 13158 3174
rect 13192 3140 13199 3174
rect 13007 3100 13199 3140
rect 13007 3066 13014 3100
rect 13048 3066 13086 3100
rect 13120 3066 13158 3100
rect 13192 3066 13199 3100
rect 13007 3026 13199 3066
rect 13007 2992 13014 3026
rect 13048 2992 13086 3026
rect 13120 2992 13158 3026
rect 13192 2992 13199 3026
rect 13007 2952 13199 2992
rect 13007 2918 13014 2952
rect 13048 2918 13086 2952
rect 13120 2918 13158 2952
rect 13192 2918 13199 2952
rect 13007 2878 13199 2918
rect 13007 2844 13014 2878
rect 13048 2844 13086 2878
rect 13120 2844 13158 2878
rect 13192 2844 13199 2878
rect 13007 2804 13199 2844
rect 13007 2770 13014 2804
rect 13048 2770 13086 2804
rect 13120 2770 13158 2804
rect 13192 2770 13199 2804
rect 13007 2730 13199 2770
rect 13007 2696 13014 2730
rect 13048 2696 13086 2730
rect 13120 2696 13158 2730
rect 13192 2696 13199 2730
rect 13007 2656 13199 2696
rect 13007 2622 13014 2656
rect 13048 2622 13086 2656
rect 13120 2622 13158 2656
rect 13192 2622 13199 2656
rect 13007 2614 13199 2622
rect 13007 1538 13013 2614
rect 13193 1538 13199 2614
rect 13007 1525 13014 1538
rect 13048 1525 13086 1538
rect 13120 1525 13158 1538
rect 13192 1525 13199 1538
rect 13007 1473 13013 1525
rect 13065 1473 13077 1525
rect 13129 1473 13141 1525
rect 13193 1473 13199 1525
rect 13007 1467 13199 1473
rect 13503 4068 13695 4074
rect 13503 2992 13509 4068
rect 13689 2992 13695 4068
rect 13503 2979 13510 2992
rect 13688 2979 13695 2992
rect 13503 2927 13509 2979
rect 13689 2927 13695 2979
rect 13503 2574 13510 2927
rect 13688 2574 13695 2927
rect 13503 2535 13695 2574
rect 13503 2501 13510 2535
rect 13544 2501 13582 2535
rect 13616 2501 13654 2535
rect 13688 2501 13695 2535
rect 13503 2461 13695 2501
rect 13503 2449 13582 2461
rect 13616 2449 13695 2461
rect 13503 1479 13510 2449
rect 13544 1479 13654 1491
rect 13688 1479 13695 2449
rect 13503 1467 13695 1479
rect 14036 4062 14226 4074
rect 14036 4028 14042 4062
rect 14076 4028 14226 4062
rect 14036 3990 14226 4028
rect 14036 3956 14042 3990
rect 14076 3956 14226 3990
rect 14036 3918 14226 3956
rect 14036 3884 14042 3918
rect 14076 3884 14226 3918
rect 14036 3846 14226 3884
rect 14036 3812 14042 3846
rect 14076 3812 14226 3846
rect 14036 3774 14226 3812
rect 14036 3740 14042 3774
rect 14076 3740 14226 3774
rect 14036 3702 14226 3740
rect 14036 3668 14042 3702
rect 14076 3668 14226 3702
rect 14036 3630 14226 3668
rect 14036 3596 14042 3630
rect 14076 3596 14226 3630
rect 14036 3558 14226 3596
rect 14036 3524 14042 3558
rect 14076 3524 14226 3558
rect 14036 3486 14226 3524
rect 14036 3452 14042 3486
rect 14076 3452 14226 3486
rect 14036 3414 14226 3452
rect 14036 3380 14042 3414
rect 14076 3380 14226 3414
rect 14036 3342 14226 3380
rect 14036 3308 14042 3342
rect 14076 3308 14226 3342
rect 14036 3270 14226 3308
rect 14036 3236 14042 3270
rect 14076 3236 14226 3270
rect 14036 3198 14226 3236
rect 14036 3164 14042 3198
rect 14076 3164 14226 3198
rect 14036 3126 14226 3164
rect 14036 3092 14042 3126
rect 14076 3092 14226 3126
rect 14036 3054 14226 3092
rect 14036 3020 14042 3054
rect 14076 3020 14226 3054
rect 14036 2982 14226 3020
rect 14036 2948 14042 2982
rect 14076 2948 14226 2982
rect 14036 2910 14226 2948
rect 14036 2876 14042 2910
rect 14076 2876 14226 2910
rect 14036 2838 14226 2876
rect 14036 2804 14042 2838
rect 14076 2804 14226 2838
rect 14036 2766 14226 2804
rect 14036 2732 14042 2766
rect 14076 2732 14226 2766
rect 14036 2693 14226 2732
rect 14036 2659 14042 2693
rect 14076 2659 14226 2693
rect 14036 2620 14226 2659
rect 14036 2614 14042 2620
rect 14076 2614 14226 2620
rect 14036 2562 14037 2614
rect 14089 2562 14105 2614
rect 14157 2562 14173 2614
rect 14225 2562 14226 2614
rect 14036 2550 14226 2562
rect 14036 2498 14037 2550
rect 14089 2498 14105 2550
rect 14157 2498 14173 2550
rect 14225 2498 14226 2550
rect 14036 2486 14226 2498
rect 14036 2434 14037 2486
rect 14089 2434 14105 2486
rect 14157 2434 14173 2486
rect 14225 2434 14226 2486
rect 14036 2422 14226 2434
rect 14036 2370 14037 2422
rect 14089 2370 14105 2422
rect 14157 2370 14173 2422
rect 14225 2370 14226 2422
rect 14036 2367 14042 2370
rect 14076 2367 14226 2370
rect 14036 2358 14226 2367
rect 14036 2306 14037 2358
rect 14089 2306 14105 2358
rect 14157 2306 14173 2358
rect 14225 2306 14226 2358
rect 14036 2294 14042 2306
rect 14076 2294 14226 2306
rect 14036 2242 14037 2294
rect 14089 2242 14105 2294
rect 14157 2242 14173 2294
rect 14225 2242 14226 2294
rect 14036 2230 14042 2242
rect 14076 2230 14226 2242
rect 14036 2178 14037 2230
rect 14089 2178 14105 2230
rect 14157 2178 14173 2230
rect 14225 2178 14226 2230
rect 14036 2166 14042 2178
rect 14076 2166 14226 2178
rect 14036 2114 14037 2166
rect 14089 2114 14105 2166
rect 14157 2114 14173 2166
rect 14225 2114 14226 2166
rect 14036 2109 14226 2114
rect 14036 2102 14042 2109
rect 14076 2102 14226 2109
rect 14036 2050 14037 2102
rect 14089 2050 14105 2102
rect 14157 2050 14173 2102
rect 14225 2050 14226 2102
rect 14036 2038 14226 2050
rect 14036 1986 14037 2038
rect 14089 1986 14105 2038
rect 14157 1986 14173 2038
rect 14225 1986 14226 2038
rect 14036 1974 14226 1986
rect 14036 1922 14037 1974
rect 14089 1922 14105 1974
rect 14157 1922 14173 1974
rect 14225 1922 14226 1974
rect 14036 1910 14226 1922
rect 14036 1858 14037 1910
rect 14089 1858 14105 1910
rect 14157 1858 14173 1910
rect 14225 1858 14226 1910
rect 14036 1856 14042 1858
rect 14076 1856 14226 1858
rect 14036 1846 14226 1856
rect 14036 1794 14037 1846
rect 14089 1794 14105 1846
rect 14157 1794 14173 1846
rect 14225 1794 14226 1846
rect 14036 1783 14042 1794
rect 14076 1783 14226 1794
rect 14036 1782 14226 1783
rect 14036 1730 14037 1782
rect 14089 1730 14105 1782
rect 14157 1730 14173 1782
rect 14225 1730 14226 1782
rect 14036 1718 14042 1730
rect 14076 1718 14226 1730
rect 14036 1666 14037 1718
rect 14089 1666 14105 1718
rect 14157 1666 14173 1718
rect 14225 1666 14226 1718
rect 14036 1654 14042 1666
rect 14076 1654 14226 1666
rect 14036 1602 14037 1654
rect 14089 1602 14105 1654
rect 14157 1602 14173 1654
rect 14225 1602 14226 1654
rect 14036 1598 14226 1602
rect 14036 1590 14042 1598
rect 14076 1590 14226 1598
rect 14036 1538 14037 1590
rect 14089 1538 14105 1590
rect 14157 1538 14173 1590
rect 14225 1538 14226 1590
rect 14036 1525 14226 1538
rect 14036 1473 14037 1525
rect 14089 1473 14105 1525
rect 14157 1473 14173 1525
rect 14225 1473 14226 1525
rect 14036 1467 14226 1473
rect 14400 4068 14510 4083
rect 14544 4068 14582 4086
rect 14616 4068 14628 4086
rect 14452 4044 14488 4068
rect 14544 4052 14576 4068
rect 14465 4016 14488 4044
rect 14540 4016 14576 4052
rect 14400 4010 14431 4016
rect 14465 4013 14628 4016
rect 14465 4010 14510 4013
rect 14400 4004 14510 4010
rect 14544 4004 14582 4013
rect 14616 4004 14628 4013
rect 14452 3971 14488 4004
rect 14544 3979 14576 4004
rect 14465 3952 14488 3971
rect 14540 3952 14576 3979
rect 14400 3940 14431 3952
rect 14465 3940 14628 3952
rect 14465 3937 14488 3940
rect 14452 3898 14488 3937
rect 14544 3906 14576 3940
rect 14465 3888 14488 3898
rect 14540 3888 14576 3906
rect 14400 3876 14431 3888
rect 14465 3876 14628 3888
rect 14465 3864 14488 3876
rect 14540 3867 14576 3876
rect 14452 3825 14488 3864
rect 14544 3833 14576 3867
rect 14465 3824 14488 3825
rect 14540 3824 14576 3833
rect 14400 3812 14431 3824
rect 14465 3812 14628 3824
rect 14465 3791 14488 3812
rect 14540 3794 14576 3812
rect 14452 3760 14488 3791
rect 14544 3760 14576 3794
rect 14400 3752 14628 3760
rect 14400 3748 14431 3752
rect 14465 3748 14628 3752
rect 14465 3718 14488 3748
rect 14540 3721 14576 3748
rect 14452 3696 14488 3718
rect 14544 3696 14576 3721
rect 14400 3687 14510 3696
rect 14544 3687 14582 3696
rect 14616 3687 14628 3696
rect 14400 3684 14628 3687
rect 14452 3679 14488 3684
rect 14465 3645 14488 3679
rect 14540 3648 14576 3684
rect 14452 3632 14488 3645
rect 14544 3632 14576 3648
rect 14400 3620 14510 3632
rect 14544 3620 14582 3632
rect 14616 3620 14628 3632
rect 14452 3606 14488 3620
rect 14544 3614 14576 3620
rect 14465 3572 14488 3606
rect 14540 3575 14576 3614
rect 14452 3568 14488 3572
rect 14544 3568 14576 3575
rect 14400 3556 14510 3568
rect 14544 3556 14582 3568
rect 14616 3556 14628 3568
rect 14452 3533 14488 3556
rect 14544 3541 14576 3556
rect 14465 3504 14488 3533
rect 14540 3504 14576 3541
rect 14400 3499 14431 3504
rect 14465 3502 14628 3504
rect 14465 3499 14510 3502
rect 14400 3492 14510 3499
rect 14544 3492 14582 3502
rect 14616 3492 14628 3502
rect 14452 3460 14488 3492
rect 14544 3468 14576 3492
rect 14465 3440 14488 3460
rect 14540 3440 14576 3468
rect 14400 3428 14431 3440
rect 14465 3429 14628 3440
rect 14465 3428 14510 3429
rect 14544 3428 14582 3429
rect 14616 3428 14628 3429
rect 14465 3426 14488 3428
rect 14452 3387 14488 3426
rect 14544 3395 14576 3428
rect 14465 3376 14488 3387
rect 14540 3376 14576 3395
rect 14400 3364 14431 3376
rect 14465 3364 14628 3376
rect 14465 3353 14488 3364
rect 14540 3356 14576 3364
rect 14452 3314 14488 3353
rect 14544 3322 14576 3356
rect 14465 3312 14488 3314
rect 14540 3312 14576 3322
rect 14400 3300 14431 3312
rect 14465 3300 14628 3312
rect 14465 3280 14488 3300
rect 14540 3283 14576 3300
rect 14452 3248 14488 3280
rect 14544 3249 14576 3283
rect 14540 3248 14576 3249
rect 14400 3241 14628 3248
rect 14400 3236 14431 3241
rect 14465 3236 14628 3241
rect 14465 3207 14488 3236
rect 14540 3210 14576 3236
rect 14452 3184 14488 3207
rect 14544 3184 14576 3210
rect 14400 3176 14510 3184
rect 14544 3176 14582 3184
rect 14616 3176 14628 3184
rect 14400 3172 14628 3176
rect 14452 3168 14488 3172
rect 14465 3134 14488 3168
rect 14540 3137 14576 3172
rect 14452 3120 14488 3134
rect 14544 3120 14576 3137
rect 14400 3108 14510 3120
rect 14544 3108 14582 3120
rect 14616 3108 14628 3120
rect 14452 3095 14488 3108
rect 14544 3103 14576 3108
rect 14465 3061 14488 3095
rect 14540 3064 14576 3103
rect 14452 3056 14488 3061
rect 14544 3056 14576 3064
rect 14400 3044 14510 3056
rect 14544 3044 14582 3056
rect 14616 3044 14628 3056
rect 14452 3022 14488 3044
rect 14544 3030 14576 3044
rect 14465 2992 14488 3022
rect 14540 2992 14576 3030
rect 14400 2988 14431 2992
rect 14465 2991 14628 2992
rect 14465 2988 14510 2991
rect 14400 2979 14510 2988
rect 14544 2979 14582 2991
rect 14616 2979 14628 2991
rect 14452 2949 14488 2979
rect 14544 2957 14576 2979
rect 14465 2927 14488 2949
rect 14540 2927 14576 2957
rect 14400 2915 14431 2927
rect 14465 2918 14628 2927
rect 14465 2915 14510 2918
rect 14400 2884 14510 2915
rect 14544 2884 14582 2918
rect 14616 2884 14628 2918
rect 14400 2876 14628 2884
rect 14400 2842 14431 2876
rect 14465 2845 14628 2876
rect 14465 2842 14510 2845
rect 14400 2811 14510 2842
rect 14544 2811 14582 2845
rect 14616 2811 14628 2845
rect 14400 2803 14628 2811
rect 14400 2769 14431 2803
rect 14465 2772 14628 2803
rect 14465 2769 14510 2772
rect 14400 2738 14510 2769
rect 14544 2738 14582 2772
rect 14616 2738 14628 2772
rect 14400 2730 14628 2738
rect 14400 2696 14431 2730
rect 14465 2699 14628 2730
rect 14465 2696 14510 2699
rect 14400 2665 14510 2696
rect 14544 2665 14582 2699
rect 14616 2665 14628 2699
rect 14400 2657 14628 2665
rect 14400 2623 14431 2657
rect 14465 2626 14628 2657
rect 14465 2623 14510 2626
rect 14400 2592 14510 2623
rect 14544 2592 14582 2626
rect 14616 2592 14628 2626
rect 14400 2584 14628 2592
rect 14400 2550 14431 2584
rect 14465 2553 14628 2584
rect 14465 2550 14510 2553
rect 14400 2519 14510 2550
rect 14544 2519 14582 2553
rect 14616 2519 14628 2553
rect 14400 2511 14628 2519
rect 14400 2477 14431 2511
rect 14465 2480 14628 2511
rect 14465 2477 14510 2480
rect 14400 2446 14510 2477
rect 14544 2446 14582 2480
rect 14616 2446 14628 2480
rect 14400 2438 14628 2446
rect 14400 2404 14431 2438
rect 14465 2407 14628 2438
rect 14465 2404 14510 2407
rect 14400 2373 14510 2404
rect 14544 2373 14582 2407
rect 14616 2373 14628 2407
rect 14400 2365 14628 2373
rect 14400 2331 14431 2365
rect 14465 2334 14628 2365
rect 14465 2331 14510 2334
rect 14400 2300 14510 2331
rect 14544 2300 14582 2334
rect 14616 2300 14628 2334
rect 14400 2292 14628 2300
rect 14400 2258 14431 2292
rect 14465 2260 14628 2292
rect 14465 2258 14510 2260
rect 14400 2226 14510 2258
rect 14544 2226 14582 2260
rect 14616 2226 14628 2260
rect 14400 2219 14628 2226
rect 14400 2185 14431 2219
rect 14465 2186 14628 2219
rect 14465 2185 14510 2186
rect 14400 2152 14510 2185
rect 14544 2152 14582 2186
rect 14616 2152 14628 2186
rect 14400 2146 14628 2152
rect 14400 2112 14431 2146
rect 14465 2112 14628 2146
rect 14400 2078 14510 2112
rect 14544 2078 14582 2112
rect 14616 2078 14628 2112
rect 14400 2073 14628 2078
rect 14400 2039 14431 2073
rect 14465 2039 14628 2073
rect 14400 2038 14628 2039
rect 14400 2004 14510 2038
rect 14544 2004 14582 2038
rect 14616 2004 14628 2038
rect 14400 2000 14628 2004
rect 14400 1966 14431 2000
rect 14465 1966 14628 2000
rect 14400 1964 14628 1966
rect 14400 1930 14510 1964
rect 14544 1930 14582 1964
rect 14616 1930 14628 1964
rect 14400 1927 14628 1930
rect 14400 1893 14431 1927
rect 14465 1893 14628 1927
rect 14400 1890 14628 1893
rect 14400 1856 14510 1890
rect 14544 1856 14582 1890
rect 14616 1856 14628 1890
rect 14400 1854 14628 1856
rect 14400 1820 14431 1854
rect 14465 1820 14628 1854
rect 14400 1816 14628 1820
rect 14400 1782 14510 1816
rect 14544 1782 14582 1816
rect 14616 1782 14628 1816
rect 14400 1781 14628 1782
rect 14400 1747 14431 1781
rect 14465 1747 14628 1781
rect 14400 1742 14628 1747
rect 14400 1708 14510 1742
rect 14544 1708 14582 1742
rect 14616 1708 14628 1742
rect 14400 1674 14431 1708
rect 14465 1674 14628 1708
rect 14400 1668 14628 1674
rect 14400 1635 14510 1668
rect 14400 1601 14431 1635
rect 14465 1634 14510 1635
rect 14544 1634 14582 1668
rect 14616 1634 14628 1668
rect 14465 1601 14628 1634
rect 14400 1594 14628 1601
rect 14400 1562 14510 1594
rect 14400 1528 14431 1562
rect 14465 1560 14510 1562
rect 14544 1560 14582 1594
rect 14616 1560 14628 1594
rect 14465 1528 14628 1560
rect 14400 1520 14628 1528
rect 14400 1489 14510 1520
rect 575 1419 803 1455
rect 575 1385 587 1419
rect 621 1385 659 1419
rect 693 1416 803 1419
rect 693 1385 733 1416
rect 575 1382 733 1385
rect 767 1382 803 1416
rect 575 1342 803 1382
rect 575 1330 733 1342
rect 575 1296 587 1330
rect 621 1296 659 1330
rect 693 1308 733 1330
rect 767 1308 803 1342
rect 14400 1455 14431 1489
rect 14465 1486 14510 1489
rect 14544 1486 14582 1520
rect 14616 1486 14628 1520
rect 14465 1455 14628 1486
rect 14400 1446 14628 1455
rect 14400 1416 14510 1446
rect 14400 1382 14431 1416
rect 14465 1412 14510 1416
rect 14544 1412 14582 1446
rect 14616 1412 14628 1446
rect 14465 1382 14628 1412
rect 14400 1372 14628 1382
rect 14400 1342 14510 1372
tri 803 1308 832 1337 sw
tri 14390 1308 14400 1318 se
rect 14400 1308 14431 1342
rect 14465 1338 14510 1342
rect 14544 1338 14582 1372
rect 14616 1338 14628 1372
rect 14465 1308 14628 1338
rect 693 1298 832 1308
tri 832 1298 842 1308 sw
tri 14380 1298 14390 1308 se
rect 14390 1298 14628 1308
rect 693 1296 842 1298
rect 575 1268 842 1296
tri 842 1268 872 1298 sw
tri 14350 1268 14380 1298 se
rect 14380 1268 14510 1298
rect 575 1241 733 1268
rect 575 1207 587 1241
rect 621 1207 659 1241
rect 693 1234 733 1241
rect 767 1234 872 1268
tri 872 1234 906 1268 sw
tri 14316 1234 14350 1268 se
rect 14350 1234 14431 1268
rect 14465 1264 14510 1268
rect 14544 1264 14582 1298
rect 14616 1264 14628 1298
rect 14465 1234 14628 1264
rect 693 1224 906 1234
tri 906 1224 916 1234 sw
tri 14306 1224 14316 1234 se
rect 14316 1224 14628 1234
rect 693 1207 916 1224
rect 575 1194 916 1207
tri 916 1194 946 1224 sw
tri 14276 1194 14306 1224 se
rect 14306 1194 14510 1224
rect 575 1160 733 1194
rect 767 1160 946 1194
tri 946 1160 980 1194 sw
tri 14242 1160 14276 1194 se
rect 14276 1160 14431 1194
rect 14465 1190 14510 1194
rect 14544 1190 14582 1224
rect 14616 1190 14628 1224
rect 14465 1160 14628 1190
rect 575 1128 980 1160
tri 980 1128 1012 1160 sw
tri 14230 1148 14242 1160 se
rect 14242 1148 14628 1160
tri 14210 1128 14230 1148 se
rect 14230 1128 14628 1148
rect 575 1116 14628 1128
rect 575 1114 767 1116
tri 575 1082 607 1114 ne
rect 607 1082 767 1114
rect 801 1082 840 1116
rect 874 1082 913 1116
rect 947 1082 986 1116
rect 1020 1082 1059 1116
rect 1093 1082 1132 1116
rect 1166 1082 1205 1116
rect 1239 1082 1278 1116
rect 1312 1082 1351 1116
rect 1385 1082 1424 1116
rect 1458 1082 1497 1116
rect 1531 1082 1570 1116
rect 1604 1082 1643 1116
rect 1677 1082 1716 1116
rect 1750 1082 1789 1116
rect 1823 1082 1862 1116
rect 1896 1082 1935 1116
rect 1969 1082 2008 1116
rect 2042 1082 2081 1116
rect 2115 1082 2154 1116
rect 2188 1082 2227 1116
rect 2261 1082 2300 1116
rect 2334 1082 2373 1116
rect 2407 1082 2446 1116
rect 2480 1082 2519 1116
rect 2553 1082 2592 1116
rect 2626 1082 2665 1116
rect 2699 1082 2738 1116
tri 607 1044 645 1082 ne
rect 645 1044 2738 1082
tri 645 1010 679 1044 ne
rect 679 1010 767 1044
rect 801 1010 840 1044
rect 874 1010 913 1044
rect 947 1010 986 1044
rect 1020 1010 1059 1044
rect 1093 1010 1132 1044
rect 1166 1010 1205 1044
rect 1239 1010 1278 1044
rect 1312 1010 1351 1044
rect 1385 1010 1424 1044
rect 1458 1010 1497 1044
rect 1531 1010 1570 1044
rect 1604 1010 1643 1044
rect 1677 1010 1716 1044
rect 1750 1010 1789 1044
rect 1823 1010 1862 1044
rect 1896 1010 1935 1044
rect 1969 1010 2008 1044
rect 2042 1010 2081 1044
rect 2115 1010 2154 1044
rect 2188 1010 2227 1044
rect 2261 1010 2300 1044
rect 2334 1010 2373 1044
rect 2407 1010 2446 1044
rect 2480 1010 2519 1044
rect 2553 1010 2592 1044
rect 2626 1010 2665 1044
rect 2699 1010 2738 1044
rect 14436 1114 14628 1116
rect 14436 1010 14512 1114
tri 679 998 691 1010 ne
rect 691 998 14512 1010
tri 14512 998 14628 1114 nw
tri 14914 862 14915 863 se
rect 14915 862 14927 4960
tri 261 680 443 862 sw
tri 14732 680 14914 862 se
rect 14914 680 14927 862
rect 249 668 14927 680
rect 249 496 308 668
rect 59 490 308 496
rect 14886 490 14927 668
rect 15105 490 15117 5420
rect 59 478 15117 490
<< via1 >>
rect 575 4050 587 4068
rect 587 4050 621 4068
rect 621 4050 627 4068
rect 663 4050 693 4068
rect 693 4050 715 4068
rect 575 4016 627 4050
rect 663 4016 715 4050
rect 751 4044 803 4068
rect 751 4016 767 4044
rect 767 4016 803 4044
rect 575 3977 587 4004
rect 587 3977 621 4004
rect 621 3977 627 4004
rect 663 3977 693 4004
rect 693 3977 715 4004
rect 575 3952 627 3977
rect 663 3952 715 3977
rect 751 3971 803 4004
rect 751 3952 767 3971
rect 767 3952 803 3971
rect 575 3938 627 3940
rect 663 3938 715 3940
rect 575 3904 587 3938
rect 587 3904 621 3938
rect 621 3904 627 3938
rect 663 3904 693 3938
rect 693 3904 715 3938
rect 751 3937 767 3940
rect 767 3937 803 3940
rect 575 3888 627 3904
rect 663 3888 715 3904
rect 751 3898 803 3937
rect 751 3888 767 3898
rect 767 3888 803 3898
rect 575 3865 627 3876
rect 663 3865 715 3876
rect 575 3831 587 3865
rect 587 3831 621 3865
rect 621 3831 627 3865
rect 663 3831 693 3865
rect 693 3831 715 3865
rect 751 3864 767 3876
rect 767 3864 803 3876
rect 575 3824 627 3831
rect 663 3824 715 3831
rect 751 3825 803 3864
rect 751 3824 767 3825
rect 767 3824 803 3825
rect 575 3792 627 3812
rect 663 3792 715 3812
rect 575 3760 587 3792
rect 587 3760 621 3792
rect 621 3760 627 3792
rect 663 3760 693 3792
rect 693 3760 715 3792
rect 751 3791 767 3812
rect 767 3791 803 3812
rect 751 3760 803 3791
rect 575 3719 627 3748
rect 663 3719 715 3748
rect 575 3696 587 3719
rect 587 3696 621 3719
rect 621 3696 627 3719
rect 663 3696 693 3719
rect 693 3696 715 3719
rect 751 3718 767 3748
rect 767 3718 803 3748
rect 751 3696 803 3718
rect 575 3646 627 3684
rect 663 3646 715 3684
rect 751 3679 803 3684
rect 575 3632 587 3646
rect 587 3632 621 3646
rect 621 3632 627 3646
rect 663 3632 693 3646
rect 693 3632 715 3646
rect 751 3645 767 3679
rect 767 3645 803 3679
rect 751 3632 803 3645
rect 575 3612 587 3620
rect 587 3612 621 3620
rect 621 3612 627 3620
rect 663 3612 693 3620
rect 693 3612 715 3620
rect 575 3573 627 3612
rect 663 3573 715 3612
rect 751 3606 803 3620
rect 575 3568 587 3573
rect 587 3568 621 3573
rect 621 3568 627 3573
rect 663 3568 693 3573
rect 693 3568 715 3573
rect 751 3572 767 3606
rect 767 3572 803 3606
rect 751 3568 803 3572
rect 575 3539 587 3556
rect 587 3539 621 3556
rect 621 3539 627 3556
rect 663 3539 693 3556
rect 693 3539 715 3556
rect 575 3504 627 3539
rect 663 3504 715 3539
rect 751 3533 803 3556
rect 751 3504 767 3533
rect 767 3504 803 3533
rect 575 3466 587 3492
rect 587 3466 621 3492
rect 621 3466 627 3492
rect 663 3466 693 3492
rect 693 3466 715 3492
rect 575 3440 627 3466
rect 663 3440 715 3466
rect 751 3460 803 3492
rect 751 3440 767 3460
rect 767 3440 803 3460
rect 575 3427 627 3428
rect 663 3427 715 3428
rect 575 3393 587 3427
rect 587 3393 621 3427
rect 621 3393 627 3427
rect 663 3393 693 3427
rect 693 3393 715 3427
rect 751 3426 767 3428
rect 767 3426 803 3428
rect 575 3376 627 3393
rect 663 3376 715 3393
rect 751 3387 803 3426
rect 751 3376 767 3387
rect 767 3376 803 3387
rect 575 3354 627 3364
rect 663 3354 715 3364
rect 575 3320 587 3354
rect 587 3320 621 3354
rect 621 3320 627 3354
rect 663 3320 693 3354
rect 693 3320 715 3354
rect 751 3353 767 3364
rect 767 3353 803 3364
rect 575 3312 627 3320
rect 663 3312 715 3320
rect 751 3314 803 3353
rect 751 3312 767 3314
rect 767 3312 803 3314
rect 575 3281 627 3300
rect 663 3281 715 3300
rect 575 3248 587 3281
rect 587 3248 621 3281
rect 621 3248 627 3281
rect 663 3248 693 3281
rect 693 3248 715 3281
rect 751 3280 767 3300
rect 767 3280 803 3300
rect 751 3248 803 3280
rect 575 3208 627 3236
rect 663 3208 715 3236
rect 575 3184 587 3208
rect 587 3184 621 3208
rect 621 3184 627 3208
rect 663 3184 693 3208
rect 693 3184 715 3208
rect 751 3207 767 3236
rect 767 3207 803 3236
rect 751 3184 803 3207
rect 575 3135 627 3172
rect 663 3135 715 3172
rect 751 3168 803 3172
rect 575 3120 587 3135
rect 587 3120 621 3135
rect 621 3120 627 3135
rect 663 3120 693 3135
rect 693 3120 715 3135
rect 751 3134 767 3168
rect 767 3134 803 3168
rect 751 3120 803 3134
rect 575 3101 587 3108
rect 587 3101 621 3108
rect 621 3101 627 3108
rect 663 3101 693 3108
rect 693 3101 715 3108
rect 575 3062 627 3101
rect 663 3062 715 3101
rect 751 3095 803 3108
rect 575 3056 587 3062
rect 587 3056 621 3062
rect 621 3056 627 3062
rect 663 3056 693 3062
rect 693 3056 715 3062
rect 751 3061 767 3095
rect 767 3061 803 3095
rect 751 3056 803 3061
rect 575 3028 587 3044
rect 587 3028 621 3044
rect 621 3028 627 3044
rect 663 3028 693 3044
rect 693 3028 715 3044
rect 575 2992 627 3028
rect 663 2992 715 3028
rect 751 3022 803 3044
rect 751 2992 767 3022
rect 767 2992 803 3022
rect 575 2955 587 2979
rect 587 2955 621 2979
rect 621 2955 627 2979
rect 663 2955 693 2979
rect 693 2955 715 2979
rect 575 2927 627 2955
rect 663 2927 715 2955
rect 751 2949 803 2979
rect 751 2927 767 2949
rect 767 2927 803 2949
rect 1109 2582 1289 2614
rect 1109 2548 1110 2582
rect 1110 2548 1144 2582
rect 1144 2548 1182 2582
rect 1182 2548 1216 2582
rect 1216 2548 1254 2582
rect 1254 2548 1288 2582
rect 1288 2548 1289 2582
rect 1109 2508 1289 2548
rect 1109 2474 1110 2508
rect 1110 2474 1144 2508
rect 1144 2474 1182 2508
rect 1182 2474 1216 2508
rect 1216 2474 1254 2508
rect 1254 2474 1288 2508
rect 1288 2474 1289 2508
rect 1109 2434 1289 2474
rect 1109 2400 1110 2434
rect 1110 2400 1144 2434
rect 1144 2400 1182 2434
rect 1182 2400 1216 2434
rect 1216 2400 1254 2434
rect 1254 2400 1288 2434
rect 1288 2400 1289 2434
rect 1109 2360 1289 2400
rect 1109 2326 1110 2360
rect 1110 2326 1144 2360
rect 1144 2326 1182 2360
rect 1182 2326 1216 2360
rect 1216 2326 1254 2360
rect 1254 2326 1288 2360
rect 1288 2326 1289 2360
rect 1109 2286 1289 2326
rect 1109 2252 1110 2286
rect 1110 2252 1144 2286
rect 1144 2252 1182 2286
rect 1182 2252 1216 2286
rect 1216 2252 1254 2286
rect 1254 2252 1288 2286
rect 1288 2252 1289 2286
rect 1109 2212 1289 2252
rect 1109 2178 1110 2212
rect 1110 2178 1144 2212
rect 1144 2178 1182 2212
rect 1182 2178 1216 2212
rect 1216 2178 1254 2212
rect 1254 2178 1288 2212
rect 1288 2178 1289 2212
rect 1109 2138 1289 2178
rect 1109 2104 1110 2138
rect 1110 2104 1144 2138
rect 1144 2104 1182 2138
rect 1182 2104 1216 2138
rect 1216 2104 1254 2138
rect 1254 2104 1288 2138
rect 1288 2104 1289 2138
rect 1109 2064 1289 2104
rect 1109 2030 1110 2064
rect 1110 2030 1144 2064
rect 1144 2030 1182 2064
rect 1182 2030 1216 2064
rect 1216 2030 1254 2064
rect 1254 2030 1288 2064
rect 1288 2030 1289 2064
rect 1109 1990 1289 2030
rect 1109 1956 1110 1990
rect 1110 1956 1144 1990
rect 1144 1956 1182 1990
rect 1182 1956 1216 1990
rect 1216 1956 1254 1990
rect 1254 1956 1288 1990
rect 1288 1956 1289 1990
rect 1109 1916 1289 1956
rect 1109 1882 1110 1916
rect 1110 1882 1144 1916
rect 1144 1882 1182 1916
rect 1182 1882 1216 1916
rect 1216 1882 1254 1916
rect 1254 1882 1288 1916
rect 1288 1882 1289 1916
rect 1109 1842 1289 1882
rect 1109 1808 1110 1842
rect 1110 1808 1144 1842
rect 1144 1808 1182 1842
rect 1182 1808 1216 1842
rect 1216 1808 1254 1842
rect 1254 1808 1288 1842
rect 1288 1808 1289 1842
rect 1109 1768 1289 1808
rect 1109 1734 1110 1768
rect 1110 1734 1144 1768
rect 1144 1734 1182 1768
rect 1182 1734 1216 1768
rect 1216 1734 1254 1768
rect 1254 1734 1288 1768
rect 1288 1734 1289 1768
rect 1109 1694 1289 1734
rect 1109 1660 1110 1694
rect 1110 1660 1144 1694
rect 1144 1660 1182 1694
rect 1182 1660 1216 1694
rect 1216 1660 1254 1694
rect 1254 1660 1288 1694
rect 1288 1660 1289 1694
rect 1109 1620 1289 1660
rect 1109 1586 1110 1620
rect 1110 1586 1144 1620
rect 1144 1586 1182 1620
rect 1182 1586 1216 1620
rect 1216 1586 1254 1620
rect 1254 1586 1288 1620
rect 1288 1586 1289 1620
rect 1109 1545 1289 1586
rect 1109 1538 1110 1545
rect 1110 1538 1144 1545
rect 1144 1538 1182 1545
rect 1182 1538 1216 1545
rect 1216 1538 1254 1545
rect 1254 1538 1288 1545
rect 1288 1538 1289 1545
rect 1109 1511 1110 1525
rect 1110 1511 1144 1525
rect 1144 1511 1161 1525
rect 1109 1473 1161 1511
rect 1173 1511 1182 1525
rect 1182 1511 1216 1525
rect 1216 1511 1225 1525
rect 1173 1473 1225 1511
rect 1237 1511 1254 1525
rect 1254 1511 1288 1525
rect 1288 1511 1289 1525
rect 1237 1473 1289 1511
rect 1605 4062 1785 4068
rect 1605 4050 1678 4062
rect 1678 4050 1712 4062
rect 1712 4050 1785 4062
rect 1605 3080 1606 4050
rect 1606 3092 1784 4050
rect 1606 3080 1640 3092
rect 1640 3080 1750 3092
rect 1750 3080 1784 3092
rect 1784 3080 1785 4050
rect 1605 3040 1785 3080
rect 1605 2992 1606 3040
rect 1606 2992 1784 3040
rect 1784 2992 1785 3040
rect 1605 2927 1606 2979
rect 1606 2927 1657 2979
rect 1669 2927 1721 2979
rect 1733 2927 1784 2979
rect 1784 2927 1785 2979
rect 2101 2582 2281 2614
rect 2101 2548 2102 2582
rect 2102 2548 2136 2582
rect 2136 2548 2174 2582
rect 2174 2548 2208 2582
rect 2208 2548 2246 2582
rect 2246 2548 2280 2582
rect 2280 2548 2281 2582
rect 2101 2508 2281 2548
rect 2101 2474 2102 2508
rect 2102 2474 2136 2508
rect 2136 2474 2174 2508
rect 2174 2474 2208 2508
rect 2208 2474 2246 2508
rect 2246 2474 2280 2508
rect 2280 2474 2281 2508
rect 2101 2434 2281 2474
rect 2101 2400 2102 2434
rect 2102 2400 2136 2434
rect 2136 2400 2174 2434
rect 2174 2400 2208 2434
rect 2208 2400 2246 2434
rect 2246 2400 2280 2434
rect 2280 2400 2281 2434
rect 2101 2360 2281 2400
rect 2101 2326 2102 2360
rect 2102 2326 2136 2360
rect 2136 2326 2174 2360
rect 2174 2326 2208 2360
rect 2208 2326 2246 2360
rect 2246 2326 2280 2360
rect 2280 2326 2281 2360
rect 2101 2286 2281 2326
rect 2101 2252 2102 2286
rect 2102 2252 2136 2286
rect 2136 2252 2174 2286
rect 2174 2252 2208 2286
rect 2208 2252 2246 2286
rect 2246 2252 2280 2286
rect 2280 2252 2281 2286
rect 2101 2212 2281 2252
rect 2101 2178 2102 2212
rect 2102 2178 2136 2212
rect 2136 2178 2174 2212
rect 2174 2178 2208 2212
rect 2208 2178 2246 2212
rect 2246 2178 2280 2212
rect 2280 2178 2281 2212
rect 2101 2138 2281 2178
rect 2101 2104 2102 2138
rect 2102 2104 2136 2138
rect 2136 2104 2174 2138
rect 2174 2104 2208 2138
rect 2208 2104 2246 2138
rect 2246 2104 2280 2138
rect 2280 2104 2281 2138
rect 2101 2064 2281 2104
rect 2101 2030 2102 2064
rect 2102 2030 2136 2064
rect 2136 2030 2174 2064
rect 2174 2030 2208 2064
rect 2208 2030 2246 2064
rect 2246 2030 2280 2064
rect 2280 2030 2281 2064
rect 2101 1990 2281 2030
rect 2101 1956 2102 1990
rect 2102 1956 2136 1990
rect 2136 1956 2174 1990
rect 2174 1956 2208 1990
rect 2208 1956 2246 1990
rect 2246 1956 2280 1990
rect 2280 1956 2281 1990
rect 2101 1916 2281 1956
rect 2101 1882 2102 1916
rect 2102 1882 2136 1916
rect 2136 1882 2174 1916
rect 2174 1882 2208 1916
rect 2208 1882 2246 1916
rect 2246 1882 2280 1916
rect 2280 1882 2281 1916
rect 2101 1842 2281 1882
rect 2101 1808 2102 1842
rect 2102 1808 2136 1842
rect 2136 1808 2174 1842
rect 2174 1808 2208 1842
rect 2208 1808 2246 1842
rect 2246 1808 2280 1842
rect 2280 1808 2281 1842
rect 2101 1768 2281 1808
rect 2101 1734 2102 1768
rect 2102 1734 2136 1768
rect 2136 1734 2174 1768
rect 2174 1734 2208 1768
rect 2208 1734 2246 1768
rect 2246 1734 2280 1768
rect 2280 1734 2281 1768
rect 2101 1694 2281 1734
rect 2101 1660 2102 1694
rect 2102 1660 2136 1694
rect 2136 1660 2174 1694
rect 2174 1660 2208 1694
rect 2208 1660 2246 1694
rect 2246 1660 2280 1694
rect 2280 1660 2281 1694
rect 2101 1620 2281 1660
rect 2101 1586 2102 1620
rect 2102 1586 2136 1620
rect 2136 1586 2174 1620
rect 2174 1586 2208 1620
rect 2208 1586 2246 1620
rect 2246 1586 2280 1620
rect 2280 1586 2281 1620
rect 2101 1545 2281 1586
rect 2101 1538 2102 1545
rect 2102 1538 2136 1545
rect 2136 1538 2174 1545
rect 2174 1538 2208 1545
rect 2208 1538 2246 1545
rect 2246 1538 2280 1545
rect 2280 1538 2281 1545
rect 2101 1511 2102 1525
rect 2102 1511 2136 1525
rect 2136 1511 2153 1525
rect 2101 1473 2153 1511
rect 2165 1511 2174 1525
rect 2174 1511 2208 1525
rect 2208 1511 2217 1525
rect 2165 1473 2217 1511
rect 2229 1511 2246 1525
rect 2246 1511 2280 1525
rect 2280 1511 2281 1525
rect 2229 1473 2281 1511
rect 2597 4062 2777 4068
rect 2597 4050 2670 4062
rect 2670 4050 2704 4062
rect 2704 4050 2777 4062
rect 2597 3080 2598 4050
rect 2598 3092 2776 4050
rect 2598 3080 2632 3092
rect 2632 3080 2742 3092
rect 2742 3080 2776 3092
rect 2776 3080 2777 4050
rect 2597 3040 2777 3080
rect 2597 2992 2598 3040
rect 2598 2992 2776 3040
rect 2776 2992 2777 3040
rect 2597 2927 2598 2979
rect 2598 2927 2649 2979
rect 2661 2927 2713 2979
rect 2725 2927 2776 2979
rect 2776 2927 2777 2979
rect 3093 2582 3273 2614
rect 3093 2548 3094 2582
rect 3094 2548 3128 2582
rect 3128 2548 3166 2582
rect 3166 2548 3200 2582
rect 3200 2548 3238 2582
rect 3238 2548 3272 2582
rect 3272 2548 3273 2582
rect 3093 2508 3273 2548
rect 3093 2474 3094 2508
rect 3094 2474 3128 2508
rect 3128 2474 3166 2508
rect 3166 2474 3200 2508
rect 3200 2474 3238 2508
rect 3238 2474 3272 2508
rect 3272 2474 3273 2508
rect 3093 2434 3273 2474
rect 3093 2400 3094 2434
rect 3094 2400 3128 2434
rect 3128 2400 3166 2434
rect 3166 2400 3200 2434
rect 3200 2400 3238 2434
rect 3238 2400 3272 2434
rect 3272 2400 3273 2434
rect 3093 2360 3273 2400
rect 3093 2326 3094 2360
rect 3094 2326 3128 2360
rect 3128 2326 3166 2360
rect 3166 2326 3200 2360
rect 3200 2326 3238 2360
rect 3238 2326 3272 2360
rect 3272 2326 3273 2360
rect 3093 2286 3273 2326
rect 3093 2252 3094 2286
rect 3094 2252 3128 2286
rect 3128 2252 3166 2286
rect 3166 2252 3200 2286
rect 3200 2252 3238 2286
rect 3238 2252 3272 2286
rect 3272 2252 3273 2286
rect 3093 2212 3273 2252
rect 3093 2178 3094 2212
rect 3094 2178 3128 2212
rect 3128 2178 3166 2212
rect 3166 2178 3200 2212
rect 3200 2178 3238 2212
rect 3238 2178 3272 2212
rect 3272 2178 3273 2212
rect 3093 2138 3273 2178
rect 3093 2104 3094 2138
rect 3094 2104 3128 2138
rect 3128 2104 3166 2138
rect 3166 2104 3200 2138
rect 3200 2104 3238 2138
rect 3238 2104 3272 2138
rect 3272 2104 3273 2138
rect 3093 2064 3273 2104
rect 3093 2030 3094 2064
rect 3094 2030 3128 2064
rect 3128 2030 3166 2064
rect 3166 2030 3200 2064
rect 3200 2030 3238 2064
rect 3238 2030 3272 2064
rect 3272 2030 3273 2064
rect 3093 1990 3273 2030
rect 3093 1956 3094 1990
rect 3094 1956 3128 1990
rect 3128 1956 3166 1990
rect 3166 1956 3200 1990
rect 3200 1956 3238 1990
rect 3238 1956 3272 1990
rect 3272 1956 3273 1990
rect 3093 1916 3273 1956
rect 3093 1882 3094 1916
rect 3094 1882 3128 1916
rect 3128 1882 3166 1916
rect 3166 1882 3200 1916
rect 3200 1882 3238 1916
rect 3238 1882 3272 1916
rect 3272 1882 3273 1916
rect 3093 1842 3273 1882
rect 3093 1808 3094 1842
rect 3094 1808 3128 1842
rect 3128 1808 3166 1842
rect 3166 1808 3200 1842
rect 3200 1808 3238 1842
rect 3238 1808 3272 1842
rect 3272 1808 3273 1842
rect 3093 1768 3273 1808
rect 3093 1734 3094 1768
rect 3094 1734 3128 1768
rect 3128 1734 3166 1768
rect 3166 1734 3200 1768
rect 3200 1734 3238 1768
rect 3238 1734 3272 1768
rect 3272 1734 3273 1768
rect 3093 1694 3273 1734
rect 3093 1660 3094 1694
rect 3094 1660 3128 1694
rect 3128 1660 3166 1694
rect 3166 1660 3200 1694
rect 3200 1660 3238 1694
rect 3238 1660 3272 1694
rect 3272 1660 3273 1694
rect 3093 1620 3273 1660
rect 3093 1586 3094 1620
rect 3094 1586 3128 1620
rect 3128 1586 3166 1620
rect 3166 1586 3200 1620
rect 3200 1586 3238 1620
rect 3238 1586 3272 1620
rect 3272 1586 3273 1620
rect 3093 1545 3273 1586
rect 3093 1538 3094 1545
rect 3094 1538 3128 1545
rect 3128 1538 3166 1545
rect 3166 1538 3200 1545
rect 3200 1538 3238 1545
rect 3238 1538 3272 1545
rect 3272 1538 3273 1545
rect 3093 1511 3094 1525
rect 3094 1511 3128 1525
rect 3128 1511 3145 1525
rect 3093 1473 3145 1511
rect 3157 1511 3166 1525
rect 3166 1511 3200 1525
rect 3200 1511 3209 1525
rect 3157 1473 3209 1511
rect 3221 1511 3238 1525
rect 3238 1511 3272 1525
rect 3272 1511 3273 1525
rect 3221 1473 3273 1511
rect 3589 4062 3769 4068
rect 3589 4050 3662 4062
rect 3662 4050 3696 4062
rect 3696 4050 3769 4062
rect 3589 3080 3590 4050
rect 3590 3092 3768 4050
rect 3590 3080 3624 3092
rect 3624 3080 3734 3092
rect 3734 3080 3768 3092
rect 3768 3080 3769 4050
rect 3589 3040 3769 3080
rect 3589 2992 3590 3040
rect 3590 2992 3768 3040
rect 3768 2992 3769 3040
rect 3589 2927 3590 2979
rect 3590 2927 3641 2979
rect 3653 2927 3705 2979
rect 3717 2927 3768 2979
rect 3768 2927 3769 2979
rect 4085 2582 4265 2614
rect 4085 2548 4086 2582
rect 4086 2548 4120 2582
rect 4120 2548 4158 2582
rect 4158 2548 4192 2582
rect 4192 2548 4230 2582
rect 4230 2548 4264 2582
rect 4264 2548 4265 2582
rect 4085 2508 4265 2548
rect 4085 2474 4086 2508
rect 4086 2474 4120 2508
rect 4120 2474 4158 2508
rect 4158 2474 4192 2508
rect 4192 2474 4230 2508
rect 4230 2474 4264 2508
rect 4264 2474 4265 2508
rect 4085 2434 4265 2474
rect 4085 2400 4086 2434
rect 4086 2400 4120 2434
rect 4120 2400 4158 2434
rect 4158 2400 4192 2434
rect 4192 2400 4230 2434
rect 4230 2400 4264 2434
rect 4264 2400 4265 2434
rect 4085 2360 4265 2400
rect 4085 2326 4086 2360
rect 4086 2326 4120 2360
rect 4120 2326 4158 2360
rect 4158 2326 4192 2360
rect 4192 2326 4230 2360
rect 4230 2326 4264 2360
rect 4264 2326 4265 2360
rect 4085 2286 4265 2326
rect 4085 2252 4086 2286
rect 4086 2252 4120 2286
rect 4120 2252 4158 2286
rect 4158 2252 4192 2286
rect 4192 2252 4230 2286
rect 4230 2252 4264 2286
rect 4264 2252 4265 2286
rect 4085 2212 4265 2252
rect 4085 2178 4086 2212
rect 4086 2178 4120 2212
rect 4120 2178 4158 2212
rect 4158 2178 4192 2212
rect 4192 2178 4230 2212
rect 4230 2178 4264 2212
rect 4264 2178 4265 2212
rect 4085 2138 4265 2178
rect 4085 2104 4086 2138
rect 4086 2104 4120 2138
rect 4120 2104 4158 2138
rect 4158 2104 4192 2138
rect 4192 2104 4230 2138
rect 4230 2104 4264 2138
rect 4264 2104 4265 2138
rect 4085 2064 4265 2104
rect 4085 2030 4086 2064
rect 4086 2030 4120 2064
rect 4120 2030 4158 2064
rect 4158 2030 4192 2064
rect 4192 2030 4230 2064
rect 4230 2030 4264 2064
rect 4264 2030 4265 2064
rect 4085 1990 4265 2030
rect 4085 1956 4086 1990
rect 4086 1956 4120 1990
rect 4120 1956 4158 1990
rect 4158 1956 4192 1990
rect 4192 1956 4230 1990
rect 4230 1956 4264 1990
rect 4264 1956 4265 1990
rect 4085 1916 4265 1956
rect 4085 1882 4086 1916
rect 4086 1882 4120 1916
rect 4120 1882 4158 1916
rect 4158 1882 4192 1916
rect 4192 1882 4230 1916
rect 4230 1882 4264 1916
rect 4264 1882 4265 1916
rect 4085 1842 4265 1882
rect 4085 1808 4086 1842
rect 4086 1808 4120 1842
rect 4120 1808 4158 1842
rect 4158 1808 4192 1842
rect 4192 1808 4230 1842
rect 4230 1808 4264 1842
rect 4264 1808 4265 1842
rect 4085 1768 4265 1808
rect 4085 1734 4086 1768
rect 4086 1734 4120 1768
rect 4120 1734 4158 1768
rect 4158 1734 4192 1768
rect 4192 1734 4230 1768
rect 4230 1734 4264 1768
rect 4264 1734 4265 1768
rect 4085 1694 4265 1734
rect 4085 1660 4086 1694
rect 4086 1660 4120 1694
rect 4120 1660 4158 1694
rect 4158 1660 4192 1694
rect 4192 1660 4230 1694
rect 4230 1660 4264 1694
rect 4264 1660 4265 1694
rect 4085 1620 4265 1660
rect 4085 1586 4086 1620
rect 4086 1586 4120 1620
rect 4120 1586 4158 1620
rect 4158 1586 4192 1620
rect 4192 1586 4230 1620
rect 4230 1586 4264 1620
rect 4264 1586 4265 1620
rect 4085 1545 4265 1586
rect 4085 1538 4086 1545
rect 4086 1538 4120 1545
rect 4120 1538 4158 1545
rect 4158 1538 4192 1545
rect 4192 1538 4230 1545
rect 4230 1538 4264 1545
rect 4264 1538 4265 1545
rect 4085 1511 4086 1525
rect 4086 1511 4120 1525
rect 4120 1511 4137 1525
rect 4085 1473 4137 1511
rect 4149 1511 4158 1525
rect 4158 1511 4192 1525
rect 4192 1511 4201 1525
rect 4149 1473 4201 1511
rect 4213 1511 4230 1525
rect 4230 1511 4264 1525
rect 4264 1511 4265 1525
rect 4213 1473 4265 1511
rect 4581 4062 4761 4068
rect 4581 4050 4654 4062
rect 4654 4050 4688 4062
rect 4688 4050 4761 4062
rect 4581 3080 4582 4050
rect 4582 3092 4760 4050
rect 4582 3080 4616 3092
rect 4616 3080 4726 3092
rect 4726 3080 4760 3092
rect 4760 3080 4761 4050
rect 4581 3040 4761 3080
rect 4581 2992 4582 3040
rect 4582 2992 4760 3040
rect 4760 2992 4761 3040
rect 4581 2927 4582 2979
rect 4582 2927 4633 2979
rect 4645 2927 4697 2979
rect 4709 2927 4760 2979
rect 4760 2927 4761 2979
rect 5077 2582 5257 2614
rect 5077 2548 5078 2582
rect 5078 2548 5112 2582
rect 5112 2548 5150 2582
rect 5150 2548 5184 2582
rect 5184 2548 5222 2582
rect 5222 2548 5256 2582
rect 5256 2548 5257 2582
rect 5077 2508 5257 2548
rect 5077 2474 5078 2508
rect 5078 2474 5112 2508
rect 5112 2474 5150 2508
rect 5150 2474 5184 2508
rect 5184 2474 5222 2508
rect 5222 2474 5256 2508
rect 5256 2474 5257 2508
rect 5077 2434 5257 2474
rect 5077 2400 5078 2434
rect 5078 2400 5112 2434
rect 5112 2400 5150 2434
rect 5150 2400 5184 2434
rect 5184 2400 5222 2434
rect 5222 2400 5256 2434
rect 5256 2400 5257 2434
rect 5077 2360 5257 2400
rect 5077 2326 5078 2360
rect 5078 2326 5112 2360
rect 5112 2326 5150 2360
rect 5150 2326 5184 2360
rect 5184 2326 5222 2360
rect 5222 2326 5256 2360
rect 5256 2326 5257 2360
rect 5077 2286 5257 2326
rect 5077 2252 5078 2286
rect 5078 2252 5112 2286
rect 5112 2252 5150 2286
rect 5150 2252 5184 2286
rect 5184 2252 5222 2286
rect 5222 2252 5256 2286
rect 5256 2252 5257 2286
rect 5077 2212 5257 2252
rect 5077 2178 5078 2212
rect 5078 2178 5112 2212
rect 5112 2178 5150 2212
rect 5150 2178 5184 2212
rect 5184 2178 5222 2212
rect 5222 2178 5256 2212
rect 5256 2178 5257 2212
rect 5077 2138 5257 2178
rect 5077 2104 5078 2138
rect 5078 2104 5112 2138
rect 5112 2104 5150 2138
rect 5150 2104 5184 2138
rect 5184 2104 5222 2138
rect 5222 2104 5256 2138
rect 5256 2104 5257 2138
rect 5077 2064 5257 2104
rect 5077 2030 5078 2064
rect 5078 2030 5112 2064
rect 5112 2030 5150 2064
rect 5150 2030 5184 2064
rect 5184 2030 5222 2064
rect 5222 2030 5256 2064
rect 5256 2030 5257 2064
rect 5077 1990 5257 2030
rect 5077 1956 5078 1990
rect 5078 1956 5112 1990
rect 5112 1956 5150 1990
rect 5150 1956 5184 1990
rect 5184 1956 5222 1990
rect 5222 1956 5256 1990
rect 5256 1956 5257 1990
rect 5077 1916 5257 1956
rect 5077 1882 5078 1916
rect 5078 1882 5112 1916
rect 5112 1882 5150 1916
rect 5150 1882 5184 1916
rect 5184 1882 5222 1916
rect 5222 1882 5256 1916
rect 5256 1882 5257 1916
rect 5077 1842 5257 1882
rect 5077 1808 5078 1842
rect 5078 1808 5112 1842
rect 5112 1808 5150 1842
rect 5150 1808 5184 1842
rect 5184 1808 5222 1842
rect 5222 1808 5256 1842
rect 5256 1808 5257 1842
rect 5077 1768 5257 1808
rect 5077 1734 5078 1768
rect 5078 1734 5112 1768
rect 5112 1734 5150 1768
rect 5150 1734 5184 1768
rect 5184 1734 5222 1768
rect 5222 1734 5256 1768
rect 5256 1734 5257 1768
rect 5077 1694 5257 1734
rect 5077 1660 5078 1694
rect 5078 1660 5112 1694
rect 5112 1660 5150 1694
rect 5150 1660 5184 1694
rect 5184 1660 5222 1694
rect 5222 1660 5256 1694
rect 5256 1660 5257 1694
rect 5077 1620 5257 1660
rect 5077 1586 5078 1620
rect 5078 1586 5112 1620
rect 5112 1586 5150 1620
rect 5150 1586 5184 1620
rect 5184 1586 5222 1620
rect 5222 1586 5256 1620
rect 5256 1586 5257 1620
rect 5077 1545 5257 1586
rect 5077 1538 5078 1545
rect 5078 1538 5112 1545
rect 5112 1538 5150 1545
rect 5150 1538 5184 1545
rect 5184 1538 5222 1545
rect 5222 1538 5256 1545
rect 5256 1538 5257 1545
rect 5077 1511 5078 1525
rect 5078 1511 5112 1525
rect 5112 1511 5129 1525
rect 5077 1473 5129 1511
rect 5141 1511 5150 1525
rect 5150 1511 5184 1525
rect 5184 1511 5193 1525
rect 5141 1473 5193 1511
rect 5205 1511 5222 1525
rect 5222 1511 5256 1525
rect 5256 1511 5257 1525
rect 5205 1473 5257 1511
rect 5573 4062 5753 4068
rect 5573 4050 5646 4062
rect 5646 4050 5680 4062
rect 5680 4050 5753 4062
rect 5573 3080 5574 4050
rect 5574 3092 5752 4050
rect 5574 3080 5608 3092
rect 5608 3080 5718 3092
rect 5718 3080 5752 3092
rect 5752 3080 5753 4050
rect 5573 3040 5753 3080
rect 5573 2992 5574 3040
rect 5574 2992 5752 3040
rect 5752 2992 5753 3040
rect 5573 2927 5574 2979
rect 5574 2927 5625 2979
rect 5637 2927 5689 2979
rect 5701 2927 5752 2979
rect 5752 2927 5753 2979
rect 6069 2582 6249 2614
rect 6069 2548 6070 2582
rect 6070 2548 6104 2582
rect 6104 2548 6142 2582
rect 6142 2548 6176 2582
rect 6176 2548 6214 2582
rect 6214 2548 6248 2582
rect 6248 2548 6249 2582
rect 6069 2508 6249 2548
rect 6069 2474 6070 2508
rect 6070 2474 6104 2508
rect 6104 2474 6142 2508
rect 6142 2474 6176 2508
rect 6176 2474 6214 2508
rect 6214 2474 6248 2508
rect 6248 2474 6249 2508
rect 6069 2434 6249 2474
rect 6069 2400 6070 2434
rect 6070 2400 6104 2434
rect 6104 2400 6142 2434
rect 6142 2400 6176 2434
rect 6176 2400 6214 2434
rect 6214 2400 6248 2434
rect 6248 2400 6249 2434
rect 6069 2360 6249 2400
rect 6069 2326 6070 2360
rect 6070 2326 6104 2360
rect 6104 2326 6142 2360
rect 6142 2326 6176 2360
rect 6176 2326 6214 2360
rect 6214 2326 6248 2360
rect 6248 2326 6249 2360
rect 6069 2286 6249 2326
rect 6069 2252 6070 2286
rect 6070 2252 6104 2286
rect 6104 2252 6142 2286
rect 6142 2252 6176 2286
rect 6176 2252 6214 2286
rect 6214 2252 6248 2286
rect 6248 2252 6249 2286
rect 6069 2212 6249 2252
rect 6069 2178 6070 2212
rect 6070 2178 6104 2212
rect 6104 2178 6142 2212
rect 6142 2178 6176 2212
rect 6176 2178 6214 2212
rect 6214 2178 6248 2212
rect 6248 2178 6249 2212
rect 6069 2138 6249 2178
rect 6069 2104 6070 2138
rect 6070 2104 6104 2138
rect 6104 2104 6142 2138
rect 6142 2104 6176 2138
rect 6176 2104 6214 2138
rect 6214 2104 6248 2138
rect 6248 2104 6249 2138
rect 6069 2064 6249 2104
rect 6069 2030 6070 2064
rect 6070 2030 6104 2064
rect 6104 2030 6142 2064
rect 6142 2030 6176 2064
rect 6176 2030 6214 2064
rect 6214 2030 6248 2064
rect 6248 2030 6249 2064
rect 6069 1990 6249 2030
rect 6069 1956 6070 1990
rect 6070 1956 6104 1990
rect 6104 1956 6142 1990
rect 6142 1956 6176 1990
rect 6176 1956 6214 1990
rect 6214 1956 6248 1990
rect 6248 1956 6249 1990
rect 6069 1916 6249 1956
rect 6069 1882 6070 1916
rect 6070 1882 6104 1916
rect 6104 1882 6142 1916
rect 6142 1882 6176 1916
rect 6176 1882 6214 1916
rect 6214 1882 6248 1916
rect 6248 1882 6249 1916
rect 6069 1842 6249 1882
rect 6069 1808 6070 1842
rect 6070 1808 6104 1842
rect 6104 1808 6142 1842
rect 6142 1808 6176 1842
rect 6176 1808 6214 1842
rect 6214 1808 6248 1842
rect 6248 1808 6249 1842
rect 6069 1768 6249 1808
rect 6069 1734 6070 1768
rect 6070 1734 6104 1768
rect 6104 1734 6142 1768
rect 6142 1734 6176 1768
rect 6176 1734 6214 1768
rect 6214 1734 6248 1768
rect 6248 1734 6249 1768
rect 6069 1694 6249 1734
rect 6069 1660 6070 1694
rect 6070 1660 6104 1694
rect 6104 1660 6142 1694
rect 6142 1660 6176 1694
rect 6176 1660 6214 1694
rect 6214 1660 6248 1694
rect 6248 1660 6249 1694
rect 6069 1620 6249 1660
rect 6069 1586 6070 1620
rect 6070 1586 6104 1620
rect 6104 1586 6142 1620
rect 6142 1586 6176 1620
rect 6176 1586 6214 1620
rect 6214 1586 6248 1620
rect 6248 1586 6249 1620
rect 6069 1545 6249 1586
rect 6069 1538 6070 1545
rect 6070 1538 6104 1545
rect 6104 1538 6142 1545
rect 6142 1538 6176 1545
rect 6176 1538 6214 1545
rect 6214 1538 6248 1545
rect 6248 1538 6249 1545
rect 6069 1511 6070 1525
rect 6070 1511 6104 1525
rect 6104 1511 6121 1525
rect 6069 1473 6121 1511
rect 6133 1511 6142 1525
rect 6142 1511 6176 1525
rect 6176 1511 6185 1525
rect 6133 1473 6185 1511
rect 6197 1511 6214 1525
rect 6214 1511 6248 1525
rect 6248 1511 6249 1525
rect 6197 1473 6249 1511
rect 6565 4062 6745 4068
rect 6565 4050 6638 4062
rect 6638 4050 6672 4062
rect 6672 4050 6745 4062
rect 6565 3080 6566 4050
rect 6566 3092 6744 4050
rect 6566 3080 6600 3092
rect 6600 3080 6710 3092
rect 6710 3080 6744 3092
rect 6744 3080 6745 4050
rect 6565 3040 6745 3080
rect 6565 2992 6566 3040
rect 6566 2992 6744 3040
rect 6744 2992 6745 3040
rect 6565 2927 6566 2979
rect 6566 2927 6617 2979
rect 6629 2927 6681 2979
rect 6693 2927 6744 2979
rect 6744 2927 6745 2979
rect 7061 2582 7241 2614
rect 7061 2548 7062 2582
rect 7062 2548 7096 2582
rect 7096 2548 7134 2582
rect 7134 2548 7168 2582
rect 7168 2548 7206 2582
rect 7206 2548 7240 2582
rect 7240 2548 7241 2582
rect 7061 2508 7241 2548
rect 7061 2474 7062 2508
rect 7062 2474 7096 2508
rect 7096 2474 7134 2508
rect 7134 2474 7168 2508
rect 7168 2474 7206 2508
rect 7206 2474 7240 2508
rect 7240 2474 7241 2508
rect 7061 2434 7241 2474
rect 7061 2400 7062 2434
rect 7062 2400 7096 2434
rect 7096 2400 7134 2434
rect 7134 2400 7168 2434
rect 7168 2400 7206 2434
rect 7206 2400 7240 2434
rect 7240 2400 7241 2434
rect 7061 2360 7241 2400
rect 7061 2326 7062 2360
rect 7062 2326 7096 2360
rect 7096 2326 7134 2360
rect 7134 2326 7168 2360
rect 7168 2326 7206 2360
rect 7206 2326 7240 2360
rect 7240 2326 7241 2360
rect 7061 2286 7241 2326
rect 7061 2252 7062 2286
rect 7062 2252 7096 2286
rect 7096 2252 7134 2286
rect 7134 2252 7168 2286
rect 7168 2252 7206 2286
rect 7206 2252 7240 2286
rect 7240 2252 7241 2286
rect 7061 2212 7241 2252
rect 7061 2178 7062 2212
rect 7062 2178 7096 2212
rect 7096 2178 7134 2212
rect 7134 2178 7168 2212
rect 7168 2178 7206 2212
rect 7206 2178 7240 2212
rect 7240 2178 7241 2212
rect 7061 2138 7241 2178
rect 7061 2104 7062 2138
rect 7062 2104 7096 2138
rect 7096 2104 7134 2138
rect 7134 2104 7168 2138
rect 7168 2104 7206 2138
rect 7206 2104 7240 2138
rect 7240 2104 7241 2138
rect 7061 2064 7241 2104
rect 7061 2030 7062 2064
rect 7062 2030 7096 2064
rect 7096 2030 7134 2064
rect 7134 2030 7168 2064
rect 7168 2030 7206 2064
rect 7206 2030 7240 2064
rect 7240 2030 7241 2064
rect 7061 1990 7241 2030
rect 7061 1956 7062 1990
rect 7062 1956 7096 1990
rect 7096 1956 7134 1990
rect 7134 1956 7168 1990
rect 7168 1956 7206 1990
rect 7206 1956 7240 1990
rect 7240 1956 7241 1990
rect 7061 1916 7241 1956
rect 7061 1882 7062 1916
rect 7062 1882 7096 1916
rect 7096 1882 7134 1916
rect 7134 1882 7168 1916
rect 7168 1882 7206 1916
rect 7206 1882 7240 1916
rect 7240 1882 7241 1916
rect 7061 1842 7241 1882
rect 7061 1808 7062 1842
rect 7062 1808 7096 1842
rect 7096 1808 7134 1842
rect 7134 1808 7168 1842
rect 7168 1808 7206 1842
rect 7206 1808 7240 1842
rect 7240 1808 7241 1842
rect 7061 1768 7241 1808
rect 7061 1734 7062 1768
rect 7062 1734 7096 1768
rect 7096 1734 7134 1768
rect 7134 1734 7168 1768
rect 7168 1734 7206 1768
rect 7206 1734 7240 1768
rect 7240 1734 7241 1768
rect 7061 1694 7241 1734
rect 7061 1660 7062 1694
rect 7062 1660 7096 1694
rect 7096 1660 7134 1694
rect 7134 1660 7168 1694
rect 7168 1660 7206 1694
rect 7206 1660 7240 1694
rect 7240 1660 7241 1694
rect 7061 1620 7241 1660
rect 7061 1586 7062 1620
rect 7062 1586 7096 1620
rect 7096 1586 7134 1620
rect 7134 1586 7168 1620
rect 7168 1586 7206 1620
rect 7206 1586 7240 1620
rect 7240 1586 7241 1620
rect 7061 1545 7241 1586
rect 7061 1538 7062 1545
rect 7062 1538 7096 1545
rect 7096 1538 7134 1545
rect 7134 1538 7168 1545
rect 7168 1538 7206 1545
rect 7206 1538 7240 1545
rect 7240 1538 7241 1545
rect 7061 1511 7062 1525
rect 7062 1511 7096 1525
rect 7096 1511 7113 1525
rect 7061 1473 7113 1511
rect 7125 1511 7134 1525
rect 7134 1511 7168 1525
rect 7168 1511 7177 1525
rect 7125 1473 7177 1511
rect 7189 1511 7206 1525
rect 7206 1511 7240 1525
rect 7240 1511 7241 1525
rect 7189 1473 7241 1511
rect 7557 4062 7737 4068
rect 7557 4050 7630 4062
rect 7630 4050 7664 4062
rect 7664 4050 7737 4062
rect 7557 3080 7558 4050
rect 7558 3092 7736 4050
rect 7558 3080 7592 3092
rect 7592 3080 7702 3092
rect 7702 3080 7736 3092
rect 7736 3080 7737 4050
rect 7557 3040 7737 3080
rect 7557 2992 7558 3040
rect 7558 2992 7736 3040
rect 7736 2992 7737 3040
rect 7557 2927 7558 2979
rect 7558 2927 7609 2979
rect 7621 2927 7673 2979
rect 7685 2927 7736 2979
rect 7736 2927 7737 2979
rect 8053 2582 8233 2614
rect 8053 2548 8054 2582
rect 8054 2548 8088 2582
rect 8088 2548 8126 2582
rect 8126 2548 8160 2582
rect 8160 2548 8198 2582
rect 8198 2548 8232 2582
rect 8232 2548 8233 2582
rect 8053 2508 8233 2548
rect 8053 2474 8054 2508
rect 8054 2474 8088 2508
rect 8088 2474 8126 2508
rect 8126 2474 8160 2508
rect 8160 2474 8198 2508
rect 8198 2474 8232 2508
rect 8232 2474 8233 2508
rect 8053 2434 8233 2474
rect 8053 2400 8054 2434
rect 8054 2400 8088 2434
rect 8088 2400 8126 2434
rect 8126 2400 8160 2434
rect 8160 2400 8198 2434
rect 8198 2400 8232 2434
rect 8232 2400 8233 2434
rect 8053 2360 8233 2400
rect 8053 2326 8054 2360
rect 8054 2326 8088 2360
rect 8088 2326 8126 2360
rect 8126 2326 8160 2360
rect 8160 2326 8198 2360
rect 8198 2326 8232 2360
rect 8232 2326 8233 2360
rect 8053 2286 8233 2326
rect 8053 2252 8054 2286
rect 8054 2252 8088 2286
rect 8088 2252 8126 2286
rect 8126 2252 8160 2286
rect 8160 2252 8198 2286
rect 8198 2252 8232 2286
rect 8232 2252 8233 2286
rect 8053 2212 8233 2252
rect 8053 2178 8054 2212
rect 8054 2178 8088 2212
rect 8088 2178 8126 2212
rect 8126 2178 8160 2212
rect 8160 2178 8198 2212
rect 8198 2178 8232 2212
rect 8232 2178 8233 2212
rect 8053 2138 8233 2178
rect 8053 2104 8054 2138
rect 8054 2104 8088 2138
rect 8088 2104 8126 2138
rect 8126 2104 8160 2138
rect 8160 2104 8198 2138
rect 8198 2104 8232 2138
rect 8232 2104 8233 2138
rect 8053 2064 8233 2104
rect 8053 2030 8054 2064
rect 8054 2030 8088 2064
rect 8088 2030 8126 2064
rect 8126 2030 8160 2064
rect 8160 2030 8198 2064
rect 8198 2030 8232 2064
rect 8232 2030 8233 2064
rect 8053 1990 8233 2030
rect 8053 1956 8054 1990
rect 8054 1956 8088 1990
rect 8088 1956 8126 1990
rect 8126 1956 8160 1990
rect 8160 1956 8198 1990
rect 8198 1956 8232 1990
rect 8232 1956 8233 1990
rect 8053 1916 8233 1956
rect 8053 1882 8054 1916
rect 8054 1882 8088 1916
rect 8088 1882 8126 1916
rect 8126 1882 8160 1916
rect 8160 1882 8198 1916
rect 8198 1882 8232 1916
rect 8232 1882 8233 1916
rect 8053 1842 8233 1882
rect 8053 1808 8054 1842
rect 8054 1808 8088 1842
rect 8088 1808 8126 1842
rect 8126 1808 8160 1842
rect 8160 1808 8198 1842
rect 8198 1808 8232 1842
rect 8232 1808 8233 1842
rect 8053 1768 8233 1808
rect 8053 1734 8054 1768
rect 8054 1734 8088 1768
rect 8088 1734 8126 1768
rect 8126 1734 8160 1768
rect 8160 1734 8198 1768
rect 8198 1734 8232 1768
rect 8232 1734 8233 1768
rect 8053 1694 8233 1734
rect 8053 1660 8054 1694
rect 8054 1660 8088 1694
rect 8088 1660 8126 1694
rect 8126 1660 8160 1694
rect 8160 1660 8198 1694
rect 8198 1660 8232 1694
rect 8232 1660 8233 1694
rect 8053 1620 8233 1660
rect 8053 1586 8054 1620
rect 8054 1586 8088 1620
rect 8088 1586 8126 1620
rect 8126 1586 8160 1620
rect 8160 1586 8198 1620
rect 8198 1586 8232 1620
rect 8232 1586 8233 1620
rect 8053 1545 8233 1586
rect 8053 1538 8054 1545
rect 8054 1538 8088 1545
rect 8088 1538 8126 1545
rect 8126 1538 8160 1545
rect 8160 1538 8198 1545
rect 8198 1538 8232 1545
rect 8232 1538 8233 1545
rect 8053 1511 8054 1525
rect 8054 1511 8088 1525
rect 8088 1511 8105 1525
rect 8053 1473 8105 1511
rect 8117 1511 8126 1525
rect 8126 1511 8160 1525
rect 8160 1511 8169 1525
rect 8117 1473 8169 1511
rect 8181 1511 8198 1525
rect 8198 1511 8232 1525
rect 8232 1511 8233 1525
rect 8181 1473 8233 1511
rect 8549 4062 8729 4068
rect 8549 4050 8622 4062
rect 8622 4050 8656 4062
rect 8656 4050 8729 4062
rect 8549 3080 8550 4050
rect 8550 3092 8728 4050
rect 8550 3080 8584 3092
rect 8584 3080 8694 3092
rect 8694 3080 8728 3092
rect 8728 3080 8729 4050
rect 8549 3040 8729 3080
rect 8549 2992 8550 3040
rect 8550 2992 8728 3040
rect 8728 2992 8729 3040
rect 8549 2927 8550 2979
rect 8550 2927 8601 2979
rect 8613 2927 8665 2979
rect 8677 2927 8728 2979
rect 8728 2927 8729 2979
rect 9045 2582 9225 2614
rect 9045 2548 9046 2582
rect 9046 2548 9080 2582
rect 9080 2548 9118 2582
rect 9118 2548 9152 2582
rect 9152 2548 9190 2582
rect 9190 2548 9224 2582
rect 9224 2548 9225 2582
rect 9045 2508 9225 2548
rect 9045 2474 9046 2508
rect 9046 2474 9080 2508
rect 9080 2474 9118 2508
rect 9118 2474 9152 2508
rect 9152 2474 9190 2508
rect 9190 2474 9224 2508
rect 9224 2474 9225 2508
rect 9045 2434 9225 2474
rect 9045 2400 9046 2434
rect 9046 2400 9080 2434
rect 9080 2400 9118 2434
rect 9118 2400 9152 2434
rect 9152 2400 9190 2434
rect 9190 2400 9224 2434
rect 9224 2400 9225 2434
rect 9045 2360 9225 2400
rect 9045 2326 9046 2360
rect 9046 2326 9080 2360
rect 9080 2326 9118 2360
rect 9118 2326 9152 2360
rect 9152 2326 9190 2360
rect 9190 2326 9224 2360
rect 9224 2326 9225 2360
rect 9045 2286 9225 2326
rect 9045 2252 9046 2286
rect 9046 2252 9080 2286
rect 9080 2252 9118 2286
rect 9118 2252 9152 2286
rect 9152 2252 9190 2286
rect 9190 2252 9224 2286
rect 9224 2252 9225 2286
rect 9045 2212 9225 2252
rect 9045 2178 9046 2212
rect 9046 2178 9080 2212
rect 9080 2178 9118 2212
rect 9118 2178 9152 2212
rect 9152 2178 9190 2212
rect 9190 2178 9224 2212
rect 9224 2178 9225 2212
rect 9045 2138 9225 2178
rect 9045 2104 9046 2138
rect 9046 2104 9080 2138
rect 9080 2104 9118 2138
rect 9118 2104 9152 2138
rect 9152 2104 9190 2138
rect 9190 2104 9224 2138
rect 9224 2104 9225 2138
rect 9045 2064 9225 2104
rect 9045 2030 9046 2064
rect 9046 2030 9080 2064
rect 9080 2030 9118 2064
rect 9118 2030 9152 2064
rect 9152 2030 9190 2064
rect 9190 2030 9224 2064
rect 9224 2030 9225 2064
rect 9045 1990 9225 2030
rect 9045 1956 9046 1990
rect 9046 1956 9080 1990
rect 9080 1956 9118 1990
rect 9118 1956 9152 1990
rect 9152 1956 9190 1990
rect 9190 1956 9224 1990
rect 9224 1956 9225 1990
rect 9045 1916 9225 1956
rect 9045 1882 9046 1916
rect 9046 1882 9080 1916
rect 9080 1882 9118 1916
rect 9118 1882 9152 1916
rect 9152 1882 9190 1916
rect 9190 1882 9224 1916
rect 9224 1882 9225 1916
rect 9045 1842 9225 1882
rect 9045 1808 9046 1842
rect 9046 1808 9080 1842
rect 9080 1808 9118 1842
rect 9118 1808 9152 1842
rect 9152 1808 9190 1842
rect 9190 1808 9224 1842
rect 9224 1808 9225 1842
rect 9045 1768 9225 1808
rect 9045 1734 9046 1768
rect 9046 1734 9080 1768
rect 9080 1734 9118 1768
rect 9118 1734 9152 1768
rect 9152 1734 9190 1768
rect 9190 1734 9224 1768
rect 9224 1734 9225 1768
rect 9045 1694 9225 1734
rect 9045 1660 9046 1694
rect 9046 1660 9080 1694
rect 9080 1660 9118 1694
rect 9118 1660 9152 1694
rect 9152 1660 9190 1694
rect 9190 1660 9224 1694
rect 9224 1660 9225 1694
rect 9045 1620 9225 1660
rect 9045 1586 9046 1620
rect 9046 1586 9080 1620
rect 9080 1586 9118 1620
rect 9118 1586 9152 1620
rect 9152 1586 9190 1620
rect 9190 1586 9224 1620
rect 9224 1586 9225 1620
rect 9045 1545 9225 1586
rect 9045 1538 9046 1545
rect 9046 1538 9080 1545
rect 9080 1538 9118 1545
rect 9118 1538 9152 1545
rect 9152 1538 9190 1545
rect 9190 1538 9224 1545
rect 9224 1538 9225 1545
rect 9045 1511 9046 1525
rect 9046 1511 9080 1525
rect 9080 1511 9097 1525
rect 9045 1473 9097 1511
rect 9109 1511 9118 1525
rect 9118 1511 9152 1525
rect 9152 1511 9161 1525
rect 9109 1473 9161 1511
rect 9173 1511 9190 1525
rect 9190 1511 9224 1525
rect 9224 1511 9225 1525
rect 9173 1473 9225 1511
rect 9541 4062 9721 4068
rect 9541 4050 9614 4062
rect 9614 4050 9648 4062
rect 9648 4050 9721 4062
rect 9541 3080 9542 4050
rect 9542 3092 9720 4050
rect 9542 3080 9576 3092
rect 9576 3080 9686 3092
rect 9686 3080 9720 3092
rect 9720 3080 9721 4050
rect 9541 3040 9721 3080
rect 9541 2992 9542 3040
rect 9542 2992 9720 3040
rect 9720 2992 9721 3040
rect 9541 2927 9542 2979
rect 9542 2927 9593 2979
rect 9605 2927 9657 2979
rect 9669 2927 9720 2979
rect 9720 2927 9721 2979
rect 10037 2582 10217 2614
rect 10037 2548 10038 2582
rect 10038 2548 10072 2582
rect 10072 2548 10110 2582
rect 10110 2548 10144 2582
rect 10144 2548 10182 2582
rect 10182 2548 10216 2582
rect 10216 2548 10217 2582
rect 10037 2508 10217 2548
rect 10037 2474 10038 2508
rect 10038 2474 10072 2508
rect 10072 2474 10110 2508
rect 10110 2474 10144 2508
rect 10144 2474 10182 2508
rect 10182 2474 10216 2508
rect 10216 2474 10217 2508
rect 10037 2434 10217 2474
rect 10037 2400 10038 2434
rect 10038 2400 10072 2434
rect 10072 2400 10110 2434
rect 10110 2400 10144 2434
rect 10144 2400 10182 2434
rect 10182 2400 10216 2434
rect 10216 2400 10217 2434
rect 10037 2360 10217 2400
rect 10037 2326 10038 2360
rect 10038 2326 10072 2360
rect 10072 2326 10110 2360
rect 10110 2326 10144 2360
rect 10144 2326 10182 2360
rect 10182 2326 10216 2360
rect 10216 2326 10217 2360
rect 10037 2286 10217 2326
rect 10037 2252 10038 2286
rect 10038 2252 10072 2286
rect 10072 2252 10110 2286
rect 10110 2252 10144 2286
rect 10144 2252 10182 2286
rect 10182 2252 10216 2286
rect 10216 2252 10217 2286
rect 10037 2212 10217 2252
rect 10037 2178 10038 2212
rect 10038 2178 10072 2212
rect 10072 2178 10110 2212
rect 10110 2178 10144 2212
rect 10144 2178 10182 2212
rect 10182 2178 10216 2212
rect 10216 2178 10217 2212
rect 10037 2138 10217 2178
rect 10037 2104 10038 2138
rect 10038 2104 10072 2138
rect 10072 2104 10110 2138
rect 10110 2104 10144 2138
rect 10144 2104 10182 2138
rect 10182 2104 10216 2138
rect 10216 2104 10217 2138
rect 10037 2064 10217 2104
rect 10037 2030 10038 2064
rect 10038 2030 10072 2064
rect 10072 2030 10110 2064
rect 10110 2030 10144 2064
rect 10144 2030 10182 2064
rect 10182 2030 10216 2064
rect 10216 2030 10217 2064
rect 10037 1990 10217 2030
rect 10037 1956 10038 1990
rect 10038 1956 10072 1990
rect 10072 1956 10110 1990
rect 10110 1956 10144 1990
rect 10144 1956 10182 1990
rect 10182 1956 10216 1990
rect 10216 1956 10217 1990
rect 10037 1916 10217 1956
rect 10037 1882 10038 1916
rect 10038 1882 10072 1916
rect 10072 1882 10110 1916
rect 10110 1882 10144 1916
rect 10144 1882 10182 1916
rect 10182 1882 10216 1916
rect 10216 1882 10217 1916
rect 10037 1842 10217 1882
rect 10037 1808 10038 1842
rect 10038 1808 10072 1842
rect 10072 1808 10110 1842
rect 10110 1808 10144 1842
rect 10144 1808 10182 1842
rect 10182 1808 10216 1842
rect 10216 1808 10217 1842
rect 10037 1768 10217 1808
rect 10037 1734 10038 1768
rect 10038 1734 10072 1768
rect 10072 1734 10110 1768
rect 10110 1734 10144 1768
rect 10144 1734 10182 1768
rect 10182 1734 10216 1768
rect 10216 1734 10217 1768
rect 10037 1694 10217 1734
rect 10037 1660 10038 1694
rect 10038 1660 10072 1694
rect 10072 1660 10110 1694
rect 10110 1660 10144 1694
rect 10144 1660 10182 1694
rect 10182 1660 10216 1694
rect 10216 1660 10217 1694
rect 10037 1620 10217 1660
rect 10037 1586 10038 1620
rect 10038 1586 10072 1620
rect 10072 1586 10110 1620
rect 10110 1586 10144 1620
rect 10144 1586 10182 1620
rect 10182 1586 10216 1620
rect 10216 1586 10217 1620
rect 10037 1545 10217 1586
rect 10037 1538 10038 1545
rect 10038 1538 10072 1545
rect 10072 1538 10110 1545
rect 10110 1538 10144 1545
rect 10144 1538 10182 1545
rect 10182 1538 10216 1545
rect 10216 1538 10217 1545
rect 10037 1511 10038 1525
rect 10038 1511 10072 1525
rect 10072 1511 10089 1525
rect 10037 1473 10089 1511
rect 10101 1511 10110 1525
rect 10110 1511 10144 1525
rect 10144 1511 10153 1525
rect 10101 1473 10153 1511
rect 10165 1511 10182 1525
rect 10182 1511 10216 1525
rect 10216 1511 10217 1525
rect 10165 1473 10217 1511
rect 10533 4062 10713 4068
rect 10533 4050 10606 4062
rect 10606 4050 10640 4062
rect 10640 4050 10713 4062
rect 10533 3080 10534 4050
rect 10534 3092 10712 4050
rect 10534 3080 10568 3092
rect 10568 3080 10678 3092
rect 10678 3080 10712 3092
rect 10712 3080 10713 4050
rect 10533 3037 10713 3080
rect 10533 3003 10534 3037
rect 10534 3003 10568 3037
rect 10568 3003 10606 3037
rect 10606 3003 10640 3037
rect 10640 3003 10678 3037
rect 10678 3003 10712 3037
rect 10712 3003 10713 3037
rect 10533 2992 10713 3003
rect 10533 2954 10585 2979
rect 10533 2927 10534 2954
rect 10534 2927 10568 2954
rect 10568 2927 10585 2954
rect 10597 2954 10649 2979
rect 10597 2927 10606 2954
rect 10606 2927 10640 2954
rect 10640 2927 10649 2954
rect 10661 2954 10713 2979
rect 10661 2927 10678 2954
rect 10678 2927 10712 2954
rect 10712 2927 10713 2954
rect 11029 2582 11209 2614
rect 11029 2548 11030 2582
rect 11030 2548 11064 2582
rect 11064 2548 11102 2582
rect 11102 2548 11136 2582
rect 11136 2548 11174 2582
rect 11174 2548 11208 2582
rect 11208 2548 11209 2582
rect 11029 2508 11209 2548
rect 11029 2474 11030 2508
rect 11030 2474 11064 2508
rect 11064 2474 11102 2508
rect 11102 2474 11136 2508
rect 11136 2474 11174 2508
rect 11174 2474 11208 2508
rect 11208 2474 11209 2508
rect 11029 2434 11209 2474
rect 11029 2400 11030 2434
rect 11030 2400 11064 2434
rect 11064 2400 11102 2434
rect 11102 2400 11136 2434
rect 11136 2400 11174 2434
rect 11174 2400 11208 2434
rect 11208 2400 11209 2434
rect 11029 2360 11209 2400
rect 11029 2326 11030 2360
rect 11030 2326 11064 2360
rect 11064 2326 11102 2360
rect 11102 2326 11136 2360
rect 11136 2326 11174 2360
rect 11174 2326 11208 2360
rect 11208 2326 11209 2360
rect 11029 2286 11209 2326
rect 11029 2252 11030 2286
rect 11030 2252 11064 2286
rect 11064 2252 11102 2286
rect 11102 2252 11136 2286
rect 11136 2252 11174 2286
rect 11174 2252 11208 2286
rect 11208 2252 11209 2286
rect 11029 2212 11209 2252
rect 11029 2178 11030 2212
rect 11030 2178 11064 2212
rect 11064 2178 11102 2212
rect 11102 2178 11136 2212
rect 11136 2178 11174 2212
rect 11174 2178 11208 2212
rect 11208 2178 11209 2212
rect 11029 2138 11209 2178
rect 11029 2104 11030 2138
rect 11030 2104 11064 2138
rect 11064 2104 11102 2138
rect 11102 2104 11136 2138
rect 11136 2104 11174 2138
rect 11174 2104 11208 2138
rect 11208 2104 11209 2138
rect 11029 2064 11209 2104
rect 11029 2030 11030 2064
rect 11030 2030 11064 2064
rect 11064 2030 11102 2064
rect 11102 2030 11136 2064
rect 11136 2030 11174 2064
rect 11174 2030 11208 2064
rect 11208 2030 11209 2064
rect 11029 1990 11209 2030
rect 11029 1956 11030 1990
rect 11030 1956 11064 1990
rect 11064 1956 11102 1990
rect 11102 1956 11136 1990
rect 11136 1956 11174 1990
rect 11174 1956 11208 1990
rect 11208 1956 11209 1990
rect 11029 1916 11209 1956
rect 11029 1882 11030 1916
rect 11030 1882 11064 1916
rect 11064 1882 11102 1916
rect 11102 1882 11136 1916
rect 11136 1882 11174 1916
rect 11174 1882 11208 1916
rect 11208 1882 11209 1916
rect 11029 1842 11209 1882
rect 11029 1808 11030 1842
rect 11030 1808 11064 1842
rect 11064 1808 11102 1842
rect 11102 1808 11136 1842
rect 11136 1808 11174 1842
rect 11174 1808 11208 1842
rect 11208 1808 11209 1842
rect 11029 1768 11209 1808
rect 11029 1734 11030 1768
rect 11030 1734 11064 1768
rect 11064 1734 11102 1768
rect 11102 1734 11136 1768
rect 11136 1734 11174 1768
rect 11174 1734 11208 1768
rect 11208 1734 11209 1768
rect 11029 1694 11209 1734
rect 11029 1660 11030 1694
rect 11030 1660 11064 1694
rect 11064 1660 11102 1694
rect 11102 1660 11136 1694
rect 11136 1660 11174 1694
rect 11174 1660 11208 1694
rect 11208 1660 11209 1694
rect 11029 1620 11209 1660
rect 11029 1586 11030 1620
rect 11030 1586 11064 1620
rect 11064 1586 11102 1620
rect 11102 1586 11136 1620
rect 11136 1586 11174 1620
rect 11174 1586 11208 1620
rect 11208 1586 11209 1620
rect 11029 1545 11209 1586
rect 11029 1538 11030 1545
rect 11030 1538 11064 1545
rect 11064 1538 11102 1545
rect 11102 1538 11136 1545
rect 11136 1538 11174 1545
rect 11174 1538 11208 1545
rect 11208 1538 11209 1545
rect 11029 1511 11030 1525
rect 11030 1511 11064 1525
rect 11064 1511 11081 1525
rect 11029 1473 11081 1511
rect 11093 1511 11102 1525
rect 11102 1511 11136 1525
rect 11136 1511 11145 1525
rect 11093 1473 11145 1511
rect 11157 1511 11174 1525
rect 11174 1511 11208 1525
rect 11208 1511 11209 1525
rect 11157 1473 11209 1511
rect 11525 4062 11705 4068
rect 11525 4050 11598 4062
rect 11598 4050 11632 4062
rect 11632 4050 11705 4062
rect 11525 3080 11526 4050
rect 11526 3092 11704 4050
rect 11526 3080 11560 3092
rect 11560 3080 11670 3092
rect 11670 3080 11704 3092
rect 11704 3080 11705 4050
rect 11525 3037 11705 3080
rect 11525 3003 11526 3037
rect 11526 3003 11560 3037
rect 11560 3003 11598 3037
rect 11598 3003 11632 3037
rect 11632 3003 11670 3037
rect 11670 3003 11704 3037
rect 11704 3003 11705 3037
rect 11525 2992 11705 3003
rect 11525 2954 11577 2979
rect 11525 2927 11526 2954
rect 11526 2927 11560 2954
rect 11560 2927 11577 2954
rect 11589 2954 11641 2979
rect 11589 2927 11598 2954
rect 11598 2927 11632 2954
rect 11632 2927 11641 2954
rect 11653 2954 11705 2979
rect 11653 2927 11670 2954
rect 11670 2927 11704 2954
rect 11704 2927 11705 2954
rect 12021 2582 12201 2614
rect 12021 2548 12022 2582
rect 12022 2548 12056 2582
rect 12056 2548 12094 2582
rect 12094 2548 12128 2582
rect 12128 2548 12166 2582
rect 12166 2548 12200 2582
rect 12200 2548 12201 2582
rect 12021 2508 12201 2548
rect 12021 2474 12022 2508
rect 12022 2474 12056 2508
rect 12056 2474 12094 2508
rect 12094 2474 12128 2508
rect 12128 2474 12166 2508
rect 12166 2474 12200 2508
rect 12200 2474 12201 2508
rect 12021 2434 12201 2474
rect 12021 2400 12022 2434
rect 12022 2400 12056 2434
rect 12056 2400 12094 2434
rect 12094 2400 12128 2434
rect 12128 2400 12166 2434
rect 12166 2400 12200 2434
rect 12200 2400 12201 2434
rect 12021 2360 12201 2400
rect 12021 2326 12022 2360
rect 12022 2326 12056 2360
rect 12056 2326 12094 2360
rect 12094 2326 12128 2360
rect 12128 2326 12166 2360
rect 12166 2326 12200 2360
rect 12200 2326 12201 2360
rect 12021 2286 12201 2326
rect 12021 2252 12022 2286
rect 12022 2252 12056 2286
rect 12056 2252 12094 2286
rect 12094 2252 12128 2286
rect 12128 2252 12166 2286
rect 12166 2252 12200 2286
rect 12200 2252 12201 2286
rect 12021 2212 12201 2252
rect 12021 2178 12022 2212
rect 12022 2178 12056 2212
rect 12056 2178 12094 2212
rect 12094 2178 12128 2212
rect 12128 2178 12166 2212
rect 12166 2178 12200 2212
rect 12200 2178 12201 2212
rect 12021 2138 12201 2178
rect 12021 2104 12022 2138
rect 12022 2104 12056 2138
rect 12056 2104 12094 2138
rect 12094 2104 12128 2138
rect 12128 2104 12166 2138
rect 12166 2104 12200 2138
rect 12200 2104 12201 2138
rect 12021 2064 12201 2104
rect 12021 2030 12022 2064
rect 12022 2030 12056 2064
rect 12056 2030 12094 2064
rect 12094 2030 12128 2064
rect 12128 2030 12166 2064
rect 12166 2030 12200 2064
rect 12200 2030 12201 2064
rect 12021 1990 12201 2030
rect 12021 1956 12022 1990
rect 12022 1956 12056 1990
rect 12056 1956 12094 1990
rect 12094 1956 12128 1990
rect 12128 1956 12166 1990
rect 12166 1956 12200 1990
rect 12200 1956 12201 1990
rect 12021 1916 12201 1956
rect 12021 1882 12022 1916
rect 12022 1882 12056 1916
rect 12056 1882 12094 1916
rect 12094 1882 12128 1916
rect 12128 1882 12166 1916
rect 12166 1882 12200 1916
rect 12200 1882 12201 1916
rect 12021 1842 12201 1882
rect 12021 1808 12022 1842
rect 12022 1808 12056 1842
rect 12056 1808 12094 1842
rect 12094 1808 12128 1842
rect 12128 1808 12166 1842
rect 12166 1808 12200 1842
rect 12200 1808 12201 1842
rect 12021 1768 12201 1808
rect 12021 1734 12022 1768
rect 12022 1734 12056 1768
rect 12056 1734 12094 1768
rect 12094 1734 12128 1768
rect 12128 1734 12166 1768
rect 12166 1734 12200 1768
rect 12200 1734 12201 1768
rect 12021 1694 12201 1734
rect 12021 1660 12022 1694
rect 12022 1660 12056 1694
rect 12056 1660 12094 1694
rect 12094 1660 12128 1694
rect 12128 1660 12166 1694
rect 12166 1660 12200 1694
rect 12200 1660 12201 1694
rect 12021 1620 12201 1660
rect 12021 1586 12022 1620
rect 12022 1586 12056 1620
rect 12056 1586 12094 1620
rect 12094 1586 12128 1620
rect 12128 1586 12166 1620
rect 12166 1586 12200 1620
rect 12200 1586 12201 1620
rect 12021 1545 12201 1586
rect 12021 1538 12022 1545
rect 12022 1538 12056 1545
rect 12056 1538 12094 1545
rect 12094 1538 12128 1545
rect 12128 1538 12166 1545
rect 12166 1538 12200 1545
rect 12200 1538 12201 1545
rect 12021 1511 12022 1525
rect 12022 1511 12056 1525
rect 12056 1511 12073 1525
rect 12021 1473 12073 1511
rect 12085 1511 12094 1525
rect 12094 1511 12128 1525
rect 12128 1511 12137 1525
rect 12085 1473 12137 1511
rect 12149 1511 12166 1525
rect 12166 1511 12200 1525
rect 12200 1511 12201 1525
rect 12149 1473 12201 1511
rect 12517 4062 12697 4068
rect 12517 4050 12590 4062
rect 12590 4050 12624 4062
rect 12624 4050 12697 4062
rect 12517 3080 12518 4050
rect 12518 3092 12696 4050
rect 12518 3080 12552 3092
rect 12552 3080 12662 3092
rect 12662 3080 12696 3092
rect 12696 3080 12697 4050
rect 12517 3038 12697 3080
rect 12517 3004 12518 3038
rect 12518 3004 12552 3038
rect 12552 3004 12590 3038
rect 12590 3004 12624 3038
rect 12624 3004 12662 3038
rect 12662 3004 12696 3038
rect 12696 3004 12697 3038
rect 12517 2992 12697 3004
rect 12517 2955 12569 2979
rect 12517 2927 12518 2955
rect 12518 2927 12552 2955
rect 12552 2927 12569 2955
rect 12581 2955 12633 2979
rect 12581 2927 12590 2955
rect 12590 2927 12624 2955
rect 12624 2927 12633 2955
rect 12645 2955 12697 2979
rect 12645 2927 12662 2955
rect 12662 2927 12696 2955
rect 12696 2927 12697 2955
rect 13013 2582 13193 2614
rect 13013 2548 13014 2582
rect 13014 2548 13048 2582
rect 13048 2548 13086 2582
rect 13086 2548 13120 2582
rect 13120 2548 13158 2582
rect 13158 2548 13192 2582
rect 13192 2548 13193 2582
rect 13013 2508 13193 2548
rect 13013 2474 13014 2508
rect 13014 2474 13048 2508
rect 13048 2474 13086 2508
rect 13086 2474 13120 2508
rect 13120 2474 13158 2508
rect 13158 2474 13192 2508
rect 13192 2474 13193 2508
rect 13013 2434 13193 2474
rect 13013 2400 13014 2434
rect 13014 2400 13048 2434
rect 13048 2400 13086 2434
rect 13086 2400 13120 2434
rect 13120 2400 13158 2434
rect 13158 2400 13192 2434
rect 13192 2400 13193 2434
rect 13013 2360 13193 2400
rect 13013 2326 13014 2360
rect 13014 2326 13048 2360
rect 13048 2326 13086 2360
rect 13086 2326 13120 2360
rect 13120 2326 13158 2360
rect 13158 2326 13192 2360
rect 13192 2326 13193 2360
rect 13013 2286 13193 2326
rect 13013 2252 13014 2286
rect 13014 2252 13048 2286
rect 13048 2252 13086 2286
rect 13086 2252 13120 2286
rect 13120 2252 13158 2286
rect 13158 2252 13192 2286
rect 13192 2252 13193 2286
rect 13013 2212 13193 2252
rect 13013 2178 13014 2212
rect 13014 2178 13048 2212
rect 13048 2178 13086 2212
rect 13086 2178 13120 2212
rect 13120 2178 13158 2212
rect 13158 2178 13192 2212
rect 13192 2178 13193 2212
rect 13013 2138 13193 2178
rect 13013 2104 13014 2138
rect 13014 2104 13048 2138
rect 13048 2104 13086 2138
rect 13086 2104 13120 2138
rect 13120 2104 13158 2138
rect 13158 2104 13192 2138
rect 13192 2104 13193 2138
rect 13013 2064 13193 2104
rect 13013 2030 13014 2064
rect 13014 2030 13048 2064
rect 13048 2030 13086 2064
rect 13086 2030 13120 2064
rect 13120 2030 13158 2064
rect 13158 2030 13192 2064
rect 13192 2030 13193 2064
rect 13013 1990 13193 2030
rect 13013 1956 13014 1990
rect 13014 1956 13048 1990
rect 13048 1956 13086 1990
rect 13086 1956 13120 1990
rect 13120 1956 13158 1990
rect 13158 1956 13192 1990
rect 13192 1956 13193 1990
rect 13013 1916 13193 1956
rect 13013 1882 13014 1916
rect 13014 1882 13048 1916
rect 13048 1882 13086 1916
rect 13086 1882 13120 1916
rect 13120 1882 13158 1916
rect 13158 1882 13192 1916
rect 13192 1882 13193 1916
rect 13013 1842 13193 1882
rect 13013 1808 13014 1842
rect 13014 1808 13048 1842
rect 13048 1808 13086 1842
rect 13086 1808 13120 1842
rect 13120 1808 13158 1842
rect 13158 1808 13192 1842
rect 13192 1808 13193 1842
rect 13013 1768 13193 1808
rect 13013 1734 13014 1768
rect 13014 1734 13048 1768
rect 13048 1734 13086 1768
rect 13086 1734 13120 1768
rect 13120 1734 13158 1768
rect 13158 1734 13192 1768
rect 13192 1734 13193 1768
rect 13013 1694 13193 1734
rect 13013 1660 13014 1694
rect 13014 1660 13048 1694
rect 13048 1660 13086 1694
rect 13086 1660 13120 1694
rect 13120 1660 13158 1694
rect 13158 1660 13192 1694
rect 13192 1660 13193 1694
rect 13013 1620 13193 1660
rect 13013 1586 13014 1620
rect 13014 1586 13048 1620
rect 13048 1586 13086 1620
rect 13086 1586 13120 1620
rect 13120 1586 13158 1620
rect 13158 1586 13192 1620
rect 13192 1586 13193 1620
rect 13013 1545 13193 1586
rect 13013 1538 13014 1545
rect 13014 1538 13048 1545
rect 13048 1538 13086 1545
rect 13086 1538 13120 1545
rect 13120 1538 13158 1545
rect 13158 1538 13192 1545
rect 13192 1538 13193 1545
rect 13013 1511 13014 1525
rect 13014 1511 13048 1525
rect 13048 1511 13065 1525
rect 13013 1473 13065 1511
rect 13077 1511 13086 1525
rect 13086 1511 13120 1525
rect 13120 1511 13129 1525
rect 13077 1473 13129 1511
rect 13141 1511 13158 1525
rect 13158 1511 13192 1525
rect 13192 1511 13193 1525
rect 13141 1473 13193 1511
rect 13509 4062 13689 4068
rect 13509 4050 13582 4062
rect 13582 4050 13616 4062
rect 13616 4050 13689 4062
rect 13509 3080 13510 4050
rect 13510 3092 13688 4050
rect 13510 3080 13544 3092
rect 13544 3080 13654 3092
rect 13654 3080 13688 3092
rect 13688 3080 13689 4050
rect 13509 3040 13689 3080
rect 13509 2992 13510 3040
rect 13510 2992 13688 3040
rect 13688 2992 13689 3040
rect 13509 2927 13510 2979
rect 13510 2927 13561 2979
rect 13573 2927 13625 2979
rect 13637 2927 13688 2979
rect 13688 2927 13689 2979
rect 14037 2586 14042 2614
rect 14042 2586 14076 2614
rect 14076 2586 14089 2614
rect 14037 2562 14089 2586
rect 14105 2562 14157 2614
rect 14173 2562 14225 2614
rect 14037 2547 14089 2550
rect 14037 2513 14042 2547
rect 14042 2513 14076 2547
rect 14076 2513 14089 2547
rect 14037 2498 14089 2513
rect 14105 2498 14157 2550
rect 14173 2498 14225 2550
rect 14037 2474 14089 2486
rect 14037 2440 14042 2474
rect 14042 2440 14076 2474
rect 14076 2440 14089 2474
rect 14037 2434 14089 2440
rect 14105 2434 14157 2486
rect 14173 2434 14225 2486
rect 14037 2401 14089 2422
rect 14037 2370 14042 2401
rect 14042 2370 14076 2401
rect 14076 2370 14089 2401
rect 14105 2370 14157 2422
rect 14173 2370 14225 2422
rect 14037 2328 14089 2358
rect 14037 2306 14042 2328
rect 14042 2306 14076 2328
rect 14076 2306 14089 2328
rect 14105 2306 14157 2358
rect 14173 2306 14225 2358
rect 14037 2255 14089 2294
rect 14037 2242 14042 2255
rect 14042 2242 14076 2255
rect 14076 2242 14089 2255
rect 14105 2242 14157 2294
rect 14173 2242 14225 2294
rect 14037 2221 14042 2230
rect 14042 2221 14076 2230
rect 14076 2221 14089 2230
rect 14037 2182 14089 2221
rect 14037 2178 14042 2182
rect 14042 2178 14076 2182
rect 14076 2178 14089 2182
rect 14105 2178 14157 2230
rect 14173 2178 14225 2230
rect 14037 2148 14042 2166
rect 14042 2148 14076 2166
rect 14076 2148 14089 2166
rect 14037 2114 14089 2148
rect 14105 2114 14157 2166
rect 14173 2114 14225 2166
rect 14037 2075 14042 2102
rect 14042 2075 14076 2102
rect 14076 2075 14089 2102
rect 14037 2050 14089 2075
rect 14105 2050 14157 2102
rect 14173 2050 14225 2102
rect 14037 2036 14089 2038
rect 14037 2002 14042 2036
rect 14042 2002 14076 2036
rect 14076 2002 14089 2036
rect 14037 1986 14089 2002
rect 14105 1986 14157 2038
rect 14173 1986 14225 2038
rect 14037 1963 14089 1974
rect 14037 1929 14042 1963
rect 14042 1929 14076 1963
rect 14076 1929 14089 1963
rect 14037 1922 14089 1929
rect 14105 1922 14157 1974
rect 14173 1922 14225 1974
rect 14037 1890 14089 1910
rect 14037 1858 14042 1890
rect 14042 1858 14076 1890
rect 14076 1858 14089 1890
rect 14105 1858 14157 1910
rect 14173 1858 14225 1910
rect 14037 1817 14089 1846
rect 14037 1794 14042 1817
rect 14042 1794 14076 1817
rect 14076 1794 14089 1817
rect 14105 1794 14157 1846
rect 14173 1794 14225 1846
rect 14037 1744 14089 1782
rect 14037 1730 14042 1744
rect 14042 1730 14076 1744
rect 14076 1730 14089 1744
rect 14105 1730 14157 1782
rect 14173 1730 14225 1782
rect 14037 1710 14042 1718
rect 14042 1710 14076 1718
rect 14076 1710 14089 1718
rect 14037 1671 14089 1710
rect 14037 1666 14042 1671
rect 14042 1666 14076 1671
rect 14076 1666 14089 1671
rect 14105 1666 14157 1718
rect 14173 1666 14225 1718
rect 14037 1637 14042 1654
rect 14042 1637 14076 1654
rect 14076 1637 14089 1654
rect 14037 1602 14089 1637
rect 14105 1602 14157 1654
rect 14173 1602 14225 1654
rect 14037 1564 14042 1590
rect 14042 1564 14076 1590
rect 14076 1564 14089 1590
rect 14037 1538 14089 1564
rect 14105 1538 14157 1590
rect 14173 1538 14225 1590
rect 14037 1491 14042 1525
rect 14042 1491 14076 1525
rect 14076 1491 14089 1525
rect 14037 1473 14089 1491
rect 14105 1473 14157 1525
rect 14173 1473 14225 1525
rect 14400 4044 14452 4068
rect 14488 4052 14510 4068
rect 14510 4052 14540 4068
rect 14576 4052 14582 4068
rect 14582 4052 14616 4068
rect 14616 4052 14628 4068
rect 14400 4016 14431 4044
rect 14431 4016 14452 4044
rect 14488 4016 14540 4052
rect 14576 4016 14628 4052
rect 14400 3971 14452 4004
rect 14488 3979 14510 4004
rect 14510 3979 14540 4004
rect 14576 3979 14582 4004
rect 14582 3979 14616 4004
rect 14616 3979 14628 4004
rect 14400 3952 14431 3971
rect 14431 3952 14452 3971
rect 14488 3952 14540 3979
rect 14576 3952 14628 3979
rect 14400 3937 14431 3940
rect 14431 3937 14452 3940
rect 14400 3898 14452 3937
rect 14488 3906 14510 3940
rect 14510 3906 14540 3940
rect 14576 3906 14582 3940
rect 14582 3906 14616 3940
rect 14616 3906 14628 3940
rect 14400 3888 14431 3898
rect 14431 3888 14452 3898
rect 14488 3888 14540 3906
rect 14576 3888 14628 3906
rect 14400 3864 14431 3876
rect 14431 3864 14452 3876
rect 14488 3867 14540 3876
rect 14576 3867 14628 3876
rect 14400 3825 14452 3864
rect 14488 3833 14510 3867
rect 14510 3833 14540 3867
rect 14576 3833 14582 3867
rect 14582 3833 14616 3867
rect 14616 3833 14628 3867
rect 14400 3824 14431 3825
rect 14431 3824 14452 3825
rect 14488 3824 14540 3833
rect 14576 3824 14628 3833
rect 14400 3791 14431 3812
rect 14431 3791 14452 3812
rect 14488 3794 14540 3812
rect 14576 3794 14628 3812
rect 14400 3760 14452 3791
rect 14488 3760 14510 3794
rect 14510 3760 14540 3794
rect 14576 3760 14582 3794
rect 14582 3760 14616 3794
rect 14616 3760 14628 3794
rect 14400 3718 14431 3748
rect 14431 3718 14452 3748
rect 14488 3721 14540 3748
rect 14576 3721 14628 3748
rect 14400 3696 14452 3718
rect 14488 3696 14510 3721
rect 14510 3696 14540 3721
rect 14576 3696 14582 3721
rect 14582 3696 14616 3721
rect 14616 3696 14628 3721
rect 14400 3679 14452 3684
rect 14400 3645 14431 3679
rect 14431 3645 14452 3679
rect 14488 3648 14540 3684
rect 14576 3648 14628 3684
rect 14400 3632 14452 3645
rect 14488 3632 14510 3648
rect 14510 3632 14540 3648
rect 14576 3632 14582 3648
rect 14582 3632 14616 3648
rect 14616 3632 14628 3648
rect 14400 3606 14452 3620
rect 14488 3614 14510 3620
rect 14510 3614 14540 3620
rect 14576 3614 14582 3620
rect 14582 3614 14616 3620
rect 14616 3614 14628 3620
rect 14400 3572 14431 3606
rect 14431 3572 14452 3606
rect 14488 3575 14540 3614
rect 14576 3575 14628 3614
rect 14400 3568 14452 3572
rect 14488 3568 14510 3575
rect 14510 3568 14540 3575
rect 14576 3568 14582 3575
rect 14582 3568 14616 3575
rect 14616 3568 14628 3575
rect 14400 3533 14452 3556
rect 14488 3541 14510 3556
rect 14510 3541 14540 3556
rect 14576 3541 14582 3556
rect 14582 3541 14616 3556
rect 14616 3541 14628 3556
rect 14400 3504 14431 3533
rect 14431 3504 14452 3533
rect 14488 3504 14540 3541
rect 14576 3504 14628 3541
rect 14400 3460 14452 3492
rect 14488 3468 14510 3492
rect 14510 3468 14540 3492
rect 14576 3468 14582 3492
rect 14582 3468 14616 3492
rect 14616 3468 14628 3492
rect 14400 3440 14431 3460
rect 14431 3440 14452 3460
rect 14488 3440 14540 3468
rect 14576 3440 14628 3468
rect 14400 3426 14431 3428
rect 14431 3426 14452 3428
rect 14400 3387 14452 3426
rect 14488 3395 14510 3428
rect 14510 3395 14540 3428
rect 14576 3395 14582 3428
rect 14582 3395 14616 3428
rect 14616 3395 14628 3428
rect 14400 3376 14431 3387
rect 14431 3376 14452 3387
rect 14488 3376 14540 3395
rect 14576 3376 14628 3395
rect 14400 3353 14431 3364
rect 14431 3353 14452 3364
rect 14488 3356 14540 3364
rect 14576 3356 14628 3364
rect 14400 3314 14452 3353
rect 14488 3322 14510 3356
rect 14510 3322 14540 3356
rect 14576 3322 14582 3356
rect 14582 3322 14616 3356
rect 14616 3322 14628 3356
rect 14400 3312 14431 3314
rect 14431 3312 14452 3314
rect 14488 3312 14540 3322
rect 14576 3312 14628 3322
rect 14400 3280 14431 3300
rect 14431 3280 14452 3300
rect 14488 3283 14540 3300
rect 14576 3283 14628 3300
rect 14400 3248 14452 3280
rect 14488 3249 14510 3283
rect 14510 3249 14540 3283
rect 14576 3249 14582 3283
rect 14582 3249 14616 3283
rect 14616 3249 14628 3283
rect 14488 3248 14540 3249
rect 14576 3248 14628 3249
rect 14400 3207 14431 3236
rect 14431 3207 14452 3236
rect 14488 3210 14540 3236
rect 14576 3210 14628 3236
rect 14400 3184 14452 3207
rect 14488 3184 14510 3210
rect 14510 3184 14540 3210
rect 14576 3184 14582 3210
rect 14582 3184 14616 3210
rect 14616 3184 14628 3210
rect 14400 3168 14452 3172
rect 14400 3134 14431 3168
rect 14431 3134 14452 3168
rect 14488 3137 14540 3172
rect 14576 3137 14628 3172
rect 14400 3120 14452 3134
rect 14488 3120 14510 3137
rect 14510 3120 14540 3137
rect 14576 3120 14582 3137
rect 14582 3120 14616 3137
rect 14616 3120 14628 3137
rect 14400 3095 14452 3108
rect 14488 3103 14510 3108
rect 14510 3103 14540 3108
rect 14576 3103 14582 3108
rect 14582 3103 14616 3108
rect 14616 3103 14628 3108
rect 14400 3061 14431 3095
rect 14431 3061 14452 3095
rect 14488 3064 14540 3103
rect 14576 3064 14628 3103
rect 14400 3056 14452 3061
rect 14488 3056 14510 3064
rect 14510 3056 14540 3064
rect 14576 3056 14582 3064
rect 14582 3056 14616 3064
rect 14616 3056 14628 3064
rect 14400 3022 14452 3044
rect 14488 3030 14510 3044
rect 14510 3030 14540 3044
rect 14576 3030 14582 3044
rect 14582 3030 14616 3044
rect 14616 3030 14628 3044
rect 14400 2992 14431 3022
rect 14431 2992 14452 3022
rect 14488 2992 14540 3030
rect 14576 2992 14628 3030
rect 14400 2949 14452 2979
rect 14488 2957 14510 2979
rect 14510 2957 14540 2979
rect 14576 2957 14582 2979
rect 14582 2957 14616 2979
rect 14616 2957 14628 2979
rect 14400 2927 14431 2949
rect 14431 2927 14452 2949
rect 14488 2927 14540 2957
rect 14576 2927 14628 2957
<< metal2 >>
rect 575 4068 14628 4074
rect 627 4016 663 4068
rect 715 4016 751 4068
rect 803 4016 1605 4068
rect 575 4004 1605 4016
rect 627 3952 663 4004
rect 715 3952 751 4004
rect 803 3952 1605 4004
rect 575 3940 1605 3952
rect 627 3888 663 3940
rect 715 3888 751 3940
rect 803 3888 1605 3940
rect 575 3876 1605 3888
rect 627 3824 663 3876
rect 715 3824 751 3876
rect 803 3824 1605 3876
rect 575 3812 1605 3824
rect 627 3760 663 3812
rect 715 3760 751 3812
rect 803 3760 1605 3812
rect 575 3748 1605 3760
rect 627 3696 663 3748
rect 715 3696 751 3748
rect 803 3696 1605 3748
rect 575 3684 1605 3696
rect 627 3632 663 3684
rect 715 3632 751 3684
rect 803 3632 1605 3684
rect 575 3620 1605 3632
rect 627 3568 663 3620
rect 715 3568 751 3620
rect 803 3568 1605 3620
rect 575 3556 1605 3568
rect 627 3504 663 3556
rect 715 3504 751 3556
rect 803 3504 1605 3556
rect 575 3492 1605 3504
rect 627 3440 663 3492
rect 715 3440 751 3492
rect 803 3440 1605 3492
rect 575 3428 1605 3440
rect 627 3376 663 3428
rect 715 3376 751 3428
rect 803 3376 1605 3428
rect 575 3364 1605 3376
rect 627 3312 663 3364
rect 715 3312 751 3364
rect 803 3312 1605 3364
rect 575 3300 1605 3312
rect 627 3248 663 3300
rect 715 3248 751 3300
rect 803 3248 1605 3300
rect 575 3236 1605 3248
rect 627 3184 663 3236
rect 715 3184 751 3236
rect 803 3184 1605 3236
rect 575 3172 1605 3184
rect 627 3120 663 3172
rect 715 3120 751 3172
rect 803 3120 1605 3172
rect 575 3108 1605 3120
rect 627 3056 663 3108
rect 715 3056 751 3108
rect 803 3056 1605 3108
rect 575 3044 1605 3056
rect 627 2992 663 3044
rect 715 2992 751 3044
rect 803 2992 1605 3044
rect 1785 2992 2597 4068
rect 2777 2992 3589 4068
rect 3769 2992 4581 4068
rect 4761 2992 5573 4068
rect 5753 2992 6565 4068
rect 6745 2992 7557 4068
rect 7737 2992 8549 4068
rect 8729 2992 9541 4068
rect 9721 2992 10533 4068
rect 10713 2992 11525 4068
rect 11705 2992 12517 4068
rect 12697 2992 13509 4068
rect 13689 4016 14400 4068
rect 14452 4016 14488 4068
rect 14540 4016 14576 4068
rect 13689 4004 14628 4016
rect 13689 3952 14400 4004
rect 14452 3952 14488 4004
rect 14540 3952 14576 4004
rect 13689 3940 14628 3952
rect 13689 3888 14400 3940
rect 14452 3888 14488 3940
rect 14540 3888 14576 3940
rect 13689 3876 14628 3888
rect 13689 3824 14400 3876
rect 14452 3824 14488 3876
rect 14540 3824 14576 3876
rect 13689 3812 14628 3824
rect 13689 3760 14400 3812
rect 14452 3760 14488 3812
rect 14540 3760 14576 3812
rect 13689 3748 14628 3760
rect 13689 3696 14400 3748
rect 14452 3696 14488 3748
rect 14540 3696 14576 3748
rect 13689 3684 14628 3696
rect 13689 3632 14400 3684
rect 14452 3632 14488 3684
rect 14540 3632 14576 3684
rect 13689 3620 14628 3632
rect 13689 3568 14400 3620
rect 14452 3568 14488 3620
rect 14540 3568 14576 3620
rect 13689 3556 14628 3568
rect 13689 3504 14400 3556
rect 14452 3504 14488 3556
rect 14540 3504 14576 3556
rect 13689 3492 14628 3504
rect 13689 3440 14400 3492
rect 14452 3440 14488 3492
rect 14540 3440 14576 3492
rect 13689 3428 14628 3440
rect 13689 3376 14400 3428
rect 14452 3376 14488 3428
rect 14540 3376 14576 3428
rect 13689 3364 14628 3376
rect 13689 3312 14400 3364
rect 14452 3312 14488 3364
rect 14540 3312 14576 3364
rect 13689 3300 14628 3312
rect 13689 3248 14400 3300
rect 14452 3248 14488 3300
rect 14540 3248 14576 3300
rect 13689 3236 14628 3248
rect 13689 3184 14400 3236
rect 14452 3184 14488 3236
rect 14540 3184 14576 3236
rect 13689 3172 14628 3184
rect 13689 3120 14400 3172
rect 14452 3120 14488 3172
rect 14540 3120 14576 3172
rect 13689 3108 14628 3120
rect 13689 3056 14400 3108
rect 14452 3056 14488 3108
rect 14540 3056 14576 3108
rect 13689 3044 14628 3056
rect 13689 2992 14400 3044
rect 14452 2992 14488 3044
rect 14540 2992 14576 3044
rect 575 2979 14628 2992
rect 627 2927 663 2979
rect 715 2927 751 2979
rect 803 2927 1605 2979
rect 1657 2927 1669 2979
rect 1721 2927 1733 2979
rect 1785 2927 2597 2979
rect 2649 2927 2661 2979
rect 2713 2927 2725 2979
rect 2777 2927 3589 2979
rect 3641 2927 3653 2979
rect 3705 2927 3717 2979
rect 3769 2927 4581 2979
rect 4633 2927 4645 2979
rect 4697 2927 4709 2979
rect 4761 2927 5573 2979
rect 5625 2927 5637 2979
rect 5689 2927 5701 2979
rect 5753 2927 6565 2979
rect 6617 2927 6629 2979
rect 6681 2927 6693 2979
rect 6745 2927 7557 2979
rect 7609 2927 7621 2979
rect 7673 2927 7685 2979
rect 7737 2927 8549 2979
rect 8601 2927 8613 2979
rect 8665 2927 8677 2979
rect 8729 2927 9541 2979
rect 9593 2927 9605 2979
rect 9657 2927 9669 2979
rect 9721 2927 10533 2979
rect 10585 2927 10597 2979
rect 10649 2927 10661 2979
rect 10713 2927 11525 2979
rect 11577 2927 11589 2979
rect 11641 2927 11653 2979
rect 11705 2927 12517 2979
rect 12569 2927 12581 2979
rect 12633 2927 12645 2979
rect 12697 2927 13509 2979
rect 13561 2927 13573 2979
rect 13625 2927 13637 2979
rect 13689 2927 14400 2979
rect 14452 2927 14488 2979
rect 14540 2927 14576 2979
rect 575 2921 14628 2927
rect 1104 2614 14226 2620
rect 1104 1538 1109 2614
rect 1289 1538 2101 2614
rect 2281 1538 3093 2614
rect 3273 1538 4085 2614
rect 4265 1538 5077 2614
rect 5257 1538 6069 2614
rect 6249 1538 7061 2614
rect 7241 1538 8053 2614
rect 8233 1538 9045 2614
rect 9225 1538 10037 2614
rect 10217 1538 11029 2614
rect 11209 1538 12021 2614
rect 12201 1538 13013 2614
rect 13193 2562 14037 2614
rect 14089 2562 14105 2614
rect 14157 2562 14173 2614
rect 14225 2562 14226 2614
rect 13193 2550 14226 2562
rect 13193 2498 14037 2550
rect 14089 2498 14105 2550
rect 14157 2498 14173 2550
rect 14225 2498 14226 2550
rect 13193 2486 14226 2498
rect 13193 2434 14037 2486
rect 14089 2434 14105 2486
rect 14157 2434 14173 2486
rect 14225 2434 14226 2486
rect 13193 2422 14226 2434
rect 13193 2370 14037 2422
rect 14089 2370 14105 2422
rect 14157 2370 14173 2422
rect 14225 2370 14226 2422
rect 13193 2358 14226 2370
rect 13193 2306 14037 2358
rect 14089 2306 14105 2358
rect 14157 2306 14173 2358
rect 14225 2306 14226 2358
rect 13193 2294 14226 2306
rect 13193 2242 14037 2294
rect 14089 2242 14105 2294
rect 14157 2242 14173 2294
rect 14225 2242 14226 2294
rect 13193 2230 14226 2242
rect 13193 2178 14037 2230
rect 14089 2178 14105 2230
rect 14157 2178 14173 2230
rect 14225 2178 14226 2230
rect 13193 2166 14226 2178
rect 13193 2114 14037 2166
rect 14089 2114 14105 2166
rect 14157 2114 14173 2166
rect 14225 2114 14226 2166
rect 13193 2102 14226 2114
rect 13193 2050 14037 2102
rect 14089 2050 14105 2102
rect 14157 2050 14173 2102
rect 14225 2050 14226 2102
rect 13193 2038 14226 2050
rect 13193 1986 14037 2038
rect 14089 1986 14105 2038
rect 14157 1986 14173 2038
rect 14225 1986 14226 2038
rect 13193 1974 14226 1986
rect 13193 1922 14037 1974
rect 14089 1922 14105 1974
rect 14157 1922 14173 1974
rect 14225 1922 14226 1974
rect 13193 1910 14226 1922
rect 13193 1858 14037 1910
rect 14089 1858 14105 1910
rect 14157 1858 14173 1910
rect 14225 1858 14226 1910
rect 13193 1846 14226 1858
rect 13193 1794 14037 1846
rect 14089 1794 14105 1846
rect 14157 1794 14173 1846
rect 14225 1794 14226 1846
rect 13193 1782 14226 1794
rect 13193 1730 14037 1782
rect 14089 1730 14105 1782
rect 14157 1730 14173 1782
rect 14225 1730 14226 1782
rect 13193 1718 14226 1730
rect 13193 1666 14037 1718
rect 14089 1666 14105 1718
rect 14157 1666 14173 1718
rect 14225 1666 14226 1718
rect 13193 1654 14226 1666
rect 13193 1602 14037 1654
rect 14089 1602 14105 1654
rect 14157 1602 14173 1654
rect 14225 1602 14226 1654
rect 13193 1590 14226 1602
rect 13193 1538 14037 1590
rect 14089 1538 14105 1590
rect 14157 1538 14173 1590
rect 14225 1538 14226 1590
rect 1104 1525 14226 1538
rect 1104 1473 1109 1525
rect 1161 1473 1173 1525
rect 1225 1473 1237 1525
rect 1289 1473 2101 1525
rect 2153 1473 2165 1525
rect 2217 1473 2229 1525
rect 2281 1473 3093 1525
rect 3145 1473 3157 1525
rect 3209 1473 3221 1525
rect 3273 1473 4085 1525
rect 4137 1473 4149 1525
rect 4201 1473 4213 1525
rect 4265 1473 5077 1525
rect 5129 1473 5141 1525
rect 5193 1473 5205 1525
rect 5257 1473 6069 1525
rect 6121 1473 6133 1525
rect 6185 1473 6197 1525
rect 6249 1473 7061 1525
rect 7113 1473 7125 1525
rect 7177 1473 7189 1525
rect 7241 1473 8053 1525
rect 8105 1473 8117 1525
rect 8169 1473 8181 1525
rect 8233 1473 9045 1525
rect 9097 1473 9109 1525
rect 9161 1473 9173 1525
rect 9225 1473 10037 1525
rect 10089 1473 10101 1525
rect 10153 1473 10165 1525
rect 10217 1473 11029 1525
rect 11081 1473 11093 1525
rect 11145 1473 11157 1525
rect 11209 1473 12021 1525
rect 12073 1473 12085 1525
rect 12137 1473 12149 1525
rect 12201 1473 13013 1525
rect 13065 1473 13077 1525
rect 13129 1473 13141 1525
rect 13193 1473 14037 1525
rect 14089 1473 14105 1525
rect 14157 1473 14173 1525
rect 14225 1473 14226 1525
rect 1104 1467 14226 1473
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_0
timestamp 1701704242
transform 1 0 14031 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_1
timestamp 1701704242
transform 1 0 14031 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_2
timestamp 1701704242
transform 1 0 8079 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_3
timestamp 1701704242
transform 1 0 9071 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_4
timestamp 1701704242
transform 1 0 10063 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_5
timestamp 1701704242
transform 1 0 11055 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_6
timestamp 1701704242
transform 1 0 12047 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_7
timestamp 1701704242
transform 1 0 13039 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_8
timestamp 1701704242
transform 1 0 8151 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_9
timestamp 1701704242
transform 1 0 9143 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_10
timestamp 1701704242
transform 1 0 10135 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_11
timestamp 1701704242
transform 1 0 11127 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_12
timestamp 1701704242
transform 1 0 12119 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_13
timestamp 1701704242
transform 1 0 13111 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_14
timestamp 1701704242
transform 1 0 13111 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_15
timestamp 1701704242
transform 1 0 12119 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_16
timestamp 1701704242
transform 1 0 11127 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_17
timestamp 1701704242
transform 1 0 10135 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_18
timestamp 1701704242
transform 1 0 9143 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_19
timestamp 1701704242
transform 1 0 8151 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_20
timestamp 1701704242
transform 1 0 13039 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_21
timestamp 1701704242
transform 1 0 12047 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_22
timestamp 1701704242
transform 1 0 11055 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_23
timestamp 1701704242
transform 1 0 10063 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_24
timestamp 1701704242
transform 1 0 9071 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_25
timestamp 1701704242
transform 1 0 8079 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_26
timestamp 1701704242
transform 1 0 1135 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_27
timestamp 1701704242
transform 1 0 1207 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_28
timestamp 1701704242
transform 1 0 2199 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_29
timestamp 1701704242
transform 1 0 2127 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_30
timestamp 1701704242
transform 1 0 1135 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_31
timestamp 1701704242
transform 1 0 1207 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_32
timestamp 1701704242
transform 1 0 2199 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_33
timestamp 1701704242
transform 1 0 2127 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_34
timestamp 1701704242
transform 1 0 3119 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_35
timestamp 1701704242
transform 1 0 4111 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_36
timestamp 1701704242
transform 1 0 5103 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_37
timestamp 1701704242
transform 1 0 6095 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_38
timestamp 1701704242
transform 1 0 7087 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_39
timestamp 1701704242
transform 1 0 3191 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_40
timestamp 1701704242
transform 1 0 4183 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_41
timestamp 1701704242
transform 1 0 5175 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_42
timestamp 1701704242
transform 1 0 6167 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_43
timestamp 1701704242
transform 1 0 7159 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_44
timestamp 1701704242
transform 1 0 7159 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_45
timestamp 1701704242
transform 1 0 6167 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_46
timestamp 1701704242
transform 1 0 5175 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_47
timestamp 1701704242
transform 1 0 4183 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_48
timestamp 1701704242
transform 1 0 3191 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_49
timestamp 1701704242
transform 1 0 7087 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_50
timestamp 1701704242
transform 1 0 6095 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_51
timestamp 1701704242
transform 1 0 5103 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_52
timestamp 1701704242
transform 1 0 4111 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_53
timestamp 1701704242
transform 1 0 3119 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808645  sky130_fd_pr__nfet_01v8__example_55959141808645_0
timestamp 1701704242
transform 1 0 924 0 -1 2457
box -78 0 -77 1
use sky130_fd_pr__nfet_01v8__example_55959141808647  sky130_fd_pr__nfet_01v8__example_55959141808647_0
timestamp 1701704242
transform 1 0 924 0 -1 4058
box -78 0 -77 1
use sky130_fd_pr__nfet_01v8__example_55959141808647  sky130_fd_pr__nfet_01v8__example_55959141808647_1
timestamp 1701704242
transform -1 0 14298 0 -1 2457
box -78 0 -77 1
use sky130_fd_pr__nfet_01v8__example_55959141808647  sky130_fd_pr__nfet_01v8__example_55959141808647_2
timestamp 1701704242
transform -1 0 14298 0 -1 4058
box -78 0 -77 1
use sky130_fd_pr__nfet_01v8__example_55959141808648  sky130_fd_pr__nfet_01v8__example_55959141808648_0
timestamp 1701704242
transform 1 0 1916 0 -1 4058
box 641 0 11554 1
use sky130_fd_pr__nfet_01v8__example_55959141808650  sky130_fd_pr__nfet_01v8__example_55959141808650_0
timestamp 1701704242
transform -1 0 1474 0 -1 2457
box -92 0 -91 1
use sky130_fd_pr__nfet_01v8__example_55959141808650  sky130_fd_pr__nfet_01v8__example_55959141808650_1
timestamp 1701704242
transform -1 0 1474 0 -1 4058
box -92 0 -91 1
use sky130_fd_pr__nfet_01v8__example_55959141808651  sky130_fd_pr__nfet_01v8__example_55959141808651_0
timestamp 1701704242
transform 1 0 1916 0 -1 2457
box 641 0 11554 1
use sky130_fd_pr__via_l1m1_centered__example_559591418082  sky130_fd_pr__via_l1m1_centered__example_559591418082_0
timestamp 1701704242
transform 1 0 15088 0 1 507
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418082  sky130_fd_pr__via_l1m1_centered__example_559591418082_1
timestamp 1701704242
transform -1 0 88 0 1 513
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418083  sky130_fd_pr__via_l1m1_centered__example_559591418083_0
timestamp 1701704242
transform 0 -1 14869 -1 0 507
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418083  sky130_fd_pr__via_l1m1_centered__example_559591418083_1
timestamp 1701704242
transform 0 -1 14869 1 0 5409
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_0
timestamp 1701704242
transform 1 0 14238 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_1
timestamp 1701704242
transform 1 0 12888 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_2
timestamp 1701704242
transform 1 0 13880 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_3
timestamp 1701704242
transform 1 0 13318 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_4
timestamp 1701704242
transform 1 0 12326 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_5
timestamp 1701704242
transform 1 0 11334 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_6
timestamp 1701704242
transform 1 0 10342 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_7
timestamp 1701704242
transform 1 0 9350 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_8
timestamp 1701704242
transform 1 0 8358 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_9
timestamp 1701704242
transform 1 0 7366 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_10
timestamp 1701704242
transform 1 0 6374 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_11
timestamp 1701704242
transform 1 0 5382 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_12
timestamp 1701704242
transform 1 0 8920 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_13
timestamp 1701704242
transform 1 0 7928 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_14
timestamp 1701704242
transform 1 0 6921 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_15
timestamp 1701704242
transform 1 0 5944 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_16
timestamp 1701704242
transform 1 0 4952 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_17
timestamp 1701704242
transform 1 0 3960 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_18
timestamp 1701704242
transform 1 0 2968 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_19
timestamp 1701704242
transform 1 0 1976 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_20
timestamp 1701704242
transform 1 0 984 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_21
timestamp 1701704242
transform 1 0 3398 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_22
timestamp 1701704242
transform 1 0 2406 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_23
timestamp 1701704242
transform 1 0 1414 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_24
timestamp 1701704242
transform 1 0 11896 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_25
timestamp 1701704242
transform 1 0 10904 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_26
timestamp 1701704242
transform 1 0 9912 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_27
timestamp 1701704242
transform 1 0 4390 0 1 4441
box 0 0 1 1
<< labels >>
flabel metal1 s 13239 5295 13646 5426 0 FreeSans 44 0 0 0 VCC_IO
port 2 nsew
flabel metal2 s 11977 2924 13386 4028 0 FreeSans 44 0 0 0 VSSIO
port 3 nsew
flabel metal2 s 11655 1819 12696 2443 0 FreeSans 44 0 0 0 PAD
port 4 nsew
<< properties >>
string GDS_END 18015922
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 17406758
<< end >>
