magic
tech sky130B
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808587  sky130_fd_pr__model__nfet_highvoltage__example_55959141808587_0
timestamp 1701704242
transform 1 0 478 0 -1 1701
box -1 0 101 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808588  sky130_fd_pr__model__pfet_highvoltage__example_55959141808588_0
timestamp 1701704242
transform 1 0 291 0 -1 3319
box -1 0 101 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808588  sky130_fd_pr__model__pfet_highvoltage__example_55959141808588_1
timestamp 1701704242
transform 1 0 447 0 -1 3319
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_0
timestamp 1701704242
transform 1 0 946 0 1 665
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_1
timestamp 1701704242
transform -1 0 890 0 1 665
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_0
timestamp 1701704242
transform 1 0 1190 0 1 1501
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_1
timestamp 1701704242
transform 1 0 910 0 1 1501
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_2
timestamp 1701704242
transform -1 0 854 0 1 1501
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808589  sky130_fd_pr__nfet_01v8__example_55959141808589_0
timestamp 1701704242
transform -1 0 1638 0 1 665
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_0
timestamp 1701704242
transform 1 0 883 0 1 3019
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_1
timestamp 1701704242
transform -1 0 827 0 1 3019
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1701704242
transform -1 0 1520 0 1 3235
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1701704242
transform 1 0 1576 0 1 3235
box -1 0 201 1
<< properties >>
string GDS_END 22042252
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22015142
<< end >>
