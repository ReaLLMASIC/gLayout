magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -68 -26 1354 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 1286 50 1328 66
rect 1320 16 1328 50
rect 1286 0 1328 16
<< ndiffc >>
rect -34 16 0 50
rect 1286 16 1320 50
<< ndiffres >>
rect 0 0 1286 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 1286 50 1320 66
rect 1286 0 1320 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 1 0 1278 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 86502650
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86502148
<< end >>
