magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 0 470 544 476
rect 0 0 544 6
<< via3 >>
rect 0 6 544 470
<< metal4 >>
rect -1 470 545 471
rect -1 6 0 470
rect 544 6 545 470
rect -1 5 545 6
<< properties >>
string GDS_END 93355782
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93352962
<< end >>
