magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2023 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1219 47 1249 177
rect 1303 47 1333 177
rect 1387 47 1417 177
rect 1471 47 1501 177
rect 1659 47 1689 177
rect 1743 47 1773 177
rect 1827 47 1857 177
rect 1911 47 1941 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 755 297 785 497
rect 839 297 869 497
rect 923 297 953 497
rect 1088 297 1118 497
rect 1219 297 1249 497
rect 1303 297 1333 497
rect 1387 297 1417 497
rect 1471 297 1501 497
rect 1659 297 1689 497
rect 1743 297 1773 497
rect 1827 297 1857 497
rect 1911 297 1941 497
<< ndiff >>
rect 27 101 79 177
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 101 247 177
rect 193 67 203 101
rect 237 67 247 101
rect 193 47 247 67
rect 277 93 331 177
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 109 415 177
rect 361 75 371 109
rect 405 75 415 109
rect 361 47 415 75
rect 445 161 499 177
rect 445 127 455 161
rect 489 127 499 161
rect 445 47 499 127
rect 529 93 583 177
rect 529 59 539 93
rect 573 59 583 93
rect 529 47 583 59
rect 613 161 667 177
rect 613 127 623 161
rect 657 127 667 161
rect 613 47 667 127
rect 697 93 749 177
rect 697 59 707 93
rect 741 59 749 93
rect 697 47 749 59
rect 803 93 855 177
rect 803 59 811 93
rect 845 59 855 93
rect 803 47 855 59
rect 885 161 939 177
rect 885 127 895 161
rect 929 127 939 161
rect 885 47 939 127
rect 969 93 1023 177
rect 969 59 979 93
rect 1013 59 1023 93
rect 969 47 1023 59
rect 1053 161 1107 177
rect 1053 127 1063 161
rect 1097 127 1107 161
rect 1053 47 1107 127
rect 1137 93 1219 177
rect 1137 59 1147 93
rect 1181 59 1219 93
rect 1137 47 1219 59
rect 1249 161 1303 177
rect 1249 127 1259 161
rect 1293 127 1303 161
rect 1249 47 1303 127
rect 1333 93 1387 177
rect 1333 59 1343 93
rect 1377 59 1387 93
rect 1333 47 1387 59
rect 1417 161 1471 177
rect 1417 127 1427 161
rect 1461 127 1471 161
rect 1417 47 1471 127
rect 1501 93 1553 177
rect 1501 59 1511 93
rect 1545 59 1553 93
rect 1501 47 1553 59
rect 1607 93 1659 177
rect 1607 59 1615 93
rect 1649 59 1659 93
rect 1607 47 1659 59
rect 1689 101 1743 177
rect 1689 67 1699 101
rect 1733 67 1743 101
rect 1689 47 1743 67
rect 1773 93 1827 177
rect 1773 59 1783 93
rect 1817 59 1827 93
rect 1773 47 1827 59
rect 1857 101 1911 177
rect 1857 67 1867 101
rect 1901 67 1911 101
rect 1857 47 1911 67
rect 1941 93 1997 177
rect 1941 59 1953 93
rect 1987 59 1997 93
rect 1941 47 1997 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 297 79 451
rect 109 417 163 497
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 297 247 451
rect 277 417 331 497
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 297 415 451
rect 445 417 499 497
rect 445 383 455 417
rect 489 383 499 417
rect 445 349 499 383
rect 445 315 455 349
rect 489 315 499 349
rect 445 297 499 315
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 297 583 451
rect 613 417 667 497
rect 613 383 623 417
rect 657 383 667 417
rect 613 349 667 383
rect 613 315 623 349
rect 657 315 667 349
rect 613 297 667 315
rect 697 469 755 497
rect 697 435 707 469
rect 741 435 755 469
rect 697 297 755 435
rect 785 485 839 497
rect 785 451 795 485
rect 829 451 839 485
rect 785 417 839 451
rect 785 383 795 417
rect 829 383 839 417
rect 785 297 839 383
rect 869 477 923 497
rect 869 443 879 477
rect 913 443 923 477
rect 869 409 923 443
rect 869 375 879 409
rect 913 375 923 409
rect 869 297 923 375
rect 953 485 1088 497
rect 953 383 970 485
rect 1072 383 1088 485
rect 953 297 1088 383
rect 1118 477 1219 497
rect 1118 443 1128 477
rect 1162 443 1219 477
rect 1118 409 1219 443
rect 1118 375 1128 409
rect 1162 375 1219 409
rect 1118 297 1219 375
rect 1249 485 1303 497
rect 1249 451 1259 485
rect 1293 451 1303 485
rect 1249 417 1303 451
rect 1249 383 1259 417
rect 1293 383 1303 417
rect 1249 297 1303 383
rect 1333 477 1387 497
rect 1333 443 1343 477
rect 1377 443 1387 477
rect 1333 409 1387 443
rect 1333 375 1343 409
rect 1377 375 1387 409
rect 1333 297 1387 375
rect 1417 485 1471 497
rect 1417 451 1427 485
rect 1461 451 1471 485
rect 1417 297 1471 451
rect 1501 477 1659 497
rect 1501 443 1511 477
rect 1545 443 1659 477
rect 1501 409 1659 443
rect 1501 375 1511 409
rect 1545 375 1659 409
rect 1501 297 1659 375
rect 1689 485 1743 497
rect 1689 451 1699 485
rect 1733 451 1743 485
rect 1689 417 1743 451
rect 1689 383 1699 417
rect 1733 383 1743 417
rect 1689 297 1743 383
rect 1773 477 1827 497
rect 1773 443 1783 477
rect 1817 443 1827 477
rect 1773 409 1827 443
rect 1773 375 1783 409
rect 1817 375 1827 409
rect 1773 297 1827 375
rect 1857 485 1911 497
rect 1857 451 1867 485
rect 1901 451 1911 485
rect 1857 417 1911 451
rect 1857 383 1867 417
rect 1901 383 1911 417
rect 1857 297 1911 383
rect 1941 477 1993 497
rect 1941 443 1951 477
rect 1985 443 1993 477
rect 1941 409 1993 443
rect 1941 375 1951 409
rect 1985 375 1993 409
rect 1941 297 1993 375
<< ndiffc >>
rect 35 67 69 101
rect 119 59 153 93
rect 203 67 237 101
rect 287 59 321 93
rect 371 75 405 109
rect 455 127 489 161
rect 539 59 573 93
rect 623 127 657 161
rect 707 59 741 93
rect 811 59 845 93
rect 895 127 929 161
rect 979 59 1013 93
rect 1063 127 1097 161
rect 1147 59 1181 93
rect 1259 127 1293 161
rect 1343 59 1377 93
rect 1427 127 1461 161
rect 1511 59 1545 93
rect 1615 59 1649 93
rect 1699 67 1733 101
rect 1783 59 1817 93
rect 1867 67 1901 101
rect 1953 59 1987 93
<< pdiffc >>
rect 35 451 69 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 455 383 489 417
rect 455 315 489 349
rect 539 451 573 485
rect 623 383 657 417
rect 623 315 657 349
rect 707 435 741 469
rect 795 451 829 485
rect 795 383 829 417
rect 879 443 913 477
rect 879 375 913 409
rect 970 383 1072 485
rect 1128 443 1162 477
rect 1128 375 1162 409
rect 1259 451 1293 485
rect 1259 383 1293 417
rect 1343 443 1377 477
rect 1343 375 1377 409
rect 1427 451 1461 485
rect 1511 443 1545 477
rect 1511 375 1545 409
rect 1699 451 1733 485
rect 1699 383 1733 417
rect 1783 443 1817 477
rect 1783 375 1817 409
rect 1867 451 1901 485
rect 1867 383 1901 417
rect 1951 443 1985 477
rect 1951 375 1985 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 755 497 785 523
rect 839 497 869 523
rect 923 497 953 523
rect 1088 497 1118 523
rect 1219 497 1249 523
rect 1303 497 1333 523
rect 1387 497 1417 523
rect 1471 497 1501 523
rect 1659 497 1689 523
rect 1743 497 1773 523
rect 1827 497 1857 523
rect 1911 497 1941 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 261 361 265
rect 22 249 361 261
rect 22 215 38 249
rect 72 215 106 249
rect 140 215 174 249
rect 208 215 242 249
rect 276 215 361 249
rect 22 203 361 215
rect 79 199 361 203
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 415 249 697 265
rect 415 215 517 249
rect 551 215 585 249
rect 619 215 653 249
rect 687 215 697 249
rect 415 199 697 215
rect 755 269 785 297
rect 839 269 869 297
rect 923 269 953 297
rect 1088 269 1118 297
rect 755 265 1118 269
rect 1219 269 1249 297
rect 1303 269 1333 297
rect 1387 269 1417 297
rect 1471 269 1501 297
rect 755 249 1137 265
rect 755 215 771 249
rect 805 215 839 249
rect 873 215 907 249
rect 941 215 975 249
rect 1009 215 1043 249
rect 1077 215 1137 249
rect 755 202 1137 215
rect 755 199 1053 202
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 202
rect 1219 249 1501 269
rect 1219 215 1235 249
rect 1269 215 1303 249
rect 1337 215 1371 249
rect 1405 215 1439 249
rect 1473 215 1501 249
rect 1219 202 1501 215
rect 1219 199 1417 202
rect 1219 177 1249 199
rect 1303 177 1333 199
rect 1387 177 1417 199
rect 1471 177 1501 202
rect 1659 265 1689 297
rect 1743 265 1773 297
rect 1827 265 1857 297
rect 1911 265 1941 297
rect 1659 261 1941 265
rect 1659 249 1997 261
rect 1659 215 1675 249
rect 1709 215 1743 249
rect 1777 215 1811 249
rect 1845 215 1879 249
rect 1913 215 1947 249
rect 1981 215 1997 249
rect 1659 203 1997 215
rect 1659 199 1941 203
rect 1659 177 1689 199
rect 1743 177 1773 199
rect 1827 177 1857 199
rect 1911 177 1941 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1219 21 1249 47
rect 1303 21 1333 47
rect 1387 21 1417 47
rect 1471 21 1501 47
rect 1659 21 1689 47
rect 1743 21 1773 47
rect 1827 21 1857 47
rect 1911 21 1941 47
<< polycont >>
rect 38 215 72 249
rect 106 215 140 249
rect 174 215 208 249
rect 242 215 276 249
rect 517 215 551 249
rect 585 215 619 249
rect 653 215 687 249
rect 771 215 805 249
rect 839 215 873 249
rect 907 215 941 249
rect 975 215 1009 249
rect 1043 215 1077 249
rect 1235 215 1269 249
rect 1303 215 1337 249
rect 1371 215 1405 249
rect 1439 215 1473 249
rect 1675 215 1709 249
rect 1743 215 1777 249
rect 1811 215 1845 249
rect 1879 215 1913 249
rect 1947 215 1981 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 779 485 845 527
rect 19 451 35 485
rect 69 451 203 485
rect 237 451 371 485
rect 405 451 539 485
rect 573 469 741 485
rect 573 451 707 469
rect 22 261 66 393
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 271 383 287 417
rect 321 383 337 417
rect 271 349 337 383
rect 395 383 455 417
rect 489 383 505 417
rect 395 349 505 383
rect 607 383 623 417
rect 657 383 673 417
rect 607 349 673 383
rect 103 315 119 349
rect 153 315 287 349
rect 321 315 455 349
rect 489 315 623 349
rect 657 315 673 349
rect 707 349 741 435
rect 779 451 795 485
rect 829 451 845 485
rect 779 417 845 451
rect 779 383 795 417
rect 829 383 845 417
rect 879 477 913 493
rect 879 409 913 443
rect 954 485 1088 527
rect 954 383 970 485
rect 1072 383 1088 485
rect 1128 477 1162 493
rect 1128 409 1162 443
rect 879 349 913 375
rect 1243 485 1309 527
rect 1243 451 1259 485
rect 1293 451 1309 485
rect 1243 417 1309 451
rect 1243 383 1259 417
rect 1293 383 1309 417
rect 1343 477 1377 493
rect 1343 409 1377 443
rect 1128 349 1162 375
rect 1411 485 1477 527
rect 1411 451 1427 485
rect 1461 451 1477 485
rect 1411 383 1477 451
rect 1511 477 1545 493
rect 1511 409 1545 443
rect 1343 349 1377 375
rect 1683 485 1749 527
rect 1683 451 1699 485
rect 1733 451 1749 485
rect 1683 417 1749 451
rect 1683 383 1699 417
rect 1733 383 1749 417
rect 1783 477 1817 493
rect 1783 409 1817 443
rect 1511 349 1545 375
rect 1851 485 1917 527
rect 1851 451 1867 485
rect 1901 451 1917 485
rect 1851 417 1917 451
rect 1851 383 1867 417
rect 1901 383 1917 417
rect 1951 477 1985 493
rect 1951 409 1985 443
rect 1783 349 1817 375
rect 1951 349 1985 375
rect 707 315 1985 349
rect 22 249 350 261
rect 22 215 38 249
rect 72 215 106 249
rect 140 215 174 249
rect 208 215 242 249
rect 276 215 350 249
rect 395 198 473 315
rect 517 249 711 265
rect 551 215 585 249
rect 619 215 653 249
rect 687 215 711 249
rect 755 249 1093 257
rect 755 215 771 249
rect 805 215 839 249
rect 873 215 907 249
rect 941 215 975 249
rect 1009 215 1043 249
rect 1077 215 1093 249
rect 1219 249 1539 260
rect 1219 215 1235 249
rect 1269 215 1303 249
rect 1337 215 1371 249
rect 1405 215 1439 249
rect 1473 215 1539 249
rect 1659 249 1997 256
rect 1659 215 1675 249
rect 1709 215 1743 249
rect 1777 215 1811 249
rect 1845 215 1879 249
rect 1913 215 1947 249
rect 1981 215 1997 249
rect 517 199 711 215
rect 439 161 473 198
rect 35 127 405 161
rect 439 127 455 161
rect 489 127 623 161
rect 657 127 895 161
rect 929 127 1063 161
rect 1097 127 1113 161
rect 1243 127 1259 161
rect 1293 127 1427 161
rect 1461 127 1901 161
rect 1961 151 1997 215
rect 35 101 69 127
rect 203 101 237 127
rect 35 51 69 67
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 371 109 405 127
rect 203 51 237 67
rect 271 59 287 93
rect 321 59 337 93
rect 1699 101 1733 127
rect 405 75 539 93
rect 371 59 539 75
rect 573 59 707 93
rect 741 59 757 93
rect 795 59 811 93
rect 845 59 979 93
rect 1013 59 1147 93
rect 1181 59 1343 93
rect 1377 59 1511 93
rect 1545 59 1561 93
rect 1599 59 1615 93
rect 1649 59 1665 93
rect 271 17 337 59
rect 1599 17 1665 59
rect 1867 101 1901 127
rect 1699 51 1733 67
rect 1767 59 1783 93
rect 1817 59 1833 93
rect 1767 17 1833 59
rect 1867 51 1901 67
rect 1937 59 1953 93
rect 1987 59 2005 93
rect 1937 17 2005 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 1962 221 1996 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1870 221 1904 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1778 221 1812 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1686 221 1720 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1498 221 1532 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1406 221 1440 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1314 221 1348 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1222 221 1256 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1962 153 1996 187 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 30 357 64 391 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1046 221 1080 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
rlabel comment s 0 0 0 0 4 a32oi_4
rlabel metal1 s 0 -48 2024 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 3501186
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3485012
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
