magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 89 233
<< metal1 >>
rect -6 233 95 236
rect -6 0 0 233
rect 89 0 95 233
rect -6 -3 95 0
<< properties >>
string GDS_END 79706572
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79705096
<< end >>
