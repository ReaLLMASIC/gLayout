magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal4 >>
rect 0 39530 9600 39593
rect 0 34814 422 39530
rect 9298 34814 9600 39530
rect 0 34750 9600 34814
rect 0 18565 9600 18593
rect 0 18329 421 18565
rect 657 18329 741 18565
rect 977 18329 1061 18565
rect 1297 18329 1381 18565
rect 1617 18329 1701 18565
rect 1937 18329 2021 18565
rect 2257 18329 2341 18565
rect 2577 18329 2661 18565
rect 2897 18329 2981 18565
rect 3217 18329 3301 18565
rect 3537 18329 3621 18565
rect 3857 18329 3941 18565
rect 4177 18329 4261 18565
rect 4497 18329 4581 18565
rect 4817 18329 4901 18565
rect 5137 18329 5221 18565
rect 5457 18329 5541 18565
rect 5777 18329 5861 18565
rect 6097 18329 6181 18565
rect 6417 18329 6501 18565
rect 6737 18329 6821 18565
rect 7057 18329 7141 18565
rect 7377 18329 7461 18565
rect 7697 18329 7781 18565
rect 8017 18329 8101 18565
rect 8337 18329 8421 18565
rect 8657 18329 8741 18565
rect 8977 18329 9061 18565
rect 9297 18329 9600 18565
rect 0 18229 9600 18329
rect 0 17993 421 18229
rect 657 17993 741 18229
rect 977 17993 1061 18229
rect 1297 17993 1381 18229
rect 1617 17993 1701 18229
rect 1937 17993 2021 18229
rect 2257 17993 2341 18229
rect 2577 17993 2661 18229
rect 2897 17993 2981 18229
rect 3217 17993 3301 18229
rect 3537 17993 3621 18229
rect 3857 17993 3941 18229
rect 4177 17993 4261 18229
rect 4497 17993 4581 18229
rect 4817 17993 4901 18229
rect 5137 17993 5221 18229
rect 5457 17993 5541 18229
rect 5777 17993 5861 18229
rect 6097 17993 6181 18229
rect 6417 17993 6501 18229
rect 6737 17993 6821 18229
rect 7057 17993 7141 18229
rect 7377 17993 7461 18229
rect 7697 17993 7781 18229
rect 8017 17993 8101 18229
rect 8337 17993 8421 18229
rect 8657 17993 8741 18229
rect 8977 17993 9061 18229
rect 9297 17993 9600 18229
rect 0 17893 9600 17993
rect 0 17657 421 17893
rect 657 17657 741 17893
rect 977 17657 1061 17893
rect 1297 17657 1381 17893
rect 1617 17657 1701 17893
rect 1937 17657 2021 17893
rect 2257 17657 2341 17893
rect 2577 17657 2661 17893
rect 2897 17657 2981 17893
rect 3217 17657 3301 17893
rect 3537 17657 3621 17893
rect 3857 17657 3941 17893
rect 4177 17657 4261 17893
rect 4497 17657 4581 17893
rect 4817 17657 4901 17893
rect 5137 17657 5221 17893
rect 5457 17657 5541 17893
rect 5777 17657 5861 17893
rect 6097 17657 6181 17893
rect 6417 17657 6501 17893
rect 6737 17657 6821 17893
rect 7057 17657 7141 17893
rect 7377 17657 7461 17893
rect 7697 17657 7781 17893
rect 8017 17657 8101 17893
rect 8337 17657 8421 17893
rect 8657 17657 8741 17893
rect 8977 17657 9061 17893
rect 9297 17657 9600 17893
rect 0 17557 9600 17657
rect 0 17321 421 17557
rect 657 17321 741 17557
rect 977 17321 1061 17557
rect 1297 17321 1381 17557
rect 1617 17321 1701 17557
rect 1937 17321 2021 17557
rect 2257 17321 2341 17557
rect 2577 17321 2661 17557
rect 2897 17321 2981 17557
rect 3217 17321 3301 17557
rect 3537 17321 3621 17557
rect 3857 17321 3941 17557
rect 4177 17321 4261 17557
rect 4497 17321 4581 17557
rect 4817 17321 4901 17557
rect 5137 17321 5221 17557
rect 5457 17321 5541 17557
rect 5777 17321 5861 17557
rect 6097 17321 6181 17557
rect 6417 17321 6501 17557
rect 6737 17321 6821 17557
rect 7057 17321 7141 17557
rect 7377 17321 7461 17557
rect 7697 17321 7781 17557
rect 8017 17321 8101 17557
rect 8337 17321 8421 17557
rect 8657 17321 8741 17557
rect 8977 17321 9061 17557
rect 9297 17321 9600 17557
rect 0 17221 9600 17321
rect 0 16985 421 17221
rect 657 16985 741 17221
rect 977 16985 1061 17221
rect 1297 16985 1381 17221
rect 1617 16985 1701 17221
rect 1937 16985 2021 17221
rect 2257 16985 2341 17221
rect 2577 16985 2661 17221
rect 2897 16985 2981 17221
rect 3217 16985 3301 17221
rect 3537 16985 3621 17221
rect 3857 16985 3941 17221
rect 4177 16985 4261 17221
rect 4497 16985 4581 17221
rect 4817 16985 4901 17221
rect 5137 16985 5221 17221
rect 5457 16985 5541 17221
rect 5777 16985 5861 17221
rect 6097 16985 6181 17221
rect 6417 16985 6501 17221
rect 6737 16985 6821 17221
rect 7057 16985 7141 17221
rect 7377 16985 7461 17221
rect 7697 16985 7781 17221
rect 8017 16985 8101 17221
rect 8337 16985 8421 17221
rect 8657 16985 8741 17221
rect 8977 16985 9061 17221
rect 9297 16985 9600 17221
rect 0 16885 9600 16985
rect 0 16649 421 16885
rect 657 16649 741 16885
rect 977 16649 1061 16885
rect 1297 16649 1381 16885
rect 1617 16649 1701 16885
rect 1937 16649 2021 16885
rect 2257 16649 2341 16885
rect 2577 16649 2661 16885
rect 2897 16649 2981 16885
rect 3217 16649 3301 16885
rect 3537 16649 3621 16885
rect 3857 16649 3941 16885
rect 4177 16649 4261 16885
rect 4497 16649 4581 16885
rect 4817 16649 4901 16885
rect 5137 16649 5221 16885
rect 5457 16649 5541 16885
rect 5777 16649 5861 16885
rect 6097 16649 6181 16885
rect 6417 16649 6501 16885
rect 6737 16649 6821 16885
rect 7057 16649 7141 16885
rect 7377 16649 7461 16885
rect 7697 16649 7781 16885
rect 8017 16649 8101 16885
rect 8337 16649 8421 16885
rect 8657 16649 8741 16885
rect 8977 16649 9061 16885
rect 9297 16649 9600 16885
rect 0 16549 9600 16649
rect 0 16313 421 16549
rect 657 16313 741 16549
rect 977 16313 1061 16549
rect 1297 16313 1381 16549
rect 1617 16313 1701 16549
rect 1937 16313 2021 16549
rect 2257 16313 2341 16549
rect 2577 16313 2661 16549
rect 2897 16313 2981 16549
rect 3217 16313 3301 16549
rect 3537 16313 3621 16549
rect 3857 16313 3941 16549
rect 4177 16313 4261 16549
rect 4497 16313 4581 16549
rect 4817 16313 4901 16549
rect 5137 16313 5221 16549
rect 5457 16313 5541 16549
rect 5777 16313 5861 16549
rect 6097 16313 6181 16549
rect 6417 16313 6501 16549
rect 6737 16313 6821 16549
rect 7057 16313 7141 16549
rect 7377 16313 7461 16549
rect 7697 16313 7781 16549
rect 8017 16313 8101 16549
rect 8337 16313 8421 16549
rect 8657 16313 8741 16549
rect 8977 16313 9061 16549
rect 9297 16313 9600 16549
rect 0 16213 9600 16313
rect 0 15977 421 16213
rect 657 15977 741 16213
rect 977 15977 1061 16213
rect 1297 15977 1381 16213
rect 1617 15977 1701 16213
rect 1937 15977 2021 16213
rect 2257 15977 2341 16213
rect 2577 15977 2661 16213
rect 2897 15977 2981 16213
rect 3217 15977 3301 16213
rect 3537 15977 3621 16213
rect 3857 15977 3941 16213
rect 4177 15977 4261 16213
rect 4497 15977 4581 16213
rect 4817 15977 4901 16213
rect 5137 15977 5221 16213
rect 5457 15977 5541 16213
rect 5777 15977 5861 16213
rect 6097 15977 6181 16213
rect 6417 15977 6501 16213
rect 6737 15977 6821 16213
rect 7057 15977 7141 16213
rect 7377 15977 7461 16213
rect 7697 15977 7781 16213
rect 8017 15977 8101 16213
rect 8337 15977 8421 16213
rect 8657 15977 8741 16213
rect 8977 15977 9061 16213
rect 9297 15977 9600 16213
rect 0 15877 9600 15977
rect 0 15641 421 15877
rect 657 15641 741 15877
rect 977 15641 1061 15877
rect 1297 15641 1381 15877
rect 1617 15641 1701 15877
rect 1937 15641 2021 15877
rect 2257 15641 2341 15877
rect 2577 15641 2661 15877
rect 2897 15641 2981 15877
rect 3217 15641 3301 15877
rect 3537 15641 3621 15877
rect 3857 15641 3941 15877
rect 4177 15641 4261 15877
rect 4497 15641 4581 15877
rect 4817 15641 4901 15877
rect 5137 15641 5221 15877
rect 5457 15641 5541 15877
rect 5777 15641 5861 15877
rect 6097 15641 6181 15877
rect 6417 15641 6501 15877
rect 6737 15641 6821 15877
rect 7057 15641 7141 15877
rect 7377 15641 7461 15877
rect 7697 15641 7781 15877
rect 8017 15641 8101 15877
rect 8337 15641 8421 15877
rect 8657 15641 8741 15877
rect 8977 15641 9061 15877
rect 9297 15641 9600 15877
rect 0 15541 9600 15641
rect 0 15305 421 15541
rect 657 15305 741 15541
rect 977 15305 1061 15541
rect 1297 15305 1381 15541
rect 1617 15305 1701 15541
rect 1937 15305 2021 15541
rect 2257 15305 2341 15541
rect 2577 15305 2661 15541
rect 2897 15305 2981 15541
rect 3217 15305 3301 15541
rect 3537 15305 3621 15541
rect 3857 15305 3941 15541
rect 4177 15305 4261 15541
rect 4497 15305 4581 15541
rect 4817 15305 4901 15541
rect 5137 15305 5221 15541
rect 5457 15305 5541 15541
rect 5777 15305 5861 15541
rect 6097 15305 6181 15541
rect 6417 15305 6501 15541
rect 6737 15305 6821 15541
rect 7057 15305 7141 15541
rect 7377 15305 7461 15541
rect 7697 15305 7781 15541
rect 8017 15305 8101 15541
rect 8337 15305 8421 15541
rect 8657 15305 8741 15541
rect 8977 15305 9061 15541
rect 9297 15305 9600 15541
rect 0 15205 9600 15305
rect 0 14969 421 15205
rect 657 14969 741 15205
rect 977 14969 1061 15205
rect 1297 14969 1381 15205
rect 1617 14969 1701 15205
rect 1937 14969 2021 15205
rect 2257 14969 2341 15205
rect 2577 14969 2661 15205
rect 2897 14969 2981 15205
rect 3217 14969 3301 15205
rect 3537 14969 3621 15205
rect 3857 14969 3941 15205
rect 4177 14969 4261 15205
rect 4497 14969 4581 15205
rect 4817 14969 4901 15205
rect 5137 14969 5221 15205
rect 5457 14969 5541 15205
rect 5777 14969 5861 15205
rect 6097 14969 6181 15205
rect 6417 14969 6501 15205
rect 6737 14969 6821 15205
rect 7057 14969 7141 15205
rect 7377 14969 7461 15205
rect 7697 14969 7781 15205
rect 8017 14969 8101 15205
rect 8337 14969 8421 15205
rect 8657 14969 8741 15205
rect 8977 14969 9061 15205
rect 9297 14969 9600 15205
rect 0 14869 9600 14969
rect 0 14633 421 14869
rect 657 14633 741 14869
rect 977 14633 1061 14869
rect 1297 14633 1381 14869
rect 1617 14633 1701 14869
rect 1937 14633 2021 14869
rect 2257 14633 2341 14869
rect 2577 14633 2661 14869
rect 2897 14633 2981 14869
rect 3217 14633 3301 14869
rect 3537 14633 3621 14869
rect 3857 14633 3941 14869
rect 4177 14633 4261 14869
rect 4497 14633 4581 14869
rect 4817 14633 4901 14869
rect 5137 14633 5221 14869
rect 5457 14633 5541 14869
rect 5777 14633 5861 14869
rect 6097 14633 6181 14869
rect 6417 14633 6501 14869
rect 6737 14633 6821 14869
rect 7057 14633 7141 14869
rect 7377 14633 7461 14869
rect 7697 14633 7781 14869
rect 8017 14633 8101 14869
rect 8337 14633 8421 14869
rect 8657 14633 8741 14869
rect 8977 14633 9061 14869
rect 9297 14633 9600 14869
rect 0 14533 9600 14633
rect 0 14297 421 14533
rect 657 14297 741 14533
rect 977 14297 1061 14533
rect 1297 14297 1381 14533
rect 1617 14297 1701 14533
rect 1937 14297 2021 14533
rect 2257 14297 2341 14533
rect 2577 14297 2661 14533
rect 2897 14297 2981 14533
rect 3217 14297 3301 14533
rect 3537 14297 3621 14533
rect 3857 14297 3941 14533
rect 4177 14297 4261 14533
rect 4497 14297 4581 14533
rect 4817 14297 4901 14533
rect 5137 14297 5221 14533
rect 5457 14297 5541 14533
rect 5777 14297 5861 14533
rect 6097 14297 6181 14533
rect 6417 14297 6501 14533
rect 6737 14297 6821 14533
rect 7057 14297 7141 14533
rect 7377 14297 7461 14533
rect 7697 14297 7781 14533
rect 8017 14297 8101 14533
rect 8337 14297 8421 14533
rect 8657 14297 8741 14533
rect 8977 14297 9061 14533
rect 9297 14297 9600 14533
rect 0 14197 9600 14297
rect 0 13961 421 14197
rect 657 13961 741 14197
rect 977 13961 1061 14197
rect 1297 13961 1381 14197
rect 1617 13961 1701 14197
rect 1937 13961 2021 14197
rect 2257 13961 2341 14197
rect 2577 13961 2661 14197
rect 2897 13961 2981 14197
rect 3217 13961 3301 14197
rect 3537 13961 3621 14197
rect 3857 13961 3941 14197
rect 4177 13961 4261 14197
rect 4497 13961 4581 14197
rect 4817 13961 4901 14197
rect 5137 13961 5221 14197
rect 5457 13961 5541 14197
rect 5777 13961 5861 14197
rect 6097 13961 6181 14197
rect 6417 13961 6501 14197
rect 6737 13961 6821 14197
rect 7057 13961 7141 14197
rect 7377 13961 7461 14197
rect 7697 13961 7781 14197
rect 8017 13961 8101 14197
rect 8337 13961 8421 14197
rect 8657 13961 8741 14197
rect 8977 13961 9061 14197
rect 9297 13961 9600 14197
rect 0 13861 9600 13961
rect 0 13625 421 13861
rect 657 13625 741 13861
rect 977 13625 1061 13861
rect 1297 13625 1381 13861
rect 1617 13625 1701 13861
rect 1937 13625 2021 13861
rect 2257 13625 2341 13861
rect 2577 13625 2661 13861
rect 2897 13625 2981 13861
rect 3217 13625 3301 13861
rect 3537 13625 3621 13861
rect 3857 13625 3941 13861
rect 4177 13625 4261 13861
rect 4497 13625 4581 13861
rect 4817 13625 4901 13861
rect 5137 13625 5221 13861
rect 5457 13625 5541 13861
rect 5777 13625 5861 13861
rect 6097 13625 6181 13861
rect 6417 13625 6501 13861
rect 6737 13625 6821 13861
rect 7057 13625 7141 13861
rect 7377 13625 7461 13861
rect 7697 13625 7781 13861
rect 8017 13625 8101 13861
rect 8337 13625 8421 13861
rect 8657 13625 8741 13861
rect 8977 13625 9061 13861
rect 9297 13625 9600 13861
rect 0 13600 9600 13625
rect 0 13256 9600 13300
rect 0 13020 422 13256
rect 658 13020 742 13256
rect 978 13020 1062 13256
rect 1298 13020 1382 13256
rect 1618 13020 1702 13256
rect 1938 13020 2022 13256
rect 2258 13020 2342 13256
rect 2578 13020 2662 13256
rect 2898 13020 2982 13256
rect 3218 13020 3302 13256
rect 3538 13020 3622 13256
rect 3858 13020 3942 13256
rect 4178 13020 4262 13256
rect 4498 13020 4582 13256
rect 4818 13020 4902 13256
rect 5138 13020 5222 13256
rect 5458 13020 5542 13256
rect 5778 13020 5862 13256
rect 6098 13020 6182 13256
rect 6418 13020 6502 13256
rect 6738 13020 6822 13256
rect 7058 13020 7142 13256
rect 7378 13020 7462 13256
rect 7698 13020 7782 13256
rect 8018 13020 8102 13256
rect 8338 13020 8422 13256
rect 8658 13020 8742 13256
rect 8978 13020 9062 13256
rect 9298 13020 9600 13256
rect 0 12690 9600 13020
rect 0 12454 422 12690
rect 658 12454 742 12690
rect 978 12454 1062 12690
rect 1298 12454 1382 12690
rect 1618 12454 1702 12690
rect 1938 12454 2022 12690
rect 2258 12454 2342 12690
rect 2578 12454 2662 12690
rect 2898 12454 2982 12690
rect 3218 12454 3302 12690
rect 3538 12454 3622 12690
rect 3858 12454 3942 12690
rect 4178 12454 4262 12690
rect 4498 12454 4582 12690
rect 4818 12454 4902 12690
rect 5138 12454 5222 12690
rect 5458 12454 5542 12690
rect 5778 12454 5862 12690
rect 6098 12454 6182 12690
rect 6418 12454 6502 12690
rect 6738 12454 6822 12690
rect 7058 12454 7142 12690
rect 7378 12454 7462 12690
rect 7698 12454 7782 12690
rect 8018 12454 8102 12690
rect 8338 12454 8422 12690
rect 8658 12454 8742 12690
rect 8978 12454 9062 12690
rect 9298 12454 9600 12690
rect 0 12410 9600 12454
rect 0 12086 9600 12130
rect 0 11850 422 12086
rect 658 11850 742 12086
rect 978 11850 1062 12086
rect 1298 11850 1382 12086
rect 1618 11850 1702 12086
rect 1938 11850 2022 12086
rect 2258 11850 2342 12086
rect 2578 11850 2662 12086
rect 2898 11850 2982 12086
rect 3218 11850 3302 12086
rect 3538 11850 3622 12086
rect 3858 11850 3942 12086
rect 4178 11850 4262 12086
rect 4498 11850 4582 12086
rect 4818 11850 4902 12086
rect 5138 11850 5222 12086
rect 5458 11850 5542 12086
rect 5778 11850 5862 12086
rect 6098 11850 6182 12086
rect 6418 11850 6502 12086
rect 6738 11850 6822 12086
rect 7058 11850 7142 12086
rect 7378 11850 7462 12086
rect 7698 11850 7782 12086
rect 8018 11850 8102 12086
rect 8338 11850 8422 12086
rect 8658 11850 8742 12086
rect 8978 11850 9062 12086
rect 9298 11850 9600 12086
rect 0 11520 9600 11850
rect 0 11284 422 11520
rect 658 11284 742 11520
rect 978 11284 1062 11520
rect 1298 11284 1382 11520
rect 1618 11284 1702 11520
rect 1938 11284 2022 11520
rect 2258 11284 2342 11520
rect 2578 11284 2662 11520
rect 2898 11284 2982 11520
rect 3218 11284 3302 11520
rect 3538 11284 3622 11520
rect 3858 11284 3942 11520
rect 4178 11284 4262 11520
rect 4498 11284 4582 11520
rect 4818 11284 4902 11520
rect 5138 11284 5222 11520
rect 5458 11284 5542 11520
rect 5778 11284 5862 11520
rect 6098 11284 6182 11520
rect 6418 11284 6502 11520
rect 6738 11284 6822 11520
rect 7058 11284 7142 11520
rect 7378 11284 7462 11520
rect 7698 11284 7782 11520
rect 8018 11284 8102 11520
rect 8338 11284 8422 11520
rect 8658 11284 8742 11520
rect 8978 11284 9062 11520
rect 9298 11284 9600 11520
rect 0 11240 9600 11284
rect 0 10874 9600 10940
rect 0 10218 3500 10814
rect 5889 10218 9600 10814
rect 0 9922 422 10158
rect 658 9922 742 10158
rect 978 9922 1062 10158
rect 1298 9922 1382 10158
rect 1618 9922 1702 10158
rect 1938 9922 2022 10158
rect 2258 9922 2342 10158
rect 2578 9922 2662 10158
rect 2898 9922 2982 10158
rect 3218 9922 3302 10158
rect 3538 9922 3622 10158
rect 3858 9922 3942 10158
rect 4178 9922 4262 10158
rect 4498 9922 4582 10158
rect 4818 9922 4902 10158
rect 5138 9922 5222 10158
rect 5458 9922 5542 10158
rect 5778 9922 5862 10158
rect 6098 9922 6182 10158
rect 6418 9922 6502 10158
rect 6738 9922 6822 10158
rect 7058 9922 7142 10158
rect 7378 9922 7462 10158
rect 7698 9922 7782 10158
rect 8018 9922 8102 10158
rect 8338 9922 8422 10158
rect 8658 9922 8742 10158
rect 8978 9922 9062 10158
rect 9298 9922 9600 10158
rect 0 9266 3500 9862
rect 5889 9266 9600 9862
rect 0 9140 9600 9206
rect 0 8796 9600 8840
rect 0 8560 422 8796
rect 658 8560 742 8796
rect 978 8560 1062 8796
rect 1298 8560 1382 8796
rect 1618 8560 1702 8796
rect 1938 8560 2022 8796
rect 2258 8560 2342 8796
rect 2578 8560 2662 8796
rect 2898 8560 2982 8796
rect 3218 8560 3302 8796
rect 3538 8560 3622 8796
rect 3858 8560 3942 8796
rect 4178 8560 4262 8796
rect 4498 8560 4582 8796
rect 4818 8560 4902 8796
rect 5138 8560 5222 8796
rect 5458 8560 5542 8796
rect 5778 8560 5862 8796
rect 6098 8560 6182 8796
rect 6418 8560 6502 8796
rect 6738 8560 6822 8796
rect 7058 8560 7142 8796
rect 7378 8560 7462 8796
rect 7698 8560 7782 8796
rect 8018 8560 8102 8796
rect 8338 8560 8422 8796
rect 8658 8560 8742 8796
rect 8978 8560 9062 8796
rect 9298 8560 9600 8796
rect 0 8190 9600 8560
rect 0 7954 422 8190
rect 658 7954 742 8190
rect 978 7954 1062 8190
rect 1298 7954 1382 8190
rect 1618 7954 1702 8190
rect 1938 7954 2022 8190
rect 2258 7954 2342 8190
rect 2578 7954 2662 8190
rect 2898 7954 2982 8190
rect 3218 7954 3302 8190
rect 3538 7954 3622 8190
rect 3858 7954 3942 8190
rect 4178 7954 4262 8190
rect 4498 7954 4582 8190
rect 4818 7954 4902 8190
rect 5138 7954 5222 8190
rect 5458 7954 5542 8190
rect 5778 7954 5862 8190
rect 6098 7954 6182 8190
rect 6418 7954 6502 8190
rect 6738 7954 6822 8190
rect 7058 7954 7142 8190
rect 7378 7954 7462 8190
rect 7698 7954 7782 8190
rect 8018 7954 8102 8190
rect 8338 7954 8422 8190
rect 8658 7954 8742 8190
rect 8978 7954 9062 8190
rect 9298 7954 9600 8190
rect 0 7910 9600 7954
rect 0 7586 9600 7630
rect 0 7350 422 7586
rect 658 7350 742 7586
rect 978 7350 1062 7586
rect 1298 7350 1382 7586
rect 1618 7350 1702 7586
rect 1938 7350 2022 7586
rect 2258 7350 2342 7586
rect 2578 7350 2662 7586
rect 2898 7350 2982 7586
rect 3218 7350 3302 7586
rect 3538 7350 3622 7586
rect 3858 7350 3942 7586
rect 4178 7350 4262 7586
rect 4498 7350 4582 7586
rect 4818 7350 4902 7586
rect 5138 7350 5222 7586
rect 5458 7350 5542 7586
rect 5778 7350 5862 7586
rect 6098 7350 6182 7586
rect 6418 7350 6502 7586
rect 6738 7350 6822 7586
rect 7058 7350 7142 7586
rect 7378 7350 7462 7586
rect 7698 7350 7782 7586
rect 8018 7350 8102 7586
rect 8338 7350 8422 7586
rect 8658 7350 8742 7586
rect 8978 7350 9062 7586
rect 9298 7350 9600 7586
rect 0 7220 9600 7350
rect 0 6984 422 7220
rect 658 6984 742 7220
rect 978 6984 1062 7220
rect 1298 6984 1382 7220
rect 1618 6984 1702 7220
rect 1938 6984 2022 7220
rect 2258 6984 2342 7220
rect 2578 6984 2662 7220
rect 2898 6984 2982 7220
rect 3218 6984 3302 7220
rect 3538 6984 3622 7220
rect 3858 6984 3942 7220
rect 4178 6984 4262 7220
rect 4498 6984 4582 7220
rect 4818 6984 4902 7220
rect 5138 6984 5222 7220
rect 5458 6984 5542 7220
rect 5778 6984 5862 7220
rect 6098 6984 6182 7220
rect 6418 6984 6502 7220
rect 6738 6984 6822 7220
rect 7058 6984 7142 7220
rect 7378 6984 7462 7220
rect 7698 6984 7782 7220
rect 8018 6984 8102 7220
rect 8338 6984 8422 7220
rect 8658 6984 8742 7220
rect 8978 6984 9062 7220
rect 9298 6984 9600 7220
rect 0 6940 9600 6984
rect 0 6616 9600 6660
rect 0 6380 422 6616
rect 658 6380 742 6616
rect 978 6380 1062 6616
rect 1298 6380 1382 6616
rect 1618 6380 1702 6616
rect 1938 6380 2022 6616
rect 2258 6380 2342 6616
rect 2578 6380 2662 6616
rect 2898 6380 2982 6616
rect 3218 6380 3302 6616
rect 3538 6380 3622 6616
rect 3858 6380 3942 6616
rect 4178 6380 4262 6616
rect 4498 6380 4582 6616
rect 4818 6380 4902 6616
rect 5138 6380 5222 6616
rect 5458 6380 5542 6616
rect 5778 6380 5862 6616
rect 6098 6380 6182 6616
rect 6418 6380 6502 6616
rect 6738 6380 6822 6616
rect 7058 6380 7142 6616
rect 7378 6380 7462 6616
rect 7698 6380 7782 6616
rect 8018 6380 8102 6616
rect 8338 6380 8422 6616
rect 8658 6380 8742 6616
rect 8978 6380 9062 6616
rect 9298 6380 9600 6616
rect 0 6250 9600 6380
rect 0 6014 422 6250
rect 658 6014 742 6250
rect 978 6014 1062 6250
rect 1298 6014 1382 6250
rect 1618 6014 1702 6250
rect 1938 6014 2022 6250
rect 2258 6014 2342 6250
rect 2578 6014 2662 6250
rect 2898 6014 2982 6250
rect 3218 6014 3302 6250
rect 3538 6014 3622 6250
rect 3858 6014 3942 6250
rect 4178 6014 4262 6250
rect 4498 6014 4582 6250
rect 4818 6014 4902 6250
rect 5138 6014 5222 6250
rect 5458 6014 5542 6250
rect 5778 6014 5862 6250
rect 6098 6014 6182 6250
rect 6418 6014 6502 6250
rect 6738 6014 6822 6250
rect 7058 6014 7142 6250
rect 7378 6014 7462 6250
rect 7698 6014 7782 6250
rect 8018 6014 8102 6250
rect 8338 6014 8422 6250
rect 8658 6014 8742 6250
rect 8978 6014 9062 6250
rect 9298 6014 9600 6250
rect 0 5970 9600 6014
rect 0 5646 9600 5690
rect 0 5410 422 5646
rect 658 5410 742 5646
rect 978 5410 1062 5646
rect 1298 5410 1382 5646
rect 1618 5410 1702 5646
rect 1938 5410 2022 5646
rect 2258 5410 2342 5646
rect 2578 5410 2662 5646
rect 2898 5410 2982 5646
rect 3218 5410 3302 5646
rect 3538 5410 3622 5646
rect 3858 5410 3942 5646
rect 4178 5410 4262 5646
rect 4498 5410 4582 5646
rect 4818 5410 4902 5646
rect 5138 5410 5222 5646
rect 5458 5410 5542 5646
rect 5778 5410 5862 5646
rect 6098 5410 6182 5646
rect 6418 5410 6502 5646
rect 6738 5410 6822 5646
rect 7058 5410 7142 5646
rect 7378 5410 7462 5646
rect 7698 5410 7782 5646
rect 8018 5410 8102 5646
rect 8338 5410 8422 5646
rect 8658 5410 8742 5646
rect 8978 5410 9062 5646
rect 9298 5410 9600 5646
rect 0 5040 9600 5410
rect 0 4804 422 5040
rect 658 4804 742 5040
rect 978 4804 1062 5040
rect 1298 4804 1382 5040
rect 1618 4804 1702 5040
rect 1938 4804 2022 5040
rect 2258 4804 2342 5040
rect 2578 4804 2662 5040
rect 2898 4804 2982 5040
rect 3218 4804 3302 5040
rect 3538 4804 3622 5040
rect 3858 4804 3942 5040
rect 4178 4804 4262 5040
rect 4498 4804 4582 5040
rect 4818 4804 4902 5040
rect 5138 4804 5222 5040
rect 5458 4804 5542 5040
rect 5778 4804 5862 5040
rect 6098 4804 6182 5040
rect 6418 4804 6502 5040
rect 6738 4804 6822 5040
rect 7058 4804 7142 5040
rect 7378 4804 7462 5040
rect 7698 4804 7782 5040
rect 8018 4804 8102 5040
rect 8338 4804 8422 5040
rect 8658 4804 8742 5040
rect 8978 4804 9062 5040
rect 9298 4804 9600 5040
rect 0 4760 9600 4804
rect 0 4436 9600 4480
rect 0 4200 422 4436
rect 658 4200 742 4436
rect 978 4200 1062 4436
rect 1298 4200 1382 4436
rect 1618 4200 1702 4436
rect 1938 4200 2022 4436
rect 2258 4200 2342 4436
rect 2578 4200 2662 4436
rect 2898 4200 2982 4436
rect 3218 4200 3302 4436
rect 3538 4200 3622 4436
rect 3858 4200 3942 4436
rect 4178 4200 4262 4436
rect 4498 4200 4582 4436
rect 4818 4200 4902 4436
rect 5138 4200 5222 4436
rect 5458 4200 5542 4436
rect 5778 4200 5862 4436
rect 6098 4200 6182 4436
rect 6418 4200 6502 4436
rect 6738 4200 6822 4436
rect 7058 4200 7142 4436
rect 7378 4200 7462 4436
rect 7698 4200 7782 4436
rect 8018 4200 8102 4436
rect 8338 4200 8422 4436
rect 8658 4200 8742 4436
rect 8978 4200 9062 4436
rect 9298 4200 9600 4436
rect 0 3830 9600 4200
rect 0 3594 422 3830
rect 658 3594 742 3830
rect 978 3594 1062 3830
rect 1298 3594 1382 3830
rect 1618 3594 1702 3830
rect 1938 3594 2022 3830
rect 2258 3594 2342 3830
rect 2578 3594 2662 3830
rect 2898 3594 2982 3830
rect 3218 3594 3302 3830
rect 3538 3594 3622 3830
rect 3858 3594 3942 3830
rect 4178 3594 4262 3830
rect 4498 3594 4582 3830
rect 4818 3594 4902 3830
rect 5138 3594 5222 3830
rect 5458 3594 5542 3830
rect 5778 3594 5862 3830
rect 6098 3594 6182 3830
rect 6418 3594 6502 3830
rect 6738 3594 6822 3830
rect 7058 3594 7142 3830
rect 7378 3594 7462 3830
rect 7698 3594 7782 3830
rect 8018 3594 8102 3830
rect 8338 3594 8422 3830
rect 8658 3594 8742 3830
rect 8978 3594 9062 3830
rect 9298 3594 9600 3830
rect 0 3550 9600 3594
rect 0 3226 9600 3270
rect 0 2990 422 3226
rect 658 2990 742 3226
rect 978 2990 1062 3226
rect 1298 2990 1382 3226
rect 1618 2990 1702 3226
rect 1938 2990 2022 3226
rect 2258 2990 2342 3226
rect 2578 2990 2662 3226
rect 2898 2990 2982 3226
rect 3218 2990 3302 3226
rect 3538 2990 3622 3226
rect 3858 2990 3942 3226
rect 4178 2990 4262 3226
rect 4498 2990 4582 3226
rect 4818 2990 4902 3226
rect 5138 2990 5222 3226
rect 5458 2990 5542 3226
rect 5778 2990 5862 3226
rect 6098 2990 6182 3226
rect 6418 2990 6502 3226
rect 6738 2990 6822 3226
rect 7058 2990 7142 3226
rect 7378 2990 7462 3226
rect 7698 2990 7782 3226
rect 8018 2990 8102 3226
rect 8338 2990 8422 3226
rect 8658 2990 8742 3226
rect 8978 2990 9062 3226
rect 9298 2990 9600 3226
rect 0 2860 9600 2990
rect 0 2624 422 2860
rect 658 2624 742 2860
rect 978 2624 1062 2860
rect 1298 2624 1382 2860
rect 1618 2624 1702 2860
rect 1938 2624 2022 2860
rect 2258 2624 2342 2860
rect 2578 2624 2662 2860
rect 2898 2624 2982 2860
rect 3218 2624 3302 2860
rect 3538 2624 3622 2860
rect 3858 2624 3942 2860
rect 4178 2624 4262 2860
rect 4498 2624 4582 2860
rect 4818 2624 4902 2860
rect 5138 2624 5222 2860
rect 5458 2624 5542 2860
rect 5778 2624 5862 2860
rect 6098 2624 6182 2860
rect 6418 2624 6502 2860
rect 6738 2624 6822 2860
rect 7058 2624 7142 2860
rect 7378 2624 7462 2860
rect 7698 2624 7782 2860
rect 8018 2624 8102 2860
rect 8338 2624 8422 2860
rect 8658 2624 8742 2860
rect 8978 2624 9062 2860
rect 9298 2624 9600 2860
rect 0 2580 9600 2624
rect 0 2256 9600 2300
rect 0 2020 422 2256
rect 658 2020 742 2256
rect 978 2020 1062 2256
rect 1298 2020 1382 2256
rect 1618 2020 1702 2256
rect 1938 2020 2022 2256
rect 2258 2020 2342 2256
rect 2578 2020 2662 2256
rect 2898 2020 2982 2256
rect 3218 2020 3302 2256
rect 3538 2020 3622 2256
rect 3858 2020 3942 2256
rect 4178 2020 4262 2256
rect 4498 2020 4582 2256
rect 4818 2020 4902 2256
rect 5138 2020 5222 2256
rect 5458 2020 5542 2256
rect 5778 2020 5862 2256
rect 6098 2020 6182 2256
rect 6418 2020 6502 2256
rect 6738 2020 6822 2256
rect 7058 2020 7142 2256
rect 7378 2020 7462 2256
rect 7698 2020 7782 2256
rect 8018 2020 8102 2256
rect 8338 2020 8422 2256
rect 8658 2020 8742 2256
rect 8978 2020 9062 2256
rect 9298 2020 9600 2256
rect 0 1650 9600 2020
rect 0 1414 422 1650
rect 658 1414 742 1650
rect 978 1414 1062 1650
rect 1298 1414 1382 1650
rect 1618 1414 1702 1650
rect 1938 1414 2022 1650
rect 2258 1414 2342 1650
rect 2578 1414 2662 1650
rect 2898 1414 2982 1650
rect 3218 1414 3302 1650
rect 3538 1414 3622 1650
rect 3858 1414 3942 1650
rect 4178 1414 4262 1650
rect 4498 1414 4582 1650
rect 4818 1414 4902 1650
rect 5138 1414 5222 1650
rect 5458 1414 5542 1650
rect 5778 1414 5862 1650
rect 6098 1414 6182 1650
rect 6418 1414 6502 1650
rect 6738 1414 6822 1650
rect 7058 1414 7142 1650
rect 7378 1414 7462 1650
rect 7698 1414 7782 1650
rect 8018 1414 8102 1650
rect 8338 1414 8422 1650
rect 8658 1414 8742 1650
rect 8978 1414 9062 1650
rect 9298 1414 9600 1650
rect 0 1370 9600 1414
rect 0 1045 9600 1090
rect 0 809 422 1045
rect 658 809 742 1045
rect 978 809 1062 1045
rect 1298 809 1382 1045
rect 1618 809 1702 1045
rect 1938 809 2022 1045
rect 2258 809 2342 1045
rect 2578 809 2662 1045
rect 2898 809 2982 1045
rect 3218 809 3302 1045
rect 3538 809 3622 1045
rect 3858 809 3942 1045
rect 4178 809 4262 1045
rect 4498 809 4582 1045
rect 4818 809 4902 1045
rect 5138 809 5222 1045
rect 5458 809 5542 1045
rect 5778 809 5862 1045
rect 6098 809 6182 1045
rect 6418 809 6502 1045
rect 6738 809 6822 1045
rect 7058 809 7142 1045
rect 7378 809 7462 1045
rect 7698 809 7782 1045
rect 8018 809 8102 1045
rect 8338 809 8422 1045
rect 8658 809 8742 1045
rect 8978 809 9062 1045
rect 9298 809 9600 1045
rect 0 663 9600 809
rect 0 427 422 663
rect 658 427 742 663
rect 978 427 1062 663
rect 1298 427 1382 663
rect 1618 427 1702 663
rect 1938 427 2022 663
rect 2258 427 2342 663
rect 2578 427 2662 663
rect 2898 427 2982 663
rect 3218 427 3302 663
rect 3538 427 3622 663
rect 3858 427 3942 663
rect 4178 427 4262 663
rect 4498 427 4582 663
rect 4818 427 4902 663
rect 5138 427 5222 663
rect 5458 427 5542 663
rect 5778 427 5862 663
rect 6098 427 6182 663
rect 6418 427 6502 663
rect 6738 427 6822 663
rect 7058 427 7142 663
rect 7378 427 7462 663
rect 7698 427 7782 663
rect 8018 427 8102 663
rect 8338 427 8422 663
rect 8658 427 8742 663
rect 8978 427 9062 663
rect 9298 427 9600 663
rect 0 281 9600 427
rect 0 45 422 281
rect 658 45 742 281
rect 978 45 1062 281
rect 1298 45 1382 281
rect 1618 45 1702 281
rect 1938 45 2022 281
rect 2258 45 2342 281
rect 2578 45 2662 281
rect 2898 45 2982 281
rect 3218 45 3302 281
rect 3538 45 3622 281
rect 3858 45 3942 281
rect 4178 45 4262 281
rect 4498 45 4582 281
rect 4818 45 4902 281
rect 5138 45 5222 281
rect 5458 45 5542 281
rect 5778 45 5862 281
rect 6098 45 6182 281
rect 6418 45 6502 281
rect 6738 45 6822 281
rect 7058 45 7142 281
rect 7378 45 7462 281
rect 7698 45 7782 281
rect 8018 45 8102 281
rect 8338 45 8422 281
rect 8658 45 8742 281
rect 8978 45 9062 281
rect 9298 45 9600 281
rect 0 0 9600 45
<< via4 >>
rect 422 34814 9298 39530
rect 421 18329 657 18565
rect 741 18329 977 18565
rect 1061 18329 1297 18565
rect 1381 18329 1617 18565
rect 1701 18329 1937 18565
rect 2021 18329 2257 18565
rect 2341 18329 2577 18565
rect 2661 18329 2897 18565
rect 2981 18329 3217 18565
rect 3301 18329 3537 18565
rect 3621 18329 3857 18565
rect 3941 18329 4177 18565
rect 4261 18329 4497 18565
rect 4581 18329 4817 18565
rect 4901 18329 5137 18565
rect 5221 18329 5457 18565
rect 5541 18329 5777 18565
rect 5861 18329 6097 18565
rect 6181 18329 6417 18565
rect 6501 18329 6737 18565
rect 6821 18329 7057 18565
rect 7141 18329 7377 18565
rect 7461 18329 7697 18565
rect 7781 18329 8017 18565
rect 8101 18329 8337 18565
rect 8421 18329 8657 18565
rect 8741 18329 8977 18565
rect 9061 18329 9297 18565
rect 421 17993 657 18229
rect 741 17993 977 18229
rect 1061 17993 1297 18229
rect 1381 17993 1617 18229
rect 1701 17993 1937 18229
rect 2021 17993 2257 18229
rect 2341 17993 2577 18229
rect 2661 17993 2897 18229
rect 2981 17993 3217 18229
rect 3301 17993 3537 18229
rect 3621 17993 3857 18229
rect 3941 17993 4177 18229
rect 4261 17993 4497 18229
rect 4581 17993 4817 18229
rect 4901 17993 5137 18229
rect 5221 17993 5457 18229
rect 5541 17993 5777 18229
rect 5861 17993 6097 18229
rect 6181 17993 6417 18229
rect 6501 17993 6737 18229
rect 6821 17993 7057 18229
rect 7141 17993 7377 18229
rect 7461 17993 7697 18229
rect 7781 17993 8017 18229
rect 8101 17993 8337 18229
rect 8421 17993 8657 18229
rect 8741 17993 8977 18229
rect 9061 17993 9297 18229
rect 421 17657 657 17893
rect 741 17657 977 17893
rect 1061 17657 1297 17893
rect 1381 17657 1617 17893
rect 1701 17657 1937 17893
rect 2021 17657 2257 17893
rect 2341 17657 2577 17893
rect 2661 17657 2897 17893
rect 2981 17657 3217 17893
rect 3301 17657 3537 17893
rect 3621 17657 3857 17893
rect 3941 17657 4177 17893
rect 4261 17657 4497 17893
rect 4581 17657 4817 17893
rect 4901 17657 5137 17893
rect 5221 17657 5457 17893
rect 5541 17657 5777 17893
rect 5861 17657 6097 17893
rect 6181 17657 6417 17893
rect 6501 17657 6737 17893
rect 6821 17657 7057 17893
rect 7141 17657 7377 17893
rect 7461 17657 7697 17893
rect 7781 17657 8017 17893
rect 8101 17657 8337 17893
rect 8421 17657 8657 17893
rect 8741 17657 8977 17893
rect 9061 17657 9297 17893
rect 421 17321 657 17557
rect 741 17321 977 17557
rect 1061 17321 1297 17557
rect 1381 17321 1617 17557
rect 1701 17321 1937 17557
rect 2021 17321 2257 17557
rect 2341 17321 2577 17557
rect 2661 17321 2897 17557
rect 2981 17321 3217 17557
rect 3301 17321 3537 17557
rect 3621 17321 3857 17557
rect 3941 17321 4177 17557
rect 4261 17321 4497 17557
rect 4581 17321 4817 17557
rect 4901 17321 5137 17557
rect 5221 17321 5457 17557
rect 5541 17321 5777 17557
rect 5861 17321 6097 17557
rect 6181 17321 6417 17557
rect 6501 17321 6737 17557
rect 6821 17321 7057 17557
rect 7141 17321 7377 17557
rect 7461 17321 7697 17557
rect 7781 17321 8017 17557
rect 8101 17321 8337 17557
rect 8421 17321 8657 17557
rect 8741 17321 8977 17557
rect 9061 17321 9297 17557
rect 421 16985 657 17221
rect 741 16985 977 17221
rect 1061 16985 1297 17221
rect 1381 16985 1617 17221
rect 1701 16985 1937 17221
rect 2021 16985 2257 17221
rect 2341 16985 2577 17221
rect 2661 16985 2897 17221
rect 2981 16985 3217 17221
rect 3301 16985 3537 17221
rect 3621 16985 3857 17221
rect 3941 16985 4177 17221
rect 4261 16985 4497 17221
rect 4581 16985 4817 17221
rect 4901 16985 5137 17221
rect 5221 16985 5457 17221
rect 5541 16985 5777 17221
rect 5861 16985 6097 17221
rect 6181 16985 6417 17221
rect 6501 16985 6737 17221
rect 6821 16985 7057 17221
rect 7141 16985 7377 17221
rect 7461 16985 7697 17221
rect 7781 16985 8017 17221
rect 8101 16985 8337 17221
rect 8421 16985 8657 17221
rect 8741 16985 8977 17221
rect 9061 16985 9297 17221
rect 421 16649 657 16885
rect 741 16649 977 16885
rect 1061 16649 1297 16885
rect 1381 16649 1617 16885
rect 1701 16649 1937 16885
rect 2021 16649 2257 16885
rect 2341 16649 2577 16885
rect 2661 16649 2897 16885
rect 2981 16649 3217 16885
rect 3301 16649 3537 16885
rect 3621 16649 3857 16885
rect 3941 16649 4177 16885
rect 4261 16649 4497 16885
rect 4581 16649 4817 16885
rect 4901 16649 5137 16885
rect 5221 16649 5457 16885
rect 5541 16649 5777 16885
rect 5861 16649 6097 16885
rect 6181 16649 6417 16885
rect 6501 16649 6737 16885
rect 6821 16649 7057 16885
rect 7141 16649 7377 16885
rect 7461 16649 7697 16885
rect 7781 16649 8017 16885
rect 8101 16649 8337 16885
rect 8421 16649 8657 16885
rect 8741 16649 8977 16885
rect 9061 16649 9297 16885
rect 421 16313 657 16549
rect 741 16313 977 16549
rect 1061 16313 1297 16549
rect 1381 16313 1617 16549
rect 1701 16313 1937 16549
rect 2021 16313 2257 16549
rect 2341 16313 2577 16549
rect 2661 16313 2897 16549
rect 2981 16313 3217 16549
rect 3301 16313 3537 16549
rect 3621 16313 3857 16549
rect 3941 16313 4177 16549
rect 4261 16313 4497 16549
rect 4581 16313 4817 16549
rect 4901 16313 5137 16549
rect 5221 16313 5457 16549
rect 5541 16313 5777 16549
rect 5861 16313 6097 16549
rect 6181 16313 6417 16549
rect 6501 16313 6737 16549
rect 6821 16313 7057 16549
rect 7141 16313 7377 16549
rect 7461 16313 7697 16549
rect 7781 16313 8017 16549
rect 8101 16313 8337 16549
rect 8421 16313 8657 16549
rect 8741 16313 8977 16549
rect 9061 16313 9297 16549
rect 421 15977 657 16213
rect 741 15977 977 16213
rect 1061 15977 1297 16213
rect 1381 15977 1617 16213
rect 1701 15977 1937 16213
rect 2021 15977 2257 16213
rect 2341 15977 2577 16213
rect 2661 15977 2897 16213
rect 2981 15977 3217 16213
rect 3301 15977 3537 16213
rect 3621 15977 3857 16213
rect 3941 15977 4177 16213
rect 4261 15977 4497 16213
rect 4581 15977 4817 16213
rect 4901 15977 5137 16213
rect 5221 15977 5457 16213
rect 5541 15977 5777 16213
rect 5861 15977 6097 16213
rect 6181 15977 6417 16213
rect 6501 15977 6737 16213
rect 6821 15977 7057 16213
rect 7141 15977 7377 16213
rect 7461 15977 7697 16213
rect 7781 15977 8017 16213
rect 8101 15977 8337 16213
rect 8421 15977 8657 16213
rect 8741 15977 8977 16213
rect 9061 15977 9297 16213
rect 421 15641 657 15877
rect 741 15641 977 15877
rect 1061 15641 1297 15877
rect 1381 15641 1617 15877
rect 1701 15641 1937 15877
rect 2021 15641 2257 15877
rect 2341 15641 2577 15877
rect 2661 15641 2897 15877
rect 2981 15641 3217 15877
rect 3301 15641 3537 15877
rect 3621 15641 3857 15877
rect 3941 15641 4177 15877
rect 4261 15641 4497 15877
rect 4581 15641 4817 15877
rect 4901 15641 5137 15877
rect 5221 15641 5457 15877
rect 5541 15641 5777 15877
rect 5861 15641 6097 15877
rect 6181 15641 6417 15877
rect 6501 15641 6737 15877
rect 6821 15641 7057 15877
rect 7141 15641 7377 15877
rect 7461 15641 7697 15877
rect 7781 15641 8017 15877
rect 8101 15641 8337 15877
rect 8421 15641 8657 15877
rect 8741 15641 8977 15877
rect 9061 15641 9297 15877
rect 421 15305 657 15541
rect 741 15305 977 15541
rect 1061 15305 1297 15541
rect 1381 15305 1617 15541
rect 1701 15305 1937 15541
rect 2021 15305 2257 15541
rect 2341 15305 2577 15541
rect 2661 15305 2897 15541
rect 2981 15305 3217 15541
rect 3301 15305 3537 15541
rect 3621 15305 3857 15541
rect 3941 15305 4177 15541
rect 4261 15305 4497 15541
rect 4581 15305 4817 15541
rect 4901 15305 5137 15541
rect 5221 15305 5457 15541
rect 5541 15305 5777 15541
rect 5861 15305 6097 15541
rect 6181 15305 6417 15541
rect 6501 15305 6737 15541
rect 6821 15305 7057 15541
rect 7141 15305 7377 15541
rect 7461 15305 7697 15541
rect 7781 15305 8017 15541
rect 8101 15305 8337 15541
rect 8421 15305 8657 15541
rect 8741 15305 8977 15541
rect 9061 15305 9297 15541
rect 421 14969 657 15205
rect 741 14969 977 15205
rect 1061 14969 1297 15205
rect 1381 14969 1617 15205
rect 1701 14969 1937 15205
rect 2021 14969 2257 15205
rect 2341 14969 2577 15205
rect 2661 14969 2897 15205
rect 2981 14969 3217 15205
rect 3301 14969 3537 15205
rect 3621 14969 3857 15205
rect 3941 14969 4177 15205
rect 4261 14969 4497 15205
rect 4581 14969 4817 15205
rect 4901 14969 5137 15205
rect 5221 14969 5457 15205
rect 5541 14969 5777 15205
rect 5861 14969 6097 15205
rect 6181 14969 6417 15205
rect 6501 14969 6737 15205
rect 6821 14969 7057 15205
rect 7141 14969 7377 15205
rect 7461 14969 7697 15205
rect 7781 14969 8017 15205
rect 8101 14969 8337 15205
rect 8421 14969 8657 15205
rect 8741 14969 8977 15205
rect 9061 14969 9297 15205
rect 421 14633 657 14869
rect 741 14633 977 14869
rect 1061 14633 1297 14869
rect 1381 14633 1617 14869
rect 1701 14633 1937 14869
rect 2021 14633 2257 14869
rect 2341 14633 2577 14869
rect 2661 14633 2897 14869
rect 2981 14633 3217 14869
rect 3301 14633 3537 14869
rect 3621 14633 3857 14869
rect 3941 14633 4177 14869
rect 4261 14633 4497 14869
rect 4581 14633 4817 14869
rect 4901 14633 5137 14869
rect 5221 14633 5457 14869
rect 5541 14633 5777 14869
rect 5861 14633 6097 14869
rect 6181 14633 6417 14869
rect 6501 14633 6737 14869
rect 6821 14633 7057 14869
rect 7141 14633 7377 14869
rect 7461 14633 7697 14869
rect 7781 14633 8017 14869
rect 8101 14633 8337 14869
rect 8421 14633 8657 14869
rect 8741 14633 8977 14869
rect 9061 14633 9297 14869
rect 421 14297 657 14533
rect 741 14297 977 14533
rect 1061 14297 1297 14533
rect 1381 14297 1617 14533
rect 1701 14297 1937 14533
rect 2021 14297 2257 14533
rect 2341 14297 2577 14533
rect 2661 14297 2897 14533
rect 2981 14297 3217 14533
rect 3301 14297 3537 14533
rect 3621 14297 3857 14533
rect 3941 14297 4177 14533
rect 4261 14297 4497 14533
rect 4581 14297 4817 14533
rect 4901 14297 5137 14533
rect 5221 14297 5457 14533
rect 5541 14297 5777 14533
rect 5861 14297 6097 14533
rect 6181 14297 6417 14533
rect 6501 14297 6737 14533
rect 6821 14297 7057 14533
rect 7141 14297 7377 14533
rect 7461 14297 7697 14533
rect 7781 14297 8017 14533
rect 8101 14297 8337 14533
rect 8421 14297 8657 14533
rect 8741 14297 8977 14533
rect 9061 14297 9297 14533
rect 421 13961 657 14197
rect 741 13961 977 14197
rect 1061 13961 1297 14197
rect 1381 13961 1617 14197
rect 1701 13961 1937 14197
rect 2021 13961 2257 14197
rect 2341 13961 2577 14197
rect 2661 13961 2897 14197
rect 2981 13961 3217 14197
rect 3301 13961 3537 14197
rect 3621 13961 3857 14197
rect 3941 13961 4177 14197
rect 4261 13961 4497 14197
rect 4581 13961 4817 14197
rect 4901 13961 5137 14197
rect 5221 13961 5457 14197
rect 5541 13961 5777 14197
rect 5861 13961 6097 14197
rect 6181 13961 6417 14197
rect 6501 13961 6737 14197
rect 6821 13961 7057 14197
rect 7141 13961 7377 14197
rect 7461 13961 7697 14197
rect 7781 13961 8017 14197
rect 8101 13961 8337 14197
rect 8421 13961 8657 14197
rect 8741 13961 8977 14197
rect 9061 13961 9297 14197
rect 421 13625 657 13861
rect 741 13625 977 13861
rect 1061 13625 1297 13861
rect 1381 13625 1617 13861
rect 1701 13625 1937 13861
rect 2021 13625 2257 13861
rect 2341 13625 2577 13861
rect 2661 13625 2897 13861
rect 2981 13625 3217 13861
rect 3301 13625 3537 13861
rect 3621 13625 3857 13861
rect 3941 13625 4177 13861
rect 4261 13625 4497 13861
rect 4581 13625 4817 13861
rect 4901 13625 5137 13861
rect 5221 13625 5457 13861
rect 5541 13625 5777 13861
rect 5861 13625 6097 13861
rect 6181 13625 6417 13861
rect 6501 13625 6737 13861
rect 6821 13625 7057 13861
rect 7141 13625 7377 13861
rect 7461 13625 7697 13861
rect 7781 13625 8017 13861
rect 8101 13625 8337 13861
rect 8421 13625 8657 13861
rect 8741 13625 8977 13861
rect 9061 13625 9297 13861
rect 422 13020 658 13256
rect 742 13020 978 13256
rect 1062 13020 1298 13256
rect 1382 13020 1618 13256
rect 1702 13020 1938 13256
rect 2022 13020 2258 13256
rect 2342 13020 2578 13256
rect 2662 13020 2898 13256
rect 2982 13020 3218 13256
rect 3302 13020 3538 13256
rect 3622 13020 3858 13256
rect 3942 13020 4178 13256
rect 4262 13020 4498 13256
rect 4582 13020 4818 13256
rect 4902 13020 5138 13256
rect 5222 13020 5458 13256
rect 5542 13020 5778 13256
rect 5862 13020 6098 13256
rect 6182 13020 6418 13256
rect 6502 13020 6738 13256
rect 6822 13020 7058 13256
rect 7142 13020 7378 13256
rect 7462 13020 7698 13256
rect 7782 13020 8018 13256
rect 8102 13020 8338 13256
rect 8422 13020 8658 13256
rect 8742 13020 8978 13256
rect 9062 13020 9298 13256
rect 422 12454 658 12690
rect 742 12454 978 12690
rect 1062 12454 1298 12690
rect 1382 12454 1618 12690
rect 1702 12454 1938 12690
rect 2022 12454 2258 12690
rect 2342 12454 2578 12690
rect 2662 12454 2898 12690
rect 2982 12454 3218 12690
rect 3302 12454 3538 12690
rect 3622 12454 3858 12690
rect 3942 12454 4178 12690
rect 4262 12454 4498 12690
rect 4582 12454 4818 12690
rect 4902 12454 5138 12690
rect 5222 12454 5458 12690
rect 5542 12454 5778 12690
rect 5862 12454 6098 12690
rect 6182 12454 6418 12690
rect 6502 12454 6738 12690
rect 6822 12454 7058 12690
rect 7142 12454 7378 12690
rect 7462 12454 7698 12690
rect 7782 12454 8018 12690
rect 8102 12454 8338 12690
rect 8422 12454 8658 12690
rect 8742 12454 8978 12690
rect 9062 12454 9298 12690
rect 422 11850 658 12086
rect 742 11850 978 12086
rect 1062 11850 1298 12086
rect 1382 11850 1618 12086
rect 1702 11850 1938 12086
rect 2022 11850 2258 12086
rect 2342 11850 2578 12086
rect 2662 11850 2898 12086
rect 2982 11850 3218 12086
rect 3302 11850 3538 12086
rect 3622 11850 3858 12086
rect 3942 11850 4178 12086
rect 4262 11850 4498 12086
rect 4582 11850 4818 12086
rect 4902 11850 5138 12086
rect 5222 11850 5458 12086
rect 5542 11850 5778 12086
rect 5862 11850 6098 12086
rect 6182 11850 6418 12086
rect 6502 11850 6738 12086
rect 6822 11850 7058 12086
rect 7142 11850 7378 12086
rect 7462 11850 7698 12086
rect 7782 11850 8018 12086
rect 8102 11850 8338 12086
rect 8422 11850 8658 12086
rect 8742 11850 8978 12086
rect 9062 11850 9298 12086
rect 422 11284 658 11520
rect 742 11284 978 11520
rect 1062 11284 1298 11520
rect 1382 11284 1618 11520
rect 1702 11284 1938 11520
rect 2022 11284 2258 11520
rect 2342 11284 2578 11520
rect 2662 11284 2898 11520
rect 2982 11284 3218 11520
rect 3302 11284 3538 11520
rect 3622 11284 3858 11520
rect 3942 11284 4178 11520
rect 4262 11284 4498 11520
rect 4582 11284 4818 11520
rect 4902 11284 5138 11520
rect 5222 11284 5458 11520
rect 5542 11284 5778 11520
rect 5862 11284 6098 11520
rect 6182 11284 6418 11520
rect 6502 11284 6738 11520
rect 6822 11284 7058 11520
rect 7142 11284 7378 11520
rect 7462 11284 7698 11520
rect 7782 11284 8018 11520
rect 8102 11284 8338 11520
rect 8422 11284 8658 11520
rect 8742 11284 8978 11520
rect 9062 11284 9298 11520
rect 422 9922 658 10158
rect 742 9922 978 10158
rect 1062 9922 1298 10158
rect 1382 9922 1618 10158
rect 1702 9922 1938 10158
rect 2022 9922 2258 10158
rect 2342 9922 2578 10158
rect 2662 9922 2898 10158
rect 2982 9922 3218 10158
rect 3302 9922 3538 10158
rect 3622 9922 3858 10158
rect 3942 9922 4178 10158
rect 4262 9922 4498 10158
rect 4582 9922 4818 10158
rect 4902 9922 5138 10158
rect 5222 9922 5458 10158
rect 5542 9922 5778 10158
rect 5862 9922 6098 10158
rect 6182 9922 6418 10158
rect 6502 9922 6738 10158
rect 6822 9922 7058 10158
rect 7142 9922 7378 10158
rect 7462 9922 7698 10158
rect 7782 9922 8018 10158
rect 8102 9922 8338 10158
rect 8422 9922 8658 10158
rect 8742 9922 8978 10158
rect 9062 9922 9298 10158
rect 422 8560 658 8796
rect 742 8560 978 8796
rect 1062 8560 1298 8796
rect 1382 8560 1618 8796
rect 1702 8560 1938 8796
rect 2022 8560 2258 8796
rect 2342 8560 2578 8796
rect 2662 8560 2898 8796
rect 2982 8560 3218 8796
rect 3302 8560 3538 8796
rect 3622 8560 3858 8796
rect 3942 8560 4178 8796
rect 4262 8560 4498 8796
rect 4582 8560 4818 8796
rect 4902 8560 5138 8796
rect 5222 8560 5458 8796
rect 5542 8560 5778 8796
rect 5862 8560 6098 8796
rect 6182 8560 6418 8796
rect 6502 8560 6738 8796
rect 6822 8560 7058 8796
rect 7142 8560 7378 8796
rect 7462 8560 7698 8796
rect 7782 8560 8018 8796
rect 8102 8560 8338 8796
rect 8422 8560 8658 8796
rect 8742 8560 8978 8796
rect 9062 8560 9298 8796
rect 422 7954 658 8190
rect 742 7954 978 8190
rect 1062 7954 1298 8190
rect 1382 7954 1618 8190
rect 1702 7954 1938 8190
rect 2022 7954 2258 8190
rect 2342 7954 2578 8190
rect 2662 7954 2898 8190
rect 2982 7954 3218 8190
rect 3302 7954 3538 8190
rect 3622 7954 3858 8190
rect 3942 7954 4178 8190
rect 4262 7954 4498 8190
rect 4582 7954 4818 8190
rect 4902 7954 5138 8190
rect 5222 7954 5458 8190
rect 5542 7954 5778 8190
rect 5862 7954 6098 8190
rect 6182 7954 6418 8190
rect 6502 7954 6738 8190
rect 6822 7954 7058 8190
rect 7142 7954 7378 8190
rect 7462 7954 7698 8190
rect 7782 7954 8018 8190
rect 8102 7954 8338 8190
rect 8422 7954 8658 8190
rect 8742 7954 8978 8190
rect 9062 7954 9298 8190
rect 422 7350 658 7586
rect 742 7350 978 7586
rect 1062 7350 1298 7586
rect 1382 7350 1618 7586
rect 1702 7350 1938 7586
rect 2022 7350 2258 7586
rect 2342 7350 2578 7586
rect 2662 7350 2898 7586
rect 2982 7350 3218 7586
rect 3302 7350 3538 7586
rect 3622 7350 3858 7586
rect 3942 7350 4178 7586
rect 4262 7350 4498 7586
rect 4582 7350 4818 7586
rect 4902 7350 5138 7586
rect 5222 7350 5458 7586
rect 5542 7350 5778 7586
rect 5862 7350 6098 7586
rect 6182 7350 6418 7586
rect 6502 7350 6738 7586
rect 6822 7350 7058 7586
rect 7142 7350 7378 7586
rect 7462 7350 7698 7586
rect 7782 7350 8018 7586
rect 8102 7350 8338 7586
rect 8422 7350 8658 7586
rect 8742 7350 8978 7586
rect 9062 7350 9298 7586
rect 422 6984 658 7220
rect 742 6984 978 7220
rect 1062 6984 1298 7220
rect 1382 6984 1618 7220
rect 1702 6984 1938 7220
rect 2022 6984 2258 7220
rect 2342 6984 2578 7220
rect 2662 6984 2898 7220
rect 2982 6984 3218 7220
rect 3302 6984 3538 7220
rect 3622 6984 3858 7220
rect 3942 6984 4178 7220
rect 4262 6984 4498 7220
rect 4582 6984 4818 7220
rect 4902 6984 5138 7220
rect 5222 6984 5458 7220
rect 5542 6984 5778 7220
rect 5862 6984 6098 7220
rect 6182 6984 6418 7220
rect 6502 6984 6738 7220
rect 6822 6984 7058 7220
rect 7142 6984 7378 7220
rect 7462 6984 7698 7220
rect 7782 6984 8018 7220
rect 8102 6984 8338 7220
rect 8422 6984 8658 7220
rect 8742 6984 8978 7220
rect 9062 6984 9298 7220
rect 422 6380 658 6616
rect 742 6380 978 6616
rect 1062 6380 1298 6616
rect 1382 6380 1618 6616
rect 1702 6380 1938 6616
rect 2022 6380 2258 6616
rect 2342 6380 2578 6616
rect 2662 6380 2898 6616
rect 2982 6380 3218 6616
rect 3302 6380 3538 6616
rect 3622 6380 3858 6616
rect 3942 6380 4178 6616
rect 4262 6380 4498 6616
rect 4582 6380 4818 6616
rect 4902 6380 5138 6616
rect 5222 6380 5458 6616
rect 5542 6380 5778 6616
rect 5862 6380 6098 6616
rect 6182 6380 6418 6616
rect 6502 6380 6738 6616
rect 6822 6380 7058 6616
rect 7142 6380 7378 6616
rect 7462 6380 7698 6616
rect 7782 6380 8018 6616
rect 8102 6380 8338 6616
rect 8422 6380 8658 6616
rect 8742 6380 8978 6616
rect 9062 6380 9298 6616
rect 422 6014 658 6250
rect 742 6014 978 6250
rect 1062 6014 1298 6250
rect 1382 6014 1618 6250
rect 1702 6014 1938 6250
rect 2022 6014 2258 6250
rect 2342 6014 2578 6250
rect 2662 6014 2898 6250
rect 2982 6014 3218 6250
rect 3302 6014 3538 6250
rect 3622 6014 3858 6250
rect 3942 6014 4178 6250
rect 4262 6014 4498 6250
rect 4582 6014 4818 6250
rect 4902 6014 5138 6250
rect 5222 6014 5458 6250
rect 5542 6014 5778 6250
rect 5862 6014 6098 6250
rect 6182 6014 6418 6250
rect 6502 6014 6738 6250
rect 6822 6014 7058 6250
rect 7142 6014 7378 6250
rect 7462 6014 7698 6250
rect 7782 6014 8018 6250
rect 8102 6014 8338 6250
rect 8422 6014 8658 6250
rect 8742 6014 8978 6250
rect 9062 6014 9298 6250
rect 422 5410 658 5646
rect 742 5410 978 5646
rect 1062 5410 1298 5646
rect 1382 5410 1618 5646
rect 1702 5410 1938 5646
rect 2022 5410 2258 5646
rect 2342 5410 2578 5646
rect 2662 5410 2898 5646
rect 2982 5410 3218 5646
rect 3302 5410 3538 5646
rect 3622 5410 3858 5646
rect 3942 5410 4178 5646
rect 4262 5410 4498 5646
rect 4582 5410 4818 5646
rect 4902 5410 5138 5646
rect 5222 5410 5458 5646
rect 5542 5410 5778 5646
rect 5862 5410 6098 5646
rect 6182 5410 6418 5646
rect 6502 5410 6738 5646
rect 6822 5410 7058 5646
rect 7142 5410 7378 5646
rect 7462 5410 7698 5646
rect 7782 5410 8018 5646
rect 8102 5410 8338 5646
rect 8422 5410 8658 5646
rect 8742 5410 8978 5646
rect 9062 5410 9298 5646
rect 422 4804 658 5040
rect 742 4804 978 5040
rect 1062 4804 1298 5040
rect 1382 4804 1618 5040
rect 1702 4804 1938 5040
rect 2022 4804 2258 5040
rect 2342 4804 2578 5040
rect 2662 4804 2898 5040
rect 2982 4804 3218 5040
rect 3302 4804 3538 5040
rect 3622 4804 3858 5040
rect 3942 4804 4178 5040
rect 4262 4804 4498 5040
rect 4582 4804 4818 5040
rect 4902 4804 5138 5040
rect 5222 4804 5458 5040
rect 5542 4804 5778 5040
rect 5862 4804 6098 5040
rect 6182 4804 6418 5040
rect 6502 4804 6738 5040
rect 6822 4804 7058 5040
rect 7142 4804 7378 5040
rect 7462 4804 7698 5040
rect 7782 4804 8018 5040
rect 8102 4804 8338 5040
rect 8422 4804 8658 5040
rect 8742 4804 8978 5040
rect 9062 4804 9298 5040
rect 422 4200 658 4436
rect 742 4200 978 4436
rect 1062 4200 1298 4436
rect 1382 4200 1618 4436
rect 1702 4200 1938 4436
rect 2022 4200 2258 4436
rect 2342 4200 2578 4436
rect 2662 4200 2898 4436
rect 2982 4200 3218 4436
rect 3302 4200 3538 4436
rect 3622 4200 3858 4436
rect 3942 4200 4178 4436
rect 4262 4200 4498 4436
rect 4582 4200 4818 4436
rect 4902 4200 5138 4436
rect 5222 4200 5458 4436
rect 5542 4200 5778 4436
rect 5862 4200 6098 4436
rect 6182 4200 6418 4436
rect 6502 4200 6738 4436
rect 6822 4200 7058 4436
rect 7142 4200 7378 4436
rect 7462 4200 7698 4436
rect 7782 4200 8018 4436
rect 8102 4200 8338 4436
rect 8422 4200 8658 4436
rect 8742 4200 8978 4436
rect 9062 4200 9298 4436
rect 422 3594 658 3830
rect 742 3594 978 3830
rect 1062 3594 1298 3830
rect 1382 3594 1618 3830
rect 1702 3594 1938 3830
rect 2022 3594 2258 3830
rect 2342 3594 2578 3830
rect 2662 3594 2898 3830
rect 2982 3594 3218 3830
rect 3302 3594 3538 3830
rect 3622 3594 3858 3830
rect 3942 3594 4178 3830
rect 4262 3594 4498 3830
rect 4582 3594 4818 3830
rect 4902 3594 5138 3830
rect 5222 3594 5458 3830
rect 5542 3594 5778 3830
rect 5862 3594 6098 3830
rect 6182 3594 6418 3830
rect 6502 3594 6738 3830
rect 6822 3594 7058 3830
rect 7142 3594 7378 3830
rect 7462 3594 7698 3830
rect 7782 3594 8018 3830
rect 8102 3594 8338 3830
rect 8422 3594 8658 3830
rect 8742 3594 8978 3830
rect 9062 3594 9298 3830
rect 422 2990 658 3226
rect 742 2990 978 3226
rect 1062 2990 1298 3226
rect 1382 2990 1618 3226
rect 1702 2990 1938 3226
rect 2022 2990 2258 3226
rect 2342 2990 2578 3226
rect 2662 2990 2898 3226
rect 2982 2990 3218 3226
rect 3302 2990 3538 3226
rect 3622 2990 3858 3226
rect 3942 2990 4178 3226
rect 4262 2990 4498 3226
rect 4582 2990 4818 3226
rect 4902 2990 5138 3226
rect 5222 2990 5458 3226
rect 5542 2990 5778 3226
rect 5862 2990 6098 3226
rect 6182 2990 6418 3226
rect 6502 2990 6738 3226
rect 6822 2990 7058 3226
rect 7142 2990 7378 3226
rect 7462 2990 7698 3226
rect 7782 2990 8018 3226
rect 8102 2990 8338 3226
rect 8422 2990 8658 3226
rect 8742 2990 8978 3226
rect 9062 2990 9298 3226
rect 422 2624 658 2860
rect 742 2624 978 2860
rect 1062 2624 1298 2860
rect 1382 2624 1618 2860
rect 1702 2624 1938 2860
rect 2022 2624 2258 2860
rect 2342 2624 2578 2860
rect 2662 2624 2898 2860
rect 2982 2624 3218 2860
rect 3302 2624 3538 2860
rect 3622 2624 3858 2860
rect 3942 2624 4178 2860
rect 4262 2624 4498 2860
rect 4582 2624 4818 2860
rect 4902 2624 5138 2860
rect 5222 2624 5458 2860
rect 5542 2624 5778 2860
rect 5862 2624 6098 2860
rect 6182 2624 6418 2860
rect 6502 2624 6738 2860
rect 6822 2624 7058 2860
rect 7142 2624 7378 2860
rect 7462 2624 7698 2860
rect 7782 2624 8018 2860
rect 8102 2624 8338 2860
rect 8422 2624 8658 2860
rect 8742 2624 8978 2860
rect 9062 2624 9298 2860
rect 422 2020 658 2256
rect 742 2020 978 2256
rect 1062 2020 1298 2256
rect 1382 2020 1618 2256
rect 1702 2020 1938 2256
rect 2022 2020 2258 2256
rect 2342 2020 2578 2256
rect 2662 2020 2898 2256
rect 2982 2020 3218 2256
rect 3302 2020 3538 2256
rect 3622 2020 3858 2256
rect 3942 2020 4178 2256
rect 4262 2020 4498 2256
rect 4582 2020 4818 2256
rect 4902 2020 5138 2256
rect 5222 2020 5458 2256
rect 5542 2020 5778 2256
rect 5862 2020 6098 2256
rect 6182 2020 6418 2256
rect 6502 2020 6738 2256
rect 6822 2020 7058 2256
rect 7142 2020 7378 2256
rect 7462 2020 7698 2256
rect 7782 2020 8018 2256
rect 8102 2020 8338 2256
rect 8422 2020 8658 2256
rect 8742 2020 8978 2256
rect 9062 2020 9298 2256
rect 422 1414 658 1650
rect 742 1414 978 1650
rect 1062 1414 1298 1650
rect 1382 1414 1618 1650
rect 1702 1414 1938 1650
rect 2022 1414 2258 1650
rect 2342 1414 2578 1650
rect 2662 1414 2898 1650
rect 2982 1414 3218 1650
rect 3302 1414 3538 1650
rect 3622 1414 3858 1650
rect 3942 1414 4178 1650
rect 4262 1414 4498 1650
rect 4582 1414 4818 1650
rect 4902 1414 5138 1650
rect 5222 1414 5458 1650
rect 5542 1414 5778 1650
rect 5862 1414 6098 1650
rect 6182 1414 6418 1650
rect 6502 1414 6738 1650
rect 6822 1414 7058 1650
rect 7142 1414 7378 1650
rect 7462 1414 7698 1650
rect 7782 1414 8018 1650
rect 8102 1414 8338 1650
rect 8422 1414 8658 1650
rect 8742 1414 8978 1650
rect 9062 1414 9298 1650
rect 422 809 658 1045
rect 742 809 978 1045
rect 1062 809 1298 1045
rect 1382 809 1618 1045
rect 1702 809 1938 1045
rect 2022 809 2258 1045
rect 2342 809 2578 1045
rect 2662 809 2898 1045
rect 2982 809 3218 1045
rect 3302 809 3538 1045
rect 3622 809 3858 1045
rect 3942 809 4178 1045
rect 4262 809 4498 1045
rect 4582 809 4818 1045
rect 4902 809 5138 1045
rect 5222 809 5458 1045
rect 5542 809 5778 1045
rect 5862 809 6098 1045
rect 6182 809 6418 1045
rect 6502 809 6738 1045
rect 6822 809 7058 1045
rect 7142 809 7378 1045
rect 7462 809 7698 1045
rect 7782 809 8018 1045
rect 8102 809 8338 1045
rect 8422 809 8658 1045
rect 8742 809 8978 1045
rect 9062 809 9298 1045
rect 422 427 658 663
rect 742 427 978 663
rect 1062 427 1298 663
rect 1382 427 1618 663
rect 1702 427 1938 663
rect 2022 427 2258 663
rect 2342 427 2578 663
rect 2662 427 2898 663
rect 2982 427 3218 663
rect 3302 427 3538 663
rect 3622 427 3858 663
rect 3942 427 4178 663
rect 4262 427 4498 663
rect 4582 427 4818 663
rect 4902 427 5138 663
rect 5222 427 5458 663
rect 5542 427 5778 663
rect 5862 427 6098 663
rect 6182 427 6418 663
rect 6502 427 6738 663
rect 6822 427 7058 663
rect 7142 427 7378 663
rect 7462 427 7698 663
rect 7782 427 8018 663
rect 8102 427 8338 663
rect 8422 427 8658 663
rect 8742 427 8978 663
rect 9062 427 9298 663
rect 422 45 658 281
rect 742 45 978 281
rect 1062 45 1298 281
rect 1382 45 1618 281
rect 1702 45 1938 281
rect 2022 45 2258 281
rect 2342 45 2578 281
rect 2662 45 2898 281
rect 2982 45 3218 281
rect 3302 45 3538 281
rect 3622 45 3858 281
rect 3942 45 4178 281
rect 4262 45 4498 281
rect 4582 45 4818 281
rect 4902 45 5138 281
rect 5222 45 5458 281
rect 5542 45 5778 281
rect 5862 45 6098 281
rect 6182 45 6418 281
rect 6502 45 6738 281
rect 6822 45 7058 281
rect 7142 45 7378 281
rect 7462 45 7698 281
rect 7782 45 8018 281
rect 8102 45 8338 281
rect 8422 45 8658 281
rect 8742 45 8978 281
rect 9062 45 9298 281
<< metal5 >>
rect 0 39530 9600 39593
rect 0 34814 422 39530
rect 9298 34814 9600 39530
rect 0 34750 9600 34814
rect 0 18565 9600 18590
rect 0 18329 421 18565
rect 657 18329 741 18565
rect 977 18329 1061 18565
rect 1297 18329 1381 18565
rect 1617 18329 1701 18565
rect 1937 18329 2021 18565
rect 2257 18329 2341 18565
rect 2577 18329 2661 18565
rect 2897 18329 2981 18565
rect 3217 18329 3301 18565
rect 3537 18329 3621 18565
rect 3857 18329 3941 18565
rect 4177 18329 4261 18565
rect 4497 18329 4581 18565
rect 4817 18329 4901 18565
rect 5137 18329 5221 18565
rect 5457 18329 5541 18565
rect 5777 18329 5861 18565
rect 6097 18329 6181 18565
rect 6417 18329 6501 18565
rect 6737 18329 6821 18565
rect 7057 18329 7141 18565
rect 7377 18329 7461 18565
rect 7697 18329 7781 18565
rect 8017 18329 8101 18565
rect 8337 18329 8421 18565
rect 8657 18329 8741 18565
rect 8977 18329 9061 18565
rect 9297 18329 9600 18565
rect 0 18229 9600 18329
rect 0 17993 421 18229
rect 657 17993 741 18229
rect 977 17993 1061 18229
rect 1297 17993 1381 18229
rect 1617 17993 1701 18229
rect 1937 17993 2021 18229
rect 2257 17993 2341 18229
rect 2577 17993 2661 18229
rect 2897 17993 2981 18229
rect 3217 17993 3301 18229
rect 3537 17993 3621 18229
rect 3857 17993 3941 18229
rect 4177 17993 4261 18229
rect 4497 17993 4581 18229
rect 4817 17993 4901 18229
rect 5137 17993 5221 18229
rect 5457 17993 5541 18229
rect 5777 17993 5861 18229
rect 6097 17993 6181 18229
rect 6417 17993 6501 18229
rect 6737 17993 6821 18229
rect 7057 17993 7141 18229
rect 7377 17993 7461 18229
rect 7697 17993 7781 18229
rect 8017 17993 8101 18229
rect 8337 17993 8421 18229
rect 8657 17993 8741 18229
rect 8977 17993 9061 18229
rect 9297 17993 9600 18229
rect 0 17893 9600 17993
rect 0 17657 421 17893
rect 657 17657 741 17893
rect 977 17657 1061 17893
rect 1297 17657 1381 17893
rect 1617 17657 1701 17893
rect 1937 17657 2021 17893
rect 2257 17657 2341 17893
rect 2577 17657 2661 17893
rect 2897 17657 2981 17893
rect 3217 17657 3301 17893
rect 3537 17657 3621 17893
rect 3857 17657 3941 17893
rect 4177 17657 4261 17893
rect 4497 17657 4581 17893
rect 4817 17657 4901 17893
rect 5137 17657 5221 17893
rect 5457 17657 5541 17893
rect 5777 17657 5861 17893
rect 6097 17657 6181 17893
rect 6417 17657 6501 17893
rect 6737 17657 6821 17893
rect 7057 17657 7141 17893
rect 7377 17657 7461 17893
rect 7697 17657 7781 17893
rect 8017 17657 8101 17893
rect 8337 17657 8421 17893
rect 8657 17657 8741 17893
rect 8977 17657 9061 17893
rect 9297 17657 9600 17893
rect 0 17557 9600 17657
rect 0 17321 421 17557
rect 657 17321 741 17557
rect 977 17321 1061 17557
rect 1297 17321 1381 17557
rect 1617 17321 1701 17557
rect 1937 17321 2021 17557
rect 2257 17321 2341 17557
rect 2577 17321 2661 17557
rect 2897 17321 2981 17557
rect 3217 17321 3301 17557
rect 3537 17321 3621 17557
rect 3857 17321 3941 17557
rect 4177 17321 4261 17557
rect 4497 17321 4581 17557
rect 4817 17321 4901 17557
rect 5137 17321 5221 17557
rect 5457 17321 5541 17557
rect 5777 17321 5861 17557
rect 6097 17321 6181 17557
rect 6417 17321 6501 17557
rect 6737 17321 6821 17557
rect 7057 17321 7141 17557
rect 7377 17321 7461 17557
rect 7697 17321 7781 17557
rect 8017 17321 8101 17557
rect 8337 17321 8421 17557
rect 8657 17321 8741 17557
rect 8977 17321 9061 17557
rect 9297 17321 9600 17557
rect 0 17221 9600 17321
rect 0 16985 421 17221
rect 657 16985 741 17221
rect 977 16985 1061 17221
rect 1297 16985 1381 17221
rect 1617 16985 1701 17221
rect 1937 16985 2021 17221
rect 2257 16985 2341 17221
rect 2577 16985 2661 17221
rect 2897 16985 2981 17221
rect 3217 16985 3301 17221
rect 3537 16985 3621 17221
rect 3857 16985 3941 17221
rect 4177 16985 4261 17221
rect 4497 16985 4581 17221
rect 4817 16985 4901 17221
rect 5137 16985 5221 17221
rect 5457 16985 5541 17221
rect 5777 16985 5861 17221
rect 6097 16985 6181 17221
rect 6417 16985 6501 17221
rect 6737 16985 6821 17221
rect 7057 16985 7141 17221
rect 7377 16985 7461 17221
rect 7697 16985 7781 17221
rect 8017 16985 8101 17221
rect 8337 16985 8421 17221
rect 8657 16985 8741 17221
rect 8977 16985 9061 17221
rect 9297 16985 9600 17221
rect 0 16885 9600 16985
rect 0 16649 421 16885
rect 657 16649 741 16885
rect 977 16649 1061 16885
rect 1297 16649 1381 16885
rect 1617 16649 1701 16885
rect 1937 16649 2021 16885
rect 2257 16649 2341 16885
rect 2577 16649 2661 16885
rect 2897 16649 2981 16885
rect 3217 16649 3301 16885
rect 3537 16649 3621 16885
rect 3857 16649 3941 16885
rect 4177 16649 4261 16885
rect 4497 16649 4581 16885
rect 4817 16649 4901 16885
rect 5137 16649 5221 16885
rect 5457 16649 5541 16885
rect 5777 16649 5861 16885
rect 6097 16649 6181 16885
rect 6417 16649 6501 16885
rect 6737 16649 6821 16885
rect 7057 16649 7141 16885
rect 7377 16649 7461 16885
rect 7697 16649 7781 16885
rect 8017 16649 8101 16885
rect 8337 16649 8421 16885
rect 8657 16649 8741 16885
rect 8977 16649 9061 16885
rect 9297 16649 9600 16885
rect 0 16549 9600 16649
rect 0 16313 421 16549
rect 657 16313 741 16549
rect 977 16313 1061 16549
rect 1297 16313 1381 16549
rect 1617 16313 1701 16549
rect 1937 16313 2021 16549
rect 2257 16313 2341 16549
rect 2577 16313 2661 16549
rect 2897 16313 2981 16549
rect 3217 16313 3301 16549
rect 3537 16313 3621 16549
rect 3857 16313 3941 16549
rect 4177 16313 4261 16549
rect 4497 16313 4581 16549
rect 4817 16313 4901 16549
rect 5137 16313 5221 16549
rect 5457 16313 5541 16549
rect 5777 16313 5861 16549
rect 6097 16313 6181 16549
rect 6417 16313 6501 16549
rect 6737 16313 6821 16549
rect 7057 16313 7141 16549
rect 7377 16313 7461 16549
rect 7697 16313 7781 16549
rect 8017 16313 8101 16549
rect 8337 16313 8421 16549
rect 8657 16313 8741 16549
rect 8977 16313 9061 16549
rect 9297 16313 9600 16549
rect 0 16213 9600 16313
rect 0 15977 421 16213
rect 657 15977 741 16213
rect 977 15977 1061 16213
rect 1297 15977 1381 16213
rect 1617 15977 1701 16213
rect 1937 15977 2021 16213
rect 2257 15977 2341 16213
rect 2577 15977 2661 16213
rect 2897 15977 2981 16213
rect 3217 15977 3301 16213
rect 3537 15977 3621 16213
rect 3857 15977 3941 16213
rect 4177 15977 4261 16213
rect 4497 15977 4581 16213
rect 4817 15977 4901 16213
rect 5137 15977 5221 16213
rect 5457 15977 5541 16213
rect 5777 15977 5861 16213
rect 6097 15977 6181 16213
rect 6417 15977 6501 16213
rect 6737 15977 6821 16213
rect 7057 15977 7141 16213
rect 7377 15977 7461 16213
rect 7697 15977 7781 16213
rect 8017 15977 8101 16213
rect 8337 15977 8421 16213
rect 8657 15977 8741 16213
rect 8977 15977 9061 16213
rect 9297 15977 9600 16213
rect 0 15877 9600 15977
rect 0 15641 421 15877
rect 657 15641 741 15877
rect 977 15641 1061 15877
rect 1297 15641 1381 15877
rect 1617 15641 1701 15877
rect 1937 15641 2021 15877
rect 2257 15641 2341 15877
rect 2577 15641 2661 15877
rect 2897 15641 2981 15877
rect 3217 15641 3301 15877
rect 3537 15641 3621 15877
rect 3857 15641 3941 15877
rect 4177 15641 4261 15877
rect 4497 15641 4581 15877
rect 4817 15641 4901 15877
rect 5137 15641 5221 15877
rect 5457 15641 5541 15877
rect 5777 15641 5861 15877
rect 6097 15641 6181 15877
rect 6417 15641 6501 15877
rect 6737 15641 6821 15877
rect 7057 15641 7141 15877
rect 7377 15641 7461 15877
rect 7697 15641 7781 15877
rect 8017 15641 8101 15877
rect 8337 15641 8421 15877
rect 8657 15641 8741 15877
rect 8977 15641 9061 15877
rect 9297 15641 9600 15877
rect 0 15541 9600 15641
rect 0 15305 421 15541
rect 657 15305 741 15541
rect 977 15305 1061 15541
rect 1297 15305 1381 15541
rect 1617 15305 1701 15541
rect 1937 15305 2021 15541
rect 2257 15305 2341 15541
rect 2577 15305 2661 15541
rect 2897 15305 2981 15541
rect 3217 15305 3301 15541
rect 3537 15305 3621 15541
rect 3857 15305 3941 15541
rect 4177 15305 4261 15541
rect 4497 15305 4581 15541
rect 4817 15305 4901 15541
rect 5137 15305 5221 15541
rect 5457 15305 5541 15541
rect 5777 15305 5861 15541
rect 6097 15305 6181 15541
rect 6417 15305 6501 15541
rect 6737 15305 6821 15541
rect 7057 15305 7141 15541
rect 7377 15305 7461 15541
rect 7697 15305 7781 15541
rect 8017 15305 8101 15541
rect 8337 15305 8421 15541
rect 8657 15305 8741 15541
rect 8977 15305 9061 15541
rect 9297 15305 9600 15541
rect 0 15205 9600 15305
rect 0 14969 421 15205
rect 657 14969 741 15205
rect 977 14969 1061 15205
rect 1297 14969 1381 15205
rect 1617 14969 1701 15205
rect 1937 14969 2021 15205
rect 2257 14969 2341 15205
rect 2577 14969 2661 15205
rect 2897 14969 2981 15205
rect 3217 14969 3301 15205
rect 3537 14969 3621 15205
rect 3857 14969 3941 15205
rect 4177 14969 4261 15205
rect 4497 14969 4581 15205
rect 4817 14969 4901 15205
rect 5137 14969 5221 15205
rect 5457 14969 5541 15205
rect 5777 14969 5861 15205
rect 6097 14969 6181 15205
rect 6417 14969 6501 15205
rect 6737 14969 6821 15205
rect 7057 14969 7141 15205
rect 7377 14969 7461 15205
rect 7697 14969 7781 15205
rect 8017 14969 8101 15205
rect 8337 14969 8421 15205
rect 8657 14969 8741 15205
rect 8977 14969 9061 15205
rect 9297 14969 9600 15205
rect 0 14869 9600 14969
rect 0 14633 421 14869
rect 657 14633 741 14869
rect 977 14633 1061 14869
rect 1297 14633 1381 14869
rect 1617 14633 1701 14869
rect 1937 14633 2021 14869
rect 2257 14633 2341 14869
rect 2577 14633 2661 14869
rect 2897 14633 2981 14869
rect 3217 14633 3301 14869
rect 3537 14633 3621 14869
rect 3857 14633 3941 14869
rect 4177 14633 4261 14869
rect 4497 14633 4581 14869
rect 4817 14633 4901 14869
rect 5137 14633 5221 14869
rect 5457 14633 5541 14869
rect 5777 14633 5861 14869
rect 6097 14633 6181 14869
rect 6417 14633 6501 14869
rect 6737 14633 6821 14869
rect 7057 14633 7141 14869
rect 7377 14633 7461 14869
rect 7697 14633 7781 14869
rect 8017 14633 8101 14869
rect 8337 14633 8421 14869
rect 8657 14633 8741 14869
rect 8977 14633 9061 14869
rect 9297 14633 9600 14869
rect 0 14533 9600 14633
rect 0 14297 421 14533
rect 657 14297 741 14533
rect 977 14297 1061 14533
rect 1297 14297 1381 14533
rect 1617 14297 1701 14533
rect 1937 14297 2021 14533
rect 2257 14297 2341 14533
rect 2577 14297 2661 14533
rect 2897 14297 2981 14533
rect 3217 14297 3301 14533
rect 3537 14297 3621 14533
rect 3857 14297 3941 14533
rect 4177 14297 4261 14533
rect 4497 14297 4581 14533
rect 4817 14297 4901 14533
rect 5137 14297 5221 14533
rect 5457 14297 5541 14533
rect 5777 14297 5861 14533
rect 6097 14297 6181 14533
rect 6417 14297 6501 14533
rect 6737 14297 6821 14533
rect 7057 14297 7141 14533
rect 7377 14297 7461 14533
rect 7697 14297 7781 14533
rect 8017 14297 8101 14533
rect 8337 14297 8421 14533
rect 8657 14297 8741 14533
rect 8977 14297 9061 14533
rect 9297 14297 9600 14533
rect 0 14197 9600 14297
rect 0 13961 421 14197
rect 657 13961 741 14197
rect 977 13961 1061 14197
rect 1297 13961 1381 14197
rect 1617 13961 1701 14197
rect 1937 13961 2021 14197
rect 2257 13961 2341 14197
rect 2577 13961 2661 14197
rect 2897 13961 2981 14197
rect 3217 13961 3301 14197
rect 3537 13961 3621 14197
rect 3857 13961 3941 14197
rect 4177 13961 4261 14197
rect 4497 13961 4581 14197
rect 4817 13961 4901 14197
rect 5137 13961 5221 14197
rect 5457 13961 5541 14197
rect 5777 13961 5861 14197
rect 6097 13961 6181 14197
rect 6417 13961 6501 14197
rect 6737 13961 6821 14197
rect 7057 13961 7141 14197
rect 7377 13961 7461 14197
rect 7697 13961 7781 14197
rect 8017 13961 8101 14197
rect 8337 13961 8421 14197
rect 8657 13961 8741 14197
rect 8977 13961 9061 14197
rect 9297 13961 9600 14197
rect 0 13861 9600 13961
rect 0 13625 421 13861
rect 657 13625 741 13861
rect 977 13625 1061 13861
rect 1297 13625 1381 13861
rect 1617 13625 1701 13861
rect 1937 13625 2021 13861
rect 2257 13625 2341 13861
rect 2577 13625 2661 13861
rect 2897 13625 2981 13861
rect 3217 13625 3301 13861
rect 3537 13625 3621 13861
rect 3857 13625 3941 13861
rect 4177 13625 4261 13861
rect 4497 13625 4581 13861
rect 4817 13625 4901 13861
rect 5137 13625 5221 13861
rect 5457 13625 5541 13861
rect 5777 13625 5861 13861
rect 6097 13625 6181 13861
rect 6417 13625 6501 13861
rect 6737 13625 6821 13861
rect 7057 13625 7141 13861
rect 7377 13625 7461 13861
rect 7697 13625 7781 13861
rect 8017 13625 8101 13861
rect 8337 13625 8421 13861
rect 8657 13625 8741 13861
rect 8977 13625 9061 13861
rect 9297 13625 9600 13861
rect 0 13600 9600 13625
rect 0 13256 9600 13280
rect 0 13020 422 13256
rect 658 13020 742 13256
rect 978 13020 1062 13256
rect 1298 13020 1382 13256
rect 1618 13020 1702 13256
rect 1938 13020 2022 13256
rect 2258 13020 2342 13256
rect 2578 13020 2662 13256
rect 2898 13020 2982 13256
rect 3218 13020 3302 13256
rect 3538 13020 3622 13256
rect 3858 13020 3942 13256
rect 4178 13020 4262 13256
rect 4498 13020 4582 13256
rect 4818 13020 4902 13256
rect 5138 13020 5222 13256
rect 5458 13020 5542 13256
rect 5778 13020 5862 13256
rect 6098 13020 6182 13256
rect 6418 13020 6502 13256
rect 6738 13020 6822 13256
rect 7058 13020 7142 13256
rect 7378 13020 7462 13256
rect 7698 13020 7782 13256
rect 8018 13020 8102 13256
rect 8338 13020 8422 13256
rect 8658 13020 8742 13256
rect 8978 13020 9062 13256
rect 9298 13020 9600 13256
rect 0 12690 9600 13020
rect 0 12454 422 12690
rect 658 12454 742 12690
rect 978 12454 1062 12690
rect 1298 12454 1382 12690
rect 1618 12454 1702 12690
rect 1938 12454 2022 12690
rect 2258 12454 2342 12690
rect 2578 12454 2662 12690
rect 2898 12454 2982 12690
rect 3218 12454 3302 12690
rect 3538 12454 3622 12690
rect 3858 12454 3942 12690
rect 4178 12454 4262 12690
rect 4498 12454 4582 12690
rect 4818 12454 4902 12690
rect 5138 12454 5222 12690
rect 5458 12454 5542 12690
rect 5778 12454 5862 12690
rect 6098 12454 6182 12690
rect 6418 12454 6502 12690
rect 6738 12454 6822 12690
rect 7058 12454 7142 12690
rect 7378 12454 7462 12690
rect 7698 12454 7782 12690
rect 8018 12454 8102 12690
rect 8338 12454 8422 12690
rect 8658 12454 8742 12690
rect 8978 12454 9062 12690
rect 9298 12454 9600 12690
rect 0 12430 9600 12454
rect 0 12086 9600 12110
rect 0 11850 422 12086
rect 658 11850 742 12086
rect 978 11850 1062 12086
rect 1298 11850 1382 12086
rect 1618 11850 1702 12086
rect 1938 11850 2022 12086
rect 2258 11850 2342 12086
rect 2578 11850 2662 12086
rect 2898 11850 2982 12086
rect 3218 11850 3302 12086
rect 3538 11850 3622 12086
rect 3858 11850 3942 12086
rect 4178 11850 4262 12086
rect 4498 11850 4582 12086
rect 4818 11850 4902 12086
rect 5138 11850 5222 12086
rect 5458 11850 5542 12086
rect 5778 11850 5862 12086
rect 6098 11850 6182 12086
rect 6418 11850 6502 12086
rect 6738 11850 6822 12086
rect 7058 11850 7142 12086
rect 7378 11850 7462 12086
rect 7698 11850 7782 12086
rect 8018 11850 8102 12086
rect 8338 11850 8422 12086
rect 8658 11850 8742 12086
rect 8978 11850 9062 12086
rect 9298 11850 9600 12086
rect 0 11520 9600 11850
rect 0 11284 422 11520
rect 658 11284 742 11520
rect 978 11284 1062 11520
rect 1298 11284 1382 11520
rect 1618 11284 1702 11520
rect 1938 11284 2022 11520
rect 2258 11284 2342 11520
rect 2578 11284 2662 11520
rect 2898 11284 2982 11520
rect 3218 11284 3302 11520
rect 3538 11284 3622 11520
rect 3858 11284 3942 11520
rect 4178 11284 4262 11520
rect 4498 11284 4582 11520
rect 4818 11284 4902 11520
rect 5138 11284 5222 11520
rect 5458 11284 5542 11520
rect 5778 11284 5862 11520
rect 6098 11284 6182 11520
rect 6418 11284 6502 11520
rect 6738 11284 6822 11520
rect 7058 11284 7142 11520
rect 7378 11284 7462 11520
rect 7698 11284 7782 11520
rect 8018 11284 8102 11520
rect 8338 11284 8422 11520
rect 8658 11284 8742 11520
rect 8978 11284 9062 11520
rect 9298 11284 9600 11520
rect 0 11260 9600 11284
rect 0 10158 9600 10940
rect 0 9922 422 10158
rect 658 9922 742 10158
rect 978 9922 1062 10158
rect 1298 9922 1382 10158
rect 1618 9922 1702 10158
rect 1938 9922 2022 10158
rect 2258 9922 2342 10158
rect 2578 9922 2662 10158
rect 2898 9922 2982 10158
rect 3218 9922 3302 10158
rect 3538 9922 3622 10158
rect 3858 9922 3942 10158
rect 4178 9922 4262 10158
rect 4498 9922 4582 10158
rect 4818 9922 4902 10158
rect 5138 9922 5222 10158
rect 5458 9922 5542 10158
rect 5778 9922 5862 10158
rect 6098 9922 6182 10158
rect 6418 9922 6502 10158
rect 6738 9922 6822 10158
rect 7058 9922 7142 10158
rect 7378 9922 7462 10158
rect 7698 9922 7782 10158
rect 8018 9922 8102 10158
rect 8338 9922 8422 10158
rect 8658 9922 8742 10158
rect 8978 9922 9062 10158
rect 9298 9922 9600 10158
rect 0 9140 9600 9922
rect 0 8796 9600 8820
rect 0 8560 422 8796
rect 658 8560 742 8796
rect 978 8560 1062 8796
rect 1298 8560 1382 8796
rect 1618 8560 1702 8796
rect 1938 8560 2022 8796
rect 2258 8560 2342 8796
rect 2578 8560 2662 8796
rect 2898 8560 2982 8796
rect 3218 8560 3302 8796
rect 3538 8560 3622 8796
rect 3858 8560 3942 8796
rect 4178 8560 4262 8796
rect 4498 8560 4582 8796
rect 4818 8560 4902 8796
rect 5138 8560 5222 8796
rect 5458 8560 5542 8796
rect 5778 8560 5862 8796
rect 6098 8560 6182 8796
rect 6418 8560 6502 8796
rect 6738 8560 6822 8796
rect 7058 8560 7142 8796
rect 7378 8560 7462 8796
rect 7698 8560 7782 8796
rect 8018 8560 8102 8796
rect 8338 8560 8422 8796
rect 8658 8560 8742 8796
rect 8978 8560 9062 8796
rect 9298 8560 9600 8796
rect 0 8190 9600 8560
rect 0 7954 422 8190
rect 658 7954 742 8190
rect 978 7954 1062 8190
rect 1298 7954 1382 8190
rect 1618 7954 1702 8190
rect 1938 7954 2022 8190
rect 2258 7954 2342 8190
rect 2578 7954 2662 8190
rect 2898 7954 2982 8190
rect 3218 7954 3302 8190
rect 3538 7954 3622 8190
rect 3858 7954 3942 8190
rect 4178 7954 4262 8190
rect 4498 7954 4582 8190
rect 4818 7954 4902 8190
rect 5138 7954 5222 8190
rect 5458 7954 5542 8190
rect 5778 7954 5862 8190
rect 6098 7954 6182 8190
rect 6418 7954 6502 8190
rect 6738 7954 6822 8190
rect 7058 7954 7142 8190
rect 7378 7954 7462 8190
rect 7698 7954 7782 8190
rect 8018 7954 8102 8190
rect 8338 7954 8422 8190
rect 8658 7954 8742 8190
rect 8978 7954 9062 8190
rect 9298 7954 9600 8190
rect 0 7930 9600 7954
rect 0 7586 9600 7610
rect 0 7350 422 7586
rect 658 7350 742 7586
rect 978 7350 1062 7586
rect 1298 7350 1382 7586
rect 1618 7350 1702 7586
rect 1938 7350 2022 7586
rect 2258 7350 2342 7586
rect 2578 7350 2662 7586
rect 2898 7350 2982 7586
rect 3218 7350 3302 7586
rect 3538 7350 3622 7586
rect 3858 7350 3942 7586
rect 4178 7350 4262 7586
rect 4498 7350 4582 7586
rect 4818 7350 4902 7586
rect 5138 7350 5222 7586
rect 5458 7350 5542 7586
rect 5778 7350 5862 7586
rect 6098 7350 6182 7586
rect 6418 7350 6502 7586
rect 6738 7350 6822 7586
rect 7058 7350 7142 7586
rect 7378 7350 7462 7586
rect 7698 7350 7782 7586
rect 8018 7350 8102 7586
rect 8338 7350 8422 7586
rect 8658 7350 8742 7586
rect 8978 7350 9062 7586
rect 9298 7350 9600 7586
rect 0 7220 9600 7350
rect 0 6984 422 7220
rect 658 6984 742 7220
rect 978 6984 1062 7220
rect 1298 6984 1382 7220
rect 1618 6984 1702 7220
rect 1938 6984 2022 7220
rect 2258 6984 2342 7220
rect 2578 6984 2662 7220
rect 2898 6984 2982 7220
rect 3218 6984 3302 7220
rect 3538 6984 3622 7220
rect 3858 6984 3942 7220
rect 4178 6984 4262 7220
rect 4498 6984 4582 7220
rect 4818 6984 4902 7220
rect 5138 6984 5222 7220
rect 5458 6984 5542 7220
rect 5778 6984 5862 7220
rect 6098 6984 6182 7220
rect 6418 6984 6502 7220
rect 6738 6984 6822 7220
rect 7058 6984 7142 7220
rect 7378 6984 7462 7220
rect 7698 6984 7782 7220
rect 8018 6984 8102 7220
rect 8338 6984 8422 7220
rect 8658 6984 8742 7220
rect 8978 6984 9062 7220
rect 9298 6984 9600 7220
rect 0 6960 9600 6984
rect 0 6616 9600 6640
rect 0 6380 422 6616
rect 658 6380 742 6616
rect 978 6380 1062 6616
rect 1298 6380 1382 6616
rect 1618 6380 1702 6616
rect 1938 6380 2022 6616
rect 2258 6380 2342 6616
rect 2578 6380 2662 6616
rect 2898 6380 2982 6616
rect 3218 6380 3302 6616
rect 3538 6380 3622 6616
rect 3858 6380 3942 6616
rect 4178 6380 4262 6616
rect 4498 6380 4582 6616
rect 4818 6380 4902 6616
rect 5138 6380 5222 6616
rect 5458 6380 5542 6616
rect 5778 6380 5862 6616
rect 6098 6380 6182 6616
rect 6418 6380 6502 6616
rect 6738 6380 6822 6616
rect 7058 6380 7142 6616
rect 7378 6380 7462 6616
rect 7698 6380 7782 6616
rect 8018 6380 8102 6616
rect 8338 6380 8422 6616
rect 8658 6380 8742 6616
rect 8978 6380 9062 6616
rect 9298 6380 9600 6616
rect 0 6250 9600 6380
rect 0 6014 422 6250
rect 658 6014 742 6250
rect 978 6014 1062 6250
rect 1298 6014 1382 6250
rect 1618 6014 1702 6250
rect 1938 6014 2022 6250
rect 2258 6014 2342 6250
rect 2578 6014 2662 6250
rect 2898 6014 2982 6250
rect 3218 6014 3302 6250
rect 3538 6014 3622 6250
rect 3858 6014 3942 6250
rect 4178 6014 4262 6250
rect 4498 6014 4582 6250
rect 4818 6014 4902 6250
rect 5138 6014 5222 6250
rect 5458 6014 5542 6250
rect 5778 6014 5862 6250
rect 6098 6014 6182 6250
rect 6418 6014 6502 6250
rect 6738 6014 6822 6250
rect 7058 6014 7142 6250
rect 7378 6014 7462 6250
rect 7698 6014 7782 6250
rect 8018 6014 8102 6250
rect 8338 6014 8422 6250
rect 8658 6014 8742 6250
rect 8978 6014 9062 6250
rect 9298 6014 9600 6250
rect 0 5990 9600 6014
rect 0 5646 9600 5670
rect 0 5410 422 5646
rect 658 5410 742 5646
rect 978 5410 1062 5646
rect 1298 5410 1382 5646
rect 1618 5410 1702 5646
rect 1938 5410 2022 5646
rect 2258 5410 2342 5646
rect 2578 5410 2662 5646
rect 2898 5410 2982 5646
rect 3218 5410 3302 5646
rect 3538 5410 3622 5646
rect 3858 5410 3942 5646
rect 4178 5410 4262 5646
rect 4498 5410 4582 5646
rect 4818 5410 4902 5646
rect 5138 5410 5222 5646
rect 5458 5410 5542 5646
rect 5778 5410 5862 5646
rect 6098 5410 6182 5646
rect 6418 5410 6502 5646
rect 6738 5410 6822 5646
rect 7058 5410 7142 5646
rect 7378 5410 7462 5646
rect 7698 5410 7782 5646
rect 8018 5410 8102 5646
rect 8338 5410 8422 5646
rect 8658 5410 8742 5646
rect 8978 5410 9062 5646
rect 9298 5410 9600 5646
rect 0 5040 9600 5410
rect 0 4804 422 5040
rect 658 4804 742 5040
rect 978 4804 1062 5040
rect 1298 4804 1382 5040
rect 1618 4804 1702 5040
rect 1938 4804 2022 5040
rect 2258 4804 2342 5040
rect 2578 4804 2662 5040
rect 2898 4804 2982 5040
rect 3218 4804 3302 5040
rect 3538 4804 3622 5040
rect 3858 4804 3942 5040
rect 4178 4804 4262 5040
rect 4498 4804 4582 5040
rect 4818 4804 4902 5040
rect 5138 4804 5222 5040
rect 5458 4804 5542 5040
rect 5778 4804 5862 5040
rect 6098 4804 6182 5040
rect 6418 4804 6502 5040
rect 6738 4804 6822 5040
rect 7058 4804 7142 5040
rect 7378 4804 7462 5040
rect 7698 4804 7782 5040
rect 8018 4804 8102 5040
rect 8338 4804 8422 5040
rect 8658 4804 8742 5040
rect 8978 4804 9062 5040
rect 9298 4804 9600 5040
rect 0 4780 9600 4804
rect 0 4436 9600 4460
rect 0 4200 422 4436
rect 658 4200 742 4436
rect 978 4200 1062 4436
rect 1298 4200 1382 4436
rect 1618 4200 1702 4436
rect 1938 4200 2022 4436
rect 2258 4200 2342 4436
rect 2578 4200 2662 4436
rect 2898 4200 2982 4436
rect 3218 4200 3302 4436
rect 3538 4200 3622 4436
rect 3858 4200 3942 4436
rect 4178 4200 4262 4436
rect 4498 4200 4582 4436
rect 4818 4200 4902 4436
rect 5138 4200 5222 4436
rect 5458 4200 5542 4436
rect 5778 4200 5862 4436
rect 6098 4200 6182 4436
rect 6418 4200 6502 4436
rect 6738 4200 6822 4436
rect 7058 4200 7142 4436
rect 7378 4200 7462 4436
rect 7698 4200 7782 4436
rect 8018 4200 8102 4436
rect 8338 4200 8422 4436
rect 8658 4200 8742 4436
rect 8978 4200 9062 4436
rect 9298 4200 9600 4436
rect 0 3830 9600 4200
rect 0 3594 422 3830
rect 658 3594 742 3830
rect 978 3594 1062 3830
rect 1298 3594 1382 3830
rect 1618 3594 1702 3830
rect 1938 3594 2022 3830
rect 2258 3594 2342 3830
rect 2578 3594 2662 3830
rect 2898 3594 2982 3830
rect 3218 3594 3302 3830
rect 3538 3594 3622 3830
rect 3858 3594 3942 3830
rect 4178 3594 4262 3830
rect 4498 3594 4582 3830
rect 4818 3594 4902 3830
rect 5138 3594 5222 3830
rect 5458 3594 5542 3830
rect 5778 3594 5862 3830
rect 6098 3594 6182 3830
rect 6418 3594 6502 3830
rect 6738 3594 6822 3830
rect 7058 3594 7142 3830
rect 7378 3594 7462 3830
rect 7698 3594 7782 3830
rect 8018 3594 8102 3830
rect 8338 3594 8422 3830
rect 8658 3594 8742 3830
rect 8978 3594 9062 3830
rect 9298 3594 9600 3830
rect 0 3570 9600 3594
rect 0 3226 9600 3250
rect 0 2990 422 3226
rect 658 2990 742 3226
rect 978 2990 1062 3226
rect 1298 2990 1382 3226
rect 1618 2990 1702 3226
rect 1938 2990 2022 3226
rect 2258 2990 2342 3226
rect 2578 2990 2662 3226
rect 2898 2990 2982 3226
rect 3218 2990 3302 3226
rect 3538 2990 3622 3226
rect 3858 2990 3942 3226
rect 4178 2990 4262 3226
rect 4498 2990 4582 3226
rect 4818 2990 4902 3226
rect 5138 2990 5222 3226
rect 5458 2990 5542 3226
rect 5778 2990 5862 3226
rect 6098 2990 6182 3226
rect 6418 2990 6502 3226
rect 6738 2990 6822 3226
rect 7058 2990 7142 3226
rect 7378 2990 7462 3226
rect 7698 2990 7782 3226
rect 8018 2990 8102 3226
rect 8338 2990 8422 3226
rect 8658 2990 8742 3226
rect 8978 2990 9062 3226
rect 9298 2990 9600 3226
rect 0 2860 9600 2990
rect 0 2624 422 2860
rect 658 2624 742 2860
rect 978 2624 1062 2860
rect 1298 2624 1382 2860
rect 1618 2624 1702 2860
rect 1938 2624 2022 2860
rect 2258 2624 2342 2860
rect 2578 2624 2662 2860
rect 2898 2624 2982 2860
rect 3218 2624 3302 2860
rect 3538 2624 3622 2860
rect 3858 2624 3942 2860
rect 4178 2624 4262 2860
rect 4498 2624 4582 2860
rect 4818 2624 4902 2860
rect 5138 2624 5222 2860
rect 5458 2624 5542 2860
rect 5778 2624 5862 2860
rect 6098 2624 6182 2860
rect 6418 2624 6502 2860
rect 6738 2624 6822 2860
rect 7058 2624 7142 2860
rect 7378 2624 7462 2860
rect 7698 2624 7782 2860
rect 8018 2624 8102 2860
rect 8338 2624 8422 2860
rect 8658 2624 8742 2860
rect 8978 2624 9062 2860
rect 9298 2624 9600 2860
rect 0 2600 9600 2624
rect 0 2256 9600 2280
rect 0 2020 422 2256
rect 658 2020 742 2256
rect 978 2020 1062 2256
rect 1298 2020 1382 2256
rect 1618 2020 1702 2256
rect 1938 2020 2022 2256
rect 2258 2020 2342 2256
rect 2578 2020 2662 2256
rect 2898 2020 2982 2256
rect 3218 2020 3302 2256
rect 3538 2020 3622 2256
rect 3858 2020 3942 2256
rect 4178 2020 4262 2256
rect 4498 2020 4582 2256
rect 4818 2020 4902 2256
rect 5138 2020 5222 2256
rect 5458 2020 5542 2256
rect 5778 2020 5862 2256
rect 6098 2020 6182 2256
rect 6418 2020 6502 2256
rect 6738 2020 6822 2256
rect 7058 2020 7142 2256
rect 7378 2020 7462 2256
rect 7698 2020 7782 2256
rect 8018 2020 8102 2256
rect 8338 2020 8422 2256
rect 8658 2020 8742 2256
rect 8978 2020 9062 2256
rect 9298 2020 9600 2256
rect 0 1650 9600 2020
rect 0 1414 422 1650
rect 658 1414 742 1650
rect 978 1414 1062 1650
rect 1298 1414 1382 1650
rect 1618 1414 1702 1650
rect 1938 1414 2022 1650
rect 2258 1414 2342 1650
rect 2578 1414 2662 1650
rect 2898 1414 2982 1650
rect 3218 1414 3302 1650
rect 3538 1414 3622 1650
rect 3858 1414 3942 1650
rect 4178 1414 4262 1650
rect 4498 1414 4582 1650
rect 4818 1414 4902 1650
rect 5138 1414 5222 1650
rect 5458 1414 5542 1650
rect 5778 1414 5862 1650
rect 6098 1414 6182 1650
rect 6418 1414 6502 1650
rect 6738 1414 6822 1650
rect 7058 1414 7142 1650
rect 7378 1414 7462 1650
rect 7698 1414 7782 1650
rect 8018 1414 8102 1650
rect 8338 1414 8422 1650
rect 8658 1414 8742 1650
rect 8978 1414 9062 1650
rect 9298 1414 9600 1650
rect 0 1390 9600 1414
rect 0 1045 9600 1070
rect 0 809 422 1045
rect 658 809 742 1045
rect 978 809 1062 1045
rect 1298 809 1382 1045
rect 1618 809 1702 1045
rect 1938 809 2022 1045
rect 2258 809 2342 1045
rect 2578 809 2662 1045
rect 2898 809 2982 1045
rect 3218 809 3302 1045
rect 3538 809 3622 1045
rect 3858 809 3942 1045
rect 4178 809 4262 1045
rect 4498 809 4582 1045
rect 4818 809 4902 1045
rect 5138 809 5222 1045
rect 5458 809 5542 1045
rect 5778 809 5862 1045
rect 6098 809 6182 1045
rect 6418 809 6502 1045
rect 6738 809 6822 1045
rect 7058 809 7142 1045
rect 7378 809 7462 1045
rect 7698 809 7782 1045
rect 8018 809 8102 1045
rect 8338 809 8422 1045
rect 8658 809 8742 1045
rect 8978 809 9062 1045
rect 9298 809 9600 1045
rect 0 663 9600 809
rect 0 427 422 663
rect 658 427 742 663
rect 978 427 1062 663
rect 1298 427 1382 663
rect 1618 427 1702 663
rect 1938 427 2022 663
rect 2258 427 2342 663
rect 2578 427 2662 663
rect 2898 427 2982 663
rect 3218 427 3302 663
rect 3538 427 3622 663
rect 3858 427 3942 663
rect 4178 427 4262 663
rect 4498 427 4582 663
rect 4818 427 4902 663
rect 5138 427 5222 663
rect 5458 427 5542 663
rect 5778 427 5862 663
rect 6098 427 6182 663
rect 6418 427 6502 663
rect 6738 427 6822 663
rect 7058 427 7142 663
rect 7378 427 7462 663
rect 7698 427 7782 663
rect 8018 427 8102 663
rect 8338 427 8422 663
rect 8658 427 8742 663
rect 8978 427 9062 663
rect 9298 427 9600 663
rect 0 281 9600 427
rect 0 45 422 281
rect 658 45 742 281
rect 978 45 1062 281
rect 1298 45 1382 281
rect 1618 45 1702 281
rect 1938 45 2022 281
rect 2258 45 2342 281
rect 2578 45 2662 281
rect 2898 45 2982 281
rect 3218 45 3302 281
rect 3538 45 3622 281
rect 3858 45 3942 281
rect 4178 45 4262 281
rect 4498 45 4582 281
rect 4818 45 4902 281
rect 5138 45 5222 281
rect 5458 45 5542 281
rect 5778 45 5862 281
rect 6098 45 6182 281
rect 6418 45 6502 281
rect 6738 45 6822 281
rect 7058 45 7142 281
rect 7378 45 7462 281
rect 7698 45 7782 281
rect 8018 45 8102 281
rect 8338 45 8422 281
rect 8658 45 8742 281
rect 8978 45 9062 281
rect 9298 45 9600 281
rect 0 20 9600 45
<< labels >>
flabel metal4 s 9346 13600 9600 18593 3 FreeSans 520 180 0 0 vddio
port 1 nsew
flabel metal4 s 9346 34750 9600 39593 3 FreeSans 520 180 0 0 vssio
port 2 nsew
flabel metal4 s 9346 1370 9600 2300 3 FreeSans 520 180 0 0 vccd
port 3 nsew
flabel metal4 s 9346 12410 9600 13300 3 FreeSans 520 180 0 0 vddio_q
port 4 nsew
flabel metal4 s 9346 6940 9600 7630 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 9346 9140 9600 9206 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 9346 3550 9600 4480 3 FreeSans 520 180 0 0 vddio
port 1 nsew
flabel metal4 s 9346 0 9600 1090 3 FreeSans 520 180 0 0 vcchib
port 6 nsew
flabel metal4 s 9346 10874 9600 10940 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 9346 9922 9600 10158 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 9346 5970 9600 6660 3 FreeSans 520 180 0 0 vswitch
port 7 nsew
flabel metal4 s 9346 4760 9600 5690 3 FreeSans 520 180 0 0 vssio
port 2 nsew
flabel metal4 s 9346 11240 9600 12130 3 FreeSans 520 180 0 0 vssio_q
port 8 nsew
flabel metal4 s 9407 2580 9600 3270 3 FreeSans 520 180 0 0 vdda
port 9 nsew
flabel metal4 s 9346 7910 9600 8840 3 FreeSans 520 180 0 0 vssd
port 10 nsew
flabel metal4 s 0 13600 254 18593 3 FreeSans 520 0 0 0 vddio
port 1 nsew
flabel metal4 s 0 34750 254 39593 3 FreeSans 520 0 0 0 vssio
port 2 nsew
flabel metal4 s 0 1370 254 2300 3 FreeSans 520 0 0 0 vccd
port 3 nsew
flabel metal4 s 0 12410 254 13300 3 FreeSans 520 0 0 0 vddio_q
port 4 nsew
flabel metal4 s 0 6940 254 7630 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 9140 254 9206 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 3550 254 4480 3 FreeSans 520 0 0 0 vddio
port 1 nsew
flabel metal4 s 0 0 254 1090 3 FreeSans 520 0 0 0 vcchib
port 6 nsew
flabel metal4 s 0 10874 254 10940 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 9922 254 10158 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 5970 254 6660 3 FreeSans 520 0 0 0 vswitch
port 7 nsew
flabel metal4 s 0 4760 254 5690 3 FreeSans 520 0 0 0 vssio
port 2 nsew
flabel metal4 s 0 11240 254 12130 3 FreeSans 520 0 0 0 vssio_q
port 8 nsew
flabel metal4 s 0 2580 193 3270 3 FreeSans 520 0 0 0 vdda
port 9 nsew
flabel metal4 s 0 7910 254 8840 3 FreeSans 520 0 0 0 vssd
port 10 nsew
flabel metal5 s 9346 3570 9600 4460 3 FreeSans 520 180 0 0 vddio
port 1 nsew
flabel metal5 s 9346 20 9600 1070 3 FreeSans 520 180 0 0 vcchib
port 6 nsew
flabel metal5 s 9346 13600 9600 18590 3 FreeSans 520 180 0 0 vddio
port 1 nsew
flabel metal5 s 9346 12430 9600 13280 3 FreeSans 520 180 0 0 vddio_q
port 4 nsew
flabel metal5 s 9346 1390 9600 2280 3 FreeSans 520 180 0 0 vccd
port 3 nsew
flabel metal5 s 9346 6961 9600 7610 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal5 s 9346 5990 9600 6640 3 FreeSans 520 180 0 0 vswitch
port 7 nsew
flabel metal5 s 9346 4780 9600 5670 3 FreeSans 520 180 0 0 vssio
port 2 nsew
flabel metal5 s 9346 11260 9600 12110 3 FreeSans 520 180 0 0 vssio_q
port 8 nsew
flabel metal5 s 9346 7930 9600 8820 3 FreeSans 520 180 0 0 vssd
port 10 nsew
flabel metal5 s 9407 2600 9600 3250 3 FreeSans 520 180 0 0 vdda
port 9 nsew
flabel metal5 s 9346 9140 9600 10940 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal5 s 9346 34750 9600 39593 3 FreeSans 520 180 0 0 vssio
port 2 nsew
flabel metal5 s 0 3570 254 4460 3 FreeSans 520 0 0 0 vddio
port 1 nsew
flabel metal5 s 0 20 254 1070 3 FreeSans 520 0 0 0 vcchib
port 6 nsew
flabel metal5 s 0 13600 254 18590 3 FreeSans 520 0 0 0 vddio
port 1 nsew
flabel metal5 s 0 12430 254 13280 3 FreeSans 520 0 0 0 vddio_q
port 4 nsew
flabel metal5 s 0 1390 254 2280 3 FreeSans 520 0 0 0 vccd
port 3 nsew
flabel metal5 s 0 6961 254 7610 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal5 s 0 5990 254 6640 3 FreeSans 520 0 0 0 vswitch
port 7 nsew
flabel metal5 s 0 4780 254 5670 3 FreeSans 520 0 0 0 vssio
port 2 nsew
flabel metal5 s 0 11260 254 12110 3 FreeSans 520 0 0 0 vssio_q
port 8 nsew
flabel metal5 s 0 7930 254 8820 3 FreeSans 520 0 0 0 vssd
port 10 nsew
flabel metal5 s 0 2600 193 3250 3 FreeSans 520 0 0 0 vdda
port 9 nsew
flabel metal5 s 0 9140 254 10940 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal5 s 0 34750 254 39593 3 FreeSans 520 0 0 0 vssio
port 2 nsew
<< properties >>
string GDS_END 644756
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 540264
<< end >>
