magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< metal3 >>
rect 99 3672 4879 3676
rect 99 3608 105 3672
rect 169 3608 187 3672
rect 251 3608 269 3672
rect 333 3608 351 3672
rect 415 3608 433 3672
rect 497 3608 515 3672
rect 579 3608 597 3672
rect 661 3608 678 3672
rect 742 3608 759 3672
rect 823 3608 840 3672
rect 904 3608 921 3672
rect 985 3608 1002 3672
rect 1066 3608 1083 3672
rect 1147 3608 1164 3672
rect 1228 3608 1245 3672
rect 1309 3608 1326 3672
rect 1390 3608 1407 3672
rect 1471 3608 1488 3672
rect 1552 3608 1569 3672
rect 1633 3608 1650 3672
rect 1714 3608 1731 3672
rect 1795 3608 1812 3672
rect 1876 3608 1893 3672
rect 1957 3608 1974 3672
rect 2038 3608 2055 3672
rect 2119 3608 2136 3672
rect 2200 3608 2217 3672
rect 2281 3608 2298 3672
rect 2362 3608 2379 3672
rect 2443 3608 2460 3672
rect 2524 3608 2541 3672
rect 2605 3608 2622 3672
rect 2686 3608 2703 3672
rect 2767 3608 2784 3672
rect 2848 3608 2865 3672
rect 2929 3608 2946 3672
rect 3010 3608 3027 3672
rect 3091 3608 3108 3672
rect 3172 3608 3189 3672
rect 3253 3608 3270 3672
rect 3334 3608 3351 3672
rect 3415 3608 3432 3672
rect 3496 3608 3513 3672
rect 3577 3608 3594 3672
rect 3658 3608 3675 3672
rect 3739 3608 3756 3672
rect 3820 3608 3837 3672
rect 3901 3608 3918 3672
rect 3982 3608 3999 3672
rect 4063 3608 4080 3672
rect 4144 3608 4161 3672
rect 4225 3608 4242 3672
rect 4306 3608 4323 3672
rect 4387 3608 4404 3672
rect 4468 3608 4485 3672
rect 4549 3608 4566 3672
rect 4630 3608 4647 3672
rect 4711 3608 4728 3672
rect 4792 3608 4809 3672
rect 4873 3608 4879 3672
rect 99 3584 4879 3608
rect 99 3520 105 3584
rect 169 3520 187 3584
rect 251 3520 269 3584
rect 333 3520 351 3584
rect 415 3520 433 3584
rect 497 3520 515 3584
rect 579 3520 597 3584
rect 661 3520 678 3584
rect 742 3520 759 3584
rect 823 3520 840 3584
rect 904 3520 921 3584
rect 985 3520 1002 3584
rect 1066 3520 1083 3584
rect 1147 3520 1164 3584
rect 1228 3520 1245 3584
rect 1309 3520 1326 3584
rect 1390 3520 1407 3584
rect 1471 3520 1488 3584
rect 1552 3520 1569 3584
rect 1633 3520 1650 3584
rect 1714 3520 1731 3584
rect 1795 3520 1812 3584
rect 1876 3520 1893 3584
rect 1957 3520 1974 3584
rect 2038 3520 2055 3584
rect 2119 3520 2136 3584
rect 2200 3520 2217 3584
rect 2281 3520 2298 3584
rect 2362 3520 2379 3584
rect 2443 3520 2460 3584
rect 2524 3520 2541 3584
rect 2605 3520 2622 3584
rect 2686 3520 2703 3584
rect 2767 3520 2784 3584
rect 2848 3520 2865 3584
rect 2929 3520 2946 3584
rect 3010 3520 3027 3584
rect 3091 3520 3108 3584
rect 3172 3520 3189 3584
rect 3253 3520 3270 3584
rect 3334 3520 3351 3584
rect 3415 3520 3432 3584
rect 3496 3520 3513 3584
rect 3577 3520 3594 3584
rect 3658 3520 3675 3584
rect 3739 3520 3756 3584
rect 3820 3520 3837 3584
rect 3901 3520 3918 3584
rect 3982 3520 3999 3584
rect 4063 3520 4080 3584
rect 4144 3520 4161 3584
rect 4225 3520 4242 3584
rect 4306 3520 4323 3584
rect 4387 3520 4404 3584
rect 4468 3520 4485 3584
rect 4549 3520 4566 3584
rect 4630 3520 4647 3584
rect 4711 3520 4728 3584
rect 4792 3520 4809 3584
rect 4873 3520 4879 3584
rect 99 3496 4879 3520
rect 99 3432 105 3496
rect 169 3432 187 3496
rect 251 3432 269 3496
rect 333 3432 351 3496
rect 415 3432 433 3496
rect 497 3432 515 3496
rect 579 3432 597 3496
rect 661 3432 678 3496
rect 742 3432 759 3496
rect 823 3432 840 3496
rect 904 3432 921 3496
rect 985 3432 1002 3496
rect 1066 3432 1083 3496
rect 1147 3432 1164 3496
rect 1228 3432 1245 3496
rect 1309 3432 1326 3496
rect 1390 3432 1407 3496
rect 1471 3432 1488 3496
rect 1552 3432 1569 3496
rect 1633 3432 1650 3496
rect 1714 3432 1731 3496
rect 1795 3432 1812 3496
rect 1876 3432 1893 3496
rect 1957 3432 1974 3496
rect 2038 3432 2055 3496
rect 2119 3432 2136 3496
rect 2200 3432 2217 3496
rect 2281 3432 2298 3496
rect 2362 3432 2379 3496
rect 2443 3432 2460 3496
rect 2524 3432 2541 3496
rect 2605 3432 2622 3496
rect 2686 3432 2703 3496
rect 2767 3432 2784 3496
rect 2848 3432 2865 3496
rect 2929 3432 2946 3496
rect 3010 3432 3027 3496
rect 3091 3432 3108 3496
rect 3172 3432 3189 3496
rect 3253 3432 3270 3496
rect 3334 3432 3351 3496
rect 3415 3432 3432 3496
rect 3496 3432 3513 3496
rect 3577 3432 3594 3496
rect 3658 3432 3675 3496
rect 3739 3432 3756 3496
rect 3820 3432 3837 3496
rect 3901 3432 3918 3496
rect 3982 3432 3999 3496
rect 4063 3432 4080 3496
rect 4144 3432 4161 3496
rect 4225 3432 4242 3496
rect 4306 3432 4323 3496
rect 4387 3432 4404 3496
rect 4468 3432 4485 3496
rect 4549 3432 4566 3496
rect 4630 3432 4647 3496
rect 4711 3432 4728 3496
rect 4792 3432 4809 3496
rect 4873 3432 4879 3496
rect 99 3408 4879 3432
rect 99 3344 105 3408
rect 169 3344 187 3408
rect 251 3344 269 3408
rect 333 3344 351 3408
rect 415 3344 433 3408
rect 497 3344 515 3408
rect 579 3344 597 3408
rect 661 3344 678 3408
rect 742 3344 759 3408
rect 823 3344 840 3408
rect 904 3344 921 3408
rect 985 3344 1002 3408
rect 1066 3344 1083 3408
rect 1147 3344 1164 3408
rect 1228 3344 1245 3408
rect 1309 3344 1326 3408
rect 1390 3344 1407 3408
rect 1471 3344 1488 3408
rect 1552 3344 1569 3408
rect 1633 3344 1650 3408
rect 1714 3344 1731 3408
rect 1795 3344 1812 3408
rect 1876 3344 1893 3408
rect 1957 3344 1974 3408
rect 2038 3344 2055 3408
rect 2119 3344 2136 3408
rect 2200 3344 2217 3408
rect 2281 3344 2298 3408
rect 2362 3344 2379 3408
rect 2443 3344 2460 3408
rect 2524 3344 2541 3408
rect 2605 3344 2622 3408
rect 2686 3344 2703 3408
rect 2767 3344 2784 3408
rect 2848 3344 2865 3408
rect 2929 3344 2946 3408
rect 3010 3344 3027 3408
rect 3091 3344 3108 3408
rect 3172 3344 3189 3408
rect 3253 3344 3270 3408
rect 3334 3344 3351 3408
rect 3415 3344 3432 3408
rect 3496 3344 3513 3408
rect 3577 3344 3594 3408
rect 3658 3344 3675 3408
rect 3739 3344 3756 3408
rect 3820 3344 3837 3408
rect 3901 3344 3918 3408
rect 3982 3344 3999 3408
rect 4063 3344 4080 3408
rect 4144 3344 4161 3408
rect 4225 3344 4242 3408
rect 4306 3344 4323 3408
rect 4387 3344 4404 3408
rect 4468 3344 4485 3408
rect 4549 3344 4566 3408
rect 4630 3344 4647 3408
rect 4711 3344 4728 3408
rect 4792 3344 4809 3408
rect 4873 3344 4879 3408
rect 99 3320 4879 3344
rect 99 3256 105 3320
rect 169 3256 187 3320
rect 251 3256 269 3320
rect 333 3256 351 3320
rect 415 3256 433 3320
rect 497 3256 515 3320
rect 579 3256 597 3320
rect 661 3256 678 3320
rect 742 3256 759 3320
rect 823 3256 840 3320
rect 904 3256 921 3320
rect 985 3256 1002 3320
rect 1066 3256 1083 3320
rect 1147 3256 1164 3320
rect 1228 3256 1245 3320
rect 1309 3256 1326 3320
rect 1390 3256 1407 3320
rect 1471 3256 1488 3320
rect 1552 3256 1569 3320
rect 1633 3256 1650 3320
rect 1714 3256 1731 3320
rect 1795 3256 1812 3320
rect 1876 3256 1893 3320
rect 1957 3256 1974 3320
rect 2038 3256 2055 3320
rect 2119 3256 2136 3320
rect 2200 3256 2217 3320
rect 2281 3256 2298 3320
rect 2362 3256 2379 3320
rect 2443 3256 2460 3320
rect 2524 3256 2541 3320
rect 2605 3256 2622 3320
rect 2686 3256 2703 3320
rect 2767 3256 2784 3320
rect 2848 3256 2865 3320
rect 2929 3256 2946 3320
rect 3010 3256 3027 3320
rect 3091 3256 3108 3320
rect 3172 3256 3189 3320
rect 3253 3256 3270 3320
rect 3334 3256 3351 3320
rect 3415 3256 3432 3320
rect 3496 3256 3513 3320
rect 3577 3256 3594 3320
rect 3658 3256 3675 3320
rect 3739 3256 3756 3320
rect 3820 3256 3837 3320
rect 3901 3256 3918 3320
rect 3982 3256 3999 3320
rect 4063 3256 4080 3320
rect 4144 3256 4161 3320
rect 4225 3256 4242 3320
rect 4306 3256 4323 3320
rect 4387 3256 4404 3320
rect 4468 3256 4485 3320
rect 4549 3256 4566 3320
rect 4630 3256 4647 3320
rect 4711 3256 4728 3320
rect 4792 3256 4809 3320
rect 4873 3256 4879 3320
rect 99 3232 4879 3256
rect 99 3168 105 3232
rect 169 3168 187 3232
rect 251 3168 269 3232
rect 333 3168 351 3232
rect 415 3168 433 3232
rect 497 3168 515 3232
rect 579 3168 597 3232
rect 661 3168 678 3232
rect 742 3168 759 3232
rect 823 3168 840 3232
rect 904 3168 921 3232
rect 985 3168 1002 3232
rect 1066 3168 1083 3232
rect 1147 3168 1164 3232
rect 1228 3168 1245 3232
rect 1309 3168 1326 3232
rect 1390 3168 1407 3232
rect 1471 3168 1488 3232
rect 1552 3168 1569 3232
rect 1633 3168 1650 3232
rect 1714 3168 1731 3232
rect 1795 3168 1812 3232
rect 1876 3168 1893 3232
rect 1957 3168 1974 3232
rect 2038 3168 2055 3232
rect 2119 3168 2136 3232
rect 2200 3168 2217 3232
rect 2281 3168 2298 3232
rect 2362 3168 2379 3232
rect 2443 3168 2460 3232
rect 2524 3168 2541 3232
rect 2605 3168 2622 3232
rect 2686 3168 2703 3232
rect 2767 3168 2784 3232
rect 2848 3168 2865 3232
rect 2929 3168 2946 3232
rect 3010 3168 3027 3232
rect 3091 3168 3108 3232
rect 3172 3168 3189 3232
rect 3253 3168 3270 3232
rect 3334 3168 3351 3232
rect 3415 3168 3432 3232
rect 3496 3168 3513 3232
rect 3577 3168 3594 3232
rect 3658 3168 3675 3232
rect 3739 3168 3756 3232
rect 3820 3168 3837 3232
rect 3901 3168 3918 3232
rect 3982 3168 3999 3232
rect 4063 3168 4080 3232
rect 4144 3168 4161 3232
rect 4225 3168 4242 3232
rect 4306 3168 4323 3232
rect 4387 3168 4404 3232
rect 4468 3168 4485 3232
rect 4549 3168 4566 3232
rect 4630 3168 4647 3232
rect 4711 3168 4728 3232
rect 4792 3168 4809 3232
rect 4873 3168 4879 3232
rect 99 3144 4879 3168
rect 99 3080 105 3144
rect 169 3080 187 3144
rect 251 3080 269 3144
rect 333 3080 351 3144
rect 415 3080 433 3144
rect 497 3080 515 3144
rect 579 3080 597 3144
rect 661 3080 678 3144
rect 742 3080 759 3144
rect 823 3080 840 3144
rect 904 3080 921 3144
rect 985 3080 1002 3144
rect 1066 3080 1083 3144
rect 1147 3080 1164 3144
rect 1228 3080 1245 3144
rect 1309 3080 1326 3144
rect 1390 3080 1407 3144
rect 1471 3080 1488 3144
rect 1552 3080 1569 3144
rect 1633 3080 1650 3144
rect 1714 3080 1731 3144
rect 1795 3080 1812 3144
rect 1876 3080 1893 3144
rect 1957 3080 1974 3144
rect 2038 3080 2055 3144
rect 2119 3080 2136 3144
rect 2200 3080 2217 3144
rect 2281 3080 2298 3144
rect 2362 3080 2379 3144
rect 2443 3080 2460 3144
rect 2524 3080 2541 3144
rect 2605 3080 2622 3144
rect 2686 3080 2703 3144
rect 2767 3080 2784 3144
rect 2848 3080 2865 3144
rect 2929 3080 2946 3144
rect 3010 3080 3027 3144
rect 3091 3080 3108 3144
rect 3172 3080 3189 3144
rect 3253 3080 3270 3144
rect 3334 3080 3351 3144
rect 3415 3080 3432 3144
rect 3496 3080 3513 3144
rect 3577 3080 3594 3144
rect 3658 3080 3675 3144
rect 3739 3080 3756 3144
rect 3820 3080 3837 3144
rect 3901 3080 3918 3144
rect 3982 3080 3999 3144
rect 4063 3080 4080 3144
rect 4144 3080 4161 3144
rect 4225 3080 4242 3144
rect 4306 3080 4323 3144
rect 4387 3080 4404 3144
rect 4468 3080 4485 3144
rect 4549 3080 4566 3144
rect 4630 3080 4647 3144
rect 4711 3080 4728 3144
rect 4792 3080 4809 3144
rect 4873 3080 4879 3144
rect 99 3056 4879 3080
rect 99 2992 105 3056
rect 169 2992 187 3056
rect 251 2992 269 3056
rect 333 2992 351 3056
rect 415 2992 433 3056
rect 497 2992 515 3056
rect 579 2992 597 3056
rect 661 2992 678 3056
rect 742 2992 759 3056
rect 823 2992 840 3056
rect 904 2992 921 3056
rect 985 2992 1002 3056
rect 1066 2992 1083 3056
rect 1147 2992 1164 3056
rect 1228 2992 1245 3056
rect 1309 2992 1326 3056
rect 1390 2992 1407 3056
rect 1471 2992 1488 3056
rect 1552 2992 1569 3056
rect 1633 2992 1650 3056
rect 1714 2992 1731 3056
rect 1795 2992 1812 3056
rect 1876 2992 1893 3056
rect 1957 2992 1974 3056
rect 2038 2992 2055 3056
rect 2119 2992 2136 3056
rect 2200 2992 2217 3056
rect 2281 2992 2298 3056
rect 2362 2992 2379 3056
rect 2443 2992 2460 3056
rect 2524 2992 2541 3056
rect 2605 2992 2622 3056
rect 2686 2992 2703 3056
rect 2767 2992 2784 3056
rect 2848 2992 2865 3056
rect 2929 2992 2946 3056
rect 3010 2992 3027 3056
rect 3091 2992 3108 3056
rect 3172 2992 3189 3056
rect 3253 2992 3270 3056
rect 3334 2992 3351 3056
rect 3415 2992 3432 3056
rect 3496 2992 3513 3056
rect 3577 2992 3594 3056
rect 3658 2992 3675 3056
rect 3739 2992 3756 3056
rect 3820 2992 3837 3056
rect 3901 2992 3918 3056
rect 3982 2992 3999 3056
rect 4063 2992 4080 3056
rect 4144 2992 4161 3056
rect 4225 2992 4242 3056
rect 4306 2992 4323 3056
rect 4387 2992 4404 3056
rect 4468 2992 4485 3056
rect 4549 2992 4566 3056
rect 4630 2992 4647 3056
rect 4711 2992 4728 3056
rect 4792 2992 4809 3056
rect 4873 2992 4879 3056
rect 99 2988 4879 2992
rect 10078 3672 14858 3676
rect 10078 3608 10084 3672
rect 10148 3608 10166 3672
rect 10230 3608 10248 3672
rect 10312 3608 10330 3672
rect 10394 3608 10412 3672
rect 10476 3608 10494 3672
rect 10558 3608 10576 3672
rect 10640 3608 10657 3672
rect 10721 3608 10738 3672
rect 10802 3608 10819 3672
rect 10883 3608 10900 3672
rect 10964 3608 10981 3672
rect 11045 3608 11062 3672
rect 11126 3608 11143 3672
rect 11207 3608 11224 3672
rect 11288 3608 11305 3672
rect 11369 3608 11386 3672
rect 11450 3608 11467 3672
rect 11531 3608 11548 3672
rect 11612 3608 11629 3672
rect 11693 3608 11710 3672
rect 11774 3608 11791 3672
rect 11855 3608 11872 3672
rect 11936 3608 11953 3672
rect 12017 3608 12034 3672
rect 12098 3608 12115 3672
rect 12179 3608 12196 3672
rect 12260 3608 12277 3672
rect 12341 3608 12358 3672
rect 12422 3608 12439 3672
rect 12503 3608 12520 3672
rect 12584 3608 12601 3672
rect 12665 3608 12682 3672
rect 12746 3608 12763 3672
rect 12827 3608 12844 3672
rect 12908 3608 12925 3672
rect 12989 3608 13006 3672
rect 13070 3608 13087 3672
rect 13151 3608 13168 3672
rect 13232 3608 13249 3672
rect 13313 3608 13330 3672
rect 13394 3608 13411 3672
rect 13475 3608 13492 3672
rect 13556 3608 13573 3672
rect 13637 3608 13654 3672
rect 13718 3608 13735 3672
rect 13799 3608 13816 3672
rect 13880 3608 13897 3672
rect 13961 3608 13978 3672
rect 14042 3608 14059 3672
rect 14123 3608 14140 3672
rect 14204 3608 14221 3672
rect 14285 3608 14302 3672
rect 14366 3608 14383 3672
rect 14447 3608 14464 3672
rect 14528 3608 14545 3672
rect 14609 3608 14626 3672
rect 14690 3608 14707 3672
rect 14771 3608 14788 3672
rect 14852 3608 14858 3672
rect 10078 3584 14858 3608
rect 10078 3520 10084 3584
rect 10148 3520 10166 3584
rect 10230 3520 10248 3584
rect 10312 3520 10330 3584
rect 10394 3520 10412 3584
rect 10476 3520 10494 3584
rect 10558 3520 10576 3584
rect 10640 3520 10657 3584
rect 10721 3520 10738 3584
rect 10802 3520 10819 3584
rect 10883 3520 10900 3584
rect 10964 3520 10981 3584
rect 11045 3520 11062 3584
rect 11126 3520 11143 3584
rect 11207 3520 11224 3584
rect 11288 3520 11305 3584
rect 11369 3520 11386 3584
rect 11450 3520 11467 3584
rect 11531 3520 11548 3584
rect 11612 3520 11629 3584
rect 11693 3520 11710 3584
rect 11774 3520 11791 3584
rect 11855 3520 11872 3584
rect 11936 3520 11953 3584
rect 12017 3520 12034 3584
rect 12098 3520 12115 3584
rect 12179 3520 12196 3584
rect 12260 3520 12277 3584
rect 12341 3520 12358 3584
rect 12422 3520 12439 3584
rect 12503 3520 12520 3584
rect 12584 3520 12601 3584
rect 12665 3520 12682 3584
rect 12746 3520 12763 3584
rect 12827 3520 12844 3584
rect 12908 3520 12925 3584
rect 12989 3520 13006 3584
rect 13070 3520 13087 3584
rect 13151 3520 13168 3584
rect 13232 3520 13249 3584
rect 13313 3520 13330 3584
rect 13394 3520 13411 3584
rect 13475 3520 13492 3584
rect 13556 3520 13573 3584
rect 13637 3520 13654 3584
rect 13718 3520 13735 3584
rect 13799 3520 13816 3584
rect 13880 3520 13897 3584
rect 13961 3520 13978 3584
rect 14042 3520 14059 3584
rect 14123 3520 14140 3584
rect 14204 3520 14221 3584
rect 14285 3520 14302 3584
rect 14366 3520 14383 3584
rect 14447 3520 14464 3584
rect 14528 3520 14545 3584
rect 14609 3520 14626 3584
rect 14690 3520 14707 3584
rect 14771 3520 14788 3584
rect 14852 3520 14858 3584
rect 10078 3496 14858 3520
rect 10078 3432 10084 3496
rect 10148 3432 10166 3496
rect 10230 3432 10248 3496
rect 10312 3432 10330 3496
rect 10394 3432 10412 3496
rect 10476 3432 10494 3496
rect 10558 3432 10576 3496
rect 10640 3432 10657 3496
rect 10721 3432 10738 3496
rect 10802 3432 10819 3496
rect 10883 3432 10900 3496
rect 10964 3432 10981 3496
rect 11045 3432 11062 3496
rect 11126 3432 11143 3496
rect 11207 3432 11224 3496
rect 11288 3432 11305 3496
rect 11369 3432 11386 3496
rect 11450 3432 11467 3496
rect 11531 3432 11548 3496
rect 11612 3432 11629 3496
rect 11693 3432 11710 3496
rect 11774 3432 11791 3496
rect 11855 3432 11872 3496
rect 11936 3432 11953 3496
rect 12017 3432 12034 3496
rect 12098 3432 12115 3496
rect 12179 3432 12196 3496
rect 12260 3432 12277 3496
rect 12341 3432 12358 3496
rect 12422 3432 12439 3496
rect 12503 3432 12520 3496
rect 12584 3432 12601 3496
rect 12665 3432 12682 3496
rect 12746 3432 12763 3496
rect 12827 3432 12844 3496
rect 12908 3432 12925 3496
rect 12989 3432 13006 3496
rect 13070 3432 13087 3496
rect 13151 3432 13168 3496
rect 13232 3432 13249 3496
rect 13313 3432 13330 3496
rect 13394 3432 13411 3496
rect 13475 3432 13492 3496
rect 13556 3432 13573 3496
rect 13637 3432 13654 3496
rect 13718 3432 13735 3496
rect 13799 3432 13816 3496
rect 13880 3432 13897 3496
rect 13961 3432 13978 3496
rect 14042 3432 14059 3496
rect 14123 3432 14140 3496
rect 14204 3432 14221 3496
rect 14285 3432 14302 3496
rect 14366 3432 14383 3496
rect 14447 3432 14464 3496
rect 14528 3432 14545 3496
rect 14609 3432 14626 3496
rect 14690 3432 14707 3496
rect 14771 3432 14788 3496
rect 14852 3432 14858 3496
rect 10078 3408 14858 3432
rect 10078 3344 10084 3408
rect 10148 3344 10166 3408
rect 10230 3344 10248 3408
rect 10312 3344 10330 3408
rect 10394 3344 10412 3408
rect 10476 3344 10494 3408
rect 10558 3344 10576 3408
rect 10640 3344 10657 3408
rect 10721 3344 10738 3408
rect 10802 3344 10819 3408
rect 10883 3344 10900 3408
rect 10964 3344 10981 3408
rect 11045 3344 11062 3408
rect 11126 3344 11143 3408
rect 11207 3344 11224 3408
rect 11288 3344 11305 3408
rect 11369 3344 11386 3408
rect 11450 3344 11467 3408
rect 11531 3344 11548 3408
rect 11612 3344 11629 3408
rect 11693 3344 11710 3408
rect 11774 3344 11791 3408
rect 11855 3344 11872 3408
rect 11936 3344 11953 3408
rect 12017 3344 12034 3408
rect 12098 3344 12115 3408
rect 12179 3344 12196 3408
rect 12260 3344 12277 3408
rect 12341 3344 12358 3408
rect 12422 3344 12439 3408
rect 12503 3344 12520 3408
rect 12584 3344 12601 3408
rect 12665 3344 12682 3408
rect 12746 3344 12763 3408
rect 12827 3344 12844 3408
rect 12908 3344 12925 3408
rect 12989 3344 13006 3408
rect 13070 3344 13087 3408
rect 13151 3344 13168 3408
rect 13232 3344 13249 3408
rect 13313 3344 13330 3408
rect 13394 3344 13411 3408
rect 13475 3344 13492 3408
rect 13556 3344 13573 3408
rect 13637 3344 13654 3408
rect 13718 3344 13735 3408
rect 13799 3344 13816 3408
rect 13880 3344 13897 3408
rect 13961 3344 13978 3408
rect 14042 3344 14059 3408
rect 14123 3344 14140 3408
rect 14204 3344 14221 3408
rect 14285 3344 14302 3408
rect 14366 3344 14383 3408
rect 14447 3344 14464 3408
rect 14528 3344 14545 3408
rect 14609 3344 14626 3408
rect 14690 3344 14707 3408
rect 14771 3344 14788 3408
rect 14852 3344 14858 3408
rect 10078 3320 14858 3344
rect 10078 3256 10084 3320
rect 10148 3256 10166 3320
rect 10230 3256 10248 3320
rect 10312 3256 10330 3320
rect 10394 3256 10412 3320
rect 10476 3256 10494 3320
rect 10558 3256 10576 3320
rect 10640 3256 10657 3320
rect 10721 3256 10738 3320
rect 10802 3256 10819 3320
rect 10883 3256 10900 3320
rect 10964 3256 10981 3320
rect 11045 3256 11062 3320
rect 11126 3256 11143 3320
rect 11207 3256 11224 3320
rect 11288 3256 11305 3320
rect 11369 3256 11386 3320
rect 11450 3256 11467 3320
rect 11531 3256 11548 3320
rect 11612 3256 11629 3320
rect 11693 3256 11710 3320
rect 11774 3256 11791 3320
rect 11855 3256 11872 3320
rect 11936 3256 11953 3320
rect 12017 3256 12034 3320
rect 12098 3256 12115 3320
rect 12179 3256 12196 3320
rect 12260 3256 12277 3320
rect 12341 3256 12358 3320
rect 12422 3256 12439 3320
rect 12503 3256 12520 3320
rect 12584 3256 12601 3320
rect 12665 3256 12682 3320
rect 12746 3256 12763 3320
rect 12827 3256 12844 3320
rect 12908 3256 12925 3320
rect 12989 3256 13006 3320
rect 13070 3256 13087 3320
rect 13151 3256 13168 3320
rect 13232 3256 13249 3320
rect 13313 3256 13330 3320
rect 13394 3256 13411 3320
rect 13475 3256 13492 3320
rect 13556 3256 13573 3320
rect 13637 3256 13654 3320
rect 13718 3256 13735 3320
rect 13799 3256 13816 3320
rect 13880 3256 13897 3320
rect 13961 3256 13978 3320
rect 14042 3256 14059 3320
rect 14123 3256 14140 3320
rect 14204 3256 14221 3320
rect 14285 3256 14302 3320
rect 14366 3256 14383 3320
rect 14447 3256 14464 3320
rect 14528 3256 14545 3320
rect 14609 3256 14626 3320
rect 14690 3256 14707 3320
rect 14771 3256 14788 3320
rect 14852 3256 14858 3320
rect 10078 3232 14858 3256
rect 10078 3168 10084 3232
rect 10148 3168 10166 3232
rect 10230 3168 10248 3232
rect 10312 3168 10330 3232
rect 10394 3168 10412 3232
rect 10476 3168 10494 3232
rect 10558 3168 10576 3232
rect 10640 3168 10657 3232
rect 10721 3168 10738 3232
rect 10802 3168 10819 3232
rect 10883 3168 10900 3232
rect 10964 3168 10981 3232
rect 11045 3168 11062 3232
rect 11126 3168 11143 3232
rect 11207 3168 11224 3232
rect 11288 3168 11305 3232
rect 11369 3168 11386 3232
rect 11450 3168 11467 3232
rect 11531 3168 11548 3232
rect 11612 3168 11629 3232
rect 11693 3168 11710 3232
rect 11774 3168 11791 3232
rect 11855 3168 11872 3232
rect 11936 3168 11953 3232
rect 12017 3168 12034 3232
rect 12098 3168 12115 3232
rect 12179 3168 12196 3232
rect 12260 3168 12277 3232
rect 12341 3168 12358 3232
rect 12422 3168 12439 3232
rect 12503 3168 12520 3232
rect 12584 3168 12601 3232
rect 12665 3168 12682 3232
rect 12746 3168 12763 3232
rect 12827 3168 12844 3232
rect 12908 3168 12925 3232
rect 12989 3168 13006 3232
rect 13070 3168 13087 3232
rect 13151 3168 13168 3232
rect 13232 3168 13249 3232
rect 13313 3168 13330 3232
rect 13394 3168 13411 3232
rect 13475 3168 13492 3232
rect 13556 3168 13573 3232
rect 13637 3168 13654 3232
rect 13718 3168 13735 3232
rect 13799 3168 13816 3232
rect 13880 3168 13897 3232
rect 13961 3168 13978 3232
rect 14042 3168 14059 3232
rect 14123 3168 14140 3232
rect 14204 3168 14221 3232
rect 14285 3168 14302 3232
rect 14366 3168 14383 3232
rect 14447 3168 14464 3232
rect 14528 3168 14545 3232
rect 14609 3168 14626 3232
rect 14690 3168 14707 3232
rect 14771 3168 14788 3232
rect 14852 3168 14858 3232
rect 10078 3144 14858 3168
rect 10078 3080 10084 3144
rect 10148 3080 10166 3144
rect 10230 3080 10248 3144
rect 10312 3080 10330 3144
rect 10394 3080 10412 3144
rect 10476 3080 10494 3144
rect 10558 3080 10576 3144
rect 10640 3080 10657 3144
rect 10721 3080 10738 3144
rect 10802 3080 10819 3144
rect 10883 3080 10900 3144
rect 10964 3080 10981 3144
rect 11045 3080 11062 3144
rect 11126 3080 11143 3144
rect 11207 3080 11224 3144
rect 11288 3080 11305 3144
rect 11369 3080 11386 3144
rect 11450 3080 11467 3144
rect 11531 3080 11548 3144
rect 11612 3080 11629 3144
rect 11693 3080 11710 3144
rect 11774 3080 11791 3144
rect 11855 3080 11872 3144
rect 11936 3080 11953 3144
rect 12017 3080 12034 3144
rect 12098 3080 12115 3144
rect 12179 3080 12196 3144
rect 12260 3080 12277 3144
rect 12341 3080 12358 3144
rect 12422 3080 12439 3144
rect 12503 3080 12520 3144
rect 12584 3080 12601 3144
rect 12665 3080 12682 3144
rect 12746 3080 12763 3144
rect 12827 3080 12844 3144
rect 12908 3080 12925 3144
rect 12989 3080 13006 3144
rect 13070 3080 13087 3144
rect 13151 3080 13168 3144
rect 13232 3080 13249 3144
rect 13313 3080 13330 3144
rect 13394 3080 13411 3144
rect 13475 3080 13492 3144
rect 13556 3080 13573 3144
rect 13637 3080 13654 3144
rect 13718 3080 13735 3144
rect 13799 3080 13816 3144
rect 13880 3080 13897 3144
rect 13961 3080 13978 3144
rect 14042 3080 14059 3144
rect 14123 3080 14140 3144
rect 14204 3080 14221 3144
rect 14285 3080 14302 3144
rect 14366 3080 14383 3144
rect 14447 3080 14464 3144
rect 14528 3080 14545 3144
rect 14609 3080 14626 3144
rect 14690 3080 14707 3144
rect 14771 3080 14788 3144
rect 14852 3080 14858 3144
rect 10078 3056 14858 3080
rect 10078 2992 10084 3056
rect 10148 2992 10166 3056
rect 10230 2992 10248 3056
rect 10312 2992 10330 3056
rect 10394 2992 10412 3056
rect 10476 2992 10494 3056
rect 10558 2992 10576 3056
rect 10640 2992 10657 3056
rect 10721 2992 10738 3056
rect 10802 2992 10819 3056
rect 10883 2992 10900 3056
rect 10964 2992 10981 3056
rect 11045 2992 11062 3056
rect 11126 2992 11143 3056
rect 11207 2992 11224 3056
rect 11288 2992 11305 3056
rect 11369 2992 11386 3056
rect 11450 2992 11467 3056
rect 11531 2992 11548 3056
rect 11612 2992 11629 3056
rect 11693 2992 11710 3056
rect 11774 2992 11791 3056
rect 11855 2992 11872 3056
rect 11936 2992 11953 3056
rect 12017 2992 12034 3056
rect 12098 2992 12115 3056
rect 12179 2992 12196 3056
rect 12260 2992 12277 3056
rect 12341 2992 12358 3056
rect 12422 2992 12439 3056
rect 12503 2992 12520 3056
rect 12584 2992 12601 3056
rect 12665 2992 12682 3056
rect 12746 2992 12763 3056
rect 12827 2992 12844 3056
rect 12908 2992 12925 3056
rect 12989 2992 13006 3056
rect 13070 2992 13087 3056
rect 13151 2992 13168 3056
rect 13232 2992 13249 3056
rect 13313 2992 13330 3056
rect 13394 2992 13411 3056
rect 13475 2992 13492 3056
rect 13556 2992 13573 3056
rect 13637 2992 13654 3056
rect 13718 2992 13735 3056
rect 13799 2992 13816 3056
rect 13880 2992 13897 3056
rect 13961 2992 13978 3056
rect 14042 2992 14059 3056
rect 14123 2992 14140 3056
rect 14204 2992 14221 3056
rect 14285 2992 14302 3056
rect 14366 2992 14383 3056
rect 14447 2992 14464 3056
rect 14528 2992 14545 3056
rect 14609 2992 14626 3056
rect 14690 2992 14707 3056
rect 14771 2992 14788 3056
rect 14852 2992 14858 3056
rect 10078 2988 14858 2992
<< via3 >>
rect 105 3608 169 3672
rect 187 3608 251 3672
rect 269 3608 333 3672
rect 351 3608 415 3672
rect 433 3608 497 3672
rect 515 3608 579 3672
rect 597 3608 661 3672
rect 678 3608 742 3672
rect 759 3608 823 3672
rect 840 3608 904 3672
rect 921 3608 985 3672
rect 1002 3608 1066 3672
rect 1083 3608 1147 3672
rect 1164 3608 1228 3672
rect 1245 3608 1309 3672
rect 1326 3608 1390 3672
rect 1407 3608 1471 3672
rect 1488 3608 1552 3672
rect 1569 3608 1633 3672
rect 1650 3608 1714 3672
rect 1731 3608 1795 3672
rect 1812 3608 1876 3672
rect 1893 3608 1957 3672
rect 1974 3608 2038 3672
rect 2055 3608 2119 3672
rect 2136 3608 2200 3672
rect 2217 3608 2281 3672
rect 2298 3608 2362 3672
rect 2379 3608 2443 3672
rect 2460 3608 2524 3672
rect 2541 3608 2605 3672
rect 2622 3608 2686 3672
rect 2703 3608 2767 3672
rect 2784 3608 2848 3672
rect 2865 3608 2929 3672
rect 2946 3608 3010 3672
rect 3027 3608 3091 3672
rect 3108 3608 3172 3672
rect 3189 3608 3253 3672
rect 3270 3608 3334 3672
rect 3351 3608 3415 3672
rect 3432 3608 3496 3672
rect 3513 3608 3577 3672
rect 3594 3608 3658 3672
rect 3675 3608 3739 3672
rect 3756 3608 3820 3672
rect 3837 3608 3901 3672
rect 3918 3608 3982 3672
rect 3999 3608 4063 3672
rect 4080 3608 4144 3672
rect 4161 3608 4225 3672
rect 4242 3608 4306 3672
rect 4323 3608 4387 3672
rect 4404 3608 4468 3672
rect 4485 3608 4549 3672
rect 4566 3608 4630 3672
rect 4647 3608 4711 3672
rect 4728 3608 4792 3672
rect 4809 3608 4873 3672
rect 105 3520 169 3584
rect 187 3520 251 3584
rect 269 3520 333 3584
rect 351 3520 415 3584
rect 433 3520 497 3584
rect 515 3520 579 3584
rect 597 3520 661 3584
rect 678 3520 742 3584
rect 759 3520 823 3584
rect 840 3520 904 3584
rect 921 3520 985 3584
rect 1002 3520 1066 3584
rect 1083 3520 1147 3584
rect 1164 3520 1228 3584
rect 1245 3520 1309 3584
rect 1326 3520 1390 3584
rect 1407 3520 1471 3584
rect 1488 3520 1552 3584
rect 1569 3520 1633 3584
rect 1650 3520 1714 3584
rect 1731 3520 1795 3584
rect 1812 3520 1876 3584
rect 1893 3520 1957 3584
rect 1974 3520 2038 3584
rect 2055 3520 2119 3584
rect 2136 3520 2200 3584
rect 2217 3520 2281 3584
rect 2298 3520 2362 3584
rect 2379 3520 2443 3584
rect 2460 3520 2524 3584
rect 2541 3520 2605 3584
rect 2622 3520 2686 3584
rect 2703 3520 2767 3584
rect 2784 3520 2848 3584
rect 2865 3520 2929 3584
rect 2946 3520 3010 3584
rect 3027 3520 3091 3584
rect 3108 3520 3172 3584
rect 3189 3520 3253 3584
rect 3270 3520 3334 3584
rect 3351 3520 3415 3584
rect 3432 3520 3496 3584
rect 3513 3520 3577 3584
rect 3594 3520 3658 3584
rect 3675 3520 3739 3584
rect 3756 3520 3820 3584
rect 3837 3520 3901 3584
rect 3918 3520 3982 3584
rect 3999 3520 4063 3584
rect 4080 3520 4144 3584
rect 4161 3520 4225 3584
rect 4242 3520 4306 3584
rect 4323 3520 4387 3584
rect 4404 3520 4468 3584
rect 4485 3520 4549 3584
rect 4566 3520 4630 3584
rect 4647 3520 4711 3584
rect 4728 3520 4792 3584
rect 4809 3520 4873 3584
rect 105 3432 169 3496
rect 187 3432 251 3496
rect 269 3432 333 3496
rect 351 3432 415 3496
rect 433 3432 497 3496
rect 515 3432 579 3496
rect 597 3432 661 3496
rect 678 3432 742 3496
rect 759 3432 823 3496
rect 840 3432 904 3496
rect 921 3432 985 3496
rect 1002 3432 1066 3496
rect 1083 3432 1147 3496
rect 1164 3432 1228 3496
rect 1245 3432 1309 3496
rect 1326 3432 1390 3496
rect 1407 3432 1471 3496
rect 1488 3432 1552 3496
rect 1569 3432 1633 3496
rect 1650 3432 1714 3496
rect 1731 3432 1795 3496
rect 1812 3432 1876 3496
rect 1893 3432 1957 3496
rect 1974 3432 2038 3496
rect 2055 3432 2119 3496
rect 2136 3432 2200 3496
rect 2217 3432 2281 3496
rect 2298 3432 2362 3496
rect 2379 3432 2443 3496
rect 2460 3432 2524 3496
rect 2541 3432 2605 3496
rect 2622 3432 2686 3496
rect 2703 3432 2767 3496
rect 2784 3432 2848 3496
rect 2865 3432 2929 3496
rect 2946 3432 3010 3496
rect 3027 3432 3091 3496
rect 3108 3432 3172 3496
rect 3189 3432 3253 3496
rect 3270 3432 3334 3496
rect 3351 3432 3415 3496
rect 3432 3432 3496 3496
rect 3513 3432 3577 3496
rect 3594 3432 3658 3496
rect 3675 3432 3739 3496
rect 3756 3432 3820 3496
rect 3837 3432 3901 3496
rect 3918 3432 3982 3496
rect 3999 3432 4063 3496
rect 4080 3432 4144 3496
rect 4161 3432 4225 3496
rect 4242 3432 4306 3496
rect 4323 3432 4387 3496
rect 4404 3432 4468 3496
rect 4485 3432 4549 3496
rect 4566 3432 4630 3496
rect 4647 3432 4711 3496
rect 4728 3432 4792 3496
rect 4809 3432 4873 3496
rect 105 3344 169 3408
rect 187 3344 251 3408
rect 269 3344 333 3408
rect 351 3344 415 3408
rect 433 3344 497 3408
rect 515 3344 579 3408
rect 597 3344 661 3408
rect 678 3344 742 3408
rect 759 3344 823 3408
rect 840 3344 904 3408
rect 921 3344 985 3408
rect 1002 3344 1066 3408
rect 1083 3344 1147 3408
rect 1164 3344 1228 3408
rect 1245 3344 1309 3408
rect 1326 3344 1390 3408
rect 1407 3344 1471 3408
rect 1488 3344 1552 3408
rect 1569 3344 1633 3408
rect 1650 3344 1714 3408
rect 1731 3344 1795 3408
rect 1812 3344 1876 3408
rect 1893 3344 1957 3408
rect 1974 3344 2038 3408
rect 2055 3344 2119 3408
rect 2136 3344 2200 3408
rect 2217 3344 2281 3408
rect 2298 3344 2362 3408
rect 2379 3344 2443 3408
rect 2460 3344 2524 3408
rect 2541 3344 2605 3408
rect 2622 3344 2686 3408
rect 2703 3344 2767 3408
rect 2784 3344 2848 3408
rect 2865 3344 2929 3408
rect 2946 3344 3010 3408
rect 3027 3344 3091 3408
rect 3108 3344 3172 3408
rect 3189 3344 3253 3408
rect 3270 3344 3334 3408
rect 3351 3344 3415 3408
rect 3432 3344 3496 3408
rect 3513 3344 3577 3408
rect 3594 3344 3658 3408
rect 3675 3344 3739 3408
rect 3756 3344 3820 3408
rect 3837 3344 3901 3408
rect 3918 3344 3982 3408
rect 3999 3344 4063 3408
rect 4080 3344 4144 3408
rect 4161 3344 4225 3408
rect 4242 3344 4306 3408
rect 4323 3344 4387 3408
rect 4404 3344 4468 3408
rect 4485 3344 4549 3408
rect 4566 3344 4630 3408
rect 4647 3344 4711 3408
rect 4728 3344 4792 3408
rect 4809 3344 4873 3408
rect 105 3256 169 3320
rect 187 3256 251 3320
rect 269 3256 333 3320
rect 351 3256 415 3320
rect 433 3256 497 3320
rect 515 3256 579 3320
rect 597 3256 661 3320
rect 678 3256 742 3320
rect 759 3256 823 3320
rect 840 3256 904 3320
rect 921 3256 985 3320
rect 1002 3256 1066 3320
rect 1083 3256 1147 3320
rect 1164 3256 1228 3320
rect 1245 3256 1309 3320
rect 1326 3256 1390 3320
rect 1407 3256 1471 3320
rect 1488 3256 1552 3320
rect 1569 3256 1633 3320
rect 1650 3256 1714 3320
rect 1731 3256 1795 3320
rect 1812 3256 1876 3320
rect 1893 3256 1957 3320
rect 1974 3256 2038 3320
rect 2055 3256 2119 3320
rect 2136 3256 2200 3320
rect 2217 3256 2281 3320
rect 2298 3256 2362 3320
rect 2379 3256 2443 3320
rect 2460 3256 2524 3320
rect 2541 3256 2605 3320
rect 2622 3256 2686 3320
rect 2703 3256 2767 3320
rect 2784 3256 2848 3320
rect 2865 3256 2929 3320
rect 2946 3256 3010 3320
rect 3027 3256 3091 3320
rect 3108 3256 3172 3320
rect 3189 3256 3253 3320
rect 3270 3256 3334 3320
rect 3351 3256 3415 3320
rect 3432 3256 3496 3320
rect 3513 3256 3577 3320
rect 3594 3256 3658 3320
rect 3675 3256 3739 3320
rect 3756 3256 3820 3320
rect 3837 3256 3901 3320
rect 3918 3256 3982 3320
rect 3999 3256 4063 3320
rect 4080 3256 4144 3320
rect 4161 3256 4225 3320
rect 4242 3256 4306 3320
rect 4323 3256 4387 3320
rect 4404 3256 4468 3320
rect 4485 3256 4549 3320
rect 4566 3256 4630 3320
rect 4647 3256 4711 3320
rect 4728 3256 4792 3320
rect 4809 3256 4873 3320
rect 105 3168 169 3232
rect 187 3168 251 3232
rect 269 3168 333 3232
rect 351 3168 415 3232
rect 433 3168 497 3232
rect 515 3168 579 3232
rect 597 3168 661 3232
rect 678 3168 742 3232
rect 759 3168 823 3232
rect 840 3168 904 3232
rect 921 3168 985 3232
rect 1002 3168 1066 3232
rect 1083 3168 1147 3232
rect 1164 3168 1228 3232
rect 1245 3168 1309 3232
rect 1326 3168 1390 3232
rect 1407 3168 1471 3232
rect 1488 3168 1552 3232
rect 1569 3168 1633 3232
rect 1650 3168 1714 3232
rect 1731 3168 1795 3232
rect 1812 3168 1876 3232
rect 1893 3168 1957 3232
rect 1974 3168 2038 3232
rect 2055 3168 2119 3232
rect 2136 3168 2200 3232
rect 2217 3168 2281 3232
rect 2298 3168 2362 3232
rect 2379 3168 2443 3232
rect 2460 3168 2524 3232
rect 2541 3168 2605 3232
rect 2622 3168 2686 3232
rect 2703 3168 2767 3232
rect 2784 3168 2848 3232
rect 2865 3168 2929 3232
rect 2946 3168 3010 3232
rect 3027 3168 3091 3232
rect 3108 3168 3172 3232
rect 3189 3168 3253 3232
rect 3270 3168 3334 3232
rect 3351 3168 3415 3232
rect 3432 3168 3496 3232
rect 3513 3168 3577 3232
rect 3594 3168 3658 3232
rect 3675 3168 3739 3232
rect 3756 3168 3820 3232
rect 3837 3168 3901 3232
rect 3918 3168 3982 3232
rect 3999 3168 4063 3232
rect 4080 3168 4144 3232
rect 4161 3168 4225 3232
rect 4242 3168 4306 3232
rect 4323 3168 4387 3232
rect 4404 3168 4468 3232
rect 4485 3168 4549 3232
rect 4566 3168 4630 3232
rect 4647 3168 4711 3232
rect 4728 3168 4792 3232
rect 4809 3168 4873 3232
rect 105 3080 169 3144
rect 187 3080 251 3144
rect 269 3080 333 3144
rect 351 3080 415 3144
rect 433 3080 497 3144
rect 515 3080 579 3144
rect 597 3080 661 3144
rect 678 3080 742 3144
rect 759 3080 823 3144
rect 840 3080 904 3144
rect 921 3080 985 3144
rect 1002 3080 1066 3144
rect 1083 3080 1147 3144
rect 1164 3080 1228 3144
rect 1245 3080 1309 3144
rect 1326 3080 1390 3144
rect 1407 3080 1471 3144
rect 1488 3080 1552 3144
rect 1569 3080 1633 3144
rect 1650 3080 1714 3144
rect 1731 3080 1795 3144
rect 1812 3080 1876 3144
rect 1893 3080 1957 3144
rect 1974 3080 2038 3144
rect 2055 3080 2119 3144
rect 2136 3080 2200 3144
rect 2217 3080 2281 3144
rect 2298 3080 2362 3144
rect 2379 3080 2443 3144
rect 2460 3080 2524 3144
rect 2541 3080 2605 3144
rect 2622 3080 2686 3144
rect 2703 3080 2767 3144
rect 2784 3080 2848 3144
rect 2865 3080 2929 3144
rect 2946 3080 3010 3144
rect 3027 3080 3091 3144
rect 3108 3080 3172 3144
rect 3189 3080 3253 3144
rect 3270 3080 3334 3144
rect 3351 3080 3415 3144
rect 3432 3080 3496 3144
rect 3513 3080 3577 3144
rect 3594 3080 3658 3144
rect 3675 3080 3739 3144
rect 3756 3080 3820 3144
rect 3837 3080 3901 3144
rect 3918 3080 3982 3144
rect 3999 3080 4063 3144
rect 4080 3080 4144 3144
rect 4161 3080 4225 3144
rect 4242 3080 4306 3144
rect 4323 3080 4387 3144
rect 4404 3080 4468 3144
rect 4485 3080 4549 3144
rect 4566 3080 4630 3144
rect 4647 3080 4711 3144
rect 4728 3080 4792 3144
rect 4809 3080 4873 3144
rect 105 2992 169 3056
rect 187 2992 251 3056
rect 269 2992 333 3056
rect 351 2992 415 3056
rect 433 2992 497 3056
rect 515 2992 579 3056
rect 597 2992 661 3056
rect 678 2992 742 3056
rect 759 2992 823 3056
rect 840 2992 904 3056
rect 921 2992 985 3056
rect 1002 2992 1066 3056
rect 1083 2992 1147 3056
rect 1164 2992 1228 3056
rect 1245 2992 1309 3056
rect 1326 2992 1390 3056
rect 1407 2992 1471 3056
rect 1488 2992 1552 3056
rect 1569 2992 1633 3056
rect 1650 2992 1714 3056
rect 1731 2992 1795 3056
rect 1812 2992 1876 3056
rect 1893 2992 1957 3056
rect 1974 2992 2038 3056
rect 2055 2992 2119 3056
rect 2136 2992 2200 3056
rect 2217 2992 2281 3056
rect 2298 2992 2362 3056
rect 2379 2992 2443 3056
rect 2460 2992 2524 3056
rect 2541 2992 2605 3056
rect 2622 2992 2686 3056
rect 2703 2992 2767 3056
rect 2784 2992 2848 3056
rect 2865 2992 2929 3056
rect 2946 2992 3010 3056
rect 3027 2992 3091 3056
rect 3108 2992 3172 3056
rect 3189 2992 3253 3056
rect 3270 2992 3334 3056
rect 3351 2992 3415 3056
rect 3432 2992 3496 3056
rect 3513 2992 3577 3056
rect 3594 2992 3658 3056
rect 3675 2992 3739 3056
rect 3756 2992 3820 3056
rect 3837 2992 3901 3056
rect 3918 2992 3982 3056
rect 3999 2992 4063 3056
rect 4080 2992 4144 3056
rect 4161 2992 4225 3056
rect 4242 2992 4306 3056
rect 4323 2992 4387 3056
rect 4404 2992 4468 3056
rect 4485 2992 4549 3056
rect 4566 2992 4630 3056
rect 4647 2992 4711 3056
rect 4728 2992 4792 3056
rect 4809 2992 4873 3056
rect 10084 3608 10148 3672
rect 10166 3608 10230 3672
rect 10248 3608 10312 3672
rect 10330 3608 10394 3672
rect 10412 3608 10476 3672
rect 10494 3608 10558 3672
rect 10576 3608 10640 3672
rect 10657 3608 10721 3672
rect 10738 3608 10802 3672
rect 10819 3608 10883 3672
rect 10900 3608 10964 3672
rect 10981 3608 11045 3672
rect 11062 3608 11126 3672
rect 11143 3608 11207 3672
rect 11224 3608 11288 3672
rect 11305 3608 11369 3672
rect 11386 3608 11450 3672
rect 11467 3608 11531 3672
rect 11548 3608 11612 3672
rect 11629 3608 11693 3672
rect 11710 3608 11774 3672
rect 11791 3608 11855 3672
rect 11872 3608 11936 3672
rect 11953 3608 12017 3672
rect 12034 3608 12098 3672
rect 12115 3608 12179 3672
rect 12196 3608 12260 3672
rect 12277 3608 12341 3672
rect 12358 3608 12422 3672
rect 12439 3608 12503 3672
rect 12520 3608 12584 3672
rect 12601 3608 12665 3672
rect 12682 3608 12746 3672
rect 12763 3608 12827 3672
rect 12844 3608 12908 3672
rect 12925 3608 12989 3672
rect 13006 3608 13070 3672
rect 13087 3608 13151 3672
rect 13168 3608 13232 3672
rect 13249 3608 13313 3672
rect 13330 3608 13394 3672
rect 13411 3608 13475 3672
rect 13492 3608 13556 3672
rect 13573 3608 13637 3672
rect 13654 3608 13718 3672
rect 13735 3608 13799 3672
rect 13816 3608 13880 3672
rect 13897 3608 13961 3672
rect 13978 3608 14042 3672
rect 14059 3608 14123 3672
rect 14140 3608 14204 3672
rect 14221 3608 14285 3672
rect 14302 3608 14366 3672
rect 14383 3608 14447 3672
rect 14464 3608 14528 3672
rect 14545 3608 14609 3672
rect 14626 3608 14690 3672
rect 14707 3608 14771 3672
rect 14788 3608 14852 3672
rect 10084 3520 10148 3584
rect 10166 3520 10230 3584
rect 10248 3520 10312 3584
rect 10330 3520 10394 3584
rect 10412 3520 10476 3584
rect 10494 3520 10558 3584
rect 10576 3520 10640 3584
rect 10657 3520 10721 3584
rect 10738 3520 10802 3584
rect 10819 3520 10883 3584
rect 10900 3520 10964 3584
rect 10981 3520 11045 3584
rect 11062 3520 11126 3584
rect 11143 3520 11207 3584
rect 11224 3520 11288 3584
rect 11305 3520 11369 3584
rect 11386 3520 11450 3584
rect 11467 3520 11531 3584
rect 11548 3520 11612 3584
rect 11629 3520 11693 3584
rect 11710 3520 11774 3584
rect 11791 3520 11855 3584
rect 11872 3520 11936 3584
rect 11953 3520 12017 3584
rect 12034 3520 12098 3584
rect 12115 3520 12179 3584
rect 12196 3520 12260 3584
rect 12277 3520 12341 3584
rect 12358 3520 12422 3584
rect 12439 3520 12503 3584
rect 12520 3520 12584 3584
rect 12601 3520 12665 3584
rect 12682 3520 12746 3584
rect 12763 3520 12827 3584
rect 12844 3520 12908 3584
rect 12925 3520 12989 3584
rect 13006 3520 13070 3584
rect 13087 3520 13151 3584
rect 13168 3520 13232 3584
rect 13249 3520 13313 3584
rect 13330 3520 13394 3584
rect 13411 3520 13475 3584
rect 13492 3520 13556 3584
rect 13573 3520 13637 3584
rect 13654 3520 13718 3584
rect 13735 3520 13799 3584
rect 13816 3520 13880 3584
rect 13897 3520 13961 3584
rect 13978 3520 14042 3584
rect 14059 3520 14123 3584
rect 14140 3520 14204 3584
rect 14221 3520 14285 3584
rect 14302 3520 14366 3584
rect 14383 3520 14447 3584
rect 14464 3520 14528 3584
rect 14545 3520 14609 3584
rect 14626 3520 14690 3584
rect 14707 3520 14771 3584
rect 14788 3520 14852 3584
rect 10084 3432 10148 3496
rect 10166 3432 10230 3496
rect 10248 3432 10312 3496
rect 10330 3432 10394 3496
rect 10412 3432 10476 3496
rect 10494 3432 10558 3496
rect 10576 3432 10640 3496
rect 10657 3432 10721 3496
rect 10738 3432 10802 3496
rect 10819 3432 10883 3496
rect 10900 3432 10964 3496
rect 10981 3432 11045 3496
rect 11062 3432 11126 3496
rect 11143 3432 11207 3496
rect 11224 3432 11288 3496
rect 11305 3432 11369 3496
rect 11386 3432 11450 3496
rect 11467 3432 11531 3496
rect 11548 3432 11612 3496
rect 11629 3432 11693 3496
rect 11710 3432 11774 3496
rect 11791 3432 11855 3496
rect 11872 3432 11936 3496
rect 11953 3432 12017 3496
rect 12034 3432 12098 3496
rect 12115 3432 12179 3496
rect 12196 3432 12260 3496
rect 12277 3432 12341 3496
rect 12358 3432 12422 3496
rect 12439 3432 12503 3496
rect 12520 3432 12584 3496
rect 12601 3432 12665 3496
rect 12682 3432 12746 3496
rect 12763 3432 12827 3496
rect 12844 3432 12908 3496
rect 12925 3432 12989 3496
rect 13006 3432 13070 3496
rect 13087 3432 13151 3496
rect 13168 3432 13232 3496
rect 13249 3432 13313 3496
rect 13330 3432 13394 3496
rect 13411 3432 13475 3496
rect 13492 3432 13556 3496
rect 13573 3432 13637 3496
rect 13654 3432 13718 3496
rect 13735 3432 13799 3496
rect 13816 3432 13880 3496
rect 13897 3432 13961 3496
rect 13978 3432 14042 3496
rect 14059 3432 14123 3496
rect 14140 3432 14204 3496
rect 14221 3432 14285 3496
rect 14302 3432 14366 3496
rect 14383 3432 14447 3496
rect 14464 3432 14528 3496
rect 14545 3432 14609 3496
rect 14626 3432 14690 3496
rect 14707 3432 14771 3496
rect 14788 3432 14852 3496
rect 10084 3344 10148 3408
rect 10166 3344 10230 3408
rect 10248 3344 10312 3408
rect 10330 3344 10394 3408
rect 10412 3344 10476 3408
rect 10494 3344 10558 3408
rect 10576 3344 10640 3408
rect 10657 3344 10721 3408
rect 10738 3344 10802 3408
rect 10819 3344 10883 3408
rect 10900 3344 10964 3408
rect 10981 3344 11045 3408
rect 11062 3344 11126 3408
rect 11143 3344 11207 3408
rect 11224 3344 11288 3408
rect 11305 3344 11369 3408
rect 11386 3344 11450 3408
rect 11467 3344 11531 3408
rect 11548 3344 11612 3408
rect 11629 3344 11693 3408
rect 11710 3344 11774 3408
rect 11791 3344 11855 3408
rect 11872 3344 11936 3408
rect 11953 3344 12017 3408
rect 12034 3344 12098 3408
rect 12115 3344 12179 3408
rect 12196 3344 12260 3408
rect 12277 3344 12341 3408
rect 12358 3344 12422 3408
rect 12439 3344 12503 3408
rect 12520 3344 12584 3408
rect 12601 3344 12665 3408
rect 12682 3344 12746 3408
rect 12763 3344 12827 3408
rect 12844 3344 12908 3408
rect 12925 3344 12989 3408
rect 13006 3344 13070 3408
rect 13087 3344 13151 3408
rect 13168 3344 13232 3408
rect 13249 3344 13313 3408
rect 13330 3344 13394 3408
rect 13411 3344 13475 3408
rect 13492 3344 13556 3408
rect 13573 3344 13637 3408
rect 13654 3344 13718 3408
rect 13735 3344 13799 3408
rect 13816 3344 13880 3408
rect 13897 3344 13961 3408
rect 13978 3344 14042 3408
rect 14059 3344 14123 3408
rect 14140 3344 14204 3408
rect 14221 3344 14285 3408
rect 14302 3344 14366 3408
rect 14383 3344 14447 3408
rect 14464 3344 14528 3408
rect 14545 3344 14609 3408
rect 14626 3344 14690 3408
rect 14707 3344 14771 3408
rect 14788 3344 14852 3408
rect 10084 3256 10148 3320
rect 10166 3256 10230 3320
rect 10248 3256 10312 3320
rect 10330 3256 10394 3320
rect 10412 3256 10476 3320
rect 10494 3256 10558 3320
rect 10576 3256 10640 3320
rect 10657 3256 10721 3320
rect 10738 3256 10802 3320
rect 10819 3256 10883 3320
rect 10900 3256 10964 3320
rect 10981 3256 11045 3320
rect 11062 3256 11126 3320
rect 11143 3256 11207 3320
rect 11224 3256 11288 3320
rect 11305 3256 11369 3320
rect 11386 3256 11450 3320
rect 11467 3256 11531 3320
rect 11548 3256 11612 3320
rect 11629 3256 11693 3320
rect 11710 3256 11774 3320
rect 11791 3256 11855 3320
rect 11872 3256 11936 3320
rect 11953 3256 12017 3320
rect 12034 3256 12098 3320
rect 12115 3256 12179 3320
rect 12196 3256 12260 3320
rect 12277 3256 12341 3320
rect 12358 3256 12422 3320
rect 12439 3256 12503 3320
rect 12520 3256 12584 3320
rect 12601 3256 12665 3320
rect 12682 3256 12746 3320
rect 12763 3256 12827 3320
rect 12844 3256 12908 3320
rect 12925 3256 12989 3320
rect 13006 3256 13070 3320
rect 13087 3256 13151 3320
rect 13168 3256 13232 3320
rect 13249 3256 13313 3320
rect 13330 3256 13394 3320
rect 13411 3256 13475 3320
rect 13492 3256 13556 3320
rect 13573 3256 13637 3320
rect 13654 3256 13718 3320
rect 13735 3256 13799 3320
rect 13816 3256 13880 3320
rect 13897 3256 13961 3320
rect 13978 3256 14042 3320
rect 14059 3256 14123 3320
rect 14140 3256 14204 3320
rect 14221 3256 14285 3320
rect 14302 3256 14366 3320
rect 14383 3256 14447 3320
rect 14464 3256 14528 3320
rect 14545 3256 14609 3320
rect 14626 3256 14690 3320
rect 14707 3256 14771 3320
rect 14788 3256 14852 3320
rect 10084 3168 10148 3232
rect 10166 3168 10230 3232
rect 10248 3168 10312 3232
rect 10330 3168 10394 3232
rect 10412 3168 10476 3232
rect 10494 3168 10558 3232
rect 10576 3168 10640 3232
rect 10657 3168 10721 3232
rect 10738 3168 10802 3232
rect 10819 3168 10883 3232
rect 10900 3168 10964 3232
rect 10981 3168 11045 3232
rect 11062 3168 11126 3232
rect 11143 3168 11207 3232
rect 11224 3168 11288 3232
rect 11305 3168 11369 3232
rect 11386 3168 11450 3232
rect 11467 3168 11531 3232
rect 11548 3168 11612 3232
rect 11629 3168 11693 3232
rect 11710 3168 11774 3232
rect 11791 3168 11855 3232
rect 11872 3168 11936 3232
rect 11953 3168 12017 3232
rect 12034 3168 12098 3232
rect 12115 3168 12179 3232
rect 12196 3168 12260 3232
rect 12277 3168 12341 3232
rect 12358 3168 12422 3232
rect 12439 3168 12503 3232
rect 12520 3168 12584 3232
rect 12601 3168 12665 3232
rect 12682 3168 12746 3232
rect 12763 3168 12827 3232
rect 12844 3168 12908 3232
rect 12925 3168 12989 3232
rect 13006 3168 13070 3232
rect 13087 3168 13151 3232
rect 13168 3168 13232 3232
rect 13249 3168 13313 3232
rect 13330 3168 13394 3232
rect 13411 3168 13475 3232
rect 13492 3168 13556 3232
rect 13573 3168 13637 3232
rect 13654 3168 13718 3232
rect 13735 3168 13799 3232
rect 13816 3168 13880 3232
rect 13897 3168 13961 3232
rect 13978 3168 14042 3232
rect 14059 3168 14123 3232
rect 14140 3168 14204 3232
rect 14221 3168 14285 3232
rect 14302 3168 14366 3232
rect 14383 3168 14447 3232
rect 14464 3168 14528 3232
rect 14545 3168 14609 3232
rect 14626 3168 14690 3232
rect 14707 3168 14771 3232
rect 14788 3168 14852 3232
rect 10084 3080 10148 3144
rect 10166 3080 10230 3144
rect 10248 3080 10312 3144
rect 10330 3080 10394 3144
rect 10412 3080 10476 3144
rect 10494 3080 10558 3144
rect 10576 3080 10640 3144
rect 10657 3080 10721 3144
rect 10738 3080 10802 3144
rect 10819 3080 10883 3144
rect 10900 3080 10964 3144
rect 10981 3080 11045 3144
rect 11062 3080 11126 3144
rect 11143 3080 11207 3144
rect 11224 3080 11288 3144
rect 11305 3080 11369 3144
rect 11386 3080 11450 3144
rect 11467 3080 11531 3144
rect 11548 3080 11612 3144
rect 11629 3080 11693 3144
rect 11710 3080 11774 3144
rect 11791 3080 11855 3144
rect 11872 3080 11936 3144
rect 11953 3080 12017 3144
rect 12034 3080 12098 3144
rect 12115 3080 12179 3144
rect 12196 3080 12260 3144
rect 12277 3080 12341 3144
rect 12358 3080 12422 3144
rect 12439 3080 12503 3144
rect 12520 3080 12584 3144
rect 12601 3080 12665 3144
rect 12682 3080 12746 3144
rect 12763 3080 12827 3144
rect 12844 3080 12908 3144
rect 12925 3080 12989 3144
rect 13006 3080 13070 3144
rect 13087 3080 13151 3144
rect 13168 3080 13232 3144
rect 13249 3080 13313 3144
rect 13330 3080 13394 3144
rect 13411 3080 13475 3144
rect 13492 3080 13556 3144
rect 13573 3080 13637 3144
rect 13654 3080 13718 3144
rect 13735 3080 13799 3144
rect 13816 3080 13880 3144
rect 13897 3080 13961 3144
rect 13978 3080 14042 3144
rect 14059 3080 14123 3144
rect 14140 3080 14204 3144
rect 14221 3080 14285 3144
rect 14302 3080 14366 3144
rect 14383 3080 14447 3144
rect 14464 3080 14528 3144
rect 14545 3080 14609 3144
rect 14626 3080 14690 3144
rect 14707 3080 14771 3144
rect 14788 3080 14852 3144
rect 10084 2992 10148 3056
rect 10166 2992 10230 3056
rect 10248 2992 10312 3056
rect 10330 2992 10394 3056
rect 10412 2992 10476 3056
rect 10494 2992 10558 3056
rect 10576 2992 10640 3056
rect 10657 2992 10721 3056
rect 10738 2992 10802 3056
rect 10819 2992 10883 3056
rect 10900 2992 10964 3056
rect 10981 2992 11045 3056
rect 11062 2992 11126 3056
rect 11143 2992 11207 3056
rect 11224 2992 11288 3056
rect 11305 2992 11369 3056
rect 11386 2992 11450 3056
rect 11467 2992 11531 3056
rect 11548 2992 11612 3056
rect 11629 2992 11693 3056
rect 11710 2992 11774 3056
rect 11791 2992 11855 3056
rect 11872 2992 11936 3056
rect 11953 2992 12017 3056
rect 12034 2992 12098 3056
rect 12115 2992 12179 3056
rect 12196 2992 12260 3056
rect 12277 2992 12341 3056
rect 12358 2992 12422 3056
rect 12439 2992 12503 3056
rect 12520 2992 12584 3056
rect 12601 2992 12665 3056
rect 12682 2992 12746 3056
rect 12763 2992 12827 3056
rect 12844 2992 12908 3056
rect 12925 2992 12989 3056
rect 13006 2992 13070 3056
rect 13087 2992 13151 3056
rect 13168 2992 13232 3056
rect 13249 2992 13313 3056
rect 13330 2992 13394 3056
rect 13411 2992 13475 3056
rect 13492 2992 13556 3056
rect 13573 2992 13637 3056
rect 13654 2992 13718 3056
rect 13735 2992 13799 3056
rect 13816 2992 13880 3056
rect 13897 2992 13961 3056
rect 13978 2992 14042 3056
rect 14059 2992 14123 3056
rect 14140 2992 14204 3056
rect 14221 2992 14285 3056
rect 14302 2992 14366 3056
rect 14383 2992 14447 3056
rect 14464 2992 14528 3056
rect 14545 2992 14609 3056
rect 14626 2992 14690 3056
rect 14707 2992 14771 3056
rect 14788 2992 14852 3056
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 254 11347
rect 14746 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 254 9613
rect 14746 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 3672 4874 3677
rect 0 3608 105 3672
rect 169 3608 187 3672
rect 251 3608 269 3672
rect 333 3608 351 3672
rect 415 3608 433 3672
rect 497 3608 515 3672
rect 579 3608 597 3672
rect 661 3608 678 3672
rect 742 3608 759 3672
rect 823 3608 840 3672
rect 904 3608 921 3672
rect 985 3608 1002 3672
rect 1066 3608 1083 3672
rect 1147 3608 1164 3672
rect 1228 3608 1245 3672
rect 1309 3608 1326 3672
rect 1390 3608 1407 3672
rect 1471 3608 1488 3672
rect 1552 3608 1569 3672
rect 1633 3608 1650 3672
rect 1714 3608 1731 3672
rect 1795 3608 1812 3672
rect 1876 3608 1893 3672
rect 1957 3608 1974 3672
rect 2038 3608 2055 3672
rect 2119 3608 2136 3672
rect 2200 3608 2217 3672
rect 2281 3608 2298 3672
rect 2362 3608 2379 3672
rect 2443 3608 2460 3672
rect 2524 3608 2541 3672
rect 2605 3608 2622 3672
rect 2686 3608 2703 3672
rect 2767 3608 2784 3672
rect 2848 3608 2865 3672
rect 2929 3608 2946 3672
rect 3010 3608 3027 3672
rect 3091 3608 3108 3672
rect 3172 3608 3189 3672
rect 3253 3608 3270 3672
rect 3334 3608 3351 3672
rect 3415 3608 3432 3672
rect 3496 3608 3513 3672
rect 3577 3608 3594 3672
rect 3658 3608 3675 3672
rect 3739 3608 3756 3672
rect 3820 3608 3837 3672
rect 3901 3608 3918 3672
rect 3982 3608 3999 3672
rect 4063 3608 4080 3672
rect 4144 3608 4161 3672
rect 4225 3608 4242 3672
rect 4306 3608 4323 3672
rect 4387 3608 4404 3672
rect 4468 3608 4485 3672
rect 4549 3608 4566 3672
rect 4630 3608 4647 3672
rect 4711 3608 4728 3672
rect 4792 3608 4809 3672
rect 4873 3608 4874 3672
rect 0 3584 4874 3608
rect 0 3520 105 3584
rect 169 3520 187 3584
rect 251 3520 269 3584
rect 333 3520 351 3584
rect 415 3520 433 3584
rect 497 3520 515 3584
rect 579 3520 597 3584
rect 661 3520 678 3584
rect 742 3520 759 3584
rect 823 3520 840 3584
rect 904 3520 921 3584
rect 985 3520 1002 3584
rect 1066 3520 1083 3584
rect 1147 3520 1164 3584
rect 1228 3520 1245 3584
rect 1309 3520 1326 3584
rect 1390 3520 1407 3584
rect 1471 3520 1488 3584
rect 1552 3520 1569 3584
rect 1633 3520 1650 3584
rect 1714 3520 1731 3584
rect 1795 3520 1812 3584
rect 1876 3520 1893 3584
rect 1957 3520 1974 3584
rect 2038 3520 2055 3584
rect 2119 3520 2136 3584
rect 2200 3520 2217 3584
rect 2281 3520 2298 3584
rect 2362 3520 2379 3584
rect 2443 3520 2460 3584
rect 2524 3520 2541 3584
rect 2605 3520 2622 3584
rect 2686 3520 2703 3584
rect 2767 3520 2784 3584
rect 2848 3520 2865 3584
rect 2929 3520 2946 3584
rect 3010 3520 3027 3584
rect 3091 3520 3108 3584
rect 3172 3520 3189 3584
rect 3253 3520 3270 3584
rect 3334 3520 3351 3584
rect 3415 3520 3432 3584
rect 3496 3520 3513 3584
rect 3577 3520 3594 3584
rect 3658 3520 3675 3584
rect 3739 3520 3756 3584
rect 3820 3520 3837 3584
rect 3901 3520 3918 3584
rect 3982 3520 3999 3584
rect 4063 3520 4080 3584
rect 4144 3520 4161 3584
rect 4225 3520 4242 3584
rect 4306 3520 4323 3584
rect 4387 3520 4404 3584
rect 4468 3520 4485 3584
rect 4549 3520 4566 3584
rect 4630 3520 4647 3584
rect 4711 3520 4728 3584
rect 4792 3520 4809 3584
rect 4873 3520 4874 3584
rect 0 3496 4874 3520
rect 0 3432 105 3496
rect 169 3432 187 3496
rect 251 3432 269 3496
rect 333 3432 351 3496
rect 415 3432 433 3496
rect 497 3432 515 3496
rect 579 3432 597 3496
rect 661 3432 678 3496
rect 742 3432 759 3496
rect 823 3432 840 3496
rect 904 3432 921 3496
rect 985 3432 1002 3496
rect 1066 3432 1083 3496
rect 1147 3432 1164 3496
rect 1228 3432 1245 3496
rect 1309 3432 1326 3496
rect 1390 3432 1407 3496
rect 1471 3432 1488 3496
rect 1552 3432 1569 3496
rect 1633 3432 1650 3496
rect 1714 3432 1731 3496
rect 1795 3432 1812 3496
rect 1876 3432 1893 3496
rect 1957 3432 1974 3496
rect 2038 3432 2055 3496
rect 2119 3432 2136 3496
rect 2200 3432 2217 3496
rect 2281 3432 2298 3496
rect 2362 3432 2379 3496
rect 2443 3432 2460 3496
rect 2524 3432 2541 3496
rect 2605 3432 2622 3496
rect 2686 3432 2703 3496
rect 2767 3432 2784 3496
rect 2848 3432 2865 3496
rect 2929 3432 2946 3496
rect 3010 3432 3027 3496
rect 3091 3432 3108 3496
rect 3172 3432 3189 3496
rect 3253 3432 3270 3496
rect 3334 3432 3351 3496
rect 3415 3432 3432 3496
rect 3496 3432 3513 3496
rect 3577 3432 3594 3496
rect 3658 3432 3675 3496
rect 3739 3432 3756 3496
rect 3820 3432 3837 3496
rect 3901 3432 3918 3496
rect 3982 3432 3999 3496
rect 4063 3432 4080 3496
rect 4144 3432 4161 3496
rect 4225 3432 4242 3496
rect 4306 3432 4323 3496
rect 4387 3432 4404 3496
rect 4468 3432 4485 3496
rect 4549 3432 4566 3496
rect 4630 3432 4647 3496
rect 4711 3432 4728 3496
rect 4792 3432 4809 3496
rect 4873 3432 4874 3496
rect 0 3408 4874 3432
rect 0 3344 105 3408
rect 169 3344 187 3408
rect 251 3344 269 3408
rect 333 3344 351 3408
rect 415 3344 433 3408
rect 497 3344 515 3408
rect 579 3344 597 3408
rect 661 3344 678 3408
rect 742 3344 759 3408
rect 823 3344 840 3408
rect 904 3344 921 3408
rect 985 3344 1002 3408
rect 1066 3344 1083 3408
rect 1147 3344 1164 3408
rect 1228 3344 1245 3408
rect 1309 3344 1326 3408
rect 1390 3344 1407 3408
rect 1471 3344 1488 3408
rect 1552 3344 1569 3408
rect 1633 3344 1650 3408
rect 1714 3344 1731 3408
rect 1795 3344 1812 3408
rect 1876 3344 1893 3408
rect 1957 3344 1974 3408
rect 2038 3344 2055 3408
rect 2119 3344 2136 3408
rect 2200 3344 2217 3408
rect 2281 3344 2298 3408
rect 2362 3344 2379 3408
rect 2443 3344 2460 3408
rect 2524 3344 2541 3408
rect 2605 3344 2622 3408
rect 2686 3344 2703 3408
rect 2767 3344 2784 3408
rect 2848 3344 2865 3408
rect 2929 3344 2946 3408
rect 3010 3344 3027 3408
rect 3091 3344 3108 3408
rect 3172 3344 3189 3408
rect 3253 3344 3270 3408
rect 3334 3344 3351 3408
rect 3415 3344 3432 3408
rect 3496 3344 3513 3408
rect 3577 3344 3594 3408
rect 3658 3344 3675 3408
rect 3739 3344 3756 3408
rect 3820 3344 3837 3408
rect 3901 3344 3918 3408
rect 3982 3344 3999 3408
rect 4063 3344 4080 3408
rect 4144 3344 4161 3408
rect 4225 3344 4242 3408
rect 4306 3344 4323 3408
rect 4387 3344 4404 3408
rect 4468 3344 4485 3408
rect 4549 3344 4566 3408
rect 4630 3344 4647 3408
rect 4711 3344 4728 3408
rect 4792 3344 4809 3408
rect 4873 3344 4874 3408
rect 0 3320 4874 3344
rect 0 3256 105 3320
rect 169 3256 187 3320
rect 251 3256 269 3320
rect 333 3256 351 3320
rect 415 3256 433 3320
rect 497 3256 515 3320
rect 579 3256 597 3320
rect 661 3256 678 3320
rect 742 3256 759 3320
rect 823 3256 840 3320
rect 904 3256 921 3320
rect 985 3256 1002 3320
rect 1066 3256 1083 3320
rect 1147 3256 1164 3320
rect 1228 3256 1245 3320
rect 1309 3256 1326 3320
rect 1390 3256 1407 3320
rect 1471 3256 1488 3320
rect 1552 3256 1569 3320
rect 1633 3256 1650 3320
rect 1714 3256 1731 3320
rect 1795 3256 1812 3320
rect 1876 3256 1893 3320
rect 1957 3256 1974 3320
rect 2038 3256 2055 3320
rect 2119 3256 2136 3320
rect 2200 3256 2217 3320
rect 2281 3256 2298 3320
rect 2362 3256 2379 3320
rect 2443 3256 2460 3320
rect 2524 3256 2541 3320
rect 2605 3256 2622 3320
rect 2686 3256 2703 3320
rect 2767 3256 2784 3320
rect 2848 3256 2865 3320
rect 2929 3256 2946 3320
rect 3010 3256 3027 3320
rect 3091 3256 3108 3320
rect 3172 3256 3189 3320
rect 3253 3256 3270 3320
rect 3334 3256 3351 3320
rect 3415 3256 3432 3320
rect 3496 3256 3513 3320
rect 3577 3256 3594 3320
rect 3658 3256 3675 3320
rect 3739 3256 3756 3320
rect 3820 3256 3837 3320
rect 3901 3256 3918 3320
rect 3982 3256 3999 3320
rect 4063 3256 4080 3320
rect 4144 3256 4161 3320
rect 4225 3256 4242 3320
rect 4306 3256 4323 3320
rect 4387 3256 4404 3320
rect 4468 3256 4485 3320
rect 4549 3256 4566 3320
rect 4630 3256 4647 3320
rect 4711 3256 4728 3320
rect 4792 3256 4809 3320
rect 4873 3256 4874 3320
rect 0 3232 4874 3256
rect 0 3168 105 3232
rect 169 3168 187 3232
rect 251 3168 269 3232
rect 333 3168 351 3232
rect 415 3168 433 3232
rect 497 3168 515 3232
rect 579 3168 597 3232
rect 661 3168 678 3232
rect 742 3168 759 3232
rect 823 3168 840 3232
rect 904 3168 921 3232
rect 985 3168 1002 3232
rect 1066 3168 1083 3232
rect 1147 3168 1164 3232
rect 1228 3168 1245 3232
rect 1309 3168 1326 3232
rect 1390 3168 1407 3232
rect 1471 3168 1488 3232
rect 1552 3168 1569 3232
rect 1633 3168 1650 3232
rect 1714 3168 1731 3232
rect 1795 3168 1812 3232
rect 1876 3168 1893 3232
rect 1957 3168 1974 3232
rect 2038 3168 2055 3232
rect 2119 3168 2136 3232
rect 2200 3168 2217 3232
rect 2281 3168 2298 3232
rect 2362 3168 2379 3232
rect 2443 3168 2460 3232
rect 2524 3168 2541 3232
rect 2605 3168 2622 3232
rect 2686 3168 2703 3232
rect 2767 3168 2784 3232
rect 2848 3168 2865 3232
rect 2929 3168 2946 3232
rect 3010 3168 3027 3232
rect 3091 3168 3108 3232
rect 3172 3168 3189 3232
rect 3253 3168 3270 3232
rect 3334 3168 3351 3232
rect 3415 3168 3432 3232
rect 3496 3168 3513 3232
rect 3577 3168 3594 3232
rect 3658 3168 3675 3232
rect 3739 3168 3756 3232
rect 3820 3168 3837 3232
rect 3901 3168 3918 3232
rect 3982 3168 3999 3232
rect 4063 3168 4080 3232
rect 4144 3168 4161 3232
rect 4225 3168 4242 3232
rect 4306 3168 4323 3232
rect 4387 3168 4404 3232
rect 4468 3168 4485 3232
rect 4549 3168 4566 3232
rect 4630 3168 4647 3232
rect 4711 3168 4728 3232
rect 4792 3168 4809 3232
rect 4873 3168 4874 3232
rect 0 3144 4874 3168
rect 0 3080 105 3144
rect 169 3080 187 3144
rect 251 3080 269 3144
rect 333 3080 351 3144
rect 415 3080 433 3144
rect 497 3080 515 3144
rect 579 3080 597 3144
rect 661 3080 678 3144
rect 742 3080 759 3144
rect 823 3080 840 3144
rect 904 3080 921 3144
rect 985 3080 1002 3144
rect 1066 3080 1083 3144
rect 1147 3080 1164 3144
rect 1228 3080 1245 3144
rect 1309 3080 1326 3144
rect 1390 3080 1407 3144
rect 1471 3080 1488 3144
rect 1552 3080 1569 3144
rect 1633 3080 1650 3144
rect 1714 3080 1731 3144
rect 1795 3080 1812 3144
rect 1876 3080 1893 3144
rect 1957 3080 1974 3144
rect 2038 3080 2055 3144
rect 2119 3080 2136 3144
rect 2200 3080 2217 3144
rect 2281 3080 2298 3144
rect 2362 3080 2379 3144
rect 2443 3080 2460 3144
rect 2524 3080 2541 3144
rect 2605 3080 2622 3144
rect 2686 3080 2703 3144
rect 2767 3080 2784 3144
rect 2848 3080 2865 3144
rect 2929 3080 2946 3144
rect 3010 3080 3027 3144
rect 3091 3080 3108 3144
rect 3172 3080 3189 3144
rect 3253 3080 3270 3144
rect 3334 3080 3351 3144
rect 3415 3080 3432 3144
rect 3496 3080 3513 3144
rect 3577 3080 3594 3144
rect 3658 3080 3675 3144
rect 3739 3080 3756 3144
rect 3820 3080 3837 3144
rect 3901 3080 3918 3144
rect 3982 3080 3999 3144
rect 4063 3080 4080 3144
rect 4144 3080 4161 3144
rect 4225 3080 4242 3144
rect 4306 3080 4323 3144
rect 4387 3080 4404 3144
rect 4468 3080 4485 3144
rect 4549 3080 4566 3144
rect 4630 3080 4647 3144
rect 4711 3080 4728 3144
rect 4792 3080 4809 3144
rect 4873 3080 4874 3144
rect 0 3056 4874 3080
rect 0 2992 105 3056
rect 169 2992 187 3056
rect 251 2992 269 3056
rect 333 2992 351 3056
rect 415 2992 433 3056
rect 497 2992 515 3056
rect 579 2992 597 3056
rect 661 2992 678 3056
rect 742 2992 759 3056
rect 823 2992 840 3056
rect 904 2992 921 3056
rect 985 2992 1002 3056
rect 1066 2992 1083 3056
rect 1147 2992 1164 3056
rect 1228 2992 1245 3056
rect 1309 2992 1326 3056
rect 1390 2992 1407 3056
rect 1471 2992 1488 3056
rect 1552 2992 1569 3056
rect 1633 2992 1650 3056
rect 1714 2992 1731 3056
rect 1795 2992 1812 3056
rect 1876 2992 1893 3056
rect 1957 2992 1974 3056
rect 2038 2992 2055 3056
rect 2119 2992 2136 3056
rect 2200 2992 2217 3056
rect 2281 2992 2298 3056
rect 2362 2992 2379 3056
rect 2443 2992 2460 3056
rect 2524 2992 2541 3056
rect 2605 2992 2622 3056
rect 2686 2992 2703 3056
rect 2767 2992 2784 3056
rect 2848 2992 2865 3056
rect 2929 2992 2946 3056
rect 3010 2992 3027 3056
rect 3091 2992 3108 3056
rect 3172 2992 3189 3056
rect 3253 2992 3270 3056
rect 3334 2992 3351 3056
rect 3415 2992 3432 3056
rect 3496 2992 3513 3056
rect 3577 2992 3594 3056
rect 3658 2992 3675 3056
rect 3739 2992 3756 3056
rect 3820 2992 3837 3056
rect 3901 2992 3918 3056
rect 3982 2992 3999 3056
rect 4063 2992 4080 3056
rect 4144 2992 4161 3056
rect 4225 2992 4242 3056
rect 4306 2992 4323 3056
rect 4387 2992 4404 3056
rect 4468 2992 4485 3056
rect 4549 2992 4566 3056
rect 4630 2992 4647 3056
rect 4711 2992 4728 3056
rect 4792 2992 4809 3056
rect 4873 2992 4874 3056
rect 0 2987 4874 2992
rect 10083 3672 15000 3677
rect 10083 3608 10084 3672
rect 10148 3608 10166 3672
rect 10230 3608 10248 3672
rect 10312 3608 10330 3672
rect 10394 3608 10412 3672
rect 10476 3608 10494 3672
rect 10558 3608 10576 3672
rect 10640 3608 10657 3672
rect 10721 3608 10738 3672
rect 10802 3608 10819 3672
rect 10883 3608 10900 3672
rect 10964 3608 10981 3672
rect 11045 3608 11062 3672
rect 11126 3608 11143 3672
rect 11207 3608 11224 3672
rect 11288 3608 11305 3672
rect 11369 3608 11386 3672
rect 11450 3608 11467 3672
rect 11531 3608 11548 3672
rect 11612 3608 11629 3672
rect 11693 3608 11710 3672
rect 11774 3608 11791 3672
rect 11855 3608 11872 3672
rect 11936 3608 11953 3672
rect 12017 3608 12034 3672
rect 12098 3608 12115 3672
rect 12179 3608 12196 3672
rect 12260 3608 12277 3672
rect 12341 3608 12358 3672
rect 12422 3608 12439 3672
rect 12503 3608 12520 3672
rect 12584 3608 12601 3672
rect 12665 3608 12682 3672
rect 12746 3608 12763 3672
rect 12827 3608 12844 3672
rect 12908 3608 12925 3672
rect 12989 3608 13006 3672
rect 13070 3608 13087 3672
rect 13151 3608 13168 3672
rect 13232 3608 13249 3672
rect 13313 3608 13330 3672
rect 13394 3608 13411 3672
rect 13475 3608 13492 3672
rect 13556 3608 13573 3672
rect 13637 3608 13654 3672
rect 13718 3608 13735 3672
rect 13799 3608 13816 3672
rect 13880 3608 13897 3672
rect 13961 3608 13978 3672
rect 14042 3608 14059 3672
rect 14123 3608 14140 3672
rect 14204 3608 14221 3672
rect 14285 3608 14302 3672
rect 14366 3608 14383 3672
rect 14447 3608 14464 3672
rect 14528 3608 14545 3672
rect 14609 3608 14626 3672
rect 14690 3608 14707 3672
rect 14771 3608 14788 3672
rect 14852 3608 15000 3672
rect 10083 3584 15000 3608
rect 10083 3520 10084 3584
rect 10148 3520 10166 3584
rect 10230 3520 10248 3584
rect 10312 3520 10330 3584
rect 10394 3520 10412 3584
rect 10476 3520 10494 3584
rect 10558 3520 10576 3584
rect 10640 3520 10657 3584
rect 10721 3520 10738 3584
rect 10802 3520 10819 3584
rect 10883 3520 10900 3584
rect 10964 3520 10981 3584
rect 11045 3520 11062 3584
rect 11126 3520 11143 3584
rect 11207 3520 11224 3584
rect 11288 3520 11305 3584
rect 11369 3520 11386 3584
rect 11450 3520 11467 3584
rect 11531 3520 11548 3584
rect 11612 3520 11629 3584
rect 11693 3520 11710 3584
rect 11774 3520 11791 3584
rect 11855 3520 11872 3584
rect 11936 3520 11953 3584
rect 12017 3520 12034 3584
rect 12098 3520 12115 3584
rect 12179 3520 12196 3584
rect 12260 3520 12277 3584
rect 12341 3520 12358 3584
rect 12422 3520 12439 3584
rect 12503 3520 12520 3584
rect 12584 3520 12601 3584
rect 12665 3520 12682 3584
rect 12746 3520 12763 3584
rect 12827 3520 12844 3584
rect 12908 3520 12925 3584
rect 12989 3520 13006 3584
rect 13070 3520 13087 3584
rect 13151 3520 13168 3584
rect 13232 3520 13249 3584
rect 13313 3520 13330 3584
rect 13394 3520 13411 3584
rect 13475 3520 13492 3584
rect 13556 3520 13573 3584
rect 13637 3520 13654 3584
rect 13718 3520 13735 3584
rect 13799 3520 13816 3584
rect 13880 3520 13897 3584
rect 13961 3520 13978 3584
rect 14042 3520 14059 3584
rect 14123 3520 14140 3584
rect 14204 3520 14221 3584
rect 14285 3520 14302 3584
rect 14366 3520 14383 3584
rect 14447 3520 14464 3584
rect 14528 3520 14545 3584
rect 14609 3520 14626 3584
rect 14690 3520 14707 3584
rect 14771 3520 14788 3584
rect 14852 3520 15000 3584
rect 10083 3496 15000 3520
rect 10083 3432 10084 3496
rect 10148 3432 10166 3496
rect 10230 3432 10248 3496
rect 10312 3432 10330 3496
rect 10394 3432 10412 3496
rect 10476 3432 10494 3496
rect 10558 3432 10576 3496
rect 10640 3432 10657 3496
rect 10721 3432 10738 3496
rect 10802 3432 10819 3496
rect 10883 3432 10900 3496
rect 10964 3432 10981 3496
rect 11045 3432 11062 3496
rect 11126 3432 11143 3496
rect 11207 3432 11224 3496
rect 11288 3432 11305 3496
rect 11369 3432 11386 3496
rect 11450 3432 11467 3496
rect 11531 3432 11548 3496
rect 11612 3432 11629 3496
rect 11693 3432 11710 3496
rect 11774 3432 11791 3496
rect 11855 3432 11872 3496
rect 11936 3432 11953 3496
rect 12017 3432 12034 3496
rect 12098 3432 12115 3496
rect 12179 3432 12196 3496
rect 12260 3432 12277 3496
rect 12341 3432 12358 3496
rect 12422 3432 12439 3496
rect 12503 3432 12520 3496
rect 12584 3432 12601 3496
rect 12665 3432 12682 3496
rect 12746 3432 12763 3496
rect 12827 3432 12844 3496
rect 12908 3432 12925 3496
rect 12989 3432 13006 3496
rect 13070 3432 13087 3496
rect 13151 3432 13168 3496
rect 13232 3432 13249 3496
rect 13313 3432 13330 3496
rect 13394 3432 13411 3496
rect 13475 3432 13492 3496
rect 13556 3432 13573 3496
rect 13637 3432 13654 3496
rect 13718 3432 13735 3496
rect 13799 3432 13816 3496
rect 13880 3432 13897 3496
rect 13961 3432 13978 3496
rect 14042 3432 14059 3496
rect 14123 3432 14140 3496
rect 14204 3432 14221 3496
rect 14285 3432 14302 3496
rect 14366 3432 14383 3496
rect 14447 3432 14464 3496
rect 14528 3432 14545 3496
rect 14609 3432 14626 3496
rect 14690 3432 14707 3496
rect 14771 3432 14788 3496
rect 14852 3432 15000 3496
rect 10083 3408 15000 3432
rect 10083 3344 10084 3408
rect 10148 3344 10166 3408
rect 10230 3344 10248 3408
rect 10312 3344 10330 3408
rect 10394 3344 10412 3408
rect 10476 3344 10494 3408
rect 10558 3344 10576 3408
rect 10640 3344 10657 3408
rect 10721 3344 10738 3408
rect 10802 3344 10819 3408
rect 10883 3344 10900 3408
rect 10964 3344 10981 3408
rect 11045 3344 11062 3408
rect 11126 3344 11143 3408
rect 11207 3344 11224 3408
rect 11288 3344 11305 3408
rect 11369 3344 11386 3408
rect 11450 3344 11467 3408
rect 11531 3344 11548 3408
rect 11612 3344 11629 3408
rect 11693 3344 11710 3408
rect 11774 3344 11791 3408
rect 11855 3344 11872 3408
rect 11936 3344 11953 3408
rect 12017 3344 12034 3408
rect 12098 3344 12115 3408
rect 12179 3344 12196 3408
rect 12260 3344 12277 3408
rect 12341 3344 12358 3408
rect 12422 3344 12439 3408
rect 12503 3344 12520 3408
rect 12584 3344 12601 3408
rect 12665 3344 12682 3408
rect 12746 3344 12763 3408
rect 12827 3344 12844 3408
rect 12908 3344 12925 3408
rect 12989 3344 13006 3408
rect 13070 3344 13087 3408
rect 13151 3344 13168 3408
rect 13232 3344 13249 3408
rect 13313 3344 13330 3408
rect 13394 3344 13411 3408
rect 13475 3344 13492 3408
rect 13556 3344 13573 3408
rect 13637 3344 13654 3408
rect 13718 3344 13735 3408
rect 13799 3344 13816 3408
rect 13880 3344 13897 3408
rect 13961 3344 13978 3408
rect 14042 3344 14059 3408
rect 14123 3344 14140 3408
rect 14204 3344 14221 3408
rect 14285 3344 14302 3408
rect 14366 3344 14383 3408
rect 14447 3344 14464 3408
rect 14528 3344 14545 3408
rect 14609 3344 14626 3408
rect 14690 3344 14707 3408
rect 14771 3344 14788 3408
rect 14852 3344 15000 3408
rect 10083 3320 15000 3344
rect 10083 3256 10084 3320
rect 10148 3256 10166 3320
rect 10230 3256 10248 3320
rect 10312 3256 10330 3320
rect 10394 3256 10412 3320
rect 10476 3256 10494 3320
rect 10558 3256 10576 3320
rect 10640 3256 10657 3320
rect 10721 3256 10738 3320
rect 10802 3256 10819 3320
rect 10883 3256 10900 3320
rect 10964 3256 10981 3320
rect 11045 3256 11062 3320
rect 11126 3256 11143 3320
rect 11207 3256 11224 3320
rect 11288 3256 11305 3320
rect 11369 3256 11386 3320
rect 11450 3256 11467 3320
rect 11531 3256 11548 3320
rect 11612 3256 11629 3320
rect 11693 3256 11710 3320
rect 11774 3256 11791 3320
rect 11855 3256 11872 3320
rect 11936 3256 11953 3320
rect 12017 3256 12034 3320
rect 12098 3256 12115 3320
rect 12179 3256 12196 3320
rect 12260 3256 12277 3320
rect 12341 3256 12358 3320
rect 12422 3256 12439 3320
rect 12503 3256 12520 3320
rect 12584 3256 12601 3320
rect 12665 3256 12682 3320
rect 12746 3256 12763 3320
rect 12827 3256 12844 3320
rect 12908 3256 12925 3320
rect 12989 3256 13006 3320
rect 13070 3256 13087 3320
rect 13151 3256 13168 3320
rect 13232 3256 13249 3320
rect 13313 3256 13330 3320
rect 13394 3256 13411 3320
rect 13475 3256 13492 3320
rect 13556 3256 13573 3320
rect 13637 3256 13654 3320
rect 13718 3256 13735 3320
rect 13799 3256 13816 3320
rect 13880 3256 13897 3320
rect 13961 3256 13978 3320
rect 14042 3256 14059 3320
rect 14123 3256 14140 3320
rect 14204 3256 14221 3320
rect 14285 3256 14302 3320
rect 14366 3256 14383 3320
rect 14447 3256 14464 3320
rect 14528 3256 14545 3320
rect 14609 3256 14626 3320
rect 14690 3256 14707 3320
rect 14771 3256 14788 3320
rect 14852 3256 15000 3320
rect 10083 3232 15000 3256
rect 10083 3168 10084 3232
rect 10148 3168 10166 3232
rect 10230 3168 10248 3232
rect 10312 3168 10330 3232
rect 10394 3168 10412 3232
rect 10476 3168 10494 3232
rect 10558 3168 10576 3232
rect 10640 3168 10657 3232
rect 10721 3168 10738 3232
rect 10802 3168 10819 3232
rect 10883 3168 10900 3232
rect 10964 3168 10981 3232
rect 11045 3168 11062 3232
rect 11126 3168 11143 3232
rect 11207 3168 11224 3232
rect 11288 3168 11305 3232
rect 11369 3168 11386 3232
rect 11450 3168 11467 3232
rect 11531 3168 11548 3232
rect 11612 3168 11629 3232
rect 11693 3168 11710 3232
rect 11774 3168 11791 3232
rect 11855 3168 11872 3232
rect 11936 3168 11953 3232
rect 12017 3168 12034 3232
rect 12098 3168 12115 3232
rect 12179 3168 12196 3232
rect 12260 3168 12277 3232
rect 12341 3168 12358 3232
rect 12422 3168 12439 3232
rect 12503 3168 12520 3232
rect 12584 3168 12601 3232
rect 12665 3168 12682 3232
rect 12746 3168 12763 3232
rect 12827 3168 12844 3232
rect 12908 3168 12925 3232
rect 12989 3168 13006 3232
rect 13070 3168 13087 3232
rect 13151 3168 13168 3232
rect 13232 3168 13249 3232
rect 13313 3168 13330 3232
rect 13394 3168 13411 3232
rect 13475 3168 13492 3232
rect 13556 3168 13573 3232
rect 13637 3168 13654 3232
rect 13718 3168 13735 3232
rect 13799 3168 13816 3232
rect 13880 3168 13897 3232
rect 13961 3168 13978 3232
rect 14042 3168 14059 3232
rect 14123 3168 14140 3232
rect 14204 3168 14221 3232
rect 14285 3168 14302 3232
rect 14366 3168 14383 3232
rect 14447 3168 14464 3232
rect 14528 3168 14545 3232
rect 14609 3168 14626 3232
rect 14690 3168 14707 3232
rect 14771 3168 14788 3232
rect 14852 3168 15000 3232
rect 10083 3144 15000 3168
rect 10083 3080 10084 3144
rect 10148 3080 10166 3144
rect 10230 3080 10248 3144
rect 10312 3080 10330 3144
rect 10394 3080 10412 3144
rect 10476 3080 10494 3144
rect 10558 3080 10576 3144
rect 10640 3080 10657 3144
rect 10721 3080 10738 3144
rect 10802 3080 10819 3144
rect 10883 3080 10900 3144
rect 10964 3080 10981 3144
rect 11045 3080 11062 3144
rect 11126 3080 11143 3144
rect 11207 3080 11224 3144
rect 11288 3080 11305 3144
rect 11369 3080 11386 3144
rect 11450 3080 11467 3144
rect 11531 3080 11548 3144
rect 11612 3080 11629 3144
rect 11693 3080 11710 3144
rect 11774 3080 11791 3144
rect 11855 3080 11872 3144
rect 11936 3080 11953 3144
rect 12017 3080 12034 3144
rect 12098 3080 12115 3144
rect 12179 3080 12196 3144
rect 12260 3080 12277 3144
rect 12341 3080 12358 3144
rect 12422 3080 12439 3144
rect 12503 3080 12520 3144
rect 12584 3080 12601 3144
rect 12665 3080 12682 3144
rect 12746 3080 12763 3144
rect 12827 3080 12844 3144
rect 12908 3080 12925 3144
rect 12989 3080 13006 3144
rect 13070 3080 13087 3144
rect 13151 3080 13168 3144
rect 13232 3080 13249 3144
rect 13313 3080 13330 3144
rect 13394 3080 13411 3144
rect 13475 3080 13492 3144
rect 13556 3080 13573 3144
rect 13637 3080 13654 3144
rect 13718 3080 13735 3144
rect 13799 3080 13816 3144
rect 13880 3080 13897 3144
rect 13961 3080 13978 3144
rect 14042 3080 14059 3144
rect 14123 3080 14140 3144
rect 14204 3080 14221 3144
rect 14285 3080 14302 3144
rect 14366 3080 14383 3144
rect 14447 3080 14464 3144
rect 14528 3080 14545 3144
rect 14609 3080 14626 3144
rect 14690 3080 14707 3144
rect 14771 3080 14788 3144
rect 14852 3080 15000 3144
rect 10083 3056 15000 3080
rect 10083 2992 10084 3056
rect 10148 2992 10166 3056
rect 10230 2992 10248 3056
rect 10312 2992 10330 3056
rect 10394 2992 10412 3056
rect 10476 2992 10494 3056
rect 10558 2992 10576 3056
rect 10640 2992 10657 3056
rect 10721 2992 10738 3056
rect 10802 2992 10819 3056
rect 10883 2992 10900 3056
rect 10964 2992 10981 3056
rect 11045 2992 11062 3056
rect 11126 2992 11143 3056
rect 11207 2992 11224 3056
rect 11288 2992 11305 3056
rect 11369 2992 11386 3056
rect 11450 2992 11467 3056
rect 11531 2992 11548 3056
rect 11612 2992 11629 3056
rect 11693 2992 11710 3056
rect 11774 2992 11791 3056
rect 11855 2992 11872 3056
rect 11936 2992 11953 3056
rect 12017 2992 12034 3056
rect 12098 2992 12115 3056
rect 12179 2992 12196 3056
rect 12260 2992 12277 3056
rect 12341 2992 12358 3056
rect 12422 2992 12439 3056
rect 12503 2992 12520 3056
rect 12584 2992 12601 3056
rect 12665 2992 12682 3056
rect 12746 2992 12763 3056
rect 12827 2992 12844 3056
rect 12908 2992 12925 3056
rect 12989 2992 13006 3056
rect 13070 2992 13087 3056
rect 13151 2992 13168 3056
rect 13232 2992 13249 3056
rect 13313 2992 13330 3056
rect 13394 2992 13411 3056
rect 13475 2992 13492 3056
rect 13556 2992 13573 3056
rect 13637 2992 13654 3056
rect 13718 2992 13735 3056
rect 13799 2992 13816 3056
rect 13880 2992 13897 3056
rect 13961 2992 13978 3056
rect 14042 2992 14059 3056
rect 14123 2992 14140 3056
rect 14204 2992 14221 3056
rect 14285 2992 14302 3056
rect 14366 2992 14383 3056
rect 14447 2992 14464 3056
rect 14528 2992 14545 3056
rect 14609 2992 14626 3056
rect 14690 2992 14707 3056
rect 14771 2992 14788 3056
rect 14852 2992 15000 3056
rect 10083 2987 15000 2992
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1701704242
transform 1 0 0 0 1 549
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 6 nsew power bidirectional
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 4 nsew power bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 3 nsew ground bidirectional
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 3 nsew ground bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 4 nsew power bidirectional
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 6 nsew power bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 10 nsew power bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 10 nsew power bidirectional
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 3 nsew ground bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 4 nsew power bidirectional
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 3 nsew ground bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 6 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 6 nsew power bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 2 nsew ground bidirectional
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 7 nsew power bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 10 nsew power bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 10 nsew power bidirectional
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 14746 10625 15000 11221 1 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 1 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 1777 15000 2707 1 VCCD
port 6 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 1 VCCD
port 6 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 1 VCCD
port 6 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 1 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 1 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 1 VCCHIB
port 7 nsew power bidirectional
rlabel metal3 s 10078 2988 14858 3676 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2987 4874 3677 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 10083 2987 15000 3677 1 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 1 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3620 14840 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3532 14840 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3444 14840 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3356 14840 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3268 14840 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3180 14840 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3092 14840 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14800 3004 14840 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3620 14759 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3532 14759 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3444 14759 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3356 14759 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3268 14759 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3180 14759 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3092 14759 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14719 3004 14759 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3620 14678 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3532 14678 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3444 14678 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3356 14678 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3268 14678 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3180 14678 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3092 14678 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14638 3004 14678 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3620 14597 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3532 14597 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3444 14597 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3356 14597 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3268 14597 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3180 14597 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3092 14597 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14557 3004 14597 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3620 14516 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3532 14516 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3444 14516 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3356 14516 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3268 14516 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3180 14516 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3092 14516 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14476 3004 14516 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3620 14435 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3532 14435 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3444 14435 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3356 14435 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3268 14435 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3180 14435 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3092 14435 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14395 3004 14435 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3620 14354 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3532 14354 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3444 14354 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3356 14354 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3268 14354 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3180 14354 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3092 14354 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14314 3004 14354 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3620 14273 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3532 14273 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3444 14273 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3356 14273 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3268 14273 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3180 14273 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3092 14273 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14233 3004 14273 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3620 14192 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3532 14192 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3444 14192 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3356 14192 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3268 14192 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3180 14192 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3092 14192 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14152 3004 14192 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3620 14111 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3532 14111 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3444 14111 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3356 14111 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3268 14111 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3180 14111 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3092 14111 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14071 3004 14111 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3620 14030 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3532 14030 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3444 14030 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3356 14030 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3268 14030 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3180 14030 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3092 14030 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13990 3004 14030 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3620 13949 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3532 13949 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3444 13949 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3356 13949 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3268 13949 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3180 13949 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3092 13949 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13909 3004 13949 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3620 13868 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3532 13868 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3444 13868 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3356 13868 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3268 13868 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3180 13868 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3092 13868 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13828 3004 13868 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3620 13787 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3532 13787 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3444 13787 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3356 13787 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3268 13787 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3180 13787 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3092 13787 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13747 3004 13787 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3620 13706 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3532 13706 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3444 13706 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3356 13706 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3268 13706 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3180 13706 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3092 13706 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13666 3004 13706 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3620 13625 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3532 13625 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3444 13625 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3356 13625 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3268 13625 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3180 13625 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3092 13625 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13585 3004 13625 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3620 13544 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3532 13544 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3444 13544 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3356 13544 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3268 13544 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3180 13544 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3092 13544 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13504 3004 13544 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3620 13463 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3532 13463 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3444 13463 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3356 13463 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3268 13463 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3180 13463 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3092 13463 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13423 3004 13463 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3620 13382 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3532 13382 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3444 13382 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3356 13382 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3268 13382 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3180 13382 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3092 13382 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13342 3004 13382 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3620 13301 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3532 13301 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3444 13301 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3356 13301 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3268 13301 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3180 13301 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3092 13301 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13261 3004 13301 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3620 13220 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3532 13220 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3444 13220 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3356 13220 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3268 13220 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3180 13220 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3092 13220 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13180 3004 13220 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3620 13139 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3532 13139 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3444 13139 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3356 13139 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3268 13139 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3180 13139 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3092 13139 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13099 3004 13139 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3620 13058 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3532 13058 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3444 13058 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3356 13058 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3268 13058 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3180 13058 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3092 13058 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13018 3004 13058 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3620 12977 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3532 12977 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3444 12977 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3356 12977 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3268 12977 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3180 12977 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3092 12977 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12937 3004 12977 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3620 12896 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3532 12896 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3444 12896 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3356 12896 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3268 12896 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3180 12896 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3092 12896 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12856 3004 12896 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3620 12815 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3532 12815 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3444 12815 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3356 12815 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3268 12815 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3180 12815 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3092 12815 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12775 3004 12815 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3620 12734 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3532 12734 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3444 12734 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3356 12734 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3268 12734 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3180 12734 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3092 12734 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12694 3004 12734 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3620 12653 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3532 12653 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3444 12653 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3356 12653 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3268 12653 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3180 12653 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3092 12653 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12613 3004 12653 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3620 12572 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3532 12572 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3444 12572 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3356 12572 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3268 12572 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3180 12572 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3092 12572 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12532 3004 12572 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3620 12491 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3532 12491 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3444 12491 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3356 12491 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3268 12491 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3180 12491 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3092 12491 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12451 3004 12491 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3620 12410 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3532 12410 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3444 12410 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3356 12410 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3268 12410 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3180 12410 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3092 12410 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12370 3004 12410 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3620 12329 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3532 12329 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3444 12329 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3356 12329 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3268 12329 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3180 12329 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3092 12329 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12289 3004 12329 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3620 12248 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3532 12248 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3444 12248 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3356 12248 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3268 12248 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3180 12248 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3092 12248 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12208 3004 12248 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3620 12167 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3532 12167 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3444 12167 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3356 12167 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3268 12167 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3180 12167 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3092 12167 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12127 3004 12167 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3620 12086 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3532 12086 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3444 12086 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3356 12086 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3268 12086 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3180 12086 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3092 12086 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12046 3004 12086 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3620 12005 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3532 12005 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3444 12005 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3356 12005 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3268 12005 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3180 12005 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3092 12005 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11965 3004 12005 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3620 11924 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3532 11924 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3444 11924 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3356 11924 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3268 11924 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3180 11924 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3092 11924 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11884 3004 11924 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3620 11843 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3532 11843 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3444 11843 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3356 11843 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3268 11843 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3180 11843 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3092 11843 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11803 3004 11843 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3620 11762 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3532 11762 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3444 11762 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3356 11762 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3268 11762 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3180 11762 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3092 11762 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11722 3004 11762 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3620 11681 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3532 11681 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3444 11681 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3356 11681 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3268 11681 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3180 11681 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3092 11681 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11641 3004 11681 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3620 11600 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3532 11600 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3444 11600 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3356 11600 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3268 11600 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3180 11600 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3092 11600 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11560 3004 11600 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3620 11519 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3532 11519 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3444 11519 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3356 11519 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3268 11519 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3180 11519 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3092 11519 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11479 3004 11519 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3620 11438 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3532 11438 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3444 11438 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3356 11438 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3268 11438 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3180 11438 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3092 11438 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11398 3004 11438 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3620 11357 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3532 11357 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3444 11357 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3356 11357 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3268 11357 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3180 11357 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3092 11357 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11317 3004 11357 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3620 11276 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3532 11276 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3444 11276 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3356 11276 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3268 11276 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3180 11276 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3092 11276 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11236 3004 11276 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3620 11195 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3532 11195 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3444 11195 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3356 11195 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3268 11195 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3180 11195 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3092 11195 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11155 3004 11195 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3620 11114 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3532 11114 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3444 11114 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3356 11114 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3268 11114 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3180 11114 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3092 11114 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11074 3004 11114 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3620 11033 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3532 11033 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3444 11033 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3356 11033 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3268 11033 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3180 11033 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3092 11033 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10993 3004 11033 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3620 10952 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3532 10952 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3444 10952 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3356 10952 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3268 10952 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3180 10952 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3092 10952 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10912 3004 10952 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3620 10871 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3532 10871 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3444 10871 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3356 10871 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3268 10871 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3180 10871 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3092 10871 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10831 3004 10871 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3620 10790 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3532 10790 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3444 10790 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3356 10790 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3268 10790 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3180 10790 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3092 10790 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10750 3004 10790 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3620 10709 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3532 10709 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3444 10709 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3356 10709 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3268 10709 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3180 10709 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3092 10709 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10669 3004 10709 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3620 10628 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3532 10628 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3444 10628 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3356 10628 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3268 10628 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3180 10628 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3092 10628 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10588 3004 10628 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3620 10546 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3532 10546 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3444 10546 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3356 10546 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3268 10546 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3180 10546 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3092 10546 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10506 3004 10546 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3620 10464 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3532 10464 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3444 10464 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3356 10464 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3268 10464 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3180 10464 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3092 10464 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10424 3004 10464 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3620 10382 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3532 10382 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3444 10382 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3356 10382 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3268 10382 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3180 10382 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3092 10382 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10342 3004 10382 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3620 10300 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3532 10300 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3444 10300 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3356 10300 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3268 10300 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3180 10300 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3092 10300 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10260 3004 10300 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3620 10218 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3532 10218 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3444 10218 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3356 10218 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3268 10218 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3180 10218 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3092 10218 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10178 3004 10218 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3620 10136 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3532 10136 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3444 10136 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3356 10136 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3268 10136 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3180 10136 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3092 10136 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10096 3004 10136 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3620 4861 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3532 4861 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3444 4861 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3356 4861 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3268 4861 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3180 4861 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3092 4861 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4821 3004 4861 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3620 4780 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3532 4780 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3444 4780 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3356 4780 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3268 4780 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3180 4780 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3092 4780 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4740 3004 4780 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3620 4699 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3532 4699 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3444 4699 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3356 4699 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3268 4699 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3180 4699 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3092 4699 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4659 3004 4699 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3620 4618 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3532 4618 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3444 4618 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3356 4618 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3268 4618 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3180 4618 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3092 4618 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4578 3004 4618 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3620 4537 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3532 4537 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3444 4537 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3356 4537 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3268 4537 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3180 4537 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3092 4537 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4497 3004 4537 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3620 4456 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3532 4456 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3444 4456 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3356 4456 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3268 4456 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3180 4456 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3092 4456 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4416 3004 4456 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3620 4375 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3532 4375 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3444 4375 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3356 4375 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3268 4375 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3180 4375 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3092 4375 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4335 3004 4375 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3620 4294 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3532 4294 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3444 4294 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3356 4294 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3268 4294 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3180 4294 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3092 4294 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4254 3004 4294 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3620 4213 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3532 4213 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3444 4213 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3356 4213 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3268 4213 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3180 4213 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3092 4213 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4173 3004 4213 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3620 4132 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3532 4132 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3444 4132 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3356 4132 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3268 4132 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3180 4132 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3092 4132 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4092 3004 4132 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3620 4051 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3532 4051 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3444 4051 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3356 4051 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3268 4051 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3180 4051 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3092 4051 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4011 3004 4051 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3620 3970 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3532 3970 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3444 3970 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3356 3970 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3268 3970 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3180 3970 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3092 3970 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3930 3004 3970 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3620 3889 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3532 3889 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3444 3889 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3356 3889 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3268 3889 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3180 3889 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3092 3889 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3849 3004 3889 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3620 3808 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3532 3808 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3444 3808 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3356 3808 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3268 3808 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3180 3808 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3092 3808 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3768 3004 3808 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3620 3727 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3532 3727 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3444 3727 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3356 3727 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3268 3727 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3180 3727 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3092 3727 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3687 3004 3727 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3620 3646 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3532 3646 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3444 3646 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3356 3646 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3268 3646 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3180 3646 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3092 3646 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3606 3004 3646 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3620 3565 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3532 3565 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3444 3565 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3356 3565 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3268 3565 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3180 3565 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3092 3565 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3525 3004 3565 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3620 3484 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3532 3484 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3444 3484 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3356 3484 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3268 3484 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3180 3484 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3092 3484 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3444 3004 3484 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3620 3403 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3532 3403 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3444 3403 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3356 3403 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3268 3403 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3180 3403 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3092 3403 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3363 3004 3403 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3620 3322 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3532 3322 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3444 3322 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3356 3322 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3268 3322 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3180 3322 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3092 3322 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3282 3004 3322 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3620 3241 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3532 3241 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3444 3241 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3356 3241 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3268 3241 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3180 3241 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3092 3241 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3201 3004 3241 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3620 3160 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3532 3160 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3444 3160 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3356 3160 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3268 3160 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3180 3160 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3092 3160 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3120 3004 3160 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3620 3079 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3532 3079 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3444 3079 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3356 3079 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3268 3079 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3180 3079 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3092 3079 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3039 3004 3079 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3620 2998 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3532 2998 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3444 2998 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3356 2998 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3268 2998 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3180 2998 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3092 2998 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2958 3004 2998 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3620 2917 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3532 2917 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3444 2917 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3356 2917 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3268 2917 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3180 2917 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3092 2917 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2877 3004 2917 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3620 2836 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3532 2836 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3444 2836 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3356 2836 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3268 2836 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3180 2836 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3092 2836 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2796 3004 2836 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3620 2755 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3532 2755 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3444 2755 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3356 2755 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3268 2755 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3180 2755 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3092 2755 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2715 3004 2755 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3620 2674 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3532 2674 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3444 2674 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3356 2674 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3268 2674 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3180 2674 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3092 2674 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2634 3004 2674 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3620 2593 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3532 2593 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3444 2593 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3356 2593 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3268 2593 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3180 2593 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3092 2593 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2553 3004 2593 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3620 2512 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3532 2512 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3444 2512 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3356 2512 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3268 2512 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3180 2512 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3092 2512 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2472 3004 2512 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3620 2431 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3532 2431 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3444 2431 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3356 2431 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3268 2431 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3180 2431 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3092 2431 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2391 3004 2431 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3620 2350 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3532 2350 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3444 2350 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3356 2350 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3268 2350 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3180 2350 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3092 2350 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2310 3004 2350 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3620 2269 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3532 2269 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3444 2269 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3356 2269 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3268 2269 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3180 2269 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3092 2269 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2229 3004 2269 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3620 2188 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3532 2188 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3444 2188 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3356 2188 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3268 2188 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3180 2188 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3092 2188 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2148 3004 2188 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3620 2107 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3532 2107 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3444 2107 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3356 2107 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3268 2107 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3180 2107 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3092 2107 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2067 3004 2107 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3620 2026 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3532 2026 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3444 2026 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3356 2026 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3268 2026 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3180 2026 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3092 2026 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1986 3004 2026 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3620 1945 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3532 1945 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3444 1945 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3356 1945 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3268 1945 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3180 1945 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3092 1945 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1905 3004 1945 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3620 1864 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3532 1864 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3444 1864 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3356 1864 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3268 1864 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3180 1864 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3092 1864 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1824 3004 1864 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3620 1783 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3532 1783 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3444 1783 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3356 1783 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3268 1783 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3180 1783 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3092 1783 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1743 3004 1783 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3620 1702 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3532 1702 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3444 1702 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3356 1702 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3268 1702 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3180 1702 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3092 1702 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1662 3004 1702 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3620 1621 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3532 1621 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3444 1621 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3356 1621 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3268 1621 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3180 1621 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3092 1621 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1581 3004 1621 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3620 1540 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3532 1540 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3444 1540 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3356 1540 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3268 1540 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3180 1540 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3092 1540 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1500 3004 1540 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3620 1459 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3532 1459 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3444 1459 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3356 1459 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3268 1459 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3180 1459 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3092 1459 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1419 3004 1459 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3620 1378 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3532 1378 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3444 1378 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3356 1378 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3268 1378 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3180 1378 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3092 1378 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1338 3004 1378 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3620 1297 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3532 1297 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3444 1297 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3356 1297 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3268 1297 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3180 1297 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3092 1297 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1257 3004 1297 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3620 1216 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3532 1216 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3444 1216 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3356 1216 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3268 1216 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3180 1216 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3092 1216 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1176 3004 1216 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3620 1135 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3532 1135 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3444 1135 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3356 1135 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3268 1135 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3180 1135 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3092 1135 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1095 3004 1135 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3620 1054 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3532 1054 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3444 1054 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3356 1054 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3268 1054 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3180 1054 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3092 1054 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1014 3004 1054 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3620 973 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3532 973 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3444 973 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3356 973 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3268 973 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3180 973 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3092 973 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 933 3004 973 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3620 892 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3532 892 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3444 892 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3356 892 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3268 892 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3180 892 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3092 892 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 852 3004 892 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3620 811 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3532 811 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3444 811 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3356 811 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3268 811 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3180 811 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3092 811 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 771 3004 811 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3620 730 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3532 730 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3444 730 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3356 730 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3268 730 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3180 730 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3092 730 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 690 3004 730 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3620 649 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3532 649 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3444 649 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3356 649 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3268 649 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3180 649 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3092 649 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 609 3004 649 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3620 567 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3532 567 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3444 567 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3356 567 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3268 567 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3180 567 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3092 567 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 527 3004 567 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3620 485 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3532 485 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3444 485 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3356 485 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3268 485 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3180 485 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3092 485 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 445 3004 485 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3620 403 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3532 403 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3444 403 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3356 403 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3268 403 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3180 403 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3092 403 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 363 3004 403 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3620 321 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3532 321 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3444 321 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3356 321 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3268 321 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3180 321 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3092 321 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 281 3004 321 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3620 239 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3532 239 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3444 239 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3356 239 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3268 239 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3180 239 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3092 239 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 199 3004 239 3044 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3620 157 3660 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3532 157 3572 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3444 157 3484 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3356 157 3396 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3268 157 3308 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3180 157 3220 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3092 157 3132 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 117 3004 157 3044 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 1 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 1 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 1 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 1 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 1 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 1 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 0 9547 254 9613 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 1 VSSD
port 3 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 1 VSSD
port 3 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 1 VSSD
port 3 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 1 VSSIO_Q
port 2 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 1 VSSIO_Q
port 2 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 1 VSSIO_Q
port 2 nsew ground bidirectional
rlabel metal4 s 14746 6377 15000 7067 1 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 1 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 1 VSWITCH
port 8 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string GDS_END 10273786
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 10204906
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
