magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 687 2066
<< mvpmos >>
rect 0 0 100 2000
rect 156 0 256 2000
rect 312 0 412 2000
rect 468 0 568 2000
<< mvpdiff >>
rect -50 0 0 2000
rect 568 0 618 2000
<< poly >>
rect 0 2000 100 2026
rect 0 -26 100 0
rect 156 2000 256 2026
rect 156 -26 256 0
rect 312 2000 412 2026
rect 312 -26 412 0
rect 468 2000 568 2026
rect 468 -26 568 0
<< locali >>
rect -45 -4 -11 1966
rect 111 -4 145 1966
rect 267 -4 301 1966
rect 423 -4 457 1966
rect 579 -4 613 1966
use hvDFL1sd2_CDNS_52468879185623  hvDFL1sd2_CDNS_52468879185623_0
timestamp 1701704242
transform 1 0 412 0 1 0
box -36 -36 92 2036
use hvDFL1sd2_CDNS_52468879185623  hvDFL1sd2_CDNS_52468879185623_1
timestamp 1701704242
transform 1 0 256 0 1 0
box -36 -36 92 2036
use hvDFL1sd2_CDNS_52468879185623  hvDFL1sd2_CDNS_52468879185623_2
timestamp 1701704242
transform 1 0 100 0 1 0
box -36 -36 92 2036
use hvDFL1sd_CDNS_52468879185624  hvDFL1sd_CDNS_52468879185624_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 2036
use hvDFL1sd_CDNS_52468879185624  hvDFL1sd_CDNS_52468879185624_1
timestamp 1701704242
transform 1 0 568 0 1 0
box -36 -36 89 2036
<< labels >>
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
flabel comment s 128 981 128 981 0 FreeSans 300 0 0 0 D
flabel comment s 284 981 284 981 0 FreeSans 300 0 0 0 S
flabel comment s 440 981 440 981 0 FreeSans 300 0 0 0 D
flabel comment s 596 981 596 981 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 90863098
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90860580
<< end >>
