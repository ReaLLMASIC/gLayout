magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 125 197
<< metal1 >>
rect -6 197 131 200
rect -6 0 0 197
rect 125 0 131 197
rect -6 -3 131 0
<< properties >>
string GDS_END 86920416
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86918748
<< end >>
