magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -91 515 1147 1337
<< pwell >>
rect 109 367 243 455
rect 813 367 947 455
<< mvpsubdiff >>
rect 135 427 217 429
rect 135 393 159 427
rect 193 393 217 427
rect 839 427 921 429
rect 839 393 863 427
rect 897 393 921 427
<< mvnsubdiff >>
rect 135 583 159 617
rect 193 583 217 617
rect 135 581 217 583
rect 839 583 863 617
rect 897 583 921 617
rect 839 581 921 583
<< mvpsubdiffcont >>
rect 159 393 193 427
rect 863 393 897 427
<< mvnsubdiffcont >>
rect 159 583 193 617
rect 863 583 897 617
<< poly >>
rect 28 1353 328 1369
rect 28 1319 210 1353
rect 244 1319 278 1353
rect 312 1319 328 1353
rect 28 1297 328 1319
rect 550 1353 684 1369
rect 550 1319 566 1353
rect 600 1319 634 1353
rect 668 1319 684 1353
rect 550 1297 684 1319
rect 728 1353 1028 1369
rect 728 1319 744 1353
rect 778 1319 812 1353
rect 846 1319 1028 1353
rect 728 1297 1028 1319
rect 28 345 124 645
rect 228 345 324 645
rect 380 579 500 645
rect 380 545 427 579
rect 461 545 500 579
rect 380 511 500 545
rect 556 589 676 645
rect 556 517 828 589
rect 380 477 427 511
rect 461 477 500 511
rect 380 461 500 477
rect 380 401 676 461
rect 556 345 676 401
rect 732 345 828 517
rect 932 345 1028 645
rect 28 71 331 93
rect 28 37 213 71
rect 247 37 281 71
rect 315 37 331 71
rect 28 21 331 37
rect 373 71 507 93
rect 373 37 389 71
rect 423 37 457 71
rect 491 37 507 71
rect 373 21 507 37
rect 901 71 1035 93
rect 901 37 917 71
rect 951 37 985 71
rect 1019 37 1035 71
rect 901 21 1035 37
<< polycont >>
rect 210 1319 244 1353
rect 278 1319 312 1353
rect 566 1319 600 1353
rect 634 1319 668 1353
rect 744 1319 778 1353
rect 812 1319 846 1353
rect 427 545 461 579
rect 427 477 461 511
rect 213 37 247 71
rect 281 37 315 71
rect 389 37 423 71
rect 457 37 491 71
rect 917 37 951 71
rect 985 37 1019 71
<< locali >>
rect 210 1353 312 1369
rect 244 1319 278 1353
rect 210 1303 312 1319
rect 566 1353 668 1369
rect 600 1319 634 1353
rect 566 1303 668 1319
rect 744 1353 846 1369
rect 778 1319 812 1353
rect 744 1303 846 1319
rect 159 785 193 823
rect 159 713 193 751
rect -17 503 17 667
rect 159 567 193 583
rect 17 469 55 503
rect -17 219 17 469
rect 159 427 193 443
rect 159 259 193 297
rect 159 187 193 225
rect 227 87 301 1303
rect 411 559 427 579
rect 461 559 477 579
rect 405 545 427 559
rect 405 525 443 545
rect 411 511 477 525
rect 411 477 427 511
rect 461 477 477 511
rect 403 87 477 162
rect 511 121 545 1270
rect 579 503 653 1303
rect 613 469 651 503
rect 213 71 315 87
rect 389 71 491 87
rect 755 71 829 1303
rect 863 785 897 823
rect 863 713 897 751
rect 863 567 897 583
rect 1039 559 1073 667
rect 1001 525 1039 559
rect 863 427 897 443
rect 863 235 897 273
rect 1039 205 1073 525
rect 931 87 1005 163
rect 917 71 1019 87
rect 247 37 281 71
rect 423 37 457 71
rect 773 37 811 71
rect 951 37 985 71
rect 213 21 315 37
rect 389 21 491 37
rect 755 21 829 37
rect 917 21 1019 37
<< viali >>
rect 159 823 193 857
rect 159 751 193 785
rect 159 679 193 713
rect 159 617 193 633
rect 159 599 193 617
rect -17 469 17 503
rect 55 469 89 503
rect 159 393 193 411
rect 159 377 193 393
rect 159 297 193 331
rect 159 225 193 259
rect 159 153 193 187
rect 371 525 405 559
rect 443 545 461 559
rect 461 545 477 559
rect 443 525 477 545
rect 579 469 613 503
rect 651 469 685 503
rect 863 823 897 857
rect 863 751 897 785
rect 863 679 897 713
rect 863 617 897 633
rect 863 599 897 617
rect 967 525 1001 559
rect 1039 525 1073 559
rect 863 393 897 411
rect 863 377 897 393
rect 863 273 897 307
rect 863 201 897 235
rect 387 37 389 71
rect 389 37 421 71
rect 459 37 491 71
rect 491 37 493 71
rect 739 37 773 71
rect 811 37 845 71
rect 917 37 951 71
rect 989 37 1019 71
rect 1019 37 1023 71
<< metal1 >>
rect -25 857 1085 869
rect -25 823 159 857
rect 193 823 863 857
rect 897 823 1085 857
rect -25 785 1085 823
rect -25 751 159 785
rect 193 751 863 785
rect 897 751 1085 785
rect -25 713 1085 751
rect -25 679 159 713
rect 193 679 863 713
rect 897 679 1085 713
rect -25 667 1085 679
rect -25 633 1085 639
rect -25 599 159 633
rect 193 599 863 633
rect 897 599 1085 633
rect -25 593 1085 599
rect 359 559 1085 565
rect 359 525 371 559
rect 405 525 443 559
rect 477 537 967 559
rect 477 525 495 537
tri 495 525 507 537 nw
tri 937 525 949 537 ne
rect 949 525 967 537
rect 1001 525 1039 559
rect 1073 525 1085 559
rect 359 519 489 525
tri 489 519 495 525 nw
tri 949 519 955 525 ne
rect 955 519 1085 525
rect -29 503 101 509
tri 101 503 107 509 sw
tri 561 503 567 509 se
rect 567 503 697 509
rect -29 469 -17 503
rect 17 469 55 503
rect 89 491 107 503
tri 107 491 119 503 sw
tri 549 491 561 503 se
rect 561 491 579 503
rect 89 469 579 491
rect 613 469 651 503
rect 685 469 697 503
rect -29 463 697 469
rect -25 411 1085 417
rect -25 377 159 411
rect 193 377 863 411
rect 897 377 1085 411
rect -25 371 1085 377
rect -25 331 1085 343
rect -25 297 159 331
rect 193 307 1085 331
rect 193 297 863 307
rect -25 273 863 297
rect 897 273 1085 307
rect -25 259 1085 273
rect -25 225 159 259
rect 193 235 1085 259
rect 193 225 863 235
rect -25 201 863 225
rect 897 201 1085 235
rect -25 187 1085 201
rect -25 153 159 187
rect 193 153 1085 187
rect -25 141 1085 153
rect 375 71 1035 77
rect 375 37 387 71
rect 421 37 459 71
rect 493 37 739 71
rect 773 37 811 71
rect 845 37 917 71
rect 951 37 989 71
rect 1023 37 1035 71
rect 375 31 1035 37
use hvnTran_CDNS_524688791851398  hvnTran_CDNS_524688791851398_0
timestamp 1701704242
transform 1 0 732 0 -1 319
box -76 -26 375 226
use hvnTran_CDNS_524688791851399  hvnTran_CDNS_524688791851399_0
timestamp 1701704242
transform 1 0 380 0 -1 319
box -76 -26 372 226
use hvnTran_CDNS_524688791851400  hvnTran_CDNS_524688791851400_0
timestamp 1701704242
transform 1 0 28 0 -1 319
box -79 -26 372 226
use hvpTran_CDNS_524688791851401  hvpTran_CDNS_524688791851401_0
timestamp 1701704242
transform 1 0 28 0 1 671
box -119 -66 1119 666
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 477 0 1 525
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 1073 0 1 525
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 1023 0 -1 71
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 89 0 -1 503
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 845 0 -1 71
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform -1 0 685 0 -1 503
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform -1 0 493 0 -1 71
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 -1 897 1 0 201
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 193 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 193 1 0 679
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 897 1 0 679
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1701704242
transform 1 0 159 0 1 377
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1701704242
transform 1 0 863 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1701704242
transform 1 0 159 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1701704242
transform 1 0 863 0 1 377
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform -1 0 331 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1701704242
transform -1 0 328 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1701704242
transform -1 0 862 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1701704242
transform -1 0 684 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1701704242
transform 0 -1 477 1 0 461
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1701704242
transform 1 0 373 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1701704242
transform 1 0 901 0 1 21
box 0 0 1 1
<< labels >>
flabel metal1 s 1044 371 1056 417 3 FreeSans 200 180 0 0 vnb
port 1 nsew
flabel metal1 s 1044 593 1056 639 3 FreeSans 200 180 0 0 vpb
port 2 nsew
flabel metal1 s 1044 141 1056 343 3 FreeSans 200 180 0 0 vgnd
port 3 nsew
flabel metal1 s 1044 667 1056 869 3 FreeSans 200 180 0 0 vpwr
port 4 nsew
flabel metal1 s 0 141 12 343 3 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 0 371 12 417 3 FreeSans 200 0 0 0 vnb
port 1 nsew
flabel metal1 s 0 593 12 639 3 FreeSans 200 0 0 0 vpb
port 2 nsew
flabel metal1 s 0 667 12 869 3 FreeSans 200 0 0 0 vpwr
port 4 nsew
flabel locali s 778 1319 812 1369 0 FreeSans 200 0 0 0 in1
port 6 nsew
flabel locali s 423 21 457 71 0 FreeSans 200 0 0 0 in1
port 6 nsew
flabel locali s 775 21 809 71 0 FreeSans 200 0 0 0 in1
port 6 nsew
flabel locali s 951 21 985 71 0 FreeSans 200 0 0 0 in1
port 6 nsew
flabel locali s 244 1319 278 1369 0 FreeSans 200 0 0 0 in0
port 7 nsew
flabel locali s 247 21 281 71 0 FreeSans 200 0 0 0 in0
port 7 nsew
flabel locali s 511 1221 545 1270 0 FreeSans 200 0 0 0 out
port 8 nsew
flabel locali s 511 121 545 171 0 FreeSans 200 0 0 0 out
port 8 nsew
<< properties >>
string GDS_END 87669752
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87662850
<< end >>
