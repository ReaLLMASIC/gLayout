magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 116 26 197 44
<< poly >>
rect 28 3236 128 3252
rect 28 3202 61 3236
rect 95 3202 128 3236
rect 28 3168 128 3202
rect 28 3134 61 3168
rect 95 3134 128 3168
rect 28 3112 128 3134
rect 184 3236 284 3252
rect 184 3202 217 3236
rect 251 3202 284 3236
rect 184 3168 284 3202
rect 184 3134 217 3168
rect 251 3134 284 3168
rect 184 3112 284 3134
<< polycont >>
rect 61 3202 95 3236
rect 61 3134 95 3168
rect 217 3202 251 3236
rect 217 3134 251 3168
<< locali >>
rect 111 3270 149 3304
rect 45 3202 61 3236
rect 95 3202 111 3236
rect 45 3168 111 3202
rect 45 3134 61 3168
rect 95 3134 111 3168
rect 201 3202 217 3236
rect 251 3202 267 3236
rect 201 3168 267 3202
rect 201 3134 217 3168
rect 251 3134 267 3168
rect 51 2830 105 3134
rect 51 2796 71 2830
rect 51 2758 105 2796
rect 51 2724 71 2758
rect 207 2400 261 3134
rect 241 2366 261 2400
rect 207 2328 261 2366
rect 241 2294 261 2328
rect 17 1970 105 2260
rect 17 1936 71 1970
rect 17 1884 105 1936
rect 17 1850 71 1884
rect 17 1798 105 1850
rect 17 1764 71 1798
rect 17 1713 105 1764
rect 17 1679 71 1713
rect 17 1628 105 1679
rect 17 1594 71 1628
rect 17 400 105 1594
rect 207 1970 295 2260
rect 241 1936 295 1970
rect 207 1884 295 1936
rect 241 1850 295 1884
rect 207 1798 295 1850
rect 241 1764 295 1798
rect 207 1713 295 1764
rect 241 1679 295 1713
rect 207 1628 295 1679
rect 241 1594 295 1628
rect 139 1193 173 1236
rect 139 1116 173 1159
rect 139 1039 173 1082
rect 139 962 173 1005
rect 139 884 173 928
rect 139 806 173 850
rect 139 728 173 772
rect 139 650 173 694
rect 139 572 173 616
rect 139 494 173 538
rect 139 416 173 460
rect 207 400 295 1594
<< viali >>
rect 77 3270 111 3304
rect 149 3270 183 3304
rect 71 2796 105 2830
rect 71 2724 105 2758
rect 207 2366 241 2400
rect 207 2294 241 2328
rect 71 1936 105 1970
rect 71 1850 105 1884
rect 71 1764 105 1798
rect 71 1679 105 1713
rect 71 1594 105 1628
rect 207 1936 241 1970
rect 207 1850 241 1884
rect 207 1764 241 1798
rect 207 1679 241 1713
rect 207 1594 241 1628
rect 139 1236 173 1270
rect 139 1159 173 1193
rect 139 1082 173 1116
rect 139 1005 173 1039
rect 139 928 173 962
rect 139 850 173 884
rect 139 772 173 806
rect 139 694 173 728
rect 139 616 173 650
rect 139 538 173 572
rect 139 460 173 494
rect 139 382 173 416
<< metal1 >>
rect 65 3304 195 3310
rect 65 3270 77 3304
rect 111 3270 149 3304
rect 183 3270 195 3304
rect 65 3264 195 3270
rect 65 3144 123 3264
tri 123 3239 148 3264 nw
rect 66 3142 122 3143
rect 65 2842 123 3142
rect 66 2841 122 2842
rect 65 2830 123 2840
rect 65 2796 71 2830
rect 105 2796 123 2830
rect 65 2758 123 2796
rect 65 2724 71 2758
rect 105 2754 123 2758
tri 123 2754 148 2779 sw
rect 105 2724 241 2754
rect 65 2714 241 2724
rect 65 2712 201 2714
rect 202 2712 240 2713
rect 202 2411 240 2412
rect 241 2410 245 2412
rect 247 2411 487 2412
rect 201 2400 245 2410
rect 201 2366 207 2400
rect 241 2366 245 2400
rect 201 2328 245 2366
rect 201 2294 207 2328
rect 241 2294 245 2328
rect 201 2282 245 2294
rect 246 2283 488 2411
rect 247 2282 487 2283
rect 489 2282 601 2412
rect -277 1982 -235 1995
rect -277 1582 -237 1982
rect -236 1583 -235 1981
rect 65 1583 66 1981
rect 67 1970 319 1982
rect 321 1981 481 1982
rect 67 1936 71 1970
rect 105 1936 207 1970
rect 241 1936 319 1970
rect 67 1884 319 1936
rect 67 1850 71 1884
rect 105 1850 207 1884
rect 241 1850 319 1884
rect 67 1798 319 1850
rect 67 1764 71 1798
rect 105 1764 207 1798
rect 241 1764 319 1798
rect 67 1713 319 1764
rect 67 1679 71 1713
rect 105 1679 207 1713
rect 241 1679 319 1713
rect 67 1628 319 1679
rect 67 1594 71 1628
rect 105 1594 207 1628
rect 241 1594 319 1628
rect 67 1582 319 1594
rect 320 1583 482 1981
rect 321 1582 481 1583
rect 483 1582 603 1982
rect -277 1569 -235 1582
rect 133 1270 179 1282
rect 133 1236 139 1270
rect 173 1236 179 1270
rect 133 1193 179 1236
rect 133 1159 139 1193
rect 173 1159 179 1193
rect 133 1116 179 1159
rect 133 1082 139 1116
rect 173 1082 179 1116
rect 133 1039 179 1082
rect 133 1005 139 1039
rect 173 1005 179 1039
rect 133 962 179 1005
rect 133 928 139 962
rect 173 928 179 962
rect 133 884 179 928
rect 133 850 139 884
rect 173 850 179 884
rect 133 806 179 850
rect 133 772 139 806
rect 173 772 179 806
rect 133 728 179 772
rect 133 694 139 728
rect 173 694 179 728
rect 133 650 179 694
rect 133 616 139 650
rect 173 616 179 650
rect 133 572 179 616
rect 133 538 139 572
rect 173 538 179 572
rect 133 494 179 538
rect 133 460 139 494
rect 173 460 179 494
rect 133 416 179 460
rect 133 382 139 416
rect 173 382 179 416
rect 133 370 179 382
<< rmetal1 >>
rect 65 3143 123 3144
rect 65 3142 66 3143
rect 122 3142 123 3143
rect 65 2841 66 2842
rect 122 2841 123 2842
rect 65 2840 123 2841
rect 201 2713 241 2714
rect 201 2712 202 2713
rect 240 2712 241 2713
rect 201 2411 202 2412
rect 240 2411 241 2412
rect 201 2410 241 2411
rect 245 2411 247 2412
rect 487 2411 489 2412
rect 245 2283 246 2411
rect 488 2283 489 2411
rect 245 2282 247 2283
rect 487 2282 489 2283
rect -237 1981 -235 1982
rect -237 1583 -236 1981
rect -237 1582 -235 1583
rect 65 1981 67 1982
rect 66 1583 67 1981
rect 319 1981 321 1982
rect 481 1981 483 1982
rect 65 1582 67 1583
rect 319 1583 320 1981
rect 482 1583 483 1981
rect 319 1582 321 1583
rect 481 1582 483 1583
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 1 0 77 0 1 3270
box 0 0 1 1
use L1M1_CDNS_524688791851450  L1M1_CDNS_524688791851450_0
timestamp 1701704242
transform -1 0 241 0 1 2294
box 0 0 1 1
use L1M1_CDNS_524688791851450  L1M1_CDNS_524688791851450_1
timestamp 1701704242
transform 1 0 71 0 1 2724
box 0 0 1 1
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_0
timestamp 1701704242
transform -1 0 284 0 -1 3086
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_1
timestamp 1701704242
transform 1 0 28 0 -1 3086
box -119 -66 219 3066
use PYL1_CDNS_524688791851449  PYL1_CDNS_524688791851449_0
timestamp 1701704242
transform -1 0 267 0 1 3118
box 0 0 1 1
use PYL1_CDNS_524688791851449  PYL1_CDNS_524688791851449_1
timestamp 1701704242
transform 1 0 45 0 1 3118
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851454  sky130_fd_io__tk_em1o_CDNS_524688791851454_0
timestamp 1701704242
transform 1 0 -289 0 1 1582
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851455  sky130_fd_io__tk_em1o_CDNS_524688791851455_0
timestamp 1701704242
transform 0 1 201 -1 0 2766
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851451  sky130_fd_io__tk_em1s_CDNS_524688791851451_0
timestamp 1701704242
transform 0 1 65 -1 0 3196
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851452  sky130_fd_io__tk_em1s_CDNS_524688791851452_0
timestamp 1701704242
transform 1 0 193 0 -1 2412
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851453  sky130_fd_io__tk_em1s_CDNS_524688791851453_0
timestamp 1701704242
transform 1 0 267 0 1 1582
box 0 0 1 1
<< labels >>
flabel comment s 221 2558 221 2558 0 FreeSans 200 90 0 0 metal open element
flabel metal1 s -275 1582 -239 1975 0 FreeSans 400 90 0 0 pad
port 3 nsew
flabel metal1 s 566 1582 601 1982 0 FreeSans 400 90 0 0 tie_hi
port 4 nsew
flabel metal1 s 73 3148 115 3256 0 FreeSans 400 90 0 0 padlo
port 2 nsew
flabel metal1 s 562 2288 601 2406 0 FreeSans 400 270 0 0 tie_hi
port 4 nsew
flabel metal1 s 133 1236 179 1282 7 FreeSans 200 90 0 0 pug_h
port 1 nsew
flabel nwell s 116 26 197 44 0 FreeSans 200 0 0 0 vpb_drvr
port 5 nsew
<< properties >>
string GDS_END 88515310
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88510856
string path 2.200 49.550 2.200 39.550 
<< end >>
