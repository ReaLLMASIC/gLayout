magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -122 -66 282 1466
<< mvpmos >>
rect 0 0 160 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 160 0 210 1400
<< poly >>
rect 0 1400 160 1432
rect 0 -32 160 0
<< locali >>
rect -45 -4 -11 1354
rect 171 -4 205 1354
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 92 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_1
timestamp 1701704242
transform 1 0 160 0 1 0
box -36 -36 92 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 D
flabel comment s 188 675 188 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85593044
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85592026
<< end >>
