magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -117 -26 196 1026
<< mvnmos >>
rect 0 0 120 1000
<< mvndiff >>
rect -91 0 0 1000
rect 120 0 170 1000
<< poly >>
rect 0 1000 120 1032
rect 0 -32 120 0
<< metal1 >>
rect -244 -16 -198 978
use hvDFTPM1s2_CDNS_5246887918513  hvDFTPM1s2_CDNS_5246887918513_0
timestamp 1701704242
transform -1 0 -91 0 1 0
box -26 -26 286 1026
<< labels >>
flabel comment s -221 481 -221 481 0 FreeSans 300 0 0 0 S
flabel comment s 145 500 145 500 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 13691996
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 13691156
<< end >>
