magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 413 53
<< metal1 >>
rect -6 53 419 56
rect -6 0 0 53
rect 413 0 419 53
rect -6 -3 419 0
<< properties >>
string GDS_END 88082842
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88081174
<< end >>
