magic
tech sky130A
timestamp 1701704242
<< metal1 >>
rect 0 0 3 58
rect 477 0 480 58
<< via1 >>
rect 3 0 477 58
<< metal2 >>
rect 0 0 3 58
rect 477 0 480 58
<< properties >>
string GDS_END 78481730
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78479678
<< end >>
