magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 3228 -69 5041 1827
<< nwell >>
rect 1025 1311 1671 1493
rect 1489 1241 1671 1311
rect 1489 1059 1992 1241
rect 1519 237 1992 1059
rect 2660 237 3354 1059
<< pwell >>
rect 4077 1351 4757 1437
<< mvpsubdiff >>
rect 4103 1377 4127 1411
rect 4161 1377 4196 1411
rect 4230 1377 4265 1411
rect 4299 1377 4333 1411
rect 4367 1377 4401 1411
rect 4435 1377 4469 1411
rect 4503 1377 4537 1411
rect 4571 1377 4605 1411
rect 4639 1377 4673 1411
rect 4707 1377 4731 1411
<< mvnsubdiff >>
rect 1091 1419 1605 1427
rect 1091 1385 1115 1419
rect 1149 1385 1183 1419
rect 1217 1385 1251 1419
rect 1285 1385 1319 1419
rect 1353 1385 1387 1419
rect 1421 1385 1455 1419
rect 1489 1403 1605 1419
rect 1489 1385 1563 1403
rect 1091 1377 1563 1385
rect 1555 1369 1563 1377
rect 1597 1369 1605 1403
rect 1555 1335 1605 1369
rect 1555 1301 1563 1335
rect 1597 1301 1605 1335
rect 1555 1267 1605 1301
rect 1555 1233 1563 1267
rect 1597 1233 1605 1267
rect 1555 1175 1605 1233
rect 1555 1167 1926 1175
rect 1555 1133 1579 1167
rect 1613 1133 1647 1167
rect 1681 1133 1715 1167
rect 1749 1133 1783 1167
rect 1817 1133 1851 1167
rect 1885 1133 1926 1167
rect 1555 1125 1926 1133
<< mvpsubdiffcont >>
rect 4127 1377 4161 1411
rect 4196 1377 4230 1411
rect 4265 1377 4299 1411
rect 4333 1377 4367 1411
rect 4401 1377 4435 1411
rect 4469 1377 4503 1411
rect 4537 1377 4571 1411
rect 4605 1377 4639 1411
rect 4673 1377 4707 1411
<< mvnsubdiffcont >>
rect 1115 1385 1149 1419
rect 1183 1385 1217 1419
rect 1251 1385 1285 1419
rect 1319 1385 1353 1419
rect 1387 1385 1421 1419
rect 1455 1385 1489 1419
rect 1563 1369 1597 1403
rect 1563 1301 1597 1335
rect 1563 1233 1597 1267
rect 1579 1133 1613 1167
rect 1647 1133 1681 1167
rect 1715 1133 1749 1167
rect 1783 1133 1817 1167
rect 1851 1133 1885 1167
<< poly >>
rect 3530 1537 3664 1553
rect 3530 1503 3546 1537
rect 3580 1503 3614 1537
rect 3648 1503 3664 1537
rect 3530 1487 3664 1503
rect 3706 1537 3840 1553
rect 3706 1503 3722 1537
rect 3756 1503 3790 1537
rect 3824 1503 3840 1537
rect 3706 1487 3840 1503
rect 3537 1481 3657 1487
rect 3713 1481 3833 1487
rect 3537 764 3657 770
rect 3713 764 3833 770
rect 3530 748 3664 764
rect 3530 714 3546 748
rect 3580 714 3614 748
rect 3648 714 3664 748
rect 3530 698 3664 714
rect 3706 748 3840 764
rect 3706 714 3722 748
rect 3756 714 3790 748
rect 3824 714 3840 748
rect 3706 698 3840 714
rect 1577 271 1697 277
rect 1753 271 1873 277
rect 2779 271 2899 277
rect 2955 271 3075 277
rect 1110 255 1244 271
rect 1110 221 1126 255
rect 1160 221 1194 255
rect 1228 221 1244 255
rect 1110 205 1244 221
rect 1300 255 1434 271
rect 1300 221 1316 255
rect 1350 221 1384 255
rect 1418 221 1434 255
rect 1300 205 1434 221
rect 1570 255 1704 271
rect 1570 221 1586 255
rect 1620 221 1654 255
rect 1688 221 1704 255
rect 1570 205 1704 221
rect 1746 255 1880 271
rect 1746 221 1762 255
rect 1796 221 1830 255
rect 1864 221 1880 255
rect 1746 205 1880 221
rect 2772 255 2906 271
rect 2772 221 2788 255
rect 2822 221 2856 255
rect 2890 221 2906 255
rect 2772 205 2906 221
rect 2948 255 3082 271
rect 2948 221 2964 255
rect 2998 221 3032 255
rect 3066 221 3082 255
rect 2948 205 3082 221
rect 4126 255 4260 271
rect 4126 221 4142 255
rect 4176 221 4210 255
rect 4244 221 4260 255
rect 4126 205 4260 221
rect 4316 255 4450 271
rect 4316 221 4332 255
rect 4366 221 4400 255
rect 4434 221 4450 255
rect 4316 205 4450 221
rect 4593 255 4727 271
rect 4593 221 4609 255
rect 4643 221 4677 255
rect 4711 221 4727 255
rect 4593 205 4727 221
<< polycont >>
rect 3546 1503 3580 1537
rect 3614 1503 3648 1537
rect 3722 1503 3756 1537
rect 3790 1503 3824 1537
rect 3546 714 3580 748
rect 3614 714 3648 748
rect 3722 714 3756 748
rect 3790 714 3824 748
rect 1126 221 1160 255
rect 1194 221 1228 255
rect 1316 221 1350 255
rect 1384 221 1418 255
rect 1586 221 1620 255
rect 1654 221 1688 255
rect 1762 221 1796 255
rect 1830 221 1864 255
rect 2788 221 2822 255
rect 2856 221 2890 255
rect 2964 221 2998 255
rect 3032 221 3066 255
rect 4142 221 4176 255
rect 4210 221 4244 255
rect 4332 221 4366 255
rect 4400 221 4434 255
rect 4609 221 4643 255
rect 4677 221 4711 255
<< locali >>
rect 3340 1537 3648 1553
rect 3340 1503 3546 1537
rect 3580 1503 3614 1537
rect 3340 1487 3648 1503
rect 3722 1537 3824 1553
rect 3756 1503 3790 1537
rect 3722 1487 3824 1503
rect 1091 1419 1605 1427
rect 1091 1385 1115 1419
rect 1149 1385 1183 1419
rect 1217 1385 1251 1419
rect 1285 1385 1319 1419
rect 1353 1385 1387 1419
rect 1421 1385 1455 1419
rect 1489 1403 1605 1419
rect 1489 1385 1563 1403
rect 1091 1377 1563 1385
rect 1555 1369 1563 1377
rect 1597 1369 1605 1403
rect 1555 1335 1605 1369
rect 1555 1301 1563 1335
rect 1597 1301 1605 1335
rect 1555 1267 1605 1301
rect 1555 1233 1563 1267
rect 1597 1233 1605 1267
rect 1555 1175 1605 1233
rect 1555 1167 1926 1175
rect 1555 1133 1579 1167
rect 1613 1133 1647 1167
rect 1681 1133 1715 1167
rect 1749 1133 1783 1167
rect 1817 1133 1851 1167
rect 1885 1133 1926 1167
rect 2696 1138 2734 1172
rect 2980 1138 3018 1172
rect 1555 1125 1926 1133
rect 1532 998 1566 1036
rect 1099 581 1133 619
rect 1366 528 1478 543
rect 1400 494 1444 528
rect 1366 479 1478 494
rect 1223 412 1335 427
rect 1257 378 1301 412
rect 1223 363 1335 378
rect 1532 304 1566 964
rect 1652 895 1742 1125
rect 1652 861 1708 895
rect 1652 823 1742 861
rect 1652 789 1708 823
rect 1652 751 1742 789
rect 1652 717 1708 751
rect 1652 327 1742 717
rect 1810 1036 1850 1070
rect 1776 998 1850 1036
rect 1810 964 1850 998
rect 1776 271 1850 964
rect 1918 980 1956 1014
rect 1884 304 1934 980
rect 2734 304 2768 1138
rect 2910 895 2944 907
rect 2910 823 2944 861
rect 2910 751 2944 789
rect 2910 705 2944 717
rect 1586 255 1688 271
rect 1110 221 1126 255
rect 1160 221 1194 255
rect 1228 221 1244 255
rect 1300 221 1310 255
rect 1350 221 1382 255
rect 1418 221 1434 255
rect 1620 221 1654 255
rect 1762 255 1864 271
rect 1796 221 1830 255
rect 1900 255 1934 304
rect 2978 271 3052 1138
rect 3086 307 3139 907
rect 3238 823 3272 861
rect 3238 751 3272 789
rect 3086 304 3105 307
rect 2788 255 2890 271
rect 1934 221 1972 255
rect 2822 221 2856 255
rect 1122 47 1228 221
rect 1156 13 1194 47
rect 1586 47 1692 221
rect 1762 205 1864 221
rect 2788 205 2890 221
rect 2964 255 3066 271
rect 2998 221 3032 255
rect 2964 205 3066 221
rect 3105 235 3139 273
rect 3340 149 3414 1487
rect 3492 1172 3526 1453
rect 3668 1349 3702 1387
rect 3668 1277 3702 1315
rect 3736 1172 3810 1487
rect 3878 1251 3969 1453
rect 4103 1377 4104 1411
rect 4161 1377 4177 1411
rect 4230 1377 4250 1411
rect 4299 1377 4323 1411
rect 4367 1377 4395 1411
rect 4435 1377 4467 1411
rect 4503 1377 4537 1411
rect 4573 1377 4605 1411
rect 4645 1377 4673 1411
rect 4717 1377 4731 1411
rect 3526 1138 3564 1172
rect 3738 1138 3776 1172
rect 3526 1059 3564 1093
rect 3738 1059 3776 1093
rect 3492 798 3526 1059
rect 3668 912 3702 996
rect 3668 840 3702 878
rect 3736 764 3810 1059
rect 3844 936 3878 974
rect 3546 748 3648 764
rect 3580 714 3614 748
rect 3546 698 3648 714
rect 3722 748 3824 764
rect 3756 714 3790 748
rect 3722 698 3824 714
rect 3556 154 3630 698
rect 3935 255 3969 1251
rect 4707 1235 4741 1273
rect 4379 644 4492 659
rect 4413 610 4458 644
rect 4379 595 4492 610
rect 4080 528 4187 543
rect 4114 494 4153 528
rect 4080 479 4187 494
rect 4234 412 4346 427
rect 4268 378 4312 412
rect 4234 363 4346 378
rect 4512 412 4624 427
rect 4546 378 4590 412
rect 4512 363 4624 378
rect 3878 221 3916 255
rect 3950 221 3969 255
rect 4126 221 4142 255
rect 4176 221 4210 255
rect 4248 221 4260 255
rect 4316 221 4332 255
rect 4366 221 4400 255
rect 4438 221 4450 255
rect 4593 221 4609 255
rect 4643 221 4677 255
rect 4715 221 4727 255
rect 3935 215 3969 221
rect 4622 154 4696 221
rect 3374 115 3412 149
rect 3340 114 3414 115
rect 3556 80 4696 154
rect 1620 13 1658 47
<< viali >>
rect 2662 1138 2696 1172
rect 2734 1138 2768 1172
rect 2946 1138 2980 1172
rect 3018 1138 3052 1172
rect 1532 1036 1566 1070
rect 1532 964 1566 998
rect 1099 619 1133 653
rect 1099 547 1133 581
rect 1366 494 1400 528
rect 1444 494 1478 528
rect 1223 378 1257 412
rect 1301 378 1335 412
rect 1708 861 1742 895
rect 1708 789 1742 823
rect 1708 717 1742 751
rect 1776 1036 1810 1070
rect 1776 964 1810 998
rect 1884 980 1918 1014
rect 1956 980 1990 1014
rect 2910 861 2944 895
rect 2910 789 2944 823
rect 2910 717 2944 751
rect 1310 221 1316 255
rect 1316 221 1344 255
rect 1382 221 1384 255
rect 1384 221 1416 255
rect 3238 861 3272 895
rect 3238 789 3272 823
rect 3238 717 3272 751
rect 3105 273 3139 307
rect 1900 221 1934 255
rect 1972 221 2006 255
rect 2784 221 2788 255
rect 2788 221 2818 255
rect 2856 221 2890 255
rect 1122 13 1156 47
rect 1194 13 1228 47
rect 3105 201 3139 235
rect 3668 1387 3702 1421
rect 3668 1315 3702 1349
rect 3668 1243 3702 1277
rect 4104 1377 4127 1411
rect 4127 1377 4138 1411
rect 4177 1377 4196 1411
rect 4196 1377 4211 1411
rect 4250 1377 4265 1411
rect 4265 1377 4284 1411
rect 4323 1377 4333 1411
rect 4333 1377 4357 1411
rect 4395 1377 4401 1411
rect 4401 1377 4429 1411
rect 4467 1377 4469 1411
rect 4469 1377 4501 1411
rect 4539 1377 4571 1411
rect 4571 1377 4573 1411
rect 4611 1377 4639 1411
rect 4639 1377 4645 1411
rect 4683 1377 4707 1411
rect 4707 1377 4717 1411
rect 3492 1138 3526 1172
rect 3564 1138 3598 1172
rect 3704 1138 3738 1172
rect 3776 1138 3810 1172
rect 3492 1059 3526 1093
rect 3564 1059 3598 1093
rect 3704 1059 3738 1093
rect 3776 1059 3810 1093
rect 3668 878 3702 912
rect 3668 806 3702 840
rect 3844 974 3878 1008
rect 3844 902 3878 936
rect 4707 1273 4741 1307
rect 4707 1201 4741 1235
rect 4379 610 4413 644
rect 4458 610 4492 644
rect 4080 494 4114 528
rect 4153 494 4187 528
rect 4234 378 4268 412
rect 4312 378 4346 412
rect 4512 378 4546 412
rect 4590 378 4624 412
rect 3844 221 3878 255
rect 3916 221 3950 255
rect 4142 221 4176 255
rect 4214 221 4244 255
rect 4244 221 4248 255
rect 4332 221 4366 255
rect 4404 221 4434 255
rect 4434 221 4438 255
rect 4609 221 4643 255
rect 4681 221 4711 255
rect 4711 221 4715 255
rect 3340 115 3374 149
rect 3412 115 3446 149
rect 1586 13 1620 47
rect 1658 13 1692 47
<< metal1 >>
rect 3328 1421 4979 1433
rect 3328 1387 3668 1421
rect 3702 1411 4979 1421
rect 3702 1387 4104 1411
rect 3328 1377 4104 1387
rect 4138 1377 4177 1411
rect 4211 1377 4250 1411
rect 4284 1377 4323 1411
rect 4357 1377 4395 1411
rect 4429 1377 4467 1411
rect 4501 1377 4539 1411
rect 4573 1377 4611 1411
rect 4645 1377 4683 1411
rect 4717 1377 4979 1411
rect 3328 1349 4979 1377
rect 3328 1315 3668 1349
rect 3702 1315 4979 1349
rect 3328 1307 4979 1315
rect 3328 1277 4707 1307
rect 3328 1243 3668 1277
rect 3702 1273 4707 1277
rect 4741 1273 4979 1307
rect 3702 1243 4979 1273
rect 3328 1235 4979 1243
rect 3328 1218 4707 1235
tri 3887 1201 3904 1218 ne
rect 3904 1201 4147 1218
tri 4147 1201 4164 1218 nw
tri 4672 1201 4689 1218 ne
rect 4689 1201 4707 1218
rect 4741 1218 4979 1235
rect 4741 1201 4747 1218
tri 3904 1178 3927 1201 ne
rect 3927 1178 4105 1201
rect 2650 1172 3822 1178
rect 2650 1138 2662 1172
rect 2696 1138 2734 1172
rect 2768 1138 2946 1172
rect 2980 1138 3018 1172
rect 3052 1138 3492 1172
rect 3526 1138 3564 1172
rect 3598 1138 3704 1172
rect 3738 1138 3776 1172
rect 3810 1138 3822 1172
tri 3927 1159 3946 1178 ne
rect 2650 1132 3822 1138
rect 1526 1093 3822 1099
rect 1526 1070 3492 1093
rect 1526 1036 1532 1070
rect 1566 1053 1776 1070
rect 1566 1036 1607 1053
tri 1607 1036 1624 1053 nw
tri 1718 1036 1735 1053 ne
rect 1735 1036 1776 1053
rect 1810 1059 3492 1070
rect 3526 1059 3564 1093
rect 3598 1059 3704 1093
rect 3738 1059 3776 1093
rect 3810 1059 3822 1093
rect 1810 1053 3822 1059
rect 1810 1036 1825 1053
rect 1526 1014 1585 1036
tri 1585 1014 1607 1036 nw
tri 1735 1014 1757 1036 ne
rect 1757 1014 1825 1036
tri 1825 1014 1864 1053 nw
rect 1872 1014 3884 1020
rect 1526 998 1572 1014
tri 1572 1001 1585 1014 nw
tri 1757 1005 1766 1014 ne
rect 1766 1005 1816 1014
tri 1816 1005 1825 1014 nw
tri 1766 1001 1770 1005 ne
rect 1526 964 1532 998
rect 1566 964 1572 998
rect 1526 952 1572 964
rect 1770 998 1816 1005
rect 1770 964 1776 998
rect 1810 964 1816 998
rect 1872 980 1884 1014
rect 1918 980 1956 1014
rect 1990 1008 3884 1014
rect 1990 980 3844 1008
rect 1872 974 3844 980
rect 3878 974 3884 1008
rect 1770 952 1816 964
tri 3786 952 3808 974 ne
rect 3808 952 3884 974
tri 3808 936 3824 952 ne
rect 3824 936 3884 952
tri 3824 924 3836 936 ne
rect 3836 924 3844 936
rect 3662 912 3708 924
tri 3836 922 3838 924 ne
rect 1529 895 1901 907
rect 1529 861 1708 895
rect 1742 861 1901 895
rect 1529 823 1901 861
rect 1529 789 1708 823
rect 1742 789 1901 823
rect 1529 751 1901 789
rect 1529 717 1708 751
rect 1742 717 1901 751
rect 1529 705 1901 717
rect 2751 895 3306 907
rect 2751 861 2910 895
rect 2944 861 3238 895
rect 3272 861 3306 895
rect 2751 823 3306 861
rect 2751 789 2910 823
rect 2944 789 3238 823
rect 3272 789 3306 823
rect 3662 878 3668 912
rect 3702 907 3708 912
tri 3708 907 3711 910 sw
rect 3702 902 3711 907
tri 3711 902 3716 907 sw
rect 3838 902 3844 924
rect 3878 902 3884 936
tri 3943 907 3946 910 se
rect 3946 907 4105 1178
tri 4105 1159 4147 1201 nw
tri 4689 1189 4701 1201 ne
rect 4701 1189 4747 1201
tri 4747 1189 4776 1218 nw
rect 3702 878 3716 902
rect 3662 858 3716 878
tri 3716 858 3760 902 sw
rect 3838 890 3884 902
tri 3926 890 3943 907 se
rect 3943 890 4105 907
tri 3894 858 3926 890 se
rect 3926 858 4105 890
rect 3662 840 4105 858
rect 3662 806 3668 840
rect 3702 806 4105 840
rect 3662 794 4105 806
rect 2751 751 3306 789
rect 2751 717 2910 751
rect 2944 717 3238 751
rect 3272 717 3306 751
rect 2751 705 3306 717
rect 1093 653 4542 665
rect 1093 619 1099 653
rect 1133 644 4542 653
rect 1133 619 4379 644
rect 1093 610 4379 619
rect 4413 610 4458 644
rect 4492 610 4542 644
rect 1093 589 4542 610
rect 1093 581 1139 589
rect 1093 547 1099 581
rect 1133 547 1139 581
rect 1093 535 1139 547
tri 1139 535 1193 589 nw
rect 1354 528 4251 549
rect 1354 494 1366 528
rect 1400 494 1444 528
rect 1478 494 4080 528
rect 4114 494 4153 528
rect 4187 494 4251 528
rect 1354 473 4251 494
rect 1211 412 4728 433
rect 1211 378 1223 412
rect 1257 378 1301 412
rect 1335 378 4234 412
rect 4268 378 4312 412
rect 4346 378 4512 412
rect 4546 378 4590 412
rect 4624 378 4728 412
rect 1211 357 4728 378
rect 3099 307 3145 319
rect 3099 273 3105 307
rect 3139 273 3145 307
rect 3099 261 3145 273
tri 3145 261 3203 319 sw
rect 1298 255 2018 261
rect 1298 221 1310 255
rect 1344 221 1382 255
rect 1416 221 1900 255
rect 1934 221 1972 255
rect 2006 221 2018 255
rect 1298 215 2018 221
rect 2772 255 2902 261
rect 2772 221 2784 255
rect 2818 221 2856 255
rect 2890 221 2902 255
tri 2769 201 2772 204 se
rect 2772 201 2902 221
rect 3099 255 4260 261
rect 3099 235 3844 255
tri 2902 201 2905 204 sw
rect 3099 201 3105 235
rect 3139 221 3844 235
rect 3878 221 3916 255
rect 3950 221 4142 255
rect 4176 221 4214 255
rect 4248 221 4260 255
rect 3139 215 4260 221
rect 4320 255 4450 261
rect 4320 221 4332 255
rect 4366 221 4404 255
rect 4438 221 4450 255
rect 3139 201 3145 215
tri 2723 155 2769 201 se
rect 2769 189 2905 201
tri 2905 189 2917 201 sw
rect 3099 189 3145 201
tri 3145 189 3171 215 nw
rect 2769 184 2917 189
tri 2917 184 2922 189 sw
rect 2769 167 2922 184
tri 2922 167 2939 184 sw
tri 4303 167 4320 184 se
rect 4320 167 4450 221
rect 4597 255 4727 261
rect 4597 221 4609 255
rect 4643 221 4681 255
rect 4715 221 4727 255
rect 4597 215 4727 221
tri 4597 167 4645 215 ne
rect 2769 155 2939 167
tri 2939 155 2951 167 sw
tri 4291 155 4303 167 se
rect 4303 155 4450 167
rect 1110 149 4450 155
rect 1110 115 3340 149
rect 3374 115 3412 149
rect 3446 115 4450 149
rect 1110 109 4450 115
tri 4597 53 4645 101 se
rect 4645 53 4691 215
tri 4691 179 4727 215 nw
rect 1110 47 4691 53
rect 1110 13 1122 47
rect 1156 13 1194 47
rect 1228 13 1586 47
rect 1620 13 1658 47
rect 1692 13 4691 47
rect 1110 7 4691 13
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_0
timestamp 1701704242
transform -1 0 3657 0 1 1255
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_1
timestamp 1701704242
transform -1 0 3657 0 -1 996
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_2
timestamp 1701704242
transform 1 0 3713 0 -1 996
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_3
timestamp 1701704242
transform 1 0 3713 0 1 1255
box -79 -26 199 226
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_0
timestamp 1701704242
transform -1 0 1697 0 -1 903
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_1
timestamp 1701704242
transform -1 0 2899 0 -1 903
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_2
timestamp 1701704242
transform 1 0 2955 0 -1 903
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_3
timestamp 1701704242
transform 1 0 1753 0 -1 903
box -119 -66 239 666
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 2944 -1 0 895
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 1 1708 -1 0 895
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 1 2910 -1 0 895
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform 0 1 3668 1 0 1243
box 0 0 1 1
use nfet_CDNS_52468879185934  nfet_CDNS_52468879185934_0
timestamp 1701704242
transform -1 0 4696 0 -1 1303
box -79 -32 179 1032
use nfet_CDNS_52468879185935  nfet_CDNS_52468879185935_0
timestamp 1701704242
transform -1 0 4416 0 -1 1303
box -79 -32 179 1032
use nfet_CDNS_52468879185935  nfet_CDNS_52468879185935_1
timestamp 1701704242
transform 1 0 4160 0 -1 1303
box -79 -32 179 1032
use pfet_CDNS_52468879185933  pfet_CDNS_52468879185933_0
timestamp 1701704242
transform 1 0 1144 0 -1 1303
box -119 -66 375 1066
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform -1 0 3082 0 1 205
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1701704242
transform -1 0 1880 0 1 205
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1701704242
transform -1 0 3840 0 1 698
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1701704242
transform -1 0 3840 0 -1 1553
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1701704242
transform 1 0 3530 0 -1 1553
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1701704242
transform 1 0 3530 0 1 698
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1701704242
transform 1 0 1570 0 1 205
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1701704242
transform 1 0 2772 0 1 205
box 0 0 1 1
<< labels >>
flabel comment s 3262 578 3262 578 0 FreeSans 200 90 0 0 lv_net
flabel comment s 1705 1148 1705 1148 0 FreeSans 200 180 0 0 lv_net
flabel metal1 s 1509 244 1509 244 0 FreeSans 520 0 0 0 sel_vdda_buf
flabel metal1 s 3623 1268 3755 1378 0 FreeSans 500 0 0 0 vssa
port 2 nsew
flabel metal1 s 2962 765 3072 855 0 FreeSans 500 0 0 0 vswitch
port 3 nsew
flabel metal1 s 1606 820 1666 866 0 FreeSans 520 0 0 0 vdda
port 5 nsew
flabel metal1 s 2513 109 2664 155 0 FreeSans 520 0 0 0 sel_vddio
port 6 nsew
flabel metal1 s 2512 7 2612 53 0 FreeSans 520 0 0 0 sel_vdda
port 7 nsew
flabel metal1 s 3235 473 3335 549 0 FreeSans 500 0 0 0 out
port 1 nsew
flabel metal1 s 3233 589 3321 665 0 FreeSans 500 0 0 0 in
port 4 nsew
<< properties >>
string GDS_END 80588872
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80568152
string path 26.625 35.050 39.500 35.050 39.500 28.750 48.800 28.750 
<< end >>
