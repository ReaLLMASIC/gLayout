magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -68 -26 4068 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 4000 50 4042 66
rect 4034 16 4042 50
rect 4000 0 4042 16
<< ndiffc >>
rect -34 16 0 50
rect 4000 16 4034 50
<< ndiffres >>
rect 0 0 4000 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 4000 50 4034 66
rect 4000 0 4034 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1701704242
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1701704242
transform 1 0 3992 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 86204744
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86204242
<< end >>
