magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 13011 30757 14335 31063
rect 14029 26640 14335 30757
rect 9725 26334 14335 26640
rect 11329 452 11435 858
rect 13345 452 13451 858
<< pwell >>
rect 9851 35709 14455 36409
rect 9851 35708 10931 35709
rect 13139 31123 14455 35709
rect 9851 30390 13969 30696
rect 9851 26998 10561 30390
rect 13677 26998 13969 30390
rect 9851 26700 13969 26998
rect 9851 24830 14455 26274
rect 9851 24183 11258 24830
rect 13969 24805 14455 24830
rect 14181 24373 14455 24805
rect 9851 23071 10851 24183
rect 14145 23071 14455 24373
rect 9851 22901 14455 23071
rect 9851 22523 12477 22901
rect 13574 22023 14455 22901
rect 13743 21471 14455 22023
rect 13575 20842 14455 21471
rect 11339 1432 11483 1518
rect 13297 1432 13441 1518
rect 11339 1008 11425 1432
rect 13355 1008 13441 1432
<< psubdiff >>
rect 11365 1468 11457 1492
rect 11399 1458 11457 1468
rect 13323 1468 13415 1492
rect 13323 1458 13381 1468
rect 11365 1393 11399 1434
rect 11365 1318 11399 1359
rect 11365 1243 11399 1284
rect 11365 1168 11399 1209
rect 11365 1092 11399 1134
rect 11365 1034 11399 1058
rect 13381 1393 13415 1434
rect 13381 1318 13415 1359
rect 13381 1243 13415 1284
rect 13381 1168 13415 1209
rect 13381 1092 13415 1134
rect 13381 1034 13415 1058
<< nsubdiff >>
rect 11365 798 11399 822
rect 11365 714 11399 764
rect 11365 630 11399 680
rect 11365 546 11399 596
rect 13381 798 13415 822
rect 13381 714 13415 764
rect 13381 630 13415 680
rect 13381 546 13415 596
rect 11399 512 11457 522
rect 11365 488 11457 512
rect 13323 512 13381 522
rect 13323 488 13415 512
<< mvpsubdiff >>
rect 9877 36349 14429 36383
rect 9877 35975 9898 36349
rect 10884 36348 14429 36349
rect 10884 36314 10939 36348
rect 10973 36314 11008 36348
rect 11042 36314 11077 36348
rect 11111 36314 11146 36348
rect 11180 36314 11215 36348
rect 11249 36314 11284 36348
rect 11318 36314 11353 36348
rect 11387 36314 11422 36348
rect 11456 36314 11491 36348
rect 11525 36314 11560 36348
rect 11594 36314 11629 36348
rect 11663 36314 11698 36348
rect 11732 36314 11767 36348
rect 11801 36314 11836 36348
rect 11870 36314 11905 36348
rect 11939 36314 11974 36348
rect 12008 36314 12043 36348
rect 12077 36314 12112 36348
rect 12146 36314 12181 36348
rect 12215 36314 12250 36348
rect 12284 36314 12319 36348
rect 12353 36314 12388 36348
rect 12422 36314 12457 36348
rect 10884 36280 12457 36314
rect 10884 36246 10939 36280
rect 10973 36246 11008 36280
rect 11042 36246 11077 36280
rect 11111 36246 11146 36280
rect 11180 36246 11215 36280
rect 11249 36246 11284 36280
rect 11318 36246 11353 36280
rect 11387 36246 11422 36280
rect 11456 36246 11491 36280
rect 11525 36246 11560 36280
rect 11594 36246 11629 36280
rect 11663 36246 11698 36280
rect 11732 36246 11767 36280
rect 11801 36246 11836 36280
rect 11870 36246 11905 36280
rect 11939 36246 11974 36280
rect 12008 36246 12043 36280
rect 12077 36246 12112 36280
rect 12146 36246 12181 36280
rect 12215 36246 12250 36280
rect 12284 36246 12319 36280
rect 12353 36246 12388 36280
rect 12422 36246 12457 36280
rect 10884 36212 12457 36246
rect 10884 36178 10939 36212
rect 10973 36178 11008 36212
rect 11042 36178 11077 36212
rect 11111 36178 11146 36212
rect 11180 36178 11215 36212
rect 11249 36178 11284 36212
rect 11318 36178 11353 36212
rect 11387 36178 11422 36212
rect 11456 36178 11491 36212
rect 11525 36178 11560 36212
rect 11594 36178 11629 36212
rect 11663 36178 11698 36212
rect 11732 36178 11767 36212
rect 11801 36178 11836 36212
rect 11870 36178 11905 36212
rect 11939 36178 11974 36212
rect 12008 36178 12043 36212
rect 12077 36178 12112 36212
rect 12146 36178 12181 36212
rect 12215 36178 12250 36212
rect 12284 36178 12319 36212
rect 12353 36178 12388 36212
rect 12422 36178 12457 36212
rect 10884 36144 12457 36178
rect 10884 36110 10939 36144
rect 10973 36110 11008 36144
rect 11042 36110 11077 36144
rect 11111 36110 11146 36144
rect 11180 36110 11215 36144
rect 11249 36110 11284 36144
rect 11318 36110 11353 36144
rect 11387 36110 11422 36144
rect 11456 36110 11491 36144
rect 11525 36110 11560 36144
rect 11594 36110 11629 36144
rect 11663 36110 11698 36144
rect 11732 36110 11767 36144
rect 11801 36110 11836 36144
rect 11870 36110 11905 36144
rect 11939 36110 11974 36144
rect 12008 36110 12043 36144
rect 12077 36110 12112 36144
rect 12146 36110 12181 36144
rect 12215 36110 12250 36144
rect 12284 36110 12319 36144
rect 12353 36110 12388 36144
rect 12422 36110 12457 36144
rect 10884 36076 12457 36110
rect 10884 36042 10939 36076
rect 10973 36042 11008 36076
rect 11042 36042 11077 36076
rect 11111 36042 11146 36076
rect 11180 36042 11215 36076
rect 11249 36042 11284 36076
rect 11318 36042 11353 36076
rect 11387 36042 11422 36076
rect 11456 36042 11491 36076
rect 11525 36042 11560 36076
rect 11594 36042 11629 36076
rect 11663 36042 11698 36076
rect 11732 36042 11767 36076
rect 11801 36042 11836 36076
rect 11870 36042 11905 36076
rect 11939 36042 11974 36076
rect 12008 36042 12043 36076
rect 12077 36042 12112 36076
rect 12146 36042 12181 36076
rect 12215 36042 12250 36076
rect 12284 36042 12319 36076
rect 12353 36042 12388 36076
rect 12422 36042 12457 36076
rect 10884 36008 12457 36042
rect 10884 35975 10939 36008
rect 9877 35974 10939 35975
rect 10973 35974 11008 36008
rect 11042 35974 11077 36008
rect 11111 35974 11146 36008
rect 11180 35974 11215 36008
rect 11249 35974 11284 36008
rect 11318 35974 11353 36008
rect 11387 35974 11422 36008
rect 11456 35974 11491 36008
rect 11525 35974 11560 36008
rect 11594 35974 11629 36008
rect 11663 35974 11698 36008
rect 11732 35974 11767 36008
rect 11801 35974 11836 36008
rect 11870 35974 11905 36008
rect 11939 35974 11974 36008
rect 12008 35974 12043 36008
rect 12077 35974 12112 36008
rect 12146 35974 12181 36008
rect 12215 35974 12250 36008
rect 12284 35974 12319 36008
rect 12353 35974 12388 36008
rect 12422 35974 12457 36008
rect 9877 35940 12457 35974
rect 9877 35906 9898 35940
rect 9932 35906 9966 35940
rect 10000 35906 10034 35940
rect 10068 35906 10102 35940
rect 10136 35906 10170 35940
rect 10204 35906 10238 35940
rect 10272 35906 10306 35940
rect 10340 35906 10374 35940
rect 10408 35906 10442 35940
rect 10476 35906 10510 35940
rect 10544 35906 10578 35940
rect 10612 35906 10646 35940
rect 10680 35906 10714 35940
rect 10748 35906 10782 35940
rect 10816 35906 10850 35940
rect 10884 35906 10939 35940
rect 10973 35906 11008 35940
rect 11042 35906 11077 35940
rect 11111 35906 11146 35940
rect 11180 35906 11215 35940
rect 11249 35906 11284 35940
rect 11318 35906 11353 35940
rect 11387 35906 11422 35940
rect 11456 35906 11491 35940
rect 11525 35906 11560 35940
rect 11594 35906 11629 35940
rect 11663 35906 11698 35940
rect 11732 35906 11767 35940
rect 11801 35906 11836 35940
rect 11870 35906 11905 35940
rect 11939 35906 11974 35940
rect 12008 35906 12043 35940
rect 12077 35906 12112 35940
rect 12146 35906 12181 35940
rect 12215 35906 12250 35940
rect 12284 35906 12319 35940
rect 12353 35906 12388 35940
rect 12422 35906 12457 35940
rect 9877 35872 12457 35906
rect 9877 35871 10939 35872
rect 9877 35837 9898 35871
rect 9932 35837 9966 35871
rect 10000 35837 10034 35871
rect 10068 35837 10102 35871
rect 10136 35837 10170 35871
rect 10204 35837 10238 35871
rect 10272 35837 10306 35871
rect 10340 35837 10374 35871
rect 10408 35837 10442 35871
rect 10476 35837 10510 35871
rect 10544 35837 10578 35871
rect 10612 35837 10646 35871
rect 10680 35837 10714 35871
rect 10748 35837 10782 35871
rect 10816 35837 10850 35871
rect 10884 35838 10939 35871
rect 10973 35838 11008 35872
rect 11042 35838 11077 35872
rect 11111 35838 11146 35872
rect 11180 35838 11215 35872
rect 11249 35838 11284 35872
rect 11318 35838 11353 35872
rect 11387 35838 11422 35872
rect 11456 35838 11491 35872
rect 11525 35838 11560 35872
rect 11594 35838 11629 35872
rect 11663 35838 11698 35872
rect 11732 35838 11767 35872
rect 11801 35838 11836 35872
rect 11870 35838 11905 35872
rect 11939 35838 11974 35872
rect 12008 35838 12043 35872
rect 12077 35838 12112 35872
rect 12146 35838 12181 35872
rect 12215 35838 12250 35872
rect 12284 35838 12319 35872
rect 12353 35838 12388 35872
rect 12422 35838 12457 35872
rect 10884 35837 12457 35838
rect 9877 35804 12457 35837
rect 9877 35802 10939 35804
rect 9877 35768 9898 35802
rect 9932 35768 9966 35802
rect 10000 35768 10034 35802
rect 10068 35768 10102 35802
rect 10136 35768 10170 35802
rect 10204 35768 10238 35802
rect 10272 35768 10306 35802
rect 10340 35768 10374 35802
rect 10408 35768 10442 35802
rect 10476 35768 10510 35802
rect 10544 35768 10578 35802
rect 10612 35768 10646 35802
rect 10680 35768 10714 35802
rect 10748 35768 10782 35802
rect 10816 35768 10850 35802
rect 10884 35770 10939 35802
rect 10973 35770 11008 35804
rect 11042 35770 11077 35804
rect 11111 35770 11146 35804
rect 11180 35770 11215 35804
rect 11249 35770 11284 35804
rect 11318 35770 11353 35804
rect 11387 35770 11422 35804
rect 11456 35770 11491 35804
rect 11525 35770 11560 35804
rect 11594 35770 11629 35804
rect 11663 35770 11698 35804
rect 11732 35770 11767 35804
rect 11801 35770 11836 35804
rect 11870 35770 11905 35804
rect 11939 35770 11974 35804
rect 12008 35770 12043 35804
rect 12077 35770 12112 35804
rect 12146 35770 12181 35804
rect 12215 35770 12250 35804
rect 12284 35770 12319 35804
rect 12353 35770 12388 35804
rect 12422 35770 12457 35804
rect 14395 35770 14429 36348
rect 10884 35768 14429 35770
rect 9877 35735 14429 35768
rect 9877 35734 10905 35735
rect 13165 35701 14429 35735
rect 13165 35599 13202 35701
rect 14392 35599 14429 35701
rect 13165 35564 14429 35599
rect 13165 35530 13202 35564
rect 13236 35530 13270 35564
rect 13304 35530 13338 35564
rect 13372 35530 13406 35564
rect 13440 35530 13474 35564
rect 13508 35530 13542 35564
rect 13576 35530 13610 35564
rect 13644 35530 13678 35564
rect 13712 35530 13746 35564
rect 13780 35530 13814 35564
rect 13848 35530 13882 35564
rect 13916 35530 13950 35564
rect 13984 35530 14018 35564
rect 14052 35530 14086 35564
rect 14120 35530 14154 35564
rect 14188 35530 14222 35564
rect 14256 35530 14290 35564
rect 14324 35530 14358 35564
rect 14392 35530 14429 35564
rect 13165 35495 14429 35530
rect 13165 35461 13202 35495
rect 13236 35461 13270 35495
rect 13304 35461 13338 35495
rect 13372 35461 13406 35495
rect 13440 35461 13474 35495
rect 13508 35461 13542 35495
rect 13576 35461 13610 35495
rect 13644 35461 13678 35495
rect 13712 35461 13746 35495
rect 13780 35461 13814 35495
rect 13848 35461 13882 35495
rect 13916 35461 13950 35495
rect 13984 35461 14018 35495
rect 14052 35461 14086 35495
rect 14120 35461 14154 35495
rect 14188 35461 14222 35495
rect 14256 35461 14290 35495
rect 14324 35461 14358 35495
rect 14392 35461 14429 35495
rect 13165 35426 14429 35461
rect 13165 35392 13202 35426
rect 13236 35392 13270 35426
rect 13304 35392 13338 35426
rect 13372 35392 13406 35426
rect 13440 35392 13474 35426
rect 13508 35392 13542 35426
rect 13576 35392 13610 35426
rect 13644 35392 13678 35426
rect 13712 35392 13746 35426
rect 13780 35392 13814 35426
rect 13848 35392 13882 35426
rect 13916 35392 13950 35426
rect 13984 35392 14018 35426
rect 14052 35392 14086 35426
rect 14120 35392 14154 35426
rect 14188 35392 14222 35426
rect 14256 35392 14290 35426
rect 14324 35392 14358 35426
rect 14392 35392 14429 35426
rect 13165 35357 14429 35392
rect 13165 35323 13202 35357
rect 13236 35323 13270 35357
rect 13304 35323 13338 35357
rect 13372 35323 13406 35357
rect 13440 35323 13474 35357
rect 13508 35323 13542 35357
rect 13576 35323 13610 35357
rect 13644 35323 13678 35357
rect 13712 35323 13746 35357
rect 13780 35323 13814 35357
rect 13848 35323 13882 35357
rect 13916 35323 13950 35357
rect 13984 35323 14018 35357
rect 14052 35323 14086 35357
rect 14120 35323 14154 35357
rect 14188 35323 14222 35357
rect 14256 35323 14290 35357
rect 14324 35323 14358 35357
rect 14392 35323 14429 35357
rect 13165 35288 14429 35323
rect 13165 35254 13202 35288
rect 13236 35254 13270 35288
rect 13304 35254 13338 35288
rect 13372 35254 13406 35288
rect 13440 35254 13474 35288
rect 13508 35254 13542 35288
rect 13576 35254 13610 35288
rect 13644 35254 13678 35288
rect 13712 35254 13746 35288
rect 13780 35254 13814 35288
rect 13848 35254 13882 35288
rect 13916 35254 13950 35288
rect 13984 35254 14018 35288
rect 14052 35254 14086 35288
rect 14120 35254 14154 35288
rect 14188 35254 14222 35288
rect 14256 35254 14290 35288
rect 14324 35254 14358 35288
rect 14392 35254 14429 35288
rect 13165 35219 14429 35254
rect 13165 35185 13202 35219
rect 13236 35185 13270 35219
rect 13304 35185 13338 35219
rect 13372 35185 13406 35219
rect 13440 35185 13474 35219
rect 13508 35185 13542 35219
rect 13576 35185 13610 35219
rect 13644 35185 13678 35219
rect 13712 35185 13746 35219
rect 13780 35185 13814 35219
rect 13848 35185 13882 35219
rect 13916 35185 13950 35219
rect 13984 35185 14018 35219
rect 14052 35185 14086 35219
rect 14120 35185 14154 35219
rect 14188 35185 14222 35219
rect 14256 35185 14290 35219
rect 14324 35185 14358 35219
rect 14392 35185 14429 35219
rect 13165 35150 14429 35185
rect 13165 35116 13202 35150
rect 13236 35116 13270 35150
rect 13304 35116 13338 35150
rect 13372 35116 13406 35150
rect 13440 35116 13474 35150
rect 13508 35116 13542 35150
rect 13576 35116 13610 35150
rect 13644 35116 13678 35150
rect 13712 35116 13746 35150
rect 13780 35116 13814 35150
rect 13848 35116 13882 35150
rect 13916 35116 13950 35150
rect 13984 35116 14018 35150
rect 14052 35116 14086 35150
rect 14120 35116 14154 35150
rect 14188 35116 14222 35150
rect 14256 35116 14290 35150
rect 14324 35116 14358 35150
rect 14392 35116 14429 35150
rect 13165 35081 14429 35116
rect 13165 35047 13202 35081
rect 13236 35047 13270 35081
rect 13304 35047 13338 35081
rect 13372 35047 13406 35081
rect 13440 35047 13474 35081
rect 13508 35047 13542 35081
rect 13576 35047 13610 35081
rect 13644 35047 13678 35081
rect 13712 35047 13746 35081
rect 13780 35047 13814 35081
rect 13848 35047 13882 35081
rect 13916 35047 13950 35081
rect 13984 35047 14018 35081
rect 14052 35047 14086 35081
rect 14120 35047 14154 35081
rect 14188 35047 14222 35081
rect 14256 35047 14290 35081
rect 14324 35047 14358 35081
rect 14392 35047 14429 35081
rect 13165 35012 14429 35047
rect 13165 34978 13202 35012
rect 13236 34978 13270 35012
rect 13304 34978 13338 35012
rect 13372 34978 13406 35012
rect 13440 34978 13474 35012
rect 13508 34978 13542 35012
rect 13576 34978 13610 35012
rect 13644 34978 13678 35012
rect 13712 34978 13746 35012
rect 13780 34978 13814 35012
rect 13848 34978 13882 35012
rect 13916 34978 13950 35012
rect 13984 34978 14018 35012
rect 14052 34978 14086 35012
rect 14120 34978 14154 35012
rect 14188 34978 14222 35012
rect 14256 34978 14290 35012
rect 14324 34978 14358 35012
rect 14392 34978 14429 35012
rect 13165 34943 14429 34978
rect 13165 34909 13202 34943
rect 13236 34909 13270 34943
rect 13304 34909 13338 34943
rect 13372 34909 13406 34943
rect 13440 34909 13474 34943
rect 13508 34909 13542 34943
rect 13576 34909 13610 34943
rect 13644 34909 13678 34943
rect 13712 34909 13746 34943
rect 13780 34909 13814 34943
rect 13848 34909 13882 34943
rect 13916 34909 13950 34943
rect 13984 34909 14018 34943
rect 14052 34909 14086 34943
rect 14120 34909 14154 34943
rect 14188 34909 14222 34943
rect 14256 34909 14290 34943
rect 14324 34909 14358 34943
rect 14392 34909 14429 34943
rect 13165 34874 14429 34909
rect 13165 34840 13202 34874
rect 13236 34840 13270 34874
rect 13304 34840 13338 34874
rect 13372 34840 13406 34874
rect 13440 34840 13474 34874
rect 13508 34840 13542 34874
rect 13576 34840 13610 34874
rect 13644 34840 13678 34874
rect 13712 34840 13746 34874
rect 13780 34840 13814 34874
rect 13848 34840 13882 34874
rect 13916 34840 13950 34874
rect 13984 34840 14018 34874
rect 14052 34840 14086 34874
rect 14120 34840 14154 34874
rect 14188 34840 14222 34874
rect 14256 34840 14290 34874
rect 14324 34840 14358 34874
rect 14392 34840 14429 34874
rect 13165 34805 14429 34840
rect 13165 34771 13202 34805
rect 13236 34771 13270 34805
rect 13304 34771 13338 34805
rect 13372 34771 13406 34805
rect 13440 34771 13474 34805
rect 13508 34771 13542 34805
rect 13576 34771 13610 34805
rect 13644 34771 13678 34805
rect 13712 34771 13746 34805
rect 13780 34771 13814 34805
rect 13848 34771 13882 34805
rect 13916 34771 13950 34805
rect 13984 34771 14018 34805
rect 14052 34771 14086 34805
rect 14120 34771 14154 34805
rect 14188 34771 14222 34805
rect 14256 34771 14290 34805
rect 14324 34771 14358 34805
rect 14392 34771 14429 34805
rect 13165 34736 14429 34771
rect 13165 34702 13202 34736
rect 13236 34702 13270 34736
rect 13304 34702 13338 34736
rect 13372 34702 13406 34736
rect 13440 34702 13474 34736
rect 13508 34702 13542 34736
rect 13576 34702 13610 34736
rect 13644 34702 13678 34736
rect 13712 34702 13746 34736
rect 13780 34702 13814 34736
rect 13848 34702 13882 34736
rect 13916 34702 13950 34736
rect 13984 34702 14018 34736
rect 14052 34702 14086 34736
rect 14120 34702 14154 34736
rect 14188 34702 14222 34736
rect 14256 34702 14290 34736
rect 14324 34702 14358 34736
rect 14392 34702 14429 34736
rect 13165 34667 14429 34702
rect 13165 34633 13202 34667
rect 13236 34633 13270 34667
rect 13304 34633 13338 34667
rect 13372 34633 13406 34667
rect 13440 34633 13474 34667
rect 13508 34633 13542 34667
rect 13576 34633 13610 34667
rect 13644 34633 13678 34667
rect 13712 34633 13746 34667
rect 13780 34633 13814 34667
rect 13848 34633 13882 34667
rect 13916 34633 13950 34667
rect 13984 34633 14018 34667
rect 14052 34633 14086 34667
rect 14120 34633 14154 34667
rect 14188 34633 14222 34667
rect 14256 34633 14290 34667
rect 14324 34633 14358 34667
rect 14392 34633 14429 34667
rect 13165 34598 14429 34633
rect 13165 34564 13202 34598
rect 13236 34564 13270 34598
rect 13304 34564 13338 34598
rect 13372 34564 13406 34598
rect 13440 34564 13474 34598
rect 13508 34564 13542 34598
rect 13576 34564 13610 34598
rect 13644 34564 13678 34598
rect 13712 34564 13746 34598
rect 13780 34564 13814 34598
rect 13848 34564 13882 34598
rect 13916 34564 13950 34598
rect 13984 34564 14018 34598
rect 14052 34564 14086 34598
rect 14120 34564 14154 34598
rect 14188 34564 14222 34598
rect 14256 34564 14290 34598
rect 14324 34564 14358 34598
rect 14392 34564 14429 34598
rect 13165 34529 14429 34564
rect 13165 34495 13202 34529
rect 13236 34495 13270 34529
rect 13304 34495 13338 34529
rect 13372 34495 13406 34529
rect 13440 34495 13474 34529
rect 13508 34495 13542 34529
rect 13576 34495 13610 34529
rect 13644 34495 13678 34529
rect 13712 34495 13746 34529
rect 13780 34495 13814 34529
rect 13848 34495 13882 34529
rect 13916 34495 13950 34529
rect 13984 34495 14018 34529
rect 14052 34495 14086 34529
rect 14120 34495 14154 34529
rect 14188 34495 14222 34529
rect 14256 34495 14290 34529
rect 14324 34495 14358 34529
rect 14392 34495 14429 34529
rect 13165 34460 14429 34495
rect 13165 34426 13202 34460
rect 13236 34426 13270 34460
rect 13304 34426 13338 34460
rect 13372 34426 13406 34460
rect 13440 34426 13474 34460
rect 13508 34426 13542 34460
rect 13576 34426 13610 34460
rect 13644 34426 13678 34460
rect 13712 34426 13746 34460
rect 13780 34426 13814 34460
rect 13848 34426 13882 34460
rect 13916 34426 13950 34460
rect 13984 34426 14018 34460
rect 14052 34426 14086 34460
rect 14120 34426 14154 34460
rect 14188 34426 14222 34460
rect 14256 34426 14290 34460
rect 14324 34426 14358 34460
rect 14392 34426 14429 34460
rect 13165 34391 14429 34426
rect 13165 34357 13202 34391
rect 13236 34357 13270 34391
rect 13304 34357 13338 34391
rect 13372 34357 13406 34391
rect 13440 34357 13474 34391
rect 13508 34357 13542 34391
rect 13576 34357 13610 34391
rect 13644 34357 13678 34391
rect 13712 34357 13746 34391
rect 13780 34357 13814 34391
rect 13848 34357 13882 34391
rect 13916 34357 13950 34391
rect 13984 34357 14018 34391
rect 14052 34357 14086 34391
rect 14120 34357 14154 34391
rect 14188 34357 14222 34391
rect 14256 34357 14290 34391
rect 14324 34357 14358 34391
rect 14392 34357 14429 34391
rect 13165 34322 14429 34357
rect 13165 34288 13202 34322
rect 13236 34288 13270 34322
rect 13304 34288 13338 34322
rect 13372 34288 13406 34322
rect 13440 34288 13474 34322
rect 13508 34288 13542 34322
rect 13576 34288 13610 34322
rect 13644 34288 13678 34322
rect 13712 34288 13746 34322
rect 13780 34288 13814 34322
rect 13848 34288 13882 34322
rect 13916 34288 13950 34322
rect 13984 34288 14018 34322
rect 14052 34288 14086 34322
rect 14120 34288 14154 34322
rect 14188 34288 14222 34322
rect 14256 34288 14290 34322
rect 14324 34288 14358 34322
rect 14392 34288 14429 34322
rect 13165 34253 14429 34288
rect 13165 34219 13202 34253
rect 13236 34219 13270 34253
rect 13304 34219 13338 34253
rect 13372 34219 13406 34253
rect 13440 34219 13474 34253
rect 13508 34219 13542 34253
rect 13576 34219 13610 34253
rect 13644 34219 13678 34253
rect 13712 34219 13746 34253
rect 13780 34219 13814 34253
rect 13848 34219 13882 34253
rect 13916 34219 13950 34253
rect 13984 34219 14018 34253
rect 14052 34219 14086 34253
rect 14120 34219 14154 34253
rect 14188 34219 14222 34253
rect 14256 34219 14290 34253
rect 14324 34219 14358 34253
rect 14392 34219 14429 34253
rect 13165 34184 14429 34219
rect 13165 34150 13202 34184
rect 13236 34150 13270 34184
rect 13304 34150 13338 34184
rect 13372 34150 13406 34184
rect 13440 34150 13474 34184
rect 13508 34150 13542 34184
rect 13576 34150 13610 34184
rect 13644 34150 13678 34184
rect 13712 34150 13746 34184
rect 13780 34150 13814 34184
rect 13848 34150 13882 34184
rect 13916 34150 13950 34184
rect 13984 34150 14018 34184
rect 14052 34150 14086 34184
rect 14120 34150 14154 34184
rect 14188 34150 14222 34184
rect 14256 34150 14290 34184
rect 14324 34150 14358 34184
rect 14392 34150 14429 34184
rect 13165 34115 14429 34150
rect 13165 34081 13202 34115
rect 13236 34081 13270 34115
rect 13304 34081 13338 34115
rect 13372 34081 13406 34115
rect 13440 34081 13474 34115
rect 13508 34081 13542 34115
rect 13576 34081 13610 34115
rect 13644 34081 13678 34115
rect 13712 34081 13746 34115
rect 13780 34081 13814 34115
rect 13848 34081 13882 34115
rect 13916 34081 13950 34115
rect 13984 34081 14018 34115
rect 14052 34081 14086 34115
rect 14120 34081 14154 34115
rect 14188 34081 14222 34115
rect 14256 34081 14290 34115
rect 14324 34081 14358 34115
rect 14392 34081 14429 34115
rect 13165 34046 14429 34081
rect 13165 34012 13202 34046
rect 13236 34012 13270 34046
rect 13304 34012 13338 34046
rect 13372 34012 13406 34046
rect 13440 34012 13474 34046
rect 13508 34012 13542 34046
rect 13576 34012 13610 34046
rect 13644 34012 13678 34046
rect 13712 34012 13746 34046
rect 13780 34012 13814 34046
rect 13848 34012 13882 34046
rect 13916 34012 13950 34046
rect 13984 34012 14018 34046
rect 14052 34012 14086 34046
rect 14120 34012 14154 34046
rect 14188 34012 14222 34046
rect 14256 34012 14290 34046
rect 14324 34012 14358 34046
rect 14392 34012 14429 34046
rect 13165 33977 14429 34012
rect 13165 33943 13202 33977
rect 13236 33943 13270 33977
rect 13304 33943 13338 33977
rect 13372 33943 13406 33977
rect 13440 33943 13474 33977
rect 13508 33943 13542 33977
rect 13576 33943 13610 33977
rect 13644 33943 13678 33977
rect 13712 33943 13746 33977
rect 13780 33943 13814 33977
rect 13848 33943 13882 33977
rect 13916 33943 13950 33977
rect 13984 33943 14018 33977
rect 14052 33943 14086 33977
rect 14120 33943 14154 33977
rect 14188 33943 14222 33977
rect 14256 33943 14290 33977
rect 14324 33943 14358 33977
rect 14392 33943 14429 33977
rect 13165 33908 14429 33943
rect 13165 33874 13202 33908
rect 13236 33874 13270 33908
rect 13304 33874 13338 33908
rect 13372 33874 13406 33908
rect 13440 33874 13474 33908
rect 13508 33874 13542 33908
rect 13576 33874 13610 33908
rect 13644 33874 13678 33908
rect 13712 33874 13746 33908
rect 13780 33874 13814 33908
rect 13848 33874 13882 33908
rect 13916 33874 13950 33908
rect 13984 33874 14018 33908
rect 14052 33874 14086 33908
rect 14120 33874 14154 33908
rect 14188 33874 14222 33908
rect 14256 33874 14290 33908
rect 14324 33874 14358 33908
rect 14392 33874 14429 33908
rect 13165 33839 14429 33874
rect 13165 33805 13202 33839
rect 13236 33805 13270 33839
rect 13304 33805 13338 33839
rect 13372 33805 13406 33839
rect 13440 33805 13474 33839
rect 13508 33805 13542 33839
rect 13576 33805 13610 33839
rect 13644 33805 13678 33839
rect 13712 33805 13746 33839
rect 13780 33805 13814 33839
rect 13848 33805 13882 33839
rect 13916 33805 13950 33839
rect 13984 33805 14018 33839
rect 14052 33805 14086 33839
rect 14120 33805 14154 33839
rect 14188 33805 14222 33839
rect 14256 33805 14290 33839
rect 14324 33805 14358 33839
rect 14392 33805 14429 33839
rect 13165 33770 14429 33805
rect 13165 33736 13202 33770
rect 13236 33736 13270 33770
rect 13304 33736 13338 33770
rect 13372 33736 13406 33770
rect 13440 33736 13474 33770
rect 13508 33736 13542 33770
rect 13576 33736 13610 33770
rect 13644 33736 13678 33770
rect 13712 33736 13746 33770
rect 13780 33736 13814 33770
rect 13848 33736 13882 33770
rect 13916 33736 13950 33770
rect 13984 33736 14018 33770
rect 14052 33736 14086 33770
rect 14120 33736 14154 33770
rect 14188 33736 14222 33770
rect 14256 33736 14290 33770
rect 14324 33736 14358 33770
rect 14392 33736 14429 33770
rect 13165 33701 14429 33736
rect 13165 33667 13202 33701
rect 13236 33667 13270 33701
rect 13304 33667 13338 33701
rect 13372 33667 13406 33701
rect 13440 33667 13474 33701
rect 13508 33667 13542 33701
rect 13576 33667 13610 33701
rect 13644 33667 13678 33701
rect 13712 33667 13746 33701
rect 13780 33667 13814 33701
rect 13848 33667 13882 33701
rect 13916 33667 13950 33701
rect 13984 33667 14018 33701
rect 14052 33667 14086 33701
rect 14120 33667 14154 33701
rect 14188 33667 14222 33701
rect 14256 33667 14290 33701
rect 14324 33667 14358 33701
rect 14392 33667 14429 33701
rect 13165 33632 14429 33667
rect 13165 33598 13202 33632
rect 13236 33598 13270 33632
rect 13304 33598 13338 33632
rect 13372 33598 13406 33632
rect 13440 33598 13474 33632
rect 13508 33598 13542 33632
rect 13576 33598 13610 33632
rect 13644 33598 13678 33632
rect 13712 33598 13746 33632
rect 13780 33598 13814 33632
rect 13848 33598 13882 33632
rect 13916 33598 13950 33632
rect 13984 33598 14018 33632
rect 14052 33598 14086 33632
rect 14120 33598 14154 33632
rect 14188 33598 14222 33632
rect 14256 33598 14290 33632
rect 14324 33598 14358 33632
rect 14392 33598 14429 33632
rect 13165 33563 14429 33598
rect 13165 33529 13202 33563
rect 13236 33529 13270 33563
rect 13304 33529 13338 33563
rect 13372 33529 13406 33563
rect 13440 33529 13474 33563
rect 13508 33529 13542 33563
rect 13576 33529 13610 33563
rect 13644 33529 13678 33563
rect 13712 33529 13746 33563
rect 13780 33529 13814 33563
rect 13848 33529 13882 33563
rect 13916 33529 13950 33563
rect 13984 33529 14018 33563
rect 14052 33529 14086 33563
rect 14120 33529 14154 33563
rect 14188 33529 14222 33563
rect 14256 33529 14290 33563
rect 14324 33529 14358 33563
rect 14392 33529 14429 33563
rect 13165 33494 14429 33529
rect 13165 33460 13202 33494
rect 13236 33460 13270 33494
rect 13304 33460 13338 33494
rect 13372 33460 13406 33494
rect 13440 33460 13474 33494
rect 13508 33460 13542 33494
rect 13576 33460 13610 33494
rect 13644 33460 13678 33494
rect 13712 33460 13746 33494
rect 13780 33460 13814 33494
rect 13848 33460 13882 33494
rect 13916 33460 13950 33494
rect 13984 33460 14018 33494
rect 14052 33460 14086 33494
rect 14120 33460 14154 33494
rect 14188 33460 14222 33494
rect 14256 33460 14290 33494
rect 14324 33460 14358 33494
rect 14392 33460 14429 33494
rect 13165 33425 14429 33460
rect 13165 33391 13202 33425
rect 13236 33391 13270 33425
rect 13304 33391 13338 33425
rect 13372 33391 13406 33425
rect 13440 33391 13474 33425
rect 13508 33391 13542 33425
rect 13576 33391 13610 33425
rect 13644 33391 13678 33425
rect 13712 33391 13746 33425
rect 13780 33391 13814 33425
rect 13848 33391 13882 33425
rect 13916 33391 13950 33425
rect 13984 33391 14018 33425
rect 14052 33391 14086 33425
rect 14120 33391 14154 33425
rect 14188 33391 14222 33425
rect 14256 33391 14290 33425
rect 14324 33391 14358 33425
rect 14392 33391 14429 33425
rect 13165 33356 14429 33391
rect 13165 33322 13202 33356
rect 13236 33322 13270 33356
rect 13304 33322 13338 33356
rect 13372 33322 13406 33356
rect 13440 33322 13474 33356
rect 13508 33322 13542 33356
rect 13576 33322 13610 33356
rect 13644 33322 13678 33356
rect 13712 33322 13746 33356
rect 13780 33322 13814 33356
rect 13848 33322 13882 33356
rect 13916 33322 13950 33356
rect 13984 33322 14018 33356
rect 14052 33322 14086 33356
rect 14120 33322 14154 33356
rect 14188 33322 14222 33356
rect 14256 33322 14290 33356
rect 14324 33322 14358 33356
rect 14392 33322 14429 33356
rect 13165 33287 14429 33322
rect 13165 33253 13202 33287
rect 13236 33253 13270 33287
rect 13304 33253 13338 33287
rect 13372 33253 13406 33287
rect 13440 33253 13474 33287
rect 13508 33253 13542 33287
rect 13576 33253 13610 33287
rect 13644 33253 13678 33287
rect 13712 33253 13746 33287
rect 13780 33253 13814 33287
rect 13848 33253 13882 33287
rect 13916 33253 13950 33287
rect 13984 33253 14018 33287
rect 14052 33253 14086 33287
rect 14120 33253 14154 33287
rect 14188 33253 14222 33287
rect 14256 33253 14290 33287
rect 14324 33253 14358 33287
rect 14392 33253 14429 33287
rect 13165 33218 14429 33253
rect 13165 33184 13202 33218
rect 13236 33184 13270 33218
rect 13304 33184 13338 33218
rect 13372 33184 13406 33218
rect 13440 33184 13474 33218
rect 13508 33184 13542 33218
rect 13576 33184 13610 33218
rect 13644 33184 13678 33218
rect 13712 33184 13746 33218
rect 13780 33184 13814 33218
rect 13848 33184 13882 33218
rect 13916 33184 13950 33218
rect 13984 33184 14018 33218
rect 14052 33184 14086 33218
rect 14120 33184 14154 33218
rect 14188 33184 14222 33218
rect 14256 33184 14290 33218
rect 14324 33184 14358 33218
rect 14392 33184 14429 33218
rect 13165 33149 14429 33184
rect 13165 33115 13202 33149
rect 13236 33115 13270 33149
rect 13304 33115 13338 33149
rect 13372 33115 13406 33149
rect 13440 33115 13474 33149
rect 13508 33115 13542 33149
rect 13576 33115 13610 33149
rect 13644 33115 13678 33149
rect 13712 33115 13746 33149
rect 13780 33115 13814 33149
rect 13848 33115 13882 33149
rect 13916 33115 13950 33149
rect 13984 33115 14018 33149
rect 14052 33115 14086 33149
rect 14120 33115 14154 33149
rect 14188 33115 14222 33149
rect 14256 33115 14290 33149
rect 14324 33115 14358 33149
rect 14392 33115 14429 33149
rect 13165 33080 14429 33115
rect 13165 33046 13202 33080
rect 13236 33046 13270 33080
rect 13304 33046 13338 33080
rect 13372 33046 13406 33080
rect 13440 33046 13474 33080
rect 13508 33046 13542 33080
rect 13576 33046 13610 33080
rect 13644 33046 13678 33080
rect 13712 33046 13746 33080
rect 13780 33046 13814 33080
rect 13848 33046 13882 33080
rect 13916 33046 13950 33080
rect 13984 33046 14018 33080
rect 14052 33046 14086 33080
rect 14120 33046 14154 33080
rect 14188 33046 14222 33080
rect 14256 33046 14290 33080
rect 14324 33046 14358 33080
rect 14392 33046 14429 33080
rect 13165 33011 14429 33046
rect 13165 32977 13202 33011
rect 13236 32977 13270 33011
rect 13304 32977 13338 33011
rect 13372 32977 13406 33011
rect 13440 32977 13474 33011
rect 13508 32977 13542 33011
rect 13576 32977 13610 33011
rect 13644 32977 13678 33011
rect 13712 32977 13746 33011
rect 13780 32977 13814 33011
rect 13848 32977 13882 33011
rect 13916 32977 13950 33011
rect 13984 32977 14018 33011
rect 14052 32977 14086 33011
rect 14120 32977 14154 33011
rect 14188 32977 14222 33011
rect 14256 32977 14290 33011
rect 14324 32977 14358 33011
rect 14392 32977 14429 33011
rect 13165 32942 14429 32977
rect 13165 32908 13202 32942
rect 13236 32908 13270 32942
rect 13304 32908 13338 32942
rect 13372 32908 13406 32942
rect 13440 32908 13474 32942
rect 13508 32908 13542 32942
rect 13576 32908 13610 32942
rect 13644 32908 13678 32942
rect 13712 32908 13746 32942
rect 13780 32908 13814 32942
rect 13848 32908 13882 32942
rect 13916 32908 13950 32942
rect 13984 32908 14018 32942
rect 14052 32908 14086 32942
rect 14120 32908 14154 32942
rect 14188 32908 14222 32942
rect 14256 32908 14290 32942
rect 14324 32908 14358 32942
rect 14392 32908 14429 32942
rect 13165 32873 14429 32908
rect 13165 32839 13202 32873
rect 13236 32839 13270 32873
rect 13304 32839 13338 32873
rect 13372 32839 13406 32873
rect 13440 32839 13474 32873
rect 13508 32839 13542 32873
rect 13576 32839 13610 32873
rect 13644 32839 13678 32873
rect 13712 32839 13746 32873
rect 13780 32839 13814 32873
rect 13848 32839 13882 32873
rect 13916 32839 13950 32873
rect 13984 32839 14018 32873
rect 14052 32839 14086 32873
rect 14120 32839 14154 32873
rect 14188 32839 14222 32873
rect 14256 32839 14290 32873
rect 14324 32839 14358 32873
rect 14392 32839 14429 32873
rect 13165 32804 14429 32839
rect 13165 32770 13202 32804
rect 13236 32770 13270 32804
rect 13304 32770 13338 32804
rect 13372 32770 13406 32804
rect 13440 32770 13474 32804
rect 13508 32770 13542 32804
rect 13576 32770 13610 32804
rect 13644 32770 13678 32804
rect 13712 32770 13746 32804
rect 13780 32770 13814 32804
rect 13848 32770 13882 32804
rect 13916 32770 13950 32804
rect 13984 32770 14018 32804
rect 14052 32770 14086 32804
rect 14120 32770 14154 32804
rect 14188 32770 14222 32804
rect 14256 32770 14290 32804
rect 14324 32770 14358 32804
rect 14392 32770 14429 32804
rect 13165 32735 14429 32770
rect 13165 32701 13202 32735
rect 13236 32701 13270 32735
rect 13304 32701 13338 32735
rect 13372 32701 13406 32735
rect 13440 32701 13474 32735
rect 13508 32701 13542 32735
rect 13576 32701 13610 32735
rect 13644 32701 13678 32735
rect 13712 32701 13746 32735
rect 13780 32701 13814 32735
rect 13848 32701 13882 32735
rect 13916 32701 13950 32735
rect 13984 32701 14018 32735
rect 14052 32701 14086 32735
rect 14120 32701 14154 32735
rect 14188 32701 14222 32735
rect 14256 32701 14290 32735
rect 14324 32701 14358 32735
rect 14392 32701 14429 32735
rect 13165 32666 14429 32701
rect 13165 32632 13202 32666
rect 13236 32632 13270 32666
rect 13304 32632 13338 32666
rect 13372 32632 13406 32666
rect 13440 32632 13474 32666
rect 13508 32632 13542 32666
rect 13576 32632 13610 32666
rect 13644 32632 13678 32666
rect 13712 32632 13746 32666
rect 13780 32632 13814 32666
rect 13848 32632 13882 32666
rect 13916 32632 13950 32666
rect 13984 32632 14018 32666
rect 14052 32632 14086 32666
rect 14120 32632 14154 32666
rect 14188 32632 14222 32666
rect 14256 32632 14290 32666
rect 14324 32632 14358 32666
rect 14392 32632 14429 32666
rect 13165 32597 14429 32632
rect 13165 32563 13202 32597
rect 13236 32563 13270 32597
rect 13304 32563 13338 32597
rect 13372 32563 13406 32597
rect 13440 32563 13474 32597
rect 13508 32563 13542 32597
rect 13576 32563 13610 32597
rect 13644 32563 13678 32597
rect 13712 32563 13746 32597
rect 13780 32563 13814 32597
rect 13848 32563 13882 32597
rect 13916 32563 13950 32597
rect 13984 32563 14018 32597
rect 14052 32563 14086 32597
rect 14120 32563 14154 32597
rect 14188 32563 14222 32597
rect 14256 32563 14290 32597
rect 14324 32563 14358 32597
rect 14392 32563 14429 32597
rect 13165 32528 14429 32563
rect 13165 32494 13202 32528
rect 13236 32494 13270 32528
rect 13304 32494 13338 32528
rect 13372 32494 13406 32528
rect 13440 32494 13474 32528
rect 13508 32494 13542 32528
rect 13576 32494 13610 32528
rect 13644 32494 13678 32528
rect 13712 32494 13746 32528
rect 13780 32494 13814 32528
rect 13848 32494 13882 32528
rect 13916 32494 13950 32528
rect 13984 32494 14018 32528
rect 14052 32494 14086 32528
rect 14120 32494 14154 32528
rect 14188 32494 14222 32528
rect 14256 32494 14290 32528
rect 14324 32494 14358 32528
rect 14392 32494 14429 32528
rect 13165 32459 14429 32494
rect 13165 32425 13202 32459
rect 13236 32425 13270 32459
rect 13304 32425 13338 32459
rect 13372 32425 13406 32459
rect 13440 32425 13474 32459
rect 13508 32425 13542 32459
rect 13576 32425 13610 32459
rect 13644 32425 13678 32459
rect 13712 32425 13746 32459
rect 13780 32425 13814 32459
rect 13848 32425 13882 32459
rect 13916 32425 13950 32459
rect 13984 32425 14018 32459
rect 14052 32425 14086 32459
rect 14120 32425 14154 32459
rect 14188 32425 14222 32459
rect 14256 32425 14290 32459
rect 14324 32425 14358 32459
rect 14392 32425 14429 32459
rect 13165 32390 14429 32425
rect 13165 32356 13202 32390
rect 13236 32356 13270 32390
rect 13304 32356 13338 32390
rect 13372 32356 13406 32390
rect 13440 32356 13474 32390
rect 13508 32356 13542 32390
rect 13576 32356 13610 32390
rect 13644 32356 13678 32390
rect 13712 32356 13746 32390
rect 13780 32356 13814 32390
rect 13848 32356 13882 32390
rect 13916 32356 13950 32390
rect 13984 32356 14018 32390
rect 14052 32356 14086 32390
rect 14120 32356 14154 32390
rect 14188 32356 14222 32390
rect 14256 32356 14290 32390
rect 14324 32356 14358 32390
rect 14392 32356 14429 32390
rect 13165 32321 14429 32356
rect 13165 32287 13202 32321
rect 13236 32287 13270 32321
rect 13304 32287 13338 32321
rect 13372 32287 13406 32321
rect 13440 32287 13474 32321
rect 13508 32287 13542 32321
rect 13576 32287 13610 32321
rect 13644 32287 13678 32321
rect 13712 32287 13746 32321
rect 13780 32287 13814 32321
rect 13848 32287 13882 32321
rect 13916 32287 13950 32321
rect 13984 32287 14018 32321
rect 14052 32287 14086 32321
rect 14120 32287 14154 32321
rect 14188 32287 14222 32321
rect 14256 32287 14290 32321
rect 14324 32287 14358 32321
rect 14392 32287 14429 32321
rect 13165 32252 14429 32287
rect 13165 32218 13202 32252
rect 13236 32218 13270 32252
rect 13304 32218 13338 32252
rect 13372 32218 13406 32252
rect 13440 32218 13474 32252
rect 13508 32218 13542 32252
rect 13576 32218 13610 32252
rect 13644 32218 13678 32252
rect 13712 32218 13746 32252
rect 13780 32218 13814 32252
rect 13848 32218 13882 32252
rect 13916 32218 13950 32252
rect 13984 32218 14018 32252
rect 14052 32218 14086 32252
rect 14120 32218 14154 32252
rect 14188 32218 14222 32252
rect 14256 32218 14290 32252
rect 14324 32218 14358 32252
rect 14392 32218 14429 32252
rect 13165 32183 14429 32218
rect 13165 32149 13202 32183
rect 13236 32149 13270 32183
rect 13304 32149 13338 32183
rect 13372 32149 13406 32183
rect 13440 32149 13474 32183
rect 13508 32149 13542 32183
rect 13576 32149 13610 32183
rect 13644 32149 13678 32183
rect 13712 32149 13746 32183
rect 13780 32149 13814 32183
rect 13848 32149 13882 32183
rect 13916 32149 13950 32183
rect 13984 32149 14018 32183
rect 14052 32149 14086 32183
rect 14120 32149 14154 32183
rect 14188 32149 14222 32183
rect 14256 32149 14290 32183
rect 14324 32149 14358 32183
rect 14392 32149 14429 32183
rect 13165 32114 14429 32149
rect 13165 32080 13202 32114
rect 13236 32080 13270 32114
rect 13304 32080 13338 32114
rect 13372 32080 13406 32114
rect 13440 32080 13474 32114
rect 13508 32080 13542 32114
rect 13576 32080 13610 32114
rect 13644 32080 13678 32114
rect 13712 32080 13746 32114
rect 13780 32080 13814 32114
rect 13848 32080 13882 32114
rect 13916 32080 13950 32114
rect 13984 32080 14018 32114
rect 14052 32080 14086 32114
rect 14120 32080 14154 32114
rect 14188 32080 14222 32114
rect 14256 32080 14290 32114
rect 14324 32080 14358 32114
rect 14392 32080 14429 32114
rect 13165 32045 14429 32080
rect 13165 32011 13202 32045
rect 13236 32011 13270 32045
rect 13304 32011 13338 32045
rect 13372 32011 13406 32045
rect 13440 32011 13474 32045
rect 13508 32011 13542 32045
rect 13576 32011 13610 32045
rect 13644 32011 13678 32045
rect 13712 32011 13746 32045
rect 13780 32011 13814 32045
rect 13848 32011 13882 32045
rect 13916 32011 13950 32045
rect 13984 32011 14018 32045
rect 14052 32011 14086 32045
rect 14120 32011 14154 32045
rect 14188 32011 14222 32045
rect 14256 32011 14290 32045
rect 14324 32011 14358 32045
rect 14392 32011 14429 32045
rect 13165 31976 14429 32011
rect 13165 31942 13202 31976
rect 13236 31942 13270 31976
rect 13304 31942 13338 31976
rect 13372 31942 13406 31976
rect 13440 31942 13474 31976
rect 13508 31942 13542 31976
rect 13576 31942 13610 31976
rect 13644 31942 13678 31976
rect 13712 31942 13746 31976
rect 13780 31942 13814 31976
rect 13848 31942 13882 31976
rect 13916 31942 13950 31976
rect 13984 31942 14018 31976
rect 14052 31942 14086 31976
rect 14120 31942 14154 31976
rect 14188 31942 14222 31976
rect 14256 31942 14290 31976
rect 14324 31942 14358 31976
rect 14392 31942 14429 31976
rect 13165 31907 14429 31942
rect 13165 31873 13202 31907
rect 13236 31873 13270 31907
rect 13304 31873 13338 31907
rect 13372 31873 13406 31907
rect 13440 31873 13474 31907
rect 13508 31873 13542 31907
rect 13576 31873 13610 31907
rect 13644 31873 13678 31907
rect 13712 31873 13746 31907
rect 13780 31873 13814 31907
rect 13848 31873 13882 31907
rect 13916 31873 13950 31907
rect 13984 31873 14018 31907
rect 14052 31873 14086 31907
rect 14120 31873 14154 31907
rect 14188 31873 14222 31907
rect 14256 31873 14290 31907
rect 14324 31873 14358 31907
rect 14392 31873 14429 31907
rect 13165 31838 14429 31873
rect 13165 31804 13202 31838
rect 13236 31804 13270 31838
rect 13304 31804 13338 31838
rect 13372 31804 13406 31838
rect 13440 31804 13474 31838
rect 13508 31804 13542 31838
rect 13576 31804 13610 31838
rect 13644 31804 13678 31838
rect 13712 31804 13746 31838
rect 13780 31804 13814 31838
rect 13848 31804 13882 31838
rect 13916 31804 13950 31838
rect 13984 31804 14018 31838
rect 14052 31804 14086 31838
rect 14120 31804 14154 31838
rect 14188 31804 14222 31838
rect 14256 31804 14290 31838
rect 14324 31804 14358 31838
rect 14392 31804 14429 31838
rect 13165 31769 14429 31804
rect 13165 31735 13202 31769
rect 13236 31735 13270 31769
rect 13304 31735 13338 31769
rect 13372 31735 13406 31769
rect 13440 31735 13474 31769
rect 13508 31735 13542 31769
rect 13576 31735 13610 31769
rect 13644 31735 13678 31769
rect 13712 31735 13746 31769
rect 13780 31735 13814 31769
rect 13848 31735 13882 31769
rect 13916 31735 13950 31769
rect 13984 31735 14018 31769
rect 14052 31735 14086 31769
rect 14120 31735 14154 31769
rect 14188 31735 14222 31769
rect 14256 31735 14290 31769
rect 14324 31735 14358 31769
rect 14392 31735 14429 31769
rect 13165 31700 14429 31735
rect 13165 31666 13202 31700
rect 13236 31666 13270 31700
rect 13304 31666 13338 31700
rect 13372 31666 13406 31700
rect 13440 31666 13474 31700
rect 13508 31666 13542 31700
rect 13576 31666 13610 31700
rect 13644 31666 13678 31700
rect 13712 31666 13746 31700
rect 13780 31666 13814 31700
rect 13848 31666 13882 31700
rect 13916 31666 13950 31700
rect 13984 31666 14018 31700
rect 14052 31666 14086 31700
rect 14120 31666 14154 31700
rect 14188 31666 14222 31700
rect 14256 31666 14290 31700
rect 14324 31666 14358 31700
rect 14392 31666 14429 31700
rect 13165 31631 14429 31666
rect 13165 31597 13202 31631
rect 13236 31597 13270 31631
rect 13304 31597 13338 31631
rect 13372 31597 13406 31631
rect 13440 31597 13474 31631
rect 13508 31597 13542 31631
rect 13576 31597 13610 31631
rect 13644 31597 13678 31631
rect 13712 31597 13746 31631
rect 13780 31597 13814 31631
rect 13848 31597 13882 31631
rect 13916 31597 13950 31631
rect 13984 31597 14018 31631
rect 14052 31597 14086 31631
rect 14120 31597 14154 31631
rect 14188 31597 14222 31631
rect 14256 31597 14290 31631
rect 14324 31597 14358 31631
rect 14392 31597 14429 31631
rect 13165 31562 14429 31597
rect 13165 31528 13202 31562
rect 13236 31528 13270 31562
rect 13304 31528 13338 31562
rect 13372 31528 13406 31562
rect 13440 31528 13474 31562
rect 13508 31528 13542 31562
rect 13576 31528 13610 31562
rect 13644 31528 13678 31562
rect 13712 31528 13746 31562
rect 13780 31528 13814 31562
rect 13848 31528 13882 31562
rect 13916 31528 13950 31562
rect 13984 31528 14018 31562
rect 14052 31528 14086 31562
rect 14120 31528 14154 31562
rect 14188 31528 14222 31562
rect 14256 31528 14290 31562
rect 14324 31528 14358 31562
rect 14392 31528 14429 31562
rect 13165 31493 14429 31528
rect 13165 31459 13202 31493
rect 13236 31459 13270 31493
rect 13304 31459 13338 31493
rect 13372 31459 13406 31493
rect 13440 31459 13474 31493
rect 13508 31459 13542 31493
rect 13576 31459 13610 31493
rect 13644 31459 13678 31493
rect 13712 31459 13746 31493
rect 13780 31459 13814 31493
rect 13848 31459 13882 31493
rect 13916 31459 13950 31493
rect 13984 31459 14018 31493
rect 14052 31459 14086 31493
rect 14120 31459 14154 31493
rect 14188 31459 14222 31493
rect 14256 31459 14290 31493
rect 14324 31459 14358 31493
rect 14392 31459 14429 31493
rect 13165 31424 14429 31459
rect 13165 31390 13202 31424
rect 13236 31390 13270 31424
rect 13304 31390 13338 31424
rect 13372 31390 13406 31424
rect 13440 31390 13474 31424
rect 13508 31390 13542 31424
rect 13576 31390 13610 31424
rect 13644 31390 13678 31424
rect 13712 31390 13746 31424
rect 13780 31390 13814 31424
rect 13848 31390 13882 31424
rect 13916 31390 13950 31424
rect 13984 31390 14018 31424
rect 14052 31390 14086 31424
rect 14120 31390 14154 31424
rect 14188 31390 14222 31424
rect 14256 31390 14290 31424
rect 14324 31390 14358 31424
rect 14392 31390 14429 31424
rect 13165 31355 14429 31390
rect 13165 31321 13202 31355
rect 13236 31321 13270 31355
rect 13304 31321 13338 31355
rect 13372 31321 13406 31355
rect 13440 31321 13474 31355
rect 13508 31321 13542 31355
rect 13576 31321 13610 31355
rect 13644 31321 13678 31355
rect 13712 31321 13746 31355
rect 13780 31321 13814 31355
rect 13848 31321 13882 31355
rect 13916 31321 13950 31355
rect 13984 31321 14018 31355
rect 14052 31321 14086 31355
rect 14120 31321 14154 31355
rect 14188 31321 14222 31355
rect 14256 31321 14290 31355
rect 14324 31321 14358 31355
rect 14392 31321 14429 31355
rect 13165 31286 14429 31321
rect 13165 31252 13202 31286
rect 13236 31252 13270 31286
rect 13304 31252 13338 31286
rect 13372 31252 13406 31286
rect 13440 31252 13474 31286
rect 13508 31252 13542 31286
rect 13576 31252 13610 31286
rect 13644 31252 13678 31286
rect 13712 31252 13746 31286
rect 13780 31252 13814 31286
rect 13848 31252 13882 31286
rect 13916 31252 13950 31286
rect 13984 31252 14018 31286
rect 14052 31252 14086 31286
rect 14120 31252 14154 31286
rect 14188 31252 14222 31286
rect 14256 31252 14290 31286
rect 14324 31252 14358 31286
rect 14392 31252 14429 31286
rect 13165 31217 14429 31252
rect 13165 31183 13202 31217
rect 13236 31183 13270 31217
rect 13304 31183 13338 31217
rect 13372 31183 13406 31217
rect 13440 31183 13474 31217
rect 13508 31183 13542 31217
rect 13576 31183 13610 31217
rect 13644 31183 13678 31217
rect 13712 31183 13746 31217
rect 13780 31183 13814 31217
rect 13848 31183 13882 31217
rect 13916 31183 13950 31217
rect 13984 31183 14018 31217
rect 14052 31183 14086 31217
rect 14120 31183 14154 31217
rect 14188 31183 14222 31217
rect 14256 31183 14290 31217
rect 14324 31183 14358 31217
rect 14392 31183 14429 31217
rect 13165 31149 14429 31183
rect 9877 30636 13943 30670
rect 9877 30602 9913 30636
rect 9947 30602 9982 30636
rect 10016 30602 10051 30636
rect 10085 30602 10120 30636
rect 10154 30602 10189 30636
rect 10223 30602 10258 30636
rect 10292 30602 10327 30636
rect 10361 30602 10396 30636
rect 10430 30602 10465 30636
rect 10499 30635 13943 30636
rect 10499 30602 10610 30635
rect 9877 30601 10610 30602
rect 10644 30601 10679 30635
rect 10713 30601 10747 30635
rect 10781 30601 10815 30635
rect 10849 30601 10883 30635
rect 10917 30601 10951 30635
rect 10985 30601 11019 30635
rect 11053 30601 11087 30635
rect 11121 30601 11155 30635
rect 11189 30601 11223 30635
rect 11257 30601 11291 30635
rect 11325 30601 11359 30635
rect 11393 30601 11427 30635
rect 11461 30601 11495 30635
rect 11529 30601 11563 30635
rect 11597 30601 11631 30635
rect 11665 30601 11699 30635
rect 11733 30601 11767 30635
rect 11801 30601 11835 30635
rect 11869 30601 11903 30635
rect 11937 30601 11971 30635
rect 12005 30601 12039 30635
rect 12073 30601 12107 30635
rect 12141 30601 12175 30635
rect 12209 30601 12243 30635
rect 12277 30601 12311 30635
rect 12345 30601 12379 30635
rect 12413 30601 12447 30635
rect 12481 30601 12515 30635
rect 12549 30601 12583 30635
rect 12617 30601 12651 30635
rect 12685 30601 12719 30635
rect 12753 30601 12787 30635
rect 12821 30601 12855 30635
rect 12889 30601 12923 30635
rect 12957 30601 12991 30635
rect 13025 30601 13059 30635
rect 13093 30601 13127 30635
rect 13161 30601 13195 30635
rect 13229 30601 13263 30635
rect 13297 30601 13331 30635
rect 13365 30601 13399 30635
rect 13433 30601 13467 30635
rect 13501 30601 13535 30635
rect 13569 30601 13603 30635
rect 13637 30601 13671 30635
rect 13705 30601 13739 30635
rect 13773 30601 13807 30635
rect 13841 30601 13875 30635
rect 13909 30601 13943 30635
rect 9877 30568 13943 30601
rect 9877 30534 9913 30568
rect 9947 30534 9982 30568
rect 10016 30534 10051 30568
rect 10085 30534 10120 30568
rect 10154 30534 10189 30568
rect 10223 30534 10258 30568
rect 10292 30534 10327 30568
rect 10361 30534 10396 30568
rect 10430 30534 10465 30568
rect 10499 30560 13943 30568
rect 10499 30534 10610 30560
rect 9877 30526 10610 30534
rect 10644 30526 10679 30560
rect 10713 30526 10747 30560
rect 10781 30526 10815 30560
rect 10849 30526 10883 30560
rect 10917 30526 10951 30560
rect 10985 30526 11019 30560
rect 11053 30526 11087 30560
rect 11121 30526 11155 30560
rect 11189 30526 11223 30560
rect 11257 30526 11291 30560
rect 11325 30526 11359 30560
rect 11393 30526 11427 30560
rect 11461 30526 11495 30560
rect 11529 30526 11563 30560
rect 11597 30526 11631 30560
rect 11665 30526 11699 30560
rect 11733 30526 11767 30560
rect 11801 30526 11835 30560
rect 11869 30526 11903 30560
rect 11937 30526 11971 30560
rect 12005 30526 12039 30560
rect 12073 30526 12107 30560
rect 12141 30526 12175 30560
rect 12209 30526 12243 30560
rect 12277 30526 12311 30560
rect 12345 30526 12379 30560
rect 12413 30526 12447 30560
rect 12481 30526 12515 30560
rect 12549 30526 12583 30560
rect 12617 30526 12651 30560
rect 12685 30526 12719 30560
rect 12753 30526 12787 30560
rect 12821 30526 12855 30560
rect 12889 30526 12923 30560
rect 12957 30526 12991 30560
rect 13025 30526 13059 30560
rect 13093 30526 13127 30560
rect 13161 30526 13195 30560
rect 13229 30526 13263 30560
rect 13297 30526 13331 30560
rect 13365 30526 13399 30560
rect 13433 30526 13467 30560
rect 13501 30526 13535 30560
rect 13569 30526 13603 30560
rect 13637 30526 13671 30560
rect 13705 30526 13739 30560
rect 13773 30526 13807 30560
rect 13841 30526 13875 30560
rect 13909 30526 13943 30560
rect 9877 30500 13943 30526
rect 9877 30466 9913 30500
rect 9947 30466 9982 30500
rect 10016 30466 10051 30500
rect 10085 30466 10120 30500
rect 10154 30466 10189 30500
rect 10223 30466 10258 30500
rect 10292 30466 10327 30500
rect 10361 30466 10396 30500
rect 10430 30466 10465 30500
rect 10499 30485 13943 30500
rect 10499 30466 10610 30485
rect 9877 30451 10610 30466
rect 10644 30451 10679 30485
rect 10713 30451 10747 30485
rect 10781 30451 10815 30485
rect 10849 30451 10883 30485
rect 10917 30451 10951 30485
rect 10985 30451 11019 30485
rect 11053 30451 11087 30485
rect 11121 30451 11155 30485
rect 11189 30451 11223 30485
rect 11257 30451 11291 30485
rect 11325 30451 11359 30485
rect 11393 30451 11427 30485
rect 11461 30451 11495 30485
rect 11529 30451 11563 30485
rect 11597 30451 11631 30485
rect 11665 30451 11699 30485
rect 11733 30451 11767 30485
rect 11801 30451 11835 30485
rect 11869 30451 11903 30485
rect 11937 30451 11971 30485
rect 12005 30451 12039 30485
rect 12073 30451 12107 30485
rect 12141 30451 12175 30485
rect 12209 30451 12243 30485
rect 12277 30451 12311 30485
rect 12345 30451 12379 30485
rect 12413 30451 12447 30485
rect 12481 30451 12515 30485
rect 12549 30451 12583 30485
rect 12617 30451 12651 30485
rect 12685 30451 12719 30485
rect 12753 30451 12787 30485
rect 12821 30451 12855 30485
rect 12889 30451 12923 30485
rect 12957 30451 12991 30485
rect 13025 30451 13059 30485
rect 13093 30451 13127 30485
rect 13161 30451 13195 30485
rect 13229 30451 13263 30485
rect 13297 30451 13331 30485
rect 13365 30451 13399 30485
rect 13433 30451 13467 30485
rect 13501 30451 13535 30485
rect 13569 30451 13603 30485
rect 13637 30451 13671 30485
rect 13705 30451 13739 30485
rect 13773 30451 13807 30485
rect 13841 30451 13875 30485
rect 13909 30451 13943 30485
rect 9877 30432 13943 30451
rect 9877 30398 9913 30432
rect 9947 30398 9982 30432
rect 10016 30398 10051 30432
rect 10085 30398 10120 30432
rect 10154 30398 10189 30432
rect 10223 30398 10258 30432
rect 10292 30398 10327 30432
rect 10361 30398 10396 30432
rect 10430 30398 10465 30432
rect 10499 30416 13943 30432
rect 10499 30398 10535 30416
rect 9877 30364 10535 30398
rect 9877 30330 9913 30364
rect 9947 30330 9982 30364
rect 10016 30330 10051 30364
rect 10085 30330 10120 30364
rect 10154 30330 10189 30364
rect 10223 30330 10258 30364
rect 10292 30330 10327 30364
rect 10361 30330 10396 30364
rect 10430 30330 10465 30364
rect 10499 30330 10535 30364
rect 9877 30296 10535 30330
rect 9877 30262 9913 30296
rect 9947 30262 9982 30296
rect 10016 30262 10051 30296
rect 10085 30262 10120 30296
rect 10154 30262 10189 30296
rect 10223 30262 10258 30296
rect 10292 30262 10327 30296
rect 10361 30262 10396 30296
rect 10430 30262 10465 30296
rect 10499 30262 10535 30296
rect 9877 30228 10535 30262
rect 9877 30194 9913 30228
rect 9947 30194 9982 30228
rect 10016 30194 10051 30228
rect 10085 30194 10120 30228
rect 10154 30194 10189 30228
rect 10223 30194 10258 30228
rect 10292 30194 10327 30228
rect 10361 30194 10396 30228
rect 10430 30194 10465 30228
rect 10499 30194 10535 30228
rect 9877 30160 10535 30194
rect 9877 30126 9913 30160
rect 9947 30126 9982 30160
rect 10016 30126 10051 30160
rect 10085 30126 10120 30160
rect 10154 30126 10189 30160
rect 10223 30126 10258 30160
rect 10292 30126 10327 30160
rect 10361 30126 10396 30160
rect 10430 30126 10465 30160
rect 10499 30126 10535 30160
rect 9877 30092 10535 30126
rect 9877 30058 9913 30092
rect 9947 30058 9982 30092
rect 10016 30058 10051 30092
rect 10085 30058 10120 30092
rect 10154 30058 10189 30092
rect 10223 30058 10258 30092
rect 10292 30058 10327 30092
rect 10361 30058 10396 30092
rect 10430 30058 10465 30092
rect 10499 30058 10535 30092
rect 9877 30024 10535 30058
rect 9877 29990 9913 30024
rect 9947 29990 9982 30024
rect 10016 29990 10051 30024
rect 10085 29990 10120 30024
rect 10154 29990 10189 30024
rect 10223 29990 10258 30024
rect 10292 29990 10327 30024
rect 10361 29990 10396 30024
rect 10430 29990 10465 30024
rect 10499 29990 10535 30024
rect 9877 29956 10535 29990
rect 9877 29922 9913 29956
rect 9947 29922 9982 29956
rect 10016 29922 10051 29956
rect 10085 29922 10120 29956
rect 10154 29922 10189 29956
rect 10223 29922 10258 29956
rect 10292 29922 10327 29956
rect 10361 29922 10396 29956
rect 10430 29922 10465 29956
rect 10499 29922 10535 29956
rect 9877 29888 10535 29922
rect 9877 29854 9913 29888
rect 9947 29854 9982 29888
rect 10016 29854 10051 29888
rect 10085 29854 10120 29888
rect 10154 29854 10189 29888
rect 10223 29854 10258 29888
rect 10292 29854 10327 29888
rect 10361 29854 10396 29888
rect 10430 29854 10465 29888
rect 10499 29854 10535 29888
rect 9877 29820 10535 29854
rect 9877 29786 9913 29820
rect 9947 29786 9982 29820
rect 10016 29786 10051 29820
rect 10085 29786 10120 29820
rect 10154 29786 10189 29820
rect 10223 29786 10258 29820
rect 10292 29786 10327 29820
rect 10361 29786 10396 29820
rect 10430 29786 10465 29820
rect 10499 29786 10535 29820
rect 9877 29752 10535 29786
rect 9877 29718 9913 29752
rect 9947 29718 9982 29752
rect 10016 29718 10051 29752
rect 10085 29718 10120 29752
rect 10154 29718 10189 29752
rect 10223 29718 10258 29752
rect 10292 29718 10327 29752
rect 10361 29718 10396 29752
rect 10430 29718 10465 29752
rect 10499 29718 10535 29752
rect 9877 29684 10535 29718
rect 9877 29650 9913 29684
rect 9947 29650 9982 29684
rect 10016 29650 10051 29684
rect 10085 29650 10120 29684
rect 10154 29650 10189 29684
rect 10223 29650 10258 29684
rect 10292 29650 10327 29684
rect 10361 29650 10396 29684
rect 10430 29650 10465 29684
rect 10499 29650 10535 29684
rect 9877 29616 10535 29650
rect 9877 29582 9913 29616
rect 9947 29582 9982 29616
rect 10016 29582 10051 29616
rect 10085 29582 10120 29616
rect 10154 29582 10189 29616
rect 10223 29582 10258 29616
rect 10292 29582 10327 29616
rect 10361 29582 10396 29616
rect 10430 29582 10465 29616
rect 10499 29582 10535 29616
rect 9877 29548 10535 29582
rect 9877 29514 9913 29548
rect 9947 29514 9982 29548
rect 10016 29514 10051 29548
rect 10085 29514 10120 29548
rect 10154 29514 10189 29548
rect 10223 29514 10258 29548
rect 10292 29514 10327 29548
rect 10361 29514 10396 29548
rect 10430 29514 10465 29548
rect 10499 29514 10535 29548
rect 9877 29480 10535 29514
rect 9877 29446 9913 29480
rect 9947 29446 9982 29480
rect 10016 29446 10051 29480
rect 10085 29446 10120 29480
rect 10154 29446 10189 29480
rect 10223 29446 10258 29480
rect 10292 29446 10327 29480
rect 10361 29446 10396 29480
rect 10430 29446 10465 29480
rect 10499 29446 10535 29480
rect 9877 29412 10535 29446
rect 9877 29378 9913 29412
rect 9947 29378 9982 29412
rect 10016 29378 10051 29412
rect 10085 29378 10120 29412
rect 10154 29378 10189 29412
rect 10223 29378 10258 29412
rect 10292 29378 10327 29412
rect 10361 29378 10396 29412
rect 10430 29378 10465 29412
rect 10499 29378 10535 29412
rect 9877 29344 10535 29378
rect 9877 29310 9913 29344
rect 9947 29310 9982 29344
rect 10016 29310 10051 29344
rect 10085 29310 10120 29344
rect 10154 29310 10189 29344
rect 10223 29310 10258 29344
rect 10292 29310 10327 29344
rect 10361 29310 10396 29344
rect 10430 29310 10465 29344
rect 10499 29310 10535 29344
rect 9877 29276 10535 29310
rect 9877 29242 9913 29276
rect 9947 29242 9982 29276
rect 10016 29242 10051 29276
rect 10085 29242 10120 29276
rect 10154 29242 10189 29276
rect 10223 29242 10258 29276
rect 10292 29242 10327 29276
rect 10361 29242 10396 29276
rect 10430 29242 10465 29276
rect 10499 29242 10535 29276
rect 9877 29208 10535 29242
rect 9877 29174 9913 29208
rect 9947 29174 9982 29208
rect 10016 29174 10051 29208
rect 10085 29174 10120 29208
rect 10154 29174 10189 29208
rect 10223 29174 10258 29208
rect 10292 29174 10327 29208
rect 10361 29174 10396 29208
rect 10430 29174 10465 29208
rect 10499 29174 10535 29208
rect 9877 29140 10535 29174
rect 9877 29106 9913 29140
rect 9947 29106 9982 29140
rect 10016 29106 10051 29140
rect 10085 29106 10120 29140
rect 10154 29106 10189 29140
rect 10223 29106 10258 29140
rect 10292 29106 10327 29140
rect 10361 29106 10396 29140
rect 10430 29106 10465 29140
rect 10499 29106 10535 29140
rect 9877 29072 10535 29106
rect 9877 29038 9913 29072
rect 9947 29038 9982 29072
rect 10016 29038 10051 29072
rect 10085 29038 10120 29072
rect 10154 29038 10189 29072
rect 10223 29038 10258 29072
rect 10292 29038 10327 29072
rect 10361 29038 10396 29072
rect 10430 29038 10465 29072
rect 10499 29038 10535 29072
rect 9877 29004 10535 29038
rect 9877 28970 9913 29004
rect 9947 28970 9982 29004
rect 10016 28970 10051 29004
rect 10085 28970 10120 29004
rect 10154 28970 10189 29004
rect 10223 28970 10258 29004
rect 10292 28970 10327 29004
rect 10361 28970 10396 29004
rect 10430 28970 10465 29004
rect 10499 28970 10535 29004
rect 9877 28936 10535 28970
rect 9877 28902 9913 28936
rect 9947 28902 9982 28936
rect 10016 28902 10051 28936
rect 10085 28902 10120 28936
rect 10154 28902 10189 28936
rect 10223 28902 10258 28936
rect 10292 28902 10327 28936
rect 10361 28902 10396 28936
rect 10430 28902 10465 28936
rect 10499 28902 10535 28936
rect 9877 28868 10535 28902
rect 9877 28834 9913 28868
rect 9947 28834 9982 28868
rect 10016 28834 10051 28868
rect 10085 28834 10120 28868
rect 10154 28834 10189 28868
rect 10223 28834 10258 28868
rect 10292 28834 10327 28868
rect 10361 28834 10396 28868
rect 10430 28834 10465 28868
rect 10499 28834 10535 28868
rect 9877 28800 10535 28834
rect 9877 28766 9913 28800
rect 9947 28766 9982 28800
rect 10016 28766 10051 28800
rect 10085 28766 10120 28800
rect 10154 28766 10189 28800
rect 10223 28766 10258 28800
rect 10292 28766 10327 28800
rect 10361 28766 10396 28800
rect 10430 28766 10465 28800
rect 10499 28766 10535 28800
rect 9877 28732 10535 28766
rect 9877 28698 9913 28732
rect 9947 28698 9982 28732
rect 10016 28698 10051 28732
rect 10085 28698 10120 28732
rect 10154 28698 10189 28732
rect 10223 28698 10258 28732
rect 10292 28698 10327 28732
rect 10361 28698 10396 28732
rect 10430 28698 10465 28732
rect 10499 28698 10535 28732
rect 9877 28664 10535 28698
rect 9877 28630 9913 28664
rect 9947 28630 9982 28664
rect 10016 28630 10051 28664
rect 10085 28630 10120 28664
rect 10154 28630 10189 28664
rect 10223 28630 10258 28664
rect 10292 28630 10327 28664
rect 10361 28630 10396 28664
rect 10430 28630 10465 28664
rect 10499 28630 10535 28664
rect 9877 28596 10535 28630
rect 9877 28562 9913 28596
rect 9947 28562 9982 28596
rect 10016 28562 10051 28596
rect 10085 28562 10120 28596
rect 10154 28562 10189 28596
rect 10223 28562 10258 28596
rect 10292 28562 10327 28596
rect 10361 28562 10396 28596
rect 10430 28562 10465 28596
rect 10499 28562 10535 28596
rect 9877 28528 10535 28562
rect 9877 28494 9913 28528
rect 9947 28494 9982 28528
rect 10016 28494 10051 28528
rect 10085 28494 10120 28528
rect 10154 28494 10189 28528
rect 10223 28494 10258 28528
rect 10292 28494 10327 28528
rect 10361 28494 10396 28528
rect 10430 28494 10465 28528
rect 10499 28494 10535 28528
rect 9877 28460 10535 28494
rect 9877 28426 9913 28460
rect 9947 28426 9982 28460
rect 10016 28426 10051 28460
rect 10085 28426 10120 28460
rect 10154 28426 10189 28460
rect 10223 28426 10258 28460
rect 10292 28426 10327 28460
rect 10361 28426 10396 28460
rect 10430 28426 10465 28460
rect 10499 28426 10535 28460
rect 9877 28392 10535 28426
rect 9877 28358 9913 28392
rect 9947 28358 9982 28392
rect 10016 28358 10051 28392
rect 10085 28358 10120 28392
rect 10154 28358 10189 28392
rect 10223 28358 10258 28392
rect 10292 28358 10327 28392
rect 10361 28358 10396 28392
rect 10430 28358 10465 28392
rect 10499 28358 10535 28392
rect 9877 28324 10535 28358
rect 9877 28290 9913 28324
rect 9947 28290 9982 28324
rect 10016 28290 10051 28324
rect 10085 28290 10120 28324
rect 10154 28290 10189 28324
rect 10223 28290 10258 28324
rect 10292 28290 10327 28324
rect 10361 28290 10396 28324
rect 10430 28290 10465 28324
rect 10499 28290 10535 28324
rect 9877 28256 10535 28290
rect 9877 28222 9913 28256
rect 9947 28222 9982 28256
rect 10016 28222 10051 28256
rect 10085 28222 10120 28256
rect 10154 28222 10189 28256
rect 10223 28222 10258 28256
rect 10292 28222 10327 28256
rect 10361 28222 10396 28256
rect 10430 28222 10465 28256
rect 10499 28222 10535 28256
rect 9877 28188 10535 28222
rect 9877 28154 9913 28188
rect 9947 28154 9982 28188
rect 10016 28154 10051 28188
rect 10085 28154 10120 28188
rect 10154 28154 10189 28188
rect 10223 28154 10258 28188
rect 10292 28154 10327 28188
rect 10361 28154 10396 28188
rect 10430 28154 10465 28188
rect 10499 28154 10535 28188
rect 9877 28120 10535 28154
rect 9877 28086 9913 28120
rect 9947 28086 9982 28120
rect 10016 28086 10051 28120
rect 10085 28086 10120 28120
rect 10154 28086 10189 28120
rect 10223 28086 10258 28120
rect 10292 28086 10327 28120
rect 10361 28086 10396 28120
rect 10430 28086 10465 28120
rect 10499 28086 10535 28120
rect 9877 28052 10535 28086
rect 9877 28018 9913 28052
rect 9947 28018 9982 28052
rect 10016 28018 10051 28052
rect 10085 28018 10120 28052
rect 10154 28018 10189 28052
rect 10223 28018 10258 28052
rect 10292 28018 10327 28052
rect 10361 28018 10396 28052
rect 10430 28018 10465 28052
rect 10499 28018 10535 28052
rect 9877 27983 10535 28018
rect 9877 27949 9913 27983
rect 9947 27949 9982 27983
rect 10016 27949 10051 27983
rect 10085 27949 10120 27983
rect 10154 27949 10189 27983
rect 10223 27949 10258 27983
rect 10292 27949 10327 27983
rect 10361 27949 10396 27983
rect 10430 27949 10465 27983
rect 10499 27949 10535 27983
rect 9877 27914 10535 27949
rect 9877 27880 9913 27914
rect 9947 27880 9982 27914
rect 10016 27880 10051 27914
rect 10085 27880 10120 27914
rect 10154 27880 10189 27914
rect 10223 27880 10258 27914
rect 10292 27880 10327 27914
rect 10361 27880 10396 27914
rect 10430 27880 10465 27914
rect 10499 27880 10535 27914
rect 9877 27845 10535 27880
rect 9877 27811 9913 27845
rect 9947 27811 9982 27845
rect 10016 27811 10051 27845
rect 10085 27811 10120 27845
rect 10154 27811 10189 27845
rect 10223 27811 10258 27845
rect 10292 27811 10327 27845
rect 10361 27811 10396 27845
rect 10430 27811 10465 27845
rect 10499 27811 10535 27845
rect 9877 27776 10535 27811
rect 9877 27742 9913 27776
rect 9947 27742 9982 27776
rect 10016 27742 10051 27776
rect 10085 27742 10120 27776
rect 10154 27742 10189 27776
rect 10223 27742 10258 27776
rect 10292 27742 10327 27776
rect 10361 27742 10396 27776
rect 10430 27742 10465 27776
rect 10499 27742 10535 27776
rect 9877 27707 10535 27742
rect 9877 27673 9913 27707
rect 9947 27673 9982 27707
rect 10016 27673 10051 27707
rect 10085 27673 10120 27707
rect 10154 27673 10189 27707
rect 10223 27673 10258 27707
rect 10292 27673 10327 27707
rect 10361 27673 10396 27707
rect 10430 27673 10465 27707
rect 10499 27673 10535 27707
rect 9877 27638 10535 27673
rect 9877 27604 9913 27638
rect 9947 27604 9982 27638
rect 10016 27604 10051 27638
rect 10085 27604 10120 27638
rect 10154 27604 10189 27638
rect 10223 27604 10258 27638
rect 10292 27604 10327 27638
rect 10361 27604 10396 27638
rect 10430 27604 10465 27638
rect 10499 27604 10535 27638
rect 9877 27569 10535 27604
rect 9877 27535 9913 27569
rect 9947 27535 9982 27569
rect 10016 27535 10051 27569
rect 10085 27535 10120 27569
rect 10154 27535 10189 27569
rect 10223 27535 10258 27569
rect 10292 27535 10327 27569
rect 10361 27535 10396 27569
rect 10430 27535 10465 27569
rect 10499 27535 10535 27569
rect 9877 27500 10535 27535
rect 9877 27466 9913 27500
rect 9947 27466 9982 27500
rect 10016 27466 10051 27500
rect 10085 27466 10120 27500
rect 10154 27466 10189 27500
rect 10223 27466 10258 27500
rect 10292 27466 10327 27500
rect 10361 27466 10396 27500
rect 10430 27466 10465 27500
rect 10499 27466 10535 27500
rect 9877 27431 10535 27466
rect 9877 27397 9913 27431
rect 9947 27397 9982 27431
rect 10016 27397 10051 27431
rect 10085 27397 10120 27431
rect 10154 27397 10189 27431
rect 10223 27397 10258 27431
rect 10292 27397 10327 27431
rect 10361 27397 10396 27431
rect 10430 27397 10465 27431
rect 10499 27397 10535 27431
rect 9877 27362 10535 27397
rect 9877 27328 9913 27362
rect 9947 27328 9982 27362
rect 10016 27328 10051 27362
rect 10085 27328 10120 27362
rect 10154 27328 10189 27362
rect 10223 27328 10258 27362
rect 10292 27328 10327 27362
rect 10361 27328 10396 27362
rect 10430 27328 10465 27362
rect 10499 27328 10535 27362
rect 9877 27293 10535 27328
rect 9877 27259 9913 27293
rect 9947 27259 9982 27293
rect 10016 27259 10051 27293
rect 10085 27259 10120 27293
rect 10154 27259 10189 27293
rect 10223 27259 10258 27293
rect 10292 27259 10327 27293
rect 10361 27259 10396 27293
rect 10430 27259 10465 27293
rect 10499 27259 10535 27293
rect 9877 27224 10535 27259
rect 9877 27190 9913 27224
rect 9947 27190 9982 27224
rect 10016 27190 10051 27224
rect 10085 27190 10120 27224
rect 10154 27190 10189 27224
rect 10223 27190 10258 27224
rect 10292 27190 10327 27224
rect 10361 27190 10396 27224
rect 10430 27190 10465 27224
rect 10499 27190 10535 27224
rect 9877 27155 10535 27190
rect 9877 27121 9913 27155
rect 9947 27121 9982 27155
rect 10016 27121 10051 27155
rect 10085 27121 10120 27155
rect 10154 27121 10189 27155
rect 10223 27121 10258 27155
rect 10292 27121 10327 27155
rect 10361 27121 10396 27155
rect 10430 27121 10465 27155
rect 10499 27121 10535 27155
rect 9877 27086 10535 27121
rect 9877 27052 9913 27086
rect 9947 27052 9982 27086
rect 10016 27052 10051 27086
rect 10085 27052 10120 27086
rect 10154 27052 10189 27086
rect 10223 27052 10258 27086
rect 10292 27052 10327 27086
rect 10361 27052 10396 27086
rect 10430 27052 10465 27086
rect 10499 27052 10535 27086
rect 9877 26972 10535 27052
rect 13703 30401 13943 30416
rect 13703 29007 13738 30401
rect 13908 29007 13943 30401
rect 13703 28972 13943 29007
rect 13703 28938 13738 28972
rect 13772 28938 13806 28972
rect 13840 28938 13874 28972
rect 13908 28938 13943 28972
rect 13703 28903 13943 28938
rect 13703 28869 13738 28903
rect 13772 28869 13806 28903
rect 13840 28869 13874 28903
rect 13908 28869 13943 28903
rect 13703 28834 13943 28869
rect 13703 28800 13738 28834
rect 13772 28800 13806 28834
rect 13840 28800 13874 28834
rect 13908 28800 13943 28834
rect 13703 28765 13943 28800
rect 13703 28731 13738 28765
rect 13772 28731 13806 28765
rect 13840 28731 13874 28765
rect 13908 28731 13943 28765
rect 13703 28696 13943 28731
rect 13703 28662 13738 28696
rect 13772 28662 13806 28696
rect 13840 28662 13874 28696
rect 13908 28662 13943 28696
rect 13703 28627 13943 28662
rect 13703 28593 13738 28627
rect 13772 28593 13806 28627
rect 13840 28593 13874 28627
rect 13908 28593 13943 28627
rect 13703 28558 13943 28593
rect 13703 28524 13738 28558
rect 13772 28524 13806 28558
rect 13840 28524 13874 28558
rect 13908 28524 13943 28558
rect 13703 28489 13943 28524
rect 13703 28455 13738 28489
rect 13772 28455 13806 28489
rect 13840 28455 13874 28489
rect 13908 28455 13943 28489
rect 13703 28420 13943 28455
rect 13703 28386 13738 28420
rect 13772 28386 13806 28420
rect 13840 28386 13874 28420
rect 13908 28386 13943 28420
rect 13703 28351 13943 28386
rect 13703 28317 13738 28351
rect 13772 28317 13806 28351
rect 13840 28317 13874 28351
rect 13908 28317 13943 28351
rect 13703 28282 13943 28317
rect 13703 28248 13738 28282
rect 13772 28248 13806 28282
rect 13840 28248 13874 28282
rect 13908 28248 13943 28282
rect 13703 28213 13943 28248
rect 13703 28179 13738 28213
rect 13772 28179 13806 28213
rect 13840 28179 13874 28213
rect 13908 28179 13943 28213
rect 13703 28144 13943 28179
rect 13703 28110 13738 28144
rect 13772 28110 13806 28144
rect 13840 28110 13874 28144
rect 13908 28110 13943 28144
rect 13703 28075 13943 28110
rect 13703 28041 13738 28075
rect 13772 28041 13806 28075
rect 13840 28041 13874 28075
rect 13908 28041 13943 28075
rect 13703 28006 13943 28041
rect 13703 27972 13738 28006
rect 13772 27972 13806 28006
rect 13840 27972 13874 28006
rect 13908 27972 13943 28006
rect 13703 27937 13943 27972
rect 13703 27903 13738 27937
rect 13772 27903 13806 27937
rect 13840 27903 13874 27937
rect 13908 27903 13943 27937
rect 13703 27868 13943 27903
rect 13703 27834 13738 27868
rect 13772 27834 13806 27868
rect 13840 27834 13874 27868
rect 13908 27834 13943 27868
rect 13703 27799 13943 27834
rect 13703 27765 13738 27799
rect 13772 27765 13806 27799
rect 13840 27765 13874 27799
rect 13908 27765 13943 27799
rect 13703 27730 13943 27765
rect 13703 27696 13738 27730
rect 13772 27696 13806 27730
rect 13840 27696 13874 27730
rect 13908 27696 13943 27730
rect 13703 27661 13943 27696
rect 13703 27627 13738 27661
rect 13772 27627 13806 27661
rect 13840 27627 13874 27661
rect 13908 27627 13943 27661
rect 13703 27592 13943 27627
rect 13703 27558 13738 27592
rect 13772 27558 13806 27592
rect 13840 27558 13874 27592
rect 13908 27558 13943 27592
rect 13703 27523 13943 27558
rect 13703 27489 13738 27523
rect 13772 27489 13806 27523
rect 13840 27489 13874 27523
rect 13908 27489 13943 27523
rect 13703 27454 13943 27489
rect 13703 27420 13738 27454
rect 13772 27420 13806 27454
rect 13840 27420 13874 27454
rect 13908 27420 13943 27454
rect 13703 27385 13943 27420
rect 13703 27351 13738 27385
rect 13772 27351 13806 27385
rect 13840 27351 13874 27385
rect 13908 27351 13943 27385
rect 13703 27316 13943 27351
rect 13703 27282 13738 27316
rect 13772 27282 13806 27316
rect 13840 27282 13874 27316
rect 13908 27282 13943 27316
rect 13703 27247 13943 27282
rect 13703 27213 13738 27247
rect 13772 27213 13806 27247
rect 13840 27213 13874 27247
rect 13908 27213 13943 27247
rect 13703 27178 13943 27213
rect 13703 27144 13738 27178
rect 13772 27144 13806 27178
rect 13840 27144 13874 27178
rect 13908 27144 13943 27178
rect 13703 27109 13943 27144
rect 13703 27075 13738 27109
rect 13772 27075 13806 27109
rect 13840 27075 13874 27109
rect 13908 27075 13943 27109
rect 13703 27040 13943 27075
rect 13703 27006 13738 27040
rect 13772 27006 13806 27040
rect 13840 27006 13874 27040
rect 13908 27006 13943 27040
rect 13703 26972 13943 27006
rect 9877 26938 13943 26972
rect 9877 26904 9911 26938
rect 9945 26904 9980 26938
rect 10014 26904 10049 26938
rect 10083 26904 10118 26938
rect 10152 26904 10187 26938
rect 10221 26904 10256 26938
rect 10290 26904 10325 26938
rect 10359 26904 10394 26938
rect 10428 26904 10463 26938
rect 10497 26904 10532 26938
rect 10566 26904 10601 26938
rect 10635 26904 10670 26938
rect 10704 26904 10739 26938
rect 10773 26904 10808 26938
rect 10842 26904 10877 26938
rect 10911 26904 10946 26938
rect 10980 26904 11015 26938
rect 11049 26904 11084 26938
rect 11118 26904 11153 26938
rect 11187 26904 11222 26938
rect 11256 26904 11291 26938
rect 11325 26904 11359 26938
rect 11393 26904 11427 26938
rect 11461 26904 11495 26938
rect 11529 26904 11563 26938
rect 11597 26904 11631 26938
rect 11665 26904 11699 26938
rect 11733 26904 11767 26938
rect 11801 26904 11835 26938
rect 11869 26904 11903 26938
rect 11937 26904 11971 26938
rect 12005 26904 12039 26938
rect 12073 26904 12107 26938
rect 12141 26904 12175 26938
rect 12209 26904 12243 26938
rect 12277 26904 12311 26938
rect 12345 26904 12379 26938
rect 12413 26904 12447 26938
rect 12481 26904 12515 26938
rect 12549 26904 12583 26938
rect 12617 26904 12651 26938
rect 12685 26904 12719 26938
rect 12753 26904 12787 26938
rect 12821 26904 12855 26938
rect 12889 26904 12923 26938
rect 12957 26904 12991 26938
rect 13025 26904 13059 26938
rect 13093 26904 13127 26938
rect 13161 26904 13195 26938
rect 13229 26904 13263 26938
rect 13297 26904 13331 26938
rect 13365 26904 13399 26938
rect 13433 26904 13467 26938
rect 13501 26904 13535 26938
rect 13569 26904 13603 26938
rect 13637 26904 13671 26938
rect 13705 26904 13739 26938
rect 13773 26904 13807 26938
rect 13841 26904 13875 26938
rect 13909 26904 13943 26938
rect 9877 26866 13943 26904
rect 9877 26832 9911 26866
rect 9945 26832 9980 26866
rect 10014 26832 10049 26866
rect 10083 26832 10118 26866
rect 10152 26832 10187 26866
rect 10221 26832 10256 26866
rect 10290 26832 10325 26866
rect 10359 26832 10394 26866
rect 10428 26832 10463 26866
rect 10497 26832 10532 26866
rect 10566 26832 10601 26866
rect 10635 26832 10670 26866
rect 10704 26832 10739 26866
rect 10773 26832 10808 26866
rect 10842 26832 10877 26866
rect 10911 26832 10946 26866
rect 10980 26832 11015 26866
rect 11049 26832 11084 26866
rect 11118 26832 11153 26866
rect 11187 26832 11222 26866
rect 11256 26832 11291 26866
rect 11325 26832 11359 26866
rect 11393 26832 11427 26866
rect 11461 26832 11495 26866
rect 11529 26832 11563 26866
rect 11597 26832 11631 26866
rect 11665 26832 11699 26866
rect 11733 26832 11767 26866
rect 11801 26832 11835 26866
rect 11869 26832 11903 26866
rect 11937 26832 11971 26866
rect 12005 26832 12039 26866
rect 12073 26832 12107 26866
rect 12141 26832 12175 26866
rect 12209 26832 12243 26866
rect 12277 26832 12311 26866
rect 12345 26832 12379 26866
rect 12413 26832 12447 26866
rect 12481 26832 12515 26866
rect 12549 26832 12583 26866
rect 12617 26832 12651 26866
rect 12685 26832 12719 26866
rect 12753 26832 12787 26866
rect 12821 26832 12855 26866
rect 12889 26832 12923 26866
rect 12957 26832 12991 26866
rect 13025 26832 13059 26866
rect 13093 26832 13127 26866
rect 13161 26832 13195 26866
rect 13229 26832 13263 26866
rect 13297 26832 13331 26866
rect 13365 26832 13399 26866
rect 13433 26832 13467 26866
rect 13501 26832 13535 26866
rect 13569 26832 13603 26866
rect 13637 26832 13671 26866
rect 13705 26832 13739 26866
rect 13773 26832 13807 26866
rect 13841 26832 13875 26866
rect 13909 26832 13943 26866
rect 9877 26794 13943 26832
rect 9877 26760 9911 26794
rect 9945 26760 9980 26794
rect 10014 26760 10049 26794
rect 10083 26760 10118 26794
rect 10152 26760 10187 26794
rect 10221 26760 10256 26794
rect 10290 26760 10325 26794
rect 10359 26760 10394 26794
rect 10428 26760 10463 26794
rect 10497 26760 10532 26794
rect 10566 26760 10601 26794
rect 10635 26760 10670 26794
rect 10704 26760 10739 26794
rect 10773 26760 10808 26794
rect 10842 26760 10877 26794
rect 10911 26760 10946 26794
rect 10980 26760 11015 26794
rect 11049 26760 11084 26794
rect 11118 26760 11153 26794
rect 11187 26760 11222 26794
rect 11256 26760 11291 26794
rect 11325 26760 11359 26794
rect 11393 26760 11427 26794
rect 11461 26760 11495 26794
rect 11529 26760 11563 26794
rect 11597 26760 11631 26794
rect 11665 26760 11699 26794
rect 11733 26760 11767 26794
rect 11801 26760 11835 26794
rect 11869 26760 11903 26794
rect 11937 26760 11971 26794
rect 12005 26760 12039 26794
rect 12073 26760 12107 26794
rect 12141 26760 12175 26794
rect 12209 26760 12243 26794
rect 12277 26760 12311 26794
rect 12345 26760 12379 26794
rect 12413 26760 12447 26794
rect 12481 26760 12515 26794
rect 12549 26760 12583 26794
rect 12617 26760 12651 26794
rect 12685 26760 12719 26794
rect 12753 26760 12787 26794
rect 12821 26760 12855 26794
rect 12889 26760 12923 26794
rect 12957 26760 12991 26794
rect 13025 26760 13059 26794
rect 13093 26760 13127 26794
rect 13161 26760 13195 26794
rect 13229 26760 13263 26794
rect 13297 26760 13331 26794
rect 13365 26760 13399 26794
rect 13433 26760 13467 26794
rect 13501 26760 13535 26794
rect 13569 26760 13603 26794
rect 13637 26760 13671 26794
rect 13705 26760 13739 26794
rect 13773 26760 13807 26794
rect 13841 26760 13875 26794
rect 13909 26760 13943 26794
rect 9877 26726 13943 26760
rect 9877 26224 14429 26248
rect 9877 26199 14233 26224
rect 9877 26165 9911 26199
rect 9945 26165 9980 26199
rect 10014 26165 10049 26199
rect 10083 26165 10118 26199
rect 10152 26165 10187 26199
rect 10221 26165 10256 26199
rect 10290 26165 10325 26199
rect 10359 26165 10394 26199
rect 10428 26165 10463 26199
rect 10497 26165 10532 26199
rect 10566 26165 10601 26199
rect 10635 26165 10670 26199
rect 10704 26165 10739 26199
rect 10773 26165 10807 26199
rect 10841 26165 10875 26199
rect 10909 26165 10943 26199
rect 10977 26165 11011 26199
rect 11045 26165 11079 26199
rect 11113 26165 11147 26199
rect 11181 26165 11215 26199
rect 11249 26165 11283 26199
rect 11317 26165 11351 26199
rect 11385 26165 11419 26199
rect 11453 26165 11487 26199
rect 11521 26165 11555 26199
rect 11589 26165 11623 26199
rect 11657 26165 11691 26199
rect 11725 26165 11759 26199
rect 11793 26165 11827 26199
rect 11861 26165 11895 26199
rect 11929 26165 11963 26199
rect 11997 26165 12031 26199
rect 12065 26165 12099 26199
rect 12133 26165 12167 26199
rect 12201 26165 12235 26199
rect 12269 26165 12303 26199
rect 12337 26165 12371 26199
rect 12405 26165 12439 26199
rect 12473 26165 12507 26199
rect 12541 26165 12575 26199
rect 12609 26165 12643 26199
rect 12677 26165 12711 26199
rect 12745 26165 12779 26199
rect 12813 26165 12847 26199
rect 12881 26165 12915 26199
rect 12949 26165 12983 26199
rect 13017 26165 13051 26199
rect 13085 26165 13119 26199
rect 13153 26165 13187 26199
rect 13221 26165 13255 26199
rect 13289 26165 13323 26199
rect 13357 26165 13391 26199
rect 13425 26165 13459 26199
rect 13493 26165 13527 26199
rect 13561 26165 13595 26199
rect 13629 26165 13663 26199
rect 13697 26165 13731 26199
rect 13765 26165 13799 26199
rect 13833 26165 13867 26199
rect 13901 26165 13935 26199
rect 13969 26165 14003 26199
rect 14037 26165 14071 26199
rect 14105 26165 14139 26199
rect 14173 26165 14233 26199
rect 9877 26129 14233 26165
rect 9877 26095 9911 26129
rect 9945 26095 9980 26129
rect 10014 26095 10049 26129
rect 10083 26095 10118 26129
rect 10152 26095 10187 26129
rect 10221 26095 10256 26129
rect 10290 26095 10325 26129
rect 10359 26095 10394 26129
rect 10428 26095 10463 26129
rect 10497 26095 10532 26129
rect 10566 26095 10601 26129
rect 10635 26095 10670 26129
rect 10704 26095 10739 26129
rect 10773 26095 10807 26129
rect 10841 26095 10875 26129
rect 10909 26095 10943 26129
rect 10977 26095 11011 26129
rect 11045 26095 11079 26129
rect 11113 26095 11147 26129
rect 11181 26095 11215 26129
rect 11249 26095 11283 26129
rect 11317 26095 11351 26129
rect 11385 26095 11419 26129
rect 11453 26095 11487 26129
rect 11521 26095 11555 26129
rect 11589 26095 11623 26129
rect 11657 26095 11691 26129
rect 11725 26095 11759 26129
rect 11793 26095 11827 26129
rect 11861 26095 11895 26129
rect 11929 26095 11963 26129
rect 11997 26095 12031 26129
rect 12065 26095 12099 26129
rect 12133 26095 12167 26129
rect 12201 26095 12235 26129
rect 12269 26095 12303 26129
rect 12337 26095 12371 26129
rect 12405 26095 12439 26129
rect 12473 26095 12507 26129
rect 12541 26095 12575 26129
rect 12609 26095 12643 26129
rect 12677 26095 12711 26129
rect 12745 26095 12779 26129
rect 12813 26095 12847 26129
rect 12881 26095 12915 26129
rect 12949 26095 12983 26129
rect 13017 26095 13051 26129
rect 13085 26095 13119 26129
rect 13153 26095 13187 26129
rect 13221 26095 13255 26129
rect 13289 26095 13323 26129
rect 13357 26095 13391 26129
rect 13425 26095 13459 26129
rect 13493 26095 13527 26129
rect 13561 26095 13595 26129
rect 13629 26095 13663 26129
rect 13697 26095 13731 26129
rect 13765 26095 13799 26129
rect 13833 26095 13867 26129
rect 13901 26095 13935 26129
rect 13969 26095 14003 26129
rect 14037 26095 14071 26129
rect 14105 26095 14139 26129
rect 14173 26095 14233 26129
rect 9877 26059 14233 26095
rect 9877 26025 9911 26059
rect 9945 26025 9980 26059
rect 10014 26025 10049 26059
rect 10083 26025 10118 26059
rect 10152 26025 10187 26059
rect 10221 26025 10256 26059
rect 10290 26025 10325 26059
rect 10359 26025 10394 26059
rect 10428 26025 10463 26059
rect 10497 26025 10532 26059
rect 10566 26025 10601 26059
rect 10635 26025 10670 26059
rect 10704 26025 10739 26059
rect 10773 26025 10807 26059
rect 10841 26025 10875 26059
rect 10909 26025 10943 26059
rect 10977 26025 11011 26059
rect 11045 26025 11079 26059
rect 11113 26025 11147 26059
rect 11181 26025 11215 26059
rect 11249 26025 11283 26059
rect 11317 26025 11351 26059
rect 11385 26025 11419 26059
rect 11453 26025 11487 26059
rect 11521 26025 11555 26059
rect 11589 26025 11623 26059
rect 11657 26025 11691 26059
rect 11725 26025 11759 26059
rect 11793 26025 11827 26059
rect 11861 26025 11895 26059
rect 11929 26025 11963 26059
rect 11997 26025 12031 26059
rect 12065 26025 12099 26059
rect 12133 26025 12167 26059
rect 12201 26025 12235 26059
rect 12269 26025 12303 26059
rect 12337 26025 12371 26059
rect 12405 26025 12439 26059
rect 12473 26025 12507 26059
rect 12541 26025 12575 26059
rect 12609 26025 12643 26059
rect 12677 26025 12711 26059
rect 12745 26025 12779 26059
rect 12813 26025 12847 26059
rect 12881 26025 12915 26059
rect 12949 26025 12983 26059
rect 13017 26025 13051 26059
rect 13085 26025 13119 26059
rect 13153 26025 13187 26059
rect 13221 26025 13255 26059
rect 13289 26025 13323 26059
rect 13357 26025 13391 26059
rect 13425 26025 13459 26059
rect 13493 26025 13527 26059
rect 13561 26025 13595 26059
rect 13629 26025 13663 26059
rect 13697 26025 13731 26059
rect 13765 26025 13799 26059
rect 13833 26025 13867 26059
rect 13901 26025 13935 26059
rect 13969 26025 14003 26059
rect 14037 26025 14071 26059
rect 14105 26025 14139 26059
rect 14173 26025 14233 26059
rect 9877 25989 14233 26025
rect 9877 25955 9911 25989
rect 9945 25955 9980 25989
rect 10014 25955 10049 25989
rect 10083 25955 10118 25989
rect 10152 25955 10187 25989
rect 10221 25955 10256 25989
rect 10290 25955 10325 25989
rect 10359 25955 10394 25989
rect 10428 25955 10463 25989
rect 10497 25955 10532 25989
rect 10566 25955 10601 25989
rect 10635 25955 10670 25989
rect 10704 25955 10739 25989
rect 10773 25955 10807 25989
rect 10841 25955 10875 25989
rect 10909 25955 10943 25989
rect 10977 25955 11011 25989
rect 11045 25955 11079 25989
rect 11113 25955 11147 25989
rect 11181 25955 11215 25989
rect 11249 25955 11283 25989
rect 11317 25955 11351 25989
rect 11385 25955 11419 25989
rect 11453 25955 11487 25989
rect 11521 25955 11555 25989
rect 11589 25955 11623 25989
rect 11657 25955 11691 25989
rect 11725 25955 11759 25989
rect 11793 25955 11827 25989
rect 11861 25955 11895 25989
rect 11929 25955 11963 25989
rect 11997 25955 12031 25989
rect 12065 25955 12099 25989
rect 12133 25955 12167 25989
rect 12201 25955 12235 25989
rect 12269 25955 12303 25989
rect 12337 25955 12371 25989
rect 12405 25955 12439 25989
rect 12473 25955 12507 25989
rect 12541 25955 12575 25989
rect 12609 25955 12643 25989
rect 12677 25955 12711 25989
rect 12745 25955 12779 25989
rect 12813 25955 12847 25989
rect 12881 25955 12915 25989
rect 12949 25955 12983 25989
rect 13017 25955 13051 25989
rect 13085 25955 13119 25989
rect 13153 25955 13187 25989
rect 13221 25955 13255 25989
rect 13289 25955 13323 25989
rect 13357 25955 13391 25989
rect 13425 25955 13459 25989
rect 13493 25955 13527 25989
rect 13561 25955 13595 25989
rect 13629 25955 13663 25989
rect 13697 25955 13731 25989
rect 13765 25955 13799 25989
rect 13833 25955 13867 25989
rect 13901 25955 13935 25989
rect 13969 25955 14003 25989
rect 14037 25955 14071 25989
rect 14105 25955 14139 25989
rect 14173 25955 14233 25989
rect 9877 25919 14233 25955
rect 9877 25885 9911 25919
rect 9945 25885 9980 25919
rect 10014 25885 10049 25919
rect 10083 25885 10118 25919
rect 10152 25885 10187 25919
rect 10221 25885 10256 25919
rect 10290 25885 10325 25919
rect 10359 25885 10394 25919
rect 10428 25885 10463 25919
rect 10497 25885 10532 25919
rect 10566 25885 10601 25919
rect 10635 25885 10670 25919
rect 10704 25885 10739 25919
rect 10773 25885 10807 25919
rect 10841 25885 10875 25919
rect 10909 25885 10943 25919
rect 10977 25885 11011 25919
rect 11045 25885 11079 25919
rect 11113 25885 11147 25919
rect 11181 25885 11215 25919
rect 11249 25885 11283 25919
rect 11317 25885 11351 25919
rect 11385 25885 11419 25919
rect 11453 25885 11487 25919
rect 11521 25885 11555 25919
rect 11589 25885 11623 25919
rect 11657 25885 11691 25919
rect 11725 25885 11759 25919
rect 11793 25885 11827 25919
rect 11861 25885 11895 25919
rect 11929 25885 11963 25919
rect 11997 25885 12031 25919
rect 12065 25885 12099 25919
rect 12133 25885 12167 25919
rect 12201 25885 12235 25919
rect 12269 25885 12303 25919
rect 12337 25885 12371 25919
rect 12405 25885 12439 25919
rect 12473 25885 12507 25919
rect 12541 25885 12575 25919
rect 12609 25885 12643 25919
rect 12677 25885 12711 25919
rect 12745 25885 12779 25919
rect 12813 25885 12847 25919
rect 12881 25885 12915 25919
rect 12949 25885 12983 25919
rect 13017 25885 13051 25919
rect 13085 25885 13119 25919
rect 13153 25885 13187 25919
rect 13221 25885 13255 25919
rect 13289 25885 13323 25919
rect 13357 25885 13391 25919
rect 13425 25885 13459 25919
rect 13493 25885 13527 25919
rect 13561 25885 13595 25919
rect 13629 25885 13663 25919
rect 13697 25885 13731 25919
rect 13765 25885 13799 25919
rect 13833 25885 13867 25919
rect 13901 25885 13935 25919
rect 13969 25885 14003 25919
rect 14037 25885 14071 25919
rect 14105 25885 14139 25919
rect 14173 25885 14233 25919
rect 9877 25849 14233 25885
rect 9877 25815 9911 25849
rect 9945 25815 9980 25849
rect 10014 25815 10049 25849
rect 10083 25815 10118 25849
rect 10152 25815 10187 25849
rect 10221 25815 10256 25849
rect 10290 25815 10325 25849
rect 10359 25815 10394 25849
rect 10428 25815 10463 25849
rect 10497 25815 10532 25849
rect 10566 25815 10601 25849
rect 10635 25815 10670 25849
rect 10704 25815 10739 25849
rect 10773 25815 10807 25849
rect 10841 25815 10875 25849
rect 10909 25815 10943 25849
rect 10977 25815 11011 25849
rect 11045 25815 11079 25849
rect 11113 25815 11147 25849
rect 11181 25815 11215 25849
rect 11249 25815 11283 25849
rect 11317 25815 11351 25849
rect 11385 25815 11419 25849
rect 11453 25815 11487 25849
rect 11521 25815 11555 25849
rect 11589 25815 11623 25849
rect 11657 25815 11691 25849
rect 11725 25815 11759 25849
rect 11793 25815 11827 25849
rect 11861 25815 11895 25849
rect 11929 25815 11963 25849
rect 11997 25815 12031 25849
rect 12065 25815 12099 25849
rect 12133 25815 12167 25849
rect 12201 25815 12235 25849
rect 12269 25815 12303 25849
rect 12337 25815 12371 25849
rect 12405 25815 12439 25849
rect 12473 25815 12507 25849
rect 12541 25815 12575 25849
rect 12609 25815 12643 25849
rect 12677 25815 12711 25849
rect 12745 25815 12779 25849
rect 12813 25815 12847 25849
rect 12881 25815 12915 25849
rect 12949 25815 12983 25849
rect 13017 25815 13051 25849
rect 13085 25815 13119 25849
rect 13153 25815 13187 25849
rect 13221 25815 13255 25849
rect 13289 25815 13323 25849
rect 13357 25815 13391 25849
rect 13425 25815 13459 25849
rect 13493 25815 13527 25849
rect 13561 25815 13595 25849
rect 13629 25815 13663 25849
rect 13697 25815 13731 25849
rect 13765 25815 13799 25849
rect 13833 25815 13867 25849
rect 13901 25815 13935 25849
rect 13969 25815 14003 25849
rect 14037 25815 14071 25849
rect 14105 25815 14139 25849
rect 14173 25815 14233 25849
rect 9877 25779 14233 25815
rect 9877 25745 9911 25779
rect 9945 25745 9980 25779
rect 10014 25745 10049 25779
rect 10083 25745 10118 25779
rect 10152 25745 10187 25779
rect 10221 25745 10256 25779
rect 10290 25745 10325 25779
rect 10359 25745 10394 25779
rect 10428 25745 10463 25779
rect 10497 25745 10532 25779
rect 10566 25745 10601 25779
rect 10635 25745 10670 25779
rect 10704 25745 10739 25779
rect 10773 25745 10807 25779
rect 10841 25745 10875 25779
rect 10909 25745 10943 25779
rect 10977 25745 11011 25779
rect 11045 25745 11079 25779
rect 11113 25745 11147 25779
rect 11181 25745 11215 25779
rect 11249 25745 11283 25779
rect 11317 25745 11351 25779
rect 11385 25745 11419 25779
rect 11453 25745 11487 25779
rect 11521 25745 11555 25779
rect 11589 25745 11623 25779
rect 11657 25745 11691 25779
rect 11725 25745 11759 25779
rect 11793 25745 11827 25779
rect 11861 25745 11895 25779
rect 11929 25745 11963 25779
rect 11997 25745 12031 25779
rect 12065 25745 12099 25779
rect 12133 25745 12167 25779
rect 12201 25745 12235 25779
rect 12269 25745 12303 25779
rect 12337 25745 12371 25779
rect 12405 25745 12439 25779
rect 12473 25745 12507 25779
rect 12541 25745 12575 25779
rect 12609 25745 12643 25779
rect 12677 25745 12711 25779
rect 12745 25745 12779 25779
rect 12813 25745 12847 25779
rect 12881 25745 12915 25779
rect 12949 25745 12983 25779
rect 13017 25745 13051 25779
rect 13085 25745 13119 25779
rect 13153 25745 13187 25779
rect 13221 25745 13255 25779
rect 13289 25745 13323 25779
rect 13357 25745 13391 25779
rect 13425 25745 13459 25779
rect 13493 25745 13527 25779
rect 13561 25745 13595 25779
rect 13629 25745 13663 25779
rect 13697 25745 13731 25779
rect 13765 25745 13799 25779
rect 13833 25745 13867 25779
rect 13901 25745 13935 25779
rect 13969 25745 14003 25779
rect 14037 25745 14071 25779
rect 14105 25745 14139 25779
rect 14173 25745 14233 25779
rect 9877 25709 14233 25745
rect 9877 25675 9911 25709
rect 9945 25675 9980 25709
rect 10014 25675 10049 25709
rect 10083 25675 10118 25709
rect 10152 25675 10187 25709
rect 10221 25675 10256 25709
rect 10290 25675 10325 25709
rect 10359 25675 10394 25709
rect 10428 25675 10463 25709
rect 10497 25675 10532 25709
rect 10566 25675 10601 25709
rect 10635 25675 10670 25709
rect 10704 25675 10739 25709
rect 10773 25675 10807 25709
rect 10841 25675 10875 25709
rect 10909 25675 10943 25709
rect 10977 25675 11011 25709
rect 11045 25675 11079 25709
rect 11113 25675 11147 25709
rect 11181 25675 11215 25709
rect 11249 25675 11283 25709
rect 11317 25675 11351 25709
rect 11385 25675 11419 25709
rect 11453 25675 11487 25709
rect 11521 25675 11555 25709
rect 11589 25675 11623 25709
rect 11657 25675 11691 25709
rect 11725 25675 11759 25709
rect 11793 25675 11827 25709
rect 11861 25675 11895 25709
rect 11929 25675 11963 25709
rect 11997 25675 12031 25709
rect 12065 25675 12099 25709
rect 12133 25675 12167 25709
rect 12201 25675 12235 25709
rect 12269 25675 12303 25709
rect 12337 25675 12371 25709
rect 12405 25675 12439 25709
rect 12473 25675 12507 25709
rect 12541 25675 12575 25709
rect 12609 25675 12643 25709
rect 12677 25675 12711 25709
rect 12745 25675 12779 25709
rect 12813 25675 12847 25709
rect 12881 25675 12915 25709
rect 12949 25675 12983 25709
rect 13017 25675 13051 25709
rect 13085 25675 13119 25709
rect 13153 25675 13187 25709
rect 13221 25675 13255 25709
rect 13289 25675 13323 25709
rect 13357 25675 13391 25709
rect 13425 25675 13459 25709
rect 13493 25675 13527 25709
rect 13561 25675 13595 25709
rect 13629 25675 13663 25709
rect 13697 25675 13731 25709
rect 13765 25675 13799 25709
rect 13833 25675 13867 25709
rect 13901 25675 13935 25709
rect 13969 25675 14003 25709
rect 14037 25675 14071 25709
rect 14105 25675 14139 25709
rect 14173 25675 14233 25709
rect 9877 25639 14233 25675
rect 9877 25605 9911 25639
rect 9945 25605 9980 25639
rect 10014 25605 10049 25639
rect 10083 25605 10118 25639
rect 10152 25605 10187 25639
rect 10221 25605 10256 25639
rect 10290 25605 10325 25639
rect 10359 25605 10394 25639
rect 10428 25605 10463 25639
rect 10497 25605 10532 25639
rect 10566 25605 10601 25639
rect 10635 25605 10670 25639
rect 10704 25605 10739 25639
rect 10773 25605 10807 25639
rect 10841 25605 10875 25639
rect 10909 25605 10943 25639
rect 10977 25605 11011 25639
rect 11045 25605 11079 25639
rect 11113 25605 11147 25639
rect 11181 25605 11215 25639
rect 11249 25605 11283 25639
rect 11317 25605 11351 25639
rect 11385 25605 11419 25639
rect 11453 25605 11487 25639
rect 11521 25605 11555 25639
rect 11589 25605 11623 25639
rect 11657 25605 11691 25639
rect 11725 25605 11759 25639
rect 11793 25605 11827 25639
rect 11861 25605 11895 25639
rect 11929 25605 11963 25639
rect 11997 25605 12031 25639
rect 12065 25605 12099 25639
rect 12133 25605 12167 25639
rect 12201 25605 12235 25639
rect 12269 25605 12303 25639
rect 12337 25605 12371 25639
rect 12405 25605 12439 25639
rect 12473 25605 12507 25639
rect 12541 25605 12575 25639
rect 12609 25605 12643 25639
rect 12677 25605 12711 25639
rect 12745 25605 12779 25639
rect 12813 25605 12847 25639
rect 12881 25605 12915 25639
rect 12949 25605 12983 25639
rect 13017 25605 13051 25639
rect 13085 25605 13119 25639
rect 13153 25605 13187 25639
rect 13221 25605 13255 25639
rect 13289 25605 13323 25639
rect 13357 25605 13391 25639
rect 13425 25605 13459 25639
rect 13493 25605 13527 25639
rect 13561 25605 13595 25639
rect 13629 25605 13663 25639
rect 13697 25605 13731 25639
rect 13765 25605 13799 25639
rect 13833 25605 13867 25639
rect 13901 25605 13935 25639
rect 13969 25605 14003 25639
rect 14037 25605 14071 25639
rect 14105 25605 14139 25639
rect 14173 25605 14233 25639
rect 9877 25569 14233 25605
rect 9877 25535 9911 25569
rect 9945 25535 9980 25569
rect 10014 25535 10049 25569
rect 10083 25535 10118 25569
rect 10152 25535 10187 25569
rect 10221 25535 10256 25569
rect 10290 25535 10325 25569
rect 10359 25535 10394 25569
rect 10428 25535 10463 25569
rect 10497 25535 10532 25569
rect 10566 25535 10601 25569
rect 10635 25535 10670 25569
rect 10704 25535 10739 25569
rect 10773 25535 10807 25569
rect 10841 25535 10875 25569
rect 10909 25535 10943 25569
rect 10977 25535 11011 25569
rect 11045 25535 11079 25569
rect 11113 25535 11147 25569
rect 11181 25535 11215 25569
rect 11249 25535 11283 25569
rect 11317 25535 11351 25569
rect 11385 25535 11419 25569
rect 11453 25535 11487 25569
rect 11521 25535 11555 25569
rect 11589 25535 11623 25569
rect 11657 25535 11691 25569
rect 11725 25535 11759 25569
rect 11793 25535 11827 25569
rect 11861 25535 11895 25569
rect 11929 25535 11963 25569
rect 11997 25535 12031 25569
rect 12065 25535 12099 25569
rect 12133 25535 12167 25569
rect 12201 25535 12235 25569
rect 12269 25535 12303 25569
rect 12337 25535 12371 25569
rect 12405 25535 12439 25569
rect 12473 25535 12507 25569
rect 12541 25535 12575 25569
rect 12609 25535 12643 25569
rect 12677 25535 12711 25569
rect 12745 25535 12779 25569
rect 12813 25535 12847 25569
rect 12881 25535 12915 25569
rect 12949 25535 12983 25569
rect 13017 25535 13051 25569
rect 13085 25535 13119 25569
rect 13153 25535 13187 25569
rect 13221 25535 13255 25569
rect 13289 25535 13323 25569
rect 13357 25535 13391 25569
rect 13425 25535 13459 25569
rect 13493 25535 13527 25569
rect 13561 25535 13595 25569
rect 13629 25535 13663 25569
rect 13697 25535 13731 25569
rect 13765 25535 13799 25569
rect 13833 25535 13867 25569
rect 13901 25535 13935 25569
rect 13969 25535 14003 25569
rect 14037 25535 14071 25569
rect 14105 25535 14139 25569
rect 14173 25535 14233 25569
rect 9877 25499 14233 25535
rect 9877 25465 9911 25499
rect 9945 25465 9980 25499
rect 10014 25465 10049 25499
rect 10083 25465 10118 25499
rect 10152 25465 10187 25499
rect 10221 25465 10256 25499
rect 10290 25465 10325 25499
rect 10359 25465 10394 25499
rect 10428 25465 10463 25499
rect 10497 25465 10532 25499
rect 10566 25465 10601 25499
rect 10635 25465 10670 25499
rect 10704 25465 10739 25499
rect 10773 25465 10807 25499
rect 10841 25465 10875 25499
rect 10909 25465 10943 25499
rect 10977 25465 11011 25499
rect 11045 25465 11079 25499
rect 11113 25465 11147 25499
rect 11181 25465 11215 25499
rect 11249 25465 11283 25499
rect 11317 25465 11351 25499
rect 11385 25465 11419 25499
rect 11453 25465 11487 25499
rect 11521 25465 11555 25499
rect 11589 25465 11623 25499
rect 11657 25465 11691 25499
rect 11725 25465 11759 25499
rect 11793 25465 11827 25499
rect 11861 25465 11895 25499
rect 11929 25465 11963 25499
rect 11997 25465 12031 25499
rect 12065 25465 12099 25499
rect 12133 25465 12167 25499
rect 12201 25465 12235 25499
rect 12269 25465 12303 25499
rect 12337 25465 12371 25499
rect 12405 25465 12439 25499
rect 12473 25465 12507 25499
rect 12541 25465 12575 25499
rect 12609 25465 12643 25499
rect 12677 25465 12711 25499
rect 12745 25465 12779 25499
rect 12813 25465 12847 25499
rect 12881 25465 12915 25499
rect 12949 25465 12983 25499
rect 13017 25465 13051 25499
rect 13085 25465 13119 25499
rect 13153 25465 13187 25499
rect 13221 25465 13255 25499
rect 13289 25465 13323 25499
rect 13357 25465 13391 25499
rect 13425 25465 13459 25499
rect 13493 25465 13527 25499
rect 13561 25465 13595 25499
rect 13629 25465 13663 25499
rect 13697 25465 13731 25499
rect 13765 25465 13799 25499
rect 13833 25465 13867 25499
rect 13901 25465 13935 25499
rect 13969 25465 14003 25499
rect 14037 25465 14071 25499
rect 14105 25465 14139 25499
rect 14173 25465 14233 25499
rect 9877 25429 14233 25465
rect 9877 25395 9911 25429
rect 9945 25395 9980 25429
rect 10014 25395 10049 25429
rect 10083 25395 10118 25429
rect 10152 25395 10187 25429
rect 10221 25395 10256 25429
rect 10290 25395 10325 25429
rect 10359 25395 10394 25429
rect 10428 25395 10463 25429
rect 10497 25395 10532 25429
rect 10566 25395 10601 25429
rect 10635 25395 10670 25429
rect 10704 25395 10739 25429
rect 10773 25395 10807 25429
rect 10841 25395 10875 25429
rect 10909 25395 10943 25429
rect 10977 25395 11011 25429
rect 11045 25395 11079 25429
rect 11113 25395 11147 25429
rect 11181 25395 11215 25429
rect 11249 25395 11283 25429
rect 11317 25395 11351 25429
rect 11385 25395 11419 25429
rect 11453 25395 11487 25429
rect 11521 25395 11555 25429
rect 11589 25395 11623 25429
rect 11657 25395 11691 25429
rect 11725 25395 11759 25429
rect 11793 25395 11827 25429
rect 11861 25395 11895 25429
rect 11929 25395 11963 25429
rect 11997 25395 12031 25429
rect 12065 25395 12099 25429
rect 12133 25395 12167 25429
rect 12201 25395 12235 25429
rect 12269 25395 12303 25429
rect 12337 25395 12371 25429
rect 12405 25395 12439 25429
rect 12473 25395 12507 25429
rect 12541 25395 12575 25429
rect 12609 25395 12643 25429
rect 12677 25395 12711 25429
rect 12745 25395 12779 25429
rect 12813 25395 12847 25429
rect 12881 25395 12915 25429
rect 12949 25395 12983 25429
rect 13017 25395 13051 25429
rect 13085 25395 13119 25429
rect 13153 25395 13187 25429
rect 13221 25395 13255 25429
rect 13289 25395 13323 25429
rect 13357 25395 13391 25429
rect 13425 25395 13459 25429
rect 13493 25395 13527 25429
rect 13561 25395 13595 25429
rect 13629 25395 13663 25429
rect 13697 25395 13731 25429
rect 13765 25395 13799 25429
rect 13833 25395 13867 25429
rect 13901 25395 13935 25429
rect 13969 25395 14003 25429
rect 14037 25395 14071 25429
rect 14105 25395 14139 25429
rect 14173 25395 14233 25429
rect 9877 25359 14233 25395
rect 9877 25325 9911 25359
rect 9945 25325 9980 25359
rect 10014 25325 10049 25359
rect 10083 25325 10118 25359
rect 10152 25325 10187 25359
rect 10221 25325 10256 25359
rect 10290 25325 10325 25359
rect 10359 25325 10394 25359
rect 10428 25325 10463 25359
rect 10497 25325 10532 25359
rect 10566 25325 10601 25359
rect 10635 25325 10670 25359
rect 10704 25325 10739 25359
rect 10773 25325 10807 25359
rect 10841 25325 10875 25359
rect 10909 25325 10943 25359
rect 10977 25325 11011 25359
rect 11045 25325 11079 25359
rect 11113 25325 11147 25359
rect 11181 25325 11215 25359
rect 11249 25325 11283 25359
rect 11317 25325 11351 25359
rect 11385 25325 11419 25359
rect 11453 25325 11487 25359
rect 11521 25325 11555 25359
rect 11589 25325 11623 25359
rect 11657 25325 11691 25359
rect 11725 25325 11759 25359
rect 11793 25325 11827 25359
rect 11861 25325 11895 25359
rect 11929 25325 11963 25359
rect 11997 25325 12031 25359
rect 12065 25325 12099 25359
rect 12133 25325 12167 25359
rect 12201 25325 12235 25359
rect 12269 25325 12303 25359
rect 12337 25325 12371 25359
rect 12405 25325 12439 25359
rect 12473 25325 12507 25359
rect 12541 25325 12575 25359
rect 12609 25325 12643 25359
rect 12677 25325 12711 25359
rect 12745 25325 12779 25359
rect 12813 25325 12847 25359
rect 12881 25325 12915 25359
rect 12949 25325 12983 25359
rect 13017 25325 13051 25359
rect 13085 25325 13119 25359
rect 13153 25325 13187 25359
rect 13221 25325 13255 25359
rect 13289 25325 13323 25359
rect 13357 25325 13391 25359
rect 13425 25325 13459 25359
rect 13493 25325 13527 25359
rect 13561 25325 13595 25359
rect 13629 25325 13663 25359
rect 13697 25325 13731 25359
rect 13765 25325 13799 25359
rect 13833 25325 13867 25359
rect 13901 25325 13935 25359
rect 13969 25325 14003 25359
rect 14037 25325 14071 25359
rect 14105 25325 14139 25359
rect 14173 25325 14233 25359
rect 9877 25289 14233 25325
rect 9877 25255 9911 25289
rect 9945 25255 9980 25289
rect 10014 25255 10049 25289
rect 10083 25255 10118 25289
rect 10152 25255 10187 25289
rect 10221 25255 10256 25289
rect 10290 25255 10325 25289
rect 10359 25255 10394 25289
rect 10428 25255 10463 25289
rect 10497 25255 10532 25289
rect 10566 25255 10601 25289
rect 10635 25255 10670 25289
rect 10704 25255 10739 25289
rect 10773 25255 10807 25289
rect 10841 25255 10875 25289
rect 10909 25255 10943 25289
rect 10977 25255 11011 25289
rect 11045 25255 11079 25289
rect 11113 25255 11147 25289
rect 11181 25255 11215 25289
rect 11249 25255 11283 25289
rect 11317 25255 11351 25289
rect 11385 25255 11419 25289
rect 11453 25255 11487 25289
rect 11521 25255 11555 25289
rect 11589 25255 11623 25289
rect 11657 25255 11691 25289
rect 11725 25255 11759 25289
rect 11793 25255 11827 25289
rect 11861 25255 11895 25289
rect 11929 25255 11963 25289
rect 11997 25255 12031 25289
rect 12065 25255 12099 25289
rect 12133 25255 12167 25289
rect 12201 25255 12235 25289
rect 12269 25255 12303 25289
rect 12337 25255 12371 25289
rect 12405 25255 12439 25289
rect 12473 25255 12507 25289
rect 12541 25255 12575 25289
rect 12609 25255 12643 25289
rect 12677 25255 12711 25289
rect 12745 25255 12779 25289
rect 12813 25255 12847 25289
rect 12881 25255 12915 25289
rect 12949 25255 12983 25289
rect 13017 25255 13051 25289
rect 13085 25255 13119 25289
rect 13153 25255 13187 25289
rect 13221 25255 13255 25289
rect 13289 25255 13323 25289
rect 13357 25255 13391 25289
rect 13425 25255 13459 25289
rect 13493 25255 13527 25289
rect 13561 25255 13595 25289
rect 13629 25255 13663 25289
rect 13697 25255 13731 25289
rect 13765 25255 13799 25289
rect 13833 25255 13867 25289
rect 13901 25255 13935 25289
rect 13969 25255 14003 25289
rect 14037 25255 14071 25289
rect 14105 25255 14139 25289
rect 14173 25255 14233 25289
rect 9877 25219 14233 25255
rect 9877 25185 9911 25219
rect 9945 25185 9980 25219
rect 10014 25185 10049 25219
rect 10083 25185 10118 25219
rect 10152 25185 10187 25219
rect 10221 25185 10256 25219
rect 10290 25185 10325 25219
rect 10359 25185 10394 25219
rect 10428 25185 10463 25219
rect 10497 25185 10532 25219
rect 10566 25185 10601 25219
rect 10635 25185 10670 25219
rect 10704 25185 10739 25219
rect 10773 25185 10807 25219
rect 10841 25185 10875 25219
rect 10909 25185 10943 25219
rect 10977 25185 11011 25219
rect 11045 25185 11079 25219
rect 11113 25185 11147 25219
rect 11181 25185 11215 25219
rect 11249 25185 11283 25219
rect 11317 25185 11351 25219
rect 11385 25185 11419 25219
rect 11453 25185 11487 25219
rect 11521 25185 11555 25219
rect 11589 25185 11623 25219
rect 11657 25185 11691 25219
rect 11725 25185 11759 25219
rect 11793 25185 11827 25219
rect 11861 25185 11895 25219
rect 11929 25185 11963 25219
rect 11997 25185 12031 25219
rect 12065 25185 12099 25219
rect 12133 25185 12167 25219
rect 12201 25185 12235 25219
rect 12269 25185 12303 25219
rect 12337 25185 12371 25219
rect 12405 25185 12439 25219
rect 12473 25185 12507 25219
rect 12541 25185 12575 25219
rect 12609 25185 12643 25219
rect 12677 25185 12711 25219
rect 12745 25185 12779 25219
rect 12813 25185 12847 25219
rect 12881 25185 12915 25219
rect 12949 25185 12983 25219
rect 13017 25185 13051 25219
rect 13085 25185 13119 25219
rect 13153 25185 13187 25219
rect 13221 25185 13255 25219
rect 13289 25185 13323 25219
rect 13357 25185 13391 25219
rect 13425 25185 13459 25219
rect 13493 25185 13527 25219
rect 13561 25185 13595 25219
rect 13629 25185 13663 25219
rect 13697 25185 13731 25219
rect 13765 25185 13799 25219
rect 13833 25185 13867 25219
rect 13901 25185 13935 25219
rect 13969 25185 14003 25219
rect 14037 25185 14071 25219
rect 14105 25185 14139 25219
rect 14173 25185 14233 25219
rect 9877 25149 14233 25185
rect 9877 25115 9911 25149
rect 9945 25115 9980 25149
rect 10014 25115 10049 25149
rect 10083 25115 10118 25149
rect 10152 25115 10187 25149
rect 10221 25115 10256 25149
rect 10290 25115 10325 25149
rect 10359 25115 10394 25149
rect 10428 25115 10463 25149
rect 10497 25115 10532 25149
rect 10566 25115 10601 25149
rect 10635 25115 10670 25149
rect 10704 25115 10739 25149
rect 10773 25115 10807 25149
rect 10841 25115 10875 25149
rect 10909 25115 10943 25149
rect 10977 25115 11011 25149
rect 11045 25115 11079 25149
rect 11113 25115 11147 25149
rect 11181 25115 11215 25149
rect 11249 25115 11283 25149
rect 11317 25115 11351 25149
rect 11385 25115 11419 25149
rect 11453 25115 11487 25149
rect 11521 25115 11555 25149
rect 11589 25115 11623 25149
rect 11657 25115 11691 25149
rect 11725 25115 11759 25149
rect 11793 25115 11827 25149
rect 11861 25115 11895 25149
rect 11929 25115 11963 25149
rect 11997 25115 12031 25149
rect 12065 25115 12099 25149
rect 12133 25115 12167 25149
rect 12201 25115 12235 25149
rect 12269 25115 12303 25149
rect 12337 25115 12371 25149
rect 12405 25115 12439 25149
rect 12473 25115 12507 25149
rect 12541 25115 12575 25149
rect 12609 25115 12643 25149
rect 12677 25115 12711 25149
rect 12745 25115 12779 25149
rect 12813 25115 12847 25149
rect 12881 25115 12915 25149
rect 12949 25115 12983 25149
rect 13017 25115 13051 25149
rect 13085 25115 13119 25149
rect 13153 25115 13187 25149
rect 13221 25115 13255 25149
rect 13289 25115 13323 25149
rect 13357 25115 13391 25149
rect 13425 25115 13459 25149
rect 13493 25115 13527 25149
rect 13561 25115 13595 25149
rect 13629 25115 13663 25149
rect 13697 25115 13731 25149
rect 13765 25115 13799 25149
rect 13833 25115 13867 25149
rect 13901 25115 13935 25149
rect 13969 25115 14003 25149
rect 14037 25115 14071 25149
rect 14105 25115 14139 25149
rect 14173 25115 14233 25149
rect 9877 25079 14233 25115
rect 9877 25045 9911 25079
rect 9945 25045 9980 25079
rect 10014 25045 10049 25079
rect 10083 25045 10118 25079
rect 10152 25045 10187 25079
rect 10221 25045 10256 25079
rect 10290 25045 10325 25079
rect 10359 25045 10394 25079
rect 10428 25045 10463 25079
rect 10497 25045 10532 25079
rect 10566 25045 10601 25079
rect 10635 25045 10670 25079
rect 10704 25045 10739 25079
rect 10773 25045 10807 25079
rect 10841 25045 10875 25079
rect 10909 25045 10943 25079
rect 10977 25045 11011 25079
rect 11045 25045 11079 25079
rect 11113 25045 11147 25079
rect 11181 25045 11215 25079
rect 11249 25045 11283 25079
rect 11317 25045 11351 25079
rect 11385 25045 11419 25079
rect 11453 25045 11487 25079
rect 11521 25045 11555 25079
rect 11589 25045 11623 25079
rect 11657 25045 11691 25079
rect 11725 25045 11759 25079
rect 11793 25045 11827 25079
rect 11861 25045 11895 25079
rect 11929 25045 11963 25079
rect 11997 25045 12031 25079
rect 12065 25045 12099 25079
rect 12133 25045 12167 25079
rect 12201 25045 12235 25079
rect 12269 25045 12303 25079
rect 12337 25045 12371 25079
rect 12405 25045 12439 25079
rect 12473 25045 12507 25079
rect 12541 25045 12575 25079
rect 12609 25045 12643 25079
rect 12677 25045 12711 25079
rect 12745 25045 12779 25079
rect 12813 25045 12847 25079
rect 12881 25045 12915 25079
rect 12949 25045 12983 25079
rect 13017 25045 13051 25079
rect 13085 25045 13119 25079
rect 13153 25045 13187 25079
rect 13221 25045 13255 25079
rect 13289 25045 13323 25079
rect 13357 25045 13391 25079
rect 13425 25045 13459 25079
rect 13493 25045 13527 25079
rect 13561 25045 13595 25079
rect 13629 25045 13663 25079
rect 13697 25045 13731 25079
rect 13765 25045 13799 25079
rect 13833 25045 13867 25079
rect 13901 25045 13935 25079
rect 13969 25045 14003 25079
rect 14037 25045 14071 25079
rect 14105 25045 14139 25079
rect 14173 25045 14233 25079
rect 9877 25009 14233 25045
rect 9877 24975 9911 25009
rect 9945 24975 9980 25009
rect 10014 24975 10049 25009
rect 10083 24975 10118 25009
rect 10152 24975 10187 25009
rect 10221 24975 10256 25009
rect 10290 24975 10325 25009
rect 10359 24975 10394 25009
rect 10428 24975 10463 25009
rect 10497 24975 10532 25009
rect 10566 24975 10601 25009
rect 10635 24975 10670 25009
rect 10704 24975 10739 25009
rect 10773 24975 10807 25009
rect 10841 24975 10875 25009
rect 10909 24975 10943 25009
rect 10977 24975 11011 25009
rect 11045 24975 11079 25009
rect 11113 24975 11147 25009
rect 11181 24975 11215 25009
rect 11249 24975 11283 25009
rect 11317 24975 11351 25009
rect 11385 24975 11419 25009
rect 11453 24975 11487 25009
rect 11521 24975 11555 25009
rect 11589 24975 11623 25009
rect 11657 24975 11691 25009
rect 11725 24975 11759 25009
rect 11793 24975 11827 25009
rect 11861 24975 11895 25009
rect 11929 24975 11963 25009
rect 11997 24975 12031 25009
rect 12065 24975 12099 25009
rect 12133 24975 12167 25009
rect 12201 24975 12235 25009
rect 12269 24975 12303 25009
rect 12337 24975 12371 25009
rect 12405 24975 12439 25009
rect 12473 24975 12507 25009
rect 12541 24975 12575 25009
rect 12609 24975 12643 25009
rect 12677 24975 12711 25009
rect 12745 24975 12779 25009
rect 12813 24975 12847 25009
rect 12881 24975 12915 25009
rect 12949 24975 12983 25009
rect 13017 24975 13051 25009
rect 13085 24975 13119 25009
rect 13153 24975 13187 25009
rect 13221 24975 13255 25009
rect 13289 24975 13323 25009
rect 13357 24975 13391 25009
rect 13425 24975 13459 25009
rect 13493 24975 13527 25009
rect 13561 24975 13595 25009
rect 13629 24975 13663 25009
rect 13697 24975 13731 25009
rect 13765 24975 13799 25009
rect 13833 24975 13867 25009
rect 13901 24975 13935 25009
rect 13969 24975 14003 25009
rect 14037 24975 14071 25009
rect 14105 24975 14139 25009
rect 14173 24975 14233 25009
rect 9877 24939 14233 24975
rect 9877 24905 9911 24939
rect 9945 24905 9980 24939
rect 10014 24905 10049 24939
rect 10083 24905 10118 24939
rect 10152 24905 10187 24939
rect 10221 24905 10256 24939
rect 10290 24905 10325 24939
rect 10359 24905 10394 24939
rect 10428 24905 10463 24939
rect 10497 24905 10532 24939
rect 10566 24905 10601 24939
rect 10635 24905 10670 24939
rect 10704 24905 10739 24939
rect 10773 24905 10807 24939
rect 10841 24905 10875 24939
rect 10909 24905 10943 24939
rect 10977 24905 11011 24939
rect 11045 24905 11079 24939
rect 11113 24905 11147 24939
rect 11181 24905 11215 24939
rect 11249 24905 11283 24939
rect 11317 24905 11351 24939
rect 11385 24905 11419 24939
rect 11453 24905 11487 24939
rect 11521 24905 11555 24939
rect 11589 24905 11623 24939
rect 11657 24905 11691 24939
rect 11725 24905 11759 24939
rect 11793 24905 11827 24939
rect 11861 24905 11895 24939
rect 11929 24905 11963 24939
rect 11997 24905 12031 24939
rect 12065 24905 12099 24939
rect 12133 24905 12167 24939
rect 12201 24905 12235 24939
rect 12269 24905 12303 24939
rect 12337 24905 12371 24939
rect 12405 24905 12439 24939
rect 12473 24905 12507 24939
rect 12541 24905 12575 24939
rect 12609 24905 12643 24939
rect 12677 24905 12711 24939
rect 12745 24905 12779 24939
rect 12813 24905 12847 24939
rect 12881 24905 12915 24939
rect 12949 24905 12983 24939
rect 13017 24905 13051 24939
rect 13085 24905 13119 24939
rect 13153 24905 13187 24939
rect 13221 24905 13255 24939
rect 13289 24905 13323 24939
rect 13357 24905 13391 24939
rect 13425 24905 13459 24939
rect 13493 24905 13527 24939
rect 13561 24905 13595 24939
rect 13629 24905 13663 24939
rect 13697 24905 13731 24939
rect 13765 24905 13799 24939
rect 13833 24905 13867 24939
rect 13901 24905 13935 24939
rect 13969 24905 14003 24939
rect 14037 24905 14071 24939
rect 14105 24905 14139 24939
rect 14173 24905 14233 24939
rect 9877 24856 14233 24905
rect 9877 24821 11232 24856
rect 13995 24831 14029 24856
rect 9877 24787 9911 24821
rect 9945 24787 9981 24821
rect 10015 24787 10051 24821
rect 10085 24787 10121 24821
rect 10155 24787 10191 24821
rect 10225 24787 10261 24821
rect 10295 24787 10331 24821
rect 10365 24787 10401 24821
rect 10435 24787 10471 24821
rect 10505 24787 10541 24821
rect 10575 24787 10611 24821
rect 10645 24787 10681 24821
rect 10715 24787 10750 24821
rect 10784 24787 10819 24821
rect 10853 24787 10888 24821
rect 10922 24787 10957 24821
rect 10991 24787 11026 24821
rect 11060 24787 11095 24821
rect 11129 24787 11164 24821
rect 11198 24787 11232 24821
rect 9877 24753 11232 24787
rect 9877 24719 9911 24753
rect 9945 24719 9981 24753
rect 10015 24719 10051 24753
rect 10085 24719 10121 24753
rect 10155 24719 10191 24753
rect 10225 24719 10261 24753
rect 10295 24719 10331 24753
rect 10365 24719 10401 24753
rect 10435 24719 10471 24753
rect 10505 24719 10541 24753
rect 10575 24719 10611 24753
rect 10645 24719 10681 24753
rect 10715 24719 10750 24753
rect 10784 24719 10819 24753
rect 10853 24719 10888 24753
rect 10922 24719 10957 24753
rect 10991 24719 11026 24753
rect 11060 24719 11095 24753
rect 11129 24719 11164 24753
rect 11198 24719 11232 24753
rect 9877 24685 11232 24719
rect 9877 24651 9911 24685
rect 9945 24651 9981 24685
rect 10015 24651 10051 24685
rect 10085 24651 10121 24685
rect 10155 24651 10191 24685
rect 10225 24651 10261 24685
rect 10295 24651 10331 24685
rect 10365 24651 10401 24685
rect 10435 24651 10471 24685
rect 10505 24651 10541 24685
rect 10575 24651 10611 24685
rect 10645 24651 10681 24685
rect 10715 24651 10750 24685
rect 10784 24651 10819 24685
rect 10853 24651 10888 24685
rect 10922 24651 10957 24685
rect 10991 24651 11026 24685
rect 11060 24651 11095 24685
rect 11129 24651 11164 24685
rect 11198 24651 11232 24685
rect 9877 24617 11232 24651
rect 9877 24583 9911 24617
rect 9945 24583 9981 24617
rect 10015 24583 10051 24617
rect 10085 24583 10121 24617
rect 10155 24583 10191 24617
rect 10225 24583 10261 24617
rect 10295 24583 10331 24617
rect 10365 24583 10401 24617
rect 10435 24583 10471 24617
rect 10505 24583 10541 24617
rect 10575 24583 10611 24617
rect 10645 24583 10681 24617
rect 10715 24583 10750 24617
rect 10784 24583 10819 24617
rect 10853 24583 10888 24617
rect 10922 24583 10957 24617
rect 10991 24583 11026 24617
rect 11060 24583 11095 24617
rect 11129 24583 11164 24617
rect 11198 24583 11232 24617
rect 9877 24549 11232 24583
rect 9877 24515 9911 24549
rect 9945 24515 9981 24549
rect 10015 24515 10051 24549
rect 10085 24515 10121 24549
rect 10155 24515 10191 24549
rect 10225 24515 10261 24549
rect 10295 24515 10331 24549
rect 10365 24515 10401 24549
rect 10435 24515 10471 24549
rect 10505 24515 10541 24549
rect 10575 24515 10611 24549
rect 10645 24515 10681 24549
rect 10715 24515 10750 24549
rect 10784 24515 10819 24549
rect 10853 24515 10888 24549
rect 10922 24515 10957 24549
rect 10991 24515 11026 24549
rect 11060 24515 11095 24549
rect 11129 24515 11164 24549
rect 11198 24515 11232 24549
rect 9877 24481 11232 24515
rect 9877 24447 9911 24481
rect 9945 24447 9981 24481
rect 10015 24447 10051 24481
rect 10085 24447 10121 24481
rect 10155 24447 10191 24481
rect 10225 24447 10261 24481
rect 10295 24447 10331 24481
rect 10365 24447 10401 24481
rect 10435 24447 10471 24481
rect 10505 24447 10541 24481
rect 10575 24447 10611 24481
rect 10645 24447 10681 24481
rect 10715 24447 10750 24481
rect 10784 24447 10819 24481
rect 10853 24447 10888 24481
rect 10922 24447 10957 24481
rect 10991 24447 11026 24481
rect 11060 24447 11095 24481
rect 11129 24447 11164 24481
rect 11198 24447 11232 24481
rect 9877 24413 11232 24447
rect 9877 24379 9911 24413
rect 9945 24379 9981 24413
rect 10015 24379 10051 24413
rect 10085 24379 10121 24413
rect 10155 24379 10191 24413
rect 10225 24379 10261 24413
rect 10295 24379 10331 24413
rect 10365 24379 10401 24413
rect 10435 24379 10471 24413
rect 10505 24379 10541 24413
rect 10575 24379 10611 24413
rect 10645 24379 10681 24413
rect 10715 24379 10750 24413
rect 10784 24379 10819 24413
rect 10853 24379 10888 24413
rect 10922 24379 10957 24413
rect 10991 24379 11026 24413
rect 11060 24379 11095 24413
rect 11129 24379 11164 24413
rect 11198 24379 11232 24413
rect 9877 24345 11232 24379
rect 14207 24347 14233 24856
rect 9877 24311 9911 24345
rect 9945 24311 9981 24345
rect 10015 24311 10051 24345
rect 10085 24311 10121 24345
rect 10155 24311 10191 24345
rect 10225 24311 10261 24345
rect 10295 24311 10331 24345
rect 10365 24311 10401 24345
rect 10435 24311 10471 24345
rect 10505 24311 10541 24345
rect 10575 24311 10611 24345
rect 10645 24311 10681 24345
rect 10715 24311 10750 24345
rect 10784 24311 10819 24345
rect 10853 24311 10888 24345
rect 10922 24311 10957 24345
rect 10991 24311 11026 24345
rect 11060 24311 11095 24345
rect 11129 24311 11164 24345
rect 11198 24311 11232 24345
rect 9877 24277 11232 24311
rect 9877 24243 9911 24277
rect 9945 24243 9981 24277
rect 10015 24243 10051 24277
rect 10085 24243 10121 24277
rect 10155 24243 10191 24277
rect 10225 24243 10261 24277
rect 10295 24243 10331 24277
rect 10365 24243 10401 24277
rect 10435 24243 10471 24277
rect 10505 24243 10541 24277
rect 10575 24243 10611 24277
rect 10645 24243 10681 24277
rect 10715 24243 10750 24277
rect 10784 24243 10819 24277
rect 10853 24243 10888 24277
rect 10922 24243 10957 24277
rect 10991 24243 11026 24277
rect 11060 24243 11095 24277
rect 11129 24243 11164 24277
rect 11198 24243 11232 24277
rect 9877 24209 11232 24243
rect 9877 24176 10825 24209
rect 9877 24142 9914 24176
rect 9948 24142 9984 24176
rect 10018 24142 10054 24176
rect 10088 24142 10124 24176
rect 10158 24142 10194 24176
rect 10228 24142 10264 24176
rect 10298 24142 10334 24176
rect 10368 24142 10404 24176
rect 10438 24142 10474 24176
rect 10508 24142 10544 24176
rect 10578 24142 10614 24176
rect 10648 24142 10684 24176
rect 10718 24142 10754 24176
rect 10788 24142 10825 24176
rect 9877 24108 10825 24142
rect 9877 24074 9914 24108
rect 9948 24074 9984 24108
rect 10018 24074 10054 24108
rect 10088 24074 10124 24108
rect 10158 24074 10194 24108
rect 10228 24074 10264 24108
rect 10298 24074 10334 24108
rect 10368 24074 10404 24108
rect 10438 24074 10474 24108
rect 10508 24074 10544 24108
rect 10578 24074 10614 24108
rect 10648 24074 10684 24108
rect 10718 24074 10754 24108
rect 10788 24074 10825 24108
rect 9877 24040 10825 24074
rect 9877 24006 9914 24040
rect 9948 24006 9984 24040
rect 10018 24006 10054 24040
rect 10088 24006 10124 24040
rect 10158 24006 10194 24040
rect 10228 24006 10264 24040
rect 10298 24006 10334 24040
rect 10368 24006 10404 24040
rect 10438 24006 10474 24040
rect 10508 24006 10544 24040
rect 10578 24006 10614 24040
rect 10648 24006 10684 24040
rect 10718 24006 10754 24040
rect 10788 24006 10825 24040
rect 9877 23971 10825 24006
rect 9877 23937 9914 23971
rect 9948 23937 9984 23971
rect 10018 23937 10054 23971
rect 10088 23937 10124 23971
rect 10158 23937 10194 23971
rect 10228 23937 10264 23971
rect 10298 23937 10334 23971
rect 10368 23937 10404 23971
rect 10438 23937 10474 23971
rect 10508 23937 10544 23971
rect 10578 23937 10614 23971
rect 10648 23937 10684 23971
rect 10718 23937 10754 23971
rect 10788 23937 10825 23971
rect 9877 23902 10825 23937
rect 9877 23868 9914 23902
rect 9948 23868 9984 23902
rect 10018 23868 10054 23902
rect 10088 23868 10124 23902
rect 10158 23868 10194 23902
rect 10228 23868 10264 23902
rect 10298 23868 10334 23902
rect 10368 23868 10404 23902
rect 10438 23868 10474 23902
rect 10508 23868 10544 23902
rect 10578 23868 10614 23902
rect 10648 23868 10684 23902
rect 10718 23868 10754 23902
rect 10788 23868 10825 23902
rect 9877 23833 10825 23868
rect 9877 23799 9914 23833
rect 9948 23799 9984 23833
rect 10018 23799 10054 23833
rect 10088 23799 10124 23833
rect 10158 23799 10194 23833
rect 10228 23799 10264 23833
rect 10298 23799 10334 23833
rect 10368 23799 10404 23833
rect 10438 23799 10474 23833
rect 10508 23799 10544 23833
rect 10578 23799 10614 23833
rect 10648 23799 10684 23833
rect 10718 23799 10754 23833
rect 10788 23799 10825 23833
rect 9877 23764 10825 23799
rect 9877 23730 9914 23764
rect 9948 23730 9984 23764
rect 10018 23730 10054 23764
rect 10088 23730 10124 23764
rect 10158 23730 10194 23764
rect 10228 23730 10264 23764
rect 10298 23730 10334 23764
rect 10368 23730 10404 23764
rect 10438 23730 10474 23764
rect 10508 23730 10544 23764
rect 10578 23730 10614 23764
rect 10648 23730 10684 23764
rect 10718 23730 10754 23764
rect 10788 23730 10825 23764
rect 9877 23695 10825 23730
rect 9877 23661 9914 23695
rect 9948 23661 9984 23695
rect 10018 23661 10054 23695
rect 10088 23661 10124 23695
rect 10158 23661 10194 23695
rect 10228 23661 10264 23695
rect 10298 23661 10334 23695
rect 10368 23661 10404 23695
rect 10438 23661 10474 23695
rect 10508 23661 10544 23695
rect 10578 23661 10614 23695
rect 10648 23661 10684 23695
rect 10718 23661 10754 23695
rect 10788 23661 10825 23695
rect 9877 23626 10825 23661
rect 9877 23592 9914 23626
rect 9948 23592 9984 23626
rect 10018 23592 10054 23626
rect 10088 23592 10124 23626
rect 10158 23592 10194 23626
rect 10228 23592 10264 23626
rect 10298 23592 10334 23626
rect 10368 23592 10404 23626
rect 10438 23592 10474 23626
rect 10508 23592 10544 23626
rect 10578 23592 10614 23626
rect 10648 23592 10684 23626
rect 10718 23592 10754 23626
rect 10788 23592 10825 23626
rect 9877 23557 10825 23592
rect 9877 23523 9914 23557
rect 9948 23523 9984 23557
rect 10018 23523 10054 23557
rect 10088 23523 10124 23557
rect 10158 23523 10194 23557
rect 10228 23523 10264 23557
rect 10298 23523 10334 23557
rect 10368 23523 10404 23557
rect 10438 23523 10474 23557
rect 10508 23523 10544 23557
rect 10578 23523 10614 23557
rect 10648 23523 10684 23557
rect 10718 23523 10754 23557
rect 10788 23523 10825 23557
rect 9877 23488 10825 23523
rect 9877 23454 9914 23488
rect 9948 23454 9984 23488
rect 10018 23454 10054 23488
rect 10088 23454 10124 23488
rect 10158 23454 10194 23488
rect 10228 23454 10264 23488
rect 10298 23454 10334 23488
rect 10368 23454 10404 23488
rect 10438 23454 10474 23488
rect 10508 23454 10544 23488
rect 10578 23454 10614 23488
rect 10648 23454 10684 23488
rect 10718 23454 10754 23488
rect 10788 23454 10825 23488
rect 9877 23419 10825 23454
rect 9877 23385 9914 23419
rect 9948 23385 9984 23419
rect 10018 23385 10054 23419
rect 10088 23385 10124 23419
rect 10158 23385 10194 23419
rect 10228 23385 10264 23419
rect 10298 23385 10334 23419
rect 10368 23385 10404 23419
rect 10438 23385 10474 23419
rect 10508 23385 10544 23419
rect 10578 23385 10614 23419
rect 10648 23385 10684 23419
rect 10718 23385 10754 23419
rect 10788 23385 10825 23419
rect 9877 23350 10825 23385
rect 9877 23316 9914 23350
rect 9948 23316 9984 23350
rect 10018 23316 10054 23350
rect 10088 23316 10124 23350
rect 10158 23316 10194 23350
rect 10228 23316 10264 23350
rect 10298 23316 10334 23350
rect 10368 23316 10404 23350
rect 10438 23316 10474 23350
rect 10508 23316 10544 23350
rect 10578 23316 10614 23350
rect 10648 23316 10684 23350
rect 10718 23316 10754 23350
rect 10788 23316 10825 23350
rect 9877 23281 10825 23316
rect 9877 23247 9914 23281
rect 9948 23247 9984 23281
rect 10018 23247 10054 23281
rect 10088 23247 10124 23281
rect 10158 23247 10194 23281
rect 10228 23247 10264 23281
rect 10298 23247 10334 23281
rect 10368 23247 10404 23281
rect 10438 23247 10474 23281
rect 10508 23247 10544 23281
rect 10578 23247 10614 23281
rect 10648 23247 10684 23281
rect 10718 23247 10754 23281
rect 10788 23247 10825 23281
rect 9877 23212 10825 23247
rect 9877 23178 9914 23212
rect 9948 23178 9984 23212
rect 10018 23178 10054 23212
rect 10088 23178 10124 23212
rect 10158 23178 10194 23212
rect 10228 23178 10264 23212
rect 10298 23178 10334 23212
rect 10368 23178 10404 23212
rect 10438 23178 10474 23212
rect 10508 23178 10544 23212
rect 10578 23178 10614 23212
rect 10648 23178 10684 23212
rect 10718 23178 10754 23212
rect 10788 23178 10825 23212
rect 9877 23143 10825 23178
rect 9877 23109 9914 23143
rect 9948 23109 9984 23143
rect 10018 23109 10054 23143
rect 10088 23109 10124 23143
rect 10158 23109 10194 23143
rect 10228 23109 10264 23143
rect 10298 23109 10334 23143
rect 10368 23109 10404 23143
rect 10438 23109 10474 23143
rect 10508 23109 10544 23143
rect 10578 23109 10614 23143
rect 10648 23109 10684 23143
rect 10718 23109 10754 23143
rect 10788 23109 10825 23143
rect 9877 23074 10825 23109
rect 9877 23040 9914 23074
rect 9948 23040 9984 23074
rect 10018 23040 10054 23074
rect 10088 23040 10124 23074
rect 10158 23040 10194 23074
rect 10228 23040 10264 23074
rect 10298 23040 10334 23074
rect 10368 23040 10404 23074
rect 10438 23040 10474 23074
rect 10508 23040 10544 23074
rect 10578 23040 10614 23074
rect 10648 23040 10684 23074
rect 10718 23040 10754 23074
rect 10788 23045 10825 23074
rect 14171 24150 14233 24347
rect 14403 24150 14429 26224
rect 14171 24115 14429 24150
rect 14171 24081 14233 24115
rect 14267 24081 14301 24115
rect 14335 24081 14369 24115
rect 14403 24081 14429 24115
rect 14171 24046 14429 24081
rect 14171 24012 14233 24046
rect 14267 24012 14301 24046
rect 14335 24012 14369 24046
rect 14403 24012 14429 24046
rect 14171 23977 14429 24012
rect 14171 23943 14233 23977
rect 14267 23943 14301 23977
rect 14335 23943 14369 23977
rect 14403 23943 14429 23977
rect 14171 23908 14429 23943
rect 14171 23874 14233 23908
rect 14267 23874 14301 23908
rect 14335 23874 14369 23908
rect 14403 23874 14429 23908
rect 14171 23839 14429 23874
rect 14171 23805 14233 23839
rect 14267 23805 14301 23839
rect 14335 23805 14369 23839
rect 14403 23805 14429 23839
rect 14171 23770 14429 23805
rect 14171 23736 14233 23770
rect 14267 23736 14301 23770
rect 14335 23736 14369 23770
rect 14403 23736 14429 23770
rect 14171 23701 14429 23736
rect 14171 23667 14233 23701
rect 14267 23667 14301 23701
rect 14335 23667 14369 23701
rect 14403 23667 14429 23701
rect 14171 23632 14429 23667
rect 14171 23598 14233 23632
rect 14267 23598 14301 23632
rect 14335 23598 14369 23632
rect 14403 23598 14429 23632
rect 14171 23563 14429 23598
rect 14171 23529 14233 23563
rect 14267 23529 14301 23563
rect 14335 23529 14369 23563
rect 14403 23529 14429 23563
rect 14171 23494 14429 23529
rect 14171 23460 14233 23494
rect 14267 23460 14301 23494
rect 14335 23460 14369 23494
rect 14403 23460 14429 23494
rect 14171 23425 14429 23460
rect 14171 23391 14233 23425
rect 14267 23391 14301 23425
rect 14335 23391 14369 23425
rect 14403 23391 14429 23425
rect 14171 23356 14429 23391
rect 14171 23322 14233 23356
rect 14267 23322 14301 23356
rect 14335 23322 14369 23356
rect 14403 23322 14429 23356
rect 14171 23287 14429 23322
rect 14171 23253 14233 23287
rect 14267 23253 14301 23287
rect 14335 23253 14369 23287
rect 14403 23253 14429 23287
rect 14171 23218 14429 23253
rect 14171 23184 14233 23218
rect 14267 23184 14301 23218
rect 14335 23184 14369 23218
rect 14403 23184 14429 23218
rect 14171 23149 14429 23184
rect 14171 23115 14233 23149
rect 14267 23115 14301 23149
rect 14335 23115 14369 23149
rect 14403 23115 14429 23149
rect 14171 23080 14429 23115
rect 14171 23046 14233 23080
rect 14267 23046 14301 23080
rect 14335 23046 14369 23080
rect 14403 23046 14429 23080
rect 14171 23045 14429 23046
rect 10788 23040 14429 23045
rect 9877 23011 14429 23040
rect 9877 23005 14233 23011
rect 9877 22971 9914 23005
rect 9948 22971 9984 23005
rect 10018 22971 10054 23005
rect 10088 22971 10124 23005
rect 10158 22971 10194 23005
rect 10228 22971 10264 23005
rect 10298 22971 10334 23005
rect 10368 22971 10404 23005
rect 10438 22971 10474 23005
rect 10508 22971 10544 23005
rect 10578 22971 10614 23005
rect 10648 22971 10684 23005
rect 10718 22971 10754 23005
rect 10788 23003 14233 23005
rect 10788 22971 10859 23003
rect 9877 22969 10859 22971
rect 10893 22969 10928 23003
rect 10962 22969 10997 23003
rect 11031 22969 11066 23003
rect 11100 22969 11135 23003
rect 11169 22969 11204 23003
rect 11238 22969 11273 23003
rect 11307 22969 11342 23003
rect 11376 22969 11411 23003
rect 11445 22969 11480 23003
rect 11514 22969 11549 23003
rect 11583 22969 11618 23003
rect 11652 22969 11687 23003
rect 11721 22969 11756 23003
rect 11790 22969 11825 23003
rect 11859 22969 11894 23003
rect 11928 22969 11963 23003
rect 11997 22969 12031 23003
rect 12065 22969 12099 23003
rect 12133 22969 12167 23003
rect 12201 22969 12235 23003
rect 12269 22969 12303 23003
rect 12337 22969 12371 23003
rect 12405 22969 12439 23003
rect 12473 22969 12507 23003
rect 12541 22969 12575 23003
rect 12609 22969 12643 23003
rect 12677 22969 12711 23003
rect 12745 22969 12779 23003
rect 12813 22969 12847 23003
rect 12881 22969 12915 23003
rect 12949 22969 12983 23003
rect 13017 22969 13051 23003
rect 13085 22969 13119 23003
rect 13153 22969 13187 23003
rect 13221 22969 13255 23003
rect 13289 22969 13323 23003
rect 13357 22969 13391 23003
rect 13425 22969 13459 23003
rect 13493 22969 13527 23003
rect 13561 22969 13595 23003
rect 13629 22969 13663 23003
rect 13697 22969 13731 23003
rect 13765 22969 13799 23003
rect 13833 22969 13867 23003
rect 13901 22998 14233 23003
rect 13901 22969 13978 22998
rect 9877 22964 13978 22969
rect 14012 22964 14048 22998
rect 14082 22964 14118 22998
rect 14152 22977 14233 22998
rect 14267 22977 14301 23011
rect 14335 22977 14369 23011
rect 14403 22977 14429 23011
rect 14152 22964 14429 22977
rect 9877 22942 14429 22964
rect 9877 22935 14233 22942
rect 9877 22901 9901 22935
rect 9935 22901 9971 22935
rect 10005 22901 10041 22935
rect 10075 22901 10111 22935
rect 10145 22901 10181 22935
rect 10215 22901 10251 22935
rect 10285 22901 10321 22935
rect 10355 22901 10391 22935
rect 10425 22901 10461 22935
rect 10495 22901 10530 22935
rect 10564 22901 10599 22935
rect 10633 22901 10668 22935
rect 10702 22901 10737 22935
rect 10771 22901 10806 22935
rect 10840 22901 10875 22935
rect 10909 22901 10944 22935
rect 10978 22901 11013 22935
rect 11047 22901 11082 22935
rect 11116 22901 11151 22935
rect 11185 22901 11220 22935
rect 11254 22901 11289 22935
rect 11323 22901 11358 22935
rect 11392 22901 11427 22935
rect 11461 22901 11496 22935
rect 11530 22901 11565 22935
rect 11599 22901 11634 22935
rect 11668 22901 11703 22935
rect 11737 22901 11772 22935
rect 11806 22901 11841 22935
rect 11875 22901 11910 22935
rect 11944 22901 11979 22935
rect 12013 22901 12048 22935
rect 12082 22901 12117 22935
rect 12151 22901 12186 22935
rect 12220 22901 12255 22935
rect 12289 22901 12324 22935
rect 12358 22901 12393 22935
rect 12427 22927 14233 22935
rect 12427 22901 12451 22927
rect 9877 22865 12451 22901
rect 9877 22831 9901 22865
rect 9935 22831 9971 22865
rect 10005 22831 10041 22865
rect 10075 22831 10111 22865
rect 10145 22831 10181 22865
rect 10215 22831 10251 22865
rect 10285 22831 10321 22865
rect 10355 22831 10391 22865
rect 10425 22831 10461 22865
rect 10495 22831 10530 22865
rect 10564 22831 10599 22865
rect 10633 22831 10668 22865
rect 10702 22831 10737 22865
rect 10771 22831 10806 22865
rect 10840 22831 10875 22865
rect 10909 22831 10944 22865
rect 10978 22831 11013 22865
rect 11047 22831 11082 22865
rect 11116 22831 11151 22865
rect 11185 22831 11220 22865
rect 11254 22831 11289 22865
rect 11323 22831 11358 22865
rect 11392 22831 11427 22865
rect 11461 22831 11496 22865
rect 11530 22831 11565 22865
rect 11599 22831 11634 22865
rect 11668 22831 11703 22865
rect 11737 22831 11772 22865
rect 11806 22831 11841 22865
rect 11875 22831 11910 22865
rect 11944 22831 11979 22865
rect 12013 22831 12048 22865
rect 12082 22831 12117 22865
rect 12151 22831 12186 22865
rect 12220 22831 12255 22865
rect 12289 22831 12324 22865
rect 12358 22831 12393 22865
rect 12427 22831 12451 22865
rect 9877 22795 12451 22831
rect 9877 22761 9901 22795
rect 9935 22761 9971 22795
rect 10005 22761 10041 22795
rect 10075 22761 10111 22795
rect 10145 22761 10181 22795
rect 10215 22761 10251 22795
rect 10285 22761 10321 22795
rect 10355 22761 10391 22795
rect 10425 22761 10461 22795
rect 10495 22761 10530 22795
rect 10564 22761 10599 22795
rect 10633 22761 10668 22795
rect 10702 22761 10737 22795
rect 10771 22761 10806 22795
rect 10840 22761 10875 22795
rect 10909 22761 10944 22795
rect 10978 22761 11013 22795
rect 11047 22761 11082 22795
rect 11116 22761 11151 22795
rect 11185 22761 11220 22795
rect 11254 22761 11289 22795
rect 11323 22761 11358 22795
rect 11392 22761 11427 22795
rect 11461 22761 11496 22795
rect 11530 22761 11565 22795
rect 11599 22761 11634 22795
rect 11668 22761 11703 22795
rect 11737 22761 11772 22795
rect 11806 22761 11841 22795
rect 11875 22761 11910 22795
rect 11944 22761 11979 22795
rect 12013 22761 12048 22795
rect 12082 22761 12117 22795
rect 12151 22761 12186 22795
rect 12220 22761 12255 22795
rect 12289 22761 12324 22795
rect 12358 22761 12393 22795
rect 12427 22761 12451 22795
rect 9877 22725 12451 22761
rect 9877 22691 9901 22725
rect 9935 22691 9971 22725
rect 10005 22691 10041 22725
rect 10075 22691 10111 22725
rect 10145 22691 10181 22725
rect 10215 22691 10251 22725
rect 10285 22691 10321 22725
rect 10355 22691 10391 22725
rect 10425 22691 10461 22725
rect 10495 22691 10530 22725
rect 10564 22691 10599 22725
rect 10633 22691 10668 22725
rect 10702 22691 10737 22725
rect 10771 22691 10806 22725
rect 10840 22691 10875 22725
rect 10909 22691 10944 22725
rect 10978 22691 11013 22725
rect 11047 22691 11082 22725
rect 11116 22691 11151 22725
rect 11185 22691 11220 22725
rect 11254 22691 11289 22725
rect 11323 22691 11358 22725
rect 11392 22691 11427 22725
rect 11461 22691 11496 22725
rect 11530 22691 11565 22725
rect 11599 22691 11634 22725
rect 11668 22691 11703 22725
rect 11737 22691 11772 22725
rect 11806 22691 11841 22725
rect 11875 22691 11910 22725
rect 11944 22691 11979 22725
rect 12013 22691 12048 22725
rect 12082 22691 12117 22725
rect 12151 22691 12186 22725
rect 12220 22691 12255 22725
rect 12289 22691 12324 22725
rect 12358 22691 12393 22725
rect 12427 22691 12451 22725
rect 9877 22655 12451 22691
rect 9877 22621 9901 22655
rect 9935 22621 9971 22655
rect 10005 22621 10041 22655
rect 10075 22621 10111 22655
rect 10145 22621 10181 22655
rect 10215 22621 10251 22655
rect 10285 22621 10321 22655
rect 10355 22621 10391 22655
rect 10425 22621 10461 22655
rect 10495 22621 10530 22655
rect 10564 22621 10599 22655
rect 10633 22621 10668 22655
rect 10702 22621 10737 22655
rect 10771 22621 10806 22655
rect 10840 22621 10875 22655
rect 10909 22621 10944 22655
rect 10978 22621 11013 22655
rect 11047 22621 11082 22655
rect 11116 22621 11151 22655
rect 11185 22621 11220 22655
rect 11254 22621 11289 22655
rect 11323 22621 11358 22655
rect 11392 22621 11427 22655
rect 11461 22621 11496 22655
rect 11530 22621 11565 22655
rect 11599 22621 11634 22655
rect 11668 22621 11703 22655
rect 11737 22621 11772 22655
rect 11806 22621 11841 22655
rect 11875 22621 11910 22655
rect 11944 22621 11979 22655
rect 12013 22621 12048 22655
rect 12082 22621 12117 22655
rect 12151 22621 12186 22655
rect 12220 22621 12255 22655
rect 12289 22621 12324 22655
rect 12358 22621 12393 22655
rect 12427 22621 12451 22655
rect 9877 22585 12451 22621
rect 9877 22551 9901 22585
rect 9935 22551 9971 22585
rect 10005 22551 10041 22585
rect 10075 22551 10111 22585
rect 10145 22551 10181 22585
rect 10215 22551 10251 22585
rect 10285 22551 10321 22585
rect 10355 22551 10391 22585
rect 10425 22551 10461 22585
rect 10495 22551 10530 22585
rect 10564 22551 10599 22585
rect 10633 22551 10668 22585
rect 10702 22551 10737 22585
rect 10771 22551 10806 22585
rect 10840 22551 10875 22585
rect 10909 22551 10944 22585
rect 10978 22551 11013 22585
rect 11047 22551 11082 22585
rect 11116 22551 11151 22585
rect 11185 22551 11220 22585
rect 11254 22551 11289 22585
rect 11323 22551 11358 22585
rect 11392 22551 11427 22585
rect 11461 22551 11496 22585
rect 11530 22551 11565 22585
rect 11599 22551 11634 22585
rect 11668 22551 11703 22585
rect 11737 22551 11772 22585
rect 11806 22551 11841 22585
rect 11875 22551 11910 22585
rect 11944 22551 11979 22585
rect 12013 22551 12048 22585
rect 12082 22551 12117 22585
rect 12151 22551 12186 22585
rect 12220 22551 12255 22585
rect 12289 22551 12324 22585
rect 12358 22551 12393 22585
rect 12427 22551 12451 22585
rect 9877 22549 12451 22551
rect 13600 22908 14233 22927
rect 14267 22908 14301 22942
rect 14335 22908 14369 22942
rect 14403 22908 14429 22942
rect 13600 22903 14429 22908
rect 13600 22869 13796 22903
rect 13830 22869 13864 22903
rect 13898 22869 13932 22903
rect 13966 22869 14000 22903
rect 14034 22869 14068 22903
rect 14102 22873 14429 22903
rect 14102 22869 14233 22873
rect 13600 22839 14233 22869
rect 14267 22839 14301 22873
rect 14335 22839 14369 22873
rect 14403 22839 14429 22873
rect 13600 22833 14429 22839
rect 13600 22799 13796 22833
rect 13830 22799 13864 22833
rect 13898 22799 13932 22833
rect 13966 22799 14000 22833
rect 14034 22799 14068 22833
rect 14102 22804 14429 22833
rect 14102 22799 14233 22804
rect 13600 22770 14233 22799
rect 14267 22770 14301 22804
rect 14335 22770 14369 22804
rect 14403 22770 14429 22804
rect 13600 22763 14429 22770
rect 13600 22729 13796 22763
rect 13830 22729 13864 22763
rect 13898 22729 13932 22763
rect 13966 22729 14000 22763
rect 14034 22729 14068 22763
rect 14102 22735 14429 22763
rect 14102 22729 14233 22735
rect 13600 22701 14233 22729
rect 14267 22701 14301 22735
rect 14335 22701 14369 22735
rect 14403 22701 14429 22735
rect 13600 22693 14429 22701
rect 13600 22659 13796 22693
rect 13830 22659 13864 22693
rect 13898 22659 13932 22693
rect 13966 22659 14000 22693
rect 14034 22659 14068 22693
rect 14102 22666 14429 22693
rect 14102 22659 14233 22666
rect 13600 22632 14233 22659
rect 14267 22632 14301 22666
rect 14335 22632 14369 22666
rect 14403 22632 14429 22666
rect 13600 22623 14429 22632
rect 13600 22589 13796 22623
rect 13830 22589 13864 22623
rect 13898 22589 13932 22623
rect 13966 22589 14000 22623
rect 14034 22589 14068 22623
rect 14102 22597 14429 22623
rect 14102 22589 14233 22597
rect 13600 22563 14233 22589
rect 14267 22563 14301 22597
rect 14335 22563 14369 22597
rect 14403 22563 14429 22597
rect 13600 22553 14429 22563
rect 13600 22519 13796 22553
rect 13830 22519 13864 22553
rect 13898 22519 13932 22553
rect 13966 22519 14000 22553
rect 14034 22519 14068 22553
rect 14102 22528 14429 22553
rect 14102 22519 14233 22528
rect 13600 22494 14233 22519
rect 14267 22494 14301 22528
rect 14335 22494 14369 22528
rect 14403 22494 14429 22528
rect 13600 22483 14429 22494
rect 13600 22449 13796 22483
rect 13830 22449 13864 22483
rect 13898 22449 13932 22483
rect 13966 22449 14000 22483
rect 14034 22449 14068 22483
rect 14102 22459 14429 22483
rect 14102 22449 14233 22459
rect 13600 22425 14233 22449
rect 14267 22425 14301 22459
rect 14335 22425 14369 22459
rect 14403 22425 14429 22459
rect 13600 22413 14429 22425
rect 13600 22379 13796 22413
rect 13830 22379 13864 22413
rect 13898 22379 13932 22413
rect 13966 22379 14000 22413
rect 14034 22379 14068 22413
rect 14102 22390 14429 22413
rect 14102 22379 14233 22390
rect 13600 22356 14233 22379
rect 14267 22356 14301 22390
rect 14335 22356 14369 22390
rect 14403 22356 14429 22390
rect 13600 22343 14429 22356
rect 13600 22309 13796 22343
rect 13830 22309 13864 22343
rect 13898 22309 13932 22343
rect 13966 22309 14000 22343
rect 14034 22309 14068 22343
rect 14102 22321 14429 22343
rect 14102 22309 14233 22321
rect 13600 22287 14233 22309
rect 14267 22287 14301 22321
rect 14335 22287 14369 22321
rect 14403 22287 14429 22321
rect 13600 22273 14429 22287
rect 13600 22239 13796 22273
rect 13830 22239 13864 22273
rect 13898 22239 13932 22273
rect 13966 22239 14000 22273
rect 14034 22239 14068 22273
rect 14102 22252 14429 22273
rect 14102 22239 14233 22252
rect 13600 22218 14233 22239
rect 14267 22218 14301 22252
rect 14335 22218 14369 22252
rect 14403 22218 14429 22252
rect 13600 22203 14429 22218
rect 13600 22169 13796 22203
rect 13830 22169 13864 22203
rect 13898 22169 13932 22203
rect 13966 22169 14000 22203
rect 14034 22169 14068 22203
rect 14102 22183 14429 22203
rect 14102 22169 14233 22183
rect 13600 22149 14233 22169
rect 14267 22149 14301 22183
rect 14335 22149 14369 22183
rect 14403 22149 14429 22183
rect 13600 22133 14429 22149
rect 13600 22099 13796 22133
rect 13830 22099 13864 22133
rect 13898 22099 13932 22133
rect 13966 22099 14000 22133
rect 14034 22099 14068 22133
rect 14102 22114 14429 22133
rect 14102 22099 14233 22114
rect 13600 22080 14233 22099
rect 14267 22080 14301 22114
rect 14335 22080 14369 22114
rect 14403 22080 14429 22114
rect 13600 22063 14429 22080
rect 13600 22049 13796 22063
rect 13769 22029 13796 22049
rect 13830 22029 13864 22063
rect 13898 22029 13932 22063
rect 13966 22029 14000 22063
rect 14034 22029 14068 22063
rect 14102 22045 14429 22063
rect 14102 22029 14233 22045
rect 13769 22011 14233 22029
rect 14267 22011 14301 22045
rect 14335 22011 14369 22045
rect 14403 22011 14429 22045
rect 13769 21993 14429 22011
rect 13769 21959 13796 21993
rect 13830 21959 13864 21993
rect 13898 21959 13932 21993
rect 13966 21959 14000 21993
rect 14034 21959 14068 21993
rect 14102 21976 14429 21993
rect 14102 21959 14233 21976
rect 13769 21942 14233 21959
rect 14267 21942 14301 21976
rect 14335 21942 14369 21976
rect 14403 21942 14429 21976
rect 13769 21923 14429 21942
rect 13769 21889 13796 21923
rect 13830 21889 13864 21923
rect 13898 21889 13932 21923
rect 13966 21889 14000 21923
rect 14034 21889 14068 21923
rect 14102 21907 14429 21923
rect 14102 21889 14233 21907
rect 13769 21873 14233 21889
rect 14267 21873 14301 21907
rect 14335 21873 14369 21907
rect 14403 21873 14429 21907
rect 13769 21853 14429 21873
rect 13769 21819 13796 21853
rect 13830 21819 13864 21853
rect 13898 21819 13932 21853
rect 13966 21819 14000 21853
rect 14034 21819 14068 21853
rect 14102 21838 14429 21853
rect 14102 21819 14233 21838
rect 13769 21804 14233 21819
rect 14267 21804 14301 21838
rect 14335 21804 14369 21838
rect 14403 21804 14429 21838
rect 13769 21783 14429 21804
rect 13769 21749 13796 21783
rect 13830 21749 13864 21783
rect 13898 21749 13932 21783
rect 13966 21749 14000 21783
rect 14034 21749 14068 21783
rect 14102 21769 14429 21783
rect 14102 21749 14233 21769
rect 13769 21735 14233 21749
rect 14267 21735 14301 21769
rect 14335 21735 14369 21769
rect 14403 21735 14429 21769
rect 13769 21713 14429 21735
rect 13769 21679 13796 21713
rect 13830 21679 13864 21713
rect 13898 21679 13932 21713
rect 13966 21679 14000 21713
rect 14034 21679 14068 21713
rect 14102 21700 14429 21713
rect 14102 21679 14233 21700
rect 13769 21666 14233 21679
rect 14267 21666 14301 21700
rect 14335 21666 14369 21700
rect 14403 21666 14429 21700
rect 13769 21643 14429 21666
rect 13769 21609 13796 21643
rect 13830 21609 13864 21643
rect 13898 21609 13932 21643
rect 13966 21609 14000 21643
rect 14034 21609 14068 21643
rect 14102 21631 14429 21643
rect 14102 21609 14233 21631
rect 13769 21597 14233 21609
rect 14267 21597 14301 21631
rect 14335 21597 14369 21631
rect 14403 21597 14429 21631
rect 13769 21573 14429 21597
rect 13769 21539 13796 21573
rect 13830 21539 13864 21573
rect 13898 21539 13932 21573
rect 13966 21539 14000 21573
rect 14034 21539 14068 21573
rect 14102 21562 14429 21573
rect 14102 21539 14233 21562
rect 13769 21528 14233 21539
rect 14267 21528 14301 21562
rect 14335 21528 14369 21562
rect 14403 21528 14429 21562
rect 13769 21503 14429 21528
rect 13769 21469 13796 21503
rect 13830 21469 13864 21503
rect 13898 21469 13932 21503
rect 13966 21469 14000 21503
rect 14034 21469 14068 21503
rect 14102 21493 14429 21503
rect 14102 21469 14233 21493
rect 13769 21459 14233 21469
rect 14267 21459 14301 21493
rect 14335 21459 14369 21493
rect 14403 21459 14429 21493
rect 13769 21445 14429 21459
rect 13601 21433 14429 21445
rect 13601 21399 13796 21433
rect 13830 21399 13864 21433
rect 13898 21399 13932 21433
rect 13966 21399 14000 21433
rect 14034 21399 14068 21433
rect 14102 21424 14429 21433
rect 14102 21399 14233 21424
rect 13601 21390 14233 21399
rect 14267 21390 14301 21424
rect 14335 21390 14369 21424
rect 14403 21390 14429 21424
rect 13601 21363 14429 21390
rect 13601 21329 13796 21363
rect 13830 21329 13864 21363
rect 13898 21329 13932 21363
rect 13966 21329 14000 21363
rect 14034 21329 14068 21363
rect 14102 21355 14429 21363
rect 14102 21329 14233 21355
rect 13601 21321 14233 21329
rect 14267 21321 14301 21355
rect 14335 21321 14369 21355
rect 14403 21321 14429 21355
rect 13601 21293 14429 21321
rect 13601 21259 13796 21293
rect 13830 21259 13864 21293
rect 13898 21259 13932 21293
rect 13966 21259 14000 21293
rect 14034 21259 14068 21293
rect 14102 21286 14429 21293
rect 14102 21259 14233 21286
rect 13601 21252 14233 21259
rect 14267 21252 14301 21286
rect 14335 21252 14369 21286
rect 14403 21252 14429 21286
rect 13601 21223 14429 21252
rect 13601 21189 13796 21223
rect 13830 21189 13864 21223
rect 13898 21189 13932 21223
rect 13966 21189 14000 21223
rect 14034 21189 14068 21223
rect 14102 21217 14429 21223
rect 14102 21189 14233 21217
rect 13601 21183 14233 21189
rect 14267 21183 14301 21217
rect 14335 21183 14369 21217
rect 14403 21183 14429 21217
rect 13601 21153 14429 21183
rect 13601 21119 13796 21153
rect 13830 21119 13864 21153
rect 13898 21119 13932 21153
rect 13966 21119 14000 21153
rect 14034 21119 14068 21153
rect 14102 21148 14429 21153
rect 14102 21119 14233 21148
rect 13601 21114 14233 21119
rect 14267 21114 14301 21148
rect 14335 21114 14369 21148
rect 14403 21114 14429 21148
rect 13601 21083 14429 21114
rect 13601 21049 13796 21083
rect 13830 21049 13864 21083
rect 13898 21049 13932 21083
rect 13966 21049 14000 21083
rect 14034 21049 14068 21083
rect 14102 21079 14429 21083
rect 14102 21049 14233 21079
rect 13601 21045 14233 21049
rect 14267 21045 14301 21079
rect 14335 21045 14369 21079
rect 14403 21045 14429 21079
rect 13601 21012 14429 21045
rect 13601 20978 13796 21012
rect 13830 20978 13864 21012
rect 13898 20978 13932 21012
rect 13966 20978 14000 21012
rect 14034 20978 14068 21012
rect 14102 21010 14429 21012
rect 14102 20978 14233 21010
rect 13601 20976 14233 20978
rect 14267 20976 14301 21010
rect 14335 20976 14369 21010
rect 14403 20976 14429 21010
rect 13601 20941 14429 20976
rect 13601 20907 13796 20941
rect 13830 20907 13864 20941
rect 13898 20907 13932 20941
rect 13966 20907 14000 20941
rect 14034 20907 14068 20941
rect 14102 20907 14233 20941
rect 14267 20907 14301 20941
rect 14335 20907 14369 20941
rect 14403 20907 14429 20941
rect 13601 20868 14429 20907
<< mvnsubdiff >>
rect 13011 30995 14268 30996
rect 13011 30927 13078 30995
rect 14200 30961 14268 30995
rect 13011 30825 13077 30927
rect 14199 30923 14268 30961
rect 14199 30893 14233 30923
rect 14131 30889 14233 30893
rect 14267 30889 14268 30923
rect 14131 30856 14268 30889
rect 14131 30825 14165 30856
rect 13011 30824 14165 30825
rect 14096 30788 14165 30824
rect 14096 26573 14097 30788
rect 9725 26572 14097 26573
rect 9725 26402 9759 26572
rect 14009 26538 14097 26572
rect 14009 26504 14165 26538
rect 14077 26470 14165 26504
rect 14077 26469 14233 26470
rect 14267 26469 14268 30856
rect 14077 26436 14268 26469
rect 14077 26402 14111 26436
rect 14145 26402 14268 26436
rect 9725 26401 14268 26402
<< psubdiffcont >>
rect 11365 1434 11399 1468
rect 11365 1359 11399 1393
rect 11365 1284 11399 1318
rect 11365 1209 11399 1243
rect 11365 1134 11399 1168
rect 11365 1058 11399 1092
rect 13381 1434 13415 1468
rect 13381 1359 13415 1393
rect 13381 1284 13415 1318
rect 13381 1209 13415 1243
rect 13381 1134 13415 1168
rect 13381 1058 13415 1092
<< nsubdiffcont >>
rect 11365 764 11399 798
rect 11365 680 11399 714
rect 11365 596 11399 630
rect 11365 512 11399 546
rect 13381 764 13415 798
rect 13381 680 13415 714
rect 13381 596 13415 630
rect 13381 512 13415 546
<< mvpsubdiffcont >>
rect 9898 35975 10884 36349
rect 10939 36314 10973 36348
rect 11008 36314 11042 36348
rect 11077 36314 11111 36348
rect 11146 36314 11180 36348
rect 11215 36314 11249 36348
rect 11284 36314 11318 36348
rect 11353 36314 11387 36348
rect 11422 36314 11456 36348
rect 11491 36314 11525 36348
rect 11560 36314 11594 36348
rect 11629 36314 11663 36348
rect 11698 36314 11732 36348
rect 11767 36314 11801 36348
rect 11836 36314 11870 36348
rect 11905 36314 11939 36348
rect 11974 36314 12008 36348
rect 12043 36314 12077 36348
rect 12112 36314 12146 36348
rect 12181 36314 12215 36348
rect 12250 36314 12284 36348
rect 12319 36314 12353 36348
rect 12388 36314 12422 36348
rect 10939 36246 10973 36280
rect 11008 36246 11042 36280
rect 11077 36246 11111 36280
rect 11146 36246 11180 36280
rect 11215 36246 11249 36280
rect 11284 36246 11318 36280
rect 11353 36246 11387 36280
rect 11422 36246 11456 36280
rect 11491 36246 11525 36280
rect 11560 36246 11594 36280
rect 11629 36246 11663 36280
rect 11698 36246 11732 36280
rect 11767 36246 11801 36280
rect 11836 36246 11870 36280
rect 11905 36246 11939 36280
rect 11974 36246 12008 36280
rect 12043 36246 12077 36280
rect 12112 36246 12146 36280
rect 12181 36246 12215 36280
rect 12250 36246 12284 36280
rect 12319 36246 12353 36280
rect 12388 36246 12422 36280
rect 10939 36178 10973 36212
rect 11008 36178 11042 36212
rect 11077 36178 11111 36212
rect 11146 36178 11180 36212
rect 11215 36178 11249 36212
rect 11284 36178 11318 36212
rect 11353 36178 11387 36212
rect 11422 36178 11456 36212
rect 11491 36178 11525 36212
rect 11560 36178 11594 36212
rect 11629 36178 11663 36212
rect 11698 36178 11732 36212
rect 11767 36178 11801 36212
rect 11836 36178 11870 36212
rect 11905 36178 11939 36212
rect 11974 36178 12008 36212
rect 12043 36178 12077 36212
rect 12112 36178 12146 36212
rect 12181 36178 12215 36212
rect 12250 36178 12284 36212
rect 12319 36178 12353 36212
rect 12388 36178 12422 36212
rect 10939 36110 10973 36144
rect 11008 36110 11042 36144
rect 11077 36110 11111 36144
rect 11146 36110 11180 36144
rect 11215 36110 11249 36144
rect 11284 36110 11318 36144
rect 11353 36110 11387 36144
rect 11422 36110 11456 36144
rect 11491 36110 11525 36144
rect 11560 36110 11594 36144
rect 11629 36110 11663 36144
rect 11698 36110 11732 36144
rect 11767 36110 11801 36144
rect 11836 36110 11870 36144
rect 11905 36110 11939 36144
rect 11974 36110 12008 36144
rect 12043 36110 12077 36144
rect 12112 36110 12146 36144
rect 12181 36110 12215 36144
rect 12250 36110 12284 36144
rect 12319 36110 12353 36144
rect 12388 36110 12422 36144
rect 10939 36042 10973 36076
rect 11008 36042 11042 36076
rect 11077 36042 11111 36076
rect 11146 36042 11180 36076
rect 11215 36042 11249 36076
rect 11284 36042 11318 36076
rect 11353 36042 11387 36076
rect 11422 36042 11456 36076
rect 11491 36042 11525 36076
rect 11560 36042 11594 36076
rect 11629 36042 11663 36076
rect 11698 36042 11732 36076
rect 11767 36042 11801 36076
rect 11836 36042 11870 36076
rect 11905 36042 11939 36076
rect 11974 36042 12008 36076
rect 12043 36042 12077 36076
rect 12112 36042 12146 36076
rect 12181 36042 12215 36076
rect 12250 36042 12284 36076
rect 12319 36042 12353 36076
rect 12388 36042 12422 36076
rect 10939 35974 10973 36008
rect 11008 35974 11042 36008
rect 11077 35974 11111 36008
rect 11146 35974 11180 36008
rect 11215 35974 11249 36008
rect 11284 35974 11318 36008
rect 11353 35974 11387 36008
rect 11422 35974 11456 36008
rect 11491 35974 11525 36008
rect 11560 35974 11594 36008
rect 11629 35974 11663 36008
rect 11698 35974 11732 36008
rect 11767 35974 11801 36008
rect 11836 35974 11870 36008
rect 11905 35974 11939 36008
rect 11974 35974 12008 36008
rect 12043 35974 12077 36008
rect 12112 35974 12146 36008
rect 12181 35974 12215 36008
rect 12250 35974 12284 36008
rect 12319 35974 12353 36008
rect 12388 35974 12422 36008
rect 9898 35906 9932 35940
rect 9966 35906 10000 35940
rect 10034 35906 10068 35940
rect 10102 35906 10136 35940
rect 10170 35906 10204 35940
rect 10238 35906 10272 35940
rect 10306 35906 10340 35940
rect 10374 35906 10408 35940
rect 10442 35906 10476 35940
rect 10510 35906 10544 35940
rect 10578 35906 10612 35940
rect 10646 35906 10680 35940
rect 10714 35906 10748 35940
rect 10782 35906 10816 35940
rect 10850 35906 10884 35940
rect 10939 35906 10973 35940
rect 11008 35906 11042 35940
rect 11077 35906 11111 35940
rect 11146 35906 11180 35940
rect 11215 35906 11249 35940
rect 11284 35906 11318 35940
rect 11353 35906 11387 35940
rect 11422 35906 11456 35940
rect 11491 35906 11525 35940
rect 11560 35906 11594 35940
rect 11629 35906 11663 35940
rect 11698 35906 11732 35940
rect 11767 35906 11801 35940
rect 11836 35906 11870 35940
rect 11905 35906 11939 35940
rect 11974 35906 12008 35940
rect 12043 35906 12077 35940
rect 12112 35906 12146 35940
rect 12181 35906 12215 35940
rect 12250 35906 12284 35940
rect 12319 35906 12353 35940
rect 12388 35906 12422 35940
rect 9898 35837 9932 35871
rect 9966 35837 10000 35871
rect 10034 35837 10068 35871
rect 10102 35837 10136 35871
rect 10170 35837 10204 35871
rect 10238 35837 10272 35871
rect 10306 35837 10340 35871
rect 10374 35837 10408 35871
rect 10442 35837 10476 35871
rect 10510 35837 10544 35871
rect 10578 35837 10612 35871
rect 10646 35837 10680 35871
rect 10714 35837 10748 35871
rect 10782 35837 10816 35871
rect 10850 35837 10884 35871
rect 10939 35838 10973 35872
rect 11008 35838 11042 35872
rect 11077 35838 11111 35872
rect 11146 35838 11180 35872
rect 11215 35838 11249 35872
rect 11284 35838 11318 35872
rect 11353 35838 11387 35872
rect 11422 35838 11456 35872
rect 11491 35838 11525 35872
rect 11560 35838 11594 35872
rect 11629 35838 11663 35872
rect 11698 35838 11732 35872
rect 11767 35838 11801 35872
rect 11836 35838 11870 35872
rect 11905 35838 11939 35872
rect 11974 35838 12008 35872
rect 12043 35838 12077 35872
rect 12112 35838 12146 35872
rect 12181 35838 12215 35872
rect 12250 35838 12284 35872
rect 12319 35838 12353 35872
rect 12388 35838 12422 35872
rect 9898 35768 9932 35802
rect 9966 35768 10000 35802
rect 10034 35768 10068 35802
rect 10102 35768 10136 35802
rect 10170 35768 10204 35802
rect 10238 35768 10272 35802
rect 10306 35768 10340 35802
rect 10374 35768 10408 35802
rect 10442 35768 10476 35802
rect 10510 35768 10544 35802
rect 10578 35768 10612 35802
rect 10646 35768 10680 35802
rect 10714 35768 10748 35802
rect 10782 35768 10816 35802
rect 10850 35768 10884 35802
rect 10939 35770 10973 35804
rect 11008 35770 11042 35804
rect 11077 35770 11111 35804
rect 11146 35770 11180 35804
rect 11215 35770 11249 35804
rect 11284 35770 11318 35804
rect 11353 35770 11387 35804
rect 11422 35770 11456 35804
rect 11491 35770 11525 35804
rect 11560 35770 11594 35804
rect 11629 35770 11663 35804
rect 11698 35770 11732 35804
rect 11767 35770 11801 35804
rect 11836 35770 11870 35804
rect 11905 35770 11939 35804
rect 11974 35770 12008 35804
rect 12043 35770 12077 35804
rect 12112 35770 12146 35804
rect 12181 35770 12215 35804
rect 12250 35770 12284 35804
rect 12319 35770 12353 35804
rect 12388 35770 12422 35804
rect 12457 35770 14395 36348
rect 13202 35599 14392 35701
rect 13202 35530 13236 35564
rect 13270 35530 13304 35564
rect 13338 35530 13372 35564
rect 13406 35530 13440 35564
rect 13474 35530 13508 35564
rect 13542 35530 13576 35564
rect 13610 35530 13644 35564
rect 13678 35530 13712 35564
rect 13746 35530 13780 35564
rect 13814 35530 13848 35564
rect 13882 35530 13916 35564
rect 13950 35530 13984 35564
rect 14018 35530 14052 35564
rect 14086 35530 14120 35564
rect 14154 35530 14188 35564
rect 14222 35530 14256 35564
rect 14290 35530 14324 35564
rect 14358 35530 14392 35564
rect 13202 35461 13236 35495
rect 13270 35461 13304 35495
rect 13338 35461 13372 35495
rect 13406 35461 13440 35495
rect 13474 35461 13508 35495
rect 13542 35461 13576 35495
rect 13610 35461 13644 35495
rect 13678 35461 13712 35495
rect 13746 35461 13780 35495
rect 13814 35461 13848 35495
rect 13882 35461 13916 35495
rect 13950 35461 13984 35495
rect 14018 35461 14052 35495
rect 14086 35461 14120 35495
rect 14154 35461 14188 35495
rect 14222 35461 14256 35495
rect 14290 35461 14324 35495
rect 14358 35461 14392 35495
rect 13202 35392 13236 35426
rect 13270 35392 13304 35426
rect 13338 35392 13372 35426
rect 13406 35392 13440 35426
rect 13474 35392 13508 35426
rect 13542 35392 13576 35426
rect 13610 35392 13644 35426
rect 13678 35392 13712 35426
rect 13746 35392 13780 35426
rect 13814 35392 13848 35426
rect 13882 35392 13916 35426
rect 13950 35392 13984 35426
rect 14018 35392 14052 35426
rect 14086 35392 14120 35426
rect 14154 35392 14188 35426
rect 14222 35392 14256 35426
rect 14290 35392 14324 35426
rect 14358 35392 14392 35426
rect 13202 35323 13236 35357
rect 13270 35323 13304 35357
rect 13338 35323 13372 35357
rect 13406 35323 13440 35357
rect 13474 35323 13508 35357
rect 13542 35323 13576 35357
rect 13610 35323 13644 35357
rect 13678 35323 13712 35357
rect 13746 35323 13780 35357
rect 13814 35323 13848 35357
rect 13882 35323 13916 35357
rect 13950 35323 13984 35357
rect 14018 35323 14052 35357
rect 14086 35323 14120 35357
rect 14154 35323 14188 35357
rect 14222 35323 14256 35357
rect 14290 35323 14324 35357
rect 14358 35323 14392 35357
rect 13202 35254 13236 35288
rect 13270 35254 13304 35288
rect 13338 35254 13372 35288
rect 13406 35254 13440 35288
rect 13474 35254 13508 35288
rect 13542 35254 13576 35288
rect 13610 35254 13644 35288
rect 13678 35254 13712 35288
rect 13746 35254 13780 35288
rect 13814 35254 13848 35288
rect 13882 35254 13916 35288
rect 13950 35254 13984 35288
rect 14018 35254 14052 35288
rect 14086 35254 14120 35288
rect 14154 35254 14188 35288
rect 14222 35254 14256 35288
rect 14290 35254 14324 35288
rect 14358 35254 14392 35288
rect 13202 35185 13236 35219
rect 13270 35185 13304 35219
rect 13338 35185 13372 35219
rect 13406 35185 13440 35219
rect 13474 35185 13508 35219
rect 13542 35185 13576 35219
rect 13610 35185 13644 35219
rect 13678 35185 13712 35219
rect 13746 35185 13780 35219
rect 13814 35185 13848 35219
rect 13882 35185 13916 35219
rect 13950 35185 13984 35219
rect 14018 35185 14052 35219
rect 14086 35185 14120 35219
rect 14154 35185 14188 35219
rect 14222 35185 14256 35219
rect 14290 35185 14324 35219
rect 14358 35185 14392 35219
rect 13202 35116 13236 35150
rect 13270 35116 13304 35150
rect 13338 35116 13372 35150
rect 13406 35116 13440 35150
rect 13474 35116 13508 35150
rect 13542 35116 13576 35150
rect 13610 35116 13644 35150
rect 13678 35116 13712 35150
rect 13746 35116 13780 35150
rect 13814 35116 13848 35150
rect 13882 35116 13916 35150
rect 13950 35116 13984 35150
rect 14018 35116 14052 35150
rect 14086 35116 14120 35150
rect 14154 35116 14188 35150
rect 14222 35116 14256 35150
rect 14290 35116 14324 35150
rect 14358 35116 14392 35150
rect 13202 35047 13236 35081
rect 13270 35047 13304 35081
rect 13338 35047 13372 35081
rect 13406 35047 13440 35081
rect 13474 35047 13508 35081
rect 13542 35047 13576 35081
rect 13610 35047 13644 35081
rect 13678 35047 13712 35081
rect 13746 35047 13780 35081
rect 13814 35047 13848 35081
rect 13882 35047 13916 35081
rect 13950 35047 13984 35081
rect 14018 35047 14052 35081
rect 14086 35047 14120 35081
rect 14154 35047 14188 35081
rect 14222 35047 14256 35081
rect 14290 35047 14324 35081
rect 14358 35047 14392 35081
rect 13202 34978 13236 35012
rect 13270 34978 13304 35012
rect 13338 34978 13372 35012
rect 13406 34978 13440 35012
rect 13474 34978 13508 35012
rect 13542 34978 13576 35012
rect 13610 34978 13644 35012
rect 13678 34978 13712 35012
rect 13746 34978 13780 35012
rect 13814 34978 13848 35012
rect 13882 34978 13916 35012
rect 13950 34978 13984 35012
rect 14018 34978 14052 35012
rect 14086 34978 14120 35012
rect 14154 34978 14188 35012
rect 14222 34978 14256 35012
rect 14290 34978 14324 35012
rect 14358 34978 14392 35012
rect 13202 34909 13236 34943
rect 13270 34909 13304 34943
rect 13338 34909 13372 34943
rect 13406 34909 13440 34943
rect 13474 34909 13508 34943
rect 13542 34909 13576 34943
rect 13610 34909 13644 34943
rect 13678 34909 13712 34943
rect 13746 34909 13780 34943
rect 13814 34909 13848 34943
rect 13882 34909 13916 34943
rect 13950 34909 13984 34943
rect 14018 34909 14052 34943
rect 14086 34909 14120 34943
rect 14154 34909 14188 34943
rect 14222 34909 14256 34943
rect 14290 34909 14324 34943
rect 14358 34909 14392 34943
rect 13202 34840 13236 34874
rect 13270 34840 13304 34874
rect 13338 34840 13372 34874
rect 13406 34840 13440 34874
rect 13474 34840 13508 34874
rect 13542 34840 13576 34874
rect 13610 34840 13644 34874
rect 13678 34840 13712 34874
rect 13746 34840 13780 34874
rect 13814 34840 13848 34874
rect 13882 34840 13916 34874
rect 13950 34840 13984 34874
rect 14018 34840 14052 34874
rect 14086 34840 14120 34874
rect 14154 34840 14188 34874
rect 14222 34840 14256 34874
rect 14290 34840 14324 34874
rect 14358 34840 14392 34874
rect 13202 34771 13236 34805
rect 13270 34771 13304 34805
rect 13338 34771 13372 34805
rect 13406 34771 13440 34805
rect 13474 34771 13508 34805
rect 13542 34771 13576 34805
rect 13610 34771 13644 34805
rect 13678 34771 13712 34805
rect 13746 34771 13780 34805
rect 13814 34771 13848 34805
rect 13882 34771 13916 34805
rect 13950 34771 13984 34805
rect 14018 34771 14052 34805
rect 14086 34771 14120 34805
rect 14154 34771 14188 34805
rect 14222 34771 14256 34805
rect 14290 34771 14324 34805
rect 14358 34771 14392 34805
rect 13202 34702 13236 34736
rect 13270 34702 13304 34736
rect 13338 34702 13372 34736
rect 13406 34702 13440 34736
rect 13474 34702 13508 34736
rect 13542 34702 13576 34736
rect 13610 34702 13644 34736
rect 13678 34702 13712 34736
rect 13746 34702 13780 34736
rect 13814 34702 13848 34736
rect 13882 34702 13916 34736
rect 13950 34702 13984 34736
rect 14018 34702 14052 34736
rect 14086 34702 14120 34736
rect 14154 34702 14188 34736
rect 14222 34702 14256 34736
rect 14290 34702 14324 34736
rect 14358 34702 14392 34736
rect 13202 34633 13236 34667
rect 13270 34633 13304 34667
rect 13338 34633 13372 34667
rect 13406 34633 13440 34667
rect 13474 34633 13508 34667
rect 13542 34633 13576 34667
rect 13610 34633 13644 34667
rect 13678 34633 13712 34667
rect 13746 34633 13780 34667
rect 13814 34633 13848 34667
rect 13882 34633 13916 34667
rect 13950 34633 13984 34667
rect 14018 34633 14052 34667
rect 14086 34633 14120 34667
rect 14154 34633 14188 34667
rect 14222 34633 14256 34667
rect 14290 34633 14324 34667
rect 14358 34633 14392 34667
rect 13202 34564 13236 34598
rect 13270 34564 13304 34598
rect 13338 34564 13372 34598
rect 13406 34564 13440 34598
rect 13474 34564 13508 34598
rect 13542 34564 13576 34598
rect 13610 34564 13644 34598
rect 13678 34564 13712 34598
rect 13746 34564 13780 34598
rect 13814 34564 13848 34598
rect 13882 34564 13916 34598
rect 13950 34564 13984 34598
rect 14018 34564 14052 34598
rect 14086 34564 14120 34598
rect 14154 34564 14188 34598
rect 14222 34564 14256 34598
rect 14290 34564 14324 34598
rect 14358 34564 14392 34598
rect 13202 34495 13236 34529
rect 13270 34495 13304 34529
rect 13338 34495 13372 34529
rect 13406 34495 13440 34529
rect 13474 34495 13508 34529
rect 13542 34495 13576 34529
rect 13610 34495 13644 34529
rect 13678 34495 13712 34529
rect 13746 34495 13780 34529
rect 13814 34495 13848 34529
rect 13882 34495 13916 34529
rect 13950 34495 13984 34529
rect 14018 34495 14052 34529
rect 14086 34495 14120 34529
rect 14154 34495 14188 34529
rect 14222 34495 14256 34529
rect 14290 34495 14324 34529
rect 14358 34495 14392 34529
rect 13202 34426 13236 34460
rect 13270 34426 13304 34460
rect 13338 34426 13372 34460
rect 13406 34426 13440 34460
rect 13474 34426 13508 34460
rect 13542 34426 13576 34460
rect 13610 34426 13644 34460
rect 13678 34426 13712 34460
rect 13746 34426 13780 34460
rect 13814 34426 13848 34460
rect 13882 34426 13916 34460
rect 13950 34426 13984 34460
rect 14018 34426 14052 34460
rect 14086 34426 14120 34460
rect 14154 34426 14188 34460
rect 14222 34426 14256 34460
rect 14290 34426 14324 34460
rect 14358 34426 14392 34460
rect 13202 34357 13236 34391
rect 13270 34357 13304 34391
rect 13338 34357 13372 34391
rect 13406 34357 13440 34391
rect 13474 34357 13508 34391
rect 13542 34357 13576 34391
rect 13610 34357 13644 34391
rect 13678 34357 13712 34391
rect 13746 34357 13780 34391
rect 13814 34357 13848 34391
rect 13882 34357 13916 34391
rect 13950 34357 13984 34391
rect 14018 34357 14052 34391
rect 14086 34357 14120 34391
rect 14154 34357 14188 34391
rect 14222 34357 14256 34391
rect 14290 34357 14324 34391
rect 14358 34357 14392 34391
rect 13202 34288 13236 34322
rect 13270 34288 13304 34322
rect 13338 34288 13372 34322
rect 13406 34288 13440 34322
rect 13474 34288 13508 34322
rect 13542 34288 13576 34322
rect 13610 34288 13644 34322
rect 13678 34288 13712 34322
rect 13746 34288 13780 34322
rect 13814 34288 13848 34322
rect 13882 34288 13916 34322
rect 13950 34288 13984 34322
rect 14018 34288 14052 34322
rect 14086 34288 14120 34322
rect 14154 34288 14188 34322
rect 14222 34288 14256 34322
rect 14290 34288 14324 34322
rect 14358 34288 14392 34322
rect 13202 34219 13236 34253
rect 13270 34219 13304 34253
rect 13338 34219 13372 34253
rect 13406 34219 13440 34253
rect 13474 34219 13508 34253
rect 13542 34219 13576 34253
rect 13610 34219 13644 34253
rect 13678 34219 13712 34253
rect 13746 34219 13780 34253
rect 13814 34219 13848 34253
rect 13882 34219 13916 34253
rect 13950 34219 13984 34253
rect 14018 34219 14052 34253
rect 14086 34219 14120 34253
rect 14154 34219 14188 34253
rect 14222 34219 14256 34253
rect 14290 34219 14324 34253
rect 14358 34219 14392 34253
rect 13202 34150 13236 34184
rect 13270 34150 13304 34184
rect 13338 34150 13372 34184
rect 13406 34150 13440 34184
rect 13474 34150 13508 34184
rect 13542 34150 13576 34184
rect 13610 34150 13644 34184
rect 13678 34150 13712 34184
rect 13746 34150 13780 34184
rect 13814 34150 13848 34184
rect 13882 34150 13916 34184
rect 13950 34150 13984 34184
rect 14018 34150 14052 34184
rect 14086 34150 14120 34184
rect 14154 34150 14188 34184
rect 14222 34150 14256 34184
rect 14290 34150 14324 34184
rect 14358 34150 14392 34184
rect 13202 34081 13236 34115
rect 13270 34081 13304 34115
rect 13338 34081 13372 34115
rect 13406 34081 13440 34115
rect 13474 34081 13508 34115
rect 13542 34081 13576 34115
rect 13610 34081 13644 34115
rect 13678 34081 13712 34115
rect 13746 34081 13780 34115
rect 13814 34081 13848 34115
rect 13882 34081 13916 34115
rect 13950 34081 13984 34115
rect 14018 34081 14052 34115
rect 14086 34081 14120 34115
rect 14154 34081 14188 34115
rect 14222 34081 14256 34115
rect 14290 34081 14324 34115
rect 14358 34081 14392 34115
rect 13202 34012 13236 34046
rect 13270 34012 13304 34046
rect 13338 34012 13372 34046
rect 13406 34012 13440 34046
rect 13474 34012 13508 34046
rect 13542 34012 13576 34046
rect 13610 34012 13644 34046
rect 13678 34012 13712 34046
rect 13746 34012 13780 34046
rect 13814 34012 13848 34046
rect 13882 34012 13916 34046
rect 13950 34012 13984 34046
rect 14018 34012 14052 34046
rect 14086 34012 14120 34046
rect 14154 34012 14188 34046
rect 14222 34012 14256 34046
rect 14290 34012 14324 34046
rect 14358 34012 14392 34046
rect 13202 33943 13236 33977
rect 13270 33943 13304 33977
rect 13338 33943 13372 33977
rect 13406 33943 13440 33977
rect 13474 33943 13508 33977
rect 13542 33943 13576 33977
rect 13610 33943 13644 33977
rect 13678 33943 13712 33977
rect 13746 33943 13780 33977
rect 13814 33943 13848 33977
rect 13882 33943 13916 33977
rect 13950 33943 13984 33977
rect 14018 33943 14052 33977
rect 14086 33943 14120 33977
rect 14154 33943 14188 33977
rect 14222 33943 14256 33977
rect 14290 33943 14324 33977
rect 14358 33943 14392 33977
rect 13202 33874 13236 33908
rect 13270 33874 13304 33908
rect 13338 33874 13372 33908
rect 13406 33874 13440 33908
rect 13474 33874 13508 33908
rect 13542 33874 13576 33908
rect 13610 33874 13644 33908
rect 13678 33874 13712 33908
rect 13746 33874 13780 33908
rect 13814 33874 13848 33908
rect 13882 33874 13916 33908
rect 13950 33874 13984 33908
rect 14018 33874 14052 33908
rect 14086 33874 14120 33908
rect 14154 33874 14188 33908
rect 14222 33874 14256 33908
rect 14290 33874 14324 33908
rect 14358 33874 14392 33908
rect 13202 33805 13236 33839
rect 13270 33805 13304 33839
rect 13338 33805 13372 33839
rect 13406 33805 13440 33839
rect 13474 33805 13508 33839
rect 13542 33805 13576 33839
rect 13610 33805 13644 33839
rect 13678 33805 13712 33839
rect 13746 33805 13780 33839
rect 13814 33805 13848 33839
rect 13882 33805 13916 33839
rect 13950 33805 13984 33839
rect 14018 33805 14052 33839
rect 14086 33805 14120 33839
rect 14154 33805 14188 33839
rect 14222 33805 14256 33839
rect 14290 33805 14324 33839
rect 14358 33805 14392 33839
rect 13202 33736 13236 33770
rect 13270 33736 13304 33770
rect 13338 33736 13372 33770
rect 13406 33736 13440 33770
rect 13474 33736 13508 33770
rect 13542 33736 13576 33770
rect 13610 33736 13644 33770
rect 13678 33736 13712 33770
rect 13746 33736 13780 33770
rect 13814 33736 13848 33770
rect 13882 33736 13916 33770
rect 13950 33736 13984 33770
rect 14018 33736 14052 33770
rect 14086 33736 14120 33770
rect 14154 33736 14188 33770
rect 14222 33736 14256 33770
rect 14290 33736 14324 33770
rect 14358 33736 14392 33770
rect 13202 33667 13236 33701
rect 13270 33667 13304 33701
rect 13338 33667 13372 33701
rect 13406 33667 13440 33701
rect 13474 33667 13508 33701
rect 13542 33667 13576 33701
rect 13610 33667 13644 33701
rect 13678 33667 13712 33701
rect 13746 33667 13780 33701
rect 13814 33667 13848 33701
rect 13882 33667 13916 33701
rect 13950 33667 13984 33701
rect 14018 33667 14052 33701
rect 14086 33667 14120 33701
rect 14154 33667 14188 33701
rect 14222 33667 14256 33701
rect 14290 33667 14324 33701
rect 14358 33667 14392 33701
rect 13202 33598 13236 33632
rect 13270 33598 13304 33632
rect 13338 33598 13372 33632
rect 13406 33598 13440 33632
rect 13474 33598 13508 33632
rect 13542 33598 13576 33632
rect 13610 33598 13644 33632
rect 13678 33598 13712 33632
rect 13746 33598 13780 33632
rect 13814 33598 13848 33632
rect 13882 33598 13916 33632
rect 13950 33598 13984 33632
rect 14018 33598 14052 33632
rect 14086 33598 14120 33632
rect 14154 33598 14188 33632
rect 14222 33598 14256 33632
rect 14290 33598 14324 33632
rect 14358 33598 14392 33632
rect 13202 33529 13236 33563
rect 13270 33529 13304 33563
rect 13338 33529 13372 33563
rect 13406 33529 13440 33563
rect 13474 33529 13508 33563
rect 13542 33529 13576 33563
rect 13610 33529 13644 33563
rect 13678 33529 13712 33563
rect 13746 33529 13780 33563
rect 13814 33529 13848 33563
rect 13882 33529 13916 33563
rect 13950 33529 13984 33563
rect 14018 33529 14052 33563
rect 14086 33529 14120 33563
rect 14154 33529 14188 33563
rect 14222 33529 14256 33563
rect 14290 33529 14324 33563
rect 14358 33529 14392 33563
rect 13202 33460 13236 33494
rect 13270 33460 13304 33494
rect 13338 33460 13372 33494
rect 13406 33460 13440 33494
rect 13474 33460 13508 33494
rect 13542 33460 13576 33494
rect 13610 33460 13644 33494
rect 13678 33460 13712 33494
rect 13746 33460 13780 33494
rect 13814 33460 13848 33494
rect 13882 33460 13916 33494
rect 13950 33460 13984 33494
rect 14018 33460 14052 33494
rect 14086 33460 14120 33494
rect 14154 33460 14188 33494
rect 14222 33460 14256 33494
rect 14290 33460 14324 33494
rect 14358 33460 14392 33494
rect 13202 33391 13236 33425
rect 13270 33391 13304 33425
rect 13338 33391 13372 33425
rect 13406 33391 13440 33425
rect 13474 33391 13508 33425
rect 13542 33391 13576 33425
rect 13610 33391 13644 33425
rect 13678 33391 13712 33425
rect 13746 33391 13780 33425
rect 13814 33391 13848 33425
rect 13882 33391 13916 33425
rect 13950 33391 13984 33425
rect 14018 33391 14052 33425
rect 14086 33391 14120 33425
rect 14154 33391 14188 33425
rect 14222 33391 14256 33425
rect 14290 33391 14324 33425
rect 14358 33391 14392 33425
rect 13202 33322 13236 33356
rect 13270 33322 13304 33356
rect 13338 33322 13372 33356
rect 13406 33322 13440 33356
rect 13474 33322 13508 33356
rect 13542 33322 13576 33356
rect 13610 33322 13644 33356
rect 13678 33322 13712 33356
rect 13746 33322 13780 33356
rect 13814 33322 13848 33356
rect 13882 33322 13916 33356
rect 13950 33322 13984 33356
rect 14018 33322 14052 33356
rect 14086 33322 14120 33356
rect 14154 33322 14188 33356
rect 14222 33322 14256 33356
rect 14290 33322 14324 33356
rect 14358 33322 14392 33356
rect 13202 33253 13236 33287
rect 13270 33253 13304 33287
rect 13338 33253 13372 33287
rect 13406 33253 13440 33287
rect 13474 33253 13508 33287
rect 13542 33253 13576 33287
rect 13610 33253 13644 33287
rect 13678 33253 13712 33287
rect 13746 33253 13780 33287
rect 13814 33253 13848 33287
rect 13882 33253 13916 33287
rect 13950 33253 13984 33287
rect 14018 33253 14052 33287
rect 14086 33253 14120 33287
rect 14154 33253 14188 33287
rect 14222 33253 14256 33287
rect 14290 33253 14324 33287
rect 14358 33253 14392 33287
rect 13202 33184 13236 33218
rect 13270 33184 13304 33218
rect 13338 33184 13372 33218
rect 13406 33184 13440 33218
rect 13474 33184 13508 33218
rect 13542 33184 13576 33218
rect 13610 33184 13644 33218
rect 13678 33184 13712 33218
rect 13746 33184 13780 33218
rect 13814 33184 13848 33218
rect 13882 33184 13916 33218
rect 13950 33184 13984 33218
rect 14018 33184 14052 33218
rect 14086 33184 14120 33218
rect 14154 33184 14188 33218
rect 14222 33184 14256 33218
rect 14290 33184 14324 33218
rect 14358 33184 14392 33218
rect 13202 33115 13236 33149
rect 13270 33115 13304 33149
rect 13338 33115 13372 33149
rect 13406 33115 13440 33149
rect 13474 33115 13508 33149
rect 13542 33115 13576 33149
rect 13610 33115 13644 33149
rect 13678 33115 13712 33149
rect 13746 33115 13780 33149
rect 13814 33115 13848 33149
rect 13882 33115 13916 33149
rect 13950 33115 13984 33149
rect 14018 33115 14052 33149
rect 14086 33115 14120 33149
rect 14154 33115 14188 33149
rect 14222 33115 14256 33149
rect 14290 33115 14324 33149
rect 14358 33115 14392 33149
rect 13202 33046 13236 33080
rect 13270 33046 13304 33080
rect 13338 33046 13372 33080
rect 13406 33046 13440 33080
rect 13474 33046 13508 33080
rect 13542 33046 13576 33080
rect 13610 33046 13644 33080
rect 13678 33046 13712 33080
rect 13746 33046 13780 33080
rect 13814 33046 13848 33080
rect 13882 33046 13916 33080
rect 13950 33046 13984 33080
rect 14018 33046 14052 33080
rect 14086 33046 14120 33080
rect 14154 33046 14188 33080
rect 14222 33046 14256 33080
rect 14290 33046 14324 33080
rect 14358 33046 14392 33080
rect 13202 32977 13236 33011
rect 13270 32977 13304 33011
rect 13338 32977 13372 33011
rect 13406 32977 13440 33011
rect 13474 32977 13508 33011
rect 13542 32977 13576 33011
rect 13610 32977 13644 33011
rect 13678 32977 13712 33011
rect 13746 32977 13780 33011
rect 13814 32977 13848 33011
rect 13882 32977 13916 33011
rect 13950 32977 13984 33011
rect 14018 32977 14052 33011
rect 14086 32977 14120 33011
rect 14154 32977 14188 33011
rect 14222 32977 14256 33011
rect 14290 32977 14324 33011
rect 14358 32977 14392 33011
rect 13202 32908 13236 32942
rect 13270 32908 13304 32942
rect 13338 32908 13372 32942
rect 13406 32908 13440 32942
rect 13474 32908 13508 32942
rect 13542 32908 13576 32942
rect 13610 32908 13644 32942
rect 13678 32908 13712 32942
rect 13746 32908 13780 32942
rect 13814 32908 13848 32942
rect 13882 32908 13916 32942
rect 13950 32908 13984 32942
rect 14018 32908 14052 32942
rect 14086 32908 14120 32942
rect 14154 32908 14188 32942
rect 14222 32908 14256 32942
rect 14290 32908 14324 32942
rect 14358 32908 14392 32942
rect 13202 32839 13236 32873
rect 13270 32839 13304 32873
rect 13338 32839 13372 32873
rect 13406 32839 13440 32873
rect 13474 32839 13508 32873
rect 13542 32839 13576 32873
rect 13610 32839 13644 32873
rect 13678 32839 13712 32873
rect 13746 32839 13780 32873
rect 13814 32839 13848 32873
rect 13882 32839 13916 32873
rect 13950 32839 13984 32873
rect 14018 32839 14052 32873
rect 14086 32839 14120 32873
rect 14154 32839 14188 32873
rect 14222 32839 14256 32873
rect 14290 32839 14324 32873
rect 14358 32839 14392 32873
rect 13202 32770 13236 32804
rect 13270 32770 13304 32804
rect 13338 32770 13372 32804
rect 13406 32770 13440 32804
rect 13474 32770 13508 32804
rect 13542 32770 13576 32804
rect 13610 32770 13644 32804
rect 13678 32770 13712 32804
rect 13746 32770 13780 32804
rect 13814 32770 13848 32804
rect 13882 32770 13916 32804
rect 13950 32770 13984 32804
rect 14018 32770 14052 32804
rect 14086 32770 14120 32804
rect 14154 32770 14188 32804
rect 14222 32770 14256 32804
rect 14290 32770 14324 32804
rect 14358 32770 14392 32804
rect 13202 32701 13236 32735
rect 13270 32701 13304 32735
rect 13338 32701 13372 32735
rect 13406 32701 13440 32735
rect 13474 32701 13508 32735
rect 13542 32701 13576 32735
rect 13610 32701 13644 32735
rect 13678 32701 13712 32735
rect 13746 32701 13780 32735
rect 13814 32701 13848 32735
rect 13882 32701 13916 32735
rect 13950 32701 13984 32735
rect 14018 32701 14052 32735
rect 14086 32701 14120 32735
rect 14154 32701 14188 32735
rect 14222 32701 14256 32735
rect 14290 32701 14324 32735
rect 14358 32701 14392 32735
rect 13202 32632 13236 32666
rect 13270 32632 13304 32666
rect 13338 32632 13372 32666
rect 13406 32632 13440 32666
rect 13474 32632 13508 32666
rect 13542 32632 13576 32666
rect 13610 32632 13644 32666
rect 13678 32632 13712 32666
rect 13746 32632 13780 32666
rect 13814 32632 13848 32666
rect 13882 32632 13916 32666
rect 13950 32632 13984 32666
rect 14018 32632 14052 32666
rect 14086 32632 14120 32666
rect 14154 32632 14188 32666
rect 14222 32632 14256 32666
rect 14290 32632 14324 32666
rect 14358 32632 14392 32666
rect 13202 32563 13236 32597
rect 13270 32563 13304 32597
rect 13338 32563 13372 32597
rect 13406 32563 13440 32597
rect 13474 32563 13508 32597
rect 13542 32563 13576 32597
rect 13610 32563 13644 32597
rect 13678 32563 13712 32597
rect 13746 32563 13780 32597
rect 13814 32563 13848 32597
rect 13882 32563 13916 32597
rect 13950 32563 13984 32597
rect 14018 32563 14052 32597
rect 14086 32563 14120 32597
rect 14154 32563 14188 32597
rect 14222 32563 14256 32597
rect 14290 32563 14324 32597
rect 14358 32563 14392 32597
rect 13202 32494 13236 32528
rect 13270 32494 13304 32528
rect 13338 32494 13372 32528
rect 13406 32494 13440 32528
rect 13474 32494 13508 32528
rect 13542 32494 13576 32528
rect 13610 32494 13644 32528
rect 13678 32494 13712 32528
rect 13746 32494 13780 32528
rect 13814 32494 13848 32528
rect 13882 32494 13916 32528
rect 13950 32494 13984 32528
rect 14018 32494 14052 32528
rect 14086 32494 14120 32528
rect 14154 32494 14188 32528
rect 14222 32494 14256 32528
rect 14290 32494 14324 32528
rect 14358 32494 14392 32528
rect 13202 32425 13236 32459
rect 13270 32425 13304 32459
rect 13338 32425 13372 32459
rect 13406 32425 13440 32459
rect 13474 32425 13508 32459
rect 13542 32425 13576 32459
rect 13610 32425 13644 32459
rect 13678 32425 13712 32459
rect 13746 32425 13780 32459
rect 13814 32425 13848 32459
rect 13882 32425 13916 32459
rect 13950 32425 13984 32459
rect 14018 32425 14052 32459
rect 14086 32425 14120 32459
rect 14154 32425 14188 32459
rect 14222 32425 14256 32459
rect 14290 32425 14324 32459
rect 14358 32425 14392 32459
rect 13202 32356 13236 32390
rect 13270 32356 13304 32390
rect 13338 32356 13372 32390
rect 13406 32356 13440 32390
rect 13474 32356 13508 32390
rect 13542 32356 13576 32390
rect 13610 32356 13644 32390
rect 13678 32356 13712 32390
rect 13746 32356 13780 32390
rect 13814 32356 13848 32390
rect 13882 32356 13916 32390
rect 13950 32356 13984 32390
rect 14018 32356 14052 32390
rect 14086 32356 14120 32390
rect 14154 32356 14188 32390
rect 14222 32356 14256 32390
rect 14290 32356 14324 32390
rect 14358 32356 14392 32390
rect 13202 32287 13236 32321
rect 13270 32287 13304 32321
rect 13338 32287 13372 32321
rect 13406 32287 13440 32321
rect 13474 32287 13508 32321
rect 13542 32287 13576 32321
rect 13610 32287 13644 32321
rect 13678 32287 13712 32321
rect 13746 32287 13780 32321
rect 13814 32287 13848 32321
rect 13882 32287 13916 32321
rect 13950 32287 13984 32321
rect 14018 32287 14052 32321
rect 14086 32287 14120 32321
rect 14154 32287 14188 32321
rect 14222 32287 14256 32321
rect 14290 32287 14324 32321
rect 14358 32287 14392 32321
rect 13202 32218 13236 32252
rect 13270 32218 13304 32252
rect 13338 32218 13372 32252
rect 13406 32218 13440 32252
rect 13474 32218 13508 32252
rect 13542 32218 13576 32252
rect 13610 32218 13644 32252
rect 13678 32218 13712 32252
rect 13746 32218 13780 32252
rect 13814 32218 13848 32252
rect 13882 32218 13916 32252
rect 13950 32218 13984 32252
rect 14018 32218 14052 32252
rect 14086 32218 14120 32252
rect 14154 32218 14188 32252
rect 14222 32218 14256 32252
rect 14290 32218 14324 32252
rect 14358 32218 14392 32252
rect 13202 32149 13236 32183
rect 13270 32149 13304 32183
rect 13338 32149 13372 32183
rect 13406 32149 13440 32183
rect 13474 32149 13508 32183
rect 13542 32149 13576 32183
rect 13610 32149 13644 32183
rect 13678 32149 13712 32183
rect 13746 32149 13780 32183
rect 13814 32149 13848 32183
rect 13882 32149 13916 32183
rect 13950 32149 13984 32183
rect 14018 32149 14052 32183
rect 14086 32149 14120 32183
rect 14154 32149 14188 32183
rect 14222 32149 14256 32183
rect 14290 32149 14324 32183
rect 14358 32149 14392 32183
rect 13202 32080 13236 32114
rect 13270 32080 13304 32114
rect 13338 32080 13372 32114
rect 13406 32080 13440 32114
rect 13474 32080 13508 32114
rect 13542 32080 13576 32114
rect 13610 32080 13644 32114
rect 13678 32080 13712 32114
rect 13746 32080 13780 32114
rect 13814 32080 13848 32114
rect 13882 32080 13916 32114
rect 13950 32080 13984 32114
rect 14018 32080 14052 32114
rect 14086 32080 14120 32114
rect 14154 32080 14188 32114
rect 14222 32080 14256 32114
rect 14290 32080 14324 32114
rect 14358 32080 14392 32114
rect 13202 32011 13236 32045
rect 13270 32011 13304 32045
rect 13338 32011 13372 32045
rect 13406 32011 13440 32045
rect 13474 32011 13508 32045
rect 13542 32011 13576 32045
rect 13610 32011 13644 32045
rect 13678 32011 13712 32045
rect 13746 32011 13780 32045
rect 13814 32011 13848 32045
rect 13882 32011 13916 32045
rect 13950 32011 13984 32045
rect 14018 32011 14052 32045
rect 14086 32011 14120 32045
rect 14154 32011 14188 32045
rect 14222 32011 14256 32045
rect 14290 32011 14324 32045
rect 14358 32011 14392 32045
rect 13202 31942 13236 31976
rect 13270 31942 13304 31976
rect 13338 31942 13372 31976
rect 13406 31942 13440 31976
rect 13474 31942 13508 31976
rect 13542 31942 13576 31976
rect 13610 31942 13644 31976
rect 13678 31942 13712 31976
rect 13746 31942 13780 31976
rect 13814 31942 13848 31976
rect 13882 31942 13916 31976
rect 13950 31942 13984 31976
rect 14018 31942 14052 31976
rect 14086 31942 14120 31976
rect 14154 31942 14188 31976
rect 14222 31942 14256 31976
rect 14290 31942 14324 31976
rect 14358 31942 14392 31976
rect 13202 31873 13236 31907
rect 13270 31873 13304 31907
rect 13338 31873 13372 31907
rect 13406 31873 13440 31907
rect 13474 31873 13508 31907
rect 13542 31873 13576 31907
rect 13610 31873 13644 31907
rect 13678 31873 13712 31907
rect 13746 31873 13780 31907
rect 13814 31873 13848 31907
rect 13882 31873 13916 31907
rect 13950 31873 13984 31907
rect 14018 31873 14052 31907
rect 14086 31873 14120 31907
rect 14154 31873 14188 31907
rect 14222 31873 14256 31907
rect 14290 31873 14324 31907
rect 14358 31873 14392 31907
rect 13202 31804 13236 31838
rect 13270 31804 13304 31838
rect 13338 31804 13372 31838
rect 13406 31804 13440 31838
rect 13474 31804 13508 31838
rect 13542 31804 13576 31838
rect 13610 31804 13644 31838
rect 13678 31804 13712 31838
rect 13746 31804 13780 31838
rect 13814 31804 13848 31838
rect 13882 31804 13916 31838
rect 13950 31804 13984 31838
rect 14018 31804 14052 31838
rect 14086 31804 14120 31838
rect 14154 31804 14188 31838
rect 14222 31804 14256 31838
rect 14290 31804 14324 31838
rect 14358 31804 14392 31838
rect 13202 31735 13236 31769
rect 13270 31735 13304 31769
rect 13338 31735 13372 31769
rect 13406 31735 13440 31769
rect 13474 31735 13508 31769
rect 13542 31735 13576 31769
rect 13610 31735 13644 31769
rect 13678 31735 13712 31769
rect 13746 31735 13780 31769
rect 13814 31735 13848 31769
rect 13882 31735 13916 31769
rect 13950 31735 13984 31769
rect 14018 31735 14052 31769
rect 14086 31735 14120 31769
rect 14154 31735 14188 31769
rect 14222 31735 14256 31769
rect 14290 31735 14324 31769
rect 14358 31735 14392 31769
rect 13202 31666 13236 31700
rect 13270 31666 13304 31700
rect 13338 31666 13372 31700
rect 13406 31666 13440 31700
rect 13474 31666 13508 31700
rect 13542 31666 13576 31700
rect 13610 31666 13644 31700
rect 13678 31666 13712 31700
rect 13746 31666 13780 31700
rect 13814 31666 13848 31700
rect 13882 31666 13916 31700
rect 13950 31666 13984 31700
rect 14018 31666 14052 31700
rect 14086 31666 14120 31700
rect 14154 31666 14188 31700
rect 14222 31666 14256 31700
rect 14290 31666 14324 31700
rect 14358 31666 14392 31700
rect 13202 31597 13236 31631
rect 13270 31597 13304 31631
rect 13338 31597 13372 31631
rect 13406 31597 13440 31631
rect 13474 31597 13508 31631
rect 13542 31597 13576 31631
rect 13610 31597 13644 31631
rect 13678 31597 13712 31631
rect 13746 31597 13780 31631
rect 13814 31597 13848 31631
rect 13882 31597 13916 31631
rect 13950 31597 13984 31631
rect 14018 31597 14052 31631
rect 14086 31597 14120 31631
rect 14154 31597 14188 31631
rect 14222 31597 14256 31631
rect 14290 31597 14324 31631
rect 14358 31597 14392 31631
rect 13202 31528 13236 31562
rect 13270 31528 13304 31562
rect 13338 31528 13372 31562
rect 13406 31528 13440 31562
rect 13474 31528 13508 31562
rect 13542 31528 13576 31562
rect 13610 31528 13644 31562
rect 13678 31528 13712 31562
rect 13746 31528 13780 31562
rect 13814 31528 13848 31562
rect 13882 31528 13916 31562
rect 13950 31528 13984 31562
rect 14018 31528 14052 31562
rect 14086 31528 14120 31562
rect 14154 31528 14188 31562
rect 14222 31528 14256 31562
rect 14290 31528 14324 31562
rect 14358 31528 14392 31562
rect 13202 31459 13236 31493
rect 13270 31459 13304 31493
rect 13338 31459 13372 31493
rect 13406 31459 13440 31493
rect 13474 31459 13508 31493
rect 13542 31459 13576 31493
rect 13610 31459 13644 31493
rect 13678 31459 13712 31493
rect 13746 31459 13780 31493
rect 13814 31459 13848 31493
rect 13882 31459 13916 31493
rect 13950 31459 13984 31493
rect 14018 31459 14052 31493
rect 14086 31459 14120 31493
rect 14154 31459 14188 31493
rect 14222 31459 14256 31493
rect 14290 31459 14324 31493
rect 14358 31459 14392 31493
rect 13202 31390 13236 31424
rect 13270 31390 13304 31424
rect 13338 31390 13372 31424
rect 13406 31390 13440 31424
rect 13474 31390 13508 31424
rect 13542 31390 13576 31424
rect 13610 31390 13644 31424
rect 13678 31390 13712 31424
rect 13746 31390 13780 31424
rect 13814 31390 13848 31424
rect 13882 31390 13916 31424
rect 13950 31390 13984 31424
rect 14018 31390 14052 31424
rect 14086 31390 14120 31424
rect 14154 31390 14188 31424
rect 14222 31390 14256 31424
rect 14290 31390 14324 31424
rect 14358 31390 14392 31424
rect 13202 31321 13236 31355
rect 13270 31321 13304 31355
rect 13338 31321 13372 31355
rect 13406 31321 13440 31355
rect 13474 31321 13508 31355
rect 13542 31321 13576 31355
rect 13610 31321 13644 31355
rect 13678 31321 13712 31355
rect 13746 31321 13780 31355
rect 13814 31321 13848 31355
rect 13882 31321 13916 31355
rect 13950 31321 13984 31355
rect 14018 31321 14052 31355
rect 14086 31321 14120 31355
rect 14154 31321 14188 31355
rect 14222 31321 14256 31355
rect 14290 31321 14324 31355
rect 14358 31321 14392 31355
rect 13202 31252 13236 31286
rect 13270 31252 13304 31286
rect 13338 31252 13372 31286
rect 13406 31252 13440 31286
rect 13474 31252 13508 31286
rect 13542 31252 13576 31286
rect 13610 31252 13644 31286
rect 13678 31252 13712 31286
rect 13746 31252 13780 31286
rect 13814 31252 13848 31286
rect 13882 31252 13916 31286
rect 13950 31252 13984 31286
rect 14018 31252 14052 31286
rect 14086 31252 14120 31286
rect 14154 31252 14188 31286
rect 14222 31252 14256 31286
rect 14290 31252 14324 31286
rect 14358 31252 14392 31286
rect 13202 31183 13236 31217
rect 13270 31183 13304 31217
rect 13338 31183 13372 31217
rect 13406 31183 13440 31217
rect 13474 31183 13508 31217
rect 13542 31183 13576 31217
rect 13610 31183 13644 31217
rect 13678 31183 13712 31217
rect 13746 31183 13780 31217
rect 13814 31183 13848 31217
rect 13882 31183 13916 31217
rect 13950 31183 13984 31217
rect 14018 31183 14052 31217
rect 14086 31183 14120 31217
rect 14154 31183 14188 31217
rect 14222 31183 14256 31217
rect 14290 31183 14324 31217
rect 14358 31183 14392 31217
rect 9913 30602 9947 30636
rect 9982 30602 10016 30636
rect 10051 30602 10085 30636
rect 10120 30602 10154 30636
rect 10189 30602 10223 30636
rect 10258 30602 10292 30636
rect 10327 30602 10361 30636
rect 10396 30602 10430 30636
rect 10465 30602 10499 30636
rect 10610 30601 10644 30635
rect 10679 30601 10713 30635
rect 10747 30601 10781 30635
rect 10815 30601 10849 30635
rect 10883 30601 10917 30635
rect 10951 30601 10985 30635
rect 11019 30601 11053 30635
rect 11087 30601 11121 30635
rect 11155 30601 11189 30635
rect 11223 30601 11257 30635
rect 11291 30601 11325 30635
rect 11359 30601 11393 30635
rect 11427 30601 11461 30635
rect 11495 30601 11529 30635
rect 11563 30601 11597 30635
rect 11631 30601 11665 30635
rect 11699 30601 11733 30635
rect 11767 30601 11801 30635
rect 11835 30601 11869 30635
rect 11903 30601 11937 30635
rect 11971 30601 12005 30635
rect 12039 30601 12073 30635
rect 12107 30601 12141 30635
rect 12175 30601 12209 30635
rect 12243 30601 12277 30635
rect 12311 30601 12345 30635
rect 12379 30601 12413 30635
rect 12447 30601 12481 30635
rect 12515 30601 12549 30635
rect 12583 30601 12617 30635
rect 12651 30601 12685 30635
rect 12719 30601 12753 30635
rect 12787 30601 12821 30635
rect 12855 30601 12889 30635
rect 12923 30601 12957 30635
rect 12991 30601 13025 30635
rect 13059 30601 13093 30635
rect 13127 30601 13161 30635
rect 13195 30601 13229 30635
rect 13263 30601 13297 30635
rect 13331 30601 13365 30635
rect 13399 30601 13433 30635
rect 13467 30601 13501 30635
rect 13535 30601 13569 30635
rect 13603 30601 13637 30635
rect 13671 30601 13705 30635
rect 13739 30601 13773 30635
rect 13807 30601 13841 30635
rect 13875 30601 13909 30635
rect 9913 30534 9947 30568
rect 9982 30534 10016 30568
rect 10051 30534 10085 30568
rect 10120 30534 10154 30568
rect 10189 30534 10223 30568
rect 10258 30534 10292 30568
rect 10327 30534 10361 30568
rect 10396 30534 10430 30568
rect 10465 30534 10499 30568
rect 10610 30526 10644 30560
rect 10679 30526 10713 30560
rect 10747 30526 10781 30560
rect 10815 30526 10849 30560
rect 10883 30526 10917 30560
rect 10951 30526 10985 30560
rect 11019 30526 11053 30560
rect 11087 30526 11121 30560
rect 11155 30526 11189 30560
rect 11223 30526 11257 30560
rect 11291 30526 11325 30560
rect 11359 30526 11393 30560
rect 11427 30526 11461 30560
rect 11495 30526 11529 30560
rect 11563 30526 11597 30560
rect 11631 30526 11665 30560
rect 11699 30526 11733 30560
rect 11767 30526 11801 30560
rect 11835 30526 11869 30560
rect 11903 30526 11937 30560
rect 11971 30526 12005 30560
rect 12039 30526 12073 30560
rect 12107 30526 12141 30560
rect 12175 30526 12209 30560
rect 12243 30526 12277 30560
rect 12311 30526 12345 30560
rect 12379 30526 12413 30560
rect 12447 30526 12481 30560
rect 12515 30526 12549 30560
rect 12583 30526 12617 30560
rect 12651 30526 12685 30560
rect 12719 30526 12753 30560
rect 12787 30526 12821 30560
rect 12855 30526 12889 30560
rect 12923 30526 12957 30560
rect 12991 30526 13025 30560
rect 13059 30526 13093 30560
rect 13127 30526 13161 30560
rect 13195 30526 13229 30560
rect 13263 30526 13297 30560
rect 13331 30526 13365 30560
rect 13399 30526 13433 30560
rect 13467 30526 13501 30560
rect 13535 30526 13569 30560
rect 13603 30526 13637 30560
rect 13671 30526 13705 30560
rect 13739 30526 13773 30560
rect 13807 30526 13841 30560
rect 13875 30526 13909 30560
rect 9913 30466 9947 30500
rect 9982 30466 10016 30500
rect 10051 30466 10085 30500
rect 10120 30466 10154 30500
rect 10189 30466 10223 30500
rect 10258 30466 10292 30500
rect 10327 30466 10361 30500
rect 10396 30466 10430 30500
rect 10465 30466 10499 30500
rect 10610 30451 10644 30485
rect 10679 30451 10713 30485
rect 10747 30451 10781 30485
rect 10815 30451 10849 30485
rect 10883 30451 10917 30485
rect 10951 30451 10985 30485
rect 11019 30451 11053 30485
rect 11087 30451 11121 30485
rect 11155 30451 11189 30485
rect 11223 30451 11257 30485
rect 11291 30451 11325 30485
rect 11359 30451 11393 30485
rect 11427 30451 11461 30485
rect 11495 30451 11529 30485
rect 11563 30451 11597 30485
rect 11631 30451 11665 30485
rect 11699 30451 11733 30485
rect 11767 30451 11801 30485
rect 11835 30451 11869 30485
rect 11903 30451 11937 30485
rect 11971 30451 12005 30485
rect 12039 30451 12073 30485
rect 12107 30451 12141 30485
rect 12175 30451 12209 30485
rect 12243 30451 12277 30485
rect 12311 30451 12345 30485
rect 12379 30451 12413 30485
rect 12447 30451 12481 30485
rect 12515 30451 12549 30485
rect 12583 30451 12617 30485
rect 12651 30451 12685 30485
rect 12719 30451 12753 30485
rect 12787 30451 12821 30485
rect 12855 30451 12889 30485
rect 12923 30451 12957 30485
rect 12991 30451 13025 30485
rect 13059 30451 13093 30485
rect 13127 30451 13161 30485
rect 13195 30451 13229 30485
rect 13263 30451 13297 30485
rect 13331 30451 13365 30485
rect 13399 30451 13433 30485
rect 13467 30451 13501 30485
rect 13535 30451 13569 30485
rect 13603 30451 13637 30485
rect 13671 30451 13705 30485
rect 13739 30451 13773 30485
rect 13807 30451 13841 30485
rect 13875 30451 13909 30485
rect 9913 30398 9947 30432
rect 9982 30398 10016 30432
rect 10051 30398 10085 30432
rect 10120 30398 10154 30432
rect 10189 30398 10223 30432
rect 10258 30398 10292 30432
rect 10327 30398 10361 30432
rect 10396 30398 10430 30432
rect 10465 30398 10499 30432
rect 9913 30330 9947 30364
rect 9982 30330 10016 30364
rect 10051 30330 10085 30364
rect 10120 30330 10154 30364
rect 10189 30330 10223 30364
rect 10258 30330 10292 30364
rect 10327 30330 10361 30364
rect 10396 30330 10430 30364
rect 10465 30330 10499 30364
rect 9913 30262 9947 30296
rect 9982 30262 10016 30296
rect 10051 30262 10085 30296
rect 10120 30262 10154 30296
rect 10189 30262 10223 30296
rect 10258 30262 10292 30296
rect 10327 30262 10361 30296
rect 10396 30262 10430 30296
rect 10465 30262 10499 30296
rect 9913 30194 9947 30228
rect 9982 30194 10016 30228
rect 10051 30194 10085 30228
rect 10120 30194 10154 30228
rect 10189 30194 10223 30228
rect 10258 30194 10292 30228
rect 10327 30194 10361 30228
rect 10396 30194 10430 30228
rect 10465 30194 10499 30228
rect 9913 30126 9947 30160
rect 9982 30126 10016 30160
rect 10051 30126 10085 30160
rect 10120 30126 10154 30160
rect 10189 30126 10223 30160
rect 10258 30126 10292 30160
rect 10327 30126 10361 30160
rect 10396 30126 10430 30160
rect 10465 30126 10499 30160
rect 9913 30058 9947 30092
rect 9982 30058 10016 30092
rect 10051 30058 10085 30092
rect 10120 30058 10154 30092
rect 10189 30058 10223 30092
rect 10258 30058 10292 30092
rect 10327 30058 10361 30092
rect 10396 30058 10430 30092
rect 10465 30058 10499 30092
rect 9913 29990 9947 30024
rect 9982 29990 10016 30024
rect 10051 29990 10085 30024
rect 10120 29990 10154 30024
rect 10189 29990 10223 30024
rect 10258 29990 10292 30024
rect 10327 29990 10361 30024
rect 10396 29990 10430 30024
rect 10465 29990 10499 30024
rect 9913 29922 9947 29956
rect 9982 29922 10016 29956
rect 10051 29922 10085 29956
rect 10120 29922 10154 29956
rect 10189 29922 10223 29956
rect 10258 29922 10292 29956
rect 10327 29922 10361 29956
rect 10396 29922 10430 29956
rect 10465 29922 10499 29956
rect 9913 29854 9947 29888
rect 9982 29854 10016 29888
rect 10051 29854 10085 29888
rect 10120 29854 10154 29888
rect 10189 29854 10223 29888
rect 10258 29854 10292 29888
rect 10327 29854 10361 29888
rect 10396 29854 10430 29888
rect 10465 29854 10499 29888
rect 9913 29786 9947 29820
rect 9982 29786 10016 29820
rect 10051 29786 10085 29820
rect 10120 29786 10154 29820
rect 10189 29786 10223 29820
rect 10258 29786 10292 29820
rect 10327 29786 10361 29820
rect 10396 29786 10430 29820
rect 10465 29786 10499 29820
rect 9913 29718 9947 29752
rect 9982 29718 10016 29752
rect 10051 29718 10085 29752
rect 10120 29718 10154 29752
rect 10189 29718 10223 29752
rect 10258 29718 10292 29752
rect 10327 29718 10361 29752
rect 10396 29718 10430 29752
rect 10465 29718 10499 29752
rect 9913 29650 9947 29684
rect 9982 29650 10016 29684
rect 10051 29650 10085 29684
rect 10120 29650 10154 29684
rect 10189 29650 10223 29684
rect 10258 29650 10292 29684
rect 10327 29650 10361 29684
rect 10396 29650 10430 29684
rect 10465 29650 10499 29684
rect 9913 29582 9947 29616
rect 9982 29582 10016 29616
rect 10051 29582 10085 29616
rect 10120 29582 10154 29616
rect 10189 29582 10223 29616
rect 10258 29582 10292 29616
rect 10327 29582 10361 29616
rect 10396 29582 10430 29616
rect 10465 29582 10499 29616
rect 9913 29514 9947 29548
rect 9982 29514 10016 29548
rect 10051 29514 10085 29548
rect 10120 29514 10154 29548
rect 10189 29514 10223 29548
rect 10258 29514 10292 29548
rect 10327 29514 10361 29548
rect 10396 29514 10430 29548
rect 10465 29514 10499 29548
rect 9913 29446 9947 29480
rect 9982 29446 10016 29480
rect 10051 29446 10085 29480
rect 10120 29446 10154 29480
rect 10189 29446 10223 29480
rect 10258 29446 10292 29480
rect 10327 29446 10361 29480
rect 10396 29446 10430 29480
rect 10465 29446 10499 29480
rect 9913 29378 9947 29412
rect 9982 29378 10016 29412
rect 10051 29378 10085 29412
rect 10120 29378 10154 29412
rect 10189 29378 10223 29412
rect 10258 29378 10292 29412
rect 10327 29378 10361 29412
rect 10396 29378 10430 29412
rect 10465 29378 10499 29412
rect 9913 29310 9947 29344
rect 9982 29310 10016 29344
rect 10051 29310 10085 29344
rect 10120 29310 10154 29344
rect 10189 29310 10223 29344
rect 10258 29310 10292 29344
rect 10327 29310 10361 29344
rect 10396 29310 10430 29344
rect 10465 29310 10499 29344
rect 9913 29242 9947 29276
rect 9982 29242 10016 29276
rect 10051 29242 10085 29276
rect 10120 29242 10154 29276
rect 10189 29242 10223 29276
rect 10258 29242 10292 29276
rect 10327 29242 10361 29276
rect 10396 29242 10430 29276
rect 10465 29242 10499 29276
rect 9913 29174 9947 29208
rect 9982 29174 10016 29208
rect 10051 29174 10085 29208
rect 10120 29174 10154 29208
rect 10189 29174 10223 29208
rect 10258 29174 10292 29208
rect 10327 29174 10361 29208
rect 10396 29174 10430 29208
rect 10465 29174 10499 29208
rect 9913 29106 9947 29140
rect 9982 29106 10016 29140
rect 10051 29106 10085 29140
rect 10120 29106 10154 29140
rect 10189 29106 10223 29140
rect 10258 29106 10292 29140
rect 10327 29106 10361 29140
rect 10396 29106 10430 29140
rect 10465 29106 10499 29140
rect 9913 29038 9947 29072
rect 9982 29038 10016 29072
rect 10051 29038 10085 29072
rect 10120 29038 10154 29072
rect 10189 29038 10223 29072
rect 10258 29038 10292 29072
rect 10327 29038 10361 29072
rect 10396 29038 10430 29072
rect 10465 29038 10499 29072
rect 9913 28970 9947 29004
rect 9982 28970 10016 29004
rect 10051 28970 10085 29004
rect 10120 28970 10154 29004
rect 10189 28970 10223 29004
rect 10258 28970 10292 29004
rect 10327 28970 10361 29004
rect 10396 28970 10430 29004
rect 10465 28970 10499 29004
rect 9913 28902 9947 28936
rect 9982 28902 10016 28936
rect 10051 28902 10085 28936
rect 10120 28902 10154 28936
rect 10189 28902 10223 28936
rect 10258 28902 10292 28936
rect 10327 28902 10361 28936
rect 10396 28902 10430 28936
rect 10465 28902 10499 28936
rect 9913 28834 9947 28868
rect 9982 28834 10016 28868
rect 10051 28834 10085 28868
rect 10120 28834 10154 28868
rect 10189 28834 10223 28868
rect 10258 28834 10292 28868
rect 10327 28834 10361 28868
rect 10396 28834 10430 28868
rect 10465 28834 10499 28868
rect 9913 28766 9947 28800
rect 9982 28766 10016 28800
rect 10051 28766 10085 28800
rect 10120 28766 10154 28800
rect 10189 28766 10223 28800
rect 10258 28766 10292 28800
rect 10327 28766 10361 28800
rect 10396 28766 10430 28800
rect 10465 28766 10499 28800
rect 9913 28698 9947 28732
rect 9982 28698 10016 28732
rect 10051 28698 10085 28732
rect 10120 28698 10154 28732
rect 10189 28698 10223 28732
rect 10258 28698 10292 28732
rect 10327 28698 10361 28732
rect 10396 28698 10430 28732
rect 10465 28698 10499 28732
rect 9913 28630 9947 28664
rect 9982 28630 10016 28664
rect 10051 28630 10085 28664
rect 10120 28630 10154 28664
rect 10189 28630 10223 28664
rect 10258 28630 10292 28664
rect 10327 28630 10361 28664
rect 10396 28630 10430 28664
rect 10465 28630 10499 28664
rect 9913 28562 9947 28596
rect 9982 28562 10016 28596
rect 10051 28562 10085 28596
rect 10120 28562 10154 28596
rect 10189 28562 10223 28596
rect 10258 28562 10292 28596
rect 10327 28562 10361 28596
rect 10396 28562 10430 28596
rect 10465 28562 10499 28596
rect 9913 28494 9947 28528
rect 9982 28494 10016 28528
rect 10051 28494 10085 28528
rect 10120 28494 10154 28528
rect 10189 28494 10223 28528
rect 10258 28494 10292 28528
rect 10327 28494 10361 28528
rect 10396 28494 10430 28528
rect 10465 28494 10499 28528
rect 9913 28426 9947 28460
rect 9982 28426 10016 28460
rect 10051 28426 10085 28460
rect 10120 28426 10154 28460
rect 10189 28426 10223 28460
rect 10258 28426 10292 28460
rect 10327 28426 10361 28460
rect 10396 28426 10430 28460
rect 10465 28426 10499 28460
rect 9913 28358 9947 28392
rect 9982 28358 10016 28392
rect 10051 28358 10085 28392
rect 10120 28358 10154 28392
rect 10189 28358 10223 28392
rect 10258 28358 10292 28392
rect 10327 28358 10361 28392
rect 10396 28358 10430 28392
rect 10465 28358 10499 28392
rect 9913 28290 9947 28324
rect 9982 28290 10016 28324
rect 10051 28290 10085 28324
rect 10120 28290 10154 28324
rect 10189 28290 10223 28324
rect 10258 28290 10292 28324
rect 10327 28290 10361 28324
rect 10396 28290 10430 28324
rect 10465 28290 10499 28324
rect 9913 28222 9947 28256
rect 9982 28222 10016 28256
rect 10051 28222 10085 28256
rect 10120 28222 10154 28256
rect 10189 28222 10223 28256
rect 10258 28222 10292 28256
rect 10327 28222 10361 28256
rect 10396 28222 10430 28256
rect 10465 28222 10499 28256
rect 9913 28154 9947 28188
rect 9982 28154 10016 28188
rect 10051 28154 10085 28188
rect 10120 28154 10154 28188
rect 10189 28154 10223 28188
rect 10258 28154 10292 28188
rect 10327 28154 10361 28188
rect 10396 28154 10430 28188
rect 10465 28154 10499 28188
rect 9913 28086 9947 28120
rect 9982 28086 10016 28120
rect 10051 28086 10085 28120
rect 10120 28086 10154 28120
rect 10189 28086 10223 28120
rect 10258 28086 10292 28120
rect 10327 28086 10361 28120
rect 10396 28086 10430 28120
rect 10465 28086 10499 28120
rect 9913 28018 9947 28052
rect 9982 28018 10016 28052
rect 10051 28018 10085 28052
rect 10120 28018 10154 28052
rect 10189 28018 10223 28052
rect 10258 28018 10292 28052
rect 10327 28018 10361 28052
rect 10396 28018 10430 28052
rect 10465 28018 10499 28052
rect 9913 27949 9947 27983
rect 9982 27949 10016 27983
rect 10051 27949 10085 27983
rect 10120 27949 10154 27983
rect 10189 27949 10223 27983
rect 10258 27949 10292 27983
rect 10327 27949 10361 27983
rect 10396 27949 10430 27983
rect 10465 27949 10499 27983
rect 9913 27880 9947 27914
rect 9982 27880 10016 27914
rect 10051 27880 10085 27914
rect 10120 27880 10154 27914
rect 10189 27880 10223 27914
rect 10258 27880 10292 27914
rect 10327 27880 10361 27914
rect 10396 27880 10430 27914
rect 10465 27880 10499 27914
rect 9913 27811 9947 27845
rect 9982 27811 10016 27845
rect 10051 27811 10085 27845
rect 10120 27811 10154 27845
rect 10189 27811 10223 27845
rect 10258 27811 10292 27845
rect 10327 27811 10361 27845
rect 10396 27811 10430 27845
rect 10465 27811 10499 27845
rect 9913 27742 9947 27776
rect 9982 27742 10016 27776
rect 10051 27742 10085 27776
rect 10120 27742 10154 27776
rect 10189 27742 10223 27776
rect 10258 27742 10292 27776
rect 10327 27742 10361 27776
rect 10396 27742 10430 27776
rect 10465 27742 10499 27776
rect 9913 27673 9947 27707
rect 9982 27673 10016 27707
rect 10051 27673 10085 27707
rect 10120 27673 10154 27707
rect 10189 27673 10223 27707
rect 10258 27673 10292 27707
rect 10327 27673 10361 27707
rect 10396 27673 10430 27707
rect 10465 27673 10499 27707
rect 9913 27604 9947 27638
rect 9982 27604 10016 27638
rect 10051 27604 10085 27638
rect 10120 27604 10154 27638
rect 10189 27604 10223 27638
rect 10258 27604 10292 27638
rect 10327 27604 10361 27638
rect 10396 27604 10430 27638
rect 10465 27604 10499 27638
rect 9913 27535 9947 27569
rect 9982 27535 10016 27569
rect 10051 27535 10085 27569
rect 10120 27535 10154 27569
rect 10189 27535 10223 27569
rect 10258 27535 10292 27569
rect 10327 27535 10361 27569
rect 10396 27535 10430 27569
rect 10465 27535 10499 27569
rect 9913 27466 9947 27500
rect 9982 27466 10016 27500
rect 10051 27466 10085 27500
rect 10120 27466 10154 27500
rect 10189 27466 10223 27500
rect 10258 27466 10292 27500
rect 10327 27466 10361 27500
rect 10396 27466 10430 27500
rect 10465 27466 10499 27500
rect 9913 27397 9947 27431
rect 9982 27397 10016 27431
rect 10051 27397 10085 27431
rect 10120 27397 10154 27431
rect 10189 27397 10223 27431
rect 10258 27397 10292 27431
rect 10327 27397 10361 27431
rect 10396 27397 10430 27431
rect 10465 27397 10499 27431
rect 9913 27328 9947 27362
rect 9982 27328 10016 27362
rect 10051 27328 10085 27362
rect 10120 27328 10154 27362
rect 10189 27328 10223 27362
rect 10258 27328 10292 27362
rect 10327 27328 10361 27362
rect 10396 27328 10430 27362
rect 10465 27328 10499 27362
rect 9913 27259 9947 27293
rect 9982 27259 10016 27293
rect 10051 27259 10085 27293
rect 10120 27259 10154 27293
rect 10189 27259 10223 27293
rect 10258 27259 10292 27293
rect 10327 27259 10361 27293
rect 10396 27259 10430 27293
rect 10465 27259 10499 27293
rect 9913 27190 9947 27224
rect 9982 27190 10016 27224
rect 10051 27190 10085 27224
rect 10120 27190 10154 27224
rect 10189 27190 10223 27224
rect 10258 27190 10292 27224
rect 10327 27190 10361 27224
rect 10396 27190 10430 27224
rect 10465 27190 10499 27224
rect 9913 27121 9947 27155
rect 9982 27121 10016 27155
rect 10051 27121 10085 27155
rect 10120 27121 10154 27155
rect 10189 27121 10223 27155
rect 10258 27121 10292 27155
rect 10327 27121 10361 27155
rect 10396 27121 10430 27155
rect 10465 27121 10499 27155
rect 9913 27052 9947 27086
rect 9982 27052 10016 27086
rect 10051 27052 10085 27086
rect 10120 27052 10154 27086
rect 10189 27052 10223 27086
rect 10258 27052 10292 27086
rect 10327 27052 10361 27086
rect 10396 27052 10430 27086
rect 10465 27052 10499 27086
rect 13738 29007 13908 30401
rect 13738 28938 13772 28972
rect 13806 28938 13840 28972
rect 13874 28938 13908 28972
rect 13738 28869 13772 28903
rect 13806 28869 13840 28903
rect 13874 28869 13908 28903
rect 13738 28800 13772 28834
rect 13806 28800 13840 28834
rect 13874 28800 13908 28834
rect 13738 28731 13772 28765
rect 13806 28731 13840 28765
rect 13874 28731 13908 28765
rect 13738 28662 13772 28696
rect 13806 28662 13840 28696
rect 13874 28662 13908 28696
rect 13738 28593 13772 28627
rect 13806 28593 13840 28627
rect 13874 28593 13908 28627
rect 13738 28524 13772 28558
rect 13806 28524 13840 28558
rect 13874 28524 13908 28558
rect 13738 28455 13772 28489
rect 13806 28455 13840 28489
rect 13874 28455 13908 28489
rect 13738 28386 13772 28420
rect 13806 28386 13840 28420
rect 13874 28386 13908 28420
rect 13738 28317 13772 28351
rect 13806 28317 13840 28351
rect 13874 28317 13908 28351
rect 13738 28248 13772 28282
rect 13806 28248 13840 28282
rect 13874 28248 13908 28282
rect 13738 28179 13772 28213
rect 13806 28179 13840 28213
rect 13874 28179 13908 28213
rect 13738 28110 13772 28144
rect 13806 28110 13840 28144
rect 13874 28110 13908 28144
rect 13738 28041 13772 28075
rect 13806 28041 13840 28075
rect 13874 28041 13908 28075
rect 13738 27972 13772 28006
rect 13806 27972 13840 28006
rect 13874 27972 13908 28006
rect 13738 27903 13772 27937
rect 13806 27903 13840 27937
rect 13874 27903 13908 27937
rect 13738 27834 13772 27868
rect 13806 27834 13840 27868
rect 13874 27834 13908 27868
rect 13738 27765 13772 27799
rect 13806 27765 13840 27799
rect 13874 27765 13908 27799
rect 13738 27696 13772 27730
rect 13806 27696 13840 27730
rect 13874 27696 13908 27730
rect 13738 27627 13772 27661
rect 13806 27627 13840 27661
rect 13874 27627 13908 27661
rect 13738 27558 13772 27592
rect 13806 27558 13840 27592
rect 13874 27558 13908 27592
rect 13738 27489 13772 27523
rect 13806 27489 13840 27523
rect 13874 27489 13908 27523
rect 13738 27420 13772 27454
rect 13806 27420 13840 27454
rect 13874 27420 13908 27454
rect 13738 27351 13772 27385
rect 13806 27351 13840 27385
rect 13874 27351 13908 27385
rect 13738 27282 13772 27316
rect 13806 27282 13840 27316
rect 13874 27282 13908 27316
rect 13738 27213 13772 27247
rect 13806 27213 13840 27247
rect 13874 27213 13908 27247
rect 13738 27144 13772 27178
rect 13806 27144 13840 27178
rect 13874 27144 13908 27178
rect 13738 27075 13772 27109
rect 13806 27075 13840 27109
rect 13874 27075 13908 27109
rect 13738 27006 13772 27040
rect 13806 27006 13840 27040
rect 13874 27006 13908 27040
rect 9911 26904 9945 26938
rect 9980 26904 10014 26938
rect 10049 26904 10083 26938
rect 10118 26904 10152 26938
rect 10187 26904 10221 26938
rect 10256 26904 10290 26938
rect 10325 26904 10359 26938
rect 10394 26904 10428 26938
rect 10463 26904 10497 26938
rect 10532 26904 10566 26938
rect 10601 26904 10635 26938
rect 10670 26904 10704 26938
rect 10739 26904 10773 26938
rect 10808 26904 10842 26938
rect 10877 26904 10911 26938
rect 10946 26904 10980 26938
rect 11015 26904 11049 26938
rect 11084 26904 11118 26938
rect 11153 26904 11187 26938
rect 11222 26904 11256 26938
rect 11291 26904 11325 26938
rect 11359 26904 11393 26938
rect 11427 26904 11461 26938
rect 11495 26904 11529 26938
rect 11563 26904 11597 26938
rect 11631 26904 11665 26938
rect 11699 26904 11733 26938
rect 11767 26904 11801 26938
rect 11835 26904 11869 26938
rect 11903 26904 11937 26938
rect 11971 26904 12005 26938
rect 12039 26904 12073 26938
rect 12107 26904 12141 26938
rect 12175 26904 12209 26938
rect 12243 26904 12277 26938
rect 12311 26904 12345 26938
rect 12379 26904 12413 26938
rect 12447 26904 12481 26938
rect 12515 26904 12549 26938
rect 12583 26904 12617 26938
rect 12651 26904 12685 26938
rect 12719 26904 12753 26938
rect 12787 26904 12821 26938
rect 12855 26904 12889 26938
rect 12923 26904 12957 26938
rect 12991 26904 13025 26938
rect 13059 26904 13093 26938
rect 13127 26904 13161 26938
rect 13195 26904 13229 26938
rect 13263 26904 13297 26938
rect 13331 26904 13365 26938
rect 13399 26904 13433 26938
rect 13467 26904 13501 26938
rect 13535 26904 13569 26938
rect 13603 26904 13637 26938
rect 13671 26904 13705 26938
rect 13739 26904 13773 26938
rect 13807 26904 13841 26938
rect 13875 26904 13909 26938
rect 9911 26832 9945 26866
rect 9980 26832 10014 26866
rect 10049 26832 10083 26866
rect 10118 26832 10152 26866
rect 10187 26832 10221 26866
rect 10256 26832 10290 26866
rect 10325 26832 10359 26866
rect 10394 26832 10428 26866
rect 10463 26832 10497 26866
rect 10532 26832 10566 26866
rect 10601 26832 10635 26866
rect 10670 26832 10704 26866
rect 10739 26832 10773 26866
rect 10808 26832 10842 26866
rect 10877 26832 10911 26866
rect 10946 26832 10980 26866
rect 11015 26832 11049 26866
rect 11084 26832 11118 26866
rect 11153 26832 11187 26866
rect 11222 26832 11256 26866
rect 11291 26832 11325 26866
rect 11359 26832 11393 26866
rect 11427 26832 11461 26866
rect 11495 26832 11529 26866
rect 11563 26832 11597 26866
rect 11631 26832 11665 26866
rect 11699 26832 11733 26866
rect 11767 26832 11801 26866
rect 11835 26832 11869 26866
rect 11903 26832 11937 26866
rect 11971 26832 12005 26866
rect 12039 26832 12073 26866
rect 12107 26832 12141 26866
rect 12175 26832 12209 26866
rect 12243 26832 12277 26866
rect 12311 26832 12345 26866
rect 12379 26832 12413 26866
rect 12447 26832 12481 26866
rect 12515 26832 12549 26866
rect 12583 26832 12617 26866
rect 12651 26832 12685 26866
rect 12719 26832 12753 26866
rect 12787 26832 12821 26866
rect 12855 26832 12889 26866
rect 12923 26832 12957 26866
rect 12991 26832 13025 26866
rect 13059 26832 13093 26866
rect 13127 26832 13161 26866
rect 13195 26832 13229 26866
rect 13263 26832 13297 26866
rect 13331 26832 13365 26866
rect 13399 26832 13433 26866
rect 13467 26832 13501 26866
rect 13535 26832 13569 26866
rect 13603 26832 13637 26866
rect 13671 26832 13705 26866
rect 13739 26832 13773 26866
rect 13807 26832 13841 26866
rect 13875 26832 13909 26866
rect 9911 26760 9945 26794
rect 9980 26760 10014 26794
rect 10049 26760 10083 26794
rect 10118 26760 10152 26794
rect 10187 26760 10221 26794
rect 10256 26760 10290 26794
rect 10325 26760 10359 26794
rect 10394 26760 10428 26794
rect 10463 26760 10497 26794
rect 10532 26760 10566 26794
rect 10601 26760 10635 26794
rect 10670 26760 10704 26794
rect 10739 26760 10773 26794
rect 10808 26760 10842 26794
rect 10877 26760 10911 26794
rect 10946 26760 10980 26794
rect 11015 26760 11049 26794
rect 11084 26760 11118 26794
rect 11153 26760 11187 26794
rect 11222 26760 11256 26794
rect 11291 26760 11325 26794
rect 11359 26760 11393 26794
rect 11427 26760 11461 26794
rect 11495 26760 11529 26794
rect 11563 26760 11597 26794
rect 11631 26760 11665 26794
rect 11699 26760 11733 26794
rect 11767 26760 11801 26794
rect 11835 26760 11869 26794
rect 11903 26760 11937 26794
rect 11971 26760 12005 26794
rect 12039 26760 12073 26794
rect 12107 26760 12141 26794
rect 12175 26760 12209 26794
rect 12243 26760 12277 26794
rect 12311 26760 12345 26794
rect 12379 26760 12413 26794
rect 12447 26760 12481 26794
rect 12515 26760 12549 26794
rect 12583 26760 12617 26794
rect 12651 26760 12685 26794
rect 12719 26760 12753 26794
rect 12787 26760 12821 26794
rect 12855 26760 12889 26794
rect 12923 26760 12957 26794
rect 12991 26760 13025 26794
rect 13059 26760 13093 26794
rect 13127 26760 13161 26794
rect 13195 26760 13229 26794
rect 13263 26760 13297 26794
rect 13331 26760 13365 26794
rect 13399 26760 13433 26794
rect 13467 26760 13501 26794
rect 13535 26760 13569 26794
rect 13603 26760 13637 26794
rect 13671 26760 13705 26794
rect 13739 26760 13773 26794
rect 13807 26760 13841 26794
rect 13875 26760 13909 26794
rect 9911 26165 9945 26199
rect 9980 26165 10014 26199
rect 10049 26165 10083 26199
rect 10118 26165 10152 26199
rect 10187 26165 10221 26199
rect 10256 26165 10290 26199
rect 10325 26165 10359 26199
rect 10394 26165 10428 26199
rect 10463 26165 10497 26199
rect 10532 26165 10566 26199
rect 10601 26165 10635 26199
rect 10670 26165 10704 26199
rect 10739 26165 10773 26199
rect 10807 26165 10841 26199
rect 10875 26165 10909 26199
rect 10943 26165 10977 26199
rect 11011 26165 11045 26199
rect 11079 26165 11113 26199
rect 11147 26165 11181 26199
rect 11215 26165 11249 26199
rect 11283 26165 11317 26199
rect 11351 26165 11385 26199
rect 11419 26165 11453 26199
rect 11487 26165 11521 26199
rect 11555 26165 11589 26199
rect 11623 26165 11657 26199
rect 11691 26165 11725 26199
rect 11759 26165 11793 26199
rect 11827 26165 11861 26199
rect 11895 26165 11929 26199
rect 11963 26165 11997 26199
rect 12031 26165 12065 26199
rect 12099 26165 12133 26199
rect 12167 26165 12201 26199
rect 12235 26165 12269 26199
rect 12303 26165 12337 26199
rect 12371 26165 12405 26199
rect 12439 26165 12473 26199
rect 12507 26165 12541 26199
rect 12575 26165 12609 26199
rect 12643 26165 12677 26199
rect 12711 26165 12745 26199
rect 12779 26165 12813 26199
rect 12847 26165 12881 26199
rect 12915 26165 12949 26199
rect 12983 26165 13017 26199
rect 13051 26165 13085 26199
rect 13119 26165 13153 26199
rect 13187 26165 13221 26199
rect 13255 26165 13289 26199
rect 13323 26165 13357 26199
rect 13391 26165 13425 26199
rect 13459 26165 13493 26199
rect 13527 26165 13561 26199
rect 13595 26165 13629 26199
rect 13663 26165 13697 26199
rect 13731 26165 13765 26199
rect 13799 26165 13833 26199
rect 13867 26165 13901 26199
rect 13935 26165 13969 26199
rect 14003 26165 14037 26199
rect 14071 26165 14105 26199
rect 14139 26165 14173 26199
rect 9911 26095 9945 26129
rect 9980 26095 10014 26129
rect 10049 26095 10083 26129
rect 10118 26095 10152 26129
rect 10187 26095 10221 26129
rect 10256 26095 10290 26129
rect 10325 26095 10359 26129
rect 10394 26095 10428 26129
rect 10463 26095 10497 26129
rect 10532 26095 10566 26129
rect 10601 26095 10635 26129
rect 10670 26095 10704 26129
rect 10739 26095 10773 26129
rect 10807 26095 10841 26129
rect 10875 26095 10909 26129
rect 10943 26095 10977 26129
rect 11011 26095 11045 26129
rect 11079 26095 11113 26129
rect 11147 26095 11181 26129
rect 11215 26095 11249 26129
rect 11283 26095 11317 26129
rect 11351 26095 11385 26129
rect 11419 26095 11453 26129
rect 11487 26095 11521 26129
rect 11555 26095 11589 26129
rect 11623 26095 11657 26129
rect 11691 26095 11725 26129
rect 11759 26095 11793 26129
rect 11827 26095 11861 26129
rect 11895 26095 11929 26129
rect 11963 26095 11997 26129
rect 12031 26095 12065 26129
rect 12099 26095 12133 26129
rect 12167 26095 12201 26129
rect 12235 26095 12269 26129
rect 12303 26095 12337 26129
rect 12371 26095 12405 26129
rect 12439 26095 12473 26129
rect 12507 26095 12541 26129
rect 12575 26095 12609 26129
rect 12643 26095 12677 26129
rect 12711 26095 12745 26129
rect 12779 26095 12813 26129
rect 12847 26095 12881 26129
rect 12915 26095 12949 26129
rect 12983 26095 13017 26129
rect 13051 26095 13085 26129
rect 13119 26095 13153 26129
rect 13187 26095 13221 26129
rect 13255 26095 13289 26129
rect 13323 26095 13357 26129
rect 13391 26095 13425 26129
rect 13459 26095 13493 26129
rect 13527 26095 13561 26129
rect 13595 26095 13629 26129
rect 13663 26095 13697 26129
rect 13731 26095 13765 26129
rect 13799 26095 13833 26129
rect 13867 26095 13901 26129
rect 13935 26095 13969 26129
rect 14003 26095 14037 26129
rect 14071 26095 14105 26129
rect 14139 26095 14173 26129
rect 9911 26025 9945 26059
rect 9980 26025 10014 26059
rect 10049 26025 10083 26059
rect 10118 26025 10152 26059
rect 10187 26025 10221 26059
rect 10256 26025 10290 26059
rect 10325 26025 10359 26059
rect 10394 26025 10428 26059
rect 10463 26025 10497 26059
rect 10532 26025 10566 26059
rect 10601 26025 10635 26059
rect 10670 26025 10704 26059
rect 10739 26025 10773 26059
rect 10807 26025 10841 26059
rect 10875 26025 10909 26059
rect 10943 26025 10977 26059
rect 11011 26025 11045 26059
rect 11079 26025 11113 26059
rect 11147 26025 11181 26059
rect 11215 26025 11249 26059
rect 11283 26025 11317 26059
rect 11351 26025 11385 26059
rect 11419 26025 11453 26059
rect 11487 26025 11521 26059
rect 11555 26025 11589 26059
rect 11623 26025 11657 26059
rect 11691 26025 11725 26059
rect 11759 26025 11793 26059
rect 11827 26025 11861 26059
rect 11895 26025 11929 26059
rect 11963 26025 11997 26059
rect 12031 26025 12065 26059
rect 12099 26025 12133 26059
rect 12167 26025 12201 26059
rect 12235 26025 12269 26059
rect 12303 26025 12337 26059
rect 12371 26025 12405 26059
rect 12439 26025 12473 26059
rect 12507 26025 12541 26059
rect 12575 26025 12609 26059
rect 12643 26025 12677 26059
rect 12711 26025 12745 26059
rect 12779 26025 12813 26059
rect 12847 26025 12881 26059
rect 12915 26025 12949 26059
rect 12983 26025 13017 26059
rect 13051 26025 13085 26059
rect 13119 26025 13153 26059
rect 13187 26025 13221 26059
rect 13255 26025 13289 26059
rect 13323 26025 13357 26059
rect 13391 26025 13425 26059
rect 13459 26025 13493 26059
rect 13527 26025 13561 26059
rect 13595 26025 13629 26059
rect 13663 26025 13697 26059
rect 13731 26025 13765 26059
rect 13799 26025 13833 26059
rect 13867 26025 13901 26059
rect 13935 26025 13969 26059
rect 14003 26025 14037 26059
rect 14071 26025 14105 26059
rect 14139 26025 14173 26059
rect 9911 25955 9945 25989
rect 9980 25955 10014 25989
rect 10049 25955 10083 25989
rect 10118 25955 10152 25989
rect 10187 25955 10221 25989
rect 10256 25955 10290 25989
rect 10325 25955 10359 25989
rect 10394 25955 10428 25989
rect 10463 25955 10497 25989
rect 10532 25955 10566 25989
rect 10601 25955 10635 25989
rect 10670 25955 10704 25989
rect 10739 25955 10773 25989
rect 10807 25955 10841 25989
rect 10875 25955 10909 25989
rect 10943 25955 10977 25989
rect 11011 25955 11045 25989
rect 11079 25955 11113 25989
rect 11147 25955 11181 25989
rect 11215 25955 11249 25989
rect 11283 25955 11317 25989
rect 11351 25955 11385 25989
rect 11419 25955 11453 25989
rect 11487 25955 11521 25989
rect 11555 25955 11589 25989
rect 11623 25955 11657 25989
rect 11691 25955 11725 25989
rect 11759 25955 11793 25989
rect 11827 25955 11861 25989
rect 11895 25955 11929 25989
rect 11963 25955 11997 25989
rect 12031 25955 12065 25989
rect 12099 25955 12133 25989
rect 12167 25955 12201 25989
rect 12235 25955 12269 25989
rect 12303 25955 12337 25989
rect 12371 25955 12405 25989
rect 12439 25955 12473 25989
rect 12507 25955 12541 25989
rect 12575 25955 12609 25989
rect 12643 25955 12677 25989
rect 12711 25955 12745 25989
rect 12779 25955 12813 25989
rect 12847 25955 12881 25989
rect 12915 25955 12949 25989
rect 12983 25955 13017 25989
rect 13051 25955 13085 25989
rect 13119 25955 13153 25989
rect 13187 25955 13221 25989
rect 13255 25955 13289 25989
rect 13323 25955 13357 25989
rect 13391 25955 13425 25989
rect 13459 25955 13493 25989
rect 13527 25955 13561 25989
rect 13595 25955 13629 25989
rect 13663 25955 13697 25989
rect 13731 25955 13765 25989
rect 13799 25955 13833 25989
rect 13867 25955 13901 25989
rect 13935 25955 13969 25989
rect 14003 25955 14037 25989
rect 14071 25955 14105 25989
rect 14139 25955 14173 25989
rect 9911 25885 9945 25919
rect 9980 25885 10014 25919
rect 10049 25885 10083 25919
rect 10118 25885 10152 25919
rect 10187 25885 10221 25919
rect 10256 25885 10290 25919
rect 10325 25885 10359 25919
rect 10394 25885 10428 25919
rect 10463 25885 10497 25919
rect 10532 25885 10566 25919
rect 10601 25885 10635 25919
rect 10670 25885 10704 25919
rect 10739 25885 10773 25919
rect 10807 25885 10841 25919
rect 10875 25885 10909 25919
rect 10943 25885 10977 25919
rect 11011 25885 11045 25919
rect 11079 25885 11113 25919
rect 11147 25885 11181 25919
rect 11215 25885 11249 25919
rect 11283 25885 11317 25919
rect 11351 25885 11385 25919
rect 11419 25885 11453 25919
rect 11487 25885 11521 25919
rect 11555 25885 11589 25919
rect 11623 25885 11657 25919
rect 11691 25885 11725 25919
rect 11759 25885 11793 25919
rect 11827 25885 11861 25919
rect 11895 25885 11929 25919
rect 11963 25885 11997 25919
rect 12031 25885 12065 25919
rect 12099 25885 12133 25919
rect 12167 25885 12201 25919
rect 12235 25885 12269 25919
rect 12303 25885 12337 25919
rect 12371 25885 12405 25919
rect 12439 25885 12473 25919
rect 12507 25885 12541 25919
rect 12575 25885 12609 25919
rect 12643 25885 12677 25919
rect 12711 25885 12745 25919
rect 12779 25885 12813 25919
rect 12847 25885 12881 25919
rect 12915 25885 12949 25919
rect 12983 25885 13017 25919
rect 13051 25885 13085 25919
rect 13119 25885 13153 25919
rect 13187 25885 13221 25919
rect 13255 25885 13289 25919
rect 13323 25885 13357 25919
rect 13391 25885 13425 25919
rect 13459 25885 13493 25919
rect 13527 25885 13561 25919
rect 13595 25885 13629 25919
rect 13663 25885 13697 25919
rect 13731 25885 13765 25919
rect 13799 25885 13833 25919
rect 13867 25885 13901 25919
rect 13935 25885 13969 25919
rect 14003 25885 14037 25919
rect 14071 25885 14105 25919
rect 14139 25885 14173 25919
rect 9911 25815 9945 25849
rect 9980 25815 10014 25849
rect 10049 25815 10083 25849
rect 10118 25815 10152 25849
rect 10187 25815 10221 25849
rect 10256 25815 10290 25849
rect 10325 25815 10359 25849
rect 10394 25815 10428 25849
rect 10463 25815 10497 25849
rect 10532 25815 10566 25849
rect 10601 25815 10635 25849
rect 10670 25815 10704 25849
rect 10739 25815 10773 25849
rect 10807 25815 10841 25849
rect 10875 25815 10909 25849
rect 10943 25815 10977 25849
rect 11011 25815 11045 25849
rect 11079 25815 11113 25849
rect 11147 25815 11181 25849
rect 11215 25815 11249 25849
rect 11283 25815 11317 25849
rect 11351 25815 11385 25849
rect 11419 25815 11453 25849
rect 11487 25815 11521 25849
rect 11555 25815 11589 25849
rect 11623 25815 11657 25849
rect 11691 25815 11725 25849
rect 11759 25815 11793 25849
rect 11827 25815 11861 25849
rect 11895 25815 11929 25849
rect 11963 25815 11997 25849
rect 12031 25815 12065 25849
rect 12099 25815 12133 25849
rect 12167 25815 12201 25849
rect 12235 25815 12269 25849
rect 12303 25815 12337 25849
rect 12371 25815 12405 25849
rect 12439 25815 12473 25849
rect 12507 25815 12541 25849
rect 12575 25815 12609 25849
rect 12643 25815 12677 25849
rect 12711 25815 12745 25849
rect 12779 25815 12813 25849
rect 12847 25815 12881 25849
rect 12915 25815 12949 25849
rect 12983 25815 13017 25849
rect 13051 25815 13085 25849
rect 13119 25815 13153 25849
rect 13187 25815 13221 25849
rect 13255 25815 13289 25849
rect 13323 25815 13357 25849
rect 13391 25815 13425 25849
rect 13459 25815 13493 25849
rect 13527 25815 13561 25849
rect 13595 25815 13629 25849
rect 13663 25815 13697 25849
rect 13731 25815 13765 25849
rect 13799 25815 13833 25849
rect 13867 25815 13901 25849
rect 13935 25815 13969 25849
rect 14003 25815 14037 25849
rect 14071 25815 14105 25849
rect 14139 25815 14173 25849
rect 9911 25745 9945 25779
rect 9980 25745 10014 25779
rect 10049 25745 10083 25779
rect 10118 25745 10152 25779
rect 10187 25745 10221 25779
rect 10256 25745 10290 25779
rect 10325 25745 10359 25779
rect 10394 25745 10428 25779
rect 10463 25745 10497 25779
rect 10532 25745 10566 25779
rect 10601 25745 10635 25779
rect 10670 25745 10704 25779
rect 10739 25745 10773 25779
rect 10807 25745 10841 25779
rect 10875 25745 10909 25779
rect 10943 25745 10977 25779
rect 11011 25745 11045 25779
rect 11079 25745 11113 25779
rect 11147 25745 11181 25779
rect 11215 25745 11249 25779
rect 11283 25745 11317 25779
rect 11351 25745 11385 25779
rect 11419 25745 11453 25779
rect 11487 25745 11521 25779
rect 11555 25745 11589 25779
rect 11623 25745 11657 25779
rect 11691 25745 11725 25779
rect 11759 25745 11793 25779
rect 11827 25745 11861 25779
rect 11895 25745 11929 25779
rect 11963 25745 11997 25779
rect 12031 25745 12065 25779
rect 12099 25745 12133 25779
rect 12167 25745 12201 25779
rect 12235 25745 12269 25779
rect 12303 25745 12337 25779
rect 12371 25745 12405 25779
rect 12439 25745 12473 25779
rect 12507 25745 12541 25779
rect 12575 25745 12609 25779
rect 12643 25745 12677 25779
rect 12711 25745 12745 25779
rect 12779 25745 12813 25779
rect 12847 25745 12881 25779
rect 12915 25745 12949 25779
rect 12983 25745 13017 25779
rect 13051 25745 13085 25779
rect 13119 25745 13153 25779
rect 13187 25745 13221 25779
rect 13255 25745 13289 25779
rect 13323 25745 13357 25779
rect 13391 25745 13425 25779
rect 13459 25745 13493 25779
rect 13527 25745 13561 25779
rect 13595 25745 13629 25779
rect 13663 25745 13697 25779
rect 13731 25745 13765 25779
rect 13799 25745 13833 25779
rect 13867 25745 13901 25779
rect 13935 25745 13969 25779
rect 14003 25745 14037 25779
rect 14071 25745 14105 25779
rect 14139 25745 14173 25779
rect 9911 25675 9945 25709
rect 9980 25675 10014 25709
rect 10049 25675 10083 25709
rect 10118 25675 10152 25709
rect 10187 25675 10221 25709
rect 10256 25675 10290 25709
rect 10325 25675 10359 25709
rect 10394 25675 10428 25709
rect 10463 25675 10497 25709
rect 10532 25675 10566 25709
rect 10601 25675 10635 25709
rect 10670 25675 10704 25709
rect 10739 25675 10773 25709
rect 10807 25675 10841 25709
rect 10875 25675 10909 25709
rect 10943 25675 10977 25709
rect 11011 25675 11045 25709
rect 11079 25675 11113 25709
rect 11147 25675 11181 25709
rect 11215 25675 11249 25709
rect 11283 25675 11317 25709
rect 11351 25675 11385 25709
rect 11419 25675 11453 25709
rect 11487 25675 11521 25709
rect 11555 25675 11589 25709
rect 11623 25675 11657 25709
rect 11691 25675 11725 25709
rect 11759 25675 11793 25709
rect 11827 25675 11861 25709
rect 11895 25675 11929 25709
rect 11963 25675 11997 25709
rect 12031 25675 12065 25709
rect 12099 25675 12133 25709
rect 12167 25675 12201 25709
rect 12235 25675 12269 25709
rect 12303 25675 12337 25709
rect 12371 25675 12405 25709
rect 12439 25675 12473 25709
rect 12507 25675 12541 25709
rect 12575 25675 12609 25709
rect 12643 25675 12677 25709
rect 12711 25675 12745 25709
rect 12779 25675 12813 25709
rect 12847 25675 12881 25709
rect 12915 25675 12949 25709
rect 12983 25675 13017 25709
rect 13051 25675 13085 25709
rect 13119 25675 13153 25709
rect 13187 25675 13221 25709
rect 13255 25675 13289 25709
rect 13323 25675 13357 25709
rect 13391 25675 13425 25709
rect 13459 25675 13493 25709
rect 13527 25675 13561 25709
rect 13595 25675 13629 25709
rect 13663 25675 13697 25709
rect 13731 25675 13765 25709
rect 13799 25675 13833 25709
rect 13867 25675 13901 25709
rect 13935 25675 13969 25709
rect 14003 25675 14037 25709
rect 14071 25675 14105 25709
rect 14139 25675 14173 25709
rect 9911 25605 9945 25639
rect 9980 25605 10014 25639
rect 10049 25605 10083 25639
rect 10118 25605 10152 25639
rect 10187 25605 10221 25639
rect 10256 25605 10290 25639
rect 10325 25605 10359 25639
rect 10394 25605 10428 25639
rect 10463 25605 10497 25639
rect 10532 25605 10566 25639
rect 10601 25605 10635 25639
rect 10670 25605 10704 25639
rect 10739 25605 10773 25639
rect 10807 25605 10841 25639
rect 10875 25605 10909 25639
rect 10943 25605 10977 25639
rect 11011 25605 11045 25639
rect 11079 25605 11113 25639
rect 11147 25605 11181 25639
rect 11215 25605 11249 25639
rect 11283 25605 11317 25639
rect 11351 25605 11385 25639
rect 11419 25605 11453 25639
rect 11487 25605 11521 25639
rect 11555 25605 11589 25639
rect 11623 25605 11657 25639
rect 11691 25605 11725 25639
rect 11759 25605 11793 25639
rect 11827 25605 11861 25639
rect 11895 25605 11929 25639
rect 11963 25605 11997 25639
rect 12031 25605 12065 25639
rect 12099 25605 12133 25639
rect 12167 25605 12201 25639
rect 12235 25605 12269 25639
rect 12303 25605 12337 25639
rect 12371 25605 12405 25639
rect 12439 25605 12473 25639
rect 12507 25605 12541 25639
rect 12575 25605 12609 25639
rect 12643 25605 12677 25639
rect 12711 25605 12745 25639
rect 12779 25605 12813 25639
rect 12847 25605 12881 25639
rect 12915 25605 12949 25639
rect 12983 25605 13017 25639
rect 13051 25605 13085 25639
rect 13119 25605 13153 25639
rect 13187 25605 13221 25639
rect 13255 25605 13289 25639
rect 13323 25605 13357 25639
rect 13391 25605 13425 25639
rect 13459 25605 13493 25639
rect 13527 25605 13561 25639
rect 13595 25605 13629 25639
rect 13663 25605 13697 25639
rect 13731 25605 13765 25639
rect 13799 25605 13833 25639
rect 13867 25605 13901 25639
rect 13935 25605 13969 25639
rect 14003 25605 14037 25639
rect 14071 25605 14105 25639
rect 14139 25605 14173 25639
rect 9911 25535 9945 25569
rect 9980 25535 10014 25569
rect 10049 25535 10083 25569
rect 10118 25535 10152 25569
rect 10187 25535 10221 25569
rect 10256 25535 10290 25569
rect 10325 25535 10359 25569
rect 10394 25535 10428 25569
rect 10463 25535 10497 25569
rect 10532 25535 10566 25569
rect 10601 25535 10635 25569
rect 10670 25535 10704 25569
rect 10739 25535 10773 25569
rect 10807 25535 10841 25569
rect 10875 25535 10909 25569
rect 10943 25535 10977 25569
rect 11011 25535 11045 25569
rect 11079 25535 11113 25569
rect 11147 25535 11181 25569
rect 11215 25535 11249 25569
rect 11283 25535 11317 25569
rect 11351 25535 11385 25569
rect 11419 25535 11453 25569
rect 11487 25535 11521 25569
rect 11555 25535 11589 25569
rect 11623 25535 11657 25569
rect 11691 25535 11725 25569
rect 11759 25535 11793 25569
rect 11827 25535 11861 25569
rect 11895 25535 11929 25569
rect 11963 25535 11997 25569
rect 12031 25535 12065 25569
rect 12099 25535 12133 25569
rect 12167 25535 12201 25569
rect 12235 25535 12269 25569
rect 12303 25535 12337 25569
rect 12371 25535 12405 25569
rect 12439 25535 12473 25569
rect 12507 25535 12541 25569
rect 12575 25535 12609 25569
rect 12643 25535 12677 25569
rect 12711 25535 12745 25569
rect 12779 25535 12813 25569
rect 12847 25535 12881 25569
rect 12915 25535 12949 25569
rect 12983 25535 13017 25569
rect 13051 25535 13085 25569
rect 13119 25535 13153 25569
rect 13187 25535 13221 25569
rect 13255 25535 13289 25569
rect 13323 25535 13357 25569
rect 13391 25535 13425 25569
rect 13459 25535 13493 25569
rect 13527 25535 13561 25569
rect 13595 25535 13629 25569
rect 13663 25535 13697 25569
rect 13731 25535 13765 25569
rect 13799 25535 13833 25569
rect 13867 25535 13901 25569
rect 13935 25535 13969 25569
rect 14003 25535 14037 25569
rect 14071 25535 14105 25569
rect 14139 25535 14173 25569
rect 9911 25465 9945 25499
rect 9980 25465 10014 25499
rect 10049 25465 10083 25499
rect 10118 25465 10152 25499
rect 10187 25465 10221 25499
rect 10256 25465 10290 25499
rect 10325 25465 10359 25499
rect 10394 25465 10428 25499
rect 10463 25465 10497 25499
rect 10532 25465 10566 25499
rect 10601 25465 10635 25499
rect 10670 25465 10704 25499
rect 10739 25465 10773 25499
rect 10807 25465 10841 25499
rect 10875 25465 10909 25499
rect 10943 25465 10977 25499
rect 11011 25465 11045 25499
rect 11079 25465 11113 25499
rect 11147 25465 11181 25499
rect 11215 25465 11249 25499
rect 11283 25465 11317 25499
rect 11351 25465 11385 25499
rect 11419 25465 11453 25499
rect 11487 25465 11521 25499
rect 11555 25465 11589 25499
rect 11623 25465 11657 25499
rect 11691 25465 11725 25499
rect 11759 25465 11793 25499
rect 11827 25465 11861 25499
rect 11895 25465 11929 25499
rect 11963 25465 11997 25499
rect 12031 25465 12065 25499
rect 12099 25465 12133 25499
rect 12167 25465 12201 25499
rect 12235 25465 12269 25499
rect 12303 25465 12337 25499
rect 12371 25465 12405 25499
rect 12439 25465 12473 25499
rect 12507 25465 12541 25499
rect 12575 25465 12609 25499
rect 12643 25465 12677 25499
rect 12711 25465 12745 25499
rect 12779 25465 12813 25499
rect 12847 25465 12881 25499
rect 12915 25465 12949 25499
rect 12983 25465 13017 25499
rect 13051 25465 13085 25499
rect 13119 25465 13153 25499
rect 13187 25465 13221 25499
rect 13255 25465 13289 25499
rect 13323 25465 13357 25499
rect 13391 25465 13425 25499
rect 13459 25465 13493 25499
rect 13527 25465 13561 25499
rect 13595 25465 13629 25499
rect 13663 25465 13697 25499
rect 13731 25465 13765 25499
rect 13799 25465 13833 25499
rect 13867 25465 13901 25499
rect 13935 25465 13969 25499
rect 14003 25465 14037 25499
rect 14071 25465 14105 25499
rect 14139 25465 14173 25499
rect 9911 25395 9945 25429
rect 9980 25395 10014 25429
rect 10049 25395 10083 25429
rect 10118 25395 10152 25429
rect 10187 25395 10221 25429
rect 10256 25395 10290 25429
rect 10325 25395 10359 25429
rect 10394 25395 10428 25429
rect 10463 25395 10497 25429
rect 10532 25395 10566 25429
rect 10601 25395 10635 25429
rect 10670 25395 10704 25429
rect 10739 25395 10773 25429
rect 10807 25395 10841 25429
rect 10875 25395 10909 25429
rect 10943 25395 10977 25429
rect 11011 25395 11045 25429
rect 11079 25395 11113 25429
rect 11147 25395 11181 25429
rect 11215 25395 11249 25429
rect 11283 25395 11317 25429
rect 11351 25395 11385 25429
rect 11419 25395 11453 25429
rect 11487 25395 11521 25429
rect 11555 25395 11589 25429
rect 11623 25395 11657 25429
rect 11691 25395 11725 25429
rect 11759 25395 11793 25429
rect 11827 25395 11861 25429
rect 11895 25395 11929 25429
rect 11963 25395 11997 25429
rect 12031 25395 12065 25429
rect 12099 25395 12133 25429
rect 12167 25395 12201 25429
rect 12235 25395 12269 25429
rect 12303 25395 12337 25429
rect 12371 25395 12405 25429
rect 12439 25395 12473 25429
rect 12507 25395 12541 25429
rect 12575 25395 12609 25429
rect 12643 25395 12677 25429
rect 12711 25395 12745 25429
rect 12779 25395 12813 25429
rect 12847 25395 12881 25429
rect 12915 25395 12949 25429
rect 12983 25395 13017 25429
rect 13051 25395 13085 25429
rect 13119 25395 13153 25429
rect 13187 25395 13221 25429
rect 13255 25395 13289 25429
rect 13323 25395 13357 25429
rect 13391 25395 13425 25429
rect 13459 25395 13493 25429
rect 13527 25395 13561 25429
rect 13595 25395 13629 25429
rect 13663 25395 13697 25429
rect 13731 25395 13765 25429
rect 13799 25395 13833 25429
rect 13867 25395 13901 25429
rect 13935 25395 13969 25429
rect 14003 25395 14037 25429
rect 14071 25395 14105 25429
rect 14139 25395 14173 25429
rect 9911 25325 9945 25359
rect 9980 25325 10014 25359
rect 10049 25325 10083 25359
rect 10118 25325 10152 25359
rect 10187 25325 10221 25359
rect 10256 25325 10290 25359
rect 10325 25325 10359 25359
rect 10394 25325 10428 25359
rect 10463 25325 10497 25359
rect 10532 25325 10566 25359
rect 10601 25325 10635 25359
rect 10670 25325 10704 25359
rect 10739 25325 10773 25359
rect 10807 25325 10841 25359
rect 10875 25325 10909 25359
rect 10943 25325 10977 25359
rect 11011 25325 11045 25359
rect 11079 25325 11113 25359
rect 11147 25325 11181 25359
rect 11215 25325 11249 25359
rect 11283 25325 11317 25359
rect 11351 25325 11385 25359
rect 11419 25325 11453 25359
rect 11487 25325 11521 25359
rect 11555 25325 11589 25359
rect 11623 25325 11657 25359
rect 11691 25325 11725 25359
rect 11759 25325 11793 25359
rect 11827 25325 11861 25359
rect 11895 25325 11929 25359
rect 11963 25325 11997 25359
rect 12031 25325 12065 25359
rect 12099 25325 12133 25359
rect 12167 25325 12201 25359
rect 12235 25325 12269 25359
rect 12303 25325 12337 25359
rect 12371 25325 12405 25359
rect 12439 25325 12473 25359
rect 12507 25325 12541 25359
rect 12575 25325 12609 25359
rect 12643 25325 12677 25359
rect 12711 25325 12745 25359
rect 12779 25325 12813 25359
rect 12847 25325 12881 25359
rect 12915 25325 12949 25359
rect 12983 25325 13017 25359
rect 13051 25325 13085 25359
rect 13119 25325 13153 25359
rect 13187 25325 13221 25359
rect 13255 25325 13289 25359
rect 13323 25325 13357 25359
rect 13391 25325 13425 25359
rect 13459 25325 13493 25359
rect 13527 25325 13561 25359
rect 13595 25325 13629 25359
rect 13663 25325 13697 25359
rect 13731 25325 13765 25359
rect 13799 25325 13833 25359
rect 13867 25325 13901 25359
rect 13935 25325 13969 25359
rect 14003 25325 14037 25359
rect 14071 25325 14105 25359
rect 14139 25325 14173 25359
rect 9911 25255 9945 25289
rect 9980 25255 10014 25289
rect 10049 25255 10083 25289
rect 10118 25255 10152 25289
rect 10187 25255 10221 25289
rect 10256 25255 10290 25289
rect 10325 25255 10359 25289
rect 10394 25255 10428 25289
rect 10463 25255 10497 25289
rect 10532 25255 10566 25289
rect 10601 25255 10635 25289
rect 10670 25255 10704 25289
rect 10739 25255 10773 25289
rect 10807 25255 10841 25289
rect 10875 25255 10909 25289
rect 10943 25255 10977 25289
rect 11011 25255 11045 25289
rect 11079 25255 11113 25289
rect 11147 25255 11181 25289
rect 11215 25255 11249 25289
rect 11283 25255 11317 25289
rect 11351 25255 11385 25289
rect 11419 25255 11453 25289
rect 11487 25255 11521 25289
rect 11555 25255 11589 25289
rect 11623 25255 11657 25289
rect 11691 25255 11725 25289
rect 11759 25255 11793 25289
rect 11827 25255 11861 25289
rect 11895 25255 11929 25289
rect 11963 25255 11997 25289
rect 12031 25255 12065 25289
rect 12099 25255 12133 25289
rect 12167 25255 12201 25289
rect 12235 25255 12269 25289
rect 12303 25255 12337 25289
rect 12371 25255 12405 25289
rect 12439 25255 12473 25289
rect 12507 25255 12541 25289
rect 12575 25255 12609 25289
rect 12643 25255 12677 25289
rect 12711 25255 12745 25289
rect 12779 25255 12813 25289
rect 12847 25255 12881 25289
rect 12915 25255 12949 25289
rect 12983 25255 13017 25289
rect 13051 25255 13085 25289
rect 13119 25255 13153 25289
rect 13187 25255 13221 25289
rect 13255 25255 13289 25289
rect 13323 25255 13357 25289
rect 13391 25255 13425 25289
rect 13459 25255 13493 25289
rect 13527 25255 13561 25289
rect 13595 25255 13629 25289
rect 13663 25255 13697 25289
rect 13731 25255 13765 25289
rect 13799 25255 13833 25289
rect 13867 25255 13901 25289
rect 13935 25255 13969 25289
rect 14003 25255 14037 25289
rect 14071 25255 14105 25289
rect 14139 25255 14173 25289
rect 9911 25185 9945 25219
rect 9980 25185 10014 25219
rect 10049 25185 10083 25219
rect 10118 25185 10152 25219
rect 10187 25185 10221 25219
rect 10256 25185 10290 25219
rect 10325 25185 10359 25219
rect 10394 25185 10428 25219
rect 10463 25185 10497 25219
rect 10532 25185 10566 25219
rect 10601 25185 10635 25219
rect 10670 25185 10704 25219
rect 10739 25185 10773 25219
rect 10807 25185 10841 25219
rect 10875 25185 10909 25219
rect 10943 25185 10977 25219
rect 11011 25185 11045 25219
rect 11079 25185 11113 25219
rect 11147 25185 11181 25219
rect 11215 25185 11249 25219
rect 11283 25185 11317 25219
rect 11351 25185 11385 25219
rect 11419 25185 11453 25219
rect 11487 25185 11521 25219
rect 11555 25185 11589 25219
rect 11623 25185 11657 25219
rect 11691 25185 11725 25219
rect 11759 25185 11793 25219
rect 11827 25185 11861 25219
rect 11895 25185 11929 25219
rect 11963 25185 11997 25219
rect 12031 25185 12065 25219
rect 12099 25185 12133 25219
rect 12167 25185 12201 25219
rect 12235 25185 12269 25219
rect 12303 25185 12337 25219
rect 12371 25185 12405 25219
rect 12439 25185 12473 25219
rect 12507 25185 12541 25219
rect 12575 25185 12609 25219
rect 12643 25185 12677 25219
rect 12711 25185 12745 25219
rect 12779 25185 12813 25219
rect 12847 25185 12881 25219
rect 12915 25185 12949 25219
rect 12983 25185 13017 25219
rect 13051 25185 13085 25219
rect 13119 25185 13153 25219
rect 13187 25185 13221 25219
rect 13255 25185 13289 25219
rect 13323 25185 13357 25219
rect 13391 25185 13425 25219
rect 13459 25185 13493 25219
rect 13527 25185 13561 25219
rect 13595 25185 13629 25219
rect 13663 25185 13697 25219
rect 13731 25185 13765 25219
rect 13799 25185 13833 25219
rect 13867 25185 13901 25219
rect 13935 25185 13969 25219
rect 14003 25185 14037 25219
rect 14071 25185 14105 25219
rect 14139 25185 14173 25219
rect 9911 25115 9945 25149
rect 9980 25115 10014 25149
rect 10049 25115 10083 25149
rect 10118 25115 10152 25149
rect 10187 25115 10221 25149
rect 10256 25115 10290 25149
rect 10325 25115 10359 25149
rect 10394 25115 10428 25149
rect 10463 25115 10497 25149
rect 10532 25115 10566 25149
rect 10601 25115 10635 25149
rect 10670 25115 10704 25149
rect 10739 25115 10773 25149
rect 10807 25115 10841 25149
rect 10875 25115 10909 25149
rect 10943 25115 10977 25149
rect 11011 25115 11045 25149
rect 11079 25115 11113 25149
rect 11147 25115 11181 25149
rect 11215 25115 11249 25149
rect 11283 25115 11317 25149
rect 11351 25115 11385 25149
rect 11419 25115 11453 25149
rect 11487 25115 11521 25149
rect 11555 25115 11589 25149
rect 11623 25115 11657 25149
rect 11691 25115 11725 25149
rect 11759 25115 11793 25149
rect 11827 25115 11861 25149
rect 11895 25115 11929 25149
rect 11963 25115 11997 25149
rect 12031 25115 12065 25149
rect 12099 25115 12133 25149
rect 12167 25115 12201 25149
rect 12235 25115 12269 25149
rect 12303 25115 12337 25149
rect 12371 25115 12405 25149
rect 12439 25115 12473 25149
rect 12507 25115 12541 25149
rect 12575 25115 12609 25149
rect 12643 25115 12677 25149
rect 12711 25115 12745 25149
rect 12779 25115 12813 25149
rect 12847 25115 12881 25149
rect 12915 25115 12949 25149
rect 12983 25115 13017 25149
rect 13051 25115 13085 25149
rect 13119 25115 13153 25149
rect 13187 25115 13221 25149
rect 13255 25115 13289 25149
rect 13323 25115 13357 25149
rect 13391 25115 13425 25149
rect 13459 25115 13493 25149
rect 13527 25115 13561 25149
rect 13595 25115 13629 25149
rect 13663 25115 13697 25149
rect 13731 25115 13765 25149
rect 13799 25115 13833 25149
rect 13867 25115 13901 25149
rect 13935 25115 13969 25149
rect 14003 25115 14037 25149
rect 14071 25115 14105 25149
rect 14139 25115 14173 25149
rect 9911 25045 9945 25079
rect 9980 25045 10014 25079
rect 10049 25045 10083 25079
rect 10118 25045 10152 25079
rect 10187 25045 10221 25079
rect 10256 25045 10290 25079
rect 10325 25045 10359 25079
rect 10394 25045 10428 25079
rect 10463 25045 10497 25079
rect 10532 25045 10566 25079
rect 10601 25045 10635 25079
rect 10670 25045 10704 25079
rect 10739 25045 10773 25079
rect 10807 25045 10841 25079
rect 10875 25045 10909 25079
rect 10943 25045 10977 25079
rect 11011 25045 11045 25079
rect 11079 25045 11113 25079
rect 11147 25045 11181 25079
rect 11215 25045 11249 25079
rect 11283 25045 11317 25079
rect 11351 25045 11385 25079
rect 11419 25045 11453 25079
rect 11487 25045 11521 25079
rect 11555 25045 11589 25079
rect 11623 25045 11657 25079
rect 11691 25045 11725 25079
rect 11759 25045 11793 25079
rect 11827 25045 11861 25079
rect 11895 25045 11929 25079
rect 11963 25045 11997 25079
rect 12031 25045 12065 25079
rect 12099 25045 12133 25079
rect 12167 25045 12201 25079
rect 12235 25045 12269 25079
rect 12303 25045 12337 25079
rect 12371 25045 12405 25079
rect 12439 25045 12473 25079
rect 12507 25045 12541 25079
rect 12575 25045 12609 25079
rect 12643 25045 12677 25079
rect 12711 25045 12745 25079
rect 12779 25045 12813 25079
rect 12847 25045 12881 25079
rect 12915 25045 12949 25079
rect 12983 25045 13017 25079
rect 13051 25045 13085 25079
rect 13119 25045 13153 25079
rect 13187 25045 13221 25079
rect 13255 25045 13289 25079
rect 13323 25045 13357 25079
rect 13391 25045 13425 25079
rect 13459 25045 13493 25079
rect 13527 25045 13561 25079
rect 13595 25045 13629 25079
rect 13663 25045 13697 25079
rect 13731 25045 13765 25079
rect 13799 25045 13833 25079
rect 13867 25045 13901 25079
rect 13935 25045 13969 25079
rect 14003 25045 14037 25079
rect 14071 25045 14105 25079
rect 14139 25045 14173 25079
rect 9911 24975 9945 25009
rect 9980 24975 10014 25009
rect 10049 24975 10083 25009
rect 10118 24975 10152 25009
rect 10187 24975 10221 25009
rect 10256 24975 10290 25009
rect 10325 24975 10359 25009
rect 10394 24975 10428 25009
rect 10463 24975 10497 25009
rect 10532 24975 10566 25009
rect 10601 24975 10635 25009
rect 10670 24975 10704 25009
rect 10739 24975 10773 25009
rect 10807 24975 10841 25009
rect 10875 24975 10909 25009
rect 10943 24975 10977 25009
rect 11011 24975 11045 25009
rect 11079 24975 11113 25009
rect 11147 24975 11181 25009
rect 11215 24975 11249 25009
rect 11283 24975 11317 25009
rect 11351 24975 11385 25009
rect 11419 24975 11453 25009
rect 11487 24975 11521 25009
rect 11555 24975 11589 25009
rect 11623 24975 11657 25009
rect 11691 24975 11725 25009
rect 11759 24975 11793 25009
rect 11827 24975 11861 25009
rect 11895 24975 11929 25009
rect 11963 24975 11997 25009
rect 12031 24975 12065 25009
rect 12099 24975 12133 25009
rect 12167 24975 12201 25009
rect 12235 24975 12269 25009
rect 12303 24975 12337 25009
rect 12371 24975 12405 25009
rect 12439 24975 12473 25009
rect 12507 24975 12541 25009
rect 12575 24975 12609 25009
rect 12643 24975 12677 25009
rect 12711 24975 12745 25009
rect 12779 24975 12813 25009
rect 12847 24975 12881 25009
rect 12915 24975 12949 25009
rect 12983 24975 13017 25009
rect 13051 24975 13085 25009
rect 13119 24975 13153 25009
rect 13187 24975 13221 25009
rect 13255 24975 13289 25009
rect 13323 24975 13357 25009
rect 13391 24975 13425 25009
rect 13459 24975 13493 25009
rect 13527 24975 13561 25009
rect 13595 24975 13629 25009
rect 13663 24975 13697 25009
rect 13731 24975 13765 25009
rect 13799 24975 13833 25009
rect 13867 24975 13901 25009
rect 13935 24975 13969 25009
rect 14003 24975 14037 25009
rect 14071 24975 14105 25009
rect 14139 24975 14173 25009
rect 9911 24905 9945 24939
rect 9980 24905 10014 24939
rect 10049 24905 10083 24939
rect 10118 24905 10152 24939
rect 10187 24905 10221 24939
rect 10256 24905 10290 24939
rect 10325 24905 10359 24939
rect 10394 24905 10428 24939
rect 10463 24905 10497 24939
rect 10532 24905 10566 24939
rect 10601 24905 10635 24939
rect 10670 24905 10704 24939
rect 10739 24905 10773 24939
rect 10807 24905 10841 24939
rect 10875 24905 10909 24939
rect 10943 24905 10977 24939
rect 11011 24905 11045 24939
rect 11079 24905 11113 24939
rect 11147 24905 11181 24939
rect 11215 24905 11249 24939
rect 11283 24905 11317 24939
rect 11351 24905 11385 24939
rect 11419 24905 11453 24939
rect 11487 24905 11521 24939
rect 11555 24905 11589 24939
rect 11623 24905 11657 24939
rect 11691 24905 11725 24939
rect 11759 24905 11793 24939
rect 11827 24905 11861 24939
rect 11895 24905 11929 24939
rect 11963 24905 11997 24939
rect 12031 24905 12065 24939
rect 12099 24905 12133 24939
rect 12167 24905 12201 24939
rect 12235 24905 12269 24939
rect 12303 24905 12337 24939
rect 12371 24905 12405 24939
rect 12439 24905 12473 24939
rect 12507 24905 12541 24939
rect 12575 24905 12609 24939
rect 12643 24905 12677 24939
rect 12711 24905 12745 24939
rect 12779 24905 12813 24939
rect 12847 24905 12881 24939
rect 12915 24905 12949 24939
rect 12983 24905 13017 24939
rect 13051 24905 13085 24939
rect 13119 24905 13153 24939
rect 13187 24905 13221 24939
rect 13255 24905 13289 24939
rect 13323 24905 13357 24939
rect 13391 24905 13425 24939
rect 13459 24905 13493 24939
rect 13527 24905 13561 24939
rect 13595 24905 13629 24939
rect 13663 24905 13697 24939
rect 13731 24905 13765 24939
rect 13799 24905 13833 24939
rect 13867 24905 13901 24939
rect 13935 24905 13969 24939
rect 14003 24905 14037 24939
rect 14071 24905 14105 24939
rect 14139 24905 14173 24939
rect 9911 24787 9945 24821
rect 9981 24787 10015 24821
rect 10051 24787 10085 24821
rect 10121 24787 10155 24821
rect 10191 24787 10225 24821
rect 10261 24787 10295 24821
rect 10331 24787 10365 24821
rect 10401 24787 10435 24821
rect 10471 24787 10505 24821
rect 10541 24787 10575 24821
rect 10611 24787 10645 24821
rect 10681 24787 10715 24821
rect 10750 24787 10784 24821
rect 10819 24787 10853 24821
rect 10888 24787 10922 24821
rect 10957 24787 10991 24821
rect 11026 24787 11060 24821
rect 11095 24787 11129 24821
rect 11164 24787 11198 24821
rect 9911 24719 9945 24753
rect 9981 24719 10015 24753
rect 10051 24719 10085 24753
rect 10121 24719 10155 24753
rect 10191 24719 10225 24753
rect 10261 24719 10295 24753
rect 10331 24719 10365 24753
rect 10401 24719 10435 24753
rect 10471 24719 10505 24753
rect 10541 24719 10575 24753
rect 10611 24719 10645 24753
rect 10681 24719 10715 24753
rect 10750 24719 10784 24753
rect 10819 24719 10853 24753
rect 10888 24719 10922 24753
rect 10957 24719 10991 24753
rect 11026 24719 11060 24753
rect 11095 24719 11129 24753
rect 11164 24719 11198 24753
rect 9911 24651 9945 24685
rect 9981 24651 10015 24685
rect 10051 24651 10085 24685
rect 10121 24651 10155 24685
rect 10191 24651 10225 24685
rect 10261 24651 10295 24685
rect 10331 24651 10365 24685
rect 10401 24651 10435 24685
rect 10471 24651 10505 24685
rect 10541 24651 10575 24685
rect 10611 24651 10645 24685
rect 10681 24651 10715 24685
rect 10750 24651 10784 24685
rect 10819 24651 10853 24685
rect 10888 24651 10922 24685
rect 10957 24651 10991 24685
rect 11026 24651 11060 24685
rect 11095 24651 11129 24685
rect 11164 24651 11198 24685
rect 9911 24583 9945 24617
rect 9981 24583 10015 24617
rect 10051 24583 10085 24617
rect 10121 24583 10155 24617
rect 10191 24583 10225 24617
rect 10261 24583 10295 24617
rect 10331 24583 10365 24617
rect 10401 24583 10435 24617
rect 10471 24583 10505 24617
rect 10541 24583 10575 24617
rect 10611 24583 10645 24617
rect 10681 24583 10715 24617
rect 10750 24583 10784 24617
rect 10819 24583 10853 24617
rect 10888 24583 10922 24617
rect 10957 24583 10991 24617
rect 11026 24583 11060 24617
rect 11095 24583 11129 24617
rect 11164 24583 11198 24617
rect 9911 24515 9945 24549
rect 9981 24515 10015 24549
rect 10051 24515 10085 24549
rect 10121 24515 10155 24549
rect 10191 24515 10225 24549
rect 10261 24515 10295 24549
rect 10331 24515 10365 24549
rect 10401 24515 10435 24549
rect 10471 24515 10505 24549
rect 10541 24515 10575 24549
rect 10611 24515 10645 24549
rect 10681 24515 10715 24549
rect 10750 24515 10784 24549
rect 10819 24515 10853 24549
rect 10888 24515 10922 24549
rect 10957 24515 10991 24549
rect 11026 24515 11060 24549
rect 11095 24515 11129 24549
rect 11164 24515 11198 24549
rect 9911 24447 9945 24481
rect 9981 24447 10015 24481
rect 10051 24447 10085 24481
rect 10121 24447 10155 24481
rect 10191 24447 10225 24481
rect 10261 24447 10295 24481
rect 10331 24447 10365 24481
rect 10401 24447 10435 24481
rect 10471 24447 10505 24481
rect 10541 24447 10575 24481
rect 10611 24447 10645 24481
rect 10681 24447 10715 24481
rect 10750 24447 10784 24481
rect 10819 24447 10853 24481
rect 10888 24447 10922 24481
rect 10957 24447 10991 24481
rect 11026 24447 11060 24481
rect 11095 24447 11129 24481
rect 11164 24447 11198 24481
rect 9911 24379 9945 24413
rect 9981 24379 10015 24413
rect 10051 24379 10085 24413
rect 10121 24379 10155 24413
rect 10191 24379 10225 24413
rect 10261 24379 10295 24413
rect 10331 24379 10365 24413
rect 10401 24379 10435 24413
rect 10471 24379 10505 24413
rect 10541 24379 10575 24413
rect 10611 24379 10645 24413
rect 10681 24379 10715 24413
rect 10750 24379 10784 24413
rect 10819 24379 10853 24413
rect 10888 24379 10922 24413
rect 10957 24379 10991 24413
rect 11026 24379 11060 24413
rect 11095 24379 11129 24413
rect 11164 24379 11198 24413
rect 9911 24311 9945 24345
rect 9981 24311 10015 24345
rect 10051 24311 10085 24345
rect 10121 24311 10155 24345
rect 10191 24311 10225 24345
rect 10261 24311 10295 24345
rect 10331 24311 10365 24345
rect 10401 24311 10435 24345
rect 10471 24311 10505 24345
rect 10541 24311 10575 24345
rect 10611 24311 10645 24345
rect 10681 24311 10715 24345
rect 10750 24311 10784 24345
rect 10819 24311 10853 24345
rect 10888 24311 10922 24345
rect 10957 24311 10991 24345
rect 11026 24311 11060 24345
rect 11095 24311 11129 24345
rect 11164 24311 11198 24345
rect 9911 24243 9945 24277
rect 9981 24243 10015 24277
rect 10051 24243 10085 24277
rect 10121 24243 10155 24277
rect 10191 24243 10225 24277
rect 10261 24243 10295 24277
rect 10331 24243 10365 24277
rect 10401 24243 10435 24277
rect 10471 24243 10505 24277
rect 10541 24243 10575 24277
rect 10611 24243 10645 24277
rect 10681 24243 10715 24277
rect 10750 24243 10784 24277
rect 10819 24243 10853 24277
rect 10888 24243 10922 24277
rect 10957 24243 10991 24277
rect 11026 24243 11060 24277
rect 11095 24243 11129 24277
rect 11164 24243 11198 24277
rect 9914 24142 9948 24176
rect 9984 24142 10018 24176
rect 10054 24142 10088 24176
rect 10124 24142 10158 24176
rect 10194 24142 10228 24176
rect 10264 24142 10298 24176
rect 10334 24142 10368 24176
rect 10404 24142 10438 24176
rect 10474 24142 10508 24176
rect 10544 24142 10578 24176
rect 10614 24142 10648 24176
rect 10684 24142 10718 24176
rect 10754 24142 10788 24176
rect 9914 24074 9948 24108
rect 9984 24074 10018 24108
rect 10054 24074 10088 24108
rect 10124 24074 10158 24108
rect 10194 24074 10228 24108
rect 10264 24074 10298 24108
rect 10334 24074 10368 24108
rect 10404 24074 10438 24108
rect 10474 24074 10508 24108
rect 10544 24074 10578 24108
rect 10614 24074 10648 24108
rect 10684 24074 10718 24108
rect 10754 24074 10788 24108
rect 9914 24006 9948 24040
rect 9984 24006 10018 24040
rect 10054 24006 10088 24040
rect 10124 24006 10158 24040
rect 10194 24006 10228 24040
rect 10264 24006 10298 24040
rect 10334 24006 10368 24040
rect 10404 24006 10438 24040
rect 10474 24006 10508 24040
rect 10544 24006 10578 24040
rect 10614 24006 10648 24040
rect 10684 24006 10718 24040
rect 10754 24006 10788 24040
rect 9914 23937 9948 23971
rect 9984 23937 10018 23971
rect 10054 23937 10088 23971
rect 10124 23937 10158 23971
rect 10194 23937 10228 23971
rect 10264 23937 10298 23971
rect 10334 23937 10368 23971
rect 10404 23937 10438 23971
rect 10474 23937 10508 23971
rect 10544 23937 10578 23971
rect 10614 23937 10648 23971
rect 10684 23937 10718 23971
rect 10754 23937 10788 23971
rect 9914 23868 9948 23902
rect 9984 23868 10018 23902
rect 10054 23868 10088 23902
rect 10124 23868 10158 23902
rect 10194 23868 10228 23902
rect 10264 23868 10298 23902
rect 10334 23868 10368 23902
rect 10404 23868 10438 23902
rect 10474 23868 10508 23902
rect 10544 23868 10578 23902
rect 10614 23868 10648 23902
rect 10684 23868 10718 23902
rect 10754 23868 10788 23902
rect 9914 23799 9948 23833
rect 9984 23799 10018 23833
rect 10054 23799 10088 23833
rect 10124 23799 10158 23833
rect 10194 23799 10228 23833
rect 10264 23799 10298 23833
rect 10334 23799 10368 23833
rect 10404 23799 10438 23833
rect 10474 23799 10508 23833
rect 10544 23799 10578 23833
rect 10614 23799 10648 23833
rect 10684 23799 10718 23833
rect 10754 23799 10788 23833
rect 9914 23730 9948 23764
rect 9984 23730 10018 23764
rect 10054 23730 10088 23764
rect 10124 23730 10158 23764
rect 10194 23730 10228 23764
rect 10264 23730 10298 23764
rect 10334 23730 10368 23764
rect 10404 23730 10438 23764
rect 10474 23730 10508 23764
rect 10544 23730 10578 23764
rect 10614 23730 10648 23764
rect 10684 23730 10718 23764
rect 10754 23730 10788 23764
rect 9914 23661 9948 23695
rect 9984 23661 10018 23695
rect 10054 23661 10088 23695
rect 10124 23661 10158 23695
rect 10194 23661 10228 23695
rect 10264 23661 10298 23695
rect 10334 23661 10368 23695
rect 10404 23661 10438 23695
rect 10474 23661 10508 23695
rect 10544 23661 10578 23695
rect 10614 23661 10648 23695
rect 10684 23661 10718 23695
rect 10754 23661 10788 23695
rect 9914 23592 9948 23626
rect 9984 23592 10018 23626
rect 10054 23592 10088 23626
rect 10124 23592 10158 23626
rect 10194 23592 10228 23626
rect 10264 23592 10298 23626
rect 10334 23592 10368 23626
rect 10404 23592 10438 23626
rect 10474 23592 10508 23626
rect 10544 23592 10578 23626
rect 10614 23592 10648 23626
rect 10684 23592 10718 23626
rect 10754 23592 10788 23626
rect 9914 23523 9948 23557
rect 9984 23523 10018 23557
rect 10054 23523 10088 23557
rect 10124 23523 10158 23557
rect 10194 23523 10228 23557
rect 10264 23523 10298 23557
rect 10334 23523 10368 23557
rect 10404 23523 10438 23557
rect 10474 23523 10508 23557
rect 10544 23523 10578 23557
rect 10614 23523 10648 23557
rect 10684 23523 10718 23557
rect 10754 23523 10788 23557
rect 9914 23454 9948 23488
rect 9984 23454 10018 23488
rect 10054 23454 10088 23488
rect 10124 23454 10158 23488
rect 10194 23454 10228 23488
rect 10264 23454 10298 23488
rect 10334 23454 10368 23488
rect 10404 23454 10438 23488
rect 10474 23454 10508 23488
rect 10544 23454 10578 23488
rect 10614 23454 10648 23488
rect 10684 23454 10718 23488
rect 10754 23454 10788 23488
rect 9914 23385 9948 23419
rect 9984 23385 10018 23419
rect 10054 23385 10088 23419
rect 10124 23385 10158 23419
rect 10194 23385 10228 23419
rect 10264 23385 10298 23419
rect 10334 23385 10368 23419
rect 10404 23385 10438 23419
rect 10474 23385 10508 23419
rect 10544 23385 10578 23419
rect 10614 23385 10648 23419
rect 10684 23385 10718 23419
rect 10754 23385 10788 23419
rect 9914 23316 9948 23350
rect 9984 23316 10018 23350
rect 10054 23316 10088 23350
rect 10124 23316 10158 23350
rect 10194 23316 10228 23350
rect 10264 23316 10298 23350
rect 10334 23316 10368 23350
rect 10404 23316 10438 23350
rect 10474 23316 10508 23350
rect 10544 23316 10578 23350
rect 10614 23316 10648 23350
rect 10684 23316 10718 23350
rect 10754 23316 10788 23350
rect 9914 23247 9948 23281
rect 9984 23247 10018 23281
rect 10054 23247 10088 23281
rect 10124 23247 10158 23281
rect 10194 23247 10228 23281
rect 10264 23247 10298 23281
rect 10334 23247 10368 23281
rect 10404 23247 10438 23281
rect 10474 23247 10508 23281
rect 10544 23247 10578 23281
rect 10614 23247 10648 23281
rect 10684 23247 10718 23281
rect 10754 23247 10788 23281
rect 9914 23178 9948 23212
rect 9984 23178 10018 23212
rect 10054 23178 10088 23212
rect 10124 23178 10158 23212
rect 10194 23178 10228 23212
rect 10264 23178 10298 23212
rect 10334 23178 10368 23212
rect 10404 23178 10438 23212
rect 10474 23178 10508 23212
rect 10544 23178 10578 23212
rect 10614 23178 10648 23212
rect 10684 23178 10718 23212
rect 10754 23178 10788 23212
rect 9914 23109 9948 23143
rect 9984 23109 10018 23143
rect 10054 23109 10088 23143
rect 10124 23109 10158 23143
rect 10194 23109 10228 23143
rect 10264 23109 10298 23143
rect 10334 23109 10368 23143
rect 10404 23109 10438 23143
rect 10474 23109 10508 23143
rect 10544 23109 10578 23143
rect 10614 23109 10648 23143
rect 10684 23109 10718 23143
rect 10754 23109 10788 23143
rect 9914 23040 9948 23074
rect 9984 23040 10018 23074
rect 10054 23040 10088 23074
rect 10124 23040 10158 23074
rect 10194 23040 10228 23074
rect 10264 23040 10298 23074
rect 10334 23040 10368 23074
rect 10404 23040 10438 23074
rect 10474 23040 10508 23074
rect 10544 23040 10578 23074
rect 10614 23040 10648 23074
rect 10684 23040 10718 23074
rect 10754 23040 10788 23074
rect 14233 24150 14403 26224
rect 14233 24081 14267 24115
rect 14301 24081 14335 24115
rect 14369 24081 14403 24115
rect 14233 24012 14267 24046
rect 14301 24012 14335 24046
rect 14369 24012 14403 24046
rect 14233 23943 14267 23977
rect 14301 23943 14335 23977
rect 14369 23943 14403 23977
rect 14233 23874 14267 23908
rect 14301 23874 14335 23908
rect 14369 23874 14403 23908
rect 14233 23805 14267 23839
rect 14301 23805 14335 23839
rect 14369 23805 14403 23839
rect 14233 23736 14267 23770
rect 14301 23736 14335 23770
rect 14369 23736 14403 23770
rect 14233 23667 14267 23701
rect 14301 23667 14335 23701
rect 14369 23667 14403 23701
rect 14233 23598 14267 23632
rect 14301 23598 14335 23632
rect 14369 23598 14403 23632
rect 14233 23529 14267 23563
rect 14301 23529 14335 23563
rect 14369 23529 14403 23563
rect 14233 23460 14267 23494
rect 14301 23460 14335 23494
rect 14369 23460 14403 23494
rect 14233 23391 14267 23425
rect 14301 23391 14335 23425
rect 14369 23391 14403 23425
rect 14233 23322 14267 23356
rect 14301 23322 14335 23356
rect 14369 23322 14403 23356
rect 14233 23253 14267 23287
rect 14301 23253 14335 23287
rect 14369 23253 14403 23287
rect 14233 23184 14267 23218
rect 14301 23184 14335 23218
rect 14369 23184 14403 23218
rect 14233 23115 14267 23149
rect 14301 23115 14335 23149
rect 14369 23115 14403 23149
rect 14233 23046 14267 23080
rect 14301 23046 14335 23080
rect 14369 23046 14403 23080
rect 9914 22971 9948 23005
rect 9984 22971 10018 23005
rect 10054 22971 10088 23005
rect 10124 22971 10158 23005
rect 10194 22971 10228 23005
rect 10264 22971 10298 23005
rect 10334 22971 10368 23005
rect 10404 22971 10438 23005
rect 10474 22971 10508 23005
rect 10544 22971 10578 23005
rect 10614 22971 10648 23005
rect 10684 22971 10718 23005
rect 10754 22971 10788 23005
rect 10859 22969 10893 23003
rect 10928 22969 10962 23003
rect 10997 22969 11031 23003
rect 11066 22969 11100 23003
rect 11135 22969 11169 23003
rect 11204 22969 11238 23003
rect 11273 22969 11307 23003
rect 11342 22969 11376 23003
rect 11411 22969 11445 23003
rect 11480 22969 11514 23003
rect 11549 22969 11583 23003
rect 11618 22969 11652 23003
rect 11687 22969 11721 23003
rect 11756 22969 11790 23003
rect 11825 22969 11859 23003
rect 11894 22969 11928 23003
rect 11963 22969 11997 23003
rect 12031 22969 12065 23003
rect 12099 22969 12133 23003
rect 12167 22969 12201 23003
rect 12235 22969 12269 23003
rect 12303 22969 12337 23003
rect 12371 22969 12405 23003
rect 12439 22969 12473 23003
rect 12507 22969 12541 23003
rect 12575 22969 12609 23003
rect 12643 22969 12677 23003
rect 12711 22969 12745 23003
rect 12779 22969 12813 23003
rect 12847 22969 12881 23003
rect 12915 22969 12949 23003
rect 12983 22969 13017 23003
rect 13051 22969 13085 23003
rect 13119 22969 13153 23003
rect 13187 22969 13221 23003
rect 13255 22969 13289 23003
rect 13323 22969 13357 23003
rect 13391 22969 13425 23003
rect 13459 22969 13493 23003
rect 13527 22969 13561 23003
rect 13595 22969 13629 23003
rect 13663 22969 13697 23003
rect 13731 22969 13765 23003
rect 13799 22969 13833 23003
rect 13867 22969 13901 23003
rect 13978 22964 14012 22998
rect 14048 22964 14082 22998
rect 14118 22964 14152 22998
rect 14233 22977 14267 23011
rect 14301 22977 14335 23011
rect 14369 22977 14403 23011
rect 9901 22901 9935 22935
rect 9971 22901 10005 22935
rect 10041 22901 10075 22935
rect 10111 22901 10145 22935
rect 10181 22901 10215 22935
rect 10251 22901 10285 22935
rect 10321 22901 10355 22935
rect 10391 22901 10425 22935
rect 10461 22901 10495 22935
rect 10530 22901 10564 22935
rect 10599 22901 10633 22935
rect 10668 22901 10702 22935
rect 10737 22901 10771 22935
rect 10806 22901 10840 22935
rect 10875 22901 10909 22935
rect 10944 22901 10978 22935
rect 11013 22901 11047 22935
rect 11082 22901 11116 22935
rect 11151 22901 11185 22935
rect 11220 22901 11254 22935
rect 11289 22901 11323 22935
rect 11358 22901 11392 22935
rect 11427 22901 11461 22935
rect 11496 22901 11530 22935
rect 11565 22901 11599 22935
rect 11634 22901 11668 22935
rect 11703 22901 11737 22935
rect 11772 22901 11806 22935
rect 11841 22901 11875 22935
rect 11910 22901 11944 22935
rect 11979 22901 12013 22935
rect 12048 22901 12082 22935
rect 12117 22901 12151 22935
rect 12186 22901 12220 22935
rect 12255 22901 12289 22935
rect 12324 22901 12358 22935
rect 12393 22901 12427 22935
rect 9901 22831 9935 22865
rect 9971 22831 10005 22865
rect 10041 22831 10075 22865
rect 10111 22831 10145 22865
rect 10181 22831 10215 22865
rect 10251 22831 10285 22865
rect 10321 22831 10355 22865
rect 10391 22831 10425 22865
rect 10461 22831 10495 22865
rect 10530 22831 10564 22865
rect 10599 22831 10633 22865
rect 10668 22831 10702 22865
rect 10737 22831 10771 22865
rect 10806 22831 10840 22865
rect 10875 22831 10909 22865
rect 10944 22831 10978 22865
rect 11013 22831 11047 22865
rect 11082 22831 11116 22865
rect 11151 22831 11185 22865
rect 11220 22831 11254 22865
rect 11289 22831 11323 22865
rect 11358 22831 11392 22865
rect 11427 22831 11461 22865
rect 11496 22831 11530 22865
rect 11565 22831 11599 22865
rect 11634 22831 11668 22865
rect 11703 22831 11737 22865
rect 11772 22831 11806 22865
rect 11841 22831 11875 22865
rect 11910 22831 11944 22865
rect 11979 22831 12013 22865
rect 12048 22831 12082 22865
rect 12117 22831 12151 22865
rect 12186 22831 12220 22865
rect 12255 22831 12289 22865
rect 12324 22831 12358 22865
rect 12393 22831 12427 22865
rect 9901 22761 9935 22795
rect 9971 22761 10005 22795
rect 10041 22761 10075 22795
rect 10111 22761 10145 22795
rect 10181 22761 10215 22795
rect 10251 22761 10285 22795
rect 10321 22761 10355 22795
rect 10391 22761 10425 22795
rect 10461 22761 10495 22795
rect 10530 22761 10564 22795
rect 10599 22761 10633 22795
rect 10668 22761 10702 22795
rect 10737 22761 10771 22795
rect 10806 22761 10840 22795
rect 10875 22761 10909 22795
rect 10944 22761 10978 22795
rect 11013 22761 11047 22795
rect 11082 22761 11116 22795
rect 11151 22761 11185 22795
rect 11220 22761 11254 22795
rect 11289 22761 11323 22795
rect 11358 22761 11392 22795
rect 11427 22761 11461 22795
rect 11496 22761 11530 22795
rect 11565 22761 11599 22795
rect 11634 22761 11668 22795
rect 11703 22761 11737 22795
rect 11772 22761 11806 22795
rect 11841 22761 11875 22795
rect 11910 22761 11944 22795
rect 11979 22761 12013 22795
rect 12048 22761 12082 22795
rect 12117 22761 12151 22795
rect 12186 22761 12220 22795
rect 12255 22761 12289 22795
rect 12324 22761 12358 22795
rect 12393 22761 12427 22795
rect 9901 22691 9935 22725
rect 9971 22691 10005 22725
rect 10041 22691 10075 22725
rect 10111 22691 10145 22725
rect 10181 22691 10215 22725
rect 10251 22691 10285 22725
rect 10321 22691 10355 22725
rect 10391 22691 10425 22725
rect 10461 22691 10495 22725
rect 10530 22691 10564 22725
rect 10599 22691 10633 22725
rect 10668 22691 10702 22725
rect 10737 22691 10771 22725
rect 10806 22691 10840 22725
rect 10875 22691 10909 22725
rect 10944 22691 10978 22725
rect 11013 22691 11047 22725
rect 11082 22691 11116 22725
rect 11151 22691 11185 22725
rect 11220 22691 11254 22725
rect 11289 22691 11323 22725
rect 11358 22691 11392 22725
rect 11427 22691 11461 22725
rect 11496 22691 11530 22725
rect 11565 22691 11599 22725
rect 11634 22691 11668 22725
rect 11703 22691 11737 22725
rect 11772 22691 11806 22725
rect 11841 22691 11875 22725
rect 11910 22691 11944 22725
rect 11979 22691 12013 22725
rect 12048 22691 12082 22725
rect 12117 22691 12151 22725
rect 12186 22691 12220 22725
rect 12255 22691 12289 22725
rect 12324 22691 12358 22725
rect 12393 22691 12427 22725
rect 9901 22621 9935 22655
rect 9971 22621 10005 22655
rect 10041 22621 10075 22655
rect 10111 22621 10145 22655
rect 10181 22621 10215 22655
rect 10251 22621 10285 22655
rect 10321 22621 10355 22655
rect 10391 22621 10425 22655
rect 10461 22621 10495 22655
rect 10530 22621 10564 22655
rect 10599 22621 10633 22655
rect 10668 22621 10702 22655
rect 10737 22621 10771 22655
rect 10806 22621 10840 22655
rect 10875 22621 10909 22655
rect 10944 22621 10978 22655
rect 11013 22621 11047 22655
rect 11082 22621 11116 22655
rect 11151 22621 11185 22655
rect 11220 22621 11254 22655
rect 11289 22621 11323 22655
rect 11358 22621 11392 22655
rect 11427 22621 11461 22655
rect 11496 22621 11530 22655
rect 11565 22621 11599 22655
rect 11634 22621 11668 22655
rect 11703 22621 11737 22655
rect 11772 22621 11806 22655
rect 11841 22621 11875 22655
rect 11910 22621 11944 22655
rect 11979 22621 12013 22655
rect 12048 22621 12082 22655
rect 12117 22621 12151 22655
rect 12186 22621 12220 22655
rect 12255 22621 12289 22655
rect 12324 22621 12358 22655
rect 12393 22621 12427 22655
rect 9901 22551 9935 22585
rect 9971 22551 10005 22585
rect 10041 22551 10075 22585
rect 10111 22551 10145 22585
rect 10181 22551 10215 22585
rect 10251 22551 10285 22585
rect 10321 22551 10355 22585
rect 10391 22551 10425 22585
rect 10461 22551 10495 22585
rect 10530 22551 10564 22585
rect 10599 22551 10633 22585
rect 10668 22551 10702 22585
rect 10737 22551 10771 22585
rect 10806 22551 10840 22585
rect 10875 22551 10909 22585
rect 10944 22551 10978 22585
rect 11013 22551 11047 22585
rect 11082 22551 11116 22585
rect 11151 22551 11185 22585
rect 11220 22551 11254 22585
rect 11289 22551 11323 22585
rect 11358 22551 11392 22585
rect 11427 22551 11461 22585
rect 11496 22551 11530 22585
rect 11565 22551 11599 22585
rect 11634 22551 11668 22585
rect 11703 22551 11737 22585
rect 11772 22551 11806 22585
rect 11841 22551 11875 22585
rect 11910 22551 11944 22585
rect 11979 22551 12013 22585
rect 12048 22551 12082 22585
rect 12117 22551 12151 22585
rect 12186 22551 12220 22585
rect 12255 22551 12289 22585
rect 12324 22551 12358 22585
rect 12393 22551 12427 22585
rect 14233 22908 14267 22942
rect 14301 22908 14335 22942
rect 14369 22908 14403 22942
rect 13796 22869 13830 22903
rect 13864 22869 13898 22903
rect 13932 22869 13966 22903
rect 14000 22869 14034 22903
rect 14068 22869 14102 22903
rect 14233 22839 14267 22873
rect 14301 22839 14335 22873
rect 14369 22839 14403 22873
rect 13796 22799 13830 22833
rect 13864 22799 13898 22833
rect 13932 22799 13966 22833
rect 14000 22799 14034 22833
rect 14068 22799 14102 22833
rect 14233 22770 14267 22804
rect 14301 22770 14335 22804
rect 14369 22770 14403 22804
rect 13796 22729 13830 22763
rect 13864 22729 13898 22763
rect 13932 22729 13966 22763
rect 14000 22729 14034 22763
rect 14068 22729 14102 22763
rect 14233 22701 14267 22735
rect 14301 22701 14335 22735
rect 14369 22701 14403 22735
rect 13796 22659 13830 22693
rect 13864 22659 13898 22693
rect 13932 22659 13966 22693
rect 14000 22659 14034 22693
rect 14068 22659 14102 22693
rect 14233 22632 14267 22666
rect 14301 22632 14335 22666
rect 14369 22632 14403 22666
rect 13796 22589 13830 22623
rect 13864 22589 13898 22623
rect 13932 22589 13966 22623
rect 14000 22589 14034 22623
rect 14068 22589 14102 22623
rect 14233 22563 14267 22597
rect 14301 22563 14335 22597
rect 14369 22563 14403 22597
rect 13796 22519 13830 22553
rect 13864 22519 13898 22553
rect 13932 22519 13966 22553
rect 14000 22519 14034 22553
rect 14068 22519 14102 22553
rect 14233 22494 14267 22528
rect 14301 22494 14335 22528
rect 14369 22494 14403 22528
rect 13796 22449 13830 22483
rect 13864 22449 13898 22483
rect 13932 22449 13966 22483
rect 14000 22449 14034 22483
rect 14068 22449 14102 22483
rect 14233 22425 14267 22459
rect 14301 22425 14335 22459
rect 14369 22425 14403 22459
rect 13796 22379 13830 22413
rect 13864 22379 13898 22413
rect 13932 22379 13966 22413
rect 14000 22379 14034 22413
rect 14068 22379 14102 22413
rect 14233 22356 14267 22390
rect 14301 22356 14335 22390
rect 14369 22356 14403 22390
rect 13796 22309 13830 22343
rect 13864 22309 13898 22343
rect 13932 22309 13966 22343
rect 14000 22309 14034 22343
rect 14068 22309 14102 22343
rect 14233 22287 14267 22321
rect 14301 22287 14335 22321
rect 14369 22287 14403 22321
rect 13796 22239 13830 22273
rect 13864 22239 13898 22273
rect 13932 22239 13966 22273
rect 14000 22239 14034 22273
rect 14068 22239 14102 22273
rect 14233 22218 14267 22252
rect 14301 22218 14335 22252
rect 14369 22218 14403 22252
rect 13796 22169 13830 22203
rect 13864 22169 13898 22203
rect 13932 22169 13966 22203
rect 14000 22169 14034 22203
rect 14068 22169 14102 22203
rect 14233 22149 14267 22183
rect 14301 22149 14335 22183
rect 14369 22149 14403 22183
rect 13796 22099 13830 22133
rect 13864 22099 13898 22133
rect 13932 22099 13966 22133
rect 14000 22099 14034 22133
rect 14068 22099 14102 22133
rect 14233 22080 14267 22114
rect 14301 22080 14335 22114
rect 14369 22080 14403 22114
rect 13796 22029 13830 22063
rect 13864 22029 13898 22063
rect 13932 22029 13966 22063
rect 14000 22029 14034 22063
rect 14068 22029 14102 22063
rect 14233 22011 14267 22045
rect 14301 22011 14335 22045
rect 14369 22011 14403 22045
rect 13796 21959 13830 21993
rect 13864 21959 13898 21993
rect 13932 21959 13966 21993
rect 14000 21959 14034 21993
rect 14068 21959 14102 21993
rect 14233 21942 14267 21976
rect 14301 21942 14335 21976
rect 14369 21942 14403 21976
rect 13796 21889 13830 21923
rect 13864 21889 13898 21923
rect 13932 21889 13966 21923
rect 14000 21889 14034 21923
rect 14068 21889 14102 21923
rect 14233 21873 14267 21907
rect 14301 21873 14335 21907
rect 14369 21873 14403 21907
rect 13796 21819 13830 21853
rect 13864 21819 13898 21853
rect 13932 21819 13966 21853
rect 14000 21819 14034 21853
rect 14068 21819 14102 21853
rect 14233 21804 14267 21838
rect 14301 21804 14335 21838
rect 14369 21804 14403 21838
rect 13796 21749 13830 21783
rect 13864 21749 13898 21783
rect 13932 21749 13966 21783
rect 14000 21749 14034 21783
rect 14068 21749 14102 21783
rect 14233 21735 14267 21769
rect 14301 21735 14335 21769
rect 14369 21735 14403 21769
rect 13796 21679 13830 21713
rect 13864 21679 13898 21713
rect 13932 21679 13966 21713
rect 14000 21679 14034 21713
rect 14068 21679 14102 21713
rect 14233 21666 14267 21700
rect 14301 21666 14335 21700
rect 14369 21666 14403 21700
rect 13796 21609 13830 21643
rect 13864 21609 13898 21643
rect 13932 21609 13966 21643
rect 14000 21609 14034 21643
rect 14068 21609 14102 21643
rect 14233 21597 14267 21631
rect 14301 21597 14335 21631
rect 14369 21597 14403 21631
rect 13796 21539 13830 21573
rect 13864 21539 13898 21573
rect 13932 21539 13966 21573
rect 14000 21539 14034 21573
rect 14068 21539 14102 21573
rect 14233 21528 14267 21562
rect 14301 21528 14335 21562
rect 14369 21528 14403 21562
rect 13796 21469 13830 21503
rect 13864 21469 13898 21503
rect 13932 21469 13966 21503
rect 14000 21469 14034 21503
rect 14068 21469 14102 21503
rect 14233 21459 14267 21493
rect 14301 21459 14335 21493
rect 14369 21459 14403 21493
rect 13796 21399 13830 21433
rect 13864 21399 13898 21433
rect 13932 21399 13966 21433
rect 14000 21399 14034 21433
rect 14068 21399 14102 21433
rect 14233 21390 14267 21424
rect 14301 21390 14335 21424
rect 14369 21390 14403 21424
rect 13796 21329 13830 21363
rect 13864 21329 13898 21363
rect 13932 21329 13966 21363
rect 14000 21329 14034 21363
rect 14068 21329 14102 21363
rect 14233 21321 14267 21355
rect 14301 21321 14335 21355
rect 14369 21321 14403 21355
rect 13796 21259 13830 21293
rect 13864 21259 13898 21293
rect 13932 21259 13966 21293
rect 14000 21259 14034 21293
rect 14068 21259 14102 21293
rect 14233 21252 14267 21286
rect 14301 21252 14335 21286
rect 14369 21252 14403 21286
rect 13796 21189 13830 21223
rect 13864 21189 13898 21223
rect 13932 21189 13966 21223
rect 14000 21189 14034 21223
rect 14068 21189 14102 21223
rect 14233 21183 14267 21217
rect 14301 21183 14335 21217
rect 14369 21183 14403 21217
rect 13796 21119 13830 21153
rect 13864 21119 13898 21153
rect 13932 21119 13966 21153
rect 14000 21119 14034 21153
rect 14068 21119 14102 21153
rect 14233 21114 14267 21148
rect 14301 21114 14335 21148
rect 14369 21114 14403 21148
rect 13796 21049 13830 21083
rect 13864 21049 13898 21083
rect 13932 21049 13966 21083
rect 14000 21049 14034 21083
rect 14068 21049 14102 21083
rect 14233 21045 14267 21079
rect 14301 21045 14335 21079
rect 14369 21045 14403 21079
rect 13796 20978 13830 21012
rect 13864 20978 13898 21012
rect 13932 20978 13966 21012
rect 14000 20978 14034 21012
rect 14068 20978 14102 21012
rect 14233 20976 14267 21010
rect 14301 20976 14335 21010
rect 14369 20976 14403 21010
rect 13796 20907 13830 20941
rect 13864 20907 13898 20941
rect 13932 20907 13966 20941
rect 14000 20907 14034 20941
rect 14068 20907 14102 20941
rect 14233 20907 14267 20941
rect 14301 20907 14335 20941
rect 14369 20907 14403 20941
<< mvnsubdiffcont >>
rect 13078 30961 14200 30995
rect 13078 30927 14199 30961
rect 13077 30893 14199 30927
rect 13077 30825 14131 30893
rect 14233 30889 14267 30923
rect 14165 30788 14267 30856
rect 9759 26504 14009 26572
rect 14097 26538 14267 30788
rect 9759 26402 14077 26504
rect 14165 26470 14267 26538
rect 14233 26469 14267 26470
rect 14111 26402 14145 26436
<< locali >>
rect 9877 36379 14429 36383
rect 9877 36351 10927 36379
rect 9877 36349 9915 36351
rect 9949 36349 9987 36351
rect 10021 36349 10059 36351
rect 10093 36349 10131 36351
rect 10165 36349 10203 36351
rect 10237 36349 10275 36351
rect 10309 36349 10347 36351
rect 10381 36349 10419 36351
rect 10453 36349 10491 36351
rect 10525 36349 10563 36351
rect 10597 36349 10635 36351
rect 10669 36349 10707 36351
rect 10741 36349 10779 36351
rect 10813 36349 10851 36351
rect 9877 35975 9898 36349
rect 10885 36345 10927 36351
rect 10961 36348 11000 36379
rect 11034 36348 11073 36379
rect 11107 36348 11146 36379
rect 11180 36348 11219 36379
rect 11253 36348 11292 36379
rect 11326 36348 11365 36379
rect 11399 36348 11438 36379
rect 11472 36348 11511 36379
rect 11545 36348 11584 36379
rect 11618 36348 11657 36379
rect 11691 36348 11730 36379
rect 11764 36348 11803 36379
rect 11837 36348 11876 36379
rect 11910 36348 11949 36379
rect 11983 36348 12022 36379
rect 12056 36348 12095 36379
rect 12129 36348 12168 36379
rect 12202 36348 12241 36379
rect 12275 36348 12314 36379
rect 12348 36348 12387 36379
rect 12421 36348 12460 36379
rect 12494 36348 12533 36379
rect 12567 36348 12606 36379
rect 12640 36348 12679 36379
rect 12713 36348 12752 36379
rect 12786 36348 12825 36379
rect 12859 36348 12898 36379
rect 12932 36348 12971 36379
rect 13005 36348 13044 36379
rect 13078 36348 13117 36379
rect 13151 36348 13190 36379
rect 13224 36348 13263 36379
rect 13297 36348 13336 36379
rect 13370 36348 13409 36379
rect 13443 36348 13482 36379
rect 13516 36348 13555 36379
rect 13589 36348 13628 36379
rect 13662 36348 13701 36379
rect 13735 36348 13774 36379
rect 13808 36348 13846 36379
rect 13880 36348 13918 36379
rect 13952 36348 13990 36379
rect 14024 36348 14062 36379
rect 14096 36348 14134 36379
rect 14168 36348 14206 36379
rect 14240 36348 14278 36379
rect 14312 36348 14350 36379
rect 14384 36348 14429 36379
rect 10973 36345 11000 36348
rect 11042 36345 11073 36348
rect 10885 36317 10939 36345
rect 10884 36314 10939 36317
rect 10973 36314 11008 36345
rect 11042 36314 11077 36345
rect 11111 36314 11146 36348
rect 11180 36314 11215 36348
rect 11253 36345 11284 36348
rect 11326 36345 11353 36348
rect 11399 36345 11422 36348
rect 11472 36345 11491 36348
rect 11545 36345 11560 36348
rect 11618 36345 11629 36348
rect 11691 36345 11698 36348
rect 11764 36345 11767 36348
rect 11249 36314 11284 36345
rect 11318 36314 11353 36345
rect 11387 36314 11422 36345
rect 11456 36314 11491 36345
rect 11525 36314 11560 36345
rect 11594 36314 11629 36345
rect 11663 36314 11698 36345
rect 11732 36314 11767 36345
rect 11801 36345 11803 36348
rect 11870 36345 11876 36348
rect 11939 36345 11949 36348
rect 12008 36345 12022 36348
rect 12077 36345 12095 36348
rect 12146 36345 12168 36348
rect 12215 36345 12241 36348
rect 12284 36345 12314 36348
rect 12353 36345 12387 36348
rect 11801 36314 11836 36345
rect 11870 36314 11905 36345
rect 11939 36314 11974 36345
rect 12008 36314 12043 36345
rect 12077 36314 12112 36345
rect 12146 36314 12181 36345
rect 12215 36314 12250 36345
rect 12284 36314 12319 36345
rect 12353 36314 12388 36345
rect 12422 36314 12457 36348
rect 10884 36303 12457 36314
rect 10884 36273 10927 36303
rect 10961 36280 11000 36303
rect 11034 36280 11073 36303
rect 11107 36280 11146 36303
rect 11180 36280 11219 36303
rect 11253 36280 11292 36303
rect 11326 36280 11365 36303
rect 11399 36280 11438 36303
rect 11472 36280 11511 36303
rect 11545 36280 11584 36303
rect 11618 36280 11657 36303
rect 11691 36280 11730 36303
rect 11764 36280 11803 36303
rect 11837 36280 11876 36303
rect 11910 36280 11949 36303
rect 11983 36280 12022 36303
rect 12056 36280 12095 36303
rect 12129 36280 12168 36303
rect 12202 36280 12241 36303
rect 12275 36280 12314 36303
rect 12348 36280 12387 36303
rect 12421 36280 12457 36303
rect 10885 36269 10927 36273
rect 10973 36269 11000 36280
rect 11042 36269 11073 36280
rect 10885 36246 10939 36269
rect 10973 36246 11008 36269
rect 11042 36246 11077 36269
rect 11111 36246 11146 36280
rect 11180 36246 11215 36280
rect 11253 36269 11284 36280
rect 11326 36269 11353 36280
rect 11399 36269 11422 36280
rect 11472 36269 11491 36280
rect 11545 36269 11560 36280
rect 11618 36269 11629 36280
rect 11691 36269 11698 36280
rect 11764 36269 11767 36280
rect 11249 36246 11284 36269
rect 11318 36246 11353 36269
rect 11387 36246 11422 36269
rect 11456 36246 11491 36269
rect 11525 36246 11560 36269
rect 11594 36246 11629 36269
rect 11663 36246 11698 36269
rect 11732 36246 11767 36269
rect 11801 36269 11803 36280
rect 11870 36269 11876 36280
rect 11939 36269 11949 36280
rect 12008 36269 12022 36280
rect 12077 36269 12095 36280
rect 12146 36269 12168 36280
rect 12215 36269 12241 36280
rect 12284 36269 12314 36280
rect 12353 36269 12387 36280
rect 11801 36246 11836 36269
rect 11870 36246 11905 36269
rect 11939 36246 11974 36269
rect 12008 36246 12043 36269
rect 12077 36246 12112 36269
rect 12146 36246 12181 36269
rect 12215 36246 12250 36269
rect 12284 36246 12319 36269
rect 12353 36246 12388 36269
rect 12422 36246 12457 36280
rect 10885 36239 12457 36246
rect 10884 36227 12457 36239
rect 10884 36195 10927 36227
rect 10961 36212 11000 36227
rect 11034 36212 11073 36227
rect 11107 36212 11146 36227
rect 11180 36212 11219 36227
rect 11253 36212 11292 36227
rect 11326 36212 11365 36227
rect 11399 36212 11438 36227
rect 11472 36212 11511 36227
rect 11545 36212 11584 36227
rect 11618 36212 11657 36227
rect 11691 36212 11730 36227
rect 11764 36212 11803 36227
rect 11837 36212 11876 36227
rect 11910 36212 11949 36227
rect 11983 36212 12022 36227
rect 12056 36212 12095 36227
rect 12129 36212 12168 36227
rect 12202 36212 12241 36227
rect 12275 36212 12314 36227
rect 12348 36212 12387 36227
rect 12421 36212 12457 36227
rect 10885 36193 10927 36195
rect 10973 36193 11000 36212
rect 11042 36193 11073 36212
rect 10885 36178 10939 36193
rect 10973 36178 11008 36193
rect 11042 36178 11077 36193
rect 11111 36178 11146 36212
rect 11180 36178 11215 36212
rect 11253 36193 11284 36212
rect 11326 36193 11353 36212
rect 11399 36193 11422 36212
rect 11472 36193 11491 36212
rect 11545 36193 11560 36212
rect 11618 36193 11629 36212
rect 11691 36193 11698 36212
rect 11764 36193 11767 36212
rect 11249 36178 11284 36193
rect 11318 36178 11353 36193
rect 11387 36178 11422 36193
rect 11456 36178 11491 36193
rect 11525 36178 11560 36193
rect 11594 36178 11629 36193
rect 11663 36178 11698 36193
rect 11732 36178 11767 36193
rect 11801 36193 11803 36212
rect 11870 36193 11876 36212
rect 11939 36193 11949 36212
rect 12008 36193 12022 36212
rect 12077 36193 12095 36212
rect 12146 36193 12168 36212
rect 12215 36193 12241 36212
rect 12284 36193 12314 36212
rect 12353 36193 12387 36212
rect 11801 36178 11836 36193
rect 11870 36178 11905 36193
rect 11939 36178 11974 36193
rect 12008 36178 12043 36193
rect 12077 36178 12112 36193
rect 12146 36178 12181 36193
rect 12215 36178 12250 36193
rect 12284 36178 12319 36193
rect 12353 36178 12388 36193
rect 12422 36178 12457 36212
rect 10885 36161 12457 36178
rect 10884 36151 12457 36161
rect 10884 36117 10927 36151
rect 10961 36144 11000 36151
rect 11034 36144 11073 36151
rect 11107 36144 11146 36151
rect 11180 36144 11219 36151
rect 11253 36144 11292 36151
rect 11326 36144 11365 36151
rect 11399 36144 11438 36151
rect 11472 36144 11511 36151
rect 11545 36144 11584 36151
rect 11618 36144 11657 36151
rect 11691 36144 11730 36151
rect 11764 36144 11803 36151
rect 11837 36144 11876 36151
rect 11910 36144 11949 36151
rect 11983 36144 12022 36151
rect 12056 36144 12095 36151
rect 12129 36144 12168 36151
rect 12202 36144 12241 36151
rect 12275 36144 12314 36151
rect 12348 36144 12387 36151
rect 12421 36144 12457 36151
rect 10973 36117 11000 36144
rect 11042 36117 11073 36144
rect 10884 36116 10939 36117
rect 10885 36110 10939 36116
rect 10973 36110 11008 36117
rect 11042 36110 11077 36117
rect 11111 36110 11146 36144
rect 11180 36110 11215 36144
rect 11253 36117 11284 36144
rect 11326 36117 11353 36144
rect 11399 36117 11422 36144
rect 11472 36117 11491 36144
rect 11545 36117 11560 36144
rect 11618 36117 11629 36144
rect 11691 36117 11698 36144
rect 11764 36117 11767 36144
rect 11249 36110 11284 36117
rect 11318 36110 11353 36117
rect 11387 36110 11422 36117
rect 11456 36110 11491 36117
rect 11525 36110 11560 36117
rect 11594 36110 11629 36117
rect 11663 36110 11698 36117
rect 11732 36110 11767 36117
rect 11801 36117 11803 36144
rect 11870 36117 11876 36144
rect 11939 36117 11949 36144
rect 12008 36117 12022 36144
rect 12077 36117 12095 36144
rect 12146 36117 12168 36144
rect 12215 36117 12241 36144
rect 12284 36117 12314 36144
rect 12353 36117 12387 36144
rect 11801 36110 11836 36117
rect 11870 36110 11905 36117
rect 11939 36110 11974 36117
rect 12008 36110 12043 36117
rect 12077 36110 12112 36117
rect 12146 36110 12181 36117
rect 12215 36110 12250 36117
rect 12284 36110 12319 36117
rect 12353 36110 12388 36117
rect 12422 36110 12457 36144
rect 10885 36082 12457 36110
rect 10884 36076 12457 36082
rect 10884 36075 10939 36076
rect 10973 36075 11008 36076
rect 11042 36075 11077 36076
rect 10884 36041 10927 36075
rect 10973 36042 11000 36075
rect 11042 36042 11073 36075
rect 11111 36042 11146 36076
rect 11180 36042 11215 36076
rect 11249 36075 11284 36076
rect 11318 36075 11353 36076
rect 11387 36075 11422 36076
rect 11456 36075 11491 36076
rect 11525 36075 11560 36076
rect 11594 36075 11629 36076
rect 11663 36075 11698 36076
rect 11732 36075 11767 36076
rect 11253 36042 11284 36075
rect 11326 36042 11353 36075
rect 11399 36042 11422 36075
rect 11472 36042 11491 36075
rect 11545 36042 11560 36075
rect 11618 36042 11629 36075
rect 11691 36042 11698 36075
rect 11764 36042 11767 36075
rect 11801 36075 11836 36076
rect 11870 36075 11905 36076
rect 11939 36075 11974 36076
rect 12008 36075 12043 36076
rect 12077 36075 12112 36076
rect 12146 36075 12181 36076
rect 12215 36075 12250 36076
rect 12284 36075 12319 36076
rect 12353 36075 12388 36076
rect 11801 36042 11803 36075
rect 11870 36042 11876 36075
rect 11939 36042 11949 36075
rect 12008 36042 12022 36075
rect 12077 36042 12095 36075
rect 12146 36042 12168 36075
rect 12215 36042 12241 36075
rect 12284 36042 12314 36075
rect 12353 36042 12387 36075
rect 12422 36042 12457 36076
rect 10961 36041 11000 36042
rect 11034 36041 11073 36042
rect 11107 36041 11146 36042
rect 11180 36041 11219 36042
rect 11253 36041 11292 36042
rect 11326 36041 11365 36042
rect 11399 36041 11438 36042
rect 11472 36041 11511 36042
rect 11545 36041 11584 36042
rect 11618 36041 11657 36042
rect 11691 36041 11730 36042
rect 11764 36041 11803 36042
rect 11837 36041 11876 36042
rect 11910 36041 11949 36042
rect 11983 36041 12022 36042
rect 12056 36041 12095 36042
rect 12129 36041 12168 36042
rect 12202 36041 12241 36042
rect 12275 36041 12314 36042
rect 12348 36041 12387 36042
rect 12421 36041 12457 36042
rect 10884 36037 12457 36041
rect 10885 36008 12457 36037
rect 10885 36003 10939 36008
rect 10884 35999 10939 36003
rect 10973 35999 11008 36008
rect 11042 35999 11077 36008
rect 10884 35975 10927 35999
rect 9877 35965 10927 35975
rect 10973 35974 11000 35999
rect 11042 35974 11073 35999
rect 11111 35974 11146 36008
rect 11180 35974 11215 36008
rect 11249 35999 11284 36008
rect 11318 35999 11353 36008
rect 11387 35999 11422 36008
rect 11456 35999 11491 36008
rect 11525 35999 11560 36008
rect 11594 35999 11629 36008
rect 11663 35999 11698 36008
rect 11732 35999 11767 36008
rect 11253 35974 11284 35999
rect 11326 35974 11353 35999
rect 11399 35974 11422 35999
rect 11472 35974 11491 35999
rect 11545 35974 11560 35999
rect 11618 35974 11629 35999
rect 11691 35974 11698 35999
rect 11764 35974 11767 35999
rect 11801 35999 11836 36008
rect 11870 35999 11905 36008
rect 11939 35999 11974 36008
rect 12008 35999 12043 36008
rect 12077 35999 12112 36008
rect 12146 35999 12181 36008
rect 12215 35999 12250 36008
rect 12284 35999 12319 36008
rect 12353 35999 12388 36008
rect 11801 35974 11803 35999
rect 11870 35974 11876 35999
rect 11939 35974 11949 35999
rect 12008 35974 12022 35999
rect 12077 35974 12095 35999
rect 12146 35974 12168 35999
rect 12215 35974 12241 35999
rect 12284 35974 12314 35999
rect 12353 35974 12387 35999
rect 12422 35974 12457 36008
rect 10961 35965 11000 35974
rect 11034 35965 11073 35974
rect 11107 35965 11146 35974
rect 11180 35965 11219 35974
rect 11253 35965 11292 35974
rect 11326 35965 11365 35974
rect 11399 35965 11438 35974
rect 11472 35965 11511 35974
rect 11545 35965 11584 35974
rect 11618 35965 11657 35974
rect 11691 35965 11730 35974
rect 11764 35965 11803 35974
rect 11837 35965 11876 35974
rect 11910 35965 11949 35974
rect 11983 35965 12022 35974
rect 12056 35965 12095 35974
rect 12129 35965 12168 35974
rect 12202 35965 12241 35974
rect 12275 35965 12314 35974
rect 12348 35965 12387 35974
rect 12421 35965 12457 35974
rect 9877 35958 12457 35965
rect 9877 35940 9915 35958
rect 9949 35940 9987 35958
rect 10021 35940 10059 35958
rect 10093 35940 10131 35958
rect 10165 35940 10203 35958
rect 10237 35940 10275 35958
rect 10309 35940 10347 35958
rect 10381 35940 10419 35958
rect 10453 35940 10491 35958
rect 10525 35940 10563 35958
rect 10597 35940 10635 35958
rect 10669 35940 10707 35958
rect 10741 35940 10779 35958
rect 10813 35940 10851 35958
rect 10885 35940 12457 35958
rect 9877 35906 9898 35940
rect 9949 35924 9966 35940
rect 10021 35924 10034 35940
rect 10093 35924 10102 35940
rect 10165 35924 10170 35940
rect 10237 35924 10238 35940
rect 9932 35906 9966 35924
rect 10000 35906 10034 35924
rect 10068 35906 10102 35924
rect 10136 35906 10170 35924
rect 10204 35906 10238 35924
rect 10272 35924 10275 35940
rect 10340 35924 10347 35940
rect 10408 35924 10419 35940
rect 10476 35924 10491 35940
rect 10544 35924 10563 35940
rect 10612 35924 10635 35940
rect 10680 35924 10707 35940
rect 10748 35924 10779 35940
rect 10272 35906 10306 35924
rect 10340 35906 10374 35924
rect 10408 35906 10442 35924
rect 10476 35906 10510 35924
rect 10544 35906 10578 35924
rect 10612 35906 10646 35924
rect 10680 35906 10714 35924
rect 10748 35906 10782 35924
rect 10816 35906 10850 35940
rect 10885 35924 10939 35940
rect 10884 35923 10939 35924
rect 10973 35923 11008 35940
rect 11042 35923 11077 35940
rect 10884 35906 10927 35923
rect 10973 35906 11000 35923
rect 11042 35906 11073 35923
rect 11111 35906 11146 35940
rect 11180 35906 11215 35940
rect 11249 35923 11284 35940
rect 11318 35923 11353 35940
rect 11387 35923 11422 35940
rect 11456 35923 11491 35940
rect 11525 35923 11560 35940
rect 11594 35923 11629 35940
rect 11663 35923 11698 35940
rect 11732 35923 11767 35940
rect 11253 35906 11284 35923
rect 11326 35906 11353 35923
rect 11399 35906 11422 35923
rect 11472 35906 11491 35923
rect 11545 35906 11560 35923
rect 11618 35906 11629 35923
rect 11691 35906 11698 35923
rect 11764 35906 11767 35923
rect 11801 35923 11836 35940
rect 11870 35923 11905 35940
rect 11939 35923 11974 35940
rect 12008 35923 12043 35940
rect 12077 35923 12112 35940
rect 12146 35923 12181 35940
rect 12215 35923 12250 35940
rect 12284 35923 12319 35940
rect 12353 35923 12388 35940
rect 11801 35906 11803 35923
rect 11870 35906 11876 35923
rect 11939 35906 11949 35923
rect 12008 35906 12022 35923
rect 12077 35906 12095 35923
rect 12146 35906 12168 35923
rect 12215 35906 12241 35923
rect 12284 35906 12314 35923
rect 12353 35906 12387 35923
rect 12422 35906 12457 35940
rect 9877 35889 10927 35906
rect 10961 35889 11000 35906
rect 11034 35889 11073 35906
rect 11107 35889 11146 35906
rect 11180 35889 11219 35906
rect 11253 35889 11292 35906
rect 11326 35889 11365 35906
rect 11399 35889 11438 35906
rect 11472 35889 11511 35906
rect 11545 35889 11584 35906
rect 11618 35889 11657 35906
rect 11691 35889 11730 35906
rect 11764 35889 11803 35906
rect 11837 35889 11876 35906
rect 11910 35889 11949 35906
rect 11983 35889 12022 35906
rect 12056 35889 12095 35906
rect 12129 35889 12168 35906
rect 12202 35889 12241 35906
rect 12275 35889 12314 35906
rect 12348 35889 12387 35906
rect 12421 35889 12457 35906
rect 9877 35879 12457 35889
rect 9877 35871 9915 35879
rect 9949 35871 9987 35879
rect 10021 35871 10059 35879
rect 10093 35871 10131 35879
rect 10165 35871 10203 35879
rect 10237 35871 10275 35879
rect 10309 35871 10347 35879
rect 10381 35871 10419 35879
rect 10453 35871 10491 35879
rect 10525 35871 10563 35879
rect 10597 35871 10635 35879
rect 10669 35871 10707 35879
rect 10741 35871 10779 35879
rect 10813 35871 10851 35879
rect 10885 35872 12457 35879
rect 9877 35837 9898 35871
rect 9949 35845 9966 35871
rect 10021 35845 10034 35871
rect 10093 35845 10102 35871
rect 10165 35845 10170 35871
rect 10237 35845 10238 35871
rect 9932 35837 9966 35845
rect 10000 35837 10034 35845
rect 10068 35837 10102 35845
rect 10136 35837 10170 35845
rect 10204 35837 10238 35845
rect 10272 35845 10275 35871
rect 10340 35845 10347 35871
rect 10408 35845 10419 35871
rect 10476 35845 10491 35871
rect 10544 35845 10563 35871
rect 10612 35845 10635 35871
rect 10680 35845 10707 35871
rect 10748 35845 10779 35871
rect 10272 35837 10306 35845
rect 10340 35837 10374 35845
rect 10408 35837 10442 35845
rect 10476 35837 10510 35845
rect 10544 35837 10578 35845
rect 10612 35837 10646 35845
rect 10680 35837 10714 35845
rect 10748 35837 10782 35845
rect 10816 35837 10850 35871
rect 10885 35847 10939 35872
rect 10973 35847 11008 35872
rect 11042 35847 11077 35872
rect 10885 35845 10927 35847
rect 10884 35837 10927 35845
rect 10973 35838 11000 35847
rect 11042 35838 11073 35847
rect 11111 35838 11146 35872
rect 11180 35838 11215 35872
rect 11249 35847 11284 35872
rect 11318 35847 11353 35872
rect 11387 35847 11422 35872
rect 11456 35847 11491 35872
rect 11525 35847 11560 35872
rect 11594 35847 11629 35872
rect 11663 35847 11698 35872
rect 11732 35847 11767 35872
rect 11253 35838 11284 35847
rect 11326 35838 11353 35847
rect 11399 35838 11422 35847
rect 11472 35838 11491 35847
rect 11545 35838 11560 35847
rect 11618 35838 11629 35847
rect 11691 35838 11698 35847
rect 11764 35838 11767 35847
rect 11801 35847 11836 35872
rect 11870 35847 11905 35872
rect 11939 35847 11974 35872
rect 12008 35847 12043 35872
rect 12077 35847 12112 35872
rect 12146 35847 12181 35872
rect 12215 35847 12250 35872
rect 12284 35847 12319 35872
rect 12353 35847 12388 35872
rect 11801 35838 11803 35847
rect 11870 35838 11876 35847
rect 11939 35838 11949 35847
rect 12008 35838 12022 35847
rect 12077 35838 12095 35847
rect 12146 35838 12168 35847
rect 12215 35838 12241 35847
rect 12284 35838 12314 35847
rect 12353 35838 12387 35847
rect 12422 35838 12457 35872
rect 9877 35813 10927 35837
rect 10961 35813 11000 35838
rect 11034 35813 11073 35838
rect 11107 35813 11146 35838
rect 11180 35813 11219 35838
rect 11253 35813 11292 35838
rect 11326 35813 11365 35838
rect 11399 35813 11438 35838
rect 11472 35813 11511 35838
rect 11545 35813 11584 35838
rect 11618 35813 11657 35838
rect 11691 35813 11730 35838
rect 11764 35813 11803 35838
rect 11837 35813 11876 35838
rect 11910 35813 11949 35838
rect 11983 35813 12022 35838
rect 12056 35813 12095 35838
rect 12129 35813 12168 35838
rect 12202 35813 12241 35838
rect 12275 35813 12314 35838
rect 12348 35813 12387 35838
rect 12421 35813 12457 35838
rect 9877 35804 12457 35813
rect 9877 35802 10939 35804
rect 9877 35768 9898 35802
rect 9932 35800 9966 35802
rect 10000 35800 10034 35802
rect 10068 35800 10102 35802
rect 10136 35800 10170 35802
rect 10204 35800 10238 35802
rect 9949 35768 9966 35800
rect 10021 35768 10034 35800
rect 10093 35768 10102 35800
rect 10165 35768 10170 35800
rect 10237 35768 10238 35800
rect 10272 35800 10306 35802
rect 10340 35800 10374 35802
rect 10408 35800 10442 35802
rect 10476 35800 10510 35802
rect 10544 35800 10578 35802
rect 10612 35800 10646 35802
rect 10680 35800 10714 35802
rect 10748 35800 10782 35802
rect 10272 35768 10275 35800
rect 10340 35768 10347 35800
rect 10408 35768 10419 35800
rect 10476 35768 10491 35800
rect 10544 35768 10563 35800
rect 10612 35768 10635 35800
rect 10680 35768 10707 35800
rect 10748 35768 10779 35800
rect 10816 35768 10850 35802
rect 10884 35800 10939 35802
rect 10885 35771 10939 35800
rect 10973 35771 11008 35804
rect 11042 35771 11077 35804
rect 9877 35766 9915 35768
rect 9949 35766 9987 35768
rect 10021 35766 10059 35768
rect 10093 35766 10131 35768
rect 10165 35766 10203 35768
rect 10237 35766 10275 35768
rect 10309 35766 10347 35768
rect 10381 35766 10419 35768
rect 10453 35766 10491 35768
rect 10525 35766 10563 35768
rect 10597 35766 10635 35768
rect 10669 35766 10707 35768
rect 10741 35766 10779 35768
rect 10813 35766 10851 35768
rect 10885 35766 10927 35771
rect 10973 35770 11000 35771
rect 11042 35770 11073 35771
rect 11111 35770 11146 35804
rect 11180 35770 11215 35804
rect 11249 35771 11284 35804
rect 11318 35771 11353 35804
rect 11387 35771 11422 35804
rect 11456 35771 11491 35804
rect 11525 35771 11560 35804
rect 11594 35771 11629 35804
rect 11663 35771 11698 35804
rect 11732 35771 11767 35804
rect 11253 35770 11284 35771
rect 11326 35770 11353 35771
rect 11399 35770 11422 35771
rect 11472 35770 11491 35771
rect 11545 35770 11560 35771
rect 11618 35770 11629 35771
rect 11691 35770 11698 35771
rect 11764 35770 11767 35771
rect 11801 35771 11836 35804
rect 11870 35771 11905 35804
rect 11939 35771 11974 35804
rect 12008 35771 12043 35804
rect 12077 35771 12112 35804
rect 12146 35771 12181 35804
rect 12215 35771 12250 35804
rect 12284 35771 12319 35804
rect 12353 35771 12388 35804
rect 11801 35770 11803 35771
rect 11870 35770 11876 35771
rect 11939 35770 11949 35771
rect 12008 35770 12022 35771
rect 12077 35770 12095 35771
rect 12146 35770 12168 35771
rect 12215 35770 12241 35771
rect 12284 35770 12314 35771
rect 12353 35770 12387 35771
rect 12422 35770 12457 35804
rect 14395 35770 14429 36348
rect 9877 35737 10927 35766
rect 10961 35737 11000 35770
rect 11034 35737 11073 35770
rect 11107 35737 11146 35770
rect 11180 35737 11219 35770
rect 11253 35737 11292 35770
rect 11326 35737 11365 35770
rect 11399 35737 11438 35770
rect 11472 35737 11511 35770
rect 11545 35737 11584 35770
rect 11618 35737 11657 35770
rect 11691 35737 11730 35770
rect 11764 35737 11803 35770
rect 11837 35737 11876 35770
rect 11910 35737 11949 35770
rect 11983 35737 12022 35770
rect 12056 35737 12095 35770
rect 12129 35737 12168 35770
rect 12202 35737 12241 35770
rect 12275 35737 12314 35770
rect 12348 35737 12387 35770
rect 12421 35737 12460 35770
rect 12494 35737 12533 35770
rect 12567 35737 12606 35770
rect 12640 35737 12679 35770
rect 12713 35737 12752 35770
rect 12786 35737 12825 35770
rect 12859 35737 12898 35770
rect 12932 35737 12971 35770
rect 13005 35737 13044 35770
rect 13078 35737 13117 35770
rect 13151 35737 13190 35770
rect 13224 35737 13263 35770
rect 13297 35737 13336 35770
rect 13370 35737 13409 35770
rect 13443 35737 13482 35770
rect 13516 35737 13555 35770
rect 13589 35737 13628 35770
rect 13662 35737 13701 35770
rect 13735 35737 13774 35770
rect 13808 35737 13846 35770
rect 13880 35737 13918 35770
rect 13952 35737 13990 35770
rect 14024 35737 14062 35770
rect 14096 35737 14134 35770
rect 14168 35737 14206 35770
rect 14240 35737 14278 35770
rect 14312 35737 14350 35770
rect 14384 35737 14429 35770
rect 9877 35734 14429 35737
rect 13165 35701 14429 35734
rect 13165 35599 13202 35701
rect 14392 35697 14429 35701
rect 14418 35663 14429 35697
rect 14392 35625 14429 35663
rect 13165 35591 13216 35599
rect 13250 35591 13289 35599
rect 13323 35591 13362 35599
rect 13396 35591 13435 35599
rect 13469 35591 13508 35599
rect 13542 35591 13581 35599
rect 13615 35591 13654 35599
rect 13688 35591 13727 35599
rect 13761 35591 13800 35599
rect 13834 35591 13873 35599
rect 13907 35591 13946 35599
rect 13980 35591 14019 35599
rect 14053 35591 14092 35599
rect 14126 35591 14165 35599
rect 14199 35591 14238 35599
rect 14272 35591 14311 35599
rect 14345 35591 14384 35599
rect 14418 35591 14429 35625
rect 13165 35564 14429 35591
rect 13165 35530 13202 35564
rect 13236 35553 13270 35564
rect 13304 35553 13338 35564
rect 13372 35553 13406 35564
rect 13440 35553 13474 35564
rect 13250 35530 13270 35553
rect 13323 35530 13338 35553
rect 13396 35530 13406 35553
rect 13469 35530 13474 35553
rect 13508 35553 13542 35564
rect 13165 35519 13216 35530
rect 13250 35519 13289 35530
rect 13323 35519 13362 35530
rect 13396 35519 13435 35530
rect 13469 35519 13508 35530
rect 13576 35553 13610 35564
rect 13644 35553 13678 35564
rect 13712 35553 13746 35564
rect 13780 35553 13814 35564
rect 13848 35553 13882 35564
rect 13916 35553 13950 35564
rect 13576 35530 13581 35553
rect 13644 35530 13654 35553
rect 13712 35530 13727 35553
rect 13780 35530 13800 35553
rect 13848 35530 13873 35553
rect 13916 35530 13946 35553
rect 13984 35530 14018 35564
rect 14052 35553 14086 35564
rect 14120 35553 14154 35564
rect 14188 35553 14222 35564
rect 14256 35553 14290 35564
rect 14324 35553 14358 35564
rect 14392 35553 14429 35564
rect 14053 35530 14086 35553
rect 14126 35530 14154 35553
rect 14199 35530 14222 35553
rect 14272 35530 14290 35553
rect 14345 35530 14358 35553
rect 13542 35519 13581 35530
rect 13615 35519 13654 35530
rect 13688 35519 13727 35530
rect 13761 35519 13800 35530
rect 13834 35519 13873 35530
rect 13907 35519 13946 35530
rect 13980 35519 14019 35530
rect 14053 35519 14092 35530
rect 14126 35519 14165 35530
rect 14199 35519 14238 35530
rect 14272 35519 14311 35530
rect 14345 35519 14384 35530
rect 14418 35519 14429 35553
rect 13165 35495 14429 35519
rect 13165 35461 13202 35495
rect 13236 35481 13270 35495
rect 13304 35481 13338 35495
rect 13372 35481 13406 35495
rect 13440 35481 13474 35495
rect 13250 35461 13270 35481
rect 13323 35461 13338 35481
rect 13396 35461 13406 35481
rect 13469 35461 13474 35481
rect 13508 35481 13542 35495
rect 13165 35447 13216 35461
rect 13250 35447 13289 35461
rect 13323 35447 13362 35461
rect 13396 35447 13435 35461
rect 13469 35447 13508 35461
rect 13576 35481 13610 35495
rect 13644 35481 13678 35495
rect 13712 35481 13746 35495
rect 13780 35481 13814 35495
rect 13848 35481 13882 35495
rect 13916 35481 13950 35495
rect 13576 35461 13581 35481
rect 13644 35461 13654 35481
rect 13712 35461 13727 35481
rect 13780 35461 13800 35481
rect 13848 35461 13873 35481
rect 13916 35461 13946 35481
rect 13984 35461 14018 35495
rect 14052 35481 14086 35495
rect 14120 35481 14154 35495
rect 14188 35481 14222 35495
rect 14256 35481 14290 35495
rect 14324 35481 14358 35495
rect 14392 35481 14429 35495
rect 14053 35461 14086 35481
rect 14126 35461 14154 35481
rect 14199 35461 14222 35481
rect 14272 35461 14290 35481
rect 14345 35461 14358 35481
rect 13542 35447 13581 35461
rect 13615 35447 13654 35461
rect 13688 35447 13727 35461
rect 13761 35447 13800 35461
rect 13834 35447 13873 35461
rect 13907 35447 13946 35461
rect 13980 35447 14019 35461
rect 14053 35447 14092 35461
rect 14126 35447 14165 35461
rect 14199 35447 14238 35461
rect 14272 35447 14311 35461
rect 14345 35447 14384 35461
rect 14418 35447 14429 35481
rect 13165 35426 14429 35447
rect 13165 35392 13202 35426
rect 13236 35409 13270 35426
rect 13304 35409 13338 35426
rect 13372 35409 13406 35426
rect 13440 35409 13474 35426
rect 13250 35392 13270 35409
rect 13323 35392 13338 35409
rect 13396 35392 13406 35409
rect 13469 35392 13474 35409
rect 13508 35409 13542 35426
rect 13165 35375 13216 35392
rect 13250 35375 13289 35392
rect 13323 35375 13362 35392
rect 13396 35375 13435 35392
rect 13469 35375 13508 35392
rect 13576 35409 13610 35426
rect 13644 35409 13678 35426
rect 13712 35409 13746 35426
rect 13780 35409 13814 35426
rect 13848 35409 13882 35426
rect 13916 35409 13950 35426
rect 13576 35392 13581 35409
rect 13644 35392 13654 35409
rect 13712 35392 13727 35409
rect 13780 35392 13800 35409
rect 13848 35392 13873 35409
rect 13916 35392 13946 35409
rect 13984 35392 14018 35426
rect 14052 35409 14086 35426
rect 14120 35409 14154 35426
rect 14188 35409 14222 35426
rect 14256 35409 14290 35426
rect 14324 35409 14358 35426
rect 14392 35409 14429 35426
rect 14053 35392 14086 35409
rect 14126 35392 14154 35409
rect 14199 35392 14222 35409
rect 14272 35392 14290 35409
rect 14345 35392 14358 35409
rect 13542 35375 13581 35392
rect 13615 35375 13654 35392
rect 13688 35375 13727 35392
rect 13761 35375 13800 35392
rect 13834 35375 13873 35392
rect 13907 35375 13946 35392
rect 13980 35375 14019 35392
rect 14053 35375 14092 35392
rect 14126 35375 14165 35392
rect 14199 35375 14238 35392
rect 14272 35375 14311 35392
rect 14345 35375 14384 35392
rect 14418 35375 14429 35409
rect 13165 35357 14429 35375
rect 13165 35323 13202 35357
rect 13236 35337 13270 35357
rect 13304 35337 13338 35357
rect 13372 35337 13406 35357
rect 13440 35337 13474 35357
rect 13250 35323 13270 35337
rect 13323 35323 13338 35337
rect 13396 35323 13406 35337
rect 13469 35323 13474 35337
rect 13508 35337 13542 35357
rect 13165 35303 13216 35323
rect 13250 35303 13289 35323
rect 13323 35303 13362 35323
rect 13396 35303 13435 35323
rect 13469 35303 13508 35323
rect 13576 35337 13610 35357
rect 13644 35337 13678 35357
rect 13712 35337 13746 35357
rect 13780 35337 13814 35357
rect 13848 35337 13882 35357
rect 13916 35337 13950 35357
rect 13576 35323 13581 35337
rect 13644 35323 13654 35337
rect 13712 35323 13727 35337
rect 13780 35323 13800 35337
rect 13848 35323 13873 35337
rect 13916 35323 13946 35337
rect 13984 35323 14018 35357
rect 14052 35337 14086 35357
rect 14120 35337 14154 35357
rect 14188 35337 14222 35357
rect 14256 35337 14290 35357
rect 14324 35337 14358 35357
rect 14392 35337 14429 35357
rect 14053 35323 14086 35337
rect 14126 35323 14154 35337
rect 14199 35323 14222 35337
rect 14272 35323 14290 35337
rect 14345 35323 14358 35337
rect 13542 35303 13581 35323
rect 13615 35303 13654 35323
rect 13688 35303 13727 35323
rect 13761 35303 13800 35323
rect 13834 35303 13873 35323
rect 13907 35303 13946 35323
rect 13980 35303 14019 35323
rect 14053 35303 14092 35323
rect 14126 35303 14165 35323
rect 14199 35303 14238 35323
rect 14272 35303 14311 35323
rect 14345 35303 14384 35323
rect 14418 35303 14429 35337
rect 13165 35288 14429 35303
rect 13165 35254 13202 35288
rect 13236 35265 13270 35288
rect 13304 35265 13338 35288
rect 13372 35265 13406 35288
rect 13440 35265 13474 35288
rect 13250 35254 13270 35265
rect 13323 35254 13338 35265
rect 13396 35254 13406 35265
rect 13469 35254 13474 35265
rect 13508 35265 13542 35288
rect 13165 35231 13216 35254
rect 13250 35231 13289 35254
rect 13323 35231 13362 35254
rect 13396 35231 13435 35254
rect 13469 35231 13508 35254
rect 13576 35265 13610 35288
rect 13644 35265 13678 35288
rect 13712 35265 13746 35288
rect 13780 35265 13814 35288
rect 13848 35265 13882 35288
rect 13916 35265 13950 35288
rect 13576 35254 13581 35265
rect 13644 35254 13654 35265
rect 13712 35254 13727 35265
rect 13780 35254 13800 35265
rect 13848 35254 13873 35265
rect 13916 35254 13946 35265
rect 13984 35254 14018 35288
rect 14052 35265 14086 35288
rect 14120 35265 14154 35288
rect 14188 35265 14222 35288
rect 14256 35265 14290 35288
rect 14324 35265 14358 35288
rect 14392 35265 14429 35288
rect 14053 35254 14086 35265
rect 14126 35254 14154 35265
rect 14199 35254 14222 35265
rect 14272 35254 14290 35265
rect 14345 35254 14358 35265
rect 13542 35231 13581 35254
rect 13615 35231 13654 35254
rect 13688 35231 13727 35254
rect 13761 35231 13800 35254
rect 13834 35231 13873 35254
rect 13907 35231 13946 35254
rect 13980 35231 14019 35254
rect 14053 35231 14092 35254
rect 14126 35231 14165 35254
rect 14199 35231 14238 35254
rect 14272 35231 14311 35254
rect 14345 35231 14384 35254
rect 14418 35231 14429 35265
rect 13165 35219 14429 35231
rect 13165 35185 13202 35219
rect 13236 35193 13270 35219
rect 13304 35193 13338 35219
rect 13372 35193 13406 35219
rect 13440 35193 13474 35219
rect 13250 35185 13270 35193
rect 13323 35185 13338 35193
rect 13396 35185 13406 35193
rect 13469 35185 13474 35193
rect 13508 35193 13542 35219
rect 13165 35159 13216 35185
rect 13250 35159 13289 35185
rect 13323 35159 13362 35185
rect 13396 35159 13435 35185
rect 13469 35159 13508 35185
rect 13576 35193 13610 35219
rect 13644 35193 13678 35219
rect 13712 35193 13746 35219
rect 13780 35193 13814 35219
rect 13848 35193 13882 35219
rect 13916 35193 13950 35219
rect 13576 35185 13581 35193
rect 13644 35185 13654 35193
rect 13712 35185 13727 35193
rect 13780 35185 13800 35193
rect 13848 35185 13873 35193
rect 13916 35185 13946 35193
rect 13984 35185 14018 35219
rect 14052 35193 14086 35219
rect 14120 35193 14154 35219
rect 14188 35193 14222 35219
rect 14256 35193 14290 35219
rect 14324 35193 14358 35219
rect 14392 35193 14429 35219
rect 14053 35185 14086 35193
rect 14126 35185 14154 35193
rect 14199 35185 14222 35193
rect 14272 35185 14290 35193
rect 14345 35185 14358 35193
rect 13542 35159 13581 35185
rect 13615 35159 13654 35185
rect 13688 35159 13727 35185
rect 13761 35159 13800 35185
rect 13834 35159 13873 35185
rect 13907 35159 13946 35185
rect 13980 35159 14019 35185
rect 14053 35159 14092 35185
rect 14126 35159 14165 35185
rect 14199 35159 14238 35185
rect 14272 35159 14311 35185
rect 14345 35159 14384 35185
rect 14418 35159 14429 35193
rect 13165 35150 14429 35159
rect 13165 35116 13202 35150
rect 13236 35121 13270 35150
rect 13304 35121 13338 35150
rect 13372 35121 13406 35150
rect 13440 35121 13474 35150
rect 13250 35116 13270 35121
rect 13323 35116 13338 35121
rect 13396 35116 13406 35121
rect 13469 35116 13474 35121
rect 13508 35121 13542 35150
rect 13165 35087 13216 35116
rect 13250 35087 13289 35116
rect 13323 35087 13362 35116
rect 13396 35087 13435 35116
rect 13469 35087 13508 35116
rect 13576 35121 13610 35150
rect 13644 35121 13678 35150
rect 13712 35121 13746 35150
rect 13780 35121 13814 35150
rect 13848 35121 13882 35150
rect 13916 35121 13950 35150
rect 13576 35116 13581 35121
rect 13644 35116 13654 35121
rect 13712 35116 13727 35121
rect 13780 35116 13800 35121
rect 13848 35116 13873 35121
rect 13916 35116 13946 35121
rect 13984 35116 14018 35150
rect 14052 35121 14086 35150
rect 14120 35121 14154 35150
rect 14188 35121 14222 35150
rect 14256 35121 14290 35150
rect 14324 35121 14358 35150
rect 14392 35121 14429 35150
rect 14053 35116 14086 35121
rect 14126 35116 14154 35121
rect 14199 35116 14222 35121
rect 14272 35116 14290 35121
rect 14345 35116 14358 35121
rect 13542 35087 13581 35116
rect 13615 35087 13654 35116
rect 13688 35087 13727 35116
rect 13761 35087 13800 35116
rect 13834 35087 13873 35116
rect 13907 35087 13946 35116
rect 13980 35087 14019 35116
rect 14053 35087 14092 35116
rect 14126 35087 14165 35116
rect 14199 35087 14238 35116
rect 14272 35087 14311 35116
rect 14345 35087 14384 35116
rect 14418 35087 14429 35121
rect 13165 35081 14429 35087
rect 13165 35047 13202 35081
rect 13236 35049 13270 35081
rect 13304 35049 13338 35081
rect 13372 35049 13406 35081
rect 13440 35049 13474 35081
rect 13250 35047 13270 35049
rect 13323 35047 13338 35049
rect 13396 35047 13406 35049
rect 13469 35047 13474 35049
rect 13508 35049 13542 35081
rect 13165 35015 13216 35047
rect 13250 35015 13289 35047
rect 13323 35015 13362 35047
rect 13396 35015 13435 35047
rect 13469 35015 13508 35047
rect 13576 35049 13610 35081
rect 13644 35049 13678 35081
rect 13712 35049 13746 35081
rect 13780 35049 13814 35081
rect 13848 35049 13882 35081
rect 13916 35049 13950 35081
rect 13576 35047 13581 35049
rect 13644 35047 13654 35049
rect 13712 35047 13727 35049
rect 13780 35047 13800 35049
rect 13848 35047 13873 35049
rect 13916 35047 13946 35049
rect 13984 35047 14018 35081
rect 14052 35049 14086 35081
rect 14120 35049 14154 35081
rect 14188 35049 14222 35081
rect 14256 35049 14290 35081
rect 14324 35049 14358 35081
rect 14392 35049 14429 35081
rect 14053 35047 14086 35049
rect 14126 35047 14154 35049
rect 14199 35047 14222 35049
rect 14272 35047 14290 35049
rect 14345 35047 14358 35049
rect 13542 35015 13581 35047
rect 13615 35015 13654 35047
rect 13688 35015 13727 35047
rect 13761 35015 13800 35047
rect 13834 35015 13873 35047
rect 13907 35015 13946 35047
rect 13980 35015 14019 35047
rect 14053 35015 14092 35047
rect 14126 35015 14165 35047
rect 14199 35015 14238 35047
rect 14272 35015 14311 35047
rect 14345 35015 14384 35047
rect 14418 35015 14429 35049
rect 13165 35012 14429 35015
rect 13165 34978 13202 35012
rect 13236 34978 13270 35012
rect 13304 34978 13338 35012
rect 13372 34978 13406 35012
rect 13440 34978 13474 35012
rect 13508 34978 13542 35012
rect 13576 34978 13610 35012
rect 13644 34978 13678 35012
rect 13712 34978 13746 35012
rect 13780 34978 13814 35012
rect 13848 34978 13882 35012
rect 13916 34978 13950 35012
rect 13984 34978 14018 35012
rect 14052 34978 14086 35012
rect 14120 34978 14154 35012
rect 14188 34978 14222 35012
rect 14256 34978 14290 35012
rect 14324 34978 14358 35012
rect 14392 34978 14429 35012
rect 13165 34977 14429 34978
rect 13165 34943 13216 34977
rect 13250 34943 13289 34977
rect 13323 34943 13362 34977
rect 13396 34943 13435 34977
rect 13469 34943 13508 34977
rect 13542 34943 13581 34977
rect 13615 34943 13654 34977
rect 13688 34943 13727 34977
rect 13761 34943 13800 34977
rect 13834 34943 13873 34977
rect 13907 34943 13946 34977
rect 13980 34943 14019 34977
rect 14053 34943 14092 34977
rect 14126 34943 14165 34977
rect 14199 34943 14238 34977
rect 14272 34943 14311 34977
rect 14345 34943 14384 34977
rect 14418 34943 14429 34977
rect 13165 34909 13202 34943
rect 13236 34909 13270 34943
rect 13304 34909 13338 34943
rect 13372 34909 13406 34943
rect 13440 34909 13474 34943
rect 13508 34909 13542 34943
rect 13576 34909 13610 34943
rect 13644 34909 13678 34943
rect 13712 34909 13746 34943
rect 13780 34909 13814 34943
rect 13848 34909 13882 34943
rect 13916 34909 13950 34943
rect 13984 34909 14018 34943
rect 14052 34909 14086 34943
rect 14120 34909 14154 34943
rect 14188 34909 14222 34943
rect 14256 34909 14290 34943
rect 14324 34909 14358 34943
rect 14392 34909 14429 34943
rect 13165 34905 14429 34909
rect 13165 34874 13216 34905
rect 13250 34874 13289 34905
rect 13323 34874 13362 34905
rect 13396 34874 13435 34905
rect 13469 34874 13508 34905
rect 13165 34840 13202 34874
rect 13250 34871 13270 34874
rect 13323 34871 13338 34874
rect 13396 34871 13406 34874
rect 13469 34871 13474 34874
rect 13236 34840 13270 34871
rect 13304 34840 13338 34871
rect 13372 34840 13406 34871
rect 13440 34840 13474 34871
rect 13542 34874 13581 34905
rect 13615 34874 13654 34905
rect 13688 34874 13727 34905
rect 13761 34874 13800 34905
rect 13834 34874 13873 34905
rect 13907 34874 13946 34905
rect 13980 34874 14019 34905
rect 14053 34874 14092 34905
rect 14126 34874 14165 34905
rect 14199 34874 14238 34905
rect 14272 34874 14311 34905
rect 14345 34874 14384 34905
rect 13508 34840 13542 34871
rect 13576 34871 13581 34874
rect 13644 34871 13654 34874
rect 13712 34871 13727 34874
rect 13780 34871 13800 34874
rect 13848 34871 13873 34874
rect 13916 34871 13946 34874
rect 13576 34840 13610 34871
rect 13644 34840 13678 34871
rect 13712 34840 13746 34871
rect 13780 34840 13814 34871
rect 13848 34840 13882 34871
rect 13916 34840 13950 34871
rect 13984 34840 14018 34874
rect 14053 34871 14086 34874
rect 14126 34871 14154 34874
rect 14199 34871 14222 34874
rect 14272 34871 14290 34874
rect 14345 34871 14358 34874
rect 14418 34871 14429 34905
rect 14052 34840 14086 34871
rect 14120 34840 14154 34871
rect 14188 34840 14222 34871
rect 14256 34840 14290 34871
rect 14324 34840 14358 34871
rect 14392 34840 14429 34871
rect 13165 34833 14429 34840
rect 13165 34805 13216 34833
rect 13250 34805 13289 34833
rect 13323 34805 13362 34833
rect 13396 34805 13435 34833
rect 13469 34805 13508 34833
rect 13165 34771 13202 34805
rect 13250 34799 13270 34805
rect 13323 34799 13338 34805
rect 13396 34799 13406 34805
rect 13469 34799 13474 34805
rect 13236 34771 13270 34799
rect 13304 34771 13338 34799
rect 13372 34771 13406 34799
rect 13440 34771 13474 34799
rect 13542 34805 13581 34833
rect 13615 34805 13654 34833
rect 13688 34805 13727 34833
rect 13761 34805 13800 34833
rect 13834 34805 13873 34833
rect 13907 34805 13946 34833
rect 13980 34805 14019 34833
rect 14053 34805 14092 34833
rect 14126 34805 14165 34833
rect 14199 34805 14238 34833
rect 14272 34805 14311 34833
rect 14345 34805 14384 34833
rect 13508 34771 13542 34799
rect 13576 34799 13581 34805
rect 13644 34799 13654 34805
rect 13712 34799 13727 34805
rect 13780 34799 13800 34805
rect 13848 34799 13873 34805
rect 13916 34799 13946 34805
rect 13576 34771 13610 34799
rect 13644 34771 13678 34799
rect 13712 34771 13746 34799
rect 13780 34771 13814 34799
rect 13848 34771 13882 34799
rect 13916 34771 13950 34799
rect 13984 34771 14018 34805
rect 14053 34799 14086 34805
rect 14126 34799 14154 34805
rect 14199 34799 14222 34805
rect 14272 34799 14290 34805
rect 14345 34799 14358 34805
rect 14418 34799 14429 34833
rect 14052 34771 14086 34799
rect 14120 34771 14154 34799
rect 14188 34771 14222 34799
rect 14256 34771 14290 34799
rect 14324 34771 14358 34799
rect 14392 34771 14429 34799
rect 13165 34760 14429 34771
rect 13165 34736 13216 34760
rect 13250 34736 13289 34760
rect 13323 34736 13362 34760
rect 13396 34736 13435 34760
rect 13469 34736 13508 34760
rect 13165 34702 13202 34736
rect 13250 34726 13270 34736
rect 13323 34726 13338 34736
rect 13396 34726 13406 34736
rect 13469 34726 13474 34736
rect 13236 34702 13270 34726
rect 13304 34702 13338 34726
rect 13372 34702 13406 34726
rect 13440 34702 13474 34726
rect 13542 34736 13581 34760
rect 13615 34736 13654 34760
rect 13688 34736 13727 34760
rect 13761 34736 13800 34760
rect 13834 34736 13873 34760
rect 13907 34736 13946 34760
rect 13980 34736 14019 34760
rect 14053 34736 14092 34760
rect 14126 34736 14165 34760
rect 14199 34736 14238 34760
rect 14272 34736 14311 34760
rect 14345 34736 14384 34760
rect 13508 34702 13542 34726
rect 13576 34726 13581 34736
rect 13644 34726 13654 34736
rect 13712 34726 13727 34736
rect 13780 34726 13800 34736
rect 13848 34726 13873 34736
rect 13916 34726 13946 34736
rect 13576 34702 13610 34726
rect 13644 34702 13678 34726
rect 13712 34702 13746 34726
rect 13780 34702 13814 34726
rect 13848 34702 13882 34726
rect 13916 34702 13950 34726
rect 13984 34702 14018 34736
rect 14053 34726 14086 34736
rect 14126 34726 14154 34736
rect 14199 34726 14222 34736
rect 14272 34726 14290 34736
rect 14345 34726 14358 34736
rect 14418 34726 14429 34760
rect 14052 34702 14086 34726
rect 14120 34702 14154 34726
rect 14188 34702 14222 34726
rect 14256 34702 14290 34726
rect 14324 34702 14358 34726
rect 14392 34702 14429 34726
rect 13165 34687 14429 34702
rect 13165 34667 13216 34687
rect 13250 34667 13289 34687
rect 13323 34667 13362 34687
rect 13396 34667 13435 34687
rect 13469 34667 13508 34687
rect 13165 34633 13202 34667
rect 13250 34653 13270 34667
rect 13323 34653 13338 34667
rect 13396 34653 13406 34667
rect 13469 34653 13474 34667
rect 13236 34633 13270 34653
rect 13304 34633 13338 34653
rect 13372 34633 13406 34653
rect 13440 34633 13474 34653
rect 13542 34667 13581 34687
rect 13615 34667 13654 34687
rect 13688 34667 13727 34687
rect 13761 34667 13800 34687
rect 13834 34667 13873 34687
rect 13907 34667 13946 34687
rect 13980 34667 14019 34687
rect 14053 34667 14092 34687
rect 14126 34667 14165 34687
rect 14199 34667 14238 34687
rect 14272 34667 14311 34687
rect 14345 34667 14384 34687
rect 13508 34633 13542 34653
rect 13576 34653 13581 34667
rect 13644 34653 13654 34667
rect 13712 34653 13727 34667
rect 13780 34653 13800 34667
rect 13848 34653 13873 34667
rect 13916 34653 13946 34667
rect 13576 34633 13610 34653
rect 13644 34633 13678 34653
rect 13712 34633 13746 34653
rect 13780 34633 13814 34653
rect 13848 34633 13882 34653
rect 13916 34633 13950 34653
rect 13984 34633 14018 34667
rect 14053 34653 14086 34667
rect 14126 34653 14154 34667
rect 14199 34653 14222 34667
rect 14272 34653 14290 34667
rect 14345 34653 14358 34667
rect 14418 34653 14429 34687
rect 14052 34633 14086 34653
rect 14120 34633 14154 34653
rect 14188 34633 14222 34653
rect 14256 34633 14290 34653
rect 14324 34633 14358 34653
rect 14392 34633 14429 34653
rect 13165 34614 14429 34633
rect 13165 34598 13216 34614
rect 13250 34598 13289 34614
rect 13323 34598 13362 34614
rect 13396 34598 13435 34614
rect 13469 34598 13508 34614
rect 13165 34564 13202 34598
rect 13250 34580 13270 34598
rect 13323 34580 13338 34598
rect 13396 34580 13406 34598
rect 13469 34580 13474 34598
rect 13236 34564 13270 34580
rect 13304 34564 13338 34580
rect 13372 34564 13406 34580
rect 13440 34564 13474 34580
rect 13542 34598 13581 34614
rect 13615 34598 13654 34614
rect 13688 34598 13727 34614
rect 13761 34598 13800 34614
rect 13834 34598 13873 34614
rect 13907 34598 13946 34614
rect 13980 34598 14019 34614
rect 14053 34598 14092 34614
rect 14126 34598 14165 34614
rect 14199 34598 14238 34614
rect 14272 34598 14311 34614
rect 14345 34598 14384 34614
rect 13508 34564 13542 34580
rect 13576 34580 13581 34598
rect 13644 34580 13654 34598
rect 13712 34580 13727 34598
rect 13780 34580 13800 34598
rect 13848 34580 13873 34598
rect 13916 34580 13946 34598
rect 13576 34564 13610 34580
rect 13644 34564 13678 34580
rect 13712 34564 13746 34580
rect 13780 34564 13814 34580
rect 13848 34564 13882 34580
rect 13916 34564 13950 34580
rect 13984 34564 14018 34598
rect 14053 34580 14086 34598
rect 14126 34580 14154 34598
rect 14199 34580 14222 34598
rect 14272 34580 14290 34598
rect 14345 34580 14358 34598
rect 14418 34580 14429 34614
rect 14052 34564 14086 34580
rect 14120 34564 14154 34580
rect 14188 34564 14222 34580
rect 14256 34564 14290 34580
rect 14324 34564 14358 34580
rect 14392 34564 14429 34580
rect 13165 34541 14429 34564
rect 13165 34529 13216 34541
rect 13250 34529 13289 34541
rect 13323 34529 13362 34541
rect 13396 34529 13435 34541
rect 13469 34529 13508 34541
rect 13165 34495 13202 34529
rect 13250 34507 13270 34529
rect 13323 34507 13338 34529
rect 13396 34507 13406 34529
rect 13469 34507 13474 34529
rect 13236 34495 13270 34507
rect 13304 34495 13338 34507
rect 13372 34495 13406 34507
rect 13440 34495 13474 34507
rect 13542 34529 13581 34541
rect 13615 34529 13654 34541
rect 13688 34529 13727 34541
rect 13761 34529 13800 34541
rect 13834 34529 13873 34541
rect 13907 34529 13946 34541
rect 13980 34529 14019 34541
rect 14053 34529 14092 34541
rect 14126 34529 14165 34541
rect 14199 34529 14238 34541
rect 14272 34529 14311 34541
rect 14345 34529 14384 34541
rect 13508 34495 13542 34507
rect 13576 34507 13581 34529
rect 13644 34507 13654 34529
rect 13712 34507 13727 34529
rect 13780 34507 13800 34529
rect 13848 34507 13873 34529
rect 13916 34507 13946 34529
rect 13576 34495 13610 34507
rect 13644 34495 13678 34507
rect 13712 34495 13746 34507
rect 13780 34495 13814 34507
rect 13848 34495 13882 34507
rect 13916 34495 13950 34507
rect 13984 34495 14018 34529
rect 14053 34507 14086 34529
rect 14126 34507 14154 34529
rect 14199 34507 14222 34529
rect 14272 34507 14290 34529
rect 14345 34507 14358 34529
rect 14418 34507 14429 34541
rect 14052 34495 14086 34507
rect 14120 34495 14154 34507
rect 14188 34495 14222 34507
rect 14256 34495 14290 34507
rect 14324 34495 14358 34507
rect 14392 34495 14429 34507
rect 13165 34468 14429 34495
rect 13165 34460 13216 34468
rect 13250 34460 13289 34468
rect 13323 34460 13362 34468
rect 13396 34460 13435 34468
rect 13469 34460 13508 34468
rect 13165 34426 13202 34460
rect 13250 34434 13270 34460
rect 13323 34434 13338 34460
rect 13396 34434 13406 34460
rect 13469 34434 13474 34460
rect 13236 34426 13270 34434
rect 13304 34426 13338 34434
rect 13372 34426 13406 34434
rect 13440 34426 13474 34434
rect 13542 34460 13581 34468
rect 13615 34460 13654 34468
rect 13688 34460 13727 34468
rect 13761 34460 13800 34468
rect 13834 34460 13873 34468
rect 13907 34460 13946 34468
rect 13980 34460 14019 34468
rect 14053 34460 14092 34468
rect 14126 34460 14165 34468
rect 14199 34460 14238 34468
rect 14272 34460 14311 34468
rect 14345 34460 14384 34468
rect 13508 34426 13542 34434
rect 13576 34434 13581 34460
rect 13644 34434 13654 34460
rect 13712 34434 13727 34460
rect 13780 34434 13800 34460
rect 13848 34434 13873 34460
rect 13916 34434 13946 34460
rect 13576 34426 13610 34434
rect 13644 34426 13678 34434
rect 13712 34426 13746 34434
rect 13780 34426 13814 34434
rect 13848 34426 13882 34434
rect 13916 34426 13950 34434
rect 13984 34426 14018 34460
rect 14053 34434 14086 34460
rect 14126 34434 14154 34460
rect 14199 34434 14222 34460
rect 14272 34434 14290 34460
rect 14345 34434 14358 34460
rect 14418 34434 14429 34468
rect 14052 34426 14086 34434
rect 14120 34426 14154 34434
rect 14188 34426 14222 34434
rect 14256 34426 14290 34434
rect 14324 34426 14358 34434
rect 14392 34426 14429 34434
rect 13165 34395 14429 34426
rect 13165 34391 13216 34395
rect 13250 34391 13289 34395
rect 13323 34391 13362 34395
rect 13396 34391 13435 34395
rect 13469 34391 13508 34395
rect 13165 34357 13202 34391
rect 13250 34361 13270 34391
rect 13323 34361 13338 34391
rect 13396 34361 13406 34391
rect 13469 34361 13474 34391
rect 13236 34357 13270 34361
rect 13304 34357 13338 34361
rect 13372 34357 13406 34361
rect 13440 34357 13474 34361
rect 13542 34391 13581 34395
rect 13615 34391 13654 34395
rect 13688 34391 13727 34395
rect 13761 34391 13800 34395
rect 13834 34391 13873 34395
rect 13907 34391 13946 34395
rect 13980 34391 14019 34395
rect 14053 34391 14092 34395
rect 14126 34391 14165 34395
rect 14199 34391 14238 34395
rect 14272 34391 14311 34395
rect 14345 34391 14384 34395
rect 13508 34357 13542 34361
rect 13576 34361 13581 34391
rect 13644 34361 13654 34391
rect 13712 34361 13727 34391
rect 13780 34361 13800 34391
rect 13848 34361 13873 34391
rect 13916 34361 13946 34391
rect 13576 34357 13610 34361
rect 13644 34357 13678 34361
rect 13712 34357 13746 34361
rect 13780 34357 13814 34361
rect 13848 34357 13882 34361
rect 13916 34357 13950 34361
rect 13984 34357 14018 34391
rect 14053 34361 14086 34391
rect 14126 34361 14154 34391
rect 14199 34361 14222 34391
rect 14272 34361 14290 34391
rect 14345 34361 14358 34391
rect 14418 34361 14429 34395
rect 14052 34357 14086 34361
rect 14120 34357 14154 34361
rect 14188 34357 14222 34361
rect 14256 34357 14290 34361
rect 14324 34357 14358 34361
rect 14392 34357 14429 34361
rect 13165 34322 14429 34357
rect 13165 34288 13202 34322
rect 13250 34288 13270 34322
rect 13323 34288 13338 34322
rect 13396 34288 13406 34322
rect 13469 34288 13474 34322
rect 13576 34288 13581 34322
rect 13644 34288 13654 34322
rect 13712 34288 13727 34322
rect 13780 34288 13800 34322
rect 13848 34288 13873 34322
rect 13916 34288 13946 34322
rect 13984 34288 14018 34322
rect 14053 34288 14086 34322
rect 14126 34288 14154 34322
rect 14199 34288 14222 34322
rect 14272 34288 14290 34322
rect 14345 34288 14358 34322
rect 14418 34288 14429 34322
rect 13165 34253 14429 34288
rect 13165 34219 13202 34253
rect 13236 34249 13270 34253
rect 13304 34249 13338 34253
rect 13372 34249 13406 34253
rect 13440 34249 13474 34253
rect 13250 34219 13270 34249
rect 13323 34219 13338 34249
rect 13396 34219 13406 34249
rect 13469 34219 13474 34249
rect 13508 34249 13542 34253
rect 13165 34215 13216 34219
rect 13250 34215 13289 34219
rect 13323 34215 13362 34219
rect 13396 34215 13435 34219
rect 13469 34215 13508 34219
rect 13576 34249 13610 34253
rect 13644 34249 13678 34253
rect 13712 34249 13746 34253
rect 13780 34249 13814 34253
rect 13848 34249 13882 34253
rect 13916 34249 13950 34253
rect 13576 34219 13581 34249
rect 13644 34219 13654 34249
rect 13712 34219 13727 34249
rect 13780 34219 13800 34249
rect 13848 34219 13873 34249
rect 13916 34219 13946 34249
rect 13984 34219 14018 34253
rect 14052 34249 14086 34253
rect 14120 34249 14154 34253
rect 14188 34249 14222 34253
rect 14256 34249 14290 34253
rect 14324 34249 14358 34253
rect 14392 34249 14429 34253
rect 14053 34219 14086 34249
rect 14126 34219 14154 34249
rect 14199 34219 14222 34249
rect 14272 34219 14290 34249
rect 14345 34219 14358 34249
rect 13542 34215 13581 34219
rect 13615 34215 13654 34219
rect 13688 34215 13727 34219
rect 13761 34215 13800 34219
rect 13834 34215 13873 34219
rect 13907 34215 13946 34219
rect 13980 34215 14019 34219
rect 14053 34215 14092 34219
rect 14126 34215 14165 34219
rect 14199 34215 14238 34219
rect 14272 34215 14311 34219
rect 14345 34215 14384 34219
rect 14418 34215 14429 34249
rect 13165 34184 14429 34215
rect 13165 34150 13202 34184
rect 13236 34176 13270 34184
rect 13304 34176 13338 34184
rect 13372 34176 13406 34184
rect 13440 34176 13474 34184
rect 13250 34150 13270 34176
rect 13323 34150 13338 34176
rect 13396 34150 13406 34176
rect 13469 34150 13474 34176
rect 13508 34176 13542 34184
rect 13165 34142 13216 34150
rect 13250 34142 13289 34150
rect 13323 34142 13362 34150
rect 13396 34142 13435 34150
rect 13469 34142 13508 34150
rect 13576 34176 13610 34184
rect 13644 34176 13678 34184
rect 13712 34176 13746 34184
rect 13780 34176 13814 34184
rect 13848 34176 13882 34184
rect 13916 34176 13950 34184
rect 13576 34150 13581 34176
rect 13644 34150 13654 34176
rect 13712 34150 13727 34176
rect 13780 34150 13800 34176
rect 13848 34150 13873 34176
rect 13916 34150 13946 34176
rect 13984 34150 14018 34184
rect 14052 34176 14086 34184
rect 14120 34176 14154 34184
rect 14188 34176 14222 34184
rect 14256 34176 14290 34184
rect 14324 34176 14358 34184
rect 14392 34176 14429 34184
rect 14053 34150 14086 34176
rect 14126 34150 14154 34176
rect 14199 34150 14222 34176
rect 14272 34150 14290 34176
rect 14345 34150 14358 34176
rect 13542 34142 13581 34150
rect 13615 34142 13654 34150
rect 13688 34142 13727 34150
rect 13761 34142 13800 34150
rect 13834 34142 13873 34150
rect 13907 34142 13946 34150
rect 13980 34142 14019 34150
rect 14053 34142 14092 34150
rect 14126 34142 14165 34150
rect 14199 34142 14238 34150
rect 14272 34142 14311 34150
rect 14345 34142 14384 34150
rect 14418 34142 14429 34176
rect 13165 34115 14429 34142
rect 13165 34081 13202 34115
rect 13236 34103 13270 34115
rect 13304 34103 13338 34115
rect 13372 34103 13406 34115
rect 13440 34103 13474 34115
rect 13250 34081 13270 34103
rect 13323 34081 13338 34103
rect 13396 34081 13406 34103
rect 13469 34081 13474 34103
rect 13508 34103 13542 34115
rect 13165 34069 13216 34081
rect 13250 34069 13289 34081
rect 13323 34069 13362 34081
rect 13396 34069 13435 34081
rect 13469 34069 13508 34081
rect 13576 34103 13610 34115
rect 13644 34103 13678 34115
rect 13712 34103 13746 34115
rect 13780 34103 13814 34115
rect 13848 34103 13882 34115
rect 13916 34103 13950 34115
rect 13576 34081 13581 34103
rect 13644 34081 13654 34103
rect 13712 34081 13727 34103
rect 13780 34081 13800 34103
rect 13848 34081 13873 34103
rect 13916 34081 13946 34103
rect 13984 34081 14018 34115
rect 14052 34103 14086 34115
rect 14120 34103 14154 34115
rect 14188 34103 14222 34115
rect 14256 34103 14290 34115
rect 14324 34103 14358 34115
rect 14392 34103 14429 34115
rect 14053 34081 14086 34103
rect 14126 34081 14154 34103
rect 14199 34081 14222 34103
rect 14272 34081 14290 34103
rect 14345 34081 14358 34103
rect 13542 34069 13581 34081
rect 13615 34069 13654 34081
rect 13688 34069 13727 34081
rect 13761 34069 13800 34081
rect 13834 34069 13873 34081
rect 13907 34069 13946 34081
rect 13980 34069 14019 34081
rect 14053 34069 14092 34081
rect 14126 34069 14165 34081
rect 14199 34069 14238 34081
rect 14272 34069 14311 34081
rect 14345 34069 14384 34081
rect 14418 34069 14429 34103
rect 13165 34046 14429 34069
rect 13165 34012 13202 34046
rect 13236 34030 13270 34046
rect 13304 34030 13338 34046
rect 13372 34030 13406 34046
rect 13440 34030 13474 34046
rect 13250 34012 13270 34030
rect 13323 34012 13338 34030
rect 13396 34012 13406 34030
rect 13469 34012 13474 34030
rect 13508 34030 13542 34046
rect 13165 33996 13216 34012
rect 13250 33996 13289 34012
rect 13323 33996 13362 34012
rect 13396 33996 13435 34012
rect 13469 33996 13508 34012
rect 13576 34030 13610 34046
rect 13644 34030 13678 34046
rect 13712 34030 13746 34046
rect 13780 34030 13814 34046
rect 13848 34030 13882 34046
rect 13916 34030 13950 34046
rect 13576 34012 13581 34030
rect 13644 34012 13654 34030
rect 13712 34012 13727 34030
rect 13780 34012 13800 34030
rect 13848 34012 13873 34030
rect 13916 34012 13946 34030
rect 13984 34012 14018 34046
rect 14052 34030 14086 34046
rect 14120 34030 14154 34046
rect 14188 34030 14222 34046
rect 14256 34030 14290 34046
rect 14324 34030 14358 34046
rect 14392 34030 14429 34046
rect 14053 34012 14086 34030
rect 14126 34012 14154 34030
rect 14199 34012 14222 34030
rect 14272 34012 14290 34030
rect 14345 34012 14358 34030
rect 13542 33996 13581 34012
rect 13615 33996 13654 34012
rect 13688 33996 13727 34012
rect 13761 33996 13800 34012
rect 13834 33996 13873 34012
rect 13907 33996 13946 34012
rect 13980 33996 14019 34012
rect 14053 33996 14092 34012
rect 14126 33996 14165 34012
rect 14199 33996 14238 34012
rect 14272 33996 14311 34012
rect 14345 33996 14384 34012
rect 14418 33996 14429 34030
rect 13165 33977 14429 33996
rect 13165 33943 13202 33977
rect 13236 33957 13270 33977
rect 13304 33957 13338 33977
rect 13372 33957 13406 33977
rect 13440 33957 13474 33977
rect 13250 33943 13270 33957
rect 13323 33943 13338 33957
rect 13396 33943 13406 33957
rect 13469 33943 13474 33957
rect 13508 33957 13542 33977
rect 13165 33923 13216 33943
rect 13250 33923 13289 33943
rect 13323 33923 13362 33943
rect 13396 33923 13435 33943
rect 13469 33923 13508 33943
rect 13576 33957 13610 33977
rect 13644 33957 13678 33977
rect 13712 33957 13746 33977
rect 13780 33957 13814 33977
rect 13848 33957 13882 33977
rect 13916 33957 13950 33977
rect 13576 33943 13581 33957
rect 13644 33943 13654 33957
rect 13712 33943 13727 33957
rect 13780 33943 13800 33957
rect 13848 33943 13873 33957
rect 13916 33943 13946 33957
rect 13984 33943 14018 33977
rect 14052 33957 14086 33977
rect 14120 33957 14154 33977
rect 14188 33957 14222 33977
rect 14256 33957 14290 33977
rect 14324 33957 14358 33977
rect 14392 33957 14429 33977
rect 14053 33943 14086 33957
rect 14126 33943 14154 33957
rect 14199 33943 14222 33957
rect 14272 33943 14290 33957
rect 14345 33943 14358 33957
rect 13542 33923 13581 33943
rect 13615 33923 13654 33943
rect 13688 33923 13727 33943
rect 13761 33923 13800 33943
rect 13834 33923 13873 33943
rect 13907 33923 13946 33943
rect 13980 33923 14019 33943
rect 14053 33923 14092 33943
rect 14126 33923 14165 33943
rect 14199 33923 14238 33943
rect 14272 33923 14311 33943
rect 14345 33923 14384 33943
rect 14418 33923 14429 33957
rect 13165 33908 14429 33923
rect 13165 33874 13202 33908
rect 13236 33884 13270 33908
rect 13304 33884 13338 33908
rect 13372 33884 13406 33908
rect 13440 33884 13474 33908
rect 13250 33874 13270 33884
rect 13323 33874 13338 33884
rect 13396 33874 13406 33884
rect 13469 33874 13474 33884
rect 13508 33884 13542 33908
rect 13165 33850 13216 33874
rect 13250 33850 13289 33874
rect 13323 33850 13362 33874
rect 13396 33850 13435 33874
rect 13469 33850 13508 33874
rect 13576 33884 13610 33908
rect 13644 33884 13678 33908
rect 13712 33884 13746 33908
rect 13780 33884 13814 33908
rect 13848 33884 13882 33908
rect 13916 33884 13950 33908
rect 13576 33874 13581 33884
rect 13644 33874 13654 33884
rect 13712 33874 13727 33884
rect 13780 33874 13800 33884
rect 13848 33874 13873 33884
rect 13916 33874 13946 33884
rect 13984 33874 14018 33908
rect 14052 33884 14086 33908
rect 14120 33884 14154 33908
rect 14188 33884 14222 33908
rect 14256 33884 14290 33908
rect 14324 33884 14358 33908
rect 14392 33884 14429 33908
rect 14053 33874 14086 33884
rect 14126 33874 14154 33884
rect 14199 33874 14222 33884
rect 14272 33874 14290 33884
rect 14345 33874 14358 33884
rect 13542 33850 13581 33874
rect 13615 33850 13654 33874
rect 13688 33850 13727 33874
rect 13761 33850 13800 33874
rect 13834 33850 13873 33874
rect 13907 33850 13946 33874
rect 13980 33850 14019 33874
rect 14053 33850 14092 33874
rect 14126 33850 14165 33874
rect 14199 33850 14238 33874
rect 14272 33850 14311 33874
rect 14345 33850 14384 33874
rect 14418 33850 14429 33884
rect 13165 33839 14429 33850
rect 13165 33805 13202 33839
rect 13236 33811 13270 33839
rect 13304 33811 13338 33839
rect 13372 33811 13406 33839
rect 13440 33811 13474 33839
rect 13250 33805 13270 33811
rect 13323 33805 13338 33811
rect 13396 33805 13406 33811
rect 13469 33805 13474 33811
rect 13508 33811 13542 33839
rect 13165 33777 13216 33805
rect 13250 33777 13289 33805
rect 13323 33777 13362 33805
rect 13396 33777 13435 33805
rect 13469 33777 13508 33805
rect 13576 33811 13610 33839
rect 13644 33811 13678 33839
rect 13712 33811 13746 33839
rect 13780 33811 13814 33839
rect 13848 33811 13882 33839
rect 13916 33811 13950 33839
rect 13576 33805 13581 33811
rect 13644 33805 13654 33811
rect 13712 33805 13727 33811
rect 13780 33805 13800 33811
rect 13848 33805 13873 33811
rect 13916 33805 13946 33811
rect 13984 33805 14018 33839
rect 14052 33811 14086 33839
rect 14120 33811 14154 33839
rect 14188 33811 14222 33839
rect 14256 33811 14290 33839
rect 14324 33811 14358 33839
rect 14392 33811 14429 33839
rect 14053 33805 14086 33811
rect 14126 33805 14154 33811
rect 14199 33805 14222 33811
rect 14272 33805 14290 33811
rect 14345 33805 14358 33811
rect 13542 33777 13581 33805
rect 13615 33777 13654 33805
rect 13688 33777 13727 33805
rect 13761 33777 13800 33805
rect 13834 33777 13873 33805
rect 13907 33777 13946 33805
rect 13980 33777 14019 33805
rect 14053 33777 14092 33805
rect 14126 33777 14165 33805
rect 14199 33777 14238 33805
rect 14272 33777 14311 33805
rect 14345 33777 14384 33805
rect 14418 33777 14429 33811
rect 13165 33770 14429 33777
rect 13165 33736 13202 33770
rect 13236 33738 13270 33770
rect 13304 33738 13338 33770
rect 13372 33738 13406 33770
rect 13440 33738 13474 33770
rect 13250 33736 13270 33738
rect 13323 33736 13338 33738
rect 13396 33736 13406 33738
rect 13469 33736 13474 33738
rect 13508 33738 13542 33770
rect 13165 33704 13216 33736
rect 13250 33704 13289 33736
rect 13323 33704 13362 33736
rect 13396 33704 13435 33736
rect 13469 33704 13508 33736
rect 13576 33738 13610 33770
rect 13644 33738 13678 33770
rect 13712 33738 13746 33770
rect 13780 33738 13814 33770
rect 13848 33738 13882 33770
rect 13916 33738 13950 33770
rect 13576 33736 13581 33738
rect 13644 33736 13654 33738
rect 13712 33736 13727 33738
rect 13780 33736 13800 33738
rect 13848 33736 13873 33738
rect 13916 33736 13946 33738
rect 13984 33736 14018 33770
rect 14052 33738 14086 33770
rect 14120 33738 14154 33770
rect 14188 33738 14222 33770
rect 14256 33738 14290 33770
rect 14324 33738 14358 33770
rect 14392 33738 14429 33770
rect 14053 33736 14086 33738
rect 14126 33736 14154 33738
rect 14199 33736 14222 33738
rect 14272 33736 14290 33738
rect 14345 33736 14358 33738
rect 13542 33704 13581 33736
rect 13615 33704 13654 33736
rect 13688 33704 13727 33736
rect 13761 33704 13800 33736
rect 13834 33704 13873 33736
rect 13907 33704 13946 33736
rect 13980 33704 14019 33736
rect 14053 33704 14092 33736
rect 14126 33704 14165 33736
rect 14199 33704 14238 33736
rect 14272 33704 14311 33736
rect 14345 33704 14384 33736
rect 14418 33704 14429 33738
rect 13165 33701 14429 33704
rect 13165 33667 13202 33701
rect 13236 33667 13270 33701
rect 13304 33667 13338 33701
rect 13372 33667 13406 33701
rect 13440 33667 13474 33701
rect 13508 33667 13542 33701
rect 13576 33667 13610 33701
rect 13644 33667 13678 33701
rect 13712 33667 13746 33701
rect 13780 33667 13814 33701
rect 13848 33667 13882 33701
rect 13916 33667 13950 33701
rect 13984 33667 14018 33701
rect 14052 33667 14086 33701
rect 14120 33667 14154 33701
rect 14188 33667 14222 33701
rect 14256 33667 14290 33701
rect 14324 33667 14358 33701
rect 14392 33667 14429 33701
rect 13165 33665 14429 33667
rect 13165 33632 13216 33665
rect 13250 33632 13289 33665
rect 13323 33632 13362 33665
rect 13396 33632 13435 33665
rect 13469 33632 13508 33665
rect 13165 33598 13202 33632
rect 13250 33631 13270 33632
rect 13323 33631 13338 33632
rect 13396 33631 13406 33632
rect 13469 33631 13474 33632
rect 13236 33598 13270 33631
rect 13304 33598 13338 33631
rect 13372 33598 13406 33631
rect 13440 33598 13474 33631
rect 13542 33632 13581 33665
rect 13615 33632 13654 33665
rect 13688 33632 13727 33665
rect 13761 33632 13800 33665
rect 13834 33632 13873 33665
rect 13907 33632 13946 33665
rect 13980 33632 14019 33665
rect 14053 33632 14092 33665
rect 14126 33632 14165 33665
rect 14199 33632 14238 33665
rect 14272 33632 14311 33665
rect 14345 33632 14384 33665
rect 13508 33598 13542 33631
rect 13576 33631 13581 33632
rect 13644 33631 13654 33632
rect 13712 33631 13727 33632
rect 13780 33631 13800 33632
rect 13848 33631 13873 33632
rect 13916 33631 13946 33632
rect 13576 33598 13610 33631
rect 13644 33598 13678 33631
rect 13712 33598 13746 33631
rect 13780 33598 13814 33631
rect 13848 33598 13882 33631
rect 13916 33598 13950 33631
rect 13984 33598 14018 33632
rect 14053 33631 14086 33632
rect 14126 33631 14154 33632
rect 14199 33631 14222 33632
rect 14272 33631 14290 33632
rect 14345 33631 14358 33632
rect 14418 33631 14429 33665
rect 14052 33598 14086 33631
rect 14120 33598 14154 33631
rect 14188 33598 14222 33631
rect 14256 33598 14290 33631
rect 14324 33598 14358 33631
rect 14392 33598 14429 33631
rect 13165 33592 14429 33598
rect 13165 33563 13216 33592
rect 13250 33563 13289 33592
rect 13323 33563 13362 33592
rect 13396 33563 13435 33592
rect 13469 33563 13508 33592
rect 13165 33529 13202 33563
rect 13250 33558 13270 33563
rect 13323 33558 13338 33563
rect 13396 33558 13406 33563
rect 13469 33558 13474 33563
rect 13236 33529 13270 33558
rect 13304 33529 13338 33558
rect 13372 33529 13406 33558
rect 13440 33529 13474 33558
rect 13542 33563 13581 33592
rect 13615 33563 13654 33592
rect 13688 33563 13727 33592
rect 13761 33563 13800 33592
rect 13834 33563 13873 33592
rect 13907 33563 13946 33592
rect 13980 33563 14019 33592
rect 14053 33563 14092 33592
rect 14126 33563 14165 33592
rect 14199 33563 14238 33592
rect 14272 33563 14311 33592
rect 14345 33563 14384 33592
rect 13508 33529 13542 33558
rect 13576 33558 13581 33563
rect 13644 33558 13654 33563
rect 13712 33558 13727 33563
rect 13780 33558 13800 33563
rect 13848 33558 13873 33563
rect 13916 33558 13946 33563
rect 13576 33529 13610 33558
rect 13644 33529 13678 33558
rect 13712 33529 13746 33558
rect 13780 33529 13814 33558
rect 13848 33529 13882 33558
rect 13916 33529 13950 33558
rect 13984 33529 14018 33563
rect 14053 33558 14086 33563
rect 14126 33558 14154 33563
rect 14199 33558 14222 33563
rect 14272 33558 14290 33563
rect 14345 33558 14358 33563
rect 14418 33558 14429 33592
rect 14052 33529 14086 33558
rect 14120 33529 14154 33558
rect 14188 33529 14222 33558
rect 14256 33529 14290 33558
rect 14324 33529 14358 33558
rect 14392 33529 14429 33558
rect 13165 33519 14429 33529
rect 13165 33494 13216 33519
rect 13250 33494 13289 33519
rect 13323 33494 13362 33519
rect 13396 33494 13435 33519
rect 13469 33494 13508 33519
rect 13165 33460 13202 33494
rect 13250 33485 13270 33494
rect 13323 33485 13338 33494
rect 13396 33485 13406 33494
rect 13469 33485 13474 33494
rect 13236 33460 13270 33485
rect 13304 33460 13338 33485
rect 13372 33460 13406 33485
rect 13440 33460 13474 33485
rect 13542 33494 13581 33519
rect 13615 33494 13654 33519
rect 13688 33494 13727 33519
rect 13761 33494 13800 33519
rect 13834 33494 13873 33519
rect 13907 33494 13946 33519
rect 13980 33494 14019 33519
rect 14053 33494 14092 33519
rect 14126 33494 14165 33519
rect 14199 33494 14238 33519
rect 14272 33494 14311 33519
rect 14345 33494 14384 33519
rect 13508 33460 13542 33485
rect 13576 33485 13581 33494
rect 13644 33485 13654 33494
rect 13712 33485 13727 33494
rect 13780 33485 13800 33494
rect 13848 33485 13873 33494
rect 13916 33485 13946 33494
rect 13576 33460 13610 33485
rect 13644 33460 13678 33485
rect 13712 33460 13746 33485
rect 13780 33460 13814 33485
rect 13848 33460 13882 33485
rect 13916 33460 13950 33485
rect 13984 33460 14018 33494
rect 14053 33485 14086 33494
rect 14126 33485 14154 33494
rect 14199 33485 14222 33494
rect 14272 33485 14290 33494
rect 14345 33485 14358 33494
rect 14418 33485 14429 33519
rect 14052 33460 14086 33485
rect 14120 33460 14154 33485
rect 14188 33460 14222 33485
rect 14256 33460 14290 33485
rect 14324 33460 14358 33485
rect 14392 33460 14429 33485
rect 13165 33446 14429 33460
rect 13165 33425 13216 33446
rect 13250 33425 13289 33446
rect 13323 33425 13362 33446
rect 13396 33425 13435 33446
rect 13469 33425 13508 33446
rect 13165 33391 13202 33425
rect 13250 33412 13270 33425
rect 13323 33412 13338 33425
rect 13396 33412 13406 33425
rect 13469 33412 13474 33425
rect 13236 33391 13270 33412
rect 13304 33391 13338 33412
rect 13372 33391 13406 33412
rect 13440 33391 13474 33412
rect 13542 33425 13581 33446
rect 13615 33425 13654 33446
rect 13688 33425 13727 33446
rect 13761 33425 13800 33446
rect 13834 33425 13873 33446
rect 13907 33425 13946 33446
rect 13980 33425 14019 33446
rect 14053 33425 14092 33446
rect 14126 33425 14165 33446
rect 14199 33425 14238 33446
rect 14272 33425 14311 33446
rect 14345 33425 14384 33446
rect 13508 33391 13542 33412
rect 13576 33412 13581 33425
rect 13644 33412 13654 33425
rect 13712 33412 13727 33425
rect 13780 33412 13800 33425
rect 13848 33412 13873 33425
rect 13916 33412 13946 33425
rect 13576 33391 13610 33412
rect 13644 33391 13678 33412
rect 13712 33391 13746 33412
rect 13780 33391 13814 33412
rect 13848 33391 13882 33412
rect 13916 33391 13950 33412
rect 13984 33391 14018 33425
rect 14053 33412 14086 33425
rect 14126 33412 14154 33425
rect 14199 33412 14222 33425
rect 14272 33412 14290 33425
rect 14345 33412 14358 33425
rect 14418 33412 14429 33446
rect 14052 33391 14086 33412
rect 14120 33391 14154 33412
rect 14188 33391 14222 33412
rect 14256 33391 14290 33412
rect 14324 33391 14358 33412
rect 14392 33391 14429 33412
rect 13165 33373 14429 33391
rect 13165 33356 13216 33373
rect 13250 33356 13289 33373
rect 13323 33356 13362 33373
rect 13396 33356 13435 33373
rect 13469 33356 13508 33373
rect 13165 33322 13202 33356
rect 13250 33339 13270 33356
rect 13323 33339 13338 33356
rect 13396 33339 13406 33356
rect 13469 33339 13474 33356
rect 13236 33322 13270 33339
rect 13304 33322 13338 33339
rect 13372 33322 13406 33339
rect 13440 33322 13474 33339
rect 13542 33356 13581 33373
rect 13615 33356 13654 33373
rect 13688 33356 13727 33373
rect 13761 33356 13800 33373
rect 13834 33356 13873 33373
rect 13907 33356 13946 33373
rect 13980 33356 14019 33373
rect 14053 33356 14092 33373
rect 14126 33356 14165 33373
rect 14199 33356 14238 33373
rect 14272 33356 14311 33373
rect 14345 33356 14384 33373
rect 13508 33322 13542 33339
rect 13576 33339 13581 33356
rect 13644 33339 13654 33356
rect 13712 33339 13727 33356
rect 13780 33339 13800 33356
rect 13848 33339 13873 33356
rect 13916 33339 13946 33356
rect 13576 33322 13610 33339
rect 13644 33322 13678 33339
rect 13712 33322 13746 33339
rect 13780 33322 13814 33339
rect 13848 33322 13882 33339
rect 13916 33322 13950 33339
rect 13984 33322 14018 33356
rect 14053 33339 14086 33356
rect 14126 33339 14154 33356
rect 14199 33339 14222 33356
rect 14272 33339 14290 33356
rect 14345 33339 14358 33356
rect 14418 33339 14429 33373
rect 14052 33322 14086 33339
rect 14120 33322 14154 33339
rect 14188 33322 14222 33339
rect 14256 33322 14290 33339
rect 14324 33322 14358 33339
rect 14392 33322 14429 33339
rect 13165 33300 14429 33322
rect 13165 33287 13216 33300
rect 13250 33287 13289 33300
rect 13323 33287 13362 33300
rect 13396 33287 13435 33300
rect 13469 33287 13508 33300
rect 13165 33253 13202 33287
rect 13250 33266 13270 33287
rect 13323 33266 13338 33287
rect 13396 33266 13406 33287
rect 13469 33266 13474 33287
rect 13236 33253 13270 33266
rect 13304 33253 13338 33266
rect 13372 33253 13406 33266
rect 13440 33253 13474 33266
rect 13542 33287 13581 33300
rect 13615 33287 13654 33300
rect 13688 33287 13727 33300
rect 13761 33287 13800 33300
rect 13834 33287 13873 33300
rect 13907 33287 13946 33300
rect 13980 33287 14019 33300
rect 14053 33287 14092 33300
rect 14126 33287 14165 33300
rect 14199 33287 14238 33300
rect 14272 33287 14311 33300
rect 14345 33287 14384 33300
rect 13508 33253 13542 33266
rect 13576 33266 13581 33287
rect 13644 33266 13654 33287
rect 13712 33266 13727 33287
rect 13780 33266 13800 33287
rect 13848 33266 13873 33287
rect 13916 33266 13946 33287
rect 13576 33253 13610 33266
rect 13644 33253 13678 33266
rect 13712 33253 13746 33266
rect 13780 33253 13814 33266
rect 13848 33253 13882 33266
rect 13916 33253 13950 33266
rect 13984 33253 14018 33287
rect 14053 33266 14086 33287
rect 14126 33266 14154 33287
rect 14199 33266 14222 33287
rect 14272 33266 14290 33287
rect 14345 33266 14358 33287
rect 14418 33266 14429 33300
rect 14052 33253 14086 33266
rect 14120 33253 14154 33266
rect 14188 33253 14222 33266
rect 14256 33253 14290 33266
rect 14324 33253 14358 33266
rect 14392 33253 14429 33266
rect 13165 33227 14429 33253
rect 13165 33218 13216 33227
rect 13250 33218 13289 33227
rect 13323 33218 13362 33227
rect 13396 33218 13435 33227
rect 13469 33218 13508 33227
rect 13165 33184 13202 33218
rect 13250 33193 13270 33218
rect 13323 33193 13338 33218
rect 13396 33193 13406 33218
rect 13469 33193 13474 33218
rect 13236 33184 13270 33193
rect 13304 33184 13338 33193
rect 13372 33184 13406 33193
rect 13440 33184 13474 33193
rect 13542 33218 13581 33227
rect 13615 33218 13654 33227
rect 13688 33218 13727 33227
rect 13761 33218 13800 33227
rect 13834 33218 13873 33227
rect 13907 33218 13946 33227
rect 13980 33218 14019 33227
rect 14053 33218 14092 33227
rect 14126 33218 14165 33227
rect 14199 33218 14238 33227
rect 14272 33218 14311 33227
rect 14345 33218 14384 33227
rect 13508 33184 13542 33193
rect 13576 33193 13581 33218
rect 13644 33193 13654 33218
rect 13712 33193 13727 33218
rect 13780 33193 13800 33218
rect 13848 33193 13873 33218
rect 13916 33193 13946 33218
rect 13576 33184 13610 33193
rect 13644 33184 13678 33193
rect 13712 33184 13746 33193
rect 13780 33184 13814 33193
rect 13848 33184 13882 33193
rect 13916 33184 13950 33193
rect 13984 33184 14018 33218
rect 14053 33193 14086 33218
rect 14126 33193 14154 33218
rect 14199 33193 14222 33218
rect 14272 33193 14290 33218
rect 14345 33193 14358 33218
rect 14418 33193 14429 33227
rect 14052 33184 14086 33193
rect 14120 33184 14154 33193
rect 14188 33184 14222 33193
rect 14256 33184 14290 33193
rect 14324 33184 14358 33193
rect 14392 33184 14429 33193
rect 13165 33154 14429 33184
rect 13165 33149 13216 33154
rect 13250 33149 13289 33154
rect 13323 33149 13362 33154
rect 13396 33149 13435 33154
rect 13469 33149 13508 33154
rect 13165 33115 13202 33149
rect 13250 33120 13270 33149
rect 13323 33120 13338 33149
rect 13396 33120 13406 33149
rect 13469 33120 13474 33149
rect 13236 33115 13270 33120
rect 13304 33115 13338 33120
rect 13372 33115 13406 33120
rect 13440 33115 13474 33120
rect 13542 33149 13581 33154
rect 13615 33149 13654 33154
rect 13688 33149 13727 33154
rect 13761 33149 13800 33154
rect 13834 33149 13873 33154
rect 13907 33149 13946 33154
rect 13980 33149 14019 33154
rect 14053 33149 14092 33154
rect 14126 33149 14165 33154
rect 14199 33149 14238 33154
rect 14272 33149 14311 33154
rect 14345 33149 14384 33154
rect 13508 33115 13542 33120
rect 13576 33120 13581 33149
rect 13644 33120 13654 33149
rect 13712 33120 13727 33149
rect 13780 33120 13800 33149
rect 13848 33120 13873 33149
rect 13916 33120 13946 33149
rect 13576 33115 13610 33120
rect 13644 33115 13678 33120
rect 13712 33115 13746 33120
rect 13780 33115 13814 33120
rect 13848 33115 13882 33120
rect 13916 33115 13950 33120
rect 13984 33115 14018 33149
rect 14053 33120 14086 33149
rect 14126 33120 14154 33149
rect 14199 33120 14222 33149
rect 14272 33120 14290 33149
rect 14345 33120 14358 33149
rect 14418 33120 14429 33154
rect 14052 33115 14086 33120
rect 14120 33115 14154 33120
rect 14188 33115 14222 33120
rect 14256 33115 14290 33120
rect 14324 33115 14358 33120
rect 14392 33115 14429 33120
rect 13165 33081 14429 33115
rect 13165 33080 13216 33081
rect 13250 33080 13289 33081
rect 13323 33080 13362 33081
rect 13396 33080 13435 33081
rect 13469 33080 13508 33081
rect 13165 33046 13202 33080
rect 13250 33047 13270 33080
rect 13323 33047 13338 33080
rect 13396 33047 13406 33080
rect 13469 33047 13474 33080
rect 13236 33046 13270 33047
rect 13304 33046 13338 33047
rect 13372 33046 13406 33047
rect 13440 33046 13474 33047
rect 13542 33080 13581 33081
rect 13615 33080 13654 33081
rect 13688 33080 13727 33081
rect 13761 33080 13800 33081
rect 13834 33080 13873 33081
rect 13907 33080 13946 33081
rect 13980 33080 14019 33081
rect 14053 33080 14092 33081
rect 14126 33080 14165 33081
rect 14199 33080 14238 33081
rect 14272 33080 14311 33081
rect 14345 33080 14384 33081
rect 13508 33046 13542 33047
rect 13576 33047 13581 33080
rect 13644 33047 13654 33080
rect 13712 33047 13727 33080
rect 13780 33047 13800 33080
rect 13848 33047 13873 33080
rect 13916 33047 13946 33080
rect 13576 33046 13610 33047
rect 13644 33046 13678 33047
rect 13712 33046 13746 33047
rect 13780 33046 13814 33047
rect 13848 33046 13882 33047
rect 13916 33046 13950 33047
rect 13984 33046 14018 33080
rect 14053 33047 14086 33080
rect 14126 33047 14154 33080
rect 14199 33047 14222 33080
rect 14272 33047 14290 33080
rect 14345 33047 14358 33080
rect 14418 33047 14429 33081
rect 14052 33046 14086 33047
rect 14120 33046 14154 33047
rect 14188 33046 14222 33047
rect 14256 33046 14290 33047
rect 14324 33046 14358 33047
rect 14392 33046 14429 33047
rect 13165 33011 14429 33046
rect 13165 32977 13202 33011
rect 13236 33008 13270 33011
rect 13304 33008 13338 33011
rect 13372 33008 13406 33011
rect 13440 33008 13474 33011
rect 13250 32977 13270 33008
rect 13323 32977 13338 33008
rect 13396 32977 13406 33008
rect 13469 32977 13474 33008
rect 13508 33008 13542 33011
rect 13165 32974 13216 32977
rect 13250 32974 13289 32977
rect 13323 32974 13362 32977
rect 13396 32974 13435 32977
rect 13469 32974 13508 32977
rect 13576 33008 13610 33011
rect 13644 33008 13678 33011
rect 13712 33008 13746 33011
rect 13780 33008 13814 33011
rect 13848 33008 13882 33011
rect 13916 33008 13950 33011
rect 13576 32977 13581 33008
rect 13644 32977 13654 33008
rect 13712 32977 13727 33008
rect 13780 32977 13800 33008
rect 13848 32977 13873 33008
rect 13916 32977 13946 33008
rect 13984 32977 14018 33011
rect 14052 33008 14086 33011
rect 14120 33008 14154 33011
rect 14188 33008 14222 33011
rect 14256 33008 14290 33011
rect 14324 33008 14358 33011
rect 14392 33008 14429 33011
rect 14053 32977 14086 33008
rect 14126 32977 14154 33008
rect 14199 32977 14222 33008
rect 14272 32977 14290 33008
rect 14345 32977 14358 33008
rect 13542 32974 13581 32977
rect 13615 32974 13654 32977
rect 13688 32974 13727 32977
rect 13761 32974 13800 32977
rect 13834 32974 13873 32977
rect 13907 32974 13946 32977
rect 13980 32974 14019 32977
rect 14053 32974 14092 32977
rect 14126 32974 14165 32977
rect 14199 32974 14238 32977
rect 14272 32974 14311 32977
rect 14345 32974 14384 32977
rect 14418 32974 14429 33008
rect 13165 32942 14429 32974
rect 13165 32908 13202 32942
rect 13236 32935 13270 32942
rect 13304 32935 13338 32942
rect 13372 32935 13406 32942
rect 13440 32935 13474 32942
rect 13250 32908 13270 32935
rect 13323 32908 13338 32935
rect 13396 32908 13406 32935
rect 13469 32908 13474 32935
rect 13508 32935 13542 32942
rect 13165 32901 13216 32908
rect 13250 32901 13289 32908
rect 13323 32901 13362 32908
rect 13396 32901 13435 32908
rect 13469 32901 13508 32908
rect 13576 32935 13610 32942
rect 13644 32935 13678 32942
rect 13712 32935 13746 32942
rect 13780 32935 13814 32942
rect 13848 32935 13882 32942
rect 13916 32935 13950 32942
rect 13576 32908 13581 32935
rect 13644 32908 13654 32935
rect 13712 32908 13727 32935
rect 13780 32908 13800 32935
rect 13848 32908 13873 32935
rect 13916 32908 13946 32935
rect 13984 32908 14018 32942
rect 14052 32935 14086 32942
rect 14120 32935 14154 32942
rect 14188 32935 14222 32942
rect 14256 32935 14290 32942
rect 14324 32935 14358 32942
rect 14392 32935 14429 32942
rect 14053 32908 14086 32935
rect 14126 32908 14154 32935
rect 14199 32908 14222 32935
rect 14272 32908 14290 32935
rect 14345 32908 14358 32935
rect 13542 32901 13581 32908
rect 13615 32901 13654 32908
rect 13688 32901 13727 32908
rect 13761 32901 13800 32908
rect 13834 32901 13873 32908
rect 13907 32901 13946 32908
rect 13980 32901 14019 32908
rect 14053 32901 14092 32908
rect 14126 32901 14165 32908
rect 14199 32901 14238 32908
rect 14272 32901 14311 32908
rect 14345 32901 14384 32908
rect 14418 32901 14429 32935
rect 13165 32873 14429 32901
rect 13165 32839 13202 32873
rect 13236 32862 13270 32873
rect 13304 32862 13338 32873
rect 13372 32862 13406 32873
rect 13440 32862 13474 32873
rect 13250 32839 13270 32862
rect 13323 32839 13338 32862
rect 13396 32839 13406 32862
rect 13469 32839 13474 32862
rect 13508 32862 13542 32873
rect 13165 32828 13216 32839
rect 13250 32828 13289 32839
rect 13323 32828 13362 32839
rect 13396 32828 13435 32839
rect 13469 32828 13508 32839
rect 13576 32862 13610 32873
rect 13644 32862 13678 32873
rect 13712 32862 13746 32873
rect 13780 32862 13814 32873
rect 13848 32862 13882 32873
rect 13916 32862 13950 32873
rect 13576 32839 13581 32862
rect 13644 32839 13654 32862
rect 13712 32839 13727 32862
rect 13780 32839 13800 32862
rect 13848 32839 13873 32862
rect 13916 32839 13946 32862
rect 13984 32839 14018 32873
rect 14052 32862 14086 32873
rect 14120 32862 14154 32873
rect 14188 32862 14222 32873
rect 14256 32862 14290 32873
rect 14324 32862 14358 32873
rect 14392 32862 14429 32873
rect 14053 32839 14086 32862
rect 14126 32839 14154 32862
rect 14199 32839 14222 32862
rect 14272 32839 14290 32862
rect 14345 32839 14358 32862
rect 13542 32828 13581 32839
rect 13615 32828 13654 32839
rect 13688 32828 13727 32839
rect 13761 32828 13800 32839
rect 13834 32828 13873 32839
rect 13907 32828 13946 32839
rect 13980 32828 14019 32839
rect 14053 32828 14092 32839
rect 14126 32828 14165 32839
rect 14199 32828 14238 32839
rect 14272 32828 14311 32839
rect 14345 32828 14384 32839
rect 14418 32828 14429 32862
rect 13165 32804 14429 32828
rect 13165 32770 13202 32804
rect 13236 32789 13270 32804
rect 13304 32789 13338 32804
rect 13372 32789 13406 32804
rect 13440 32789 13474 32804
rect 13250 32770 13270 32789
rect 13323 32770 13338 32789
rect 13396 32770 13406 32789
rect 13469 32770 13474 32789
rect 13508 32789 13542 32804
rect 13165 32755 13216 32770
rect 13250 32755 13289 32770
rect 13323 32755 13362 32770
rect 13396 32755 13435 32770
rect 13469 32755 13508 32770
rect 13576 32789 13610 32804
rect 13644 32789 13678 32804
rect 13712 32789 13746 32804
rect 13780 32789 13814 32804
rect 13848 32789 13882 32804
rect 13916 32789 13950 32804
rect 13576 32770 13581 32789
rect 13644 32770 13654 32789
rect 13712 32770 13727 32789
rect 13780 32770 13800 32789
rect 13848 32770 13873 32789
rect 13916 32770 13946 32789
rect 13984 32770 14018 32804
rect 14052 32789 14086 32804
rect 14120 32789 14154 32804
rect 14188 32789 14222 32804
rect 14256 32789 14290 32804
rect 14324 32789 14358 32804
rect 14392 32789 14429 32804
rect 14053 32770 14086 32789
rect 14126 32770 14154 32789
rect 14199 32770 14222 32789
rect 14272 32770 14290 32789
rect 14345 32770 14358 32789
rect 13542 32755 13581 32770
rect 13615 32755 13654 32770
rect 13688 32755 13727 32770
rect 13761 32755 13800 32770
rect 13834 32755 13873 32770
rect 13907 32755 13946 32770
rect 13980 32755 14019 32770
rect 14053 32755 14092 32770
rect 14126 32755 14165 32770
rect 14199 32755 14238 32770
rect 14272 32755 14311 32770
rect 14345 32755 14384 32770
rect 14418 32755 14429 32789
rect 13165 32735 14429 32755
rect 13165 32701 13202 32735
rect 13236 32716 13270 32735
rect 13304 32716 13338 32735
rect 13372 32716 13406 32735
rect 13440 32716 13474 32735
rect 13250 32701 13270 32716
rect 13323 32701 13338 32716
rect 13396 32701 13406 32716
rect 13469 32701 13474 32716
rect 13508 32716 13542 32735
rect 13165 32682 13216 32701
rect 13250 32682 13289 32701
rect 13323 32682 13362 32701
rect 13396 32682 13435 32701
rect 13469 32682 13508 32701
rect 13576 32716 13610 32735
rect 13644 32716 13678 32735
rect 13712 32716 13746 32735
rect 13780 32716 13814 32735
rect 13848 32716 13882 32735
rect 13916 32716 13950 32735
rect 13576 32701 13581 32716
rect 13644 32701 13654 32716
rect 13712 32701 13727 32716
rect 13780 32701 13800 32716
rect 13848 32701 13873 32716
rect 13916 32701 13946 32716
rect 13984 32701 14018 32735
rect 14052 32716 14086 32735
rect 14120 32716 14154 32735
rect 14188 32716 14222 32735
rect 14256 32716 14290 32735
rect 14324 32716 14358 32735
rect 14392 32716 14429 32735
rect 14053 32701 14086 32716
rect 14126 32701 14154 32716
rect 14199 32701 14222 32716
rect 14272 32701 14290 32716
rect 14345 32701 14358 32716
rect 13542 32682 13581 32701
rect 13615 32682 13654 32701
rect 13688 32682 13727 32701
rect 13761 32682 13800 32701
rect 13834 32682 13873 32701
rect 13907 32682 13946 32701
rect 13980 32682 14019 32701
rect 14053 32682 14092 32701
rect 14126 32682 14165 32701
rect 14199 32682 14238 32701
rect 14272 32682 14311 32701
rect 14345 32682 14384 32701
rect 14418 32682 14429 32716
rect 13165 32666 14429 32682
rect 13165 32632 13202 32666
rect 13236 32643 13270 32666
rect 13304 32643 13338 32666
rect 13372 32643 13406 32666
rect 13440 32643 13474 32666
rect 13250 32632 13270 32643
rect 13323 32632 13338 32643
rect 13396 32632 13406 32643
rect 13469 32632 13474 32643
rect 13508 32643 13542 32666
rect 13165 32609 13216 32632
rect 13250 32609 13289 32632
rect 13323 32609 13362 32632
rect 13396 32609 13435 32632
rect 13469 32609 13508 32632
rect 13576 32643 13610 32666
rect 13644 32643 13678 32666
rect 13712 32643 13746 32666
rect 13780 32643 13814 32666
rect 13848 32643 13882 32666
rect 13916 32643 13950 32666
rect 13576 32632 13581 32643
rect 13644 32632 13654 32643
rect 13712 32632 13727 32643
rect 13780 32632 13800 32643
rect 13848 32632 13873 32643
rect 13916 32632 13946 32643
rect 13984 32632 14018 32666
rect 14052 32643 14086 32666
rect 14120 32643 14154 32666
rect 14188 32643 14222 32666
rect 14256 32643 14290 32666
rect 14324 32643 14358 32666
rect 14392 32643 14429 32666
rect 14053 32632 14086 32643
rect 14126 32632 14154 32643
rect 14199 32632 14222 32643
rect 14272 32632 14290 32643
rect 14345 32632 14358 32643
rect 13542 32609 13581 32632
rect 13615 32609 13654 32632
rect 13688 32609 13727 32632
rect 13761 32609 13800 32632
rect 13834 32609 13873 32632
rect 13907 32609 13946 32632
rect 13980 32609 14019 32632
rect 14053 32609 14092 32632
rect 14126 32609 14165 32632
rect 14199 32609 14238 32632
rect 14272 32609 14311 32632
rect 14345 32609 14384 32632
rect 14418 32609 14429 32643
rect 13165 32597 14429 32609
rect 13165 32563 13202 32597
rect 13236 32570 13270 32597
rect 13304 32570 13338 32597
rect 13372 32570 13406 32597
rect 13440 32570 13474 32597
rect 13250 32563 13270 32570
rect 13323 32563 13338 32570
rect 13396 32563 13406 32570
rect 13469 32563 13474 32570
rect 13508 32570 13542 32597
rect 13165 32536 13216 32563
rect 13250 32536 13289 32563
rect 13323 32536 13362 32563
rect 13396 32536 13435 32563
rect 13469 32536 13508 32563
rect 13576 32570 13610 32597
rect 13644 32570 13678 32597
rect 13712 32570 13746 32597
rect 13780 32570 13814 32597
rect 13848 32570 13882 32597
rect 13916 32570 13950 32597
rect 13576 32563 13581 32570
rect 13644 32563 13654 32570
rect 13712 32563 13727 32570
rect 13780 32563 13800 32570
rect 13848 32563 13873 32570
rect 13916 32563 13946 32570
rect 13984 32563 14018 32597
rect 14052 32570 14086 32597
rect 14120 32570 14154 32597
rect 14188 32570 14222 32597
rect 14256 32570 14290 32597
rect 14324 32570 14358 32597
rect 14392 32570 14429 32597
rect 14053 32563 14086 32570
rect 14126 32563 14154 32570
rect 14199 32563 14222 32570
rect 14272 32563 14290 32570
rect 14345 32563 14358 32570
rect 13542 32536 13581 32563
rect 13615 32536 13654 32563
rect 13688 32536 13727 32563
rect 13761 32536 13800 32563
rect 13834 32536 13873 32563
rect 13907 32536 13946 32563
rect 13980 32536 14019 32563
rect 14053 32536 14092 32563
rect 14126 32536 14165 32563
rect 14199 32536 14238 32563
rect 14272 32536 14311 32563
rect 14345 32536 14384 32563
rect 14418 32536 14429 32570
rect 13165 32528 14429 32536
rect 13165 32494 13202 32528
rect 13236 32497 13270 32528
rect 13304 32497 13338 32528
rect 13372 32497 13406 32528
rect 13440 32497 13474 32528
rect 13250 32494 13270 32497
rect 13323 32494 13338 32497
rect 13396 32494 13406 32497
rect 13469 32494 13474 32497
rect 13508 32497 13542 32528
rect 13165 32463 13216 32494
rect 13250 32463 13289 32494
rect 13323 32463 13362 32494
rect 13396 32463 13435 32494
rect 13469 32463 13508 32494
rect 13576 32497 13610 32528
rect 13644 32497 13678 32528
rect 13712 32497 13746 32528
rect 13780 32497 13814 32528
rect 13848 32497 13882 32528
rect 13916 32497 13950 32528
rect 13576 32494 13581 32497
rect 13644 32494 13654 32497
rect 13712 32494 13727 32497
rect 13780 32494 13800 32497
rect 13848 32494 13873 32497
rect 13916 32494 13946 32497
rect 13984 32494 14018 32528
rect 14052 32497 14086 32528
rect 14120 32497 14154 32528
rect 14188 32497 14222 32528
rect 14256 32497 14290 32528
rect 14324 32497 14358 32528
rect 14392 32497 14429 32528
rect 14053 32494 14086 32497
rect 14126 32494 14154 32497
rect 14199 32494 14222 32497
rect 14272 32494 14290 32497
rect 14345 32494 14358 32497
rect 13542 32463 13581 32494
rect 13615 32463 13654 32494
rect 13688 32463 13727 32494
rect 13761 32463 13800 32494
rect 13834 32463 13873 32494
rect 13907 32463 13946 32494
rect 13980 32463 14019 32494
rect 14053 32463 14092 32494
rect 14126 32463 14165 32494
rect 14199 32463 14238 32494
rect 14272 32463 14311 32494
rect 14345 32463 14384 32494
rect 14418 32463 14429 32497
rect 13165 32459 14429 32463
rect 13165 32425 13202 32459
rect 13236 32425 13270 32459
rect 13304 32425 13338 32459
rect 13372 32425 13406 32459
rect 13440 32425 13474 32459
rect 13508 32425 13542 32459
rect 13576 32425 13610 32459
rect 13644 32425 13678 32459
rect 13712 32425 13746 32459
rect 13780 32425 13814 32459
rect 13848 32425 13882 32459
rect 13916 32425 13950 32459
rect 13984 32425 14018 32459
rect 14052 32425 14086 32459
rect 14120 32425 14154 32459
rect 14188 32425 14222 32459
rect 14256 32425 14290 32459
rect 14324 32425 14358 32459
rect 14392 32425 14429 32459
rect 13165 32424 14429 32425
rect 13165 32390 13216 32424
rect 13250 32390 13289 32424
rect 13323 32390 13362 32424
rect 13396 32390 13435 32424
rect 13469 32390 13508 32424
rect 13542 32390 13581 32424
rect 13615 32390 13654 32424
rect 13688 32390 13727 32424
rect 13761 32390 13800 32424
rect 13834 32390 13873 32424
rect 13907 32390 13946 32424
rect 13980 32390 14019 32424
rect 14053 32390 14092 32424
rect 14126 32390 14165 32424
rect 14199 32390 14238 32424
rect 14272 32390 14311 32424
rect 14345 32390 14384 32424
rect 14418 32390 14429 32424
rect 13165 32356 13202 32390
rect 13236 32356 13270 32390
rect 13304 32356 13338 32390
rect 13372 32356 13406 32390
rect 13440 32356 13474 32390
rect 13508 32356 13542 32390
rect 13576 32356 13610 32390
rect 13644 32356 13678 32390
rect 13712 32356 13746 32390
rect 13780 32356 13814 32390
rect 13848 32356 13882 32390
rect 13916 32356 13950 32390
rect 13984 32356 14018 32390
rect 14052 32356 14086 32390
rect 14120 32356 14154 32390
rect 14188 32356 14222 32390
rect 14256 32356 14290 32390
rect 14324 32356 14358 32390
rect 14392 32356 14429 32390
rect 13165 32351 14429 32356
rect 13165 32321 13216 32351
rect 13250 32321 13289 32351
rect 13323 32321 13362 32351
rect 13396 32321 13435 32351
rect 13469 32321 13508 32351
rect 13165 32287 13202 32321
rect 13250 32317 13270 32321
rect 13323 32317 13338 32321
rect 13396 32317 13406 32321
rect 13469 32317 13474 32321
rect 13236 32287 13270 32317
rect 13304 32287 13338 32317
rect 13372 32287 13406 32317
rect 13440 32287 13474 32317
rect 13542 32321 13581 32351
rect 13615 32321 13654 32351
rect 13688 32321 13727 32351
rect 13761 32321 13800 32351
rect 13834 32321 13873 32351
rect 13907 32321 13946 32351
rect 13980 32321 14019 32351
rect 14053 32321 14092 32351
rect 14126 32321 14165 32351
rect 14199 32321 14238 32351
rect 14272 32321 14311 32351
rect 14345 32321 14384 32351
rect 13508 32287 13542 32317
rect 13576 32317 13581 32321
rect 13644 32317 13654 32321
rect 13712 32317 13727 32321
rect 13780 32317 13800 32321
rect 13848 32317 13873 32321
rect 13916 32317 13946 32321
rect 13576 32287 13610 32317
rect 13644 32287 13678 32317
rect 13712 32287 13746 32317
rect 13780 32287 13814 32317
rect 13848 32287 13882 32317
rect 13916 32287 13950 32317
rect 13984 32287 14018 32321
rect 14053 32317 14086 32321
rect 14126 32317 14154 32321
rect 14199 32317 14222 32321
rect 14272 32317 14290 32321
rect 14345 32317 14358 32321
rect 14418 32317 14429 32351
rect 14052 32287 14086 32317
rect 14120 32287 14154 32317
rect 14188 32287 14222 32317
rect 14256 32287 14290 32317
rect 14324 32287 14358 32317
rect 14392 32287 14429 32317
rect 13165 32278 14429 32287
rect 13165 32252 13216 32278
rect 13250 32252 13289 32278
rect 13323 32252 13362 32278
rect 13396 32252 13435 32278
rect 13469 32252 13508 32278
rect 13165 32218 13202 32252
rect 13250 32244 13270 32252
rect 13323 32244 13338 32252
rect 13396 32244 13406 32252
rect 13469 32244 13474 32252
rect 13236 32218 13270 32244
rect 13304 32218 13338 32244
rect 13372 32218 13406 32244
rect 13440 32218 13474 32244
rect 13542 32252 13581 32278
rect 13615 32252 13654 32278
rect 13688 32252 13727 32278
rect 13761 32252 13800 32278
rect 13834 32252 13873 32278
rect 13907 32252 13946 32278
rect 13980 32252 14019 32278
rect 14053 32252 14092 32278
rect 14126 32252 14165 32278
rect 14199 32252 14238 32278
rect 14272 32252 14311 32278
rect 14345 32252 14384 32278
rect 13508 32218 13542 32244
rect 13576 32244 13581 32252
rect 13644 32244 13654 32252
rect 13712 32244 13727 32252
rect 13780 32244 13800 32252
rect 13848 32244 13873 32252
rect 13916 32244 13946 32252
rect 13576 32218 13610 32244
rect 13644 32218 13678 32244
rect 13712 32218 13746 32244
rect 13780 32218 13814 32244
rect 13848 32218 13882 32244
rect 13916 32218 13950 32244
rect 13984 32218 14018 32252
rect 14053 32244 14086 32252
rect 14126 32244 14154 32252
rect 14199 32244 14222 32252
rect 14272 32244 14290 32252
rect 14345 32244 14358 32252
rect 14418 32244 14429 32278
rect 14052 32218 14086 32244
rect 14120 32218 14154 32244
rect 14188 32218 14222 32244
rect 14256 32218 14290 32244
rect 14324 32218 14358 32244
rect 14392 32218 14429 32244
rect 13165 32205 14429 32218
rect 13165 32183 13216 32205
rect 13250 32183 13289 32205
rect 13323 32183 13362 32205
rect 13396 32183 13435 32205
rect 13469 32183 13508 32205
rect 13165 32149 13202 32183
rect 13250 32171 13270 32183
rect 13323 32171 13338 32183
rect 13396 32171 13406 32183
rect 13469 32171 13474 32183
rect 13236 32149 13270 32171
rect 13304 32149 13338 32171
rect 13372 32149 13406 32171
rect 13440 32149 13474 32171
rect 13542 32183 13581 32205
rect 13615 32183 13654 32205
rect 13688 32183 13727 32205
rect 13761 32183 13800 32205
rect 13834 32183 13873 32205
rect 13907 32183 13946 32205
rect 13980 32183 14019 32205
rect 14053 32183 14092 32205
rect 14126 32183 14165 32205
rect 14199 32183 14238 32205
rect 14272 32183 14311 32205
rect 14345 32183 14384 32205
rect 13508 32149 13542 32171
rect 13576 32171 13581 32183
rect 13644 32171 13654 32183
rect 13712 32171 13727 32183
rect 13780 32171 13800 32183
rect 13848 32171 13873 32183
rect 13916 32171 13946 32183
rect 13576 32149 13610 32171
rect 13644 32149 13678 32171
rect 13712 32149 13746 32171
rect 13780 32149 13814 32171
rect 13848 32149 13882 32171
rect 13916 32149 13950 32171
rect 13984 32149 14018 32183
rect 14053 32171 14086 32183
rect 14126 32171 14154 32183
rect 14199 32171 14222 32183
rect 14272 32171 14290 32183
rect 14345 32171 14358 32183
rect 14418 32171 14429 32205
rect 14052 32149 14086 32171
rect 14120 32149 14154 32171
rect 14188 32149 14222 32171
rect 14256 32149 14290 32171
rect 14324 32149 14358 32171
rect 14392 32149 14429 32171
rect 13165 32132 14429 32149
rect 13165 32114 13216 32132
rect 13250 32114 13289 32132
rect 13323 32114 13362 32132
rect 13396 32114 13435 32132
rect 13469 32114 13508 32132
rect 13165 32080 13202 32114
rect 13250 32098 13270 32114
rect 13323 32098 13338 32114
rect 13396 32098 13406 32114
rect 13469 32098 13474 32114
rect 13236 32080 13270 32098
rect 13304 32080 13338 32098
rect 13372 32080 13406 32098
rect 13440 32080 13474 32098
rect 13542 32114 13581 32132
rect 13615 32114 13654 32132
rect 13688 32114 13727 32132
rect 13761 32114 13800 32132
rect 13834 32114 13873 32132
rect 13907 32114 13946 32132
rect 13980 32114 14019 32132
rect 14053 32114 14092 32132
rect 14126 32114 14165 32132
rect 14199 32114 14238 32132
rect 14272 32114 14311 32132
rect 14345 32114 14384 32132
rect 13508 32080 13542 32098
rect 13576 32098 13581 32114
rect 13644 32098 13654 32114
rect 13712 32098 13727 32114
rect 13780 32098 13800 32114
rect 13848 32098 13873 32114
rect 13916 32098 13946 32114
rect 13576 32080 13610 32098
rect 13644 32080 13678 32098
rect 13712 32080 13746 32098
rect 13780 32080 13814 32098
rect 13848 32080 13882 32098
rect 13916 32080 13950 32098
rect 13984 32080 14018 32114
rect 14053 32098 14086 32114
rect 14126 32098 14154 32114
rect 14199 32098 14222 32114
rect 14272 32098 14290 32114
rect 14345 32098 14358 32114
rect 14418 32098 14429 32132
rect 14052 32080 14086 32098
rect 14120 32080 14154 32098
rect 14188 32080 14222 32098
rect 14256 32080 14290 32098
rect 14324 32080 14358 32098
rect 14392 32080 14429 32098
rect 13165 32059 14429 32080
rect 13165 32045 13216 32059
rect 13250 32045 13289 32059
rect 13323 32045 13362 32059
rect 13396 32045 13435 32059
rect 13469 32045 13508 32059
rect 13165 32011 13202 32045
rect 13250 32025 13270 32045
rect 13323 32025 13338 32045
rect 13396 32025 13406 32045
rect 13469 32025 13474 32045
rect 13236 32011 13270 32025
rect 13304 32011 13338 32025
rect 13372 32011 13406 32025
rect 13440 32011 13474 32025
rect 13542 32045 13581 32059
rect 13615 32045 13654 32059
rect 13688 32045 13727 32059
rect 13761 32045 13800 32059
rect 13834 32045 13873 32059
rect 13907 32045 13946 32059
rect 13980 32045 14019 32059
rect 14053 32045 14092 32059
rect 14126 32045 14165 32059
rect 14199 32045 14238 32059
rect 14272 32045 14311 32059
rect 14345 32045 14384 32059
rect 13508 32011 13542 32025
rect 13576 32025 13581 32045
rect 13644 32025 13654 32045
rect 13712 32025 13727 32045
rect 13780 32025 13800 32045
rect 13848 32025 13873 32045
rect 13916 32025 13946 32045
rect 13576 32011 13610 32025
rect 13644 32011 13678 32025
rect 13712 32011 13746 32025
rect 13780 32011 13814 32025
rect 13848 32011 13882 32025
rect 13916 32011 13950 32025
rect 13984 32011 14018 32045
rect 14053 32025 14086 32045
rect 14126 32025 14154 32045
rect 14199 32025 14222 32045
rect 14272 32025 14290 32045
rect 14345 32025 14358 32045
rect 14418 32025 14429 32059
rect 14052 32011 14086 32025
rect 14120 32011 14154 32025
rect 14188 32011 14222 32025
rect 14256 32011 14290 32025
rect 14324 32011 14358 32025
rect 14392 32011 14429 32025
rect 13165 31986 14429 32011
rect 13165 31976 13216 31986
rect 13250 31976 13289 31986
rect 13323 31976 13362 31986
rect 13396 31976 13435 31986
rect 13469 31976 13508 31986
rect 13165 31942 13202 31976
rect 13250 31952 13270 31976
rect 13323 31952 13338 31976
rect 13396 31952 13406 31976
rect 13469 31952 13474 31976
rect 13236 31942 13270 31952
rect 13304 31942 13338 31952
rect 13372 31942 13406 31952
rect 13440 31942 13474 31952
rect 13542 31976 13581 31986
rect 13615 31976 13654 31986
rect 13688 31976 13727 31986
rect 13761 31976 13800 31986
rect 13834 31976 13873 31986
rect 13907 31976 13946 31986
rect 13980 31976 14019 31986
rect 14053 31976 14092 31986
rect 14126 31976 14165 31986
rect 14199 31976 14238 31986
rect 14272 31976 14311 31986
rect 14345 31976 14384 31986
rect 13508 31942 13542 31952
rect 13576 31952 13581 31976
rect 13644 31952 13654 31976
rect 13712 31952 13727 31976
rect 13780 31952 13800 31976
rect 13848 31952 13873 31976
rect 13916 31952 13946 31976
rect 13576 31942 13610 31952
rect 13644 31942 13678 31952
rect 13712 31942 13746 31952
rect 13780 31942 13814 31952
rect 13848 31942 13882 31952
rect 13916 31942 13950 31952
rect 13984 31942 14018 31976
rect 14053 31952 14086 31976
rect 14126 31952 14154 31976
rect 14199 31952 14222 31976
rect 14272 31952 14290 31976
rect 14345 31952 14358 31976
rect 14418 31952 14429 31986
rect 14052 31942 14086 31952
rect 14120 31942 14154 31952
rect 14188 31942 14222 31952
rect 14256 31942 14290 31952
rect 14324 31942 14358 31952
rect 14392 31942 14429 31952
rect 13165 31913 14429 31942
rect 13165 31907 13216 31913
rect 13250 31907 13289 31913
rect 13323 31907 13362 31913
rect 13396 31907 13435 31913
rect 13469 31907 13508 31913
rect 13165 31873 13202 31907
rect 13250 31879 13270 31907
rect 13323 31879 13338 31907
rect 13396 31879 13406 31907
rect 13469 31879 13474 31907
rect 13236 31873 13270 31879
rect 13304 31873 13338 31879
rect 13372 31873 13406 31879
rect 13440 31873 13474 31879
rect 13542 31907 13581 31913
rect 13615 31907 13654 31913
rect 13688 31907 13727 31913
rect 13761 31907 13800 31913
rect 13834 31907 13873 31913
rect 13907 31907 13946 31913
rect 13980 31907 14019 31913
rect 14053 31907 14092 31913
rect 14126 31907 14165 31913
rect 14199 31907 14238 31913
rect 14272 31907 14311 31913
rect 14345 31907 14384 31913
rect 13508 31873 13542 31879
rect 13576 31879 13581 31907
rect 13644 31879 13654 31907
rect 13712 31879 13727 31907
rect 13780 31879 13800 31907
rect 13848 31879 13873 31907
rect 13916 31879 13946 31907
rect 13576 31873 13610 31879
rect 13644 31873 13678 31879
rect 13712 31873 13746 31879
rect 13780 31873 13814 31879
rect 13848 31873 13882 31879
rect 13916 31873 13950 31879
rect 13984 31873 14018 31907
rect 14053 31879 14086 31907
rect 14126 31879 14154 31907
rect 14199 31879 14222 31907
rect 14272 31879 14290 31907
rect 14345 31879 14358 31907
rect 14418 31879 14429 31913
rect 14052 31873 14086 31879
rect 14120 31873 14154 31879
rect 14188 31873 14222 31879
rect 14256 31873 14290 31879
rect 14324 31873 14358 31879
rect 14392 31873 14429 31879
rect 13165 31840 14429 31873
rect 13165 31838 13216 31840
rect 13250 31838 13289 31840
rect 13323 31838 13362 31840
rect 13396 31838 13435 31840
rect 13469 31838 13508 31840
rect 13165 31804 13202 31838
rect 13250 31806 13270 31838
rect 13323 31806 13338 31838
rect 13396 31806 13406 31838
rect 13469 31806 13474 31838
rect 13236 31804 13270 31806
rect 13304 31804 13338 31806
rect 13372 31804 13406 31806
rect 13440 31804 13474 31806
rect 13542 31838 13581 31840
rect 13615 31838 13654 31840
rect 13688 31838 13727 31840
rect 13761 31838 13800 31840
rect 13834 31838 13873 31840
rect 13907 31838 13946 31840
rect 13980 31838 14019 31840
rect 14053 31838 14092 31840
rect 14126 31838 14165 31840
rect 14199 31838 14238 31840
rect 14272 31838 14311 31840
rect 14345 31838 14384 31840
rect 13508 31804 13542 31806
rect 13576 31806 13581 31838
rect 13644 31806 13654 31838
rect 13712 31806 13727 31838
rect 13780 31806 13800 31838
rect 13848 31806 13873 31838
rect 13916 31806 13946 31838
rect 13576 31804 13610 31806
rect 13644 31804 13678 31806
rect 13712 31804 13746 31806
rect 13780 31804 13814 31806
rect 13848 31804 13882 31806
rect 13916 31804 13950 31806
rect 13984 31804 14018 31838
rect 14053 31806 14086 31838
rect 14126 31806 14154 31838
rect 14199 31806 14222 31838
rect 14272 31806 14290 31838
rect 14345 31806 14358 31838
rect 14418 31806 14429 31840
rect 14052 31804 14086 31806
rect 14120 31804 14154 31806
rect 14188 31804 14222 31806
rect 14256 31804 14290 31806
rect 14324 31804 14358 31806
rect 14392 31804 14429 31806
rect 13165 31769 14429 31804
rect 13165 31735 13202 31769
rect 13236 31767 13270 31769
rect 13304 31767 13338 31769
rect 13372 31767 13406 31769
rect 13440 31767 13474 31769
rect 13250 31735 13270 31767
rect 13323 31735 13338 31767
rect 13396 31735 13406 31767
rect 13469 31735 13474 31767
rect 13508 31767 13542 31769
rect 13165 31733 13216 31735
rect 13250 31733 13289 31735
rect 13323 31733 13362 31735
rect 13396 31733 13435 31735
rect 13469 31733 13508 31735
rect 13576 31767 13610 31769
rect 13644 31767 13678 31769
rect 13712 31767 13746 31769
rect 13780 31767 13814 31769
rect 13848 31767 13882 31769
rect 13916 31767 13950 31769
rect 13576 31735 13581 31767
rect 13644 31735 13654 31767
rect 13712 31735 13727 31767
rect 13780 31735 13800 31767
rect 13848 31735 13873 31767
rect 13916 31735 13946 31767
rect 13984 31735 14018 31769
rect 14052 31767 14086 31769
rect 14120 31767 14154 31769
rect 14188 31767 14222 31769
rect 14256 31767 14290 31769
rect 14324 31767 14358 31769
rect 14392 31767 14429 31769
rect 14053 31735 14086 31767
rect 14126 31735 14154 31767
rect 14199 31735 14222 31767
rect 14272 31735 14290 31767
rect 14345 31735 14358 31767
rect 13542 31733 13581 31735
rect 13615 31733 13654 31735
rect 13688 31733 13727 31735
rect 13761 31733 13800 31735
rect 13834 31733 13873 31735
rect 13907 31733 13946 31735
rect 13980 31733 14019 31735
rect 14053 31733 14092 31735
rect 14126 31733 14165 31735
rect 14199 31733 14238 31735
rect 14272 31733 14311 31735
rect 14345 31733 14384 31735
rect 14418 31733 14429 31767
rect 13165 31700 14429 31733
rect 13165 31666 13202 31700
rect 13236 31694 13270 31700
rect 13304 31694 13338 31700
rect 13372 31694 13406 31700
rect 13440 31694 13474 31700
rect 13250 31666 13270 31694
rect 13323 31666 13338 31694
rect 13396 31666 13406 31694
rect 13469 31666 13474 31694
rect 13508 31694 13542 31700
rect 13165 31660 13216 31666
rect 13250 31660 13289 31666
rect 13323 31660 13362 31666
rect 13396 31660 13435 31666
rect 13469 31660 13508 31666
rect 13576 31694 13610 31700
rect 13644 31694 13678 31700
rect 13712 31694 13746 31700
rect 13780 31694 13814 31700
rect 13848 31694 13882 31700
rect 13916 31694 13950 31700
rect 13576 31666 13581 31694
rect 13644 31666 13654 31694
rect 13712 31666 13727 31694
rect 13780 31666 13800 31694
rect 13848 31666 13873 31694
rect 13916 31666 13946 31694
rect 13984 31666 14018 31700
rect 14052 31694 14086 31700
rect 14120 31694 14154 31700
rect 14188 31694 14222 31700
rect 14256 31694 14290 31700
rect 14324 31694 14358 31700
rect 14392 31694 14429 31700
rect 14053 31666 14086 31694
rect 14126 31666 14154 31694
rect 14199 31666 14222 31694
rect 14272 31666 14290 31694
rect 14345 31666 14358 31694
rect 13542 31660 13581 31666
rect 13615 31660 13654 31666
rect 13688 31660 13727 31666
rect 13761 31660 13800 31666
rect 13834 31660 13873 31666
rect 13907 31660 13946 31666
rect 13980 31660 14019 31666
rect 14053 31660 14092 31666
rect 14126 31660 14165 31666
rect 14199 31660 14238 31666
rect 14272 31660 14311 31666
rect 14345 31660 14384 31666
rect 14418 31660 14429 31694
rect 13165 31631 14429 31660
rect 13165 31597 13202 31631
rect 13236 31621 13270 31631
rect 13304 31621 13338 31631
rect 13372 31621 13406 31631
rect 13440 31621 13474 31631
rect 13250 31597 13270 31621
rect 13323 31597 13338 31621
rect 13396 31597 13406 31621
rect 13469 31597 13474 31621
rect 13508 31621 13542 31631
rect 13165 31587 13216 31597
rect 13250 31587 13289 31597
rect 13323 31587 13362 31597
rect 13396 31587 13435 31597
rect 13469 31587 13508 31597
rect 13576 31621 13610 31631
rect 13644 31621 13678 31631
rect 13712 31621 13746 31631
rect 13780 31621 13814 31631
rect 13848 31621 13882 31631
rect 13916 31621 13950 31631
rect 13576 31597 13581 31621
rect 13644 31597 13654 31621
rect 13712 31597 13727 31621
rect 13780 31597 13800 31621
rect 13848 31597 13873 31621
rect 13916 31597 13946 31621
rect 13984 31597 14018 31631
rect 14052 31621 14086 31631
rect 14120 31621 14154 31631
rect 14188 31621 14222 31631
rect 14256 31621 14290 31631
rect 14324 31621 14358 31631
rect 14392 31621 14429 31631
rect 14053 31597 14086 31621
rect 14126 31597 14154 31621
rect 14199 31597 14222 31621
rect 14272 31597 14290 31621
rect 14345 31597 14358 31621
rect 13542 31587 13581 31597
rect 13615 31587 13654 31597
rect 13688 31587 13727 31597
rect 13761 31587 13800 31597
rect 13834 31587 13873 31597
rect 13907 31587 13946 31597
rect 13980 31587 14019 31597
rect 14053 31587 14092 31597
rect 14126 31587 14165 31597
rect 14199 31587 14238 31597
rect 14272 31587 14311 31597
rect 14345 31587 14384 31597
rect 14418 31587 14429 31621
rect 13165 31562 14429 31587
rect 13165 31528 13202 31562
rect 13236 31548 13270 31562
rect 13304 31548 13338 31562
rect 13372 31548 13406 31562
rect 13440 31548 13474 31562
rect 13250 31528 13270 31548
rect 13323 31528 13338 31548
rect 13396 31528 13406 31548
rect 13469 31528 13474 31548
rect 13508 31548 13542 31562
rect 13165 31514 13216 31528
rect 13250 31514 13289 31528
rect 13323 31514 13362 31528
rect 13396 31514 13435 31528
rect 13469 31514 13508 31528
rect 13576 31548 13610 31562
rect 13644 31548 13678 31562
rect 13712 31548 13746 31562
rect 13780 31548 13814 31562
rect 13848 31548 13882 31562
rect 13916 31548 13950 31562
rect 13576 31528 13581 31548
rect 13644 31528 13654 31548
rect 13712 31528 13727 31548
rect 13780 31528 13800 31548
rect 13848 31528 13873 31548
rect 13916 31528 13946 31548
rect 13984 31528 14018 31562
rect 14052 31548 14086 31562
rect 14120 31548 14154 31562
rect 14188 31548 14222 31562
rect 14256 31548 14290 31562
rect 14324 31548 14358 31562
rect 14392 31548 14429 31562
rect 14053 31528 14086 31548
rect 14126 31528 14154 31548
rect 14199 31528 14222 31548
rect 14272 31528 14290 31548
rect 14345 31528 14358 31548
rect 13542 31514 13581 31528
rect 13615 31514 13654 31528
rect 13688 31514 13727 31528
rect 13761 31514 13800 31528
rect 13834 31514 13873 31528
rect 13907 31514 13946 31528
rect 13980 31514 14019 31528
rect 14053 31514 14092 31528
rect 14126 31514 14165 31528
rect 14199 31514 14238 31528
rect 14272 31514 14311 31528
rect 14345 31514 14384 31528
rect 14418 31514 14429 31548
rect 13165 31493 14429 31514
rect 13165 31459 13202 31493
rect 13236 31475 13270 31493
rect 13304 31475 13338 31493
rect 13372 31475 13406 31493
rect 13440 31475 13474 31493
rect 13250 31459 13270 31475
rect 13323 31459 13338 31475
rect 13396 31459 13406 31475
rect 13469 31459 13474 31475
rect 13508 31475 13542 31493
rect 13165 31441 13216 31459
rect 13250 31441 13289 31459
rect 13323 31441 13362 31459
rect 13396 31441 13435 31459
rect 13469 31441 13508 31459
rect 13576 31475 13610 31493
rect 13644 31475 13678 31493
rect 13712 31475 13746 31493
rect 13780 31475 13814 31493
rect 13848 31475 13882 31493
rect 13916 31475 13950 31493
rect 13576 31459 13581 31475
rect 13644 31459 13654 31475
rect 13712 31459 13727 31475
rect 13780 31459 13800 31475
rect 13848 31459 13873 31475
rect 13916 31459 13946 31475
rect 13984 31459 14018 31493
rect 14052 31475 14086 31493
rect 14120 31475 14154 31493
rect 14188 31475 14222 31493
rect 14256 31475 14290 31493
rect 14324 31475 14358 31493
rect 14392 31475 14429 31493
rect 14053 31459 14086 31475
rect 14126 31459 14154 31475
rect 14199 31459 14222 31475
rect 14272 31459 14290 31475
rect 14345 31459 14358 31475
rect 13542 31441 13581 31459
rect 13615 31441 13654 31459
rect 13688 31441 13727 31459
rect 13761 31441 13800 31459
rect 13834 31441 13873 31459
rect 13907 31441 13946 31459
rect 13980 31441 14019 31459
rect 14053 31441 14092 31459
rect 14126 31441 14165 31459
rect 14199 31441 14238 31459
rect 14272 31441 14311 31459
rect 14345 31441 14384 31459
rect 14418 31441 14429 31475
rect 13165 31424 14429 31441
rect 13165 31390 13202 31424
rect 13236 31402 13270 31424
rect 13304 31402 13338 31424
rect 13372 31402 13406 31424
rect 13440 31402 13474 31424
rect 13250 31390 13270 31402
rect 13323 31390 13338 31402
rect 13396 31390 13406 31402
rect 13469 31390 13474 31402
rect 13508 31402 13542 31424
rect 13165 31368 13216 31390
rect 13250 31368 13289 31390
rect 13323 31368 13362 31390
rect 13396 31368 13435 31390
rect 13469 31368 13508 31390
rect 13576 31402 13610 31424
rect 13644 31402 13678 31424
rect 13712 31402 13746 31424
rect 13780 31402 13814 31424
rect 13848 31402 13882 31424
rect 13916 31402 13950 31424
rect 13576 31390 13581 31402
rect 13644 31390 13654 31402
rect 13712 31390 13727 31402
rect 13780 31390 13800 31402
rect 13848 31390 13873 31402
rect 13916 31390 13946 31402
rect 13984 31390 14018 31424
rect 14052 31402 14086 31424
rect 14120 31402 14154 31424
rect 14188 31402 14222 31424
rect 14256 31402 14290 31424
rect 14324 31402 14358 31424
rect 14392 31402 14429 31424
rect 14053 31390 14086 31402
rect 14126 31390 14154 31402
rect 14199 31390 14222 31402
rect 14272 31390 14290 31402
rect 14345 31390 14358 31402
rect 13542 31368 13581 31390
rect 13615 31368 13654 31390
rect 13688 31368 13727 31390
rect 13761 31368 13800 31390
rect 13834 31368 13873 31390
rect 13907 31368 13946 31390
rect 13980 31368 14019 31390
rect 14053 31368 14092 31390
rect 14126 31368 14165 31390
rect 14199 31368 14238 31390
rect 14272 31368 14311 31390
rect 14345 31368 14384 31390
rect 14418 31368 14429 31402
rect 13165 31355 14429 31368
rect 13165 31321 13202 31355
rect 13236 31329 13270 31355
rect 13304 31329 13338 31355
rect 13372 31329 13406 31355
rect 13440 31329 13474 31355
rect 13250 31321 13270 31329
rect 13323 31321 13338 31329
rect 13396 31321 13406 31329
rect 13469 31321 13474 31329
rect 13508 31329 13542 31355
rect 13165 31295 13216 31321
rect 13250 31295 13289 31321
rect 13323 31295 13362 31321
rect 13396 31295 13435 31321
rect 13469 31295 13508 31321
rect 13576 31329 13610 31355
rect 13644 31329 13678 31355
rect 13712 31329 13746 31355
rect 13780 31329 13814 31355
rect 13848 31329 13882 31355
rect 13916 31329 13950 31355
rect 13576 31321 13581 31329
rect 13644 31321 13654 31329
rect 13712 31321 13727 31329
rect 13780 31321 13800 31329
rect 13848 31321 13873 31329
rect 13916 31321 13946 31329
rect 13984 31321 14018 31355
rect 14052 31329 14086 31355
rect 14120 31329 14154 31355
rect 14188 31329 14222 31355
rect 14256 31329 14290 31355
rect 14324 31329 14358 31355
rect 14392 31329 14429 31355
rect 14053 31321 14086 31329
rect 14126 31321 14154 31329
rect 14199 31321 14222 31329
rect 14272 31321 14290 31329
rect 14345 31321 14358 31329
rect 13542 31295 13581 31321
rect 13615 31295 13654 31321
rect 13688 31295 13727 31321
rect 13761 31295 13800 31321
rect 13834 31295 13873 31321
rect 13907 31295 13946 31321
rect 13980 31295 14019 31321
rect 14053 31295 14092 31321
rect 14126 31295 14165 31321
rect 14199 31295 14238 31321
rect 14272 31295 14311 31321
rect 14345 31295 14384 31321
rect 14418 31295 14429 31329
rect 13165 31286 14429 31295
rect 13165 31252 13202 31286
rect 13236 31256 13270 31286
rect 13304 31256 13338 31286
rect 13372 31256 13406 31286
rect 13440 31256 13474 31286
rect 13250 31252 13270 31256
rect 13323 31252 13338 31256
rect 13396 31252 13406 31256
rect 13469 31252 13474 31256
rect 13508 31256 13542 31286
rect 13165 31222 13216 31252
rect 13250 31222 13289 31252
rect 13323 31222 13362 31252
rect 13396 31222 13435 31252
rect 13469 31222 13508 31252
rect 13576 31256 13610 31286
rect 13644 31256 13678 31286
rect 13712 31256 13746 31286
rect 13780 31256 13814 31286
rect 13848 31256 13882 31286
rect 13916 31256 13950 31286
rect 13576 31252 13581 31256
rect 13644 31252 13654 31256
rect 13712 31252 13727 31256
rect 13780 31252 13800 31256
rect 13848 31252 13873 31256
rect 13916 31252 13946 31256
rect 13984 31252 14018 31286
rect 14052 31256 14086 31286
rect 14120 31256 14154 31286
rect 14188 31256 14222 31286
rect 14256 31256 14290 31286
rect 14324 31256 14358 31286
rect 14392 31256 14429 31286
rect 14053 31252 14086 31256
rect 14126 31252 14154 31256
rect 14199 31252 14222 31256
rect 14272 31252 14290 31256
rect 14345 31252 14358 31256
rect 13542 31222 13581 31252
rect 13615 31222 13654 31252
rect 13688 31222 13727 31252
rect 13761 31222 13800 31252
rect 13834 31222 13873 31252
rect 13907 31222 13946 31252
rect 13980 31222 14019 31252
rect 14053 31222 14092 31252
rect 14126 31222 14165 31252
rect 14199 31222 14238 31252
rect 14272 31222 14311 31252
rect 14345 31222 14384 31252
rect 14418 31222 14429 31256
rect 13165 31217 14429 31222
rect 13165 31183 13202 31217
rect 13236 31183 13270 31217
rect 13304 31183 13338 31217
rect 13372 31183 13406 31217
rect 13440 31183 13474 31217
rect 13508 31183 13542 31217
rect 13576 31183 13610 31217
rect 13644 31183 13678 31217
rect 13712 31183 13746 31217
rect 13780 31183 13814 31217
rect 13848 31183 13882 31217
rect 13916 31183 13950 31217
rect 13984 31183 14018 31217
rect 14052 31183 14086 31217
rect 14120 31183 14154 31217
rect 14188 31183 14222 31217
rect 14256 31183 14290 31217
rect 14324 31183 14358 31217
rect 14392 31183 14429 31217
rect 13165 31149 13216 31183
rect 13250 31149 13289 31183
rect 13323 31149 13362 31183
rect 13396 31149 13435 31183
rect 13469 31149 13508 31183
rect 13542 31149 13581 31183
rect 13615 31149 13654 31183
rect 13688 31149 13727 31183
rect 13761 31149 13800 31183
rect 13834 31149 13873 31183
rect 13907 31149 13946 31183
rect 13980 31149 14019 31183
rect 14053 31149 14092 31183
rect 14126 31149 14165 31183
rect 14199 31149 14238 31183
rect 14272 31149 14311 31183
rect 14345 31149 14384 31183
rect 14418 31149 14429 31183
rect 13011 30995 14268 30996
rect 13011 30991 13078 30995
rect 13011 30957 13051 30991
rect 14200 30961 14268 30995
rect 13011 30927 13078 30957
rect 13011 30863 13077 30927
rect 14199 30923 14268 30961
rect 14199 30919 14233 30923
rect 14199 30893 14230 30919
rect 14131 30885 14230 30893
rect 14267 30889 14268 30923
rect 14264 30885 14268 30889
rect 14131 30863 14268 30885
rect 13011 30829 13051 30863
rect 14136 30856 14268 30863
rect 14136 30829 14165 30856
rect 13011 30825 13077 30829
rect 14131 30825 14165 30829
rect 13011 30824 14165 30825
rect 14096 30791 14165 30824
rect 14096 30788 14102 30791
rect 14136 30788 14165 30791
rect 9877 30664 13943 30670
rect 9877 30636 10246 30664
rect 10280 30636 10320 30664
rect 10354 30636 10394 30664
rect 10428 30636 10467 30664
rect 9877 30602 9913 30636
rect 9947 30602 9982 30636
rect 10016 30602 10051 30636
rect 10085 30602 10120 30636
rect 10154 30602 10189 30636
rect 10223 30630 10246 30636
rect 10292 30630 10320 30636
rect 10361 30630 10394 30636
rect 10223 30602 10258 30630
rect 10292 30602 10327 30630
rect 10361 30602 10396 30630
rect 10430 30602 10465 30636
rect 10501 30630 10540 30664
rect 10574 30635 10613 30664
rect 10647 30635 10686 30664
rect 10720 30635 10759 30664
rect 10793 30635 10832 30664
rect 10866 30635 10905 30664
rect 10939 30635 10978 30664
rect 11012 30635 11051 30664
rect 11085 30635 11124 30664
rect 11158 30635 11197 30664
rect 11231 30635 11270 30664
rect 11304 30635 11343 30664
rect 11377 30635 11416 30664
rect 11450 30635 11489 30664
rect 11523 30635 11562 30664
rect 11596 30635 11635 30664
rect 11669 30635 11708 30664
rect 11742 30635 11781 30664
rect 11815 30635 11854 30664
rect 11888 30635 11927 30664
rect 11961 30635 12000 30664
rect 12034 30635 12073 30664
rect 10574 30630 10610 30635
rect 10647 30630 10679 30635
rect 10720 30630 10747 30635
rect 10793 30630 10815 30635
rect 10866 30630 10883 30635
rect 10939 30630 10951 30635
rect 11012 30630 11019 30635
rect 11085 30630 11087 30635
rect 10499 30602 10610 30630
rect 9877 30601 10610 30602
rect 10644 30601 10679 30630
rect 10713 30601 10747 30630
rect 10781 30601 10815 30630
rect 10849 30601 10883 30630
rect 10917 30601 10951 30630
rect 10985 30601 11019 30630
rect 11053 30601 11087 30630
rect 11121 30630 11124 30635
rect 11189 30630 11197 30635
rect 11257 30630 11270 30635
rect 11325 30630 11343 30635
rect 11393 30630 11416 30635
rect 11461 30630 11489 30635
rect 11529 30630 11562 30635
rect 11121 30601 11155 30630
rect 11189 30601 11223 30630
rect 11257 30601 11291 30630
rect 11325 30601 11359 30630
rect 11393 30601 11427 30630
rect 11461 30601 11495 30630
rect 11529 30601 11563 30630
rect 11597 30601 11631 30635
rect 11669 30630 11699 30635
rect 11742 30630 11767 30635
rect 11815 30630 11835 30635
rect 11888 30630 11903 30635
rect 11961 30630 11971 30635
rect 12034 30630 12039 30635
rect 11665 30601 11699 30630
rect 11733 30601 11767 30630
rect 11801 30601 11835 30630
rect 11869 30601 11903 30630
rect 11937 30601 11971 30630
rect 12005 30601 12039 30630
rect 12107 30635 12146 30664
rect 12180 30635 12219 30664
rect 12253 30635 12292 30664
rect 12326 30635 12365 30664
rect 12399 30635 12438 30664
rect 12472 30635 12511 30664
rect 12545 30635 12584 30664
rect 12618 30635 12657 30664
rect 12691 30635 12730 30664
rect 12764 30635 12803 30664
rect 12837 30635 12876 30664
rect 12910 30635 12949 30664
rect 12983 30635 13022 30664
rect 13056 30635 13095 30664
rect 13129 30635 13168 30664
rect 13202 30635 13241 30664
rect 13275 30635 13314 30664
rect 13348 30635 13387 30664
rect 13421 30635 13460 30664
rect 13494 30635 13533 30664
rect 13567 30635 13606 30664
rect 13640 30635 13679 30664
rect 13713 30635 13752 30664
rect 13786 30635 13825 30664
rect 13859 30635 13898 30664
rect 12073 30601 12107 30630
rect 12141 30630 12146 30635
rect 12209 30630 12219 30635
rect 12277 30630 12292 30635
rect 12345 30630 12365 30635
rect 12413 30630 12438 30635
rect 12481 30630 12511 30635
rect 12141 30601 12175 30630
rect 12209 30601 12243 30630
rect 12277 30601 12311 30630
rect 12345 30601 12379 30630
rect 12413 30601 12447 30630
rect 12481 30601 12515 30630
rect 12549 30601 12583 30635
rect 12618 30630 12651 30635
rect 12691 30630 12719 30635
rect 12764 30630 12787 30635
rect 12837 30630 12855 30635
rect 12910 30630 12923 30635
rect 12983 30630 12991 30635
rect 13056 30630 13059 30635
rect 12617 30601 12651 30630
rect 12685 30601 12719 30630
rect 12753 30601 12787 30630
rect 12821 30601 12855 30630
rect 12889 30601 12923 30630
rect 12957 30601 12991 30630
rect 13025 30601 13059 30630
rect 13093 30630 13095 30635
rect 13161 30630 13168 30635
rect 13229 30630 13241 30635
rect 13297 30630 13314 30635
rect 13365 30630 13387 30635
rect 13433 30630 13460 30635
rect 13501 30630 13533 30635
rect 13093 30601 13127 30630
rect 13161 30601 13195 30630
rect 13229 30601 13263 30630
rect 13297 30601 13331 30630
rect 13365 30601 13399 30630
rect 13433 30601 13467 30630
rect 13501 30601 13535 30630
rect 13569 30601 13603 30635
rect 13640 30630 13671 30635
rect 13713 30630 13739 30635
rect 13786 30630 13807 30635
rect 13859 30630 13875 30635
rect 13932 30630 13943 30664
rect 13637 30601 13671 30630
rect 13705 30601 13739 30630
rect 13773 30601 13807 30630
rect 13841 30601 13875 30630
rect 13909 30601 13943 30630
rect 9877 30568 13943 30601
rect 9877 30534 9913 30568
rect 9947 30534 9982 30568
rect 10016 30534 10051 30568
rect 10085 30534 10120 30568
rect 10154 30534 10189 30568
rect 10223 30557 10258 30568
rect 10292 30557 10327 30568
rect 10361 30557 10396 30568
rect 10223 30534 10246 30557
rect 10292 30534 10320 30557
rect 10361 30534 10394 30557
rect 10430 30534 10465 30568
rect 10499 30560 13943 30568
rect 10499 30557 10610 30560
rect 10644 30557 10679 30560
rect 10713 30557 10747 30560
rect 10781 30557 10815 30560
rect 10849 30557 10883 30560
rect 10917 30557 10951 30560
rect 10985 30557 11019 30560
rect 11053 30557 11087 30560
rect 9877 30523 10246 30534
rect 10280 30523 10320 30534
rect 10354 30523 10394 30534
rect 10428 30523 10467 30534
rect 10501 30523 10540 30557
rect 10574 30526 10610 30557
rect 10647 30526 10679 30557
rect 10720 30526 10747 30557
rect 10793 30526 10815 30557
rect 10866 30526 10883 30557
rect 10939 30526 10951 30557
rect 11012 30526 11019 30557
rect 11085 30526 11087 30557
rect 11121 30557 11155 30560
rect 11189 30557 11223 30560
rect 11257 30557 11291 30560
rect 11325 30557 11359 30560
rect 11393 30557 11427 30560
rect 11461 30557 11495 30560
rect 11529 30557 11563 30560
rect 11121 30526 11124 30557
rect 11189 30526 11197 30557
rect 11257 30526 11270 30557
rect 11325 30526 11343 30557
rect 11393 30526 11416 30557
rect 11461 30526 11489 30557
rect 11529 30526 11562 30557
rect 11597 30526 11631 30560
rect 11665 30557 11699 30560
rect 11733 30557 11767 30560
rect 11801 30557 11835 30560
rect 11869 30557 11903 30560
rect 11937 30557 11971 30560
rect 12005 30557 12039 30560
rect 11669 30526 11699 30557
rect 11742 30526 11767 30557
rect 11815 30526 11835 30557
rect 11888 30526 11903 30557
rect 11961 30526 11971 30557
rect 12034 30526 12039 30557
rect 12073 30557 12107 30560
rect 10574 30523 10613 30526
rect 10647 30523 10686 30526
rect 10720 30523 10759 30526
rect 10793 30523 10832 30526
rect 10866 30523 10905 30526
rect 10939 30523 10978 30526
rect 11012 30523 11051 30526
rect 11085 30523 11124 30526
rect 11158 30523 11197 30526
rect 11231 30523 11270 30526
rect 11304 30523 11343 30526
rect 11377 30523 11416 30526
rect 11450 30523 11489 30526
rect 11523 30523 11562 30526
rect 11596 30523 11635 30526
rect 11669 30523 11708 30526
rect 11742 30523 11781 30526
rect 11815 30523 11854 30526
rect 11888 30523 11927 30526
rect 11961 30523 12000 30526
rect 12034 30523 12073 30526
rect 12141 30557 12175 30560
rect 12209 30557 12243 30560
rect 12277 30557 12311 30560
rect 12345 30557 12379 30560
rect 12413 30557 12447 30560
rect 12481 30557 12515 30560
rect 12141 30526 12146 30557
rect 12209 30526 12219 30557
rect 12277 30526 12292 30557
rect 12345 30526 12365 30557
rect 12413 30526 12438 30557
rect 12481 30526 12511 30557
rect 12549 30526 12583 30560
rect 12617 30557 12651 30560
rect 12685 30557 12719 30560
rect 12753 30557 12787 30560
rect 12821 30557 12855 30560
rect 12889 30557 12923 30560
rect 12957 30557 12991 30560
rect 13025 30557 13059 30560
rect 12618 30526 12651 30557
rect 12691 30526 12719 30557
rect 12764 30526 12787 30557
rect 12837 30526 12855 30557
rect 12910 30526 12923 30557
rect 12983 30526 12991 30557
rect 13056 30526 13059 30557
rect 13093 30557 13127 30560
rect 13161 30557 13195 30560
rect 13229 30557 13263 30560
rect 13297 30557 13331 30560
rect 13365 30557 13399 30560
rect 13433 30557 13467 30560
rect 13501 30557 13535 30560
rect 13093 30526 13095 30557
rect 13161 30526 13168 30557
rect 13229 30526 13241 30557
rect 13297 30526 13314 30557
rect 13365 30526 13387 30557
rect 13433 30526 13460 30557
rect 13501 30526 13533 30557
rect 13569 30526 13603 30560
rect 13637 30557 13671 30560
rect 13705 30557 13739 30560
rect 13773 30557 13807 30560
rect 13841 30557 13875 30560
rect 13909 30557 13943 30560
rect 13640 30526 13671 30557
rect 13713 30526 13739 30557
rect 13786 30526 13807 30557
rect 13859 30526 13875 30557
rect 12107 30523 12146 30526
rect 12180 30523 12219 30526
rect 12253 30523 12292 30526
rect 12326 30523 12365 30526
rect 12399 30523 12438 30526
rect 12472 30523 12511 30526
rect 12545 30523 12584 30526
rect 12618 30523 12657 30526
rect 12691 30523 12730 30526
rect 12764 30523 12803 30526
rect 12837 30523 12876 30526
rect 12910 30523 12949 30526
rect 12983 30523 13022 30526
rect 13056 30523 13095 30526
rect 13129 30523 13168 30526
rect 13202 30523 13241 30526
rect 13275 30523 13314 30526
rect 13348 30523 13387 30526
rect 13421 30523 13460 30526
rect 13494 30523 13533 30526
rect 13567 30523 13606 30526
rect 13640 30523 13679 30526
rect 13713 30523 13752 30526
rect 13786 30523 13825 30526
rect 13859 30523 13898 30526
rect 13932 30523 13943 30557
rect 9877 30500 13943 30523
rect 9877 30466 9913 30500
rect 9947 30466 9982 30500
rect 10016 30466 10051 30500
rect 10085 30466 10120 30500
rect 10154 30466 10189 30500
rect 10223 30466 10258 30500
rect 10292 30466 10327 30500
rect 10361 30466 10396 30500
rect 10430 30466 10465 30500
rect 10499 30485 13943 30500
rect 10499 30466 10610 30485
rect 9877 30451 10610 30466
rect 10644 30451 10679 30485
rect 10713 30451 10747 30485
rect 10781 30451 10815 30485
rect 10849 30451 10883 30485
rect 10917 30451 10951 30485
rect 10985 30451 11019 30485
rect 11053 30451 11087 30485
rect 11121 30451 11155 30485
rect 11189 30451 11223 30485
rect 11257 30451 11291 30485
rect 11325 30451 11359 30485
rect 11393 30451 11427 30485
rect 11461 30451 11495 30485
rect 11529 30451 11563 30485
rect 11597 30451 11631 30485
rect 11665 30451 11699 30485
rect 11733 30451 11767 30485
rect 11801 30451 11835 30485
rect 11869 30451 11903 30485
rect 11937 30451 11971 30485
rect 12005 30451 12039 30485
rect 12073 30451 12107 30485
rect 12141 30451 12175 30485
rect 12209 30451 12243 30485
rect 12277 30451 12311 30485
rect 12345 30451 12379 30485
rect 12413 30451 12447 30485
rect 12481 30451 12515 30485
rect 12549 30451 12583 30485
rect 12617 30451 12651 30485
rect 12685 30451 12719 30485
rect 12753 30451 12787 30485
rect 12821 30451 12855 30485
rect 12889 30451 12923 30485
rect 12957 30451 12991 30485
rect 13025 30451 13059 30485
rect 13093 30451 13127 30485
rect 13161 30451 13195 30485
rect 13229 30451 13263 30485
rect 13297 30451 13331 30485
rect 13365 30451 13399 30485
rect 13433 30451 13467 30485
rect 13501 30451 13535 30485
rect 13569 30451 13603 30485
rect 13637 30451 13671 30485
rect 13705 30451 13739 30485
rect 13773 30451 13807 30485
rect 13841 30451 13875 30485
rect 13909 30451 13943 30485
rect 9877 30450 13943 30451
rect 9877 30432 10246 30450
rect 10280 30432 10320 30450
rect 10354 30432 10394 30450
rect 10428 30432 10467 30450
rect 9877 30398 9913 30432
rect 9947 30398 9982 30432
rect 10016 30398 10051 30432
rect 10085 30398 10120 30432
rect 10154 30398 10189 30432
rect 10223 30416 10246 30432
rect 10292 30416 10320 30432
rect 10361 30416 10394 30432
rect 10223 30398 10258 30416
rect 10292 30398 10327 30416
rect 10361 30398 10396 30416
rect 10430 30398 10465 30432
rect 10501 30416 10540 30450
rect 10574 30416 10613 30450
rect 10647 30416 10686 30450
rect 10720 30416 10759 30450
rect 10793 30416 10832 30450
rect 10866 30416 10905 30450
rect 10939 30416 10978 30450
rect 11012 30416 11051 30450
rect 11085 30416 11124 30450
rect 11158 30416 11197 30450
rect 11231 30416 11270 30450
rect 11304 30416 11343 30450
rect 11377 30416 11416 30450
rect 11450 30416 11489 30450
rect 11523 30416 11562 30450
rect 11596 30416 11635 30450
rect 11669 30416 11708 30450
rect 11742 30416 11781 30450
rect 11815 30416 11854 30450
rect 11888 30416 11927 30450
rect 11961 30416 12000 30450
rect 12034 30416 12073 30450
rect 12107 30416 12146 30450
rect 12180 30416 12219 30450
rect 12253 30416 12292 30450
rect 12326 30416 12365 30450
rect 12399 30416 12438 30450
rect 12472 30416 12511 30450
rect 12545 30416 12584 30450
rect 12618 30416 12657 30450
rect 12691 30416 12730 30450
rect 12764 30416 12803 30450
rect 12837 30416 12876 30450
rect 12910 30416 12949 30450
rect 12983 30416 13022 30450
rect 13056 30416 13095 30450
rect 13129 30416 13168 30450
rect 13202 30416 13241 30450
rect 13275 30416 13314 30450
rect 13348 30416 13387 30450
rect 13421 30416 13460 30450
rect 13494 30416 13533 30450
rect 13567 30416 13606 30450
rect 13640 30416 13679 30450
rect 13713 30416 13752 30450
rect 13786 30416 13825 30450
rect 13859 30416 13898 30450
rect 13932 30416 13943 30450
rect 10499 30398 10535 30416
rect 9877 30364 10535 30398
rect 9877 30330 9913 30364
rect 9947 30330 9982 30364
rect 10016 30330 10051 30364
rect 10085 30330 10120 30364
rect 10154 30330 10189 30364
rect 10223 30330 10258 30364
rect 10292 30330 10327 30364
rect 10361 30330 10396 30364
rect 10430 30330 10465 30364
rect 10499 30330 10535 30364
rect 9877 30296 10535 30330
rect 9877 30262 9913 30296
rect 9947 30262 9982 30296
rect 10016 30262 10051 30296
rect 10085 30262 10120 30296
rect 10154 30262 10189 30296
rect 10223 30262 10258 30296
rect 10292 30262 10327 30296
rect 10361 30262 10396 30296
rect 10430 30262 10465 30296
rect 10499 30262 10535 30296
rect 9877 30228 10535 30262
rect 9877 30194 9913 30228
rect 9947 30194 9982 30228
rect 10016 30194 10051 30228
rect 10085 30194 10120 30228
rect 10154 30194 10189 30228
rect 10223 30194 10258 30228
rect 10292 30194 10327 30228
rect 10361 30194 10396 30228
rect 10430 30194 10465 30228
rect 10499 30194 10535 30228
rect 9877 30160 10535 30194
rect 9877 30126 9913 30160
rect 9947 30126 9982 30160
rect 10016 30126 10051 30160
rect 10085 30126 10120 30160
rect 10154 30126 10189 30160
rect 10223 30126 10258 30160
rect 10292 30126 10327 30160
rect 10361 30126 10396 30160
rect 10430 30126 10465 30160
rect 10499 30126 10535 30160
rect 9877 30092 10535 30126
rect 9877 30058 9913 30092
rect 9947 30058 9982 30092
rect 10016 30058 10051 30092
rect 10085 30058 10120 30092
rect 10154 30058 10189 30092
rect 10223 30058 10258 30092
rect 10292 30058 10327 30092
rect 10361 30058 10396 30092
rect 10430 30058 10465 30092
rect 10499 30058 10535 30092
rect 9877 30024 10535 30058
rect 9877 29990 9913 30024
rect 9947 29990 9982 30024
rect 10016 29990 10051 30024
rect 10085 29990 10120 30024
rect 10154 29990 10189 30024
rect 10223 29990 10258 30024
rect 10292 29990 10327 30024
rect 10361 29990 10396 30024
rect 10430 29990 10465 30024
rect 10499 29990 10535 30024
rect 9877 29956 10535 29990
rect 9877 29922 9913 29956
rect 9947 29922 9982 29956
rect 10016 29922 10051 29956
rect 10085 29922 10120 29956
rect 10154 29922 10189 29956
rect 10223 29922 10258 29956
rect 10292 29922 10327 29956
rect 10361 29922 10396 29956
rect 10430 29922 10465 29956
rect 10499 29922 10535 29956
rect 9877 29888 10535 29922
rect 9877 29854 9913 29888
rect 9947 29854 9982 29888
rect 10016 29854 10051 29888
rect 10085 29854 10120 29888
rect 10154 29854 10189 29888
rect 10223 29854 10258 29888
rect 10292 29854 10327 29888
rect 10361 29854 10396 29888
rect 10430 29854 10465 29888
rect 10499 29854 10535 29888
rect 9877 29820 10535 29854
rect 9877 29786 9913 29820
rect 9947 29786 9982 29820
rect 10016 29786 10051 29820
rect 10085 29786 10120 29820
rect 10154 29786 10189 29820
rect 10223 29786 10258 29820
rect 10292 29786 10327 29820
rect 10361 29786 10396 29820
rect 10430 29786 10465 29820
rect 10499 29786 10535 29820
rect 9877 29752 10535 29786
rect 9877 29718 9913 29752
rect 9947 29718 9982 29752
rect 10016 29718 10051 29752
rect 10085 29718 10120 29752
rect 10154 29718 10189 29752
rect 10223 29718 10258 29752
rect 10292 29718 10327 29752
rect 10361 29718 10396 29752
rect 10430 29718 10465 29752
rect 10499 29718 10535 29752
rect 9877 29684 10535 29718
rect 9877 29650 9913 29684
rect 9947 29650 9982 29684
rect 10016 29650 10051 29684
rect 10085 29650 10120 29684
rect 10154 29650 10189 29684
rect 10223 29650 10258 29684
rect 10292 29650 10327 29684
rect 10361 29650 10396 29684
rect 10430 29650 10465 29684
rect 10499 29650 10535 29684
rect 9877 29616 10535 29650
rect 9877 29582 9913 29616
rect 9947 29582 9982 29616
rect 10016 29582 10051 29616
rect 10085 29582 10120 29616
rect 10154 29582 10189 29616
rect 10223 29582 10258 29616
rect 10292 29582 10327 29616
rect 10361 29582 10396 29616
rect 10430 29582 10465 29616
rect 10499 29582 10535 29616
rect 9877 29548 10535 29582
rect 9877 29514 9913 29548
rect 9947 29514 9982 29548
rect 10016 29514 10051 29548
rect 10085 29514 10120 29548
rect 10154 29514 10189 29548
rect 10223 29514 10258 29548
rect 10292 29514 10327 29548
rect 10361 29514 10396 29548
rect 10430 29514 10465 29548
rect 10499 29514 10535 29548
rect 9877 29480 10535 29514
rect 9877 29446 9913 29480
rect 9947 29446 9982 29480
rect 10016 29446 10051 29480
rect 10085 29446 10120 29480
rect 10154 29446 10189 29480
rect 10223 29446 10258 29480
rect 10292 29446 10327 29480
rect 10361 29446 10396 29480
rect 10430 29446 10465 29480
rect 10499 29446 10535 29480
rect 9877 29412 10535 29446
rect 9877 29378 9913 29412
rect 9947 29378 9982 29412
rect 10016 29378 10051 29412
rect 10085 29378 10120 29412
rect 10154 29378 10189 29412
rect 10223 29378 10258 29412
rect 10292 29378 10327 29412
rect 10361 29378 10396 29412
rect 10430 29378 10465 29412
rect 10499 29378 10535 29412
rect 9877 29344 10535 29378
rect 9877 29310 9913 29344
rect 9947 29310 9982 29344
rect 10016 29310 10051 29344
rect 10085 29310 10120 29344
rect 10154 29310 10189 29344
rect 10223 29310 10258 29344
rect 10292 29310 10327 29344
rect 10361 29310 10396 29344
rect 10430 29310 10465 29344
rect 10499 29310 10535 29344
rect 9877 29276 10535 29310
rect 9877 29242 9913 29276
rect 9947 29242 9982 29276
rect 10016 29242 10051 29276
rect 10085 29242 10120 29276
rect 10154 29242 10189 29276
rect 10223 29242 10258 29276
rect 10292 29242 10327 29276
rect 10361 29242 10396 29276
rect 10430 29242 10465 29276
rect 10499 29242 10535 29276
rect 9877 29208 10535 29242
rect 9877 29174 9913 29208
rect 9947 29174 9982 29208
rect 10016 29174 10051 29208
rect 10085 29174 10120 29208
rect 10154 29174 10189 29208
rect 10223 29175 10258 29208
rect 10223 29174 10248 29175
rect 10292 29174 10327 29208
rect 10361 29175 10396 29208
rect 10430 29175 10465 29208
rect 10499 29175 10535 29208
rect 13703 30401 13943 30416
rect 13703 30374 13738 30401
rect 13908 30374 13943 30401
rect 13703 30340 13705 30374
rect 13908 30340 13909 30374
rect 13943 30340 13944 30374
rect 13703 30301 13738 30340
rect 13908 30301 13944 30340
rect 13703 30267 13705 30301
rect 13703 30228 13738 30267
rect 13908 30267 13909 30301
rect 13943 30267 13944 30301
rect 13908 30228 13944 30267
rect 13703 30194 13705 30228
rect 13703 30155 13738 30194
rect 13908 30194 13909 30228
rect 13943 30194 13944 30228
rect 13908 30155 13944 30194
rect 13703 30121 13705 30155
rect 13703 30082 13738 30121
rect 13908 30121 13909 30155
rect 13943 30121 13944 30155
rect 13908 30082 13944 30121
rect 13703 30048 13705 30082
rect 13703 30009 13738 30048
rect 13908 30048 13909 30082
rect 13943 30048 13944 30082
rect 13908 30009 13944 30048
rect 13703 29975 13705 30009
rect 13703 29936 13738 29975
rect 13908 29975 13909 30009
rect 13943 29975 13944 30009
rect 13908 29936 13944 29975
rect 13703 29902 13705 29936
rect 13703 29863 13738 29902
rect 13908 29902 13909 29936
rect 13943 29902 13944 29936
rect 13908 29863 13944 29902
rect 13703 29829 13705 29863
rect 13703 29790 13738 29829
rect 13908 29829 13909 29863
rect 13943 29829 13944 29863
rect 13908 29790 13944 29829
rect 13703 29756 13705 29790
rect 13703 29717 13738 29756
rect 13908 29756 13909 29790
rect 13943 29756 13944 29790
rect 13908 29717 13944 29756
rect 13703 29683 13705 29717
rect 13703 29644 13738 29683
rect 13908 29683 13909 29717
rect 13943 29683 13944 29717
rect 13908 29644 13944 29683
rect 13703 29610 13705 29644
rect 13703 29571 13738 29610
rect 13908 29610 13909 29644
rect 13943 29610 13944 29644
rect 13908 29572 13944 29610
rect 13703 29537 13705 29571
rect 13703 29498 13738 29537
rect 13908 29538 13909 29572
rect 13943 29538 13944 29572
rect 13908 29500 13944 29538
rect 13703 29464 13705 29498
rect 13703 29425 13738 29464
rect 13908 29466 13909 29500
rect 13943 29466 13944 29500
rect 13908 29428 13944 29466
rect 13703 29391 13705 29425
rect 13703 29352 13738 29391
rect 13908 29394 13909 29428
rect 13943 29394 13944 29428
rect 13908 29356 13944 29394
rect 13703 29318 13705 29352
rect 13703 29279 13738 29318
rect 13908 29322 13909 29356
rect 13943 29322 13944 29356
rect 13908 29284 13944 29322
rect 13703 29245 13705 29279
rect 13703 29206 13738 29245
rect 13908 29250 13909 29284
rect 13943 29250 13944 29284
rect 13908 29212 13944 29250
rect 10365 29174 10396 29175
rect 10448 29174 10465 29175
rect 9877 29141 10248 29174
rect 10282 29141 10331 29174
rect 10365 29141 10414 29174
rect 10448 29141 10497 29174
rect 10531 29141 10580 29175
rect 10614 29141 10615 29175
rect 9877 29140 10615 29141
rect 9877 29106 9913 29140
rect 9947 29106 9982 29140
rect 10016 29106 10051 29140
rect 10085 29106 10120 29140
rect 10154 29106 10189 29140
rect 10223 29106 10258 29140
rect 10292 29106 10327 29140
rect 10361 29106 10396 29140
rect 10430 29106 10465 29140
rect 10499 29106 10615 29140
rect 9877 29102 10615 29106
rect 9877 29072 10248 29102
rect 10282 29072 10331 29102
rect 10365 29072 10414 29102
rect 10448 29072 10497 29102
rect 9877 29038 9913 29072
rect 9947 29038 9982 29072
rect 10016 29038 10051 29072
rect 10085 29038 10120 29072
rect 10154 29038 10189 29072
rect 10223 29068 10248 29072
rect 10223 29038 10258 29068
rect 10292 29038 10327 29072
rect 10365 29068 10396 29072
rect 10448 29068 10465 29072
rect 10531 29068 10580 29102
rect 10614 29068 10615 29102
rect 10361 29038 10396 29068
rect 10430 29038 10465 29068
rect 10499 29038 10615 29068
rect 9877 29029 10615 29038
rect 9877 29004 10248 29029
rect 10282 29004 10331 29029
rect 10365 29004 10414 29029
rect 10448 29004 10497 29029
rect 9877 28970 9913 29004
rect 9947 28970 9982 29004
rect 10016 28970 10051 29004
rect 10085 28970 10120 29004
rect 10154 28970 10189 29004
rect 10223 28995 10248 29004
rect 10223 28970 10258 28995
rect 10292 28970 10327 29004
rect 10365 28995 10396 29004
rect 10448 28995 10465 29004
rect 10531 28995 10580 29029
rect 10614 28995 10615 29029
rect 10361 28970 10396 28995
rect 10430 28970 10465 28995
rect 10499 28970 10615 28995
rect 9877 28956 10615 28970
rect 9877 28936 10248 28956
rect 10282 28936 10331 28956
rect 10365 28936 10414 28956
rect 10448 28936 10497 28956
rect 9877 28902 9913 28936
rect 9947 28902 9982 28936
rect 10016 28902 10051 28936
rect 10085 28902 10120 28936
rect 10154 28902 10189 28936
rect 10223 28922 10248 28936
rect 10223 28902 10258 28922
rect 10292 28902 10327 28936
rect 10365 28922 10396 28936
rect 10448 28922 10465 28936
rect 10531 28922 10580 28956
rect 10614 28922 10615 28956
rect 10361 28902 10396 28922
rect 10430 28902 10465 28922
rect 10499 28902 10615 28922
rect 9877 28883 10615 28902
rect 9877 28868 10248 28883
rect 10282 28868 10331 28883
rect 10365 28868 10414 28883
rect 10448 28868 10497 28883
rect 9877 28834 9913 28868
rect 9947 28834 9982 28868
rect 10016 28834 10051 28868
rect 10085 28834 10120 28868
rect 10154 28834 10189 28868
rect 10223 28849 10248 28868
rect 10223 28834 10258 28849
rect 10292 28834 10327 28868
rect 10365 28849 10396 28868
rect 10448 28849 10465 28868
rect 10531 28849 10580 28883
rect 10614 28849 10615 28883
rect 10361 28834 10396 28849
rect 10430 28834 10465 28849
rect 10499 28834 10615 28849
rect 9877 28810 10615 28834
rect 9877 28800 10248 28810
rect 10282 28800 10331 28810
rect 10365 28800 10414 28810
rect 10448 28800 10497 28810
rect 9877 28766 9913 28800
rect 9947 28766 9982 28800
rect 10016 28766 10051 28800
rect 10085 28766 10120 28800
rect 10154 28766 10189 28800
rect 10223 28776 10248 28800
rect 10223 28766 10258 28776
rect 10292 28766 10327 28800
rect 10365 28776 10396 28800
rect 10448 28776 10465 28800
rect 10531 28776 10580 28810
rect 10614 28776 10615 28810
rect 10361 28766 10396 28776
rect 10430 28766 10465 28776
rect 10499 28766 10615 28776
rect 9877 28737 10615 28766
rect 9877 28732 10248 28737
rect 10282 28732 10331 28737
rect 10365 28732 10414 28737
rect 10448 28732 10497 28737
rect 9877 28698 9913 28732
rect 9947 28698 9982 28732
rect 10016 28698 10051 28732
rect 10085 28698 10120 28732
rect 10154 28698 10189 28732
rect 10223 28703 10248 28732
rect 10223 28698 10258 28703
rect 10292 28698 10327 28732
rect 10365 28703 10396 28732
rect 10448 28703 10465 28732
rect 10531 28703 10580 28737
rect 10614 28703 10615 28737
rect 10361 28698 10396 28703
rect 10430 28698 10465 28703
rect 10499 28698 10615 28703
rect 9877 28664 10615 28698
rect 9877 28630 9913 28664
rect 9947 28630 9982 28664
rect 10016 28630 10051 28664
rect 10085 28630 10120 28664
rect 10154 28630 10189 28664
rect 10223 28630 10248 28664
rect 10292 28630 10327 28664
rect 10365 28630 10396 28664
rect 10448 28630 10465 28664
rect 10531 28630 10580 28664
rect 10614 28630 10615 28664
rect 9877 28596 10615 28630
rect 9877 28562 9913 28596
rect 9947 28562 9982 28596
rect 10016 28562 10051 28596
rect 10085 28562 10120 28596
rect 10154 28562 10189 28596
rect 10223 28591 10258 28596
rect 10223 28562 10248 28591
rect 10292 28562 10327 28596
rect 10361 28591 10396 28596
rect 10430 28591 10465 28596
rect 10499 28591 10615 28596
rect 10365 28562 10396 28591
rect 10448 28562 10465 28591
rect 9877 28557 10248 28562
rect 10282 28557 10331 28562
rect 10365 28557 10414 28562
rect 10448 28557 10497 28562
rect 10531 28557 10580 28591
rect 10614 28557 10615 28591
rect 9877 28528 10615 28557
rect 9877 28494 9913 28528
rect 9947 28494 9982 28528
rect 10016 28494 10051 28528
rect 10085 28494 10120 28528
rect 10154 28494 10189 28528
rect 10223 28518 10258 28528
rect 10223 28494 10248 28518
rect 10292 28494 10327 28528
rect 10361 28518 10396 28528
rect 10430 28518 10465 28528
rect 10499 28518 10615 28528
rect 10365 28494 10396 28518
rect 10448 28494 10465 28518
rect 9877 28484 10248 28494
rect 10282 28484 10331 28494
rect 10365 28484 10414 28494
rect 10448 28484 10497 28494
rect 10531 28484 10580 28518
rect 10614 28484 10615 28518
rect 9877 28460 10615 28484
rect 9877 28426 9913 28460
rect 9947 28426 9982 28460
rect 10016 28426 10051 28460
rect 10085 28426 10120 28460
rect 10154 28426 10189 28460
rect 10223 28445 10258 28460
rect 10223 28426 10248 28445
rect 10292 28426 10327 28460
rect 10361 28445 10396 28460
rect 10430 28445 10465 28460
rect 10499 28445 10615 28460
rect 10365 28426 10396 28445
rect 10448 28426 10465 28445
rect 9877 28411 10248 28426
rect 10282 28411 10331 28426
rect 10365 28411 10414 28426
rect 10448 28411 10497 28426
rect 10531 28411 10580 28445
rect 10614 28411 10615 28445
rect 9877 28392 10615 28411
rect 9877 28358 9913 28392
rect 9947 28358 9982 28392
rect 10016 28358 10051 28392
rect 10085 28358 10120 28392
rect 10154 28358 10189 28392
rect 10223 28372 10258 28392
rect 10223 28358 10248 28372
rect 10292 28358 10327 28392
rect 10361 28372 10396 28392
rect 10430 28372 10465 28392
rect 10499 28372 10615 28392
rect 10365 28358 10396 28372
rect 10448 28358 10465 28372
rect 9877 28338 10248 28358
rect 10282 28338 10331 28358
rect 10365 28338 10414 28358
rect 10448 28338 10497 28358
rect 10531 28338 10580 28372
rect 10614 28338 10615 28372
rect 9877 28324 10615 28338
rect 9877 28290 9913 28324
rect 9947 28290 9982 28324
rect 10016 28290 10051 28324
rect 10085 28290 10120 28324
rect 10154 28290 10189 28324
rect 10223 28299 10258 28324
rect 10223 28290 10248 28299
rect 10292 28290 10327 28324
rect 10361 28299 10396 28324
rect 10430 28299 10465 28324
rect 10499 28299 10615 28324
rect 10365 28290 10396 28299
rect 10448 28290 10465 28299
rect 9877 28265 10248 28290
rect 10282 28265 10331 28290
rect 10365 28265 10414 28290
rect 10448 28265 10497 28290
rect 10531 28265 10580 28299
rect 10614 28265 10615 28299
rect 9877 28256 10615 28265
rect 9877 28222 9913 28256
rect 9947 28222 9982 28256
rect 10016 28222 10051 28256
rect 10085 28222 10120 28256
rect 10154 28222 10189 28256
rect 10223 28226 10258 28256
rect 10223 28222 10248 28226
rect 10292 28222 10327 28256
rect 10361 28226 10396 28256
rect 10430 28226 10465 28256
rect 10499 28226 10615 28256
rect 10365 28222 10396 28226
rect 10448 28222 10465 28226
rect 9877 28192 10248 28222
rect 10282 28192 10331 28222
rect 10365 28192 10414 28222
rect 10448 28192 10497 28222
rect 10531 28192 10580 28226
rect 10614 28192 10615 28226
rect 9877 28188 10615 28192
rect 9877 28154 9913 28188
rect 9947 28154 9982 28188
rect 10016 28154 10051 28188
rect 10085 28154 10120 28188
rect 10154 28154 10189 28188
rect 10223 28154 10258 28188
rect 10292 28154 10327 28188
rect 10361 28154 10396 28188
rect 10430 28154 10465 28188
rect 10499 28154 10615 28188
rect 9877 28153 10615 28154
rect 9877 28120 10248 28153
rect 10282 28120 10331 28153
rect 10365 28120 10414 28153
rect 10448 28120 10497 28153
rect 9877 28086 9913 28120
rect 9947 28086 9982 28120
rect 10016 28086 10051 28120
rect 10085 28086 10120 28120
rect 10154 28086 10189 28120
rect 10223 28119 10248 28120
rect 10223 28086 10258 28119
rect 10292 28086 10327 28120
rect 10365 28119 10396 28120
rect 10448 28119 10465 28120
rect 10531 28119 10580 28153
rect 10614 28119 10615 28153
rect 10361 28086 10396 28119
rect 10430 28086 10465 28119
rect 10499 28086 10615 28119
rect 9877 28080 10615 28086
rect 9877 28052 10248 28080
rect 10282 28052 10331 28080
rect 10365 28052 10414 28080
rect 10448 28052 10497 28080
rect 9877 28018 9913 28052
rect 9947 28018 9982 28052
rect 10016 28018 10051 28052
rect 10085 28018 10120 28052
rect 10154 28018 10189 28052
rect 10223 28046 10248 28052
rect 10223 28018 10258 28046
rect 10292 28018 10327 28052
rect 10365 28046 10396 28052
rect 10448 28046 10465 28052
rect 10531 28046 10580 28080
rect 10614 28046 10615 28080
rect 10361 28018 10396 28046
rect 10430 28018 10465 28046
rect 10499 28018 10615 28046
rect 9877 28007 10615 28018
rect 9877 27983 10248 28007
rect 10282 27983 10331 28007
rect 10365 27983 10414 28007
rect 10448 27983 10497 28007
rect 9877 27949 9913 27983
rect 9947 27949 9982 27983
rect 10016 27949 10051 27983
rect 10085 27949 10120 27983
rect 10154 27949 10189 27983
rect 10223 27973 10248 27983
rect 10223 27949 10258 27973
rect 10292 27949 10327 27983
rect 10365 27973 10396 27983
rect 10448 27973 10465 27983
rect 10531 27973 10580 28007
rect 10614 27973 10615 28007
rect 10361 27949 10396 27973
rect 10430 27949 10465 27973
rect 10499 27949 10615 27973
rect 9877 27934 10615 27949
rect 9877 27914 10248 27934
rect 10282 27914 10331 27934
rect 10365 27914 10414 27934
rect 10448 27914 10497 27934
rect 9877 27880 9913 27914
rect 9947 27880 9982 27914
rect 10016 27880 10051 27914
rect 10085 27880 10120 27914
rect 10154 27880 10189 27914
rect 10223 27900 10248 27914
rect 10223 27880 10258 27900
rect 10292 27880 10327 27914
rect 10365 27900 10396 27914
rect 10448 27900 10465 27914
rect 10531 27900 10580 27934
rect 10614 27900 10615 27934
rect 10361 27880 10396 27900
rect 10430 27880 10465 27900
rect 10499 27880 10615 27900
rect 9877 27861 10615 27880
rect 9877 27845 10248 27861
rect 10282 27845 10331 27861
rect 10365 27845 10414 27861
rect 10448 27845 10497 27861
rect 9877 27811 9913 27845
rect 9947 27811 9982 27845
rect 10016 27811 10051 27845
rect 10085 27811 10120 27845
rect 10154 27811 10189 27845
rect 10223 27827 10248 27845
rect 10223 27811 10258 27827
rect 10292 27811 10327 27845
rect 10365 27827 10396 27845
rect 10448 27827 10465 27845
rect 10531 27827 10580 27861
rect 10614 27827 10615 27861
rect 10361 27811 10396 27827
rect 10430 27811 10465 27827
rect 10499 27811 10615 27827
rect 9877 27788 10615 27811
rect 9877 27776 10248 27788
rect 10282 27776 10331 27788
rect 10365 27776 10414 27788
rect 10448 27776 10497 27788
rect 9877 27742 9913 27776
rect 9947 27742 9982 27776
rect 10016 27742 10051 27776
rect 10085 27742 10120 27776
rect 10154 27742 10189 27776
rect 10223 27754 10248 27776
rect 10223 27742 10258 27754
rect 10292 27742 10327 27776
rect 10365 27754 10396 27776
rect 10448 27754 10465 27776
rect 10531 27754 10580 27788
rect 10614 27754 10615 27788
rect 10361 27742 10396 27754
rect 10430 27742 10465 27754
rect 10499 27742 10615 27754
rect 9877 27715 10615 27742
rect 9877 27707 10248 27715
rect 10282 27707 10331 27715
rect 10365 27707 10414 27715
rect 10448 27707 10497 27715
rect 9877 27673 9913 27707
rect 9947 27673 9982 27707
rect 10016 27673 10051 27707
rect 10085 27673 10120 27707
rect 10154 27673 10189 27707
rect 10223 27681 10248 27707
rect 10223 27673 10258 27681
rect 10292 27673 10327 27707
rect 10365 27681 10396 27707
rect 10448 27681 10465 27707
rect 10531 27681 10580 27715
rect 10614 27681 10615 27715
rect 10361 27673 10396 27681
rect 10430 27673 10465 27681
rect 10499 27673 10615 27681
rect 9877 27642 10615 27673
rect 9877 27638 10248 27642
rect 10282 27638 10331 27642
rect 10365 27638 10414 27642
rect 10448 27638 10497 27642
rect 9877 27604 9913 27638
rect 9947 27604 9982 27638
rect 10016 27604 10051 27638
rect 10085 27604 10120 27638
rect 10154 27604 10189 27638
rect 10223 27608 10248 27638
rect 10223 27604 10258 27608
rect 10292 27604 10327 27638
rect 10365 27608 10396 27638
rect 10448 27608 10465 27638
rect 10531 27608 10580 27642
rect 10614 27608 10615 27642
rect 10361 27604 10396 27608
rect 10430 27604 10465 27608
rect 10499 27604 10615 27608
rect 9877 27569 10615 27604
rect 9877 27535 9913 27569
rect 9947 27535 9982 27569
rect 10016 27535 10051 27569
rect 10085 27535 10120 27569
rect 10154 27535 10189 27569
rect 10223 27568 10258 27569
rect 10223 27535 10248 27568
rect 10292 27535 10327 27569
rect 10361 27568 10396 27569
rect 10430 27568 10465 27569
rect 10499 27568 10615 27569
rect 10365 27535 10396 27568
rect 10448 27535 10465 27568
rect 9877 27534 10248 27535
rect 10282 27534 10331 27535
rect 10365 27534 10414 27535
rect 10448 27534 10497 27535
rect 10531 27534 10580 27568
rect 10614 27534 10615 27568
rect 9877 27500 10615 27534
rect 9877 27466 9913 27500
rect 9947 27466 9982 27500
rect 10016 27466 10051 27500
rect 10085 27466 10120 27500
rect 10154 27466 10189 27500
rect 10223 27494 10258 27500
rect 10223 27466 10248 27494
rect 10292 27466 10327 27500
rect 10361 27494 10396 27500
rect 10430 27494 10465 27500
rect 10499 27494 10615 27500
rect 10365 27466 10396 27494
rect 10448 27466 10465 27494
rect 9877 27460 10248 27466
rect 10282 27460 10331 27466
rect 10365 27460 10414 27466
rect 10448 27460 10497 27466
rect 10531 27460 10580 27494
rect 10614 27460 10615 27494
rect 9877 27431 10615 27460
rect 9877 27397 9913 27431
rect 9947 27397 9982 27431
rect 10016 27397 10051 27431
rect 10085 27397 10120 27431
rect 10154 27397 10189 27431
rect 10223 27420 10258 27431
rect 10223 27397 10248 27420
rect 10292 27397 10327 27431
rect 10361 27420 10396 27431
rect 10430 27420 10465 27431
rect 10499 27420 10615 27431
rect 10365 27397 10396 27420
rect 10448 27397 10465 27420
rect 9877 27386 10248 27397
rect 10282 27386 10331 27397
rect 10365 27386 10414 27397
rect 10448 27386 10497 27397
rect 10531 27386 10580 27420
rect 10614 27386 10615 27420
rect 9877 27362 10615 27386
rect 9877 27328 9913 27362
rect 9947 27328 9982 27362
rect 10016 27328 10051 27362
rect 10085 27328 10120 27362
rect 10154 27328 10189 27362
rect 10223 27346 10258 27362
rect 10223 27328 10248 27346
rect 10292 27328 10327 27362
rect 10361 27346 10396 27362
rect 10430 27346 10465 27362
rect 10499 27346 10615 27362
rect 10365 27328 10396 27346
rect 10448 27328 10465 27346
rect 9877 27312 10248 27328
rect 10282 27312 10331 27328
rect 10365 27312 10414 27328
rect 10448 27312 10497 27328
rect 10531 27312 10580 27346
rect 10614 27312 10615 27346
rect 9877 27293 10615 27312
rect 9877 27259 9913 27293
rect 9947 27259 9982 27293
rect 10016 27259 10051 27293
rect 10085 27259 10120 27293
rect 10154 27259 10189 27293
rect 10223 27272 10258 27293
rect 10223 27259 10248 27272
rect 10292 27259 10327 27293
rect 10361 27272 10396 27293
rect 10430 27272 10465 27293
rect 10499 27272 10615 27293
rect 10365 27259 10396 27272
rect 10448 27259 10465 27272
rect 9877 27238 10248 27259
rect 10282 27238 10331 27259
rect 10365 27238 10414 27259
rect 10448 27238 10497 27259
rect 10531 27238 10580 27272
rect 10614 27238 10615 27272
rect 9877 27224 10615 27238
rect 9877 27190 9913 27224
rect 9947 27190 9982 27224
rect 10016 27190 10051 27224
rect 10085 27190 10120 27224
rect 10154 27190 10189 27224
rect 10223 27198 10258 27224
rect 10223 27190 10248 27198
rect 10292 27190 10327 27224
rect 10361 27198 10396 27224
rect 10430 27198 10465 27224
rect 10499 27198 10615 27224
rect 10365 27190 10396 27198
rect 10448 27190 10465 27198
rect 9877 27164 10248 27190
rect 10282 27164 10331 27190
rect 10365 27164 10414 27190
rect 10448 27164 10497 27190
rect 10531 27164 10580 27198
rect 10614 27164 10615 27198
rect 9877 27155 10615 27164
rect 9877 27121 9913 27155
rect 9947 27121 9982 27155
rect 10016 27121 10051 27155
rect 10085 27121 10120 27155
rect 10154 27121 10189 27155
rect 10223 27124 10258 27155
rect 10223 27121 10248 27124
rect 10292 27121 10327 27155
rect 10361 27124 10396 27155
rect 10430 27124 10465 27155
rect 10499 27124 10615 27155
rect 10365 27121 10396 27124
rect 10448 27121 10465 27124
rect 9877 27090 10248 27121
rect 10282 27090 10331 27121
rect 10365 27090 10414 27121
rect 10448 27090 10497 27121
rect 10531 27090 10580 27124
rect 10614 27090 10615 27124
rect 9877 27086 10615 27090
rect 9877 27052 9913 27086
rect 9947 27052 9982 27086
rect 10016 27052 10051 27086
rect 10085 27052 10120 27086
rect 10154 27052 10189 27086
rect 10223 27052 10258 27086
rect 10292 27052 10327 27086
rect 10361 27052 10396 27086
rect 10430 27052 10465 27086
rect 10499 27052 10615 27086
rect 9877 27050 10615 27052
rect 9877 27016 10248 27050
rect 10282 27016 10331 27050
rect 10365 27016 10414 27050
rect 10448 27016 10497 27050
rect 10531 27016 10580 27050
rect 10614 27016 10615 27050
rect 9877 26976 10615 27016
rect 9877 26942 10248 26976
rect 10282 26942 10331 26976
rect 10365 26942 10414 26976
rect 10448 26942 10497 26976
rect 10531 26942 10580 26976
rect 10614 26972 10615 26976
rect 13703 29172 13705 29206
rect 13703 29133 13738 29172
rect 13908 29178 13909 29212
rect 13943 29178 13944 29212
rect 13908 29140 13944 29178
rect 13703 29099 13705 29133
rect 13703 29060 13738 29099
rect 13908 29106 13909 29140
rect 13943 29106 13944 29140
rect 13908 29068 13944 29106
rect 13703 29026 13705 29060
rect 13703 29007 13738 29026
rect 13908 29034 13909 29068
rect 13943 29034 13944 29068
rect 13908 29007 13944 29034
rect 13703 28996 13944 29007
rect 13703 28987 13909 28996
rect 13703 28953 13705 28987
rect 13739 28984 13909 28987
rect 13739 28972 13807 28984
rect 13841 28972 13909 28984
rect 13703 28938 13738 28953
rect 13772 28938 13806 28972
rect 13841 28950 13874 28972
rect 13840 28938 13874 28950
rect 13908 28962 13909 28972
rect 13943 28962 13944 28996
rect 13908 28938 13944 28962
rect 13703 28924 13944 28938
rect 13703 28914 13909 28924
rect 13703 28880 13705 28914
rect 13739 28911 13909 28914
rect 13739 28903 13807 28911
rect 13841 28903 13909 28911
rect 13703 28869 13738 28880
rect 13772 28869 13806 28903
rect 13841 28877 13874 28903
rect 13840 28869 13874 28877
rect 13908 28890 13909 28903
rect 13943 28890 13944 28924
rect 13908 28869 13944 28890
rect 13703 28852 13944 28869
rect 13703 28841 13909 28852
rect 13703 28807 13705 28841
rect 13739 28838 13909 28841
rect 13739 28834 13807 28838
rect 13841 28834 13909 28838
rect 13703 28800 13738 28807
rect 13772 28800 13806 28834
rect 13841 28804 13874 28834
rect 13840 28800 13874 28804
rect 13908 28818 13909 28834
rect 13943 28818 13944 28852
rect 13908 28800 13944 28818
rect 13703 28780 13944 28800
rect 13703 28769 13909 28780
rect 13703 28735 13705 28769
rect 13739 28765 13909 28769
rect 13703 28731 13738 28735
rect 13772 28731 13806 28765
rect 13841 28731 13874 28765
rect 13908 28746 13909 28765
rect 13943 28746 13944 28780
rect 13908 28731 13944 28746
rect 13703 28708 13944 28731
rect 13703 28697 13909 28708
rect 13703 28663 13705 28697
rect 13739 28696 13909 28697
rect 13703 28662 13738 28663
rect 13772 28662 13806 28696
rect 13840 28692 13874 28696
rect 13841 28662 13874 28692
rect 13908 28674 13909 28696
rect 13943 28674 13944 28708
rect 13908 28662 13944 28674
rect 13703 28658 13807 28662
rect 13841 28658 13944 28662
rect 13703 28636 13944 28658
rect 13703 28627 13909 28636
rect 13703 28625 13738 28627
rect 13703 28591 13705 28625
rect 13772 28593 13806 28627
rect 13840 28619 13874 28627
rect 13841 28593 13874 28619
rect 13908 28602 13909 28627
rect 13943 28602 13944 28636
rect 13908 28593 13944 28602
rect 13739 28591 13807 28593
rect 13703 28585 13807 28591
rect 13841 28585 13944 28593
rect 13703 28564 13944 28585
rect 13703 28558 13909 28564
rect 13703 28553 13738 28558
rect 13703 28519 13705 28553
rect 13772 28524 13806 28558
rect 13840 28546 13874 28558
rect 13841 28524 13874 28546
rect 13908 28530 13909 28558
rect 13943 28530 13944 28564
rect 13908 28524 13944 28530
rect 13739 28519 13807 28524
rect 13703 28512 13807 28519
rect 13841 28512 13944 28524
rect 13703 28492 13944 28512
rect 13703 28489 13909 28492
rect 13703 28481 13738 28489
rect 13703 28447 13705 28481
rect 13772 28455 13806 28489
rect 13840 28473 13874 28489
rect 13841 28455 13874 28473
rect 13908 28458 13909 28489
rect 13943 28458 13944 28492
rect 13908 28455 13944 28458
rect 13739 28447 13807 28455
rect 13703 28439 13807 28447
rect 13841 28439 13944 28455
rect 13703 28420 13944 28439
rect 13703 28409 13738 28420
rect 13703 28375 13705 28409
rect 13772 28386 13806 28420
rect 13840 28400 13874 28420
rect 13841 28386 13874 28400
rect 13908 28386 13909 28420
rect 13943 28386 13944 28420
rect 13739 28375 13807 28386
rect 13703 28366 13807 28375
rect 13841 28366 13944 28386
rect 13703 28351 13944 28366
rect 13703 28337 13738 28351
rect 13703 28303 13705 28337
rect 13772 28317 13806 28351
rect 13840 28327 13874 28351
rect 13841 28317 13874 28327
rect 13908 28348 13944 28351
rect 13908 28317 13909 28348
rect 13739 28303 13807 28317
rect 13703 28293 13807 28303
rect 13841 28314 13909 28317
rect 13943 28314 13944 28348
rect 13841 28293 13944 28314
rect 13703 28282 13944 28293
rect 13703 28265 13738 28282
rect 13703 28231 13705 28265
rect 13772 28248 13806 28282
rect 13840 28254 13874 28282
rect 13841 28248 13874 28254
rect 13908 28276 13944 28282
rect 13908 28248 13909 28276
rect 13739 28231 13807 28248
rect 13703 28220 13807 28231
rect 13841 28242 13909 28248
rect 13943 28242 13944 28276
rect 13841 28220 13944 28242
rect 13703 28213 13944 28220
rect 13703 28193 13738 28213
rect 13703 28159 13705 28193
rect 13772 28179 13806 28213
rect 13840 28181 13874 28213
rect 13841 28179 13874 28181
rect 13908 28204 13944 28213
rect 13908 28179 13909 28204
rect 13739 28159 13807 28179
rect 13703 28147 13807 28159
rect 13841 28170 13909 28179
rect 13943 28170 13944 28204
rect 13841 28147 13944 28170
rect 13703 28144 13944 28147
rect 13703 28121 13738 28144
rect 13703 28087 13705 28121
rect 13772 28110 13806 28144
rect 13840 28110 13874 28144
rect 13908 28132 13944 28144
rect 13908 28110 13909 28132
rect 13739 28108 13909 28110
rect 13739 28087 13807 28108
rect 13703 28075 13807 28087
rect 13841 28098 13909 28108
rect 13943 28098 13944 28132
rect 13841 28075 13944 28098
rect 13703 28049 13738 28075
rect 13703 28015 13705 28049
rect 13772 28041 13806 28075
rect 13841 28074 13874 28075
rect 13840 28041 13874 28074
rect 13908 28060 13944 28075
rect 13908 28041 13909 28060
rect 13739 28035 13909 28041
rect 13739 28015 13807 28035
rect 13703 28006 13807 28015
rect 13841 28026 13909 28035
rect 13943 28026 13944 28060
rect 13841 28006 13944 28026
rect 13703 27977 13738 28006
rect 13703 27943 13705 27977
rect 13772 27972 13806 28006
rect 13841 28001 13874 28006
rect 13840 27972 13874 28001
rect 13908 27988 13944 28006
rect 13908 27972 13909 27988
rect 13739 27962 13909 27972
rect 13739 27943 13807 27962
rect 13703 27937 13807 27943
rect 13841 27954 13909 27962
rect 13943 27954 13944 27988
rect 13841 27937 13944 27954
rect 13703 27905 13738 27937
rect 13703 27871 13705 27905
rect 13772 27903 13806 27937
rect 13841 27928 13874 27937
rect 13840 27903 13874 27928
rect 13908 27916 13944 27937
rect 13908 27903 13909 27916
rect 13739 27889 13909 27903
rect 13739 27871 13807 27889
rect 13703 27868 13807 27871
rect 13841 27882 13909 27889
rect 13943 27882 13944 27916
rect 13841 27868 13944 27882
rect 13703 27834 13738 27868
rect 13772 27834 13806 27868
rect 13841 27855 13874 27868
rect 13840 27834 13874 27855
rect 13908 27844 13944 27868
rect 13908 27834 13909 27844
rect 13703 27833 13909 27834
rect 13703 27799 13705 27833
rect 13739 27816 13909 27833
rect 13739 27799 13807 27816
rect 13841 27810 13909 27816
rect 13943 27810 13944 27844
rect 13841 27799 13944 27810
rect 13703 27765 13738 27799
rect 13772 27765 13806 27799
rect 13841 27782 13874 27799
rect 13840 27765 13874 27782
rect 13908 27772 13944 27799
rect 13908 27765 13909 27772
rect 13703 27761 13909 27765
rect 13703 27727 13705 27761
rect 13739 27743 13909 27761
rect 13739 27730 13807 27743
rect 13841 27738 13909 27743
rect 13943 27738 13944 27772
rect 13841 27730 13944 27738
rect 13703 27696 13738 27727
rect 13772 27696 13806 27730
rect 13841 27709 13874 27730
rect 13840 27696 13874 27709
rect 13908 27700 13944 27730
rect 13908 27696 13909 27700
rect 13703 27689 13909 27696
rect 13703 27655 13705 27689
rect 13739 27670 13909 27689
rect 13739 27661 13807 27670
rect 13841 27666 13909 27670
rect 13943 27666 13944 27700
rect 13841 27661 13944 27666
rect 13703 27627 13738 27655
rect 13772 27627 13806 27661
rect 13841 27636 13874 27661
rect 13840 27627 13874 27636
rect 13908 27628 13944 27661
rect 13908 27627 13909 27628
rect 13703 27617 13909 27627
rect 13703 27583 13705 27617
rect 13739 27597 13909 27617
rect 13739 27592 13807 27597
rect 13841 27594 13909 27597
rect 13943 27594 13944 27628
rect 13841 27592 13944 27594
rect 13703 27558 13738 27583
rect 13772 27558 13806 27592
rect 13841 27563 13874 27592
rect 13840 27558 13874 27563
rect 13908 27558 13944 27592
rect 13703 27556 13944 27558
rect 13703 27545 13909 27556
rect 13703 27511 13705 27545
rect 13739 27524 13909 27545
rect 13739 27523 13807 27524
rect 13841 27523 13909 27524
rect 13703 27489 13738 27511
rect 13772 27489 13806 27523
rect 13841 27490 13874 27523
rect 13840 27489 13874 27490
rect 13908 27522 13909 27523
rect 13943 27522 13944 27556
rect 13908 27489 13944 27522
rect 13703 27484 13944 27489
rect 13703 27473 13909 27484
rect 13703 27439 13705 27473
rect 13739 27454 13909 27473
rect 13703 27420 13738 27439
rect 13772 27420 13806 27454
rect 13840 27451 13874 27454
rect 13841 27420 13874 27451
rect 13908 27450 13909 27454
rect 13943 27450 13944 27484
rect 13908 27420 13944 27450
rect 13703 27417 13807 27420
rect 13841 27417 13944 27420
rect 13703 27412 13944 27417
rect 13703 27401 13909 27412
rect 13703 27367 13705 27401
rect 13739 27385 13909 27401
rect 13703 27351 13738 27367
rect 13772 27351 13806 27385
rect 13840 27378 13874 27385
rect 13841 27351 13874 27378
rect 13908 27378 13909 27385
rect 13943 27378 13944 27412
rect 13908 27351 13944 27378
rect 13703 27344 13807 27351
rect 13841 27344 13944 27351
rect 13703 27340 13944 27344
rect 13703 27329 13909 27340
rect 13703 27295 13705 27329
rect 13739 27316 13909 27329
rect 13703 27282 13738 27295
rect 13772 27282 13806 27316
rect 13840 27305 13874 27316
rect 13841 27282 13874 27305
rect 13908 27306 13909 27316
rect 13943 27306 13944 27340
rect 13908 27282 13944 27306
rect 13703 27271 13807 27282
rect 13841 27271 13944 27282
rect 13703 27268 13944 27271
rect 13703 27257 13909 27268
rect 13703 27223 13705 27257
rect 13739 27247 13909 27257
rect 13703 27213 13738 27223
rect 13772 27213 13806 27247
rect 13840 27232 13874 27247
rect 13841 27213 13874 27232
rect 13908 27234 13909 27247
rect 13943 27234 13944 27268
rect 13908 27213 13944 27234
rect 13703 27198 13807 27213
rect 13841 27198 13944 27213
rect 13703 27196 13944 27198
rect 13703 27185 13909 27196
rect 13703 27151 13705 27185
rect 13739 27178 13909 27185
rect 13703 27144 13738 27151
rect 13772 27144 13806 27178
rect 13840 27159 13874 27178
rect 13841 27144 13874 27159
rect 13908 27162 13909 27178
rect 13943 27162 13944 27196
rect 13908 27144 13944 27162
rect 13703 27125 13807 27144
rect 13841 27125 13944 27144
rect 13703 27124 13944 27125
rect 13703 27113 13909 27124
rect 13703 27079 13705 27113
rect 13739 27109 13909 27113
rect 13703 27075 13738 27079
rect 13772 27075 13806 27109
rect 13840 27086 13874 27109
rect 13841 27075 13874 27086
rect 13908 27090 13909 27109
rect 13943 27090 13944 27124
rect 13908 27075 13944 27090
rect 13703 27052 13807 27075
rect 13841 27052 13944 27075
rect 13703 27041 13909 27052
rect 13703 27007 13705 27041
rect 13739 27040 13909 27041
rect 13703 27006 13738 27007
rect 13772 27006 13806 27040
rect 13840 27013 13874 27040
rect 13841 27006 13874 27013
rect 13908 27018 13909 27040
rect 13943 27018 13944 27052
rect 13908 27006 13944 27018
rect 13703 26979 13807 27006
rect 13841 26980 13944 27006
rect 13841 26979 13909 26980
rect 13703 26972 13909 26979
rect 10614 26969 13909 26972
rect 10614 26942 10659 26969
rect 9877 26938 10659 26942
rect 10693 26938 10731 26969
rect 10765 26938 10803 26969
rect 10837 26938 10875 26969
rect 10909 26938 10947 26969
rect 10981 26938 11019 26969
rect 11053 26938 11091 26969
rect 11125 26938 11163 26969
rect 11197 26938 11235 26969
rect 11269 26938 11307 26969
rect 11341 26938 11379 26969
rect 11413 26938 11451 26969
rect 11485 26938 11523 26969
rect 11557 26938 11595 26969
rect 11629 26938 11667 26969
rect 11701 26938 11739 26969
rect 11773 26938 11811 26969
rect 11845 26938 11883 26969
rect 11917 26938 11955 26969
rect 11989 26938 12027 26969
rect 12061 26938 12099 26969
rect 12133 26938 12172 26969
rect 12206 26938 12245 26969
rect 12279 26938 12318 26969
rect 12352 26938 12391 26969
rect 12425 26938 12464 26969
rect 12498 26938 12537 26969
rect 12571 26938 12610 26969
rect 12644 26938 12683 26969
rect 12717 26938 12756 26969
rect 12790 26938 12829 26969
rect 12863 26938 12902 26969
rect 12936 26938 12975 26969
rect 13009 26938 13048 26969
rect 13082 26938 13121 26969
rect 13155 26938 13194 26969
rect 13228 26938 13267 26969
rect 13301 26938 13340 26969
rect 13374 26938 13413 26969
rect 13447 26938 13486 26969
rect 13520 26938 13559 26969
rect 13593 26938 13632 26969
rect 13666 26938 13705 26969
rect 9877 26904 9911 26938
rect 9945 26904 9980 26938
rect 10014 26904 10049 26938
rect 10083 26904 10118 26938
rect 10152 26904 10187 26938
rect 10221 26904 10256 26938
rect 10290 26904 10325 26938
rect 10359 26904 10394 26938
rect 10428 26904 10463 26938
rect 10497 26904 10532 26938
rect 10566 26904 10601 26938
rect 10635 26935 10659 26938
rect 10704 26935 10731 26938
rect 10773 26935 10803 26938
rect 10842 26935 10875 26938
rect 10635 26904 10670 26935
rect 10704 26904 10739 26935
rect 10773 26904 10808 26935
rect 10842 26904 10877 26935
rect 10911 26904 10946 26938
rect 10981 26935 11015 26938
rect 11053 26935 11084 26938
rect 11125 26935 11153 26938
rect 11197 26935 11222 26938
rect 11269 26935 11291 26938
rect 11341 26935 11359 26938
rect 11413 26935 11427 26938
rect 11485 26935 11495 26938
rect 11557 26935 11563 26938
rect 11629 26935 11631 26938
rect 10980 26904 11015 26935
rect 11049 26904 11084 26935
rect 11118 26904 11153 26935
rect 11187 26904 11222 26935
rect 11256 26904 11291 26935
rect 11325 26904 11359 26935
rect 11393 26904 11427 26935
rect 11461 26904 11495 26935
rect 11529 26904 11563 26935
rect 11597 26904 11631 26935
rect 11665 26935 11667 26938
rect 11733 26935 11739 26938
rect 11801 26935 11811 26938
rect 11869 26935 11883 26938
rect 11937 26935 11955 26938
rect 12005 26935 12027 26938
rect 12073 26935 12099 26938
rect 12141 26935 12172 26938
rect 11665 26904 11699 26935
rect 11733 26904 11767 26935
rect 11801 26904 11835 26935
rect 11869 26904 11903 26935
rect 11937 26904 11971 26935
rect 12005 26904 12039 26935
rect 12073 26904 12107 26935
rect 12141 26904 12175 26935
rect 12209 26904 12243 26938
rect 12279 26935 12311 26938
rect 12352 26935 12379 26938
rect 12425 26935 12447 26938
rect 12498 26935 12515 26938
rect 12571 26935 12583 26938
rect 12644 26935 12651 26938
rect 12717 26935 12719 26938
rect 12277 26904 12311 26935
rect 12345 26904 12379 26935
rect 12413 26904 12447 26935
rect 12481 26904 12515 26935
rect 12549 26904 12583 26935
rect 12617 26904 12651 26935
rect 12685 26904 12719 26935
rect 12753 26935 12756 26938
rect 12821 26935 12829 26938
rect 12889 26935 12902 26938
rect 12957 26935 12975 26938
rect 13025 26935 13048 26938
rect 13093 26935 13121 26938
rect 13161 26935 13194 26938
rect 12753 26904 12787 26935
rect 12821 26904 12855 26935
rect 12889 26904 12923 26935
rect 12957 26904 12991 26935
rect 13025 26904 13059 26935
rect 13093 26904 13127 26935
rect 13161 26904 13195 26935
rect 13229 26904 13263 26938
rect 13301 26935 13331 26938
rect 13374 26935 13399 26938
rect 13447 26935 13467 26938
rect 13520 26935 13535 26938
rect 13593 26935 13603 26938
rect 13666 26935 13671 26938
rect 13297 26904 13331 26935
rect 13365 26904 13399 26935
rect 13433 26904 13467 26935
rect 13501 26904 13535 26935
rect 13569 26904 13603 26935
rect 13637 26904 13671 26935
rect 13739 26946 13909 26969
rect 13943 26946 13944 26980
rect 13739 26940 13944 26946
rect 13739 26938 13807 26940
rect 13841 26938 13944 26940
rect 13705 26904 13739 26935
rect 13773 26904 13807 26938
rect 13841 26904 13875 26938
rect 13909 26908 13944 26938
rect 9877 26902 13909 26904
rect 9877 26868 10248 26902
rect 10282 26868 10331 26902
rect 10365 26868 10414 26902
rect 10448 26868 10497 26902
rect 10531 26868 10580 26902
rect 10614 26874 13909 26902
rect 13943 26874 13944 26908
rect 10614 26868 13944 26874
rect 9877 26867 13944 26868
rect 9877 26866 10659 26867
rect 10693 26866 10732 26867
rect 10766 26866 10805 26867
rect 10839 26866 10878 26867
rect 10912 26866 10951 26867
rect 10985 26866 11024 26867
rect 11058 26866 11097 26867
rect 11131 26866 11170 26867
rect 11204 26866 11243 26867
rect 11277 26866 11316 26867
rect 11350 26866 11389 26867
rect 11423 26866 11462 26867
rect 11496 26866 11535 26867
rect 11569 26866 11608 26867
rect 11642 26866 11681 26867
rect 11715 26866 11754 26867
rect 11788 26866 11827 26867
rect 11861 26866 11900 26867
rect 11934 26866 11973 26867
rect 12007 26866 12046 26867
rect 12080 26866 12119 26867
rect 12153 26866 12192 26867
rect 12226 26866 12265 26867
rect 12299 26866 12338 26867
rect 12372 26866 12411 26867
rect 12445 26866 12484 26867
rect 12518 26866 12557 26867
rect 12591 26866 12630 26867
rect 12664 26866 12703 26867
rect 12737 26866 12776 26867
rect 12810 26866 12849 26867
rect 12883 26866 12922 26867
rect 12956 26866 12995 26867
rect 13029 26866 13068 26867
rect 13102 26866 13141 26867
rect 13175 26866 13215 26867
rect 13249 26866 13289 26867
rect 13323 26866 13363 26867
rect 13397 26866 13437 26867
rect 13471 26866 13511 26867
rect 13545 26866 13585 26867
rect 13619 26866 13659 26867
rect 13693 26866 13733 26867
rect 13767 26866 13807 26867
rect 13841 26866 13944 26867
rect 9877 26832 9911 26866
rect 9945 26832 9980 26866
rect 10014 26832 10049 26866
rect 10083 26832 10118 26866
rect 10152 26832 10187 26866
rect 10221 26832 10256 26866
rect 10290 26832 10325 26866
rect 10359 26832 10394 26866
rect 10428 26832 10463 26866
rect 10497 26832 10532 26866
rect 10566 26832 10601 26866
rect 10635 26833 10659 26866
rect 10704 26833 10732 26866
rect 10773 26833 10805 26866
rect 10635 26832 10670 26833
rect 10704 26832 10739 26833
rect 10773 26832 10808 26833
rect 10842 26832 10877 26866
rect 10912 26833 10946 26866
rect 10985 26833 11015 26866
rect 11058 26833 11084 26866
rect 11131 26833 11153 26866
rect 11204 26833 11222 26866
rect 11277 26833 11291 26866
rect 11350 26833 11359 26866
rect 11423 26833 11427 26866
rect 10911 26832 10946 26833
rect 10980 26832 11015 26833
rect 11049 26832 11084 26833
rect 11118 26832 11153 26833
rect 11187 26832 11222 26833
rect 11256 26832 11291 26833
rect 11325 26832 11359 26833
rect 11393 26832 11427 26833
rect 11461 26833 11462 26866
rect 11529 26833 11535 26866
rect 11597 26833 11608 26866
rect 11665 26833 11681 26866
rect 11733 26833 11754 26866
rect 11801 26833 11827 26866
rect 11869 26833 11900 26866
rect 11461 26832 11495 26833
rect 11529 26832 11563 26833
rect 11597 26832 11631 26833
rect 11665 26832 11699 26833
rect 11733 26832 11767 26833
rect 11801 26832 11835 26833
rect 11869 26832 11903 26833
rect 11937 26832 11971 26866
rect 12007 26833 12039 26866
rect 12080 26833 12107 26866
rect 12153 26833 12175 26866
rect 12226 26833 12243 26866
rect 12299 26833 12311 26866
rect 12372 26833 12379 26866
rect 12445 26833 12447 26866
rect 12005 26832 12039 26833
rect 12073 26832 12107 26833
rect 12141 26832 12175 26833
rect 12209 26832 12243 26833
rect 12277 26832 12311 26833
rect 12345 26832 12379 26833
rect 12413 26832 12447 26833
rect 12481 26833 12484 26866
rect 12549 26833 12557 26866
rect 12617 26833 12630 26866
rect 12685 26833 12703 26866
rect 12753 26833 12776 26866
rect 12821 26833 12849 26866
rect 12889 26833 12922 26866
rect 12481 26832 12515 26833
rect 12549 26832 12583 26833
rect 12617 26832 12651 26833
rect 12685 26832 12719 26833
rect 12753 26832 12787 26833
rect 12821 26832 12855 26833
rect 12889 26832 12923 26833
rect 12957 26832 12991 26866
rect 13029 26833 13059 26866
rect 13102 26833 13127 26866
rect 13175 26833 13195 26866
rect 13249 26833 13263 26866
rect 13323 26833 13331 26866
rect 13397 26833 13399 26866
rect 13025 26832 13059 26833
rect 13093 26832 13127 26833
rect 13161 26832 13195 26833
rect 13229 26832 13263 26833
rect 13297 26832 13331 26833
rect 13365 26832 13399 26833
rect 13433 26833 13437 26866
rect 13501 26833 13511 26866
rect 13569 26833 13585 26866
rect 13637 26833 13659 26866
rect 13705 26833 13733 26866
rect 13433 26832 13467 26833
rect 13501 26832 13535 26833
rect 13569 26832 13603 26833
rect 13637 26832 13671 26833
rect 13705 26832 13739 26833
rect 13773 26832 13807 26866
rect 13841 26832 13875 26866
rect 13909 26836 13944 26866
rect 9877 26828 13909 26832
rect 9877 26794 10248 26828
rect 10282 26794 10331 26828
rect 10365 26794 10414 26828
rect 10448 26794 10497 26828
rect 10531 26794 10580 26828
rect 10614 26802 13909 26828
rect 13943 26802 13944 26836
rect 10614 26794 13944 26802
rect 9877 26760 9911 26794
rect 9945 26760 9980 26794
rect 10014 26760 10049 26794
rect 10083 26760 10118 26794
rect 10152 26760 10187 26794
rect 10221 26760 10256 26794
rect 10290 26760 10325 26794
rect 10359 26760 10394 26794
rect 10428 26760 10463 26794
rect 10497 26760 10532 26794
rect 10566 26760 10601 26794
rect 10635 26765 10670 26794
rect 10704 26765 10739 26794
rect 10773 26765 10808 26794
rect 10842 26765 10877 26794
rect 10635 26760 10659 26765
rect 10704 26760 10731 26765
rect 10773 26760 10803 26765
rect 10842 26760 10875 26765
rect 10911 26760 10946 26794
rect 10980 26765 11015 26794
rect 11049 26765 11084 26794
rect 11118 26765 11153 26794
rect 11187 26765 11222 26794
rect 11256 26765 11291 26794
rect 11325 26765 11359 26794
rect 11393 26765 11427 26794
rect 11461 26765 11495 26794
rect 11529 26765 11563 26794
rect 11597 26765 11631 26794
rect 10981 26760 11015 26765
rect 11053 26760 11084 26765
rect 11125 26760 11153 26765
rect 11197 26760 11222 26765
rect 11269 26760 11291 26765
rect 11341 26760 11359 26765
rect 11413 26760 11427 26765
rect 11485 26760 11495 26765
rect 11557 26760 11563 26765
rect 11629 26760 11631 26765
rect 11665 26765 11699 26794
rect 11733 26765 11767 26794
rect 11801 26765 11835 26794
rect 11869 26765 11903 26794
rect 11937 26765 11971 26794
rect 12005 26765 12039 26794
rect 12073 26765 12107 26794
rect 12141 26765 12175 26794
rect 11665 26760 11667 26765
rect 11733 26760 11739 26765
rect 11801 26760 11811 26765
rect 11869 26760 11883 26765
rect 11937 26760 11955 26765
rect 12005 26760 12027 26765
rect 12073 26760 12099 26765
rect 12141 26760 12171 26765
rect 12209 26760 12243 26794
rect 12277 26760 12311 26794
rect 12345 26765 12379 26794
rect 12413 26765 12447 26794
rect 12481 26765 12515 26794
rect 12549 26765 12583 26794
rect 12617 26765 12651 26794
rect 12685 26765 12719 26794
rect 12753 26765 12787 26794
rect 12821 26765 12855 26794
rect 12349 26760 12379 26765
rect 12421 26760 12447 26765
rect 12493 26760 12515 26765
rect 12565 26760 12583 26765
rect 12637 26760 12651 26765
rect 12709 26760 12719 26765
rect 12781 26760 12787 26765
rect 12853 26760 12855 26765
rect 12889 26765 12923 26794
rect 12957 26765 12991 26794
rect 13025 26765 13059 26794
rect 13093 26765 13127 26794
rect 13161 26765 13195 26794
rect 13229 26765 13263 26794
rect 13297 26765 13331 26794
rect 12889 26760 12891 26765
rect 12957 26760 12963 26765
rect 13025 26760 13035 26765
rect 13093 26760 13108 26765
rect 13161 26760 13181 26765
rect 13229 26760 13254 26765
rect 13297 26760 13327 26765
rect 13365 26760 13399 26794
rect 13433 26765 13467 26794
rect 13501 26765 13535 26794
rect 13569 26765 13603 26794
rect 13637 26765 13671 26794
rect 13705 26765 13739 26794
rect 13773 26765 13807 26794
rect 13841 26765 13875 26794
rect 13434 26760 13467 26765
rect 13507 26760 13535 26765
rect 13580 26760 13603 26765
rect 13653 26760 13671 26765
rect 13726 26760 13739 26765
rect 13799 26760 13807 26765
rect 13872 26760 13875 26765
rect 13909 26760 13944 26794
rect 9877 26754 10659 26760
rect 9877 26726 10248 26754
rect 10176 26720 10248 26726
rect 10282 26720 10331 26754
rect 10365 26720 10414 26754
rect 10448 26720 10497 26754
rect 10531 26720 10580 26754
rect 10614 26731 10659 26754
rect 10693 26731 10731 26760
rect 10765 26731 10803 26760
rect 10837 26731 10875 26760
rect 10909 26731 10947 26760
rect 10981 26731 11019 26760
rect 11053 26731 11091 26760
rect 11125 26731 11163 26760
rect 11197 26731 11235 26760
rect 11269 26731 11307 26760
rect 11341 26731 11379 26760
rect 11413 26731 11451 26760
rect 11485 26731 11523 26760
rect 11557 26731 11595 26760
rect 11629 26731 11667 26760
rect 11701 26731 11739 26760
rect 11773 26731 11811 26760
rect 11845 26731 11883 26760
rect 11917 26731 11955 26760
rect 11989 26731 12027 26760
rect 12061 26731 12099 26760
rect 12133 26731 12171 26760
rect 12205 26731 12243 26760
rect 12277 26731 12315 26760
rect 12349 26731 12387 26760
rect 12421 26731 12459 26760
rect 12493 26731 12531 26760
rect 12565 26731 12603 26760
rect 12637 26731 12675 26760
rect 12709 26731 12747 26760
rect 12781 26731 12819 26760
rect 12853 26731 12891 26760
rect 12925 26731 12963 26760
rect 12997 26731 13035 26760
rect 13069 26731 13108 26760
rect 13142 26731 13181 26760
rect 13215 26731 13254 26760
rect 13288 26731 13327 26760
rect 13361 26731 13400 26760
rect 13434 26731 13473 26760
rect 13507 26731 13546 26760
rect 13580 26731 13619 26760
rect 13653 26731 13692 26760
rect 13726 26731 13765 26760
rect 13799 26731 13838 26760
rect 13872 26731 13944 26760
rect 10614 26730 13944 26731
rect 10614 26726 13943 26730
rect 10614 26720 10615 26726
rect 14096 26573 14097 30788
rect 9725 26572 14097 26573
rect 9725 26402 9759 26572
rect 14009 26568 14097 26572
rect 14009 26534 14030 26568
rect 14064 26538 14097 26568
rect 14064 26534 14102 26538
rect 14136 26534 14165 26538
rect 14009 26504 14165 26534
rect 14077 26470 14165 26504
rect 14077 26469 14233 26470
rect 14267 26469 14268 30856
rect 14077 26440 14268 26469
rect 14077 26406 14086 26440
rect 14120 26436 14158 26440
rect 14145 26406 14158 26436
rect 14192 26406 14268 26440
rect 14077 26402 14111 26406
rect 14145 26402 14268 26406
rect 9725 26401 14268 26402
rect 9877 26214 9909 26248
rect 9943 26214 9981 26248
rect 10015 26214 10053 26248
rect 10087 26214 10125 26248
rect 10159 26214 10197 26248
rect 10231 26214 10269 26248
rect 10303 26214 10341 26248
rect 10375 26214 10413 26248
rect 10447 26214 10485 26248
rect 10519 26214 10557 26248
rect 10591 26214 10629 26248
rect 10663 26214 10701 26248
rect 10735 26214 10773 26248
rect 10807 26214 10845 26248
rect 10879 26214 10917 26248
rect 10951 26214 10989 26248
rect 11023 26214 11061 26248
rect 11095 26214 11133 26248
rect 11167 26214 11205 26248
rect 11239 26214 11277 26248
rect 11311 26214 11349 26248
rect 11383 26214 11421 26248
rect 11455 26214 11493 26248
rect 11527 26214 11565 26248
rect 11599 26214 11637 26248
rect 11671 26214 11709 26248
rect 11743 26214 11781 26248
rect 11815 26214 11853 26248
rect 11887 26214 11925 26248
rect 11959 26214 11997 26248
rect 12031 26214 12069 26248
rect 12103 26214 12141 26248
rect 12175 26214 12213 26248
rect 12247 26214 12285 26248
rect 12319 26214 12357 26248
rect 12391 26214 12429 26248
rect 12463 26214 12501 26248
rect 12535 26214 12573 26248
rect 12607 26214 12645 26248
rect 12679 26214 12717 26248
rect 12751 26214 12789 26248
rect 12823 26214 12861 26248
rect 12895 26214 12933 26248
rect 12967 26214 13005 26248
rect 13039 26214 13077 26248
rect 13111 26214 13149 26248
rect 13183 26214 13221 26248
rect 13255 26214 13293 26248
rect 13327 26214 13365 26248
rect 13399 26214 13437 26248
rect 13471 26214 13509 26248
rect 13543 26214 13581 26248
rect 13615 26214 13653 26248
rect 13687 26214 13756 26248
rect 13790 26214 13828 26248
rect 13862 26214 13900 26248
rect 13934 26214 13972 26248
rect 14006 26214 14044 26248
rect 14078 26214 14116 26248
rect 14150 26224 14429 26248
rect 14150 26214 14233 26224
rect 9877 26199 14233 26214
rect 9877 26174 9911 26199
rect 9877 26140 9909 26174
rect 9945 26165 9980 26199
rect 10014 26174 10049 26199
rect 10083 26174 10118 26199
rect 10152 26174 10187 26199
rect 10221 26174 10256 26199
rect 10290 26174 10325 26199
rect 10359 26174 10394 26199
rect 10428 26174 10463 26199
rect 10497 26174 10532 26199
rect 10566 26174 10601 26199
rect 10635 26174 10670 26199
rect 10704 26174 10739 26199
rect 10015 26165 10049 26174
rect 10087 26165 10118 26174
rect 10159 26165 10187 26174
rect 10231 26165 10256 26174
rect 10303 26165 10325 26174
rect 10375 26165 10394 26174
rect 10447 26165 10463 26174
rect 10519 26165 10532 26174
rect 10591 26165 10601 26174
rect 10663 26165 10670 26174
rect 10735 26165 10739 26174
rect 10773 26174 10807 26199
rect 9943 26140 9981 26165
rect 10015 26140 10053 26165
rect 10087 26140 10125 26165
rect 10159 26140 10197 26165
rect 10231 26140 10269 26165
rect 10303 26140 10341 26165
rect 10375 26140 10413 26165
rect 10447 26140 10485 26165
rect 10519 26140 10557 26165
rect 10591 26140 10629 26165
rect 10663 26140 10701 26165
rect 10735 26140 10773 26165
rect 10841 26174 10875 26199
rect 10909 26174 10943 26199
rect 10977 26174 11011 26199
rect 11045 26174 11079 26199
rect 11113 26174 11147 26199
rect 11181 26174 11215 26199
rect 11249 26174 11283 26199
rect 11317 26174 11351 26199
rect 10841 26165 10845 26174
rect 10909 26165 10917 26174
rect 10977 26165 10989 26174
rect 11045 26165 11061 26174
rect 11113 26165 11133 26174
rect 11181 26165 11205 26174
rect 11249 26165 11277 26174
rect 11317 26165 11349 26174
rect 11385 26165 11419 26199
rect 11453 26174 11487 26199
rect 11521 26174 11555 26199
rect 11589 26174 11623 26199
rect 11657 26174 11691 26199
rect 11725 26174 11759 26199
rect 11793 26174 11827 26199
rect 11861 26174 11895 26199
rect 11929 26174 11963 26199
rect 11455 26165 11487 26174
rect 11527 26165 11555 26174
rect 11599 26165 11623 26174
rect 11671 26165 11691 26174
rect 11743 26165 11759 26174
rect 11815 26165 11827 26174
rect 11887 26165 11895 26174
rect 11959 26165 11963 26174
rect 11997 26174 12031 26199
rect 10807 26140 10845 26165
rect 10879 26140 10917 26165
rect 10951 26140 10989 26165
rect 11023 26140 11061 26165
rect 11095 26140 11133 26165
rect 11167 26140 11205 26165
rect 11239 26140 11277 26165
rect 11311 26140 11349 26165
rect 11383 26140 11421 26165
rect 11455 26140 11493 26165
rect 11527 26140 11565 26165
rect 11599 26140 11637 26165
rect 11671 26140 11709 26165
rect 11743 26140 11781 26165
rect 11815 26140 11853 26165
rect 11887 26140 11925 26165
rect 11959 26140 11997 26165
rect 12065 26174 12099 26199
rect 12133 26174 12167 26199
rect 12201 26174 12235 26199
rect 12269 26174 12303 26199
rect 12337 26174 12371 26199
rect 12405 26174 12439 26199
rect 12473 26174 12507 26199
rect 12541 26174 12575 26199
rect 12065 26165 12069 26174
rect 12133 26165 12141 26174
rect 12201 26165 12213 26174
rect 12269 26165 12285 26174
rect 12337 26165 12357 26174
rect 12405 26165 12429 26174
rect 12473 26165 12501 26174
rect 12541 26165 12573 26174
rect 12609 26165 12643 26199
rect 12677 26174 12711 26199
rect 12745 26174 12779 26199
rect 12813 26174 12847 26199
rect 12881 26174 12915 26199
rect 12949 26174 12983 26199
rect 13017 26174 13051 26199
rect 13085 26174 13119 26199
rect 13153 26174 13187 26199
rect 12679 26165 12711 26174
rect 12751 26165 12779 26174
rect 12823 26165 12847 26174
rect 12895 26165 12915 26174
rect 12967 26165 12983 26174
rect 13039 26165 13051 26174
rect 13111 26165 13119 26174
rect 13183 26165 13187 26174
rect 13221 26174 13255 26199
rect 12031 26140 12069 26165
rect 12103 26140 12141 26165
rect 12175 26140 12213 26165
rect 12247 26140 12285 26165
rect 12319 26140 12357 26165
rect 12391 26140 12429 26165
rect 12463 26140 12501 26165
rect 12535 26140 12573 26165
rect 12607 26140 12645 26165
rect 12679 26140 12717 26165
rect 12751 26140 12789 26165
rect 12823 26140 12861 26165
rect 12895 26140 12933 26165
rect 12967 26140 13005 26165
rect 13039 26140 13077 26165
rect 13111 26140 13149 26165
rect 13183 26140 13221 26165
rect 13289 26174 13323 26199
rect 13357 26174 13391 26199
rect 13425 26174 13459 26199
rect 13493 26174 13527 26199
rect 13561 26174 13595 26199
rect 13629 26174 13663 26199
rect 13289 26165 13293 26174
rect 13357 26165 13365 26174
rect 13425 26165 13437 26174
rect 13493 26165 13509 26174
rect 13561 26165 13581 26174
rect 13629 26165 13653 26174
rect 13697 26165 13731 26199
rect 13765 26175 13799 26199
rect 13833 26175 13867 26199
rect 13901 26175 13935 26199
rect 13790 26165 13799 26175
rect 13862 26165 13867 26175
rect 13934 26165 13935 26175
rect 13969 26175 14003 26199
rect 14037 26175 14071 26199
rect 14105 26175 14139 26199
rect 13969 26165 13972 26175
rect 14037 26165 14044 26175
rect 14105 26165 14116 26175
rect 14173 26165 14233 26199
rect 13255 26140 13293 26165
rect 13327 26140 13365 26165
rect 13399 26140 13437 26165
rect 13471 26140 13509 26165
rect 13543 26140 13581 26165
rect 13615 26140 13653 26165
rect 13687 26141 13756 26165
rect 13790 26141 13828 26165
rect 13862 26141 13900 26165
rect 13934 26141 13972 26165
rect 14006 26141 14044 26165
rect 14078 26141 14116 26165
rect 14150 26141 14233 26165
rect 13687 26140 14233 26141
rect 9877 26129 14233 26140
rect 9877 26100 9911 26129
rect 9877 26066 9909 26100
rect 9945 26095 9980 26129
rect 10014 26100 10049 26129
rect 10083 26100 10118 26129
rect 10152 26100 10187 26129
rect 10221 26100 10256 26129
rect 10290 26100 10325 26129
rect 10359 26100 10394 26129
rect 10428 26100 10463 26129
rect 10497 26100 10532 26129
rect 10566 26100 10601 26129
rect 10635 26100 10670 26129
rect 10704 26100 10739 26129
rect 10015 26095 10049 26100
rect 10087 26095 10118 26100
rect 10159 26095 10187 26100
rect 10231 26095 10256 26100
rect 10303 26095 10325 26100
rect 10375 26095 10394 26100
rect 10447 26095 10463 26100
rect 10519 26095 10532 26100
rect 10591 26095 10601 26100
rect 10663 26095 10670 26100
rect 10735 26095 10739 26100
rect 10773 26100 10807 26129
rect 9943 26066 9981 26095
rect 10015 26066 10053 26095
rect 10087 26066 10125 26095
rect 10159 26066 10197 26095
rect 10231 26066 10269 26095
rect 10303 26066 10341 26095
rect 10375 26066 10413 26095
rect 10447 26066 10485 26095
rect 10519 26066 10557 26095
rect 10591 26066 10629 26095
rect 10663 26066 10701 26095
rect 10735 26066 10773 26095
rect 10841 26100 10875 26129
rect 10909 26100 10943 26129
rect 10977 26100 11011 26129
rect 11045 26100 11079 26129
rect 11113 26100 11147 26129
rect 11181 26100 11215 26129
rect 11249 26100 11283 26129
rect 11317 26100 11351 26129
rect 10841 26095 10845 26100
rect 10909 26095 10917 26100
rect 10977 26095 10989 26100
rect 11045 26095 11061 26100
rect 11113 26095 11133 26100
rect 11181 26095 11205 26100
rect 11249 26095 11277 26100
rect 11317 26095 11349 26100
rect 11385 26095 11419 26129
rect 11453 26100 11487 26129
rect 11521 26100 11555 26129
rect 11589 26100 11623 26129
rect 11657 26100 11691 26129
rect 11725 26100 11759 26129
rect 11793 26100 11827 26129
rect 11861 26100 11895 26129
rect 11929 26100 11963 26129
rect 11455 26095 11487 26100
rect 11527 26095 11555 26100
rect 11599 26095 11623 26100
rect 11671 26095 11691 26100
rect 11743 26095 11759 26100
rect 11815 26095 11827 26100
rect 11887 26095 11895 26100
rect 11959 26095 11963 26100
rect 11997 26100 12031 26129
rect 10807 26066 10845 26095
rect 10879 26066 10917 26095
rect 10951 26066 10989 26095
rect 11023 26066 11061 26095
rect 11095 26066 11133 26095
rect 11167 26066 11205 26095
rect 11239 26066 11277 26095
rect 11311 26066 11349 26095
rect 11383 26066 11421 26095
rect 11455 26066 11493 26095
rect 11527 26066 11565 26095
rect 11599 26066 11637 26095
rect 11671 26066 11709 26095
rect 11743 26066 11781 26095
rect 11815 26066 11853 26095
rect 11887 26066 11925 26095
rect 11959 26066 11997 26095
rect 12065 26100 12099 26129
rect 12133 26100 12167 26129
rect 12201 26100 12235 26129
rect 12269 26100 12303 26129
rect 12337 26100 12371 26129
rect 12405 26100 12439 26129
rect 12473 26100 12507 26129
rect 12541 26100 12575 26129
rect 12065 26095 12069 26100
rect 12133 26095 12141 26100
rect 12201 26095 12213 26100
rect 12269 26095 12285 26100
rect 12337 26095 12357 26100
rect 12405 26095 12429 26100
rect 12473 26095 12501 26100
rect 12541 26095 12573 26100
rect 12609 26095 12643 26129
rect 12677 26100 12711 26129
rect 12745 26100 12779 26129
rect 12813 26100 12847 26129
rect 12881 26100 12915 26129
rect 12949 26100 12983 26129
rect 13017 26100 13051 26129
rect 13085 26100 13119 26129
rect 13153 26100 13187 26129
rect 12679 26095 12711 26100
rect 12751 26095 12779 26100
rect 12823 26095 12847 26100
rect 12895 26095 12915 26100
rect 12967 26095 12983 26100
rect 13039 26095 13051 26100
rect 13111 26095 13119 26100
rect 13183 26095 13187 26100
rect 13221 26100 13255 26129
rect 12031 26066 12069 26095
rect 12103 26066 12141 26095
rect 12175 26066 12213 26095
rect 12247 26066 12285 26095
rect 12319 26066 12357 26095
rect 12391 26066 12429 26095
rect 12463 26066 12501 26095
rect 12535 26066 12573 26095
rect 12607 26066 12645 26095
rect 12679 26066 12717 26095
rect 12751 26066 12789 26095
rect 12823 26066 12861 26095
rect 12895 26066 12933 26095
rect 12967 26066 13005 26095
rect 13039 26066 13077 26095
rect 13111 26066 13149 26095
rect 13183 26066 13221 26095
rect 13289 26100 13323 26129
rect 13357 26100 13391 26129
rect 13425 26100 13459 26129
rect 13493 26100 13527 26129
rect 13561 26100 13595 26129
rect 13629 26100 13663 26129
rect 13289 26095 13293 26100
rect 13357 26095 13365 26100
rect 13425 26095 13437 26100
rect 13493 26095 13509 26100
rect 13561 26095 13581 26100
rect 13629 26095 13653 26100
rect 13697 26095 13731 26129
rect 13765 26102 13799 26129
rect 13833 26102 13867 26129
rect 13901 26102 13935 26129
rect 13790 26095 13799 26102
rect 13862 26095 13867 26102
rect 13934 26095 13935 26102
rect 13969 26102 14003 26129
rect 14037 26102 14071 26129
rect 14105 26102 14139 26129
rect 13969 26095 13972 26102
rect 14037 26095 14044 26102
rect 14105 26095 14116 26102
rect 14173 26095 14233 26129
rect 13255 26066 13293 26095
rect 13327 26066 13365 26095
rect 13399 26066 13437 26095
rect 13471 26066 13509 26095
rect 13543 26066 13581 26095
rect 13615 26066 13653 26095
rect 13687 26068 13756 26095
rect 13790 26068 13828 26095
rect 13862 26068 13900 26095
rect 13934 26068 13972 26095
rect 14006 26068 14044 26095
rect 14078 26068 14116 26095
rect 14150 26068 14233 26095
rect 13687 26066 14233 26068
rect 9877 26059 14233 26066
rect 9877 26026 9911 26059
rect 9877 25992 9909 26026
rect 9945 26025 9980 26059
rect 10014 26026 10049 26059
rect 10083 26026 10118 26059
rect 10152 26026 10187 26059
rect 10221 26026 10256 26059
rect 10290 26026 10325 26059
rect 10359 26026 10394 26059
rect 10428 26026 10463 26059
rect 10497 26026 10532 26059
rect 10566 26026 10601 26059
rect 10635 26026 10670 26059
rect 10704 26026 10739 26059
rect 10015 26025 10049 26026
rect 10087 26025 10118 26026
rect 10159 26025 10187 26026
rect 10231 26025 10256 26026
rect 10303 26025 10325 26026
rect 10375 26025 10394 26026
rect 10447 26025 10463 26026
rect 10519 26025 10532 26026
rect 10591 26025 10601 26026
rect 10663 26025 10670 26026
rect 10735 26025 10739 26026
rect 10773 26026 10807 26059
rect 9943 25992 9981 26025
rect 10015 25992 10053 26025
rect 10087 25992 10125 26025
rect 10159 25992 10197 26025
rect 10231 25992 10269 26025
rect 10303 25992 10341 26025
rect 10375 25992 10413 26025
rect 10447 25992 10485 26025
rect 10519 25992 10557 26025
rect 10591 25992 10629 26025
rect 10663 25992 10701 26025
rect 10735 25992 10773 26025
rect 10841 26026 10875 26059
rect 10909 26026 10943 26059
rect 10977 26026 11011 26059
rect 11045 26026 11079 26059
rect 11113 26026 11147 26059
rect 11181 26026 11215 26059
rect 11249 26026 11283 26059
rect 11317 26026 11351 26059
rect 10841 26025 10845 26026
rect 10909 26025 10917 26026
rect 10977 26025 10989 26026
rect 11045 26025 11061 26026
rect 11113 26025 11133 26026
rect 11181 26025 11205 26026
rect 11249 26025 11277 26026
rect 11317 26025 11349 26026
rect 11385 26025 11419 26059
rect 11453 26026 11487 26059
rect 11521 26026 11555 26059
rect 11589 26026 11623 26059
rect 11657 26026 11691 26059
rect 11725 26026 11759 26059
rect 11793 26026 11827 26059
rect 11861 26026 11895 26059
rect 11929 26026 11963 26059
rect 11455 26025 11487 26026
rect 11527 26025 11555 26026
rect 11599 26025 11623 26026
rect 11671 26025 11691 26026
rect 11743 26025 11759 26026
rect 11815 26025 11827 26026
rect 11887 26025 11895 26026
rect 11959 26025 11963 26026
rect 11997 26026 12031 26059
rect 10807 25992 10845 26025
rect 10879 25992 10917 26025
rect 10951 25992 10989 26025
rect 11023 25992 11061 26025
rect 11095 25992 11133 26025
rect 11167 25992 11205 26025
rect 11239 25992 11277 26025
rect 11311 25992 11349 26025
rect 11383 25992 11421 26025
rect 11455 25992 11493 26025
rect 11527 25992 11565 26025
rect 11599 25992 11637 26025
rect 11671 25992 11709 26025
rect 11743 25992 11781 26025
rect 11815 25992 11853 26025
rect 11887 25992 11925 26025
rect 11959 25992 11997 26025
rect 12065 26026 12099 26059
rect 12133 26026 12167 26059
rect 12201 26026 12235 26059
rect 12269 26026 12303 26059
rect 12337 26026 12371 26059
rect 12405 26026 12439 26059
rect 12473 26026 12507 26059
rect 12541 26026 12575 26059
rect 12065 26025 12069 26026
rect 12133 26025 12141 26026
rect 12201 26025 12213 26026
rect 12269 26025 12285 26026
rect 12337 26025 12357 26026
rect 12405 26025 12429 26026
rect 12473 26025 12501 26026
rect 12541 26025 12573 26026
rect 12609 26025 12643 26059
rect 12677 26026 12711 26059
rect 12745 26026 12779 26059
rect 12813 26026 12847 26059
rect 12881 26026 12915 26059
rect 12949 26026 12983 26059
rect 13017 26026 13051 26059
rect 13085 26026 13119 26059
rect 13153 26026 13187 26059
rect 12679 26025 12711 26026
rect 12751 26025 12779 26026
rect 12823 26025 12847 26026
rect 12895 26025 12915 26026
rect 12967 26025 12983 26026
rect 13039 26025 13051 26026
rect 13111 26025 13119 26026
rect 13183 26025 13187 26026
rect 13221 26026 13255 26059
rect 12031 25992 12069 26025
rect 12103 25992 12141 26025
rect 12175 25992 12213 26025
rect 12247 25992 12285 26025
rect 12319 25992 12357 26025
rect 12391 25992 12429 26025
rect 12463 25992 12501 26025
rect 12535 25992 12573 26025
rect 12607 25992 12645 26025
rect 12679 25992 12717 26025
rect 12751 25992 12789 26025
rect 12823 25992 12861 26025
rect 12895 25992 12933 26025
rect 12967 25992 13005 26025
rect 13039 25992 13077 26025
rect 13111 25992 13149 26025
rect 13183 25992 13221 26025
rect 13289 26026 13323 26059
rect 13357 26026 13391 26059
rect 13425 26026 13459 26059
rect 13493 26026 13527 26059
rect 13561 26026 13595 26059
rect 13629 26026 13663 26059
rect 13289 26025 13293 26026
rect 13357 26025 13365 26026
rect 13425 26025 13437 26026
rect 13493 26025 13509 26026
rect 13561 26025 13581 26026
rect 13629 26025 13653 26026
rect 13697 26025 13731 26059
rect 13765 26029 13799 26059
rect 13833 26029 13867 26059
rect 13901 26029 13935 26059
rect 13790 26025 13799 26029
rect 13862 26025 13867 26029
rect 13934 26025 13935 26029
rect 13969 26029 14003 26059
rect 14037 26029 14071 26059
rect 14105 26029 14139 26059
rect 13969 26025 13972 26029
rect 14037 26025 14044 26029
rect 14105 26025 14116 26029
rect 14173 26025 14233 26059
rect 13255 25992 13293 26025
rect 13327 25992 13365 26025
rect 13399 25992 13437 26025
rect 13471 25992 13509 26025
rect 13543 25992 13581 26025
rect 13615 25992 13653 26025
rect 13687 25995 13756 26025
rect 13790 25995 13828 26025
rect 13862 25995 13900 26025
rect 13934 25995 13972 26025
rect 14006 25995 14044 26025
rect 14078 25995 14116 26025
rect 14150 25995 14233 26025
rect 13687 25992 14233 25995
rect 9877 25989 14233 25992
rect 9877 25955 9911 25989
rect 9945 25955 9980 25989
rect 10014 25955 10049 25989
rect 10083 25955 10118 25989
rect 10152 25955 10187 25989
rect 10221 25955 10256 25989
rect 10290 25955 10325 25989
rect 10359 25955 10394 25989
rect 10428 25955 10463 25989
rect 10497 25955 10532 25989
rect 10566 25955 10601 25989
rect 10635 25955 10670 25989
rect 10704 25955 10739 25989
rect 10773 25955 10807 25989
rect 10841 25955 10875 25989
rect 10909 25955 10943 25989
rect 10977 25955 11011 25989
rect 11045 25955 11079 25989
rect 11113 25955 11147 25989
rect 11181 25955 11215 25989
rect 11249 25955 11283 25989
rect 11317 25955 11351 25989
rect 11385 25955 11419 25989
rect 11453 25955 11487 25989
rect 11521 25955 11555 25989
rect 11589 25955 11623 25989
rect 11657 25955 11691 25989
rect 11725 25955 11759 25989
rect 11793 25955 11827 25989
rect 11861 25955 11895 25989
rect 11929 25955 11963 25989
rect 11997 25955 12031 25989
rect 12065 25955 12099 25989
rect 12133 25955 12167 25989
rect 12201 25955 12235 25989
rect 12269 25955 12303 25989
rect 12337 25955 12371 25989
rect 12405 25955 12439 25989
rect 12473 25955 12507 25989
rect 12541 25955 12575 25989
rect 12609 25955 12643 25989
rect 12677 25955 12711 25989
rect 12745 25955 12779 25989
rect 12813 25955 12847 25989
rect 12881 25955 12915 25989
rect 12949 25955 12983 25989
rect 13017 25955 13051 25989
rect 13085 25955 13119 25989
rect 13153 25955 13187 25989
rect 13221 25955 13255 25989
rect 13289 25955 13323 25989
rect 13357 25955 13391 25989
rect 13425 25955 13459 25989
rect 13493 25955 13527 25989
rect 13561 25955 13595 25989
rect 13629 25955 13663 25989
rect 13697 25955 13731 25989
rect 13765 25955 13799 25989
rect 13833 25955 13867 25989
rect 13901 25955 13935 25989
rect 13969 25955 14003 25989
rect 14037 25955 14071 25989
rect 14105 25955 14139 25989
rect 14173 25955 14233 25989
rect 9877 25953 13756 25955
rect 9877 25919 9909 25953
rect 9943 25919 9981 25953
rect 10015 25919 10053 25953
rect 10087 25919 10125 25953
rect 10159 25919 10197 25953
rect 10231 25919 10269 25953
rect 10303 25919 10341 25953
rect 10375 25919 10413 25953
rect 10447 25919 10485 25953
rect 10519 25919 10557 25953
rect 10591 25919 10629 25953
rect 10663 25919 10701 25953
rect 10735 25919 10773 25953
rect 10807 25919 10845 25953
rect 10879 25919 10917 25953
rect 10951 25919 10989 25953
rect 11023 25919 11061 25953
rect 11095 25919 11133 25953
rect 11167 25919 11205 25953
rect 11239 25919 11277 25953
rect 11311 25919 11349 25953
rect 11383 25919 11421 25953
rect 11455 25919 11493 25953
rect 11527 25919 11565 25953
rect 11599 25919 11637 25953
rect 11671 25919 11709 25953
rect 11743 25919 11781 25953
rect 11815 25919 11853 25953
rect 11887 25919 11925 25953
rect 11959 25919 11997 25953
rect 12031 25919 12069 25953
rect 12103 25919 12141 25953
rect 12175 25919 12213 25953
rect 12247 25919 12285 25953
rect 12319 25919 12357 25953
rect 12391 25919 12429 25953
rect 12463 25919 12501 25953
rect 12535 25919 12573 25953
rect 12607 25919 12645 25953
rect 12679 25919 12717 25953
rect 12751 25919 12789 25953
rect 12823 25919 12861 25953
rect 12895 25919 12933 25953
rect 12967 25919 13005 25953
rect 13039 25919 13077 25953
rect 13111 25919 13149 25953
rect 13183 25919 13221 25953
rect 13255 25919 13293 25953
rect 13327 25919 13365 25953
rect 13399 25919 13437 25953
rect 13471 25919 13509 25953
rect 13543 25919 13581 25953
rect 13615 25919 13653 25953
rect 13687 25921 13756 25953
rect 13790 25921 13828 25955
rect 13862 25921 13900 25955
rect 13934 25921 13972 25955
rect 14006 25921 14044 25955
rect 14078 25921 14116 25955
rect 14150 25921 14233 25955
rect 13687 25919 14233 25921
rect 9877 25885 9911 25919
rect 9945 25885 9980 25919
rect 10014 25885 10049 25919
rect 10083 25885 10118 25919
rect 10152 25885 10187 25919
rect 10221 25885 10256 25919
rect 10290 25885 10325 25919
rect 10359 25885 10394 25919
rect 10428 25885 10463 25919
rect 10497 25885 10532 25919
rect 10566 25885 10601 25919
rect 10635 25885 10670 25919
rect 10704 25885 10739 25919
rect 10773 25885 10807 25919
rect 10841 25885 10875 25919
rect 10909 25885 10943 25919
rect 10977 25885 11011 25919
rect 11045 25885 11079 25919
rect 11113 25885 11147 25919
rect 11181 25885 11215 25919
rect 11249 25885 11283 25919
rect 11317 25885 11351 25919
rect 11385 25885 11419 25919
rect 11453 25885 11487 25919
rect 11521 25885 11555 25919
rect 11589 25885 11623 25919
rect 11657 25885 11691 25919
rect 11725 25885 11759 25919
rect 11793 25885 11827 25919
rect 11861 25885 11895 25919
rect 11929 25885 11963 25919
rect 11997 25885 12031 25919
rect 12065 25885 12099 25919
rect 12133 25885 12167 25919
rect 12201 25885 12235 25919
rect 12269 25885 12303 25919
rect 12337 25885 12371 25919
rect 12405 25885 12439 25919
rect 12473 25885 12507 25919
rect 12541 25885 12575 25919
rect 12609 25885 12643 25919
rect 12677 25885 12711 25919
rect 12745 25885 12779 25919
rect 12813 25885 12847 25919
rect 12881 25885 12915 25919
rect 12949 25885 12983 25919
rect 13017 25885 13051 25919
rect 13085 25885 13119 25919
rect 13153 25885 13187 25919
rect 13221 25885 13255 25919
rect 13289 25885 13323 25919
rect 13357 25885 13391 25919
rect 13425 25885 13459 25919
rect 13493 25885 13527 25919
rect 13561 25885 13595 25919
rect 13629 25885 13663 25919
rect 13697 25885 13731 25919
rect 13765 25885 13799 25919
rect 13833 25885 13867 25919
rect 13901 25885 13935 25919
rect 13969 25885 14003 25919
rect 14037 25885 14071 25919
rect 14105 25885 14139 25919
rect 14173 25885 14233 25919
rect 9877 25881 14233 25885
rect 9877 25880 13756 25881
rect 9877 25846 9909 25880
rect 9943 25849 9981 25880
rect 10015 25849 10053 25880
rect 10087 25849 10125 25880
rect 10159 25849 10197 25880
rect 10231 25849 10269 25880
rect 10303 25849 10341 25880
rect 10375 25849 10413 25880
rect 10447 25849 10485 25880
rect 10519 25849 10557 25880
rect 10591 25849 10629 25880
rect 10663 25849 10701 25880
rect 10735 25849 10773 25880
rect 9877 25815 9911 25846
rect 9945 25815 9980 25849
rect 10015 25846 10049 25849
rect 10087 25846 10118 25849
rect 10159 25846 10187 25849
rect 10231 25846 10256 25849
rect 10303 25846 10325 25849
rect 10375 25846 10394 25849
rect 10447 25846 10463 25849
rect 10519 25846 10532 25849
rect 10591 25846 10601 25849
rect 10663 25846 10670 25849
rect 10735 25846 10739 25849
rect 10014 25815 10049 25846
rect 10083 25815 10118 25846
rect 10152 25815 10187 25846
rect 10221 25815 10256 25846
rect 10290 25815 10325 25846
rect 10359 25815 10394 25846
rect 10428 25815 10463 25846
rect 10497 25815 10532 25846
rect 10566 25815 10601 25846
rect 10635 25815 10670 25846
rect 10704 25815 10739 25846
rect 10807 25849 10845 25880
rect 10879 25849 10917 25880
rect 10951 25849 10989 25880
rect 11023 25849 11061 25880
rect 11095 25849 11133 25880
rect 11167 25849 11205 25880
rect 11239 25849 11277 25880
rect 11311 25849 11349 25880
rect 11383 25849 11421 25880
rect 11455 25849 11493 25880
rect 11527 25849 11565 25880
rect 11599 25849 11637 25880
rect 11671 25849 11709 25880
rect 11743 25849 11781 25880
rect 11815 25849 11853 25880
rect 11887 25849 11925 25880
rect 11959 25849 11997 25880
rect 10773 25815 10807 25846
rect 10841 25846 10845 25849
rect 10909 25846 10917 25849
rect 10977 25846 10989 25849
rect 11045 25846 11061 25849
rect 11113 25846 11133 25849
rect 11181 25846 11205 25849
rect 11249 25846 11277 25849
rect 11317 25846 11349 25849
rect 10841 25815 10875 25846
rect 10909 25815 10943 25846
rect 10977 25815 11011 25846
rect 11045 25815 11079 25846
rect 11113 25815 11147 25846
rect 11181 25815 11215 25846
rect 11249 25815 11283 25846
rect 11317 25815 11351 25846
rect 11385 25815 11419 25849
rect 11455 25846 11487 25849
rect 11527 25846 11555 25849
rect 11599 25846 11623 25849
rect 11671 25846 11691 25849
rect 11743 25846 11759 25849
rect 11815 25846 11827 25849
rect 11887 25846 11895 25849
rect 11959 25846 11963 25849
rect 11453 25815 11487 25846
rect 11521 25815 11555 25846
rect 11589 25815 11623 25846
rect 11657 25815 11691 25846
rect 11725 25815 11759 25846
rect 11793 25815 11827 25846
rect 11861 25815 11895 25846
rect 11929 25815 11963 25846
rect 12031 25849 12069 25880
rect 12103 25849 12141 25880
rect 12175 25849 12213 25880
rect 12247 25849 12285 25880
rect 12319 25849 12357 25880
rect 12391 25849 12429 25880
rect 12463 25849 12501 25880
rect 12535 25849 12573 25880
rect 12607 25849 12645 25880
rect 12679 25849 12717 25880
rect 12751 25849 12789 25880
rect 12823 25849 12861 25880
rect 12895 25849 12933 25880
rect 12967 25849 13005 25880
rect 13039 25849 13077 25880
rect 13111 25849 13149 25880
rect 13183 25849 13221 25880
rect 11997 25815 12031 25846
rect 12065 25846 12069 25849
rect 12133 25846 12141 25849
rect 12201 25846 12213 25849
rect 12269 25846 12285 25849
rect 12337 25846 12357 25849
rect 12405 25846 12429 25849
rect 12473 25846 12501 25849
rect 12541 25846 12573 25849
rect 12065 25815 12099 25846
rect 12133 25815 12167 25846
rect 12201 25815 12235 25846
rect 12269 25815 12303 25846
rect 12337 25815 12371 25846
rect 12405 25815 12439 25846
rect 12473 25815 12507 25846
rect 12541 25815 12575 25846
rect 12609 25815 12643 25849
rect 12679 25846 12711 25849
rect 12751 25846 12779 25849
rect 12823 25846 12847 25849
rect 12895 25846 12915 25849
rect 12967 25846 12983 25849
rect 13039 25846 13051 25849
rect 13111 25846 13119 25849
rect 13183 25846 13187 25849
rect 12677 25815 12711 25846
rect 12745 25815 12779 25846
rect 12813 25815 12847 25846
rect 12881 25815 12915 25846
rect 12949 25815 12983 25846
rect 13017 25815 13051 25846
rect 13085 25815 13119 25846
rect 13153 25815 13187 25846
rect 13255 25849 13293 25880
rect 13327 25849 13365 25880
rect 13399 25849 13437 25880
rect 13471 25849 13509 25880
rect 13543 25849 13581 25880
rect 13615 25849 13653 25880
rect 13687 25849 13756 25880
rect 13790 25849 13828 25881
rect 13862 25849 13900 25881
rect 13934 25849 13972 25881
rect 14006 25849 14044 25881
rect 14078 25849 14116 25881
rect 14150 25849 14233 25881
rect 13221 25815 13255 25846
rect 13289 25846 13293 25849
rect 13357 25846 13365 25849
rect 13425 25846 13437 25849
rect 13493 25846 13509 25849
rect 13561 25846 13581 25849
rect 13629 25846 13653 25849
rect 13289 25815 13323 25846
rect 13357 25815 13391 25846
rect 13425 25815 13459 25846
rect 13493 25815 13527 25846
rect 13561 25815 13595 25846
rect 13629 25815 13663 25846
rect 13697 25815 13731 25849
rect 13790 25847 13799 25849
rect 13862 25847 13867 25849
rect 13934 25847 13935 25849
rect 13765 25815 13799 25847
rect 13833 25815 13867 25847
rect 13901 25815 13935 25847
rect 13969 25847 13972 25849
rect 14037 25847 14044 25849
rect 14105 25847 14116 25849
rect 13969 25815 14003 25847
rect 14037 25815 14071 25847
rect 14105 25815 14139 25847
rect 14173 25815 14233 25849
rect 9877 25807 14233 25815
rect 9877 25773 9909 25807
rect 9943 25779 9981 25807
rect 10015 25779 10053 25807
rect 10087 25779 10125 25807
rect 10159 25779 10197 25807
rect 10231 25779 10269 25807
rect 10303 25779 10341 25807
rect 10375 25779 10413 25807
rect 10447 25779 10485 25807
rect 10519 25779 10557 25807
rect 10591 25779 10629 25807
rect 10663 25779 10701 25807
rect 10735 25779 10773 25807
rect 9877 25745 9911 25773
rect 9945 25745 9980 25779
rect 10015 25773 10049 25779
rect 10087 25773 10118 25779
rect 10159 25773 10187 25779
rect 10231 25773 10256 25779
rect 10303 25773 10325 25779
rect 10375 25773 10394 25779
rect 10447 25773 10463 25779
rect 10519 25773 10532 25779
rect 10591 25773 10601 25779
rect 10663 25773 10670 25779
rect 10735 25773 10739 25779
rect 10014 25745 10049 25773
rect 10083 25745 10118 25773
rect 10152 25745 10187 25773
rect 10221 25745 10256 25773
rect 10290 25745 10325 25773
rect 10359 25745 10394 25773
rect 10428 25745 10463 25773
rect 10497 25745 10532 25773
rect 10566 25745 10601 25773
rect 10635 25745 10670 25773
rect 10704 25745 10739 25773
rect 10807 25779 10845 25807
rect 10879 25779 10917 25807
rect 10951 25779 10989 25807
rect 11023 25779 11061 25807
rect 11095 25779 11133 25807
rect 11167 25779 11205 25807
rect 11239 25779 11277 25807
rect 11311 25779 11349 25807
rect 11383 25779 11421 25807
rect 11455 25779 11493 25807
rect 11527 25779 11565 25807
rect 11599 25779 11637 25807
rect 11671 25779 11709 25807
rect 11743 25779 11781 25807
rect 11815 25779 11853 25807
rect 11887 25779 11925 25807
rect 11959 25779 11997 25807
rect 10773 25745 10807 25773
rect 10841 25773 10845 25779
rect 10909 25773 10917 25779
rect 10977 25773 10989 25779
rect 11045 25773 11061 25779
rect 11113 25773 11133 25779
rect 11181 25773 11205 25779
rect 11249 25773 11277 25779
rect 11317 25773 11349 25779
rect 10841 25745 10875 25773
rect 10909 25745 10943 25773
rect 10977 25745 11011 25773
rect 11045 25745 11079 25773
rect 11113 25745 11147 25773
rect 11181 25745 11215 25773
rect 11249 25745 11283 25773
rect 11317 25745 11351 25773
rect 11385 25745 11419 25779
rect 11455 25773 11487 25779
rect 11527 25773 11555 25779
rect 11599 25773 11623 25779
rect 11671 25773 11691 25779
rect 11743 25773 11759 25779
rect 11815 25773 11827 25779
rect 11887 25773 11895 25779
rect 11959 25773 11963 25779
rect 11453 25745 11487 25773
rect 11521 25745 11555 25773
rect 11589 25745 11623 25773
rect 11657 25745 11691 25773
rect 11725 25745 11759 25773
rect 11793 25745 11827 25773
rect 11861 25745 11895 25773
rect 11929 25745 11963 25773
rect 12031 25779 12069 25807
rect 12103 25779 12141 25807
rect 12175 25779 12213 25807
rect 12247 25779 12285 25807
rect 12319 25779 12357 25807
rect 12391 25779 12429 25807
rect 12463 25779 12501 25807
rect 12535 25779 12573 25807
rect 12607 25779 12645 25807
rect 12679 25779 12717 25807
rect 12751 25779 12789 25807
rect 12823 25779 12861 25807
rect 12895 25779 12933 25807
rect 12967 25779 13005 25807
rect 13039 25779 13077 25807
rect 13111 25779 13149 25807
rect 13183 25779 13221 25807
rect 11997 25745 12031 25773
rect 12065 25773 12069 25779
rect 12133 25773 12141 25779
rect 12201 25773 12213 25779
rect 12269 25773 12285 25779
rect 12337 25773 12357 25779
rect 12405 25773 12429 25779
rect 12473 25773 12501 25779
rect 12541 25773 12573 25779
rect 12065 25745 12099 25773
rect 12133 25745 12167 25773
rect 12201 25745 12235 25773
rect 12269 25745 12303 25773
rect 12337 25745 12371 25773
rect 12405 25745 12439 25773
rect 12473 25745 12507 25773
rect 12541 25745 12575 25773
rect 12609 25745 12643 25779
rect 12679 25773 12711 25779
rect 12751 25773 12779 25779
rect 12823 25773 12847 25779
rect 12895 25773 12915 25779
rect 12967 25773 12983 25779
rect 13039 25773 13051 25779
rect 13111 25773 13119 25779
rect 13183 25773 13187 25779
rect 12677 25745 12711 25773
rect 12745 25745 12779 25773
rect 12813 25745 12847 25773
rect 12881 25745 12915 25773
rect 12949 25745 12983 25773
rect 13017 25745 13051 25773
rect 13085 25745 13119 25773
rect 13153 25745 13187 25773
rect 13255 25779 13293 25807
rect 13327 25779 13365 25807
rect 13399 25779 13437 25807
rect 13471 25779 13509 25807
rect 13543 25779 13581 25807
rect 13615 25779 13653 25807
rect 13687 25779 13756 25807
rect 13790 25779 13828 25807
rect 13862 25779 13900 25807
rect 13934 25779 13972 25807
rect 14006 25779 14044 25807
rect 14078 25779 14116 25807
rect 14150 25779 14233 25807
rect 13221 25745 13255 25773
rect 13289 25773 13293 25779
rect 13357 25773 13365 25779
rect 13425 25773 13437 25779
rect 13493 25773 13509 25779
rect 13561 25773 13581 25779
rect 13629 25773 13653 25779
rect 13289 25745 13323 25773
rect 13357 25745 13391 25773
rect 13425 25745 13459 25773
rect 13493 25745 13527 25773
rect 13561 25745 13595 25773
rect 13629 25745 13663 25773
rect 13697 25745 13731 25779
rect 13790 25773 13799 25779
rect 13862 25773 13867 25779
rect 13934 25773 13935 25779
rect 13765 25745 13799 25773
rect 13833 25745 13867 25773
rect 13901 25745 13935 25773
rect 13969 25773 13972 25779
rect 14037 25773 14044 25779
rect 14105 25773 14116 25779
rect 13969 25745 14003 25773
rect 14037 25745 14071 25773
rect 14105 25745 14139 25773
rect 14173 25745 14233 25779
rect 9877 25734 14233 25745
rect 9877 25700 9909 25734
rect 9943 25709 9981 25734
rect 10015 25709 10053 25734
rect 10087 25709 10125 25734
rect 10159 25709 10197 25734
rect 10231 25709 10269 25734
rect 10303 25709 10341 25734
rect 10375 25709 10413 25734
rect 10447 25709 10485 25734
rect 10519 25709 10557 25734
rect 10591 25709 10629 25734
rect 10663 25709 10701 25734
rect 10735 25709 10773 25734
rect 9877 25675 9911 25700
rect 9945 25675 9980 25709
rect 10015 25700 10049 25709
rect 10087 25700 10118 25709
rect 10159 25700 10187 25709
rect 10231 25700 10256 25709
rect 10303 25700 10325 25709
rect 10375 25700 10394 25709
rect 10447 25700 10463 25709
rect 10519 25700 10532 25709
rect 10591 25700 10601 25709
rect 10663 25700 10670 25709
rect 10735 25700 10739 25709
rect 10014 25675 10049 25700
rect 10083 25675 10118 25700
rect 10152 25675 10187 25700
rect 10221 25675 10256 25700
rect 10290 25675 10325 25700
rect 10359 25675 10394 25700
rect 10428 25675 10463 25700
rect 10497 25675 10532 25700
rect 10566 25675 10601 25700
rect 10635 25675 10670 25700
rect 10704 25675 10739 25700
rect 10807 25709 10845 25734
rect 10879 25709 10917 25734
rect 10951 25709 10989 25734
rect 11023 25709 11061 25734
rect 11095 25709 11133 25734
rect 11167 25709 11205 25734
rect 11239 25709 11277 25734
rect 11311 25709 11349 25734
rect 11383 25709 11421 25734
rect 11455 25709 11493 25734
rect 11527 25709 11565 25734
rect 11599 25709 11637 25734
rect 11671 25709 11709 25734
rect 11743 25709 11781 25734
rect 11815 25709 11853 25734
rect 11887 25709 11925 25734
rect 11959 25709 11997 25734
rect 10773 25675 10807 25700
rect 10841 25700 10845 25709
rect 10909 25700 10917 25709
rect 10977 25700 10989 25709
rect 11045 25700 11061 25709
rect 11113 25700 11133 25709
rect 11181 25700 11205 25709
rect 11249 25700 11277 25709
rect 11317 25700 11349 25709
rect 10841 25675 10875 25700
rect 10909 25675 10943 25700
rect 10977 25675 11011 25700
rect 11045 25675 11079 25700
rect 11113 25675 11147 25700
rect 11181 25675 11215 25700
rect 11249 25675 11283 25700
rect 11317 25675 11351 25700
rect 11385 25675 11419 25709
rect 11455 25700 11487 25709
rect 11527 25700 11555 25709
rect 11599 25700 11623 25709
rect 11671 25700 11691 25709
rect 11743 25700 11759 25709
rect 11815 25700 11827 25709
rect 11887 25700 11895 25709
rect 11959 25700 11963 25709
rect 11453 25675 11487 25700
rect 11521 25675 11555 25700
rect 11589 25675 11623 25700
rect 11657 25675 11691 25700
rect 11725 25675 11759 25700
rect 11793 25675 11827 25700
rect 11861 25675 11895 25700
rect 11929 25675 11963 25700
rect 12031 25709 12069 25734
rect 12103 25709 12141 25734
rect 12175 25709 12213 25734
rect 12247 25709 12285 25734
rect 12319 25709 12357 25734
rect 12391 25709 12429 25734
rect 12463 25709 12501 25734
rect 12535 25709 12573 25734
rect 12607 25709 12645 25734
rect 12679 25709 12717 25734
rect 12751 25709 12789 25734
rect 12823 25709 12861 25734
rect 12895 25709 12933 25734
rect 12967 25709 13005 25734
rect 13039 25709 13077 25734
rect 13111 25709 13149 25734
rect 13183 25709 13221 25734
rect 11997 25675 12031 25700
rect 12065 25700 12069 25709
rect 12133 25700 12141 25709
rect 12201 25700 12213 25709
rect 12269 25700 12285 25709
rect 12337 25700 12357 25709
rect 12405 25700 12429 25709
rect 12473 25700 12501 25709
rect 12541 25700 12573 25709
rect 12065 25675 12099 25700
rect 12133 25675 12167 25700
rect 12201 25675 12235 25700
rect 12269 25675 12303 25700
rect 12337 25675 12371 25700
rect 12405 25675 12439 25700
rect 12473 25675 12507 25700
rect 12541 25675 12575 25700
rect 12609 25675 12643 25709
rect 12679 25700 12711 25709
rect 12751 25700 12779 25709
rect 12823 25700 12847 25709
rect 12895 25700 12915 25709
rect 12967 25700 12983 25709
rect 13039 25700 13051 25709
rect 13111 25700 13119 25709
rect 13183 25700 13187 25709
rect 12677 25675 12711 25700
rect 12745 25675 12779 25700
rect 12813 25675 12847 25700
rect 12881 25675 12915 25700
rect 12949 25675 12983 25700
rect 13017 25675 13051 25700
rect 13085 25675 13119 25700
rect 13153 25675 13187 25700
rect 13255 25709 13293 25734
rect 13327 25709 13365 25734
rect 13399 25709 13437 25734
rect 13471 25709 13509 25734
rect 13543 25709 13581 25734
rect 13615 25709 13653 25734
rect 13687 25733 14233 25734
rect 13687 25709 13756 25733
rect 13790 25709 13828 25733
rect 13862 25709 13900 25733
rect 13934 25709 13972 25733
rect 14006 25709 14044 25733
rect 14078 25709 14116 25733
rect 14150 25709 14233 25733
rect 13221 25675 13255 25700
rect 13289 25700 13293 25709
rect 13357 25700 13365 25709
rect 13425 25700 13437 25709
rect 13493 25700 13509 25709
rect 13561 25700 13581 25709
rect 13629 25700 13653 25709
rect 13289 25675 13323 25700
rect 13357 25675 13391 25700
rect 13425 25675 13459 25700
rect 13493 25675 13527 25700
rect 13561 25675 13595 25700
rect 13629 25675 13663 25700
rect 13697 25675 13731 25709
rect 13790 25699 13799 25709
rect 13862 25699 13867 25709
rect 13934 25699 13935 25709
rect 13765 25675 13799 25699
rect 13833 25675 13867 25699
rect 13901 25675 13935 25699
rect 13969 25699 13972 25709
rect 14037 25699 14044 25709
rect 14105 25699 14116 25709
rect 13969 25675 14003 25699
rect 14037 25675 14071 25699
rect 14105 25675 14139 25699
rect 14173 25675 14233 25709
rect 9877 25661 14233 25675
rect 9877 25627 9909 25661
rect 9943 25639 9981 25661
rect 10015 25639 10053 25661
rect 10087 25639 10125 25661
rect 10159 25639 10197 25661
rect 10231 25639 10269 25661
rect 10303 25639 10341 25661
rect 10375 25639 10413 25661
rect 10447 25639 10485 25661
rect 10519 25639 10557 25661
rect 10591 25639 10629 25661
rect 10663 25639 10701 25661
rect 10735 25639 10773 25661
rect 9877 25605 9911 25627
rect 9945 25605 9980 25639
rect 10015 25627 10049 25639
rect 10087 25627 10118 25639
rect 10159 25627 10187 25639
rect 10231 25627 10256 25639
rect 10303 25627 10325 25639
rect 10375 25627 10394 25639
rect 10447 25627 10463 25639
rect 10519 25627 10532 25639
rect 10591 25627 10601 25639
rect 10663 25627 10670 25639
rect 10735 25627 10739 25639
rect 10014 25605 10049 25627
rect 10083 25605 10118 25627
rect 10152 25605 10187 25627
rect 10221 25605 10256 25627
rect 10290 25605 10325 25627
rect 10359 25605 10394 25627
rect 10428 25605 10463 25627
rect 10497 25605 10532 25627
rect 10566 25605 10601 25627
rect 10635 25605 10670 25627
rect 10704 25605 10739 25627
rect 10807 25639 10845 25661
rect 10879 25639 10917 25661
rect 10951 25639 10989 25661
rect 11023 25639 11061 25661
rect 11095 25639 11133 25661
rect 11167 25639 11205 25661
rect 11239 25639 11277 25661
rect 11311 25639 11349 25661
rect 11383 25639 11421 25661
rect 11455 25639 11493 25661
rect 11527 25639 11565 25661
rect 11599 25639 11637 25661
rect 11671 25639 11709 25661
rect 11743 25639 11781 25661
rect 11815 25639 11853 25661
rect 11887 25639 11925 25661
rect 11959 25639 11997 25661
rect 10773 25605 10807 25627
rect 10841 25627 10845 25639
rect 10909 25627 10917 25639
rect 10977 25627 10989 25639
rect 11045 25627 11061 25639
rect 11113 25627 11133 25639
rect 11181 25627 11205 25639
rect 11249 25627 11277 25639
rect 11317 25627 11349 25639
rect 10841 25605 10875 25627
rect 10909 25605 10943 25627
rect 10977 25605 11011 25627
rect 11045 25605 11079 25627
rect 11113 25605 11147 25627
rect 11181 25605 11215 25627
rect 11249 25605 11283 25627
rect 11317 25605 11351 25627
rect 11385 25605 11419 25639
rect 11455 25627 11487 25639
rect 11527 25627 11555 25639
rect 11599 25627 11623 25639
rect 11671 25627 11691 25639
rect 11743 25627 11759 25639
rect 11815 25627 11827 25639
rect 11887 25627 11895 25639
rect 11959 25627 11963 25639
rect 11453 25605 11487 25627
rect 11521 25605 11555 25627
rect 11589 25605 11623 25627
rect 11657 25605 11691 25627
rect 11725 25605 11759 25627
rect 11793 25605 11827 25627
rect 11861 25605 11895 25627
rect 11929 25605 11963 25627
rect 12031 25639 12069 25661
rect 12103 25639 12141 25661
rect 12175 25639 12213 25661
rect 12247 25639 12285 25661
rect 12319 25639 12357 25661
rect 12391 25639 12429 25661
rect 12463 25639 12501 25661
rect 12535 25639 12573 25661
rect 12607 25639 12645 25661
rect 12679 25639 12717 25661
rect 12751 25639 12789 25661
rect 12823 25639 12861 25661
rect 12895 25639 12933 25661
rect 12967 25639 13005 25661
rect 13039 25639 13077 25661
rect 13111 25639 13149 25661
rect 13183 25639 13221 25661
rect 11997 25605 12031 25627
rect 12065 25627 12069 25639
rect 12133 25627 12141 25639
rect 12201 25627 12213 25639
rect 12269 25627 12285 25639
rect 12337 25627 12357 25639
rect 12405 25627 12429 25639
rect 12473 25627 12501 25639
rect 12541 25627 12573 25639
rect 12065 25605 12099 25627
rect 12133 25605 12167 25627
rect 12201 25605 12235 25627
rect 12269 25605 12303 25627
rect 12337 25605 12371 25627
rect 12405 25605 12439 25627
rect 12473 25605 12507 25627
rect 12541 25605 12575 25627
rect 12609 25605 12643 25639
rect 12679 25627 12711 25639
rect 12751 25627 12779 25639
rect 12823 25627 12847 25639
rect 12895 25627 12915 25639
rect 12967 25627 12983 25639
rect 13039 25627 13051 25639
rect 13111 25627 13119 25639
rect 13183 25627 13187 25639
rect 12677 25605 12711 25627
rect 12745 25605 12779 25627
rect 12813 25605 12847 25627
rect 12881 25605 12915 25627
rect 12949 25605 12983 25627
rect 13017 25605 13051 25627
rect 13085 25605 13119 25627
rect 13153 25605 13187 25627
rect 13255 25639 13293 25661
rect 13327 25639 13365 25661
rect 13399 25639 13437 25661
rect 13471 25639 13509 25661
rect 13543 25639 13581 25661
rect 13615 25639 13653 25661
rect 13687 25659 14233 25661
rect 13687 25639 13756 25659
rect 13790 25639 13828 25659
rect 13862 25639 13900 25659
rect 13934 25639 13972 25659
rect 14006 25639 14044 25659
rect 14078 25639 14116 25659
rect 14150 25639 14233 25659
rect 13221 25605 13255 25627
rect 13289 25627 13293 25639
rect 13357 25627 13365 25639
rect 13425 25627 13437 25639
rect 13493 25627 13509 25639
rect 13561 25627 13581 25639
rect 13629 25627 13653 25639
rect 13289 25605 13323 25627
rect 13357 25605 13391 25627
rect 13425 25605 13459 25627
rect 13493 25605 13527 25627
rect 13561 25605 13595 25627
rect 13629 25605 13663 25627
rect 13697 25605 13731 25639
rect 13790 25625 13799 25639
rect 13862 25625 13867 25639
rect 13934 25625 13935 25639
rect 13765 25605 13799 25625
rect 13833 25605 13867 25625
rect 13901 25605 13935 25625
rect 13969 25625 13972 25639
rect 14037 25625 14044 25639
rect 14105 25625 14116 25639
rect 13969 25605 14003 25625
rect 14037 25605 14071 25625
rect 14105 25605 14139 25625
rect 14173 25605 14233 25639
rect 9877 25588 14233 25605
rect 9877 25554 9909 25588
rect 9943 25569 9981 25588
rect 10015 25569 10053 25588
rect 10087 25569 10125 25588
rect 10159 25569 10197 25588
rect 10231 25569 10269 25588
rect 10303 25569 10341 25588
rect 10375 25569 10413 25588
rect 10447 25569 10485 25588
rect 10519 25569 10557 25588
rect 10591 25569 10629 25588
rect 10663 25569 10701 25588
rect 10735 25569 10773 25588
rect 9877 25535 9911 25554
rect 9945 25535 9980 25569
rect 10015 25554 10049 25569
rect 10087 25554 10118 25569
rect 10159 25554 10187 25569
rect 10231 25554 10256 25569
rect 10303 25554 10325 25569
rect 10375 25554 10394 25569
rect 10447 25554 10463 25569
rect 10519 25554 10532 25569
rect 10591 25554 10601 25569
rect 10663 25554 10670 25569
rect 10735 25554 10739 25569
rect 10014 25535 10049 25554
rect 10083 25535 10118 25554
rect 10152 25535 10187 25554
rect 10221 25535 10256 25554
rect 10290 25535 10325 25554
rect 10359 25535 10394 25554
rect 10428 25535 10463 25554
rect 10497 25535 10532 25554
rect 10566 25535 10601 25554
rect 10635 25535 10670 25554
rect 10704 25535 10739 25554
rect 10807 25569 10845 25588
rect 10879 25569 10917 25588
rect 10951 25569 10989 25588
rect 11023 25569 11061 25588
rect 11095 25569 11133 25588
rect 11167 25569 11205 25588
rect 11239 25569 11277 25588
rect 11311 25569 11349 25588
rect 11383 25569 11421 25588
rect 11455 25569 11493 25588
rect 11527 25569 11565 25588
rect 11599 25569 11637 25588
rect 11671 25569 11709 25588
rect 11743 25569 11781 25588
rect 11815 25569 11853 25588
rect 11887 25569 11925 25588
rect 11959 25569 11997 25588
rect 10773 25535 10807 25554
rect 10841 25554 10845 25569
rect 10909 25554 10917 25569
rect 10977 25554 10989 25569
rect 11045 25554 11061 25569
rect 11113 25554 11133 25569
rect 11181 25554 11205 25569
rect 11249 25554 11277 25569
rect 11317 25554 11349 25569
rect 10841 25535 10875 25554
rect 10909 25535 10943 25554
rect 10977 25535 11011 25554
rect 11045 25535 11079 25554
rect 11113 25535 11147 25554
rect 11181 25535 11215 25554
rect 11249 25535 11283 25554
rect 11317 25535 11351 25554
rect 11385 25535 11419 25569
rect 11455 25554 11487 25569
rect 11527 25554 11555 25569
rect 11599 25554 11623 25569
rect 11671 25554 11691 25569
rect 11743 25554 11759 25569
rect 11815 25554 11827 25569
rect 11887 25554 11895 25569
rect 11959 25554 11963 25569
rect 11453 25535 11487 25554
rect 11521 25535 11555 25554
rect 11589 25535 11623 25554
rect 11657 25535 11691 25554
rect 11725 25535 11759 25554
rect 11793 25535 11827 25554
rect 11861 25535 11895 25554
rect 11929 25535 11963 25554
rect 12031 25569 12069 25588
rect 12103 25569 12141 25588
rect 12175 25569 12213 25588
rect 12247 25569 12285 25588
rect 12319 25569 12357 25588
rect 12391 25569 12429 25588
rect 12463 25569 12501 25588
rect 12535 25569 12573 25588
rect 12607 25569 12645 25588
rect 12679 25569 12717 25588
rect 12751 25569 12789 25588
rect 12823 25569 12861 25588
rect 12895 25569 12933 25588
rect 12967 25569 13005 25588
rect 13039 25569 13077 25588
rect 13111 25569 13149 25588
rect 13183 25569 13221 25588
rect 11997 25535 12031 25554
rect 12065 25554 12069 25569
rect 12133 25554 12141 25569
rect 12201 25554 12213 25569
rect 12269 25554 12285 25569
rect 12337 25554 12357 25569
rect 12405 25554 12429 25569
rect 12473 25554 12501 25569
rect 12541 25554 12573 25569
rect 12065 25535 12099 25554
rect 12133 25535 12167 25554
rect 12201 25535 12235 25554
rect 12269 25535 12303 25554
rect 12337 25535 12371 25554
rect 12405 25535 12439 25554
rect 12473 25535 12507 25554
rect 12541 25535 12575 25554
rect 12609 25535 12643 25569
rect 12679 25554 12711 25569
rect 12751 25554 12779 25569
rect 12823 25554 12847 25569
rect 12895 25554 12915 25569
rect 12967 25554 12983 25569
rect 13039 25554 13051 25569
rect 13111 25554 13119 25569
rect 13183 25554 13187 25569
rect 12677 25535 12711 25554
rect 12745 25535 12779 25554
rect 12813 25535 12847 25554
rect 12881 25535 12915 25554
rect 12949 25535 12983 25554
rect 13017 25535 13051 25554
rect 13085 25535 13119 25554
rect 13153 25535 13187 25554
rect 13255 25569 13293 25588
rect 13327 25569 13365 25588
rect 13399 25569 13437 25588
rect 13471 25569 13509 25588
rect 13543 25569 13581 25588
rect 13615 25569 13653 25588
rect 13687 25585 14233 25588
rect 13687 25569 13756 25585
rect 13790 25569 13828 25585
rect 13862 25569 13900 25585
rect 13934 25569 13972 25585
rect 14006 25569 14044 25585
rect 14078 25569 14116 25585
rect 14150 25569 14233 25585
rect 13221 25535 13255 25554
rect 13289 25554 13293 25569
rect 13357 25554 13365 25569
rect 13425 25554 13437 25569
rect 13493 25554 13509 25569
rect 13561 25554 13581 25569
rect 13629 25554 13653 25569
rect 13289 25535 13323 25554
rect 13357 25535 13391 25554
rect 13425 25535 13459 25554
rect 13493 25535 13527 25554
rect 13561 25535 13595 25554
rect 13629 25535 13663 25554
rect 13697 25535 13731 25569
rect 13790 25551 13799 25569
rect 13862 25551 13867 25569
rect 13934 25551 13935 25569
rect 13765 25535 13799 25551
rect 13833 25535 13867 25551
rect 13901 25535 13935 25551
rect 13969 25551 13972 25569
rect 14037 25551 14044 25569
rect 14105 25551 14116 25569
rect 13969 25535 14003 25551
rect 14037 25535 14071 25551
rect 14105 25535 14139 25551
rect 14173 25535 14233 25569
rect 9877 25515 14233 25535
rect 9877 25481 9909 25515
rect 9943 25499 9981 25515
rect 10015 25499 10053 25515
rect 10087 25499 10125 25515
rect 10159 25499 10197 25515
rect 10231 25499 10269 25515
rect 10303 25499 10341 25515
rect 10375 25499 10413 25515
rect 10447 25499 10485 25515
rect 10519 25499 10557 25515
rect 10591 25499 10629 25515
rect 10663 25499 10701 25515
rect 10735 25499 10773 25515
rect 9877 25465 9911 25481
rect 9945 25465 9980 25499
rect 10015 25481 10049 25499
rect 10087 25481 10118 25499
rect 10159 25481 10187 25499
rect 10231 25481 10256 25499
rect 10303 25481 10325 25499
rect 10375 25481 10394 25499
rect 10447 25481 10463 25499
rect 10519 25481 10532 25499
rect 10591 25481 10601 25499
rect 10663 25481 10670 25499
rect 10735 25481 10739 25499
rect 10014 25465 10049 25481
rect 10083 25465 10118 25481
rect 10152 25465 10187 25481
rect 10221 25465 10256 25481
rect 10290 25465 10325 25481
rect 10359 25465 10394 25481
rect 10428 25465 10463 25481
rect 10497 25465 10532 25481
rect 10566 25465 10601 25481
rect 10635 25465 10670 25481
rect 10704 25465 10739 25481
rect 10807 25499 10845 25515
rect 10879 25499 10917 25515
rect 10951 25499 10989 25515
rect 11023 25499 11061 25515
rect 11095 25499 11133 25515
rect 11167 25499 11205 25515
rect 11239 25499 11277 25515
rect 11311 25499 11349 25515
rect 11383 25499 11421 25515
rect 11455 25499 11493 25515
rect 11527 25499 11565 25515
rect 11599 25499 11637 25515
rect 11671 25499 11709 25515
rect 11743 25499 11781 25515
rect 11815 25499 11853 25515
rect 11887 25499 11925 25515
rect 11959 25499 11997 25515
rect 10773 25465 10807 25481
rect 10841 25481 10845 25499
rect 10909 25481 10917 25499
rect 10977 25481 10989 25499
rect 11045 25481 11061 25499
rect 11113 25481 11133 25499
rect 11181 25481 11205 25499
rect 11249 25481 11277 25499
rect 11317 25481 11349 25499
rect 10841 25465 10875 25481
rect 10909 25465 10943 25481
rect 10977 25465 11011 25481
rect 11045 25465 11079 25481
rect 11113 25465 11147 25481
rect 11181 25465 11215 25481
rect 11249 25465 11283 25481
rect 11317 25465 11351 25481
rect 11385 25465 11419 25499
rect 11455 25481 11487 25499
rect 11527 25481 11555 25499
rect 11599 25481 11623 25499
rect 11671 25481 11691 25499
rect 11743 25481 11759 25499
rect 11815 25481 11827 25499
rect 11887 25481 11895 25499
rect 11959 25481 11963 25499
rect 11453 25465 11487 25481
rect 11521 25465 11555 25481
rect 11589 25465 11623 25481
rect 11657 25465 11691 25481
rect 11725 25465 11759 25481
rect 11793 25465 11827 25481
rect 11861 25465 11895 25481
rect 11929 25465 11963 25481
rect 12031 25499 12069 25515
rect 12103 25499 12141 25515
rect 12175 25499 12213 25515
rect 12247 25499 12285 25515
rect 12319 25499 12357 25515
rect 12391 25499 12429 25515
rect 12463 25499 12501 25515
rect 12535 25499 12573 25515
rect 12607 25499 12645 25515
rect 12679 25499 12717 25515
rect 12751 25499 12789 25515
rect 12823 25499 12861 25515
rect 12895 25499 12933 25515
rect 12967 25499 13005 25515
rect 13039 25499 13077 25515
rect 13111 25499 13149 25515
rect 13183 25499 13221 25515
rect 11997 25465 12031 25481
rect 12065 25481 12069 25499
rect 12133 25481 12141 25499
rect 12201 25481 12213 25499
rect 12269 25481 12285 25499
rect 12337 25481 12357 25499
rect 12405 25481 12429 25499
rect 12473 25481 12501 25499
rect 12541 25481 12573 25499
rect 12065 25465 12099 25481
rect 12133 25465 12167 25481
rect 12201 25465 12235 25481
rect 12269 25465 12303 25481
rect 12337 25465 12371 25481
rect 12405 25465 12439 25481
rect 12473 25465 12507 25481
rect 12541 25465 12575 25481
rect 12609 25465 12643 25499
rect 12679 25481 12711 25499
rect 12751 25481 12779 25499
rect 12823 25481 12847 25499
rect 12895 25481 12915 25499
rect 12967 25481 12983 25499
rect 13039 25481 13051 25499
rect 13111 25481 13119 25499
rect 13183 25481 13187 25499
rect 12677 25465 12711 25481
rect 12745 25465 12779 25481
rect 12813 25465 12847 25481
rect 12881 25465 12915 25481
rect 12949 25465 12983 25481
rect 13017 25465 13051 25481
rect 13085 25465 13119 25481
rect 13153 25465 13187 25481
rect 13255 25499 13293 25515
rect 13327 25499 13365 25515
rect 13399 25499 13437 25515
rect 13471 25499 13509 25515
rect 13543 25499 13581 25515
rect 13615 25499 13653 25515
rect 13687 25511 14233 25515
rect 13687 25499 13756 25511
rect 13790 25499 13828 25511
rect 13862 25499 13900 25511
rect 13934 25499 13972 25511
rect 14006 25499 14044 25511
rect 14078 25499 14116 25511
rect 14150 25499 14233 25511
rect 13221 25465 13255 25481
rect 13289 25481 13293 25499
rect 13357 25481 13365 25499
rect 13425 25481 13437 25499
rect 13493 25481 13509 25499
rect 13561 25481 13581 25499
rect 13629 25481 13653 25499
rect 13289 25465 13323 25481
rect 13357 25465 13391 25481
rect 13425 25465 13459 25481
rect 13493 25465 13527 25481
rect 13561 25465 13595 25481
rect 13629 25465 13663 25481
rect 13697 25465 13731 25499
rect 13790 25477 13799 25499
rect 13862 25477 13867 25499
rect 13934 25477 13935 25499
rect 13765 25465 13799 25477
rect 13833 25465 13867 25477
rect 13901 25465 13935 25477
rect 13969 25477 13972 25499
rect 14037 25477 14044 25499
rect 14105 25477 14116 25499
rect 13969 25465 14003 25477
rect 14037 25465 14071 25477
rect 14105 25465 14139 25477
rect 14173 25465 14233 25499
rect 9877 25442 14233 25465
rect 9877 25408 9909 25442
rect 9943 25429 9981 25442
rect 10015 25429 10053 25442
rect 10087 25429 10125 25442
rect 10159 25429 10197 25442
rect 10231 25429 10269 25442
rect 10303 25429 10341 25442
rect 10375 25429 10413 25442
rect 10447 25429 10485 25442
rect 10519 25429 10557 25442
rect 10591 25429 10629 25442
rect 10663 25429 10701 25442
rect 10735 25429 10773 25442
rect 9877 25395 9911 25408
rect 9945 25395 9980 25429
rect 10015 25408 10049 25429
rect 10087 25408 10118 25429
rect 10159 25408 10187 25429
rect 10231 25408 10256 25429
rect 10303 25408 10325 25429
rect 10375 25408 10394 25429
rect 10447 25408 10463 25429
rect 10519 25408 10532 25429
rect 10591 25408 10601 25429
rect 10663 25408 10670 25429
rect 10735 25408 10739 25429
rect 10014 25395 10049 25408
rect 10083 25395 10118 25408
rect 10152 25395 10187 25408
rect 10221 25395 10256 25408
rect 10290 25395 10325 25408
rect 10359 25395 10394 25408
rect 10428 25395 10463 25408
rect 10497 25395 10532 25408
rect 10566 25395 10601 25408
rect 10635 25395 10670 25408
rect 10704 25395 10739 25408
rect 10807 25429 10845 25442
rect 10879 25429 10917 25442
rect 10951 25429 10989 25442
rect 11023 25429 11061 25442
rect 11095 25429 11133 25442
rect 11167 25429 11205 25442
rect 11239 25429 11277 25442
rect 11311 25429 11349 25442
rect 11383 25429 11421 25442
rect 11455 25429 11493 25442
rect 11527 25429 11565 25442
rect 11599 25429 11637 25442
rect 11671 25429 11709 25442
rect 11743 25429 11781 25442
rect 11815 25429 11853 25442
rect 11887 25429 11925 25442
rect 11959 25429 11997 25442
rect 10773 25395 10807 25408
rect 10841 25408 10845 25429
rect 10909 25408 10917 25429
rect 10977 25408 10989 25429
rect 11045 25408 11061 25429
rect 11113 25408 11133 25429
rect 11181 25408 11205 25429
rect 11249 25408 11277 25429
rect 11317 25408 11349 25429
rect 10841 25395 10875 25408
rect 10909 25395 10943 25408
rect 10977 25395 11011 25408
rect 11045 25395 11079 25408
rect 11113 25395 11147 25408
rect 11181 25395 11215 25408
rect 11249 25395 11283 25408
rect 11317 25395 11351 25408
rect 11385 25395 11419 25429
rect 11455 25408 11487 25429
rect 11527 25408 11555 25429
rect 11599 25408 11623 25429
rect 11671 25408 11691 25429
rect 11743 25408 11759 25429
rect 11815 25408 11827 25429
rect 11887 25408 11895 25429
rect 11959 25408 11963 25429
rect 11453 25395 11487 25408
rect 11521 25395 11555 25408
rect 11589 25395 11623 25408
rect 11657 25395 11691 25408
rect 11725 25395 11759 25408
rect 11793 25395 11827 25408
rect 11861 25395 11895 25408
rect 11929 25395 11963 25408
rect 12031 25429 12069 25442
rect 12103 25429 12141 25442
rect 12175 25429 12213 25442
rect 12247 25429 12285 25442
rect 12319 25429 12357 25442
rect 12391 25429 12429 25442
rect 12463 25429 12501 25442
rect 12535 25429 12573 25442
rect 12607 25429 12645 25442
rect 12679 25429 12717 25442
rect 12751 25429 12789 25442
rect 12823 25429 12861 25442
rect 12895 25429 12933 25442
rect 12967 25429 13005 25442
rect 13039 25429 13077 25442
rect 13111 25429 13149 25442
rect 13183 25429 13221 25442
rect 11997 25395 12031 25408
rect 12065 25408 12069 25429
rect 12133 25408 12141 25429
rect 12201 25408 12213 25429
rect 12269 25408 12285 25429
rect 12337 25408 12357 25429
rect 12405 25408 12429 25429
rect 12473 25408 12501 25429
rect 12541 25408 12573 25429
rect 12065 25395 12099 25408
rect 12133 25395 12167 25408
rect 12201 25395 12235 25408
rect 12269 25395 12303 25408
rect 12337 25395 12371 25408
rect 12405 25395 12439 25408
rect 12473 25395 12507 25408
rect 12541 25395 12575 25408
rect 12609 25395 12643 25429
rect 12679 25408 12711 25429
rect 12751 25408 12779 25429
rect 12823 25408 12847 25429
rect 12895 25408 12915 25429
rect 12967 25408 12983 25429
rect 13039 25408 13051 25429
rect 13111 25408 13119 25429
rect 13183 25408 13187 25429
rect 12677 25395 12711 25408
rect 12745 25395 12779 25408
rect 12813 25395 12847 25408
rect 12881 25395 12915 25408
rect 12949 25395 12983 25408
rect 13017 25395 13051 25408
rect 13085 25395 13119 25408
rect 13153 25395 13187 25408
rect 13255 25429 13293 25442
rect 13327 25429 13365 25442
rect 13399 25429 13437 25442
rect 13471 25429 13509 25442
rect 13543 25429 13581 25442
rect 13615 25429 13653 25442
rect 13687 25437 14233 25442
rect 13687 25429 13756 25437
rect 13790 25429 13828 25437
rect 13862 25429 13900 25437
rect 13934 25429 13972 25437
rect 14006 25429 14044 25437
rect 14078 25429 14116 25437
rect 14150 25429 14233 25437
rect 13221 25395 13255 25408
rect 13289 25408 13293 25429
rect 13357 25408 13365 25429
rect 13425 25408 13437 25429
rect 13493 25408 13509 25429
rect 13561 25408 13581 25429
rect 13629 25408 13653 25429
rect 13289 25395 13323 25408
rect 13357 25395 13391 25408
rect 13425 25395 13459 25408
rect 13493 25395 13527 25408
rect 13561 25395 13595 25408
rect 13629 25395 13663 25408
rect 13697 25395 13731 25429
rect 13790 25403 13799 25429
rect 13862 25403 13867 25429
rect 13934 25403 13935 25429
rect 13765 25395 13799 25403
rect 13833 25395 13867 25403
rect 13901 25395 13935 25403
rect 13969 25403 13972 25429
rect 14037 25403 14044 25429
rect 14105 25403 14116 25429
rect 13969 25395 14003 25403
rect 14037 25395 14071 25403
rect 14105 25395 14139 25403
rect 14173 25395 14233 25429
rect 9877 25369 14233 25395
rect 9877 25335 9909 25369
rect 9943 25359 9981 25369
rect 10015 25359 10053 25369
rect 10087 25359 10125 25369
rect 10159 25359 10197 25369
rect 10231 25359 10269 25369
rect 10303 25359 10341 25369
rect 10375 25359 10413 25369
rect 10447 25359 10485 25369
rect 10519 25359 10557 25369
rect 10591 25359 10629 25369
rect 10663 25359 10701 25369
rect 10735 25359 10773 25369
rect 9877 25325 9911 25335
rect 9945 25325 9980 25359
rect 10015 25335 10049 25359
rect 10087 25335 10118 25359
rect 10159 25335 10187 25359
rect 10231 25335 10256 25359
rect 10303 25335 10325 25359
rect 10375 25335 10394 25359
rect 10447 25335 10463 25359
rect 10519 25335 10532 25359
rect 10591 25335 10601 25359
rect 10663 25335 10670 25359
rect 10735 25335 10739 25359
rect 10014 25325 10049 25335
rect 10083 25325 10118 25335
rect 10152 25325 10187 25335
rect 10221 25325 10256 25335
rect 10290 25325 10325 25335
rect 10359 25325 10394 25335
rect 10428 25325 10463 25335
rect 10497 25325 10532 25335
rect 10566 25325 10601 25335
rect 10635 25325 10670 25335
rect 10704 25325 10739 25335
rect 10807 25359 10845 25369
rect 10879 25359 10917 25369
rect 10951 25359 10989 25369
rect 11023 25359 11061 25369
rect 11095 25359 11133 25369
rect 11167 25359 11205 25369
rect 11239 25359 11277 25369
rect 11311 25359 11349 25369
rect 11383 25359 11421 25369
rect 11455 25359 11493 25369
rect 11527 25359 11565 25369
rect 11599 25359 11637 25369
rect 11671 25359 11709 25369
rect 11743 25359 11781 25369
rect 11815 25359 11853 25369
rect 11887 25359 11925 25369
rect 11959 25359 11997 25369
rect 10773 25325 10807 25335
rect 10841 25335 10845 25359
rect 10909 25335 10917 25359
rect 10977 25335 10989 25359
rect 11045 25335 11061 25359
rect 11113 25335 11133 25359
rect 11181 25335 11205 25359
rect 11249 25335 11277 25359
rect 11317 25335 11349 25359
rect 10841 25325 10875 25335
rect 10909 25325 10943 25335
rect 10977 25325 11011 25335
rect 11045 25325 11079 25335
rect 11113 25325 11147 25335
rect 11181 25325 11215 25335
rect 11249 25325 11283 25335
rect 11317 25325 11351 25335
rect 11385 25325 11419 25359
rect 11455 25335 11487 25359
rect 11527 25335 11555 25359
rect 11599 25335 11623 25359
rect 11671 25335 11691 25359
rect 11743 25335 11759 25359
rect 11815 25335 11827 25359
rect 11887 25335 11895 25359
rect 11959 25335 11963 25359
rect 11453 25325 11487 25335
rect 11521 25325 11555 25335
rect 11589 25325 11623 25335
rect 11657 25325 11691 25335
rect 11725 25325 11759 25335
rect 11793 25325 11827 25335
rect 11861 25325 11895 25335
rect 11929 25325 11963 25335
rect 12031 25359 12069 25369
rect 12103 25359 12141 25369
rect 12175 25359 12213 25369
rect 12247 25359 12285 25369
rect 12319 25359 12357 25369
rect 12391 25359 12429 25369
rect 12463 25359 12501 25369
rect 12535 25359 12573 25369
rect 12607 25359 12645 25369
rect 12679 25359 12717 25369
rect 12751 25359 12789 25369
rect 12823 25359 12861 25369
rect 12895 25359 12933 25369
rect 12967 25359 13005 25369
rect 13039 25359 13077 25369
rect 13111 25359 13149 25369
rect 13183 25359 13221 25369
rect 11997 25325 12031 25335
rect 12065 25335 12069 25359
rect 12133 25335 12141 25359
rect 12201 25335 12213 25359
rect 12269 25335 12285 25359
rect 12337 25335 12357 25359
rect 12405 25335 12429 25359
rect 12473 25335 12501 25359
rect 12541 25335 12573 25359
rect 12065 25325 12099 25335
rect 12133 25325 12167 25335
rect 12201 25325 12235 25335
rect 12269 25325 12303 25335
rect 12337 25325 12371 25335
rect 12405 25325 12439 25335
rect 12473 25325 12507 25335
rect 12541 25325 12575 25335
rect 12609 25325 12643 25359
rect 12679 25335 12711 25359
rect 12751 25335 12779 25359
rect 12823 25335 12847 25359
rect 12895 25335 12915 25359
rect 12967 25335 12983 25359
rect 13039 25335 13051 25359
rect 13111 25335 13119 25359
rect 13183 25335 13187 25359
rect 12677 25325 12711 25335
rect 12745 25325 12779 25335
rect 12813 25325 12847 25335
rect 12881 25325 12915 25335
rect 12949 25325 12983 25335
rect 13017 25325 13051 25335
rect 13085 25325 13119 25335
rect 13153 25325 13187 25335
rect 13255 25359 13293 25369
rect 13327 25359 13365 25369
rect 13399 25359 13437 25369
rect 13471 25359 13509 25369
rect 13543 25359 13581 25369
rect 13615 25359 13653 25369
rect 13687 25363 14233 25369
rect 13687 25359 13756 25363
rect 13790 25359 13828 25363
rect 13862 25359 13900 25363
rect 13934 25359 13972 25363
rect 14006 25359 14044 25363
rect 14078 25359 14116 25363
rect 14150 25359 14233 25363
rect 13221 25325 13255 25335
rect 13289 25335 13293 25359
rect 13357 25335 13365 25359
rect 13425 25335 13437 25359
rect 13493 25335 13509 25359
rect 13561 25335 13581 25359
rect 13629 25335 13653 25359
rect 13289 25325 13323 25335
rect 13357 25325 13391 25335
rect 13425 25325 13459 25335
rect 13493 25325 13527 25335
rect 13561 25325 13595 25335
rect 13629 25325 13663 25335
rect 13697 25325 13731 25359
rect 13790 25329 13799 25359
rect 13862 25329 13867 25359
rect 13934 25329 13935 25359
rect 13765 25325 13799 25329
rect 13833 25325 13867 25329
rect 13901 25325 13935 25329
rect 13969 25329 13972 25359
rect 14037 25329 14044 25359
rect 14105 25329 14116 25359
rect 13969 25325 14003 25329
rect 14037 25325 14071 25329
rect 14105 25325 14139 25329
rect 14173 25325 14233 25359
rect 9877 25296 14233 25325
rect 9877 25262 9909 25296
rect 9943 25289 9981 25296
rect 10015 25289 10053 25296
rect 10087 25289 10125 25296
rect 10159 25289 10197 25296
rect 10231 25289 10269 25296
rect 10303 25289 10341 25296
rect 10375 25289 10413 25296
rect 10447 25289 10485 25296
rect 10519 25289 10557 25296
rect 10591 25289 10629 25296
rect 10663 25289 10701 25296
rect 10735 25289 10773 25296
rect 9877 25255 9911 25262
rect 9945 25255 9980 25289
rect 10015 25262 10049 25289
rect 10087 25262 10118 25289
rect 10159 25262 10187 25289
rect 10231 25262 10256 25289
rect 10303 25262 10325 25289
rect 10375 25262 10394 25289
rect 10447 25262 10463 25289
rect 10519 25262 10532 25289
rect 10591 25262 10601 25289
rect 10663 25262 10670 25289
rect 10735 25262 10739 25289
rect 10014 25255 10049 25262
rect 10083 25255 10118 25262
rect 10152 25255 10187 25262
rect 10221 25255 10256 25262
rect 10290 25255 10325 25262
rect 10359 25255 10394 25262
rect 10428 25255 10463 25262
rect 10497 25255 10532 25262
rect 10566 25255 10601 25262
rect 10635 25255 10670 25262
rect 10704 25255 10739 25262
rect 10807 25289 10845 25296
rect 10879 25289 10917 25296
rect 10951 25289 10989 25296
rect 11023 25289 11061 25296
rect 11095 25289 11133 25296
rect 11167 25289 11205 25296
rect 11239 25289 11277 25296
rect 11311 25289 11349 25296
rect 11383 25289 11421 25296
rect 11455 25289 11493 25296
rect 11527 25289 11565 25296
rect 11599 25289 11637 25296
rect 11671 25289 11709 25296
rect 11743 25289 11781 25296
rect 11815 25289 11853 25296
rect 11887 25289 11925 25296
rect 11959 25289 11997 25296
rect 10773 25255 10807 25262
rect 10841 25262 10845 25289
rect 10909 25262 10917 25289
rect 10977 25262 10989 25289
rect 11045 25262 11061 25289
rect 11113 25262 11133 25289
rect 11181 25262 11205 25289
rect 11249 25262 11277 25289
rect 11317 25262 11349 25289
rect 10841 25255 10875 25262
rect 10909 25255 10943 25262
rect 10977 25255 11011 25262
rect 11045 25255 11079 25262
rect 11113 25255 11147 25262
rect 11181 25255 11215 25262
rect 11249 25255 11283 25262
rect 11317 25255 11351 25262
rect 11385 25255 11419 25289
rect 11455 25262 11487 25289
rect 11527 25262 11555 25289
rect 11599 25262 11623 25289
rect 11671 25262 11691 25289
rect 11743 25262 11759 25289
rect 11815 25262 11827 25289
rect 11887 25262 11895 25289
rect 11959 25262 11963 25289
rect 11453 25255 11487 25262
rect 11521 25255 11555 25262
rect 11589 25255 11623 25262
rect 11657 25255 11691 25262
rect 11725 25255 11759 25262
rect 11793 25255 11827 25262
rect 11861 25255 11895 25262
rect 11929 25255 11963 25262
rect 12031 25289 12069 25296
rect 12103 25289 12141 25296
rect 12175 25289 12213 25296
rect 12247 25289 12285 25296
rect 12319 25289 12357 25296
rect 12391 25289 12429 25296
rect 12463 25289 12501 25296
rect 12535 25289 12573 25296
rect 12607 25289 12645 25296
rect 12679 25289 12717 25296
rect 12751 25289 12789 25296
rect 12823 25289 12861 25296
rect 12895 25289 12933 25296
rect 12967 25289 13005 25296
rect 13039 25289 13077 25296
rect 13111 25289 13149 25296
rect 13183 25289 13221 25296
rect 11997 25255 12031 25262
rect 12065 25262 12069 25289
rect 12133 25262 12141 25289
rect 12201 25262 12213 25289
rect 12269 25262 12285 25289
rect 12337 25262 12357 25289
rect 12405 25262 12429 25289
rect 12473 25262 12501 25289
rect 12541 25262 12573 25289
rect 12065 25255 12099 25262
rect 12133 25255 12167 25262
rect 12201 25255 12235 25262
rect 12269 25255 12303 25262
rect 12337 25255 12371 25262
rect 12405 25255 12439 25262
rect 12473 25255 12507 25262
rect 12541 25255 12575 25262
rect 12609 25255 12643 25289
rect 12679 25262 12711 25289
rect 12751 25262 12779 25289
rect 12823 25262 12847 25289
rect 12895 25262 12915 25289
rect 12967 25262 12983 25289
rect 13039 25262 13051 25289
rect 13111 25262 13119 25289
rect 13183 25262 13187 25289
rect 12677 25255 12711 25262
rect 12745 25255 12779 25262
rect 12813 25255 12847 25262
rect 12881 25255 12915 25262
rect 12949 25255 12983 25262
rect 13017 25255 13051 25262
rect 13085 25255 13119 25262
rect 13153 25255 13187 25262
rect 13255 25289 13293 25296
rect 13327 25289 13365 25296
rect 13399 25289 13437 25296
rect 13471 25289 13509 25296
rect 13543 25289 13581 25296
rect 13615 25289 13653 25296
rect 13687 25289 14233 25296
rect 13221 25255 13255 25262
rect 13289 25262 13293 25289
rect 13357 25262 13365 25289
rect 13425 25262 13437 25289
rect 13493 25262 13509 25289
rect 13561 25262 13581 25289
rect 13629 25262 13653 25289
rect 13289 25255 13323 25262
rect 13357 25255 13391 25262
rect 13425 25255 13459 25262
rect 13493 25255 13527 25262
rect 13561 25255 13595 25262
rect 13629 25255 13663 25262
rect 13697 25255 13731 25289
rect 13790 25255 13799 25289
rect 13862 25255 13867 25289
rect 13934 25255 13935 25289
rect 13969 25255 13972 25289
rect 14037 25255 14044 25289
rect 14105 25255 14116 25289
rect 14173 25255 14233 25289
rect 9877 25223 14233 25255
rect 9877 25189 9909 25223
rect 9943 25219 9981 25223
rect 10015 25219 10053 25223
rect 10087 25219 10125 25223
rect 10159 25219 10197 25223
rect 10231 25219 10269 25223
rect 10303 25219 10341 25223
rect 10375 25219 10413 25223
rect 10447 25219 10485 25223
rect 10519 25219 10557 25223
rect 10591 25219 10629 25223
rect 10663 25219 10701 25223
rect 10735 25219 10773 25223
rect 9877 25185 9911 25189
rect 9945 25185 9980 25219
rect 10015 25189 10049 25219
rect 10087 25189 10118 25219
rect 10159 25189 10187 25219
rect 10231 25189 10256 25219
rect 10303 25189 10325 25219
rect 10375 25189 10394 25219
rect 10447 25189 10463 25219
rect 10519 25189 10532 25219
rect 10591 25189 10601 25219
rect 10663 25189 10670 25219
rect 10735 25189 10739 25219
rect 10014 25185 10049 25189
rect 10083 25185 10118 25189
rect 10152 25185 10187 25189
rect 10221 25185 10256 25189
rect 10290 25185 10325 25189
rect 10359 25185 10394 25189
rect 10428 25185 10463 25189
rect 10497 25185 10532 25189
rect 10566 25185 10601 25189
rect 10635 25185 10670 25189
rect 10704 25185 10739 25189
rect 10807 25219 10845 25223
rect 10879 25219 10917 25223
rect 10951 25219 10989 25223
rect 11023 25219 11061 25223
rect 11095 25219 11133 25223
rect 11167 25219 11205 25223
rect 11239 25219 11277 25223
rect 11311 25219 11349 25223
rect 11383 25219 11421 25223
rect 11455 25219 11493 25223
rect 11527 25219 11565 25223
rect 11599 25219 11637 25223
rect 11671 25219 11709 25223
rect 11743 25219 11781 25223
rect 11815 25219 11853 25223
rect 11887 25219 11925 25223
rect 11959 25219 11997 25223
rect 10773 25185 10807 25189
rect 10841 25189 10845 25219
rect 10909 25189 10917 25219
rect 10977 25189 10989 25219
rect 11045 25189 11061 25219
rect 11113 25189 11133 25219
rect 11181 25189 11205 25219
rect 11249 25189 11277 25219
rect 11317 25189 11349 25219
rect 10841 25185 10875 25189
rect 10909 25185 10943 25189
rect 10977 25185 11011 25189
rect 11045 25185 11079 25189
rect 11113 25185 11147 25189
rect 11181 25185 11215 25189
rect 11249 25185 11283 25189
rect 11317 25185 11351 25189
rect 11385 25185 11419 25219
rect 11455 25189 11487 25219
rect 11527 25189 11555 25219
rect 11599 25189 11623 25219
rect 11671 25189 11691 25219
rect 11743 25189 11759 25219
rect 11815 25189 11827 25219
rect 11887 25189 11895 25219
rect 11959 25189 11963 25219
rect 11453 25185 11487 25189
rect 11521 25185 11555 25189
rect 11589 25185 11623 25189
rect 11657 25185 11691 25189
rect 11725 25185 11759 25189
rect 11793 25185 11827 25189
rect 11861 25185 11895 25189
rect 11929 25185 11963 25189
rect 12031 25219 12069 25223
rect 12103 25219 12141 25223
rect 12175 25219 12213 25223
rect 12247 25219 12285 25223
rect 12319 25219 12357 25223
rect 12391 25219 12429 25223
rect 12463 25219 12501 25223
rect 12535 25219 12573 25223
rect 12607 25219 12645 25223
rect 12679 25219 12717 25223
rect 12751 25219 12789 25223
rect 12823 25219 12861 25223
rect 12895 25219 12933 25223
rect 12967 25219 13005 25223
rect 13039 25219 13077 25223
rect 13111 25219 13149 25223
rect 13183 25219 13221 25223
rect 11997 25185 12031 25189
rect 12065 25189 12069 25219
rect 12133 25189 12141 25219
rect 12201 25189 12213 25219
rect 12269 25189 12285 25219
rect 12337 25189 12357 25219
rect 12405 25189 12429 25219
rect 12473 25189 12501 25219
rect 12541 25189 12573 25219
rect 12065 25185 12099 25189
rect 12133 25185 12167 25189
rect 12201 25185 12235 25189
rect 12269 25185 12303 25189
rect 12337 25185 12371 25189
rect 12405 25185 12439 25189
rect 12473 25185 12507 25189
rect 12541 25185 12575 25189
rect 12609 25185 12643 25219
rect 12679 25189 12711 25219
rect 12751 25189 12779 25219
rect 12823 25189 12847 25219
rect 12895 25189 12915 25219
rect 12967 25189 12983 25219
rect 13039 25189 13051 25219
rect 13111 25189 13119 25219
rect 13183 25189 13187 25219
rect 12677 25185 12711 25189
rect 12745 25185 12779 25189
rect 12813 25185 12847 25189
rect 12881 25185 12915 25189
rect 12949 25185 12983 25189
rect 13017 25185 13051 25189
rect 13085 25185 13119 25189
rect 13153 25185 13187 25189
rect 13255 25219 13293 25223
rect 13327 25219 13365 25223
rect 13399 25219 13437 25223
rect 13471 25219 13509 25223
rect 13543 25219 13581 25223
rect 13615 25219 13653 25223
rect 13687 25219 14233 25223
rect 13221 25185 13255 25189
rect 13289 25189 13293 25219
rect 13357 25189 13365 25219
rect 13425 25189 13437 25219
rect 13493 25189 13509 25219
rect 13561 25189 13581 25219
rect 13629 25189 13653 25219
rect 13289 25185 13323 25189
rect 13357 25185 13391 25189
rect 13425 25185 13459 25189
rect 13493 25185 13527 25189
rect 13561 25185 13595 25189
rect 13629 25185 13663 25189
rect 13697 25185 13731 25219
rect 13765 25215 13799 25219
rect 13833 25215 13867 25219
rect 13901 25215 13935 25219
rect 13790 25185 13799 25215
rect 13862 25185 13867 25215
rect 13934 25185 13935 25215
rect 13969 25215 14003 25219
rect 14037 25215 14071 25219
rect 14105 25215 14139 25219
rect 13969 25185 13972 25215
rect 14037 25185 14044 25215
rect 14105 25185 14116 25215
rect 14173 25185 14233 25219
rect 9877 25181 13756 25185
rect 13790 25181 13828 25185
rect 13862 25181 13900 25185
rect 13934 25181 13972 25185
rect 14006 25181 14044 25185
rect 14078 25181 14116 25185
rect 14150 25181 14233 25185
rect 9877 25150 14233 25181
rect 9877 25116 9909 25150
rect 9943 25149 9981 25150
rect 10015 25149 10053 25150
rect 10087 25149 10125 25150
rect 10159 25149 10197 25150
rect 10231 25149 10269 25150
rect 10303 25149 10341 25150
rect 10375 25149 10413 25150
rect 10447 25149 10485 25150
rect 10519 25149 10557 25150
rect 10591 25149 10629 25150
rect 10663 25149 10701 25150
rect 10735 25149 10773 25150
rect 9877 25115 9911 25116
rect 9945 25115 9980 25149
rect 10015 25116 10049 25149
rect 10087 25116 10118 25149
rect 10159 25116 10187 25149
rect 10231 25116 10256 25149
rect 10303 25116 10325 25149
rect 10375 25116 10394 25149
rect 10447 25116 10463 25149
rect 10519 25116 10532 25149
rect 10591 25116 10601 25149
rect 10663 25116 10670 25149
rect 10735 25116 10739 25149
rect 10014 25115 10049 25116
rect 10083 25115 10118 25116
rect 10152 25115 10187 25116
rect 10221 25115 10256 25116
rect 10290 25115 10325 25116
rect 10359 25115 10394 25116
rect 10428 25115 10463 25116
rect 10497 25115 10532 25116
rect 10566 25115 10601 25116
rect 10635 25115 10670 25116
rect 10704 25115 10739 25116
rect 10807 25149 10845 25150
rect 10879 25149 10917 25150
rect 10951 25149 10989 25150
rect 11023 25149 11061 25150
rect 11095 25149 11133 25150
rect 11167 25149 11205 25150
rect 11239 25149 11277 25150
rect 11311 25149 11349 25150
rect 11383 25149 11421 25150
rect 11455 25149 11493 25150
rect 11527 25149 11565 25150
rect 11599 25149 11637 25150
rect 11671 25149 11709 25150
rect 11743 25149 11781 25150
rect 11815 25149 11853 25150
rect 11887 25149 11925 25150
rect 11959 25149 11997 25150
rect 10773 25115 10807 25116
rect 10841 25116 10845 25149
rect 10909 25116 10917 25149
rect 10977 25116 10989 25149
rect 11045 25116 11061 25149
rect 11113 25116 11133 25149
rect 11181 25116 11205 25149
rect 11249 25116 11277 25149
rect 11317 25116 11349 25149
rect 10841 25115 10875 25116
rect 10909 25115 10943 25116
rect 10977 25115 11011 25116
rect 11045 25115 11079 25116
rect 11113 25115 11147 25116
rect 11181 25115 11215 25116
rect 11249 25115 11283 25116
rect 11317 25115 11351 25116
rect 11385 25115 11419 25149
rect 11455 25116 11487 25149
rect 11527 25116 11555 25149
rect 11599 25116 11623 25149
rect 11671 25116 11691 25149
rect 11743 25116 11759 25149
rect 11815 25116 11827 25149
rect 11887 25116 11895 25149
rect 11959 25116 11963 25149
rect 11453 25115 11487 25116
rect 11521 25115 11555 25116
rect 11589 25115 11623 25116
rect 11657 25115 11691 25116
rect 11725 25115 11759 25116
rect 11793 25115 11827 25116
rect 11861 25115 11895 25116
rect 11929 25115 11963 25116
rect 12031 25149 12069 25150
rect 12103 25149 12141 25150
rect 12175 25149 12213 25150
rect 12247 25149 12285 25150
rect 12319 25149 12357 25150
rect 12391 25149 12429 25150
rect 12463 25149 12501 25150
rect 12535 25149 12573 25150
rect 12607 25149 12645 25150
rect 12679 25149 12717 25150
rect 12751 25149 12789 25150
rect 12823 25149 12861 25150
rect 12895 25149 12933 25150
rect 12967 25149 13005 25150
rect 13039 25149 13077 25150
rect 13111 25149 13149 25150
rect 13183 25149 13221 25150
rect 11997 25115 12031 25116
rect 12065 25116 12069 25149
rect 12133 25116 12141 25149
rect 12201 25116 12213 25149
rect 12269 25116 12285 25149
rect 12337 25116 12357 25149
rect 12405 25116 12429 25149
rect 12473 25116 12501 25149
rect 12541 25116 12573 25149
rect 12065 25115 12099 25116
rect 12133 25115 12167 25116
rect 12201 25115 12235 25116
rect 12269 25115 12303 25116
rect 12337 25115 12371 25116
rect 12405 25115 12439 25116
rect 12473 25115 12507 25116
rect 12541 25115 12575 25116
rect 12609 25115 12643 25149
rect 12679 25116 12711 25149
rect 12751 25116 12779 25149
rect 12823 25116 12847 25149
rect 12895 25116 12915 25149
rect 12967 25116 12983 25149
rect 13039 25116 13051 25149
rect 13111 25116 13119 25149
rect 13183 25116 13187 25149
rect 12677 25115 12711 25116
rect 12745 25115 12779 25116
rect 12813 25115 12847 25116
rect 12881 25115 12915 25116
rect 12949 25115 12983 25116
rect 13017 25115 13051 25116
rect 13085 25115 13119 25116
rect 13153 25115 13187 25116
rect 13255 25149 13293 25150
rect 13327 25149 13365 25150
rect 13399 25149 13437 25150
rect 13471 25149 13509 25150
rect 13543 25149 13581 25150
rect 13615 25149 13653 25150
rect 13687 25149 14233 25150
rect 13221 25115 13255 25116
rect 13289 25116 13293 25149
rect 13357 25116 13365 25149
rect 13425 25116 13437 25149
rect 13493 25116 13509 25149
rect 13561 25116 13581 25149
rect 13629 25116 13653 25149
rect 13289 25115 13323 25116
rect 13357 25115 13391 25116
rect 13425 25115 13459 25116
rect 13493 25115 13527 25116
rect 13561 25115 13595 25116
rect 13629 25115 13663 25116
rect 13697 25115 13731 25149
rect 13765 25141 13799 25149
rect 13833 25141 13867 25149
rect 13901 25141 13935 25149
rect 13790 25115 13799 25141
rect 13862 25115 13867 25141
rect 13934 25115 13935 25141
rect 13969 25141 14003 25149
rect 14037 25141 14071 25149
rect 14105 25141 14139 25149
rect 13969 25115 13972 25141
rect 14037 25115 14044 25141
rect 14105 25115 14116 25141
rect 14173 25115 14233 25149
rect 9877 25107 13756 25115
rect 13790 25107 13828 25115
rect 13862 25107 13900 25115
rect 13934 25107 13972 25115
rect 14006 25107 14044 25115
rect 14078 25107 14116 25115
rect 14150 25107 14233 25115
rect 9877 25079 14233 25107
rect 9877 25045 9911 25079
rect 9945 25045 9980 25079
rect 10014 25045 10049 25079
rect 10083 25045 10118 25079
rect 10152 25045 10187 25079
rect 10221 25045 10256 25079
rect 10290 25045 10325 25079
rect 10359 25045 10394 25079
rect 10428 25045 10463 25079
rect 10497 25045 10532 25079
rect 10566 25045 10601 25079
rect 10635 25045 10670 25079
rect 10704 25045 10739 25079
rect 10773 25045 10807 25079
rect 10841 25045 10875 25079
rect 10909 25045 10943 25079
rect 10977 25045 11011 25079
rect 11045 25045 11079 25079
rect 11113 25045 11147 25079
rect 11181 25045 11215 25079
rect 11249 25045 11283 25079
rect 11317 25045 11351 25079
rect 11385 25045 11419 25079
rect 11453 25045 11487 25079
rect 11521 25045 11555 25079
rect 11589 25045 11623 25079
rect 11657 25045 11691 25079
rect 11725 25045 11759 25079
rect 11793 25045 11827 25079
rect 11861 25045 11895 25079
rect 11929 25045 11963 25079
rect 11997 25045 12031 25079
rect 12065 25045 12099 25079
rect 12133 25045 12167 25079
rect 12201 25045 12235 25079
rect 12269 25045 12303 25079
rect 12337 25045 12371 25079
rect 12405 25045 12439 25079
rect 12473 25045 12507 25079
rect 12541 25045 12575 25079
rect 12609 25045 12643 25079
rect 12677 25045 12711 25079
rect 12745 25045 12779 25079
rect 12813 25045 12847 25079
rect 12881 25045 12915 25079
rect 12949 25045 12983 25079
rect 13017 25045 13051 25079
rect 13085 25045 13119 25079
rect 13153 25045 13187 25079
rect 13221 25045 13255 25079
rect 13289 25045 13323 25079
rect 13357 25045 13391 25079
rect 13425 25045 13459 25079
rect 13493 25045 13527 25079
rect 13561 25045 13595 25079
rect 13629 25045 13663 25079
rect 13697 25045 13731 25079
rect 13765 25067 13799 25079
rect 13833 25067 13867 25079
rect 13901 25067 13935 25079
rect 13790 25045 13799 25067
rect 13862 25045 13867 25067
rect 13934 25045 13935 25067
rect 13969 25067 14003 25079
rect 14037 25067 14071 25079
rect 14105 25067 14139 25079
rect 13969 25045 13972 25067
rect 14037 25045 14044 25067
rect 14105 25045 14116 25067
rect 14173 25045 14233 25079
rect 9877 25033 13756 25045
rect 13790 25033 13828 25045
rect 13862 25033 13900 25045
rect 13934 25033 13972 25045
rect 14006 25033 14044 25045
rect 14078 25033 14116 25045
rect 14150 25033 14233 25045
rect 9877 25009 14233 25033
rect 9877 24975 9911 25009
rect 9945 24975 9980 25009
rect 10014 24975 10049 25009
rect 10083 24975 10118 25009
rect 10152 24975 10187 25009
rect 10221 24975 10256 25009
rect 10290 24975 10325 25009
rect 10359 24975 10394 25009
rect 10428 24975 10463 25009
rect 10497 24975 10532 25009
rect 10566 24975 10601 25009
rect 10635 24975 10670 25009
rect 10704 24975 10739 25009
rect 10773 24975 10807 25009
rect 10841 24975 10875 25009
rect 10909 24975 10943 25009
rect 10977 24975 11011 25009
rect 11045 24975 11079 25009
rect 11113 24975 11147 25009
rect 11181 24975 11215 25009
rect 11249 24975 11283 25009
rect 11317 24975 11351 25009
rect 11385 24975 11419 25009
rect 11453 24975 11487 25009
rect 11521 24975 11555 25009
rect 11589 24975 11623 25009
rect 11657 24975 11691 25009
rect 11725 24975 11759 25009
rect 11793 24975 11827 25009
rect 11861 24975 11895 25009
rect 11929 24975 11963 25009
rect 11997 24975 12031 25009
rect 12065 24975 12099 25009
rect 12133 24975 12167 25009
rect 12201 24975 12235 25009
rect 12269 24975 12303 25009
rect 12337 24975 12371 25009
rect 12405 24975 12439 25009
rect 12473 24975 12507 25009
rect 12541 24975 12575 25009
rect 12609 24975 12643 25009
rect 12677 24975 12711 25009
rect 12745 24975 12779 25009
rect 12813 24975 12847 25009
rect 12881 24975 12915 25009
rect 12949 24975 12983 25009
rect 13017 24975 13051 25009
rect 13085 24975 13119 25009
rect 13153 24975 13187 25009
rect 13221 24975 13255 25009
rect 13289 24975 13323 25009
rect 13357 24975 13391 25009
rect 13425 24975 13459 25009
rect 13493 24975 13527 25009
rect 13561 24975 13595 25009
rect 13629 24975 13663 25009
rect 13697 24975 13731 25009
rect 13765 24975 13799 25009
rect 13833 24975 13867 25009
rect 13901 24975 13935 25009
rect 13969 24975 14003 25009
rect 14037 24975 14071 25009
rect 14105 24975 14139 25009
rect 14173 24975 14233 25009
rect 9877 24939 14233 24975
rect 9877 24905 9911 24939
rect 9945 24905 9980 24939
rect 10014 24905 10049 24939
rect 10083 24905 10118 24939
rect 10152 24905 10187 24939
rect 10221 24905 10256 24939
rect 10290 24905 10325 24939
rect 10359 24905 10394 24939
rect 10428 24905 10463 24939
rect 10497 24905 10532 24939
rect 10566 24905 10601 24939
rect 10635 24905 10670 24939
rect 10704 24905 10739 24939
rect 10773 24905 10807 24939
rect 10841 24905 10875 24939
rect 10909 24905 10943 24939
rect 10977 24905 11011 24939
rect 11045 24905 11079 24939
rect 11113 24905 11147 24939
rect 11181 24905 11215 24939
rect 11249 24905 11283 24939
rect 11317 24905 11351 24939
rect 11385 24905 11419 24939
rect 11453 24905 11487 24939
rect 11521 24905 11555 24939
rect 11589 24905 11623 24939
rect 11657 24905 11691 24939
rect 11725 24905 11759 24939
rect 11793 24905 11827 24939
rect 11861 24905 11895 24939
rect 11929 24905 11963 24939
rect 11997 24905 12031 24939
rect 12065 24905 12099 24939
rect 12133 24905 12167 24939
rect 12201 24905 12235 24939
rect 12269 24905 12303 24939
rect 12337 24905 12371 24939
rect 12405 24905 12439 24939
rect 12473 24905 12507 24939
rect 12541 24905 12575 24939
rect 12609 24905 12643 24939
rect 12677 24905 12711 24939
rect 12745 24905 12779 24939
rect 12813 24905 12847 24939
rect 12881 24905 12915 24939
rect 12949 24905 12983 24939
rect 13017 24905 13051 24939
rect 13085 24905 13119 24939
rect 13153 24905 13187 24939
rect 13221 24905 13255 24939
rect 13289 24905 13323 24939
rect 13357 24905 13391 24939
rect 13425 24905 13459 24939
rect 13493 24905 13527 24939
rect 13561 24905 13595 24939
rect 13629 24905 13663 24939
rect 13697 24905 13731 24939
rect 13765 24905 13799 24939
rect 13833 24905 13867 24939
rect 13901 24905 13935 24939
rect 13969 24905 14003 24939
rect 14037 24905 14071 24939
rect 14105 24905 14139 24939
rect 14173 24905 14233 24939
rect 9877 24822 14233 24905
rect 9877 24821 11232 24822
rect 9877 24787 9911 24821
rect 9945 24787 9981 24821
rect 10015 24787 10051 24821
rect 10085 24787 10121 24821
rect 10155 24787 10191 24821
rect 10225 24787 10261 24821
rect 10295 24787 10331 24821
rect 10365 24787 10401 24821
rect 10435 24787 10471 24821
rect 10505 24787 10541 24821
rect 10575 24787 10611 24821
rect 10645 24787 10681 24821
rect 10715 24787 10750 24821
rect 10784 24787 10819 24821
rect 10853 24787 10888 24821
rect 10922 24787 10957 24821
rect 10991 24787 11026 24821
rect 11060 24787 11095 24821
rect 11129 24787 11164 24821
rect 11198 24787 11232 24821
rect 9877 24753 11232 24787
rect 9877 24719 9911 24753
rect 9945 24719 9981 24753
rect 10015 24719 10051 24753
rect 10085 24719 10121 24753
rect 10155 24719 10191 24753
rect 10225 24719 10261 24753
rect 10295 24719 10331 24753
rect 10365 24719 10401 24753
rect 10435 24719 10471 24753
rect 10505 24719 10541 24753
rect 10575 24719 10611 24753
rect 10645 24719 10681 24753
rect 10715 24719 10750 24753
rect 10784 24719 10819 24753
rect 10853 24719 10888 24753
rect 10922 24719 10957 24753
rect 10991 24719 11026 24753
rect 11060 24719 11095 24753
rect 11129 24719 11164 24753
rect 11198 24719 11232 24753
rect 9877 24685 11232 24719
rect 9877 24651 9911 24685
rect 9945 24651 9981 24685
rect 10015 24651 10051 24685
rect 10085 24651 10121 24685
rect 10155 24651 10191 24685
rect 10225 24651 10261 24685
rect 10295 24651 10331 24685
rect 10365 24651 10401 24685
rect 10435 24651 10471 24685
rect 10505 24651 10541 24685
rect 10575 24651 10611 24685
rect 10645 24651 10681 24685
rect 10715 24651 10750 24685
rect 10784 24651 10819 24685
rect 10853 24651 10888 24685
rect 10922 24651 10957 24685
rect 10991 24651 11026 24685
rect 11060 24651 11095 24685
rect 11129 24651 11164 24685
rect 11198 24651 11232 24685
rect 9877 24617 11232 24651
rect 9877 24583 9911 24617
rect 9945 24583 9981 24617
rect 10015 24583 10051 24617
rect 10085 24583 10121 24617
rect 10155 24583 10191 24617
rect 10225 24583 10261 24617
rect 10295 24583 10331 24617
rect 10365 24583 10401 24617
rect 10435 24583 10471 24617
rect 10505 24583 10541 24617
rect 10575 24583 10611 24617
rect 10645 24583 10681 24617
rect 10715 24583 10750 24617
rect 10784 24583 10819 24617
rect 10853 24583 10888 24617
rect 10922 24583 10957 24617
rect 10991 24583 11026 24617
rect 11060 24583 11095 24617
rect 11129 24583 11164 24617
rect 11198 24583 11232 24617
rect 9877 24562 11232 24583
rect 9877 24549 9914 24562
rect 9948 24549 9990 24562
rect 10024 24549 10066 24562
rect 10100 24549 10142 24562
rect 10176 24549 10218 24562
rect 10252 24549 10294 24562
rect 10328 24549 10369 24562
rect 10403 24549 10444 24562
rect 10478 24549 10519 24562
rect 10553 24549 10594 24562
rect 10628 24549 10669 24562
rect 10703 24549 10744 24562
rect 10778 24549 10819 24562
rect 10853 24549 10894 24562
rect 10928 24549 10969 24562
rect 11003 24549 11044 24562
rect 11078 24549 11119 24562
rect 11153 24549 11194 24562
rect 9877 24515 9911 24549
rect 9948 24528 9981 24549
rect 10024 24528 10051 24549
rect 10100 24528 10121 24549
rect 10176 24528 10191 24549
rect 10252 24528 10261 24549
rect 10328 24528 10331 24549
rect 9945 24515 9981 24528
rect 10015 24515 10051 24528
rect 10085 24515 10121 24528
rect 10155 24515 10191 24528
rect 10225 24515 10261 24528
rect 10295 24515 10331 24528
rect 10365 24528 10369 24549
rect 10435 24528 10444 24549
rect 10505 24528 10519 24549
rect 10575 24528 10594 24549
rect 10645 24528 10669 24549
rect 10715 24528 10744 24549
rect 10365 24515 10401 24528
rect 10435 24515 10471 24528
rect 10505 24515 10541 24528
rect 10575 24515 10611 24528
rect 10645 24515 10681 24528
rect 10715 24515 10750 24528
rect 10784 24515 10819 24549
rect 10853 24515 10888 24549
rect 10928 24528 10957 24549
rect 11003 24528 11026 24549
rect 11078 24528 11095 24549
rect 11153 24528 11164 24549
rect 11228 24528 11232 24562
rect 10922 24515 10957 24528
rect 10991 24515 11026 24528
rect 11060 24515 11095 24528
rect 11129 24515 11164 24528
rect 11198 24515 11232 24528
rect 9877 24490 11232 24515
rect 9877 24481 9914 24490
rect 9948 24481 9990 24490
rect 10024 24481 10066 24490
rect 10100 24481 10142 24490
rect 10176 24481 10218 24490
rect 10252 24481 10294 24490
rect 10328 24481 10369 24490
rect 10403 24481 10444 24490
rect 10478 24481 10519 24490
rect 10553 24481 10594 24490
rect 10628 24481 10669 24490
rect 10703 24481 10744 24490
rect 10778 24481 10819 24490
rect 10853 24481 10894 24490
rect 10928 24481 10969 24490
rect 11003 24481 11044 24490
rect 11078 24481 11119 24490
rect 11153 24481 11194 24490
rect 9877 24447 9911 24481
rect 9948 24456 9981 24481
rect 10024 24456 10051 24481
rect 10100 24456 10121 24481
rect 10176 24456 10191 24481
rect 10252 24456 10261 24481
rect 10328 24456 10331 24481
rect 9945 24447 9981 24456
rect 10015 24447 10051 24456
rect 10085 24447 10121 24456
rect 10155 24447 10191 24456
rect 10225 24447 10261 24456
rect 10295 24447 10331 24456
rect 10365 24456 10369 24481
rect 10435 24456 10444 24481
rect 10505 24456 10519 24481
rect 10575 24456 10594 24481
rect 10645 24456 10669 24481
rect 10715 24456 10744 24481
rect 10365 24447 10401 24456
rect 10435 24447 10471 24456
rect 10505 24447 10541 24456
rect 10575 24447 10611 24456
rect 10645 24447 10681 24456
rect 10715 24447 10750 24456
rect 10784 24447 10819 24481
rect 10853 24447 10888 24481
rect 10928 24456 10957 24481
rect 11003 24456 11026 24481
rect 11078 24456 11095 24481
rect 11153 24456 11164 24481
rect 11228 24456 11232 24490
rect 10922 24447 10957 24456
rect 10991 24447 11026 24456
rect 11060 24447 11095 24456
rect 11129 24447 11164 24456
rect 11198 24447 11232 24456
rect 9877 24418 11232 24447
rect 9877 24413 9914 24418
rect 9948 24413 9990 24418
rect 10024 24413 10066 24418
rect 10100 24413 10142 24418
rect 10176 24413 10218 24418
rect 10252 24413 10294 24418
rect 10328 24413 10369 24418
rect 10403 24413 10444 24418
rect 10478 24413 10519 24418
rect 10553 24413 10594 24418
rect 10628 24413 10669 24418
rect 10703 24413 10744 24418
rect 10778 24413 10819 24418
rect 10853 24413 10894 24418
rect 10928 24413 10969 24418
rect 11003 24413 11044 24418
rect 11078 24413 11119 24418
rect 11153 24413 11194 24418
rect 9877 24379 9911 24413
rect 9948 24384 9981 24413
rect 10024 24384 10051 24413
rect 10100 24384 10121 24413
rect 10176 24384 10191 24413
rect 10252 24384 10261 24413
rect 10328 24384 10331 24413
rect 9945 24379 9981 24384
rect 10015 24379 10051 24384
rect 10085 24379 10121 24384
rect 10155 24379 10191 24384
rect 10225 24379 10261 24384
rect 10295 24379 10331 24384
rect 10365 24384 10369 24413
rect 10435 24384 10444 24413
rect 10505 24384 10519 24413
rect 10575 24384 10594 24413
rect 10645 24384 10669 24413
rect 10715 24384 10744 24413
rect 10365 24379 10401 24384
rect 10435 24379 10471 24384
rect 10505 24379 10541 24384
rect 10575 24379 10611 24384
rect 10645 24379 10681 24384
rect 10715 24379 10750 24384
rect 10784 24379 10819 24413
rect 10853 24379 10888 24413
rect 10928 24384 10957 24413
rect 11003 24384 11026 24413
rect 11078 24384 11095 24413
rect 11153 24384 11164 24413
rect 11228 24384 11232 24418
rect 10922 24379 10957 24384
rect 10991 24379 11026 24384
rect 11060 24379 11095 24384
rect 11129 24379 11164 24384
rect 11198 24379 11232 24384
rect 9877 24346 11232 24379
rect 9877 24345 9914 24346
rect 9948 24345 9990 24346
rect 10024 24345 10066 24346
rect 10100 24345 10142 24346
rect 10176 24345 10218 24346
rect 10252 24345 10294 24346
rect 10328 24345 10369 24346
rect 10403 24345 10444 24346
rect 10478 24345 10519 24346
rect 10553 24345 10594 24346
rect 10628 24345 10669 24346
rect 10703 24345 10744 24346
rect 10778 24345 10819 24346
rect 10853 24345 10894 24346
rect 10928 24345 10969 24346
rect 11003 24345 11044 24346
rect 11078 24345 11119 24346
rect 11153 24345 11194 24346
rect 9877 24311 9911 24345
rect 9948 24312 9981 24345
rect 10024 24312 10051 24345
rect 10100 24312 10121 24345
rect 10176 24312 10191 24345
rect 10252 24312 10261 24345
rect 10328 24312 10331 24345
rect 9945 24311 9981 24312
rect 10015 24311 10051 24312
rect 10085 24311 10121 24312
rect 10155 24311 10191 24312
rect 10225 24311 10261 24312
rect 10295 24311 10331 24312
rect 10365 24312 10369 24345
rect 10435 24312 10444 24345
rect 10505 24312 10519 24345
rect 10575 24312 10594 24345
rect 10645 24312 10669 24345
rect 10715 24312 10744 24345
rect 10365 24311 10401 24312
rect 10435 24311 10471 24312
rect 10505 24311 10541 24312
rect 10575 24311 10611 24312
rect 10645 24311 10681 24312
rect 10715 24311 10750 24312
rect 10784 24311 10819 24345
rect 10853 24311 10888 24345
rect 10928 24312 10957 24345
rect 11003 24312 11026 24345
rect 11078 24312 11095 24345
rect 11153 24312 11164 24345
rect 11228 24312 11232 24346
rect 10922 24311 10957 24312
rect 10991 24311 11026 24312
rect 11060 24311 11095 24312
rect 11129 24311 11164 24312
rect 11198 24311 11232 24312
rect 9877 24277 11232 24311
rect 9877 24243 9911 24277
rect 9945 24274 9981 24277
rect 10015 24274 10051 24277
rect 10085 24274 10121 24277
rect 10155 24274 10191 24277
rect 10225 24274 10261 24277
rect 10295 24274 10331 24277
rect 9948 24243 9981 24274
rect 10024 24243 10051 24274
rect 10100 24243 10121 24274
rect 10176 24243 10191 24274
rect 10252 24243 10261 24274
rect 10328 24243 10331 24274
rect 10365 24274 10401 24277
rect 10435 24274 10471 24277
rect 10505 24274 10541 24277
rect 10575 24274 10611 24277
rect 10645 24274 10681 24277
rect 10715 24274 10750 24277
rect 10365 24243 10369 24274
rect 10435 24243 10444 24274
rect 10505 24243 10519 24274
rect 10575 24243 10594 24274
rect 10645 24243 10669 24274
rect 10715 24243 10744 24274
rect 10784 24243 10819 24277
rect 10853 24243 10888 24277
rect 10922 24274 10957 24277
rect 10991 24274 11026 24277
rect 11060 24274 11095 24277
rect 11129 24274 11164 24277
rect 11198 24274 11232 24277
rect 10928 24243 10957 24274
rect 11003 24243 11026 24274
rect 11078 24243 11095 24274
rect 11153 24243 11164 24274
rect 9877 24240 9914 24243
rect 9948 24240 9990 24243
rect 10024 24240 10066 24243
rect 10100 24240 10142 24243
rect 10176 24240 10218 24243
rect 10252 24240 10294 24243
rect 10328 24240 10369 24243
rect 10403 24240 10444 24243
rect 10478 24240 10519 24243
rect 10553 24240 10594 24243
rect 10628 24240 10669 24243
rect 10703 24240 10744 24243
rect 10778 24240 10819 24243
rect 10853 24240 10894 24243
rect 10928 24240 10969 24243
rect 11003 24240 11044 24243
rect 11078 24240 11119 24243
rect 11153 24240 11194 24243
rect 11228 24240 11232 24274
rect 9877 24209 11232 24240
rect 9877 24176 10825 24209
rect 9877 24171 9914 24176
rect 9948 24171 9984 24176
rect 9877 24137 9905 24171
rect 9948 24142 9981 24171
rect 10018 24142 10054 24176
rect 10088 24171 10124 24176
rect 10158 24171 10194 24176
rect 10228 24171 10264 24176
rect 10298 24171 10334 24176
rect 10368 24171 10404 24176
rect 10438 24171 10474 24176
rect 10091 24142 10124 24171
rect 10167 24142 10194 24171
rect 10243 24142 10264 24171
rect 10319 24142 10334 24171
rect 10395 24142 10404 24171
rect 10471 24142 10474 24171
rect 10508 24171 10544 24176
rect 10578 24171 10614 24176
rect 10648 24171 10684 24176
rect 10508 24142 10513 24171
rect 10578 24142 10589 24171
rect 10648 24142 10665 24171
rect 10718 24142 10754 24176
rect 10788 24142 10825 24176
rect 9939 24137 9981 24142
rect 10015 24137 10057 24142
rect 10091 24137 10133 24142
rect 10167 24137 10209 24142
rect 10243 24137 10285 24142
rect 10319 24137 10361 24142
rect 10395 24137 10437 24142
rect 10471 24137 10513 24142
rect 10547 24137 10589 24142
rect 10623 24137 10665 24142
rect 10699 24137 10825 24142
rect 9877 24108 10825 24137
rect 9877 24097 9914 24108
rect 9948 24097 9984 24108
rect 9877 24063 9905 24097
rect 9948 24074 9981 24097
rect 10018 24074 10054 24108
rect 10088 24097 10124 24108
rect 10158 24097 10194 24108
rect 10228 24097 10264 24108
rect 10298 24097 10334 24108
rect 10368 24097 10404 24108
rect 10438 24097 10474 24108
rect 10091 24074 10124 24097
rect 10167 24074 10194 24097
rect 10243 24074 10264 24097
rect 10319 24074 10334 24097
rect 10395 24074 10404 24097
rect 10471 24074 10474 24097
rect 10508 24097 10544 24108
rect 10578 24097 10614 24108
rect 10648 24097 10684 24108
rect 10508 24074 10513 24097
rect 10578 24074 10589 24097
rect 10648 24074 10665 24097
rect 10718 24074 10754 24108
rect 10788 24074 10825 24108
rect 9939 24063 9981 24074
rect 10015 24063 10057 24074
rect 10091 24063 10133 24074
rect 10167 24063 10209 24074
rect 10243 24063 10285 24074
rect 10319 24063 10361 24074
rect 10395 24063 10437 24074
rect 10471 24063 10513 24074
rect 10547 24063 10589 24074
rect 10623 24063 10665 24074
rect 10699 24063 10825 24074
rect 9877 24040 10825 24063
rect 9877 24023 9914 24040
rect 9948 24023 9984 24040
rect 9877 23989 9905 24023
rect 9948 24006 9981 24023
rect 10018 24006 10054 24040
rect 10088 24023 10124 24040
rect 10158 24023 10194 24040
rect 10228 24023 10264 24040
rect 10298 24023 10334 24040
rect 10368 24023 10404 24040
rect 10438 24023 10474 24040
rect 10091 24006 10124 24023
rect 10167 24006 10194 24023
rect 10243 24006 10264 24023
rect 10319 24006 10334 24023
rect 10395 24006 10404 24023
rect 10471 24006 10474 24023
rect 10508 24023 10544 24040
rect 10578 24023 10614 24040
rect 10648 24023 10684 24040
rect 10508 24006 10513 24023
rect 10578 24006 10589 24023
rect 10648 24006 10665 24023
rect 10718 24006 10754 24040
rect 10788 24006 10825 24040
rect 9939 23989 9981 24006
rect 10015 23989 10057 24006
rect 10091 23989 10133 24006
rect 10167 23989 10209 24006
rect 10243 23989 10285 24006
rect 10319 23989 10361 24006
rect 10395 23989 10437 24006
rect 10471 23989 10513 24006
rect 10547 23989 10589 24006
rect 10623 23989 10665 24006
rect 10699 23989 10825 24006
rect 9877 23971 10825 23989
rect 9877 23949 9914 23971
rect 9948 23949 9984 23971
rect 9877 23915 9905 23949
rect 9948 23937 9981 23949
rect 10018 23937 10054 23971
rect 10088 23949 10124 23971
rect 10158 23949 10194 23971
rect 10228 23949 10264 23971
rect 10298 23949 10334 23971
rect 10368 23949 10404 23971
rect 10438 23949 10474 23971
rect 10091 23937 10124 23949
rect 10167 23937 10194 23949
rect 10243 23937 10264 23949
rect 10319 23937 10334 23949
rect 10395 23937 10404 23949
rect 10471 23937 10474 23949
rect 10508 23949 10544 23971
rect 10578 23949 10614 23971
rect 10648 23949 10684 23971
rect 10508 23937 10513 23949
rect 10578 23937 10589 23949
rect 10648 23937 10665 23949
rect 10718 23937 10754 23971
rect 10788 23937 10825 23971
rect 9939 23915 9981 23937
rect 10015 23915 10057 23937
rect 10091 23915 10133 23937
rect 10167 23915 10209 23937
rect 10243 23915 10285 23937
rect 10319 23915 10361 23937
rect 10395 23915 10437 23937
rect 10471 23915 10513 23937
rect 10547 23915 10589 23937
rect 10623 23915 10665 23937
rect 10699 23915 10825 23937
rect 9877 23902 10825 23915
rect 9877 23875 9914 23902
rect 9948 23875 9984 23902
rect 9877 23841 9905 23875
rect 9948 23868 9981 23875
rect 10018 23868 10054 23902
rect 10088 23875 10124 23902
rect 10158 23875 10194 23902
rect 10228 23875 10264 23902
rect 10298 23875 10334 23902
rect 10368 23875 10404 23902
rect 10438 23875 10474 23902
rect 10091 23868 10124 23875
rect 10167 23868 10194 23875
rect 10243 23868 10264 23875
rect 10319 23868 10334 23875
rect 10395 23868 10404 23875
rect 10471 23868 10474 23875
rect 10508 23875 10544 23902
rect 10578 23875 10614 23902
rect 10648 23875 10684 23902
rect 10508 23868 10513 23875
rect 10578 23868 10589 23875
rect 10648 23868 10665 23875
rect 10718 23868 10754 23902
rect 10788 23868 10825 23902
rect 9939 23841 9981 23868
rect 10015 23841 10057 23868
rect 10091 23841 10133 23868
rect 10167 23841 10209 23868
rect 10243 23841 10285 23868
rect 10319 23841 10361 23868
rect 10395 23841 10437 23868
rect 10471 23841 10513 23868
rect 10547 23841 10589 23868
rect 10623 23841 10665 23868
rect 10699 23841 10825 23868
rect 9877 23833 10825 23841
rect 9877 23801 9914 23833
rect 9948 23801 9984 23833
rect 9877 23767 9905 23801
rect 9948 23799 9981 23801
rect 10018 23799 10054 23833
rect 10088 23801 10124 23833
rect 10158 23801 10194 23833
rect 10228 23801 10264 23833
rect 10298 23801 10334 23833
rect 10368 23801 10404 23833
rect 10438 23801 10474 23833
rect 10091 23799 10124 23801
rect 10167 23799 10194 23801
rect 10243 23799 10264 23801
rect 10319 23799 10334 23801
rect 10395 23799 10404 23801
rect 10471 23799 10474 23801
rect 10508 23801 10544 23833
rect 10578 23801 10614 23833
rect 10648 23801 10684 23833
rect 10508 23799 10513 23801
rect 10578 23799 10589 23801
rect 10648 23799 10665 23801
rect 10718 23799 10754 23833
rect 10788 23799 10825 23833
rect 9939 23767 9981 23799
rect 10015 23767 10057 23799
rect 10091 23767 10133 23799
rect 10167 23767 10209 23799
rect 10243 23767 10285 23799
rect 10319 23767 10361 23799
rect 10395 23767 10437 23799
rect 10471 23767 10513 23799
rect 10547 23767 10589 23799
rect 10623 23767 10665 23799
rect 10699 23767 10825 23799
rect 9877 23764 10825 23767
rect 9877 23730 9914 23764
rect 9948 23730 9984 23764
rect 10018 23730 10054 23764
rect 10088 23730 10124 23764
rect 10158 23730 10194 23764
rect 10228 23730 10264 23764
rect 10298 23730 10334 23764
rect 10368 23730 10404 23764
rect 10438 23730 10474 23764
rect 10508 23730 10544 23764
rect 10578 23730 10614 23764
rect 10648 23730 10684 23764
rect 10718 23730 10754 23764
rect 10788 23730 10825 23764
rect 9877 23727 10825 23730
rect 9877 23693 9905 23727
rect 9939 23695 9981 23727
rect 10015 23695 10057 23727
rect 10091 23695 10133 23727
rect 10167 23695 10209 23727
rect 10243 23695 10285 23727
rect 10319 23695 10361 23727
rect 10395 23695 10437 23727
rect 10471 23695 10513 23727
rect 10547 23695 10589 23727
rect 10623 23695 10665 23727
rect 10699 23695 10825 23727
rect 9948 23693 9981 23695
rect 9877 23661 9914 23693
rect 9948 23661 9984 23693
rect 10018 23661 10054 23695
rect 10091 23693 10124 23695
rect 10167 23693 10194 23695
rect 10243 23693 10264 23695
rect 10319 23693 10334 23695
rect 10395 23693 10404 23695
rect 10471 23693 10474 23695
rect 10088 23661 10124 23693
rect 10158 23661 10194 23693
rect 10228 23661 10264 23693
rect 10298 23661 10334 23693
rect 10368 23661 10404 23693
rect 10438 23661 10474 23693
rect 10508 23693 10513 23695
rect 10578 23693 10589 23695
rect 10648 23693 10665 23695
rect 10508 23661 10544 23693
rect 10578 23661 10614 23693
rect 10648 23661 10684 23693
rect 10718 23661 10754 23695
rect 10788 23661 10825 23695
rect 9877 23653 10825 23661
rect 9877 23619 9905 23653
rect 9939 23626 9981 23653
rect 10015 23626 10057 23653
rect 10091 23626 10133 23653
rect 10167 23626 10209 23653
rect 10243 23626 10285 23653
rect 10319 23626 10361 23653
rect 10395 23626 10437 23653
rect 10471 23626 10513 23653
rect 10547 23626 10589 23653
rect 10623 23626 10665 23653
rect 10699 23626 10825 23653
rect 9948 23619 9981 23626
rect 9877 23592 9914 23619
rect 9948 23592 9984 23619
rect 10018 23592 10054 23626
rect 10091 23619 10124 23626
rect 10167 23619 10194 23626
rect 10243 23619 10264 23626
rect 10319 23619 10334 23626
rect 10395 23619 10404 23626
rect 10471 23619 10474 23626
rect 10088 23592 10124 23619
rect 10158 23592 10194 23619
rect 10228 23592 10264 23619
rect 10298 23592 10334 23619
rect 10368 23592 10404 23619
rect 10438 23592 10474 23619
rect 10508 23619 10513 23626
rect 10578 23619 10589 23626
rect 10648 23619 10665 23626
rect 10508 23592 10544 23619
rect 10578 23592 10614 23619
rect 10648 23592 10684 23619
rect 10718 23592 10754 23626
rect 10788 23592 10825 23626
rect 9877 23579 10825 23592
rect 9877 23545 9905 23579
rect 9939 23557 9981 23579
rect 10015 23557 10057 23579
rect 10091 23557 10133 23579
rect 10167 23557 10209 23579
rect 10243 23557 10285 23579
rect 10319 23557 10361 23579
rect 10395 23557 10437 23579
rect 10471 23557 10513 23579
rect 10547 23557 10589 23579
rect 10623 23557 10665 23579
rect 10699 23557 10825 23579
rect 9948 23545 9981 23557
rect 9877 23523 9914 23545
rect 9948 23523 9984 23545
rect 10018 23523 10054 23557
rect 10091 23545 10124 23557
rect 10167 23545 10194 23557
rect 10243 23545 10264 23557
rect 10319 23545 10334 23557
rect 10395 23545 10404 23557
rect 10471 23545 10474 23557
rect 10088 23523 10124 23545
rect 10158 23523 10194 23545
rect 10228 23523 10264 23545
rect 10298 23523 10334 23545
rect 10368 23523 10404 23545
rect 10438 23523 10474 23545
rect 10508 23545 10513 23557
rect 10578 23545 10589 23557
rect 10648 23545 10665 23557
rect 10508 23523 10544 23545
rect 10578 23523 10614 23545
rect 10648 23523 10684 23545
rect 10718 23523 10754 23557
rect 10788 23523 10825 23557
rect 9877 23505 10825 23523
rect 9877 23471 9905 23505
rect 9939 23488 9981 23505
rect 10015 23488 10057 23505
rect 10091 23488 10133 23505
rect 10167 23488 10209 23505
rect 10243 23488 10285 23505
rect 10319 23488 10361 23505
rect 10395 23488 10437 23505
rect 10471 23488 10513 23505
rect 10547 23488 10589 23505
rect 10623 23488 10665 23505
rect 10699 23488 10825 23505
rect 9948 23471 9981 23488
rect 9877 23454 9914 23471
rect 9948 23454 9984 23471
rect 10018 23454 10054 23488
rect 10091 23471 10124 23488
rect 10167 23471 10194 23488
rect 10243 23471 10264 23488
rect 10319 23471 10334 23488
rect 10395 23471 10404 23488
rect 10471 23471 10474 23488
rect 10088 23454 10124 23471
rect 10158 23454 10194 23471
rect 10228 23454 10264 23471
rect 10298 23454 10334 23471
rect 10368 23454 10404 23471
rect 10438 23454 10474 23471
rect 10508 23471 10513 23488
rect 10578 23471 10589 23488
rect 10648 23471 10665 23488
rect 10508 23454 10544 23471
rect 10578 23454 10614 23471
rect 10648 23454 10684 23471
rect 10718 23454 10754 23488
rect 10788 23454 10825 23488
rect 9877 23431 10825 23454
rect 9877 23397 9905 23431
rect 9939 23419 9981 23431
rect 10015 23419 10057 23431
rect 10091 23419 10133 23431
rect 10167 23419 10209 23431
rect 10243 23419 10285 23431
rect 10319 23419 10361 23431
rect 10395 23419 10437 23431
rect 10471 23419 10513 23431
rect 10547 23419 10589 23431
rect 10623 23419 10665 23431
rect 10699 23419 10825 23431
rect 9948 23397 9981 23419
rect 9877 23385 9914 23397
rect 9948 23385 9984 23397
rect 10018 23385 10054 23419
rect 10091 23397 10124 23419
rect 10167 23397 10194 23419
rect 10243 23397 10264 23419
rect 10319 23397 10334 23419
rect 10395 23397 10404 23419
rect 10471 23397 10474 23419
rect 10088 23385 10124 23397
rect 10158 23385 10194 23397
rect 10228 23385 10264 23397
rect 10298 23385 10334 23397
rect 10368 23385 10404 23397
rect 10438 23385 10474 23397
rect 10508 23397 10513 23419
rect 10578 23397 10589 23419
rect 10648 23397 10665 23419
rect 10508 23385 10544 23397
rect 10578 23385 10614 23397
rect 10648 23385 10684 23397
rect 10718 23385 10754 23419
rect 10788 23385 10825 23419
rect 9877 23357 10825 23385
rect 9877 23323 9905 23357
rect 9939 23350 9981 23357
rect 10015 23350 10057 23357
rect 10091 23350 10133 23357
rect 10167 23350 10209 23357
rect 10243 23350 10285 23357
rect 10319 23350 10361 23357
rect 10395 23350 10437 23357
rect 10471 23350 10513 23357
rect 10547 23350 10589 23357
rect 10623 23350 10665 23357
rect 10699 23350 10825 23357
rect 9948 23323 9981 23350
rect 9877 23316 9914 23323
rect 9948 23316 9984 23323
rect 10018 23316 10054 23350
rect 10091 23323 10124 23350
rect 10167 23323 10194 23350
rect 10243 23323 10264 23350
rect 10319 23323 10334 23350
rect 10395 23323 10404 23350
rect 10471 23323 10474 23350
rect 10088 23316 10124 23323
rect 10158 23316 10194 23323
rect 10228 23316 10264 23323
rect 10298 23316 10334 23323
rect 10368 23316 10404 23323
rect 10438 23316 10474 23323
rect 10508 23323 10513 23350
rect 10578 23323 10589 23350
rect 10648 23323 10665 23350
rect 10508 23316 10544 23323
rect 10578 23316 10614 23323
rect 10648 23316 10684 23323
rect 10718 23316 10754 23350
rect 10788 23316 10825 23350
rect 9877 23283 10825 23316
rect 9877 23249 9905 23283
rect 9939 23281 9981 23283
rect 10015 23281 10057 23283
rect 10091 23281 10133 23283
rect 10167 23281 10209 23283
rect 10243 23281 10285 23283
rect 10319 23281 10361 23283
rect 10395 23281 10437 23283
rect 10471 23281 10513 23283
rect 10547 23281 10589 23283
rect 10623 23281 10665 23283
rect 10699 23281 10825 23283
rect 9948 23249 9981 23281
rect 9877 23247 9914 23249
rect 9948 23247 9984 23249
rect 10018 23247 10054 23281
rect 10091 23249 10124 23281
rect 10167 23249 10194 23281
rect 10243 23249 10264 23281
rect 10319 23249 10334 23281
rect 10395 23249 10404 23281
rect 10471 23249 10474 23281
rect 10088 23247 10124 23249
rect 10158 23247 10194 23249
rect 10228 23247 10264 23249
rect 10298 23247 10334 23249
rect 10368 23247 10404 23249
rect 10438 23247 10474 23249
rect 10508 23249 10513 23281
rect 10578 23249 10589 23281
rect 10648 23249 10665 23281
rect 10508 23247 10544 23249
rect 10578 23247 10614 23249
rect 10648 23247 10684 23249
rect 10718 23247 10754 23281
rect 10788 23247 10825 23281
rect 9877 23212 10825 23247
rect 9877 23209 9914 23212
rect 9948 23209 9984 23212
rect 9877 23175 9905 23209
rect 9948 23178 9981 23209
rect 10018 23178 10054 23212
rect 10088 23209 10124 23212
rect 10158 23209 10194 23212
rect 10228 23209 10264 23212
rect 10298 23209 10334 23212
rect 10368 23209 10404 23212
rect 10438 23209 10474 23212
rect 10091 23178 10124 23209
rect 10167 23178 10194 23209
rect 10243 23178 10264 23209
rect 10319 23178 10334 23209
rect 10395 23178 10404 23209
rect 10471 23178 10474 23209
rect 10508 23209 10544 23212
rect 10578 23209 10614 23212
rect 10648 23209 10684 23212
rect 10508 23178 10513 23209
rect 10578 23178 10589 23209
rect 10648 23178 10665 23209
rect 10718 23178 10754 23212
rect 10788 23178 10825 23212
rect 9939 23175 9981 23178
rect 10015 23175 10057 23178
rect 10091 23175 10133 23178
rect 10167 23175 10209 23178
rect 10243 23175 10285 23178
rect 10319 23175 10361 23178
rect 10395 23175 10437 23178
rect 10471 23175 10513 23178
rect 10547 23175 10589 23178
rect 10623 23175 10665 23178
rect 10699 23175 10825 23178
rect 9877 23143 10825 23175
rect 9877 23135 9914 23143
rect 9948 23135 9984 23143
rect 9877 23101 9905 23135
rect 9948 23109 9981 23135
rect 10018 23109 10054 23143
rect 10088 23135 10124 23143
rect 10158 23135 10194 23143
rect 10228 23135 10264 23143
rect 10298 23135 10334 23143
rect 10368 23135 10404 23143
rect 10438 23135 10474 23143
rect 10091 23109 10124 23135
rect 10167 23109 10194 23135
rect 10243 23109 10264 23135
rect 10319 23109 10334 23135
rect 10395 23109 10404 23135
rect 10471 23109 10474 23135
rect 10508 23135 10544 23143
rect 10578 23135 10614 23143
rect 10648 23135 10684 23143
rect 10508 23109 10513 23135
rect 10578 23109 10589 23135
rect 10648 23109 10665 23135
rect 10718 23109 10754 23143
rect 10788 23109 10825 23143
rect 9939 23101 9981 23109
rect 10015 23101 10057 23109
rect 10091 23101 10133 23109
rect 10167 23101 10209 23109
rect 10243 23101 10285 23109
rect 10319 23101 10361 23109
rect 10395 23101 10437 23109
rect 10471 23101 10513 23109
rect 10547 23101 10589 23109
rect 10623 23101 10665 23109
rect 10699 23101 10825 23109
rect 9877 23074 10825 23101
rect 9877 23061 9914 23074
rect 9948 23061 9984 23074
rect 9877 23027 9905 23061
rect 9948 23040 9981 23061
rect 10018 23040 10054 23074
rect 10088 23061 10124 23074
rect 10158 23061 10194 23074
rect 10228 23061 10264 23074
rect 10298 23061 10334 23074
rect 10368 23061 10404 23074
rect 10438 23061 10474 23074
rect 10091 23040 10124 23061
rect 10167 23040 10194 23061
rect 10243 23040 10264 23061
rect 10319 23040 10334 23061
rect 10395 23040 10404 23061
rect 10471 23040 10474 23061
rect 10508 23061 10544 23074
rect 10578 23061 10614 23074
rect 10648 23061 10684 23074
rect 10508 23040 10513 23061
rect 10578 23040 10589 23061
rect 10648 23040 10665 23061
rect 10718 23040 10754 23074
rect 10788 23045 10825 23074
rect 14146 24150 14233 24822
rect 14403 24150 14429 26224
rect 14146 24146 14429 24150
rect 14146 24115 14252 24146
rect 14286 24115 14324 24146
rect 14358 24115 14429 24146
rect 14146 24081 14233 24115
rect 14286 24112 14301 24115
rect 14358 24112 14369 24115
rect 14267 24081 14301 24112
rect 14335 24081 14369 24112
rect 14403 24081 14429 24115
rect 14146 24073 14429 24081
rect 14146 24046 14252 24073
rect 14286 24046 14324 24073
rect 14358 24046 14429 24073
rect 14146 24012 14233 24046
rect 14286 24039 14301 24046
rect 14358 24039 14369 24046
rect 14267 24012 14301 24039
rect 14335 24012 14369 24039
rect 14403 24012 14429 24046
rect 14146 24000 14429 24012
rect 14146 23977 14252 24000
rect 14286 23977 14324 24000
rect 14358 23977 14429 24000
rect 14146 23943 14233 23977
rect 14286 23966 14301 23977
rect 14358 23966 14369 23977
rect 14267 23943 14301 23966
rect 14335 23943 14369 23966
rect 14403 23943 14429 23977
rect 14146 23927 14429 23943
rect 14146 23908 14252 23927
rect 14286 23908 14324 23927
rect 14358 23908 14429 23927
rect 14146 23874 14233 23908
rect 14286 23893 14301 23908
rect 14358 23893 14369 23908
rect 14267 23874 14301 23893
rect 14335 23874 14369 23893
rect 14403 23874 14429 23908
rect 14146 23854 14429 23874
rect 14146 23839 14252 23854
rect 14286 23839 14324 23854
rect 14358 23839 14429 23854
rect 14146 23805 14233 23839
rect 14286 23820 14301 23839
rect 14358 23820 14369 23839
rect 14267 23805 14301 23820
rect 14335 23805 14369 23820
rect 14403 23805 14429 23839
rect 14146 23781 14429 23805
rect 14146 23770 14252 23781
rect 14286 23770 14324 23781
rect 14358 23770 14429 23781
rect 14146 23736 14233 23770
rect 14286 23747 14301 23770
rect 14358 23747 14369 23770
rect 14267 23736 14301 23747
rect 14335 23736 14369 23747
rect 14403 23736 14429 23770
rect 14146 23708 14429 23736
rect 14146 23701 14252 23708
rect 14286 23701 14324 23708
rect 14358 23701 14429 23708
rect 14146 23667 14233 23701
rect 14286 23674 14301 23701
rect 14358 23674 14369 23701
rect 14267 23667 14301 23674
rect 14335 23667 14369 23674
rect 14403 23667 14429 23701
rect 14146 23635 14429 23667
rect 14146 23632 14252 23635
rect 14286 23632 14324 23635
rect 14358 23632 14429 23635
rect 14146 23598 14233 23632
rect 14286 23601 14301 23632
rect 14358 23601 14369 23632
rect 14267 23598 14301 23601
rect 14335 23598 14369 23601
rect 14403 23598 14429 23632
rect 14146 23563 14429 23598
rect 14146 23529 14233 23563
rect 14267 23562 14301 23563
rect 14335 23562 14369 23563
rect 14286 23529 14301 23562
rect 14358 23529 14369 23562
rect 14403 23529 14429 23563
rect 14146 23528 14252 23529
rect 14286 23528 14324 23529
rect 14358 23528 14429 23529
rect 14146 23494 14429 23528
rect 14146 23460 14233 23494
rect 14267 23489 14301 23494
rect 14335 23489 14369 23494
rect 14286 23460 14301 23489
rect 14358 23460 14369 23489
rect 14403 23460 14429 23494
rect 14146 23455 14252 23460
rect 14286 23455 14324 23460
rect 14358 23455 14429 23460
rect 14146 23425 14429 23455
rect 14146 23391 14233 23425
rect 14267 23416 14301 23425
rect 14335 23416 14369 23425
rect 14286 23391 14301 23416
rect 14358 23391 14369 23416
rect 14403 23391 14429 23425
rect 14146 23382 14252 23391
rect 14286 23382 14324 23391
rect 14358 23382 14429 23391
rect 14146 23356 14429 23382
rect 14146 23322 14233 23356
rect 14267 23343 14301 23356
rect 14335 23343 14369 23356
rect 14286 23322 14301 23343
rect 14358 23322 14369 23343
rect 14403 23322 14429 23356
rect 14146 23309 14252 23322
rect 14286 23309 14324 23322
rect 14358 23309 14429 23322
rect 14146 23287 14429 23309
rect 14146 23253 14233 23287
rect 14267 23270 14301 23287
rect 14335 23270 14369 23287
rect 14286 23253 14301 23270
rect 14358 23253 14369 23270
rect 14403 23253 14429 23287
rect 14146 23236 14252 23253
rect 14286 23236 14324 23253
rect 14358 23236 14429 23253
rect 14146 23218 14429 23236
rect 14146 23184 14233 23218
rect 14267 23197 14301 23218
rect 14335 23197 14369 23218
rect 14286 23184 14301 23197
rect 14358 23184 14369 23197
rect 14403 23184 14429 23218
rect 14146 23163 14252 23184
rect 14286 23163 14324 23184
rect 14358 23163 14429 23184
rect 14146 23149 14429 23163
rect 14146 23115 14233 23149
rect 14267 23124 14301 23149
rect 14335 23124 14369 23149
rect 14286 23115 14301 23124
rect 14358 23115 14369 23124
rect 14403 23115 14429 23149
rect 14146 23090 14252 23115
rect 14286 23090 14324 23115
rect 14358 23090 14429 23115
rect 14146 23080 14429 23090
rect 14146 23046 14233 23080
rect 14267 23051 14301 23080
rect 14335 23051 14369 23080
rect 14286 23046 14301 23051
rect 14358 23046 14369 23051
rect 14403 23046 14429 23080
rect 14146 23045 14252 23046
rect 10788 23040 14252 23045
rect 9939 23027 9981 23040
rect 10015 23027 10057 23040
rect 10091 23027 10133 23040
rect 10167 23027 10209 23040
rect 10243 23027 10285 23040
rect 10319 23027 10361 23040
rect 10395 23027 10437 23040
rect 10471 23027 10513 23040
rect 10547 23027 10589 23040
rect 10623 23027 10665 23040
rect 10699 23027 14252 23040
rect 9877 23017 14252 23027
rect 14286 23017 14324 23046
rect 14358 23017 14429 23046
rect 9877 23011 14429 23017
rect 9877 23005 14233 23011
rect 9877 22987 9914 23005
rect 9948 22987 9984 23005
rect 9877 22953 9905 22987
rect 9948 22971 9981 22987
rect 10018 22971 10054 23005
rect 10088 22987 10124 23005
rect 10158 22987 10194 23005
rect 10228 22987 10264 23005
rect 10298 22987 10334 23005
rect 10368 22987 10404 23005
rect 10438 22987 10474 23005
rect 10091 22971 10124 22987
rect 10167 22971 10194 22987
rect 10243 22971 10264 22987
rect 10319 22971 10334 22987
rect 10395 22971 10404 22987
rect 10471 22971 10474 22987
rect 10508 22987 10544 23005
rect 10578 22987 10614 23005
rect 10648 22987 10684 23005
rect 10508 22971 10513 22987
rect 10578 22971 10589 22987
rect 10648 22971 10665 22987
rect 10718 22971 10754 23005
rect 10788 23003 14233 23005
rect 10788 23000 10859 23003
rect 10893 23000 10928 23003
rect 10962 23000 10997 23003
rect 11031 23000 11066 23003
rect 11100 23000 11135 23003
rect 11169 23000 11204 23003
rect 11238 23000 11273 23003
rect 9939 22953 9981 22971
rect 10015 22953 10057 22971
rect 10091 22953 10133 22971
rect 10167 22953 10209 22971
rect 10243 22953 10285 22971
rect 10319 22953 10361 22971
rect 10395 22953 10437 22971
rect 10471 22953 10513 22971
rect 10547 22953 10589 22971
rect 10623 22953 10665 22971
rect 10699 22966 10759 22971
rect 10793 22966 10832 23000
rect 10893 22969 10905 23000
rect 10962 22969 10978 23000
rect 11031 22969 11051 23000
rect 11100 22969 11124 23000
rect 11169 22969 11197 23000
rect 11238 22969 11270 23000
rect 11307 22969 11342 23003
rect 11376 23000 11411 23003
rect 11445 23000 11480 23003
rect 11514 23000 11549 23003
rect 11583 23000 11618 23003
rect 11652 23000 11687 23003
rect 11721 23000 11756 23003
rect 11790 23000 11825 23003
rect 11859 23000 11894 23003
rect 11928 23000 11963 23003
rect 11997 23000 12031 23003
rect 11377 22969 11411 23000
rect 11450 22969 11480 23000
rect 11523 22969 11549 23000
rect 11596 22969 11618 23000
rect 11669 22969 11687 23000
rect 11741 22969 11756 23000
rect 11813 22969 11825 23000
rect 11885 22969 11894 23000
rect 11957 22969 11963 23000
rect 12029 22969 12031 23000
rect 12065 23000 12099 23003
rect 12133 23000 12167 23003
rect 12201 23000 12235 23003
rect 12065 22969 12067 23000
rect 12133 22969 12139 23000
rect 12201 22969 12211 23000
rect 12269 22969 12303 23003
rect 12337 22969 12371 23003
rect 12405 22969 12439 23003
rect 12473 22984 12507 23003
rect 12541 22984 12575 23003
rect 12609 22984 12643 23003
rect 12677 22984 12711 23003
rect 12745 22984 12779 23003
rect 12813 22984 12847 23003
rect 12473 22969 12476 22984
rect 12541 22969 12550 22984
rect 12609 22969 12624 22984
rect 12677 22969 12698 22984
rect 12745 22969 12772 22984
rect 12813 22969 12846 22984
rect 12881 22969 12915 23003
rect 12949 22984 12983 23003
rect 13017 22984 13051 23003
rect 13085 22984 13119 23003
rect 13153 22984 13187 23003
rect 13221 22984 13255 23003
rect 13289 22984 13323 23003
rect 12954 22969 12983 22984
rect 13028 22969 13051 22984
rect 13102 22969 13119 22984
rect 13175 22969 13187 22984
rect 13248 22969 13255 22984
rect 13321 22969 13323 22984
rect 13357 22984 13391 23003
rect 13425 22984 13459 23003
rect 13493 22984 13527 23003
rect 13561 22984 13595 23003
rect 13629 22984 13663 23003
rect 13357 22969 13360 22984
rect 13425 22969 13433 22984
rect 13493 22969 13506 22984
rect 13561 22969 13579 22984
rect 13629 22969 13652 22984
rect 13697 22969 13731 23003
rect 13765 22999 13799 23003
rect 13833 22999 13867 23003
rect 13901 22999 14233 23003
rect 13790 22969 13799 22999
rect 13862 22969 13867 22999
rect 10866 22966 10905 22969
rect 10939 22966 10978 22969
rect 11012 22966 11051 22969
rect 11085 22966 11124 22969
rect 11158 22966 11197 22969
rect 11231 22966 11270 22969
rect 11304 22966 11343 22969
rect 11377 22966 11416 22969
rect 11450 22966 11489 22969
rect 11523 22966 11562 22969
rect 11596 22966 11635 22969
rect 11669 22966 11707 22969
rect 11741 22966 11779 22969
rect 11813 22966 11851 22969
rect 11885 22966 11923 22969
rect 11957 22966 11995 22969
rect 12029 22966 12067 22969
rect 12101 22966 12139 22969
rect 12173 22966 12211 22969
rect 12245 22966 12476 22969
rect 10699 22953 12476 22966
rect 9877 22950 12476 22953
rect 12510 22950 12550 22969
rect 12584 22950 12624 22969
rect 12658 22950 12698 22969
rect 12732 22950 12772 22969
rect 12806 22950 12846 22969
rect 12880 22950 12920 22969
rect 12954 22950 12994 22969
rect 13028 22950 13068 22969
rect 13102 22950 13141 22969
rect 13175 22950 13214 22969
rect 13248 22950 13287 22969
rect 13321 22950 13360 22969
rect 13394 22950 13433 22969
rect 13467 22950 13506 22969
rect 13540 22950 13579 22969
rect 13613 22950 13652 22969
rect 13686 22965 13756 22969
rect 13790 22965 13828 22969
rect 13862 22965 13900 22969
rect 13934 22965 13972 22999
rect 14006 22998 14044 22999
rect 14078 22998 14116 22999
rect 14150 22998 14233 22999
rect 14012 22965 14044 22998
rect 14082 22965 14116 22998
rect 14152 22977 14233 22998
rect 14267 22978 14301 23011
rect 14335 22978 14369 23011
rect 14286 22977 14301 22978
rect 14358 22977 14369 22978
rect 14403 22977 14429 23011
rect 13686 22964 13978 22965
rect 14012 22964 14048 22965
rect 14082 22964 14118 22965
rect 14152 22964 14252 22977
rect 13686 22950 14252 22964
rect 9877 22944 14252 22950
rect 14286 22944 14324 22977
rect 14358 22944 14429 22977
rect 9877 22942 14429 22944
rect 9877 22935 14233 22942
rect 9877 22901 9901 22935
rect 9935 22913 9971 22935
rect 10005 22913 10041 22935
rect 10075 22913 10111 22935
rect 10145 22913 10181 22935
rect 10215 22913 10251 22935
rect 9939 22901 9971 22913
rect 10015 22901 10041 22913
rect 10091 22901 10111 22913
rect 10167 22901 10181 22913
rect 10243 22901 10251 22913
rect 10285 22913 10321 22935
rect 9877 22879 9905 22901
rect 9939 22879 9981 22901
rect 10015 22879 10057 22901
rect 10091 22879 10133 22901
rect 10167 22879 10209 22901
rect 10243 22879 10285 22901
rect 10319 22901 10321 22913
rect 10355 22913 10391 22935
rect 10425 22913 10461 22935
rect 10495 22913 10530 22935
rect 10564 22913 10599 22935
rect 10633 22913 10668 22935
rect 10355 22901 10361 22913
rect 10425 22901 10437 22913
rect 10495 22901 10513 22913
rect 10564 22901 10589 22913
rect 10633 22901 10665 22913
rect 10702 22901 10737 22935
rect 10771 22914 10806 22935
rect 10840 22914 10875 22935
rect 10909 22914 10944 22935
rect 10793 22901 10806 22914
rect 10866 22901 10875 22914
rect 10939 22901 10944 22914
rect 10978 22914 11013 22935
rect 10319 22879 10361 22901
rect 10395 22879 10437 22901
rect 10471 22879 10513 22901
rect 10547 22879 10589 22901
rect 10623 22879 10665 22901
rect 10699 22880 10759 22901
rect 10793 22880 10832 22901
rect 10866 22880 10905 22901
rect 10939 22880 10978 22901
rect 11012 22901 11013 22914
rect 11047 22914 11082 22935
rect 11116 22914 11151 22935
rect 11185 22914 11220 22935
rect 11254 22914 11289 22935
rect 11323 22914 11358 22935
rect 11392 22914 11427 22935
rect 11461 22914 11496 22935
rect 11530 22914 11565 22935
rect 11047 22901 11051 22914
rect 11116 22901 11124 22914
rect 11185 22901 11197 22914
rect 11254 22901 11270 22914
rect 11323 22901 11343 22914
rect 11392 22901 11416 22914
rect 11461 22901 11489 22914
rect 11530 22901 11562 22914
rect 11599 22901 11634 22935
rect 11668 22914 11703 22935
rect 11737 22914 11772 22935
rect 11806 22914 11841 22935
rect 11875 22914 11910 22935
rect 11944 22914 11979 22935
rect 12013 22914 12048 22935
rect 12082 22914 12117 22935
rect 12151 22914 12186 22935
rect 12220 22914 12255 22935
rect 11669 22901 11703 22914
rect 11741 22901 11772 22914
rect 11813 22901 11841 22914
rect 11885 22901 11910 22914
rect 11957 22901 11979 22914
rect 12029 22901 12048 22914
rect 12101 22901 12117 22914
rect 12173 22901 12186 22914
rect 12245 22901 12255 22914
rect 12289 22901 12324 22935
rect 12358 22901 12393 22935
rect 12427 22927 14233 22935
rect 12427 22901 12451 22927
rect 11012 22880 11051 22901
rect 11085 22880 11124 22901
rect 11158 22880 11197 22901
rect 11231 22880 11270 22901
rect 11304 22880 11343 22901
rect 11377 22880 11416 22901
rect 11450 22880 11489 22901
rect 11523 22880 11562 22901
rect 11596 22880 11635 22901
rect 11669 22880 11707 22901
rect 11741 22880 11779 22901
rect 11813 22880 11851 22901
rect 11885 22880 11923 22901
rect 11957 22880 11995 22901
rect 12029 22880 12067 22901
rect 12101 22880 12139 22901
rect 12173 22880 12211 22901
rect 12245 22880 12451 22901
rect 10699 22879 12451 22880
rect 9877 22865 12451 22879
rect 9877 22831 9901 22865
rect 9935 22839 9971 22865
rect 10005 22839 10041 22865
rect 10075 22839 10111 22865
rect 10145 22839 10181 22865
rect 10215 22839 10251 22865
rect 9939 22831 9971 22839
rect 10015 22831 10041 22839
rect 10091 22831 10111 22839
rect 10167 22831 10181 22839
rect 10243 22831 10251 22839
rect 10285 22839 10321 22865
rect 9877 22805 9905 22831
rect 9939 22805 9981 22831
rect 10015 22805 10057 22831
rect 10091 22805 10133 22831
rect 10167 22805 10209 22831
rect 10243 22805 10285 22831
rect 10319 22831 10321 22839
rect 10355 22839 10391 22865
rect 10425 22839 10461 22865
rect 10495 22839 10530 22865
rect 10564 22839 10599 22865
rect 10633 22839 10668 22865
rect 10355 22831 10361 22839
rect 10425 22831 10437 22839
rect 10495 22831 10513 22839
rect 10564 22831 10589 22839
rect 10633 22831 10665 22839
rect 10702 22831 10737 22865
rect 10771 22831 10806 22865
rect 10840 22831 10875 22865
rect 10909 22831 10944 22865
rect 10978 22831 11013 22865
rect 11047 22831 11082 22865
rect 11116 22831 11151 22865
rect 11185 22831 11220 22865
rect 11254 22831 11289 22865
rect 11323 22831 11358 22865
rect 11392 22831 11427 22865
rect 11461 22831 11496 22865
rect 11530 22831 11565 22865
rect 11599 22831 11634 22865
rect 11668 22831 11703 22865
rect 11737 22831 11772 22865
rect 11806 22831 11841 22865
rect 11875 22831 11910 22865
rect 11944 22831 11979 22865
rect 12013 22831 12048 22865
rect 12082 22831 12117 22865
rect 12151 22831 12186 22865
rect 12220 22831 12255 22865
rect 12289 22831 12324 22865
rect 12358 22831 12393 22865
rect 12427 22831 12451 22865
rect 10319 22805 10361 22831
rect 10395 22805 10437 22831
rect 10471 22805 10513 22831
rect 10547 22805 10589 22831
rect 10623 22805 10665 22831
rect 10699 22828 12451 22831
rect 10699 22805 10759 22828
rect 9877 22795 10759 22805
rect 10793 22795 10832 22828
rect 10866 22795 10905 22828
rect 10939 22795 10978 22828
rect 9877 22761 9901 22795
rect 9935 22765 9971 22795
rect 10005 22765 10041 22795
rect 10075 22765 10111 22795
rect 10145 22765 10181 22795
rect 10215 22765 10251 22795
rect 9939 22761 9971 22765
rect 10015 22761 10041 22765
rect 10091 22761 10111 22765
rect 10167 22761 10181 22765
rect 10243 22761 10251 22765
rect 10285 22765 10321 22795
rect 9877 22731 9905 22761
rect 9939 22731 9981 22761
rect 10015 22731 10057 22761
rect 10091 22731 10133 22761
rect 10167 22731 10209 22761
rect 10243 22731 10285 22761
rect 10319 22761 10321 22765
rect 10355 22765 10391 22795
rect 10425 22765 10461 22795
rect 10495 22765 10530 22795
rect 10564 22765 10599 22795
rect 10633 22765 10668 22795
rect 10355 22761 10361 22765
rect 10425 22761 10437 22765
rect 10495 22761 10513 22765
rect 10564 22761 10589 22765
rect 10633 22761 10665 22765
rect 10702 22761 10737 22795
rect 10793 22794 10806 22795
rect 10866 22794 10875 22795
rect 10939 22794 10944 22795
rect 10771 22761 10806 22794
rect 10840 22761 10875 22794
rect 10909 22761 10944 22794
rect 11012 22795 11051 22828
rect 11085 22795 11124 22828
rect 11158 22795 11197 22828
rect 11231 22795 11270 22828
rect 11304 22795 11343 22828
rect 11377 22795 11416 22828
rect 11450 22795 11489 22828
rect 11523 22795 11562 22828
rect 11596 22795 11635 22828
rect 11669 22795 11707 22828
rect 11741 22795 11779 22828
rect 11813 22795 11851 22828
rect 11885 22795 11923 22828
rect 11957 22795 11995 22828
rect 12029 22795 12067 22828
rect 12101 22795 12139 22828
rect 12173 22795 12211 22828
rect 12245 22795 12451 22828
rect 11012 22794 11013 22795
rect 10978 22761 11013 22794
rect 11047 22794 11051 22795
rect 11116 22794 11124 22795
rect 11185 22794 11197 22795
rect 11254 22794 11270 22795
rect 11323 22794 11343 22795
rect 11392 22794 11416 22795
rect 11461 22794 11489 22795
rect 11530 22794 11562 22795
rect 11047 22761 11082 22794
rect 11116 22761 11151 22794
rect 11185 22761 11220 22794
rect 11254 22761 11289 22794
rect 11323 22761 11358 22794
rect 11392 22761 11427 22794
rect 11461 22761 11496 22794
rect 11530 22761 11565 22794
rect 11599 22761 11634 22795
rect 11669 22794 11703 22795
rect 11741 22794 11772 22795
rect 11813 22794 11841 22795
rect 11885 22794 11910 22795
rect 11957 22794 11979 22795
rect 12029 22794 12048 22795
rect 12101 22794 12117 22795
rect 12173 22794 12186 22795
rect 12245 22794 12255 22795
rect 11668 22761 11703 22794
rect 11737 22761 11772 22794
rect 11806 22761 11841 22794
rect 11875 22761 11910 22794
rect 11944 22761 11979 22794
rect 12013 22761 12048 22794
rect 12082 22761 12117 22794
rect 12151 22761 12186 22794
rect 12220 22761 12255 22794
rect 12289 22761 12324 22795
rect 12358 22761 12393 22795
rect 12427 22761 12451 22795
rect 10319 22731 10361 22761
rect 10395 22731 10437 22761
rect 10471 22731 10513 22761
rect 10547 22731 10589 22761
rect 10623 22731 10665 22761
rect 10699 22742 12451 22761
rect 10699 22731 10759 22742
rect 9877 22725 10759 22731
rect 10793 22725 10832 22742
rect 10866 22725 10905 22742
rect 10939 22725 10978 22742
rect 9877 22691 9901 22725
rect 9935 22691 9971 22725
rect 10005 22691 10041 22725
rect 10075 22691 10111 22725
rect 10145 22691 10181 22725
rect 10215 22691 10251 22725
rect 10285 22691 10321 22725
rect 10355 22691 10391 22725
rect 10425 22691 10461 22725
rect 10495 22691 10530 22725
rect 10564 22691 10599 22725
rect 10633 22691 10668 22725
rect 10702 22691 10737 22725
rect 10793 22708 10806 22725
rect 10866 22708 10875 22725
rect 10939 22708 10944 22725
rect 10771 22691 10806 22708
rect 10840 22691 10875 22708
rect 10909 22691 10944 22708
rect 11012 22725 11051 22742
rect 11085 22725 11124 22742
rect 11158 22725 11197 22742
rect 11231 22725 11270 22742
rect 11304 22725 11343 22742
rect 11377 22725 11416 22742
rect 11450 22725 11489 22742
rect 11523 22725 11562 22742
rect 11596 22725 11635 22742
rect 11669 22725 11707 22742
rect 11741 22725 11779 22742
rect 11813 22725 11851 22742
rect 11885 22725 11923 22742
rect 11957 22725 11995 22742
rect 12029 22725 12067 22742
rect 12101 22725 12139 22742
rect 12173 22725 12211 22742
rect 12245 22725 12451 22742
rect 11012 22708 11013 22725
rect 10978 22691 11013 22708
rect 11047 22708 11051 22725
rect 11116 22708 11124 22725
rect 11185 22708 11197 22725
rect 11254 22708 11270 22725
rect 11323 22708 11343 22725
rect 11392 22708 11416 22725
rect 11461 22708 11489 22725
rect 11530 22708 11562 22725
rect 11047 22691 11082 22708
rect 11116 22691 11151 22708
rect 11185 22691 11220 22708
rect 11254 22691 11289 22708
rect 11323 22691 11358 22708
rect 11392 22691 11427 22708
rect 11461 22691 11496 22708
rect 11530 22691 11565 22708
rect 11599 22691 11634 22725
rect 11669 22708 11703 22725
rect 11741 22708 11772 22725
rect 11813 22708 11841 22725
rect 11885 22708 11910 22725
rect 11957 22708 11979 22725
rect 12029 22708 12048 22725
rect 12101 22708 12117 22725
rect 12173 22708 12186 22725
rect 12245 22708 12255 22725
rect 11668 22691 11703 22708
rect 11737 22691 11772 22708
rect 11806 22691 11841 22708
rect 11875 22691 11910 22708
rect 11944 22691 11979 22708
rect 12013 22691 12048 22708
rect 12082 22691 12117 22708
rect 12151 22691 12186 22708
rect 12220 22691 12255 22708
rect 12289 22691 12324 22725
rect 12358 22691 12393 22725
rect 12427 22691 12451 22725
rect 9877 22657 9905 22691
rect 9939 22657 9981 22691
rect 10015 22657 10057 22691
rect 10091 22657 10133 22691
rect 10167 22657 10209 22691
rect 10243 22657 10285 22691
rect 10319 22657 10361 22691
rect 10395 22657 10437 22691
rect 10471 22657 10513 22691
rect 10547 22657 10589 22691
rect 10623 22657 10665 22691
rect 10699 22657 12451 22691
rect 9877 22656 12451 22657
rect 9877 22655 10759 22656
rect 10793 22655 10832 22656
rect 10866 22655 10905 22656
rect 10939 22655 10978 22656
rect 9877 22621 9901 22655
rect 9935 22621 9971 22655
rect 10005 22621 10041 22655
rect 10075 22621 10111 22655
rect 10145 22621 10181 22655
rect 10215 22621 10251 22655
rect 10285 22621 10321 22655
rect 10355 22621 10391 22655
rect 10425 22621 10461 22655
rect 10495 22621 10530 22655
rect 10564 22621 10599 22655
rect 10633 22621 10668 22655
rect 10702 22621 10737 22655
rect 10793 22622 10806 22655
rect 10866 22622 10875 22655
rect 10939 22622 10944 22655
rect 10771 22621 10806 22622
rect 10840 22621 10875 22622
rect 10909 22621 10944 22622
rect 11012 22655 11051 22656
rect 11085 22655 11124 22656
rect 11158 22655 11197 22656
rect 11231 22655 11270 22656
rect 11304 22655 11343 22656
rect 11377 22655 11416 22656
rect 11450 22655 11489 22656
rect 11523 22655 11562 22656
rect 11596 22655 11635 22656
rect 11669 22655 11707 22656
rect 11741 22655 11779 22656
rect 11813 22655 11851 22656
rect 11885 22655 11923 22656
rect 11957 22655 11995 22656
rect 12029 22655 12067 22656
rect 12101 22655 12139 22656
rect 12173 22655 12211 22656
rect 12245 22655 12451 22656
rect 11012 22622 11013 22655
rect 10978 22621 11013 22622
rect 11047 22622 11051 22655
rect 11116 22622 11124 22655
rect 11185 22622 11197 22655
rect 11254 22622 11270 22655
rect 11323 22622 11343 22655
rect 11392 22622 11416 22655
rect 11461 22622 11489 22655
rect 11530 22622 11562 22655
rect 11047 22621 11082 22622
rect 11116 22621 11151 22622
rect 11185 22621 11220 22622
rect 11254 22621 11289 22622
rect 11323 22621 11358 22622
rect 11392 22621 11427 22622
rect 11461 22621 11496 22622
rect 11530 22621 11565 22622
rect 11599 22621 11634 22655
rect 11669 22622 11703 22655
rect 11741 22622 11772 22655
rect 11813 22622 11841 22655
rect 11885 22622 11910 22655
rect 11957 22622 11979 22655
rect 12029 22622 12048 22655
rect 12101 22622 12117 22655
rect 12173 22622 12186 22655
rect 12245 22622 12255 22655
rect 11668 22621 11703 22622
rect 11737 22621 11772 22622
rect 11806 22621 11841 22622
rect 11875 22621 11910 22622
rect 11944 22621 11979 22622
rect 12013 22621 12048 22622
rect 12082 22621 12117 22622
rect 12151 22621 12186 22622
rect 12220 22621 12255 22622
rect 12289 22621 12324 22655
rect 12358 22621 12393 22655
rect 12427 22621 12451 22655
rect 9877 22617 12451 22621
rect 9877 22585 9905 22617
rect 9939 22585 9981 22617
rect 10015 22585 10057 22617
rect 10091 22585 10133 22617
rect 10167 22585 10209 22617
rect 10243 22585 10285 22617
rect 9877 22551 9901 22585
rect 9939 22583 9971 22585
rect 10015 22583 10041 22585
rect 10091 22583 10111 22585
rect 10167 22583 10181 22585
rect 10243 22583 10251 22585
rect 9935 22551 9971 22583
rect 10005 22551 10041 22583
rect 10075 22551 10111 22583
rect 10145 22551 10181 22583
rect 10215 22551 10251 22583
rect 10319 22585 10361 22617
rect 10395 22585 10437 22617
rect 10471 22585 10513 22617
rect 10547 22585 10589 22617
rect 10623 22585 10665 22617
rect 10699 22585 12451 22617
rect 10319 22583 10321 22585
rect 10285 22551 10321 22583
rect 10355 22583 10361 22585
rect 10425 22583 10437 22585
rect 10495 22583 10513 22585
rect 10564 22583 10589 22585
rect 10633 22583 10665 22585
rect 10355 22551 10391 22583
rect 10425 22551 10461 22583
rect 10495 22551 10530 22583
rect 10564 22551 10599 22583
rect 10633 22551 10668 22583
rect 10702 22551 10737 22585
rect 10771 22551 10806 22585
rect 10840 22551 10875 22585
rect 10909 22551 10944 22585
rect 10978 22551 11013 22585
rect 11047 22551 11082 22585
rect 11116 22551 11151 22585
rect 11185 22551 11220 22585
rect 11254 22551 11289 22585
rect 11323 22551 11358 22585
rect 11392 22551 11427 22585
rect 11461 22551 11496 22585
rect 11530 22551 11565 22585
rect 11599 22551 11634 22585
rect 11668 22551 11703 22585
rect 11737 22551 11772 22585
rect 11806 22551 11841 22585
rect 11875 22551 11910 22585
rect 11944 22551 11979 22585
rect 12013 22551 12048 22585
rect 12082 22551 12117 22585
rect 12151 22551 12186 22585
rect 12220 22551 12255 22585
rect 12289 22551 12324 22585
rect 12358 22551 12393 22585
rect 12427 22551 12451 22585
rect 9877 22549 12451 22551
rect 13600 22925 14233 22927
rect 13600 22891 13756 22925
rect 13790 22903 13828 22925
rect 13862 22903 13900 22925
rect 13934 22903 13972 22925
rect 14006 22903 14044 22925
rect 14078 22903 14116 22925
rect 13790 22891 13796 22903
rect 13862 22891 13864 22903
rect 13600 22869 13796 22891
rect 13830 22869 13864 22891
rect 13898 22891 13900 22903
rect 13966 22891 13972 22903
rect 14034 22891 14044 22903
rect 14102 22891 14116 22903
rect 14150 22908 14233 22925
rect 14267 22908 14301 22942
rect 14335 22908 14369 22942
rect 14403 22908 14429 22942
rect 14150 22905 14429 22908
rect 14150 22891 14252 22905
rect 13898 22869 13932 22891
rect 13966 22869 14000 22891
rect 14034 22869 14068 22891
rect 14102 22873 14252 22891
rect 14286 22873 14324 22905
rect 14358 22873 14429 22905
rect 14102 22869 14233 22873
rect 14286 22871 14301 22873
rect 14358 22871 14369 22873
rect 13600 22851 14233 22869
rect 13600 22817 13756 22851
rect 13790 22833 13828 22851
rect 13862 22833 13900 22851
rect 13934 22833 13972 22851
rect 14006 22833 14044 22851
rect 14078 22833 14116 22851
rect 13790 22817 13796 22833
rect 13862 22817 13864 22833
rect 13600 22799 13796 22817
rect 13830 22799 13864 22817
rect 13898 22817 13900 22833
rect 13966 22817 13972 22833
rect 14034 22817 14044 22833
rect 14102 22817 14116 22833
rect 14150 22839 14233 22851
rect 14267 22839 14301 22871
rect 14335 22839 14369 22871
rect 14403 22839 14429 22873
rect 14150 22832 14429 22839
rect 14150 22817 14252 22832
rect 13898 22799 13932 22817
rect 13966 22799 14000 22817
rect 14034 22799 14068 22817
rect 14102 22804 14252 22817
rect 14286 22804 14324 22832
rect 14358 22804 14429 22832
rect 14102 22799 14233 22804
rect 13600 22777 14233 22799
rect 14286 22798 14301 22804
rect 14358 22798 14369 22804
rect 13600 22743 13756 22777
rect 13790 22763 13828 22777
rect 13862 22763 13900 22777
rect 13934 22763 13972 22777
rect 14006 22763 14044 22777
rect 14078 22763 14116 22777
rect 13790 22743 13796 22763
rect 13862 22743 13864 22763
rect 13600 22729 13796 22743
rect 13830 22729 13864 22743
rect 13898 22743 13900 22763
rect 13966 22743 13972 22763
rect 14034 22743 14044 22763
rect 14102 22743 14116 22763
rect 14150 22770 14233 22777
rect 14267 22770 14301 22798
rect 14335 22770 14369 22798
rect 14403 22770 14429 22804
rect 14150 22759 14429 22770
rect 14150 22743 14252 22759
rect 13898 22729 13932 22743
rect 13966 22729 14000 22743
rect 14034 22729 14068 22743
rect 14102 22735 14252 22743
rect 14286 22735 14324 22759
rect 14358 22735 14429 22759
rect 14102 22729 14233 22735
rect 13600 22703 14233 22729
rect 14286 22725 14301 22735
rect 14358 22725 14369 22735
rect 13600 22669 13756 22703
rect 13790 22693 13828 22703
rect 13862 22693 13900 22703
rect 13934 22693 13972 22703
rect 14006 22693 14044 22703
rect 14078 22693 14116 22703
rect 13790 22669 13796 22693
rect 13862 22669 13864 22693
rect 13600 22659 13796 22669
rect 13830 22659 13864 22669
rect 13898 22669 13900 22693
rect 13966 22669 13972 22693
rect 14034 22669 14044 22693
rect 14102 22669 14116 22693
rect 14150 22701 14233 22703
rect 14267 22701 14301 22725
rect 14335 22701 14369 22725
rect 14403 22701 14429 22735
rect 14150 22686 14429 22701
rect 14150 22669 14252 22686
rect 13898 22659 13932 22669
rect 13966 22659 14000 22669
rect 14034 22659 14068 22669
rect 14102 22666 14252 22669
rect 14286 22666 14324 22686
rect 14358 22666 14429 22686
rect 14102 22659 14233 22666
rect 13600 22632 14233 22659
rect 14286 22652 14301 22666
rect 14358 22652 14369 22666
rect 14267 22632 14301 22652
rect 14335 22632 14369 22652
rect 14403 22632 14429 22666
rect 13600 22629 14429 22632
rect 13600 22595 13756 22629
rect 13790 22623 13828 22629
rect 13862 22623 13900 22629
rect 13934 22623 13972 22629
rect 14006 22623 14044 22629
rect 14078 22623 14116 22629
rect 13790 22595 13796 22623
rect 13862 22595 13864 22623
rect 13600 22589 13796 22595
rect 13830 22589 13864 22595
rect 13898 22595 13900 22623
rect 13966 22595 13972 22623
rect 14034 22595 14044 22623
rect 14102 22595 14116 22623
rect 14150 22613 14429 22629
rect 14150 22597 14252 22613
rect 14286 22597 14324 22613
rect 14358 22597 14429 22613
rect 14150 22595 14233 22597
rect 13898 22589 13932 22595
rect 13966 22589 14000 22595
rect 14034 22589 14068 22595
rect 14102 22589 14233 22595
rect 13600 22563 14233 22589
rect 14286 22579 14301 22597
rect 14358 22579 14369 22597
rect 14267 22563 14301 22579
rect 14335 22563 14369 22579
rect 14403 22563 14429 22597
rect 13600 22555 14429 22563
rect 13600 22521 13756 22555
rect 13790 22553 13828 22555
rect 13862 22553 13900 22555
rect 13934 22553 13972 22555
rect 14006 22553 14044 22555
rect 14078 22553 14116 22555
rect 13790 22521 13796 22553
rect 13862 22521 13864 22553
rect 13600 22519 13796 22521
rect 13830 22519 13864 22521
rect 13898 22521 13900 22553
rect 13966 22521 13972 22553
rect 14034 22521 14044 22553
rect 14102 22521 14116 22553
rect 14150 22540 14429 22555
rect 14150 22528 14252 22540
rect 14286 22528 14324 22540
rect 14358 22528 14429 22540
rect 14150 22521 14233 22528
rect 13898 22519 13932 22521
rect 13966 22519 14000 22521
rect 14034 22519 14068 22521
rect 14102 22519 14233 22521
rect 13600 22494 14233 22519
rect 14286 22506 14301 22528
rect 14358 22506 14369 22528
rect 14267 22494 14301 22506
rect 14335 22494 14369 22506
rect 14403 22494 14429 22528
rect 13600 22483 14429 22494
rect 13600 22481 13796 22483
rect 13830 22481 13864 22483
rect 13600 22447 13756 22481
rect 13790 22449 13796 22481
rect 13862 22449 13864 22481
rect 13898 22481 13932 22483
rect 13966 22481 14000 22483
rect 14034 22481 14068 22483
rect 14102 22481 14429 22483
rect 13898 22449 13900 22481
rect 13966 22449 13972 22481
rect 14034 22449 14044 22481
rect 14102 22449 14116 22481
rect 13790 22447 13828 22449
rect 13862 22447 13900 22449
rect 13934 22447 13972 22449
rect 14006 22447 14044 22449
rect 14078 22447 14116 22449
rect 14150 22467 14429 22481
rect 14150 22459 14252 22467
rect 14286 22459 14324 22467
rect 14358 22459 14429 22467
rect 14150 22447 14233 22459
rect 13600 22425 14233 22447
rect 14286 22433 14301 22459
rect 14358 22433 14369 22459
rect 14267 22425 14301 22433
rect 14335 22425 14369 22433
rect 14403 22425 14429 22459
rect 13600 22413 14429 22425
rect 13600 22407 13796 22413
rect 13830 22407 13864 22413
rect 13600 22373 13756 22407
rect 13790 22379 13796 22407
rect 13862 22379 13864 22407
rect 13898 22407 13932 22413
rect 13966 22407 14000 22413
rect 14034 22407 14068 22413
rect 14102 22407 14429 22413
rect 13898 22379 13900 22407
rect 13966 22379 13972 22407
rect 14034 22379 14044 22407
rect 14102 22379 14116 22407
rect 13790 22373 13828 22379
rect 13862 22373 13900 22379
rect 13934 22373 13972 22379
rect 14006 22373 14044 22379
rect 14078 22373 14116 22379
rect 14150 22394 14429 22407
rect 14150 22390 14252 22394
rect 14286 22390 14324 22394
rect 14358 22390 14429 22394
rect 14150 22373 14233 22390
rect 13600 22356 14233 22373
rect 14286 22360 14301 22390
rect 14358 22360 14369 22390
rect 14267 22356 14301 22360
rect 14335 22356 14369 22360
rect 14403 22356 14429 22390
rect 13600 22343 14429 22356
rect 13600 22333 13796 22343
rect 13830 22333 13864 22343
rect 13600 22299 13756 22333
rect 13790 22309 13796 22333
rect 13862 22309 13864 22333
rect 13898 22333 13932 22343
rect 13966 22333 14000 22343
rect 14034 22333 14068 22343
rect 14102 22333 14429 22343
rect 13898 22309 13900 22333
rect 13966 22309 13972 22333
rect 14034 22309 14044 22333
rect 14102 22309 14116 22333
rect 13790 22299 13828 22309
rect 13862 22299 13900 22309
rect 13934 22299 13972 22309
rect 14006 22299 14044 22309
rect 14078 22299 14116 22309
rect 14150 22321 14429 22333
rect 14150 22299 14233 22321
rect 13600 22287 14233 22299
rect 14286 22287 14301 22321
rect 14358 22287 14369 22321
rect 14403 22287 14429 22321
rect 13600 22273 14429 22287
rect 13600 22259 13796 22273
rect 13830 22259 13864 22273
rect 13600 22225 13756 22259
rect 13790 22239 13796 22259
rect 13862 22239 13864 22259
rect 13898 22259 13932 22273
rect 13966 22259 14000 22273
rect 14034 22259 14068 22273
rect 14102 22259 14429 22273
rect 13898 22239 13900 22259
rect 13966 22239 13972 22259
rect 14034 22239 14044 22259
rect 14102 22239 14116 22259
rect 13790 22225 13828 22239
rect 13862 22225 13900 22239
rect 13934 22225 13972 22239
rect 14006 22225 14044 22239
rect 14078 22225 14116 22239
rect 14150 22252 14429 22259
rect 14150 22225 14233 22252
rect 14267 22248 14301 22252
rect 14335 22248 14369 22252
rect 13600 22218 14233 22225
rect 14286 22218 14301 22248
rect 14358 22218 14369 22248
rect 14403 22218 14429 22252
rect 13600 22214 14252 22218
rect 14286 22214 14324 22218
rect 14358 22214 14429 22218
rect 13600 22203 14429 22214
rect 13600 22185 13796 22203
rect 13830 22185 13864 22203
rect 13600 22151 13756 22185
rect 13790 22169 13796 22185
rect 13862 22169 13864 22185
rect 13898 22185 13932 22203
rect 13966 22185 14000 22203
rect 14034 22185 14068 22203
rect 14102 22185 14429 22203
rect 13898 22169 13900 22185
rect 13966 22169 13972 22185
rect 14034 22169 14044 22185
rect 14102 22169 14116 22185
rect 13790 22151 13828 22169
rect 13862 22151 13900 22169
rect 13934 22151 13972 22169
rect 14006 22151 14044 22169
rect 14078 22151 14116 22169
rect 14150 22183 14429 22185
rect 14150 22151 14233 22183
rect 14267 22175 14301 22183
rect 14335 22175 14369 22183
rect 13600 22149 14233 22151
rect 14286 22149 14301 22175
rect 14358 22149 14369 22175
rect 14403 22149 14429 22183
rect 13600 22141 14252 22149
rect 14286 22141 14324 22149
rect 14358 22141 14429 22149
rect 13600 22133 14429 22141
rect 13600 22111 13796 22133
rect 13830 22111 13864 22133
rect 13600 22077 13756 22111
rect 13790 22099 13796 22111
rect 13862 22099 13864 22111
rect 13898 22111 13932 22133
rect 13966 22111 14000 22133
rect 14034 22111 14068 22133
rect 14102 22114 14429 22133
rect 14102 22111 14233 22114
rect 13898 22099 13900 22111
rect 13966 22099 13972 22111
rect 14034 22099 14044 22111
rect 14102 22099 14116 22111
rect 13790 22077 13828 22099
rect 13862 22077 13900 22099
rect 13934 22077 13972 22099
rect 14006 22077 14044 22099
rect 14078 22077 14116 22099
rect 14150 22080 14233 22111
rect 14267 22102 14301 22114
rect 14335 22102 14369 22114
rect 14286 22080 14301 22102
rect 14358 22080 14369 22102
rect 14403 22080 14429 22114
rect 14150 22077 14252 22080
rect 13600 22068 14252 22077
rect 14286 22068 14324 22080
rect 14358 22068 14429 22080
rect 13600 22063 14429 22068
rect 13600 22037 13796 22063
rect 13830 22037 13864 22063
rect 13600 22032 13756 22037
rect 13750 22003 13756 22032
rect 13790 22029 13796 22037
rect 13862 22029 13864 22037
rect 13898 22037 13932 22063
rect 13966 22037 14000 22063
rect 14034 22037 14068 22063
rect 14102 22045 14429 22063
rect 14102 22037 14233 22045
rect 13898 22029 13900 22037
rect 13966 22029 13972 22037
rect 14034 22029 14044 22037
rect 14102 22029 14116 22037
rect 13790 22003 13828 22029
rect 13862 22003 13900 22029
rect 13934 22003 13972 22029
rect 14006 22003 14044 22029
rect 14078 22003 14116 22029
rect 14150 22011 14233 22037
rect 14267 22029 14301 22045
rect 14335 22029 14369 22045
rect 14286 22011 14301 22029
rect 14358 22011 14369 22029
rect 14403 22011 14429 22045
rect 14150 22003 14252 22011
rect 13750 21995 14252 22003
rect 14286 21995 14324 22011
rect 14358 21995 14429 22011
rect 13750 21993 14429 21995
rect 13750 21963 13796 21993
rect 13830 21963 13864 21993
rect 13750 21929 13756 21963
rect 13790 21959 13796 21963
rect 13862 21959 13864 21963
rect 13898 21963 13932 21993
rect 13966 21963 14000 21993
rect 14034 21963 14068 21993
rect 14102 21976 14429 21993
rect 14102 21963 14233 21976
rect 13898 21959 13900 21963
rect 13966 21959 13972 21963
rect 14034 21959 14044 21963
rect 14102 21959 14116 21963
rect 13790 21929 13828 21959
rect 13862 21929 13900 21959
rect 13934 21929 13972 21959
rect 14006 21929 14044 21959
rect 14078 21929 14116 21959
rect 14150 21942 14233 21963
rect 14267 21956 14301 21976
rect 14335 21956 14369 21976
rect 14286 21942 14301 21956
rect 14358 21942 14369 21956
rect 14403 21942 14429 21976
rect 14150 21929 14252 21942
rect 13750 21923 14252 21929
rect 13750 21889 13796 21923
rect 13830 21889 13864 21923
rect 13898 21889 13932 21923
rect 13966 21889 14000 21923
rect 14034 21889 14068 21923
rect 14102 21922 14252 21923
rect 14286 21922 14324 21942
rect 14358 21922 14429 21942
rect 14102 21907 14429 21922
rect 14102 21889 14233 21907
rect 13750 21855 13756 21889
rect 13790 21855 13828 21889
rect 13862 21855 13900 21889
rect 13934 21855 13972 21889
rect 14006 21855 14044 21889
rect 14078 21855 14116 21889
rect 14150 21873 14233 21889
rect 14267 21883 14301 21907
rect 14335 21883 14369 21907
rect 14286 21873 14301 21883
rect 14358 21873 14369 21883
rect 14403 21873 14429 21907
rect 14150 21855 14252 21873
rect 13750 21853 14252 21855
rect 13750 21819 13796 21853
rect 13830 21819 13864 21853
rect 13898 21819 13932 21853
rect 13966 21819 14000 21853
rect 14034 21819 14068 21853
rect 14102 21849 14252 21853
rect 14286 21849 14324 21873
rect 14358 21849 14429 21873
rect 14102 21838 14429 21849
rect 14102 21819 14233 21838
rect 13750 21815 14233 21819
rect 13750 21781 13756 21815
rect 13790 21783 13828 21815
rect 13862 21783 13900 21815
rect 13934 21783 13972 21815
rect 14006 21783 14044 21815
rect 14078 21783 14116 21815
rect 13790 21781 13796 21783
rect 13862 21781 13864 21783
rect 13750 21749 13796 21781
rect 13830 21749 13864 21781
rect 13898 21781 13900 21783
rect 13966 21781 13972 21783
rect 14034 21781 14044 21783
rect 14102 21781 14116 21783
rect 14150 21804 14233 21815
rect 14267 21810 14301 21838
rect 14335 21810 14369 21838
rect 14286 21804 14301 21810
rect 14358 21804 14369 21810
rect 14403 21804 14429 21838
rect 14150 21781 14252 21804
rect 13898 21749 13932 21781
rect 13966 21749 14000 21781
rect 14034 21749 14068 21781
rect 14102 21776 14252 21781
rect 14286 21776 14324 21804
rect 14358 21776 14429 21804
rect 14102 21769 14429 21776
rect 14102 21749 14233 21769
rect 13750 21741 14233 21749
rect 13750 21707 13756 21741
rect 13790 21713 13828 21741
rect 13862 21713 13900 21741
rect 13934 21713 13972 21741
rect 14006 21713 14044 21741
rect 14078 21713 14116 21741
rect 13790 21707 13796 21713
rect 13862 21707 13864 21713
rect 13750 21679 13796 21707
rect 13830 21679 13864 21707
rect 13898 21707 13900 21713
rect 13966 21707 13972 21713
rect 14034 21707 14044 21713
rect 14102 21707 14116 21713
rect 14150 21735 14233 21741
rect 14267 21737 14301 21769
rect 14335 21737 14369 21769
rect 14286 21735 14301 21737
rect 14358 21735 14369 21737
rect 14403 21735 14429 21769
rect 14150 21707 14252 21735
rect 13898 21679 13932 21707
rect 13966 21679 14000 21707
rect 14034 21679 14068 21707
rect 14102 21703 14252 21707
rect 14286 21703 14324 21735
rect 14358 21703 14429 21735
rect 14102 21700 14429 21703
rect 14102 21679 14233 21700
rect 13750 21666 14233 21679
rect 14267 21666 14301 21700
rect 14335 21666 14369 21700
rect 14403 21666 14429 21700
rect 13750 21632 13756 21666
rect 13790 21643 13828 21666
rect 13862 21643 13900 21666
rect 13934 21643 13972 21666
rect 14006 21643 14044 21666
rect 14078 21643 14116 21666
rect 13790 21632 13796 21643
rect 13862 21632 13864 21643
rect 13750 21609 13796 21632
rect 13830 21609 13864 21632
rect 13898 21632 13900 21643
rect 13966 21632 13972 21643
rect 14034 21632 14044 21643
rect 14102 21632 14116 21643
rect 14150 21664 14429 21666
rect 14150 21632 14252 21664
rect 13898 21609 13932 21632
rect 13966 21609 14000 21632
rect 14034 21609 14068 21632
rect 14102 21631 14252 21632
rect 14286 21631 14324 21664
rect 14358 21631 14429 21664
rect 14102 21609 14233 21631
rect 14286 21630 14301 21631
rect 14358 21630 14369 21631
rect 13750 21597 14233 21609
rect 14267 21597 14301 21630
rect 14335 21597 14369 21630
rect 14403 21597 14429 21631
rect 13750 21591 14429 21597
rect 13750 21557 13756 21591
rect 13790 21573 13828 21591
rect 13862 21573 13900 21591
rect 13934 21573 13972 21591
rect 14006 21573 14044 21591
rect 14078 21573 14116 21591
rect 13790 21557 13796 21573
rect 13862 21557 13864 21573
rect 13750 21539 13796 21557
rect 13830 21539 13864 21557
rect 13898 21557 13900 21573
rect 13966 21557 13972 21573
rect 14034 21557 14044 21573
rect 14102 21557 14116 21573
rect 14150 21562 14252 21591
rect 14286 21562 14324 21591
rect 14358 21562 14429 21591
rect 14150 21557 14233 21562
rect 14286 21557 14301 21562
rect 14358 21557 14369 21562
rect 13898 21539 13932 21557
rect 13966 21539 14000 21557
rect 14034 21539 14068 21557
rect 14102 21539 14233 21557
rect 13750 21528 14233 21539
rect 14267 21528 14301 21557
rect 14335 21528 14369 21557
rect 14403 21528 14429 21562
rect 13750 21518 14429 21528
rect 13750 21516 14252 21518
rect 13750 21482 13756 21516
rect 13790 21503 13828 21516
rect 13862 21503 13900 21516
rect 13934 21503 13972 21516
rect 14006 21503 14044 21516
rect 14078 21503 14116 21516
rect 13790 21482 13796 21503
rect 13862 21482 13864 21503
rect 13750 21469 13796 21482
rect 13830 21469 13864 21482
rect 13898 21482 13900 21503
rect 13966 21482 13972 21503
rect 14034 21482 14044 21503
rect 14102 21482 14116 21503
rect 14150 21493 14252 21516
rect 14286 21493 14324 21518
rect 14358 21493 14429 21518
rect 14150 21482 14233 21493
rect 14286 21484 14301 21493
rect 14358 21484 14369 21493
rect 13898 21469 13932 21482
rect 13966 21469 14000 21482
rect 14034 21469 14068 21482
rect 14102 21469 14233 21482
rect 13750 21459 14233 21469
rect 14267 21459 14301 21484
rect 14335 21459 14369 21484
rect 14403 21459 14429 21493
rect 13750 21445 14429 21459
rect 13750 21441 14252 21445
rect 13750 21407 13756 21441
rect 13790 21433 13828 21441
rect 13862 21433 13900 21441
rect 13934 21433 13972 21441
rect 14006 21433 14044 21441
rect 14078 21433 14116 21441
rect 13790 21407 13796 21433
rect 13862 21407 13864 21433
rect 13750 21399 13796 21407
rect 13830 21399 13864 21407
rect 13898 21407 13900 21433
rect 13966 21407 13972 21433
rect 14034 21407 14044 21433
rect 14102 21407 14116 21433
rect 14150 21424 14252 21441
rect 14286 21424 14324 21445
rect 14358 21424 14429 21445
rect 14150 21407 14233 21424
rect 14286 21411 14301 21424
rect 14358 21411 14369 21424
rect 13898 21399 13932 21407
rect 13966 21399 14000 21407
rect 14034 21399 14068 21407
rect 14102 21399 14233 21407
rect 13750 21390 14233 21399
rect 14267 21390 14301 21411
rect 14335 21390 14369 21411
rect 14403 21390 14429 21424
rect 13750 21371 14429 21390
rect 13750 21366 14252 21371
rect 13750 21332 13756 21366
rect 13790 21363 13828 21366
rect 13862 21363 13900 21366
rect 13934 21363 13972 21366
rect 14006 21363 14044 21366
rect 14078 21363 14116 21366
rect 13790 21332 13796 21363
rect 13862 21332 13864 21363
rect 13750 21329 13796 21332
rect 13830 21329 13864 21332
rect 13898 21332 13900 21363
rect 13966 21332 13972 21363
rect 14034 21332 14044 21363
rect 14102 21332 14116 21363
rect 14150 21355 14252 21366
rect 14286 21355 14324 21371
rect 14358 21355 14429 21371
rect 14150 21332 14233 21355
rect 14286 21337 14301 21355
rect 14358 21337 14369 21355
rect 13898 21329 13932 21332
rect 13966 21329 14000 21332
rect 14034 21329 14068 21332
rect 14102 21329 14233 21332
rect 13750 21321 14233 21329
rect 14267 21321 14301 21337
rect 14335 21321 14369 21337
rect 14403 21321 14429 21355
rect 13750 21297 14429 21321
rect 13750 21293 14252 21297
rect 13750 21291 13796 21293
rect 13830 21291 13864 21293
rect 13750 21257 13756 21291
rect 13790 21259 13796 21291
rect 13862 21259 13864 21291
rect 13898 21291 13932 21293
rect 13966 21291 14000 21293
rect 14034 21291 14068 21293
rect 14102 21291 14252 21293
rect 13898 21259 13900 21291
rect 13966 21259 13972 21291
rect 14034 21259 14044 21291
rect 14102 21259 14116 21291
rect 13790 21257 13828 21259
rect 13862 21257 13900 21259
rect 13934 21257 13972 21259
rect 14006 21257 14044 21259
rect 14078 21257 14116 21259
rect 14150 21286 14252 21291
rect 14286 21286 14324 21297
rect 14358 21286 14429 21297
rect 14150 21257 14233 21286
rect 14286 21263 14301 21286
rect 14358 21263 14369 21286
rect 13750 21252 14233 21257
rect 14267 21252 14301 21263
rect 14335 21252 14369 21263
rect 14403 21252 14429 21286
rect 13750 21223 14429 21252
rect 13750 21216 13796 21223
rect 13830 21216 13864 21223
rect 13750 21182 13756 21216
rect 13790 21189 13796 21216
rect 13862 21189 13864 21216
rect 13898 21216 13932 21223
rect 13966 21216 14000 21223
rect 14034 21216 14068 21223
rect 14102 21217 14252 21223
rect 14286 21217 14324 21223
rect 14358 21217 14429 21223
rect 14102 21216 14233 21217
rect 13898 21189 13900 21216
rect 13966 21189 13972 21216
rect 14034 21189 14044 21216
rect 14102 21189 14116 21216
rect 13790 21182 13828 21189
rect 13862 21182 13900 21189
rect 13934 21182 13972 21189
rect 14006 21182 14044 21189
rect 14078 21182 14116 21189
rect 14150 21183 14233 21216
rect 14286 21189 14301 21217
rect 14358 21189 14369 21217
rect 14267 21183 14301 21189
rect 14335 21183 14369 21189
rect 14403 21183 14429 21217
rect 14150 21182 14429 21183
rect 13750 21153 14429 21182
rect 13750 21141 13796 21153
rect 13830 21141 13864 21153
rect 13750 21107 13756 21141
rect 13790 21119 13796 21141
rect 13862 21119 13864 21141
rect 13898 21141 13932 21153
rect 13966 21141 14000 21153
rect 14034 21141 14068 21153
rect 14102 21149 14429 21153
rect 14102 21148 14252 21149
rect 14286 21148 14324 21149
rect 14358 21148 14429 21149
rect 14102 21141 14233 21148
rect 13898 21119 13900 21141
rect 13966 21119 13972 21141
rect 14034 21119 14044 21141
rect 14102 21119 14116 21141
rect 13790 21107 13828 21119
rect 13862 21107 13900 21119
rect 13934 21107 13972 21119
rect 14006 21107 14044 21119
rect 14078 21107 14116 21119
rect 14150 21114 14233 21141
rect 14286 21115 14301 21148
rect 14358 21115 14369 21148
rect 14267 21114 14301 21115
rect 14335 21114 14369 21115
rect 14403 21114 14429 21148
rect 14150 21107 14429 21114
rect 13750 21083 14429 21107
rect 13750 21066 13796 21083
rect 13830 21066 13864 21083
rect 13750 21032 13756 21066
rect 13790 21049 13796 21066
rect 13862 21049 13864 21066
rect 13898 21066 13932 21083
rect 13966 21066 14000 21083
rect 14034 21066 14068 21083
rect 14102 21079 14429 21083
rect 14102 21066 14233 21079
rect 14267 21075 14301 21079
rect 14335 21075 14369 21079
rect 13898 21049 13900 21066
rect 13966 21049 13972 21066
rect 14034 21049 14044 21066
rect 14102 21049 14116 21066
rect 13790 21032 13828 21049
rect 13862 21032 13900 21049
rect 13934 21032 13972 21049
rect 14006 21032 14044 21049
rect 14078 21032 14116 21049
rect 14150 21045 14233 21066
rect 14286 21045 14301 21075
rect 14358 21045 14369 21075
rect 14403 21045 14429 21079
rect 14150 21041 14252 21045
rect 14286 21041 14324 21045
rect 14358 21041 14429 21045
rect 14150 21032 14429 21041
rect 13750 21012 14429 21032
rect 13750 20978 13796 21012
rect 13830 20978 13864 21012
rect 13898 20978 13932 21012
rect 13966 20978 14000 21012
rect 14034 20978 14068 21012
rect 14102 21010 14429 21012
rect 14102 20978 14233 21010
rect 13750 20976 14233 20978
rect 14267 20976 14301 21010
rect 14335 20976 14369 21010
rect 14403 20976 14429 21010
rect 13750 20941 14429 20976
rect 13750 20907 13796 20941
rect 13830 20907 13864 20941
rect 13898 20907 13932 20941
rect 13966 20907 14000 20941
rect 14034 20907 14068 20941
rect 14102 20907 14233 20941
rect 14267 20907 14301 20941
rect 14335 20907 14369 20941
rect 14403 20907 14429 20941
rect 13750 20874 14429 20907
rect 10911 17287 10945 17325
rect 1807 10943 1841 10981
rect 1807 10871 1841 10909
rect 1807 10799 1841 10837
rect 1923 10943 1957 10981
rect 1923 10871 1957 10909
rect 1923 10799 1957 10837
rect 517 10594 567 10628
rect 517 10182 567 10216
rect 846 5383 1592 5414
rect 880 5349 926 5383
rect 960 5349 1005 5383
rect 1039 5349 1084 5383
rect 1118 5349 1163 5383
rect 1197 5349 1242 5383
rect 1276 5349 1321 5383
rect 1355 5349 1400 5383
rect 1434 5349 1479 5383
rect 1513 5349 1558 5383
rect 846 5318 1592 5349
rect 517 3700 567 3734
rect 517 3288 567 3322
rect 951 3233 985 3271
rect 517 3178 567 3212
rect 1807 3260 1841 3298
rect 1807 3188 1841 3226
rect 1807 3116 1841 3154
rect 1923 3260 1957 3298
rect 1923 3188 1957 3226
rect 1923 3116 1957 3154
rect 11365 1486 11437 1492
rect 11399 1458 11437 1486
rect 11471 1458 11509 1492
rect 11543 1458 11581 1492
rect 11615 1458 11653 1492
rect 11687 1458 11725 1492
rect 11759 1458 11797 1492
rect 11831 1458 11869 1492
rect 11903 1458 11941 1492
rect 11975 1458 12013 1492
rect 12047 1458 12085 1492
rect 12119 1458 12157 1492
rect 12191 1458 12229 1492
rect 12263 1458 12301 1492
rect 12335 1458 12373 1492
rect 12407 1458 12445 1492
rect 12479 1458 12517 1492
rect 12551 1458 12589 1492
rect 12623 1458 12661 1492
rect 12695 1458 12733 1492
rect 12767 1458 12805 1492
rect 12839 1458 12877 1492
rect 12911 1458 12949 1492
rect 12983 1458 13021 1492
rect 13055 1458 13093 1492
rect 13127 1458 13165 1492
rect 13199 1458 13237 1492
rect 13271 1458 13309 1492
rect 13343 1486 13415 1492
rect 13343 1458 13381 1486
rect 11365 1406 11399 1434
rect 13381 1406 13415 1434
rect 11365 1325 11399 1359
rect 11365 1244 11399 1284
rect 12243 1226 12277 1376
rect 12503 1226 12537 1376
rect 13381 1325 13415 1359
rect 13381 1244 13415 1284
rect 11365 1168 11399 1209
rect 11365 1092 11399 1129
rect 11481 1154 11515 1192
rect 11481 1082 11515 1120
rect 11737 1154 11771 1192
rect 11737 1082 11771 1120
rect 11861 1154 11895 1192
rect 11861 1082 11895 1120
rect 12117 1154 12151 1192
rect 12243 1154 12277 1192
rect 12373 1154 12407 1192
rect 12503 1154 12537 1192
rect 12629 1154 12663 1192
rect 12117 1082 12151 1120
rect 12373 1082 12407 1120
rect 12629 1082 12663 1120
rect 12885 1154 12919 1192
rect 12885 1082 12919 1120
rect 13009 1154 13043 1192
rect 13009 1082 13043 1120
rect 13265 1154 13299 1192
rect 13265 1082 13299 1120
rect 13381 1168 13415 1209
rect 13381 1092 13415 1129
rect 11365 1034 11399 1048
rect 13381 1034 13415 1048
rect 11365 814 11399 822
rect 13381 814 13415 822
rect 11365 719 11399 764
rect 11365 630 11399 680
rect 11481 742 11515 780
rect 11481 670 11515 708
rect 11737 742 11771 780
rect 11737 670 11771 708
rect 11993 742 12027 780
rect 11993 670 12027 708
rect 12753 742 12787 780
rect 12127 624 12165 658
rect 12199 624 12237 658
rect 12753 670 12787 708
rect 11365 546 11399 590
rect 12369 594 12403 644
rect 12543 624 12581 658
rect 12615 624 12653 658
rect 13009 742 13043 780
rect 13009 670 13043 708
rect 13265 742 13299 780
rect 13265 670 13299 708
rect 13381 719 13415 764
rect 13381 630 13415 680
rect 13381 546 13415 590
rect 11399 494 11437 522
rect 11365 488 11437 494
rect 11471 488 11509 522
rect 11543 488 11581 522
rect 11615 488 11653 522
rect 11687 488 11725 522
rect 11759 488 11797 522
rect 11831 488 11869 522
rect 11903 488 11941 522
rect 11975 488 12013 522
rect 12047 488 12085 522
rect 12119 488 12157 522
rect 12191 488 12229 522
rect 12263 488 12301 522
rect 12335 488 12373 522
rect 12407 488 12445 522
rect 12479 488 12517 522
rect 12551 488 12589 522
rect 12623 488 12661 522
rect 12695 488 12733 522
rect 12767 488 12805 522
rect 12839 488 12877 522
rect 12911 488 12949 522
rect 12983 488 13021 522
rect 13055 488 13093 522
rect 13127 488 13165 522
rect 13199 488 13237 522
rect 13271 488 13309 522
rect 13343 494 13381 522
rect 13343 488 13415 494
<< viali >>
rect 9915 36349 9949 36351
rect 9987 36349 10021 36351
rect 10059 36349 10093 36351
rect 10131 36349 10165 36351
rect 10203 36349 10237 36351
rect 10275 36349 10309 36351
rect 10347 36349 10381 36351
rect 10419 36349 10453 36351
rect 10491 36349 10525 36351
rect 10563 36349 10597 36351
rect 10635 36349 10669 36351
rect 10707 36349 10741 36351
rect 10779 36349 10813 36351
rect 10851 36349 10885 36351
rect 9915 36317 9949 36349
rect 9987 36317 10021 36349
rect 10059 36317 10093 36349
rect 10131 36317 10165 36349
rect 10203 36317 10237 36349
rect 10275 36317 10309 36349
rect 10347 36317 10381 36349
rect 10419 36317 10453 36349
rect 10491 36317 10525 36349
rect 10563 36317 10597 36349
rect 10635 36317 10669 36349
rect 10707 36317 10741 36349
rect 10779 36317 10813 36349
rect 10851 36317 10884 36349
rect 10884 36317 10885 36349
rect 10927 36348 10961 36379
rect 11000 36348 11034 36379
rect 11073 36348 11107 36379
rect 11146 36348 11180 36379
rect 11219 36348 11253 36379
rect 11292 36348 11326 36379
rect 11365 36348 11399 36379
rect 11438 36348 11472 36379
rect 11511 36348 11545 36379
rect 11584 36348 11618 36379
rect 11657 36348 11691 36379
rect 11730 36348 11764 36379
rect 11803 36348 11837 36379
rect 11876 36348 11910 36379
rect 11949 36348 11983 36379
rect 12022 36348 12056 36379
rect 12095 36348 12129 36379
rect 12168 36348 12202 36379
rect 12241 36348 12275 36379
rect 12314 36348 12348 36379
rect 12387 36348 12421 36379
rect 12460 36348 12494 36379
rect 12533 36348 12567 36379
rect 12606 36348 12640 36379
rect 12679 36348 12713 36379
rect 12752 36348 12786 36379
rect 12825 36348 12859 36379
rect 12898 36348 12932 36379
rect 12971 36348 13005 36379
rect 13044 36348 13078 36379
rect 13117 36348 13151 36379
rect 13190 36348 13224 36379
rect 13263 36348 13297 36379
rect 13336 36348 13370 36379
rect 13409 36348 13443 36379
rect 13482 36348 13516 36379
rect 13555 36348 13589 36379
rect 13628 36348 13662 36379
rect 13701 36348 13735 36379
rect 13774 36348 13808 36379
rect 13846 36348 13880 36379
rect 13918 36348 13952 36379
rect 13990 36348 14024 36379
rect 14062 36348 14096 36379
rect 14134 36348 14168 36379
rect 14206 36348 14240 36379
rect 14278 36348 14312 36379
rect 14350 36348 14384 36379
rect 10927 36345 10939 36348
rect 10939 36345 10961 36348
rect 11000 36345 11008 36348
rect 11008 36345 11034 36348
rect 11073 36345 11077 36348
rect 11077 36345 11107 36348
rect 11146 36345 11180 36348
rect 11219 36345 11249 36348
rect 11249 36345 11253 36348
rect 11292 36345 11318 36348
rect 11318 36345 11326 36348
rect 11365 36345 11387 36348
rect 11387 36345 11399 36348
rect 11438 36345 11456 36348
rect 11456 36345 11472 36348
rect 11511 36345 11525 36348
rect 11525 36345 11545 36348
rect 11584 36345 11594 36348
rect 11594 36345 11618 36348
rect 11657 36345 11663 36348
rect 11663 36345 11691 36348
rect 11730 36345 11732 36348
rect 11732 36345 11764 36348
rect 11803 36345 11836 36348
rect 11836 36345 11837 36348
rect 11876 36345 11905 36348
rect 11905 36345 11910 36348
rect 11949 36345 11974 36348
rect 11974 36345 11983 36348
rect 12022 36345 12043 36348
rect 12043 36345 12056 36348
rect 12095 36345 12112 36348
rect 12112 36345 12129 36348
rect 12168 36345 12181 36348
rect 12181 36345 12202 36348
rect 12241 36345 12250 36348
rect 12250 36345 12275 36348
rect 12314 36345 12319 36348
rect 12319 36345 12348 36348
rect 12387 36345 12388 36348
rect 12388 36345 12421 36348
rect 12460 36345 12494 36348
rect 12533 36345 12567 36348
rect 12606 36345 12640 36348
rect 12679 36345 12713 36348
rect 12752 36345 12786 36348
rect 12825 36345 12859 36348
rect 12898 36345 12932 36348
rect 12971 36345 13005 36348
rect 13044 36345 13078 36348
rect 13117 36345 13151 36348
rect 13190 36345 13224 36348
rect 13263 36345 13297 36348
rect 13336 36345 13370 36348
rect 13409 36345 13443 36348
rect 13482 36345 13516 36348
rect 13555 36345 13589 36348
rect 13628 36345 13662 36348
rect 13701 36345 13735 36348
rect 13774 36345 13808 36348
rect 13846 36345 13880 36348
rect 13918 36345 13952 36348
rect 13990 36345 14024 36348
rect 14062 36345 14096 36348
rect 14134 36345 14168 36348
rect 14206 36345 14240 36348
rect 14278 36345 14312 36348
rect 14350 36345 14384 36348
rect 10927 36280 10961 36303
rect 11000 36280 11034 36303
rect 11073 36280 11107 36303
rect 11146 36280 11180 36303
rect 11219 36280 11253 36303
rect 11292 36280 11326 36303
rect 11365 36280 11399 36303
rect 11438 36280 11472 36303
rect 11511 36280 11545 36303
rect 11584 36280 11618 36303
rect 11657 36280 11691 36303
rect 11730 36280 11764 36303
rect 11803 36280 11837 36303
rect 11876 36280 11910 36303
rect 11949 36280 11983 36303
rect 12022 36280 12056 36303
rect 12095 36280 12129 36303
rect 12168 36280 12202 36303
rect 12241 36280 12275 36303
rect 12314 36280 12348 36303
rect 12387 36280 12421 36303
rect 9915 36239 9949 36273
rect 9987 36239 10021 36273
rect 10059 36239 10093 36273
rect 10131 36239 10165 36273
rect 10203 36239 10237 36273
rect 10275 36239 10309 36273
rect 10347 36239 10381 36273
rect 10419 36239 10453 36273
rect 10491 36239 10525 36273
rect 10563 36239 10597 36273
rect 10635 36239 10669 36273
rect 10707 36239 10741 36273
rect 10779 36239 10813 36273
rect 10851 36239 10884 36273
rect 10884 36239 10885 36273
rect 10927 36269 10939 36280
rect 10939 36269 10961 36280
rect 11000 36269 11008 36280
rect 11008 36269 11034 36280
rect 11073 36269 11077 36280
rect 11077 36269 11107 36280
rect 11146 36269 11180 36280
rect 11219 36269 11249 36280
rect 11249 36269 11253 36280
rect 11292 36269 11318 36280
rect 11318 36269 11326 36280
rect 11365 36269 11387 36280
rect 11387 36269 11399 36280
rect 11438 36269 11456 36280
rect 11456 36269 11472 36280
rect 11511 36269 11525 36280
rect 11525 36269 11545 36280
rect 11584 36269 11594 36280
rect 11594 36269 11618 36280
rect 11657 36269 11663 36280
rect 11663 36269 11691 36280
rect 11730 36269 11732 36280
rect 11732 36269 11764 36280
rect 11803 36269 11836 36280
rect 11836 36269 11837 36280
rect 11876 36269 11905 36280
rect 11905 36269 11910 36280
rect 11949 36269 11974 36280
rect 11974 36269 11983 36280
rect 12022 36269 12043 36280
rect 12043 36269 12056 36280
rect 12095 36269 12112 36280
rect 12112 36269 12129 36280
rect 12168 36269 12181 36280
rect 12181 36269 12202 36280
rect 12241 36269 12250 36280
rect 12250 36269 12275 36280
rect 12314 36269 12319 36280
rect 12319 36269 12348 36280
rect 12387 36269 12388 36280
rect 12388 36269 12421 36280
rect 12460 36269 12494 36303
rect 12533 36269 12567 36303
rect 12606 36269 12640 36303
rect 12679 36269 12713 36303
rect 12752 36269 12786 36303
rect 12825 36269 12859 36303
rect 12898 36269 12932 36303
rect 12971 36269 13005 36303
rect 13044 36269 13078 36303
rect 13117 36269 13151 36303
rect 13190 36269 13224 36303
rect 13263 36269 13297 36303
rect 13336 36269 13370 36303
rect 13409 36269 13443 36303
rect 13482 36269 13516 36303
rect 13555 36269 13589 36303
rect 13628 36269 13662 36303
rect 13701 36269 13735 36303
rect 13774 36269 13808 36303
rect 13846 36269 13880 36303
rect 13918 36269 13952 36303
rect 13990 36269 14024 36303
rect 14062 36269 14096 36303
rect 14134 36269 14168 36303
rect 14206 36269 14240 36303
rect 14278 36269 14312 36303
rect 14350 36269 14384 36303
rect 10927 36212 10961 36227
rect 11000 36212 11034 36227
rect 11073 36212 11107 36227
rect 11146 36212 11180 36227
rect 11219 36212 11253 36227
rect 11292 36212 11326 36227
rect 11365 36212 11399 36227
rect 11438 36212 11472 36227
rect 11511 36212 11545 36227
rect 11584 36212 11618 36227
rect 11657 36212 11691 36227
rect 11730 36212 11764 36227
rect 11803 36212 11837 36227
rect 11876 36212 11910 36227
rect 11949 36212 11983 36227
rect 12022 36212 12056 36227
rect 12095 36212 12129 36227
rect 12168 36212 12202 36227
rect 12241 36212 12275 36227
rect 12314 36212 12348 36227
rect 12387 36212 12421 36227
rect 9915 36161 9949 36195
rect 9987 36161 10021 36195
rect 10059 36161 10093 36195
rect 10131 36161 10165 36195
rect 10203 36161 10237 36195
rect 10275 36161 10309 36195
rect 10347 36161 10381 36195
rect 10419 36161 10453 36195
rect 10491 36161 10525 36195
rect 10563 36161 10597 36195
rect 10635 36161 10669 36195
rect 10707 36161 10741 36195
rect 10779 36161 10813 36195
rect 10851 36161 10884 36195
rect 10884 36161 10885 36195
rect 10927 36193 10939 36212
rect 10939 36193 10961 36212
rect 11000 36193 11008 36212
rect 11008 36193 11034 36212
rect 11073 36193 11077 36212
rect 11077 36193 11107 36212
rect 11146 36193 11180 36212
rect 11219 36193 11249 36212
rect 11249 36193 11253 36212
rect 11292 36193 11318 36212
rect 11318 36193 11326 36212
rect 11365 36193 11387 36212
rect 11387 36193 11399 36212
rect 11438 36193 11456 36212
rect 11456 36193 11472 36212
rect 11511 36193 11525 36212
rect 11525 36193 11545 36212
rect 11584 36193 11594 36212
rect 11594 36193 11618 36212
rect 11657 36193 11663 36212
rect 11663 36193 11691 36212
rect 11730 36193 11732 36212
rect 11732 36193 11764 36212
rect 11803 36193 11836 36212
rect 11836 36193 11837 36212
rect 11876 36193 11905 36212
rect 11905 36193 11910 36212
rect 11949 36193 11974 36212
rect 11974 36193 11983 36212
rect 12022 36193 12043 36212
rect 12043 36193 12056 36212
rect 12095 36193 12112 36212
rect 12112 36193 12129 36212
rect 12168 36193 12181 36212
rect 12181 36193 12202 36212
rect 12241 36193 12250 36212
rect 12250 36193 12275 36212
rect 12314 36193 12319 36212
rect 12319 36193 12348 36212
rect 12387 36193 12388 36212
rect 12388 36193 12421 36212
rect 12460 36193 12494 36227
rect 12533 36193 12567 36227
rect 12606 36193 12640 36227
rect 12679 36193 12713 36227
rect 12752 36193 12786 36227
rect 12825 36193 12859 36227
rect 12898 36193 12932 36227
rect 12971 36193 13005 36227
rect 13044 36193 13078 36227
rect 13117 36193 13151 36227
rect 13190 36193 13224 36227
rect 13263 36193 13297 36227
rect 13336 36193 13370 36227
rect 13409 36193 13443 36227
rect 13482 36193 13516 36227
rect 13555 36193 13589 36227
rect 13628 36193 13662 36227
rect 13701 36193 13735 36227
rect 13774 36193 13808 36227
rect 13846 36193 13880 36227
rect 13918 36193 13952 36227
rect 13990 36193 14024 36227
rect 14062 36193 14096 36227
rect 14134 36193 14168 36227
rect 14206 36193 14240 36227
rect 14278 36193 14312 36227
rect 14350 36193 14384 36227
rect 10927 36144 10961 36151
rect 11000 36144 11034 36151
rect 11073 36144 11107 36151
rect 11146 36144 11180 36151
rect 11219 36144 11253 36151
rect 11292 36144 11326 36151
rect 11365 36144 11399 36151
rect 11438 36144 11472 36151
rect 11511 36144 11545 36151
rect 11584 36144 11618 36151
rect 11657 36144 11691 36151
rect 11730 36144 11764 36151
rect 11803 36144 11837 36151
rect 11876 36144 11910 36151
rect 11949 36144 11983 36151
rect 12022 36144 12056 36151
rect 12095 36144 12129 36151
rect 12168 36144 12202 36151
rect 12241 36144 12275 36151
rect 12314 36144 12348 36151
rect 12387 36144 12421 36151
rect 10927 36117 10939 36144
rect 10939 36117 10961 36144
rect 11000 36117 11008 36144
rect 11008 36117 11034 36144
rect 11073 36117 11077 36144
rect 11077 36117 11107 36144
rect 9915 36082 9949 36116
rect 9987 36082 10021 36116
rect 10059 36082 10093 36116
rect 10131 36082 10165 36116
rect 10203 36082 10237 36116
rect 10275 36082 10309 36116
rect 10347 36082 10381 36116
rect 10419 36082 10453 36116
rect 10491 36082 10525 36116
rect 10563 36082 10597 36116
rect 10635 36082 10669 36116
rect 10707 36082 10741 36116
rect 10779 36082 10813 36116
rect 10851 36082 10884 36116
rect 10884 36082 10885 36116
rect 11146 36117 11180 36144
rect 11219 36117 11249 36144
rect 11249 36117 11253 36144
rect 11292 36117 11318 36144
rect 11318 36117 11326 36144
rect 11365 36117 11387 36144
rect 11387 36117 11399 36144
rect 11438 36117 11456 36144
rect 11456 36117 11472 36144
rect 11511 36117 11525 36144
rect 11525 36117 11545 36144
rect 11584 36117 11594 36144
rect 11594 36117 11618 36144
rect 11657 36117 11663 36144
rect 11663 36117 11691 36144
rect 11730 36117 11732 36144
rect 11732 36117 11764 36144
rect 11803 36117 11836 36144
rect 11836 36117 11837 36144
rect 11876 36117 11905 36144
rect 11905 36117 11910 36144
rect 11949 36117 11974 36144
rect 11974 36117 11983 36144
rect 12022 36117 12043 36144
rect 12043 36117 12056 36144
rect 12095 36117 12112 36144
rect 12112 36117 12129 36144
rect 12168 36117 12181 36144
rect 12181 36117 12202 36144
rect 12241 36117 12250 36144
rect 12250 36117 12275 36144
rect 12314 36117 12319 36144
rect 12319 36117 12348 36144
rect 12387 36117 12388 36144
rect 12388 36117 12421 36144
rect 12460 36117 12494 36151
rect 12533 36117 12567 36151
rect 12606 36117 12640 36151
rect 12679 36117 12713 36151
rect 12752 36117 12786 36151
rect 12825 36117 12859 36151
rect 12898 36117 12932 36151
rect 12971 36117 13005 36151
rect 13044 36117 13078 36151
rect 13117 36117 13151 36151
rect 13190 36117 13224 36151
rect 13263 36117 13297 36151
rect 13336 36117 13370 36151
rect 13409 36117 13443 36151
rect 13482 36117 13516 36151
rect 13555 36117 13589 36151
rect 13628 36117 13662 36151
rect 13701 36117 13735 36151
rect 13774 36117 13808 36151
rect 13846 36117 13880 36151
rect 13918 36117 13952 36151
rect 13990 36117 14024 36151
rect 14062 36117 14096 36151
rect 14134 36117 14168 36151
rect 14206 36117 14240 36151
rect 14278 36117 14312 36151
rect 14350 36117 14384 36151
rect 10927 36042 10939 36075
rect 10939 36042 10961 36075
rect 11000 36042 11008 36075
rect 11008 36042 11034 36075
rect 11073 36042 11077 36075
rect 11077 36042 11107 36075
rect 11146 36042 11180 36075
rect 11219 36042 11249 36075
rect 11249 36042 11253 36075
rect 11292 36042 11318 36075
rect 11318 36042 11326 36075
rect 11365 36042 11387 36075
rect 11387 36042 11399 36075
rect 11438 36042 11456 36075
rect 11456 36042 11472 36075
rect 11511 36042 11525 36075
rect 11525 36042 11545 36075
rect 11584 36042 11594 36075
rect 11594 36042 11618 36075
rect 11657 36042 11663 36075
rect 11663 36042 11691 36075
rect 11730 36042 11732 36075
rect 11732 36042 11764 36075
rect 11803 36042 11836 36075
rect 11836 36042 11837 36075
rect 11876 36042 11905 36075
rect 11905 36042 11910 36075
rect 11949 36042 11974 36075
rect 11974 36042 11983 36075
rect 12022 36042 12043 36075
rect 12043 36042 12056 36075
rect 12095 36042 12112 36075
rect 12112 36042 12129 36075
rect 12168 36042 12181 36075
rect 12181 36042 12202 36075
rect 12241 36042 12250 36075
rect 12250 36042 12275 36075
rect 12314 36042 12319 36075
rect 12319 36042 12348 36075
rect 12387 36042 12388 36075
rect 12388 36042 12421 36075
rect 10927 36041 10961 36042
rect 11000 36041 11034 36042
rect 11073 36041 11107 36042
rect 11146 36041 11180 36042
rect 11219 36041 11253 36042
rect 11292 36041 11326 36042
rect 11365 36041 11399 36042
rect 11438 36041 11472 36042
rect 11511 36041 11545 36042
rect 11584 36041 11618 36042
rect 11657 36041 11691 36042
rect 11730 36041 11764 36042
rect 11803 36041 11837 36042
rect 11876 36041 11910 36042
rect 11949 36041 11983 36042
rect 12022 36041 12056 36042
rect 12095 36041 12129 36042
rect 12168 36041 12202 36042
rect 12241 36041 12275 36042
rect 12314 36041 12348 36042
rect 12387 36041 12421 36042
rect 12460 36041 12494 36075
rect 12533 36041 12567 36075
rect 12606 36041 12640 36075
rect 12679 36041 12713 36075
rect 12752 36041 12786 36075
rect 12825 36041 12859 36075
rect 12898 36041 12932 36075
rect 12971 36041 13005 36075
rect 13044 36041 13078 36075
rect 13117 36041 13151 36075
rect 13190 36041 13224 36075
rect 13263 36041 13297 36075
rect 13336 36041 13370 36075
rect 13409 36041 13443 36075
rect 13482 36041 13516 36075
rect 13555 36041 13589 36075
rect 13628 36041 13662 36075
rect 13701 36041 13735 36075
rect 13774 36041 13808 36075
rect 13846 36041 13880 36075
rect 13918 36041 13952 36075
rect 13990 36041 14024 36075
rect 14062 36041 14096 36075
rect 14134 36041 14168 36075
rect 14206 36041 14240 36075
rect 14278 36041 14312 36075
rect 14350 36041 14384 36075
rect 9915 36003 9949 36037
rect 9987 36003 10021 36037
rect 10059 36003 10093 36037
rect 10131 36003 10165 36037
rect 10203 36003 10237 36037
rect 10275 36003 10309 36037
rect 10347 36003 10381 36037
rect 10419 36003 10453 36037
rect 10491 36003 10525 36037
rect 10563 36003 10597 36037
rect 10635 36003 10669 36037
rect 10707 36003 10741 36037
rect 10779 36003 10813 36037
rect 10851 36003 10884 36037
rect 10884 36003 10885 36037
rect 10927 35974 10939 35999
rect 10939 35974 10961 35999
rect 11000 35974 11008 35999
rect 11008 35974 11034 35999
rect 11073 35974 11077 35999
rect 11077 35974 11107 35999
rect 11146 35974 11180 35999
rect 11219 35974 11249 35999
rect 11249 35974 11253 35999
rect 11292 35974 11318 35999
rect 11318 35974 11326 35999
rect 11365 35974 11387 35999
rect 11387 35974 11399 35999
rect 11438 35974 11456 35999
rect 11456 35974 11472 35999
rect 11511 35974 11525 35999
rect 11525 35974 11545 35999
rect 11584 35974 11594 35999
rect 11594 35974 11618 35999
rect 11657 35974 11663 35999
rect 11663 35974 11691 35999
rect 11730 35974 11732 35999
rect 11732 35974 11764 35999
rect 11803 35974 11836 35999
rect 11836 35974 11837 35999
rect 11876 35974 11905 35999
rect 11905 35974 11910 35999
rect 11949 35974 11974 35999
rect 11974 35974 11983 35999
rect 12022 35974 12043 35999
rect 12043 35974 12056 35999
rect 12095 35974 12112 35999
rect 12112 35974 12129 35999
rect 12168 35974 12181 35999
rect 12181 35974 12202 35999
rect 12241 35974 12250 35999
rect 12250 35974 12275 35999
rect 12314 35974 12319 35999
rect 12319 35974 12348 35999
rect 12387 35974 12388 35999
rect 12388 35974 12421 35999
rect 10927 35965 10961 35974
rect 11000 35965 11034 35974
rect 11073 35965 11107 35974
rect 11146 35965 11180 35974
rect 11219 35965 11253 35974
rect 11292 35965 11326 35974
rect 11365 35965 11399 35974
rect 11438 35965 11472 35974
rect 11511 35965 11545 35974
rect 11584 35965 11618 35974
rect 11657 35965 11691 35974
rect 11730 35965 11764 35974
rect 11803 35965 11837 35974
rect 11876 35965 11910 35974
rect 11949 35965 11983 35974
rect 12022 35965 12056 35974
rect 12095 35965 12129 35974
rect 12168 35965 12202 35974
rect 12241 35965 12275 35974
rect 12314 35965 12348 35974
rect 12387 35965 12421 35974
rect 12460 35965 12494 35999
rect 12533 35965 12567 35999
rect 12606 35965 12640 35999
rect 12679 35965 12713 35999
rect 12752 35965 12786 35999
rect 12825 35965 12859 35999
rect 12898 35965 12932 35999
rect 12971 35965 13005 35999
rect 13044 35965 13078 35999
rect 13117 35965 13151 35999
rect 13190 35965 13224 35999
rect 13263 35965 13297 35999
rect 13336 35965 13370 35999
rect 13409 35965 13443 35999
rect 13482 35965 13516 35999
rect 13555 35965 13589 35999
rect 13628 35965 13662 35999
rect 13701 35965 13735 35999
rect 13774 35965 13808 35999
rect 13846 35965 13880 35999
rect 13918 35965 13952 35999
rect 13990 35965 14024 35999
rect 14062 35965 14096 35999
rect 14134 35965 14168 35999
rect 14206 35965 14240 35999
rect 14278 35965 14312 35999
rect 14350 35965 14384 35999
rect 9915 35940 9949 35958
rect 9987 35940 10021 35958
rect 10059 35940 10093 35958
rect 10131 35940 10165 35958
rect 10203 35940 10237 35958
rect 10275 35940 10309 35958
rect 10347 35940 10381 35958
rect 10419 35940 10453 35958
rect 10491 35940 10525 35958
rect 10563 35940 10597 35958
rect 10635 35940 10669 35958
rect 10707 35940 10741 35958
rect 10779 35940 10813 35958
rect 10851 35940 10885 35958
rect 9915 35924 9932 35940
rect 9932 35924 9949 35940
rect 9987 35924 10000 35940
rect 10000 35924 10021 35940
rect 10059 35924 10068 35940
rect 10068 35924 10093 35940
rect 10131 35924 10136 35940
rect 10136 35924 10165 35940
rect 10203 35924 10204 35940
rect 10204 35924 10237 35940
rect 10275 35924 10306 35940
rect 10306 35924 10309 35940
rect 10347 35924 10374 35940
rect 10374 35924 10381 35940
rect 10419 35924 10442 35940
rect 10442 35924 10453 35940
rect 10491 35924 10510 35940
rect 10510 35924 10525 35940
rect 10563 35924 10578 35940
rect 10578 35924 10597 35940
rect 10635 35924 10646 35940
rect 10646 35924 10669 35940
rect 10707 35924 10714 35940
rect 10714 35924 10741 35940
rect 10779 35924 10782 35940
rect 10782 35924 10813 35940
rect 10851 35924 10884 35940
rect 10884 35924 10885 35940
rect 10927 35906 10939 35923
rect 10939 35906 10961 35923
rect 11000 35906 11008 35923
rect 11008 35906 11034 35923
rect 11073 35906 11077 35923
rect 11077 35906 11107 35923
rect 11146 35906 11180 35923
rect 11219 35906 11249 35923
rect 11249 35906 11253 35923
rect 11292 35906 11318 35923
rect 11318 35906 11326 35923
rect 11365 35906 11387 35923
rect 11387 35906 11399 35923
rect 11438 35906 11456 35923
rect 11456 35906 11472 35923
rect 11511 35906 11525 35923
rect 11525 35906 11545 35923
rect 11584 35906 11594 35923
rect 11594 35906 11618 35923
rect 11657 35906 11663 35923
rect 11663 35906 11691 35923
rect 11730 35906 11732 35923
rect 11732 35906 11764 35923
rect 11803 35906 11836 35923
rect 11836 35906 11837 35923
rect 11876 35906 11905 35923
rect 11905 35906 11910 35923
rect 11949 35906 11974 35923
rect 11974 35906 11983 35923
rect 12022 35906 12043 35923
rect 12043 35906 12056 35923
rect 12095 35906 12112 35923
rect 12112 35906 12129 35923
rect 12168 35906 12181 35923
rect 12181 35906 12202 35923
rect 12241 35906 12250 35923
rect 12250 35906 12275 35923
rect 12314 35906 12319 35923
rect 12319 35906 12348 35923
rect 12387 35906 12388 35923
rect 12388 35906 12421 35923
rect 10927 35889 10961 35906
rect 11000 35889 11034 35906
rect 11073 35889 11107 35906
rect 11146 35889 11180 35906
rect 11219 35889 11253 35906
rect 11292 35889 11326 35906
rect 11365 35889 11399 35906
rect 11438 35889 11472 35906
rect 11511 35889 11545 35906
rect 11584 35889 11618 35906
rect 11657 35889 11691 35906
rect 11730 35889 11764 35906
rect 11803 35889 11837 35906
rect 11876 35889 11910 35906
rect 11949 35889 11983 35906
rect 12022 35889 12056 35906
rect 12095 35889 12129 35906
rect 12168 35889 12202 35906
rect 12241 35889 12275 35906
rect 12314 35889 12348 35906
rect 12387 35889 12421 35906
rect 12460 35889 12494 35923
rect 12533 35889 12567 35923
rect 12606 35889 12640 35923
rect 12679 35889 12713 35923
rect 12752 35889 12786 35923
rect 12825 35889 12859 35923
rect 12898 35889 12932 35923
rect 12971 35889 13005 35923
rect 13044 35889 13078 35923
rect 13117 35889 13151 35923
rect 13190 35889 13224 35923
rect 13263 35889 13297 35923
rect 13336 35889 13370 35923
rect 13409 35889 13443 35923
rect 13482 35889 13516 35923
rect 13555 35889 13589 35923
rect 13628 35889 13662 35923
rect 13701 35889 13735 35923
rect 13774 35889 13808 35923
rect 13846 35889 13880 35923
rect 13918 35889 13952 35923
rect 13990 35889 14024 35923
rect 14062 35889 14096 35923
rect 14134 35889 14168 35923
rect 14206 35889 14240 35923
rect 14278 35889 14312 35923
rect 14350 35889 14384 35923
rect 9915 35871 9949 35879
rect 9987 35871 10021 35879
rect 10059 35871 10093 35879
rect 10131 35871 10165 35879
rect 10203 35871 10237 35879
rect 10275 35871 10309 35879
rect 10347 35871 10381 35879
rect 10419 35871 10453 35879
rect 10491 35871 10525 35879
rect 10563 35871 10597 35879
rect 10635 35871 10669 35879
rect 10707 35871 10741 35879
rect 10779 35871 10813 35879
rect 10851 35871 10885 35879
rect 9915 35845 9932 35871
rect 9932 35845 9949 35871
rect 9987 35845 10000 35871
rect 10000 35845 10021 35871
rect 10059 35845 10068 35871
rect 10068 35845 10093 35871
rect 10131 35845 10136 35871
rect 10136 35845 10165 35871
rect 10203 35845 10204 35871
rect 10204 35845 10237 35871
rect 10275 35845 10306 35871
rect 10306 35845 10309 35871
rect 10347 35845 10374 35871
rect 10374 35845 10381 35871
rect 10419 35845 10442 35871
rect 10442 35845 10453 35871
rect 10491 35845 10510 35871
rect 10510 35845 10525 35871
rect 10563 35845 10578 35871
rect 10578 35845 10597 35871
rect 10635 35845 10646 35871
rect 10646 35845 10669 35871
rect 10707 35845 10714 35871
rect 10714 35845 10741 35871
rect 10779 35845 10782 35871
rect 10782 35845 10813 35871
rect 10851 35845 10884 35871
rect 10884 35845 10885 35871
rect 10927 35838 10939 35847
rect 10939 35838 10961 35847
rect 11000 35838 11008 35847
rect 11008 35838 11034 35847
rect 11073 35838 11077 35847
rect 11077 35838 11107 35847
rect 11146 35838 11180 35847
rect 11219 35838 11249 35847
rect 11249 35838 11253 35847
rect 11292 35838 11318 35847
rect 11318 35838 11326 35847
rect 11365 35838 11387 35847
rect 11387 35838 11399 35847
rect 11438 35838 11456 35847
rect 11456 35838 11472 35847
rect 11511 35838 11525 35847
rect 11525 35838 11545 35847
rect 11584 35838 11594 35847
rect 11594 35838 11618 35847
rect 11657 35838 11663 35847
rect 11663 35838 11691 35847
rect 11730 35838 11732 35847
rect 11732 35838 11764 35847
rect 11803 35838 11836 35847
rect 11836 35838 11837 35847
rect 11876 35838 11905 35847
rect 11905 35838 11910 35847
rect 11949 35838 11974 35847
rect 11974 35838 11983 35847
rect 12022 35838 12043 35847
rect 12043 35838 12056 35847
rect 12095 35838 12112 35847
rect 12112 35838 12129 35847
rect 12168 35838 12181 35847
rect 12181 35838 12202 35847
rect 12241 35838 12250 35847
rect 12250 35838 12275 35847
rect 12314 35838 12319 35847
rect 12319 35838 12348 35847
rect 12387 35838 12388 35847
rect 12388 35838 12421 35847
rect 10927 35813 10961 35838
rect 11000 35813 11034 35838
rect 11073 35813 11107 35838
rect 11146 35813 11180 35838
rect 11219 35813 11253 35838
rect 11292 35813 11326 35838
rect 11365 35813 11399 35838
rect 11438 35813 11472 35838
rect 11511 35813 11545 35838
rect 11584 35813 11618 35838
rect 11657 35813 11691 35838
rect 11730 35813 11764 35838
rect 11803 35813 11837 35838
rect 11876 35813 11910 35838
rect 11949 35813 11983 35838
rect 12022 35813 12056 35838
rect 12095 35813 12129 35838
rect 12168 35813 12202 35838
rect 12241 35813 12275 35838
rect 12314 35813 12348 35838
rect 12387 35813 12421 35838
rect 12460 35813 12494 35847
rect 12533 35813 12567 35847
rect 12606 35813 12640 35847
rect 12679 35813 12713 35847
rect 12752 35813 12786 35847
rect 12825 35813 12859 35847
rect 12898 35813 12932 35847
rect 12971 35813 13005 35847
rect 13044 35813 13078 35847
rect 13117 35813 13151 35847
rect 13190 35813 13224 35847
rect 13263 35813 13297 35847
rect 13336 35813 13370 35847
rect 13409 35813 13443 35847
rect 13482 35813 13516 35847
rect 13555 35813 13589 35847
rect 13628 35813 13662 35847
rect 13701 35813 13735 35847
rect 13774 35813 13808 35847
rect 13846 35813 13880 35847
rect 13918 35813 13952 35847
rect 13990 35813 14024 35847
rect 14062 35813 14096 35847
rect 14134 35813 14168 35847
rect 14206 35813 14240 35847
rect 14278 35813 14312 35847
rect 14350 35813 14384 35847
rect 9915 35768 9932 35800
rect 9932 35768 9949 35800
rect 9987 35768 10000 35800
rect 10000 35768 10021 35800
rect 10059 35768 10068 35800
rect 10068 35768 10093 35800
rect 10131 35768 10136 35800
rect 10136 35768 10165 35800
rect 10203 35768 10204 35800
rect 10204 35768 10237 35800
rect 10275 35768 10306 35800
rect 10306 35768 10309 35800
rect 10347 35768 10374 35800
rect 10374 35768 10381 35800
rect 10419 35768 10442 35800
rect 10442 35768 10453 35800
rect 10491 35768 10510 35800
rect 10510 35768 10525 35800
rect 10563 35768 10578 35800
rect 10578 35768 10597 35800
rect 10635 35768 10646 35800
rect 10646 35768 10669 35800
rect 10707 35768 10714 35800
rect 10714 35768 10741 35800
rect 10779 35768 10782 35800
rect 10782 35768 10813 35800
rect 10851 35768 10884 35800
rect 10884 35768 10885 35800
rect 9915 35766 9949 35768
rect 9987 35766 10021 35768
rect 10059 35766 10093 35768
rect 10131 35766 10165 35768
rect 10203 35766 10237 35768
rect 10275 35766 10309 35768
rect 10347 35766 10381 35768
rect 10419 35766 10453 35768
rect 10491 35766 10525 35768
rect 10563 35766 10597 35768
rect 10635 35766 10669 35768
rect 10707 35766 10741 35768
rect 10779 35766 10813 35768
rect 10851 35766 10885 35768
rect 10927 35770 10939 35771
rect 10939 35770 10961 35771
rect 11000 35770 11008 35771
rect 11008 35770 11034 35771
rect 11073 35770 11077 35771
rect 11077 35770 11107 35771
rect 11146 35770 11180 35771
rect 11219 35770 11249 35771
rect 11249 35770 11253 35771
rect 11292 35770 11318 35771
rect 11318 35770 11326 35771
rect 11365 35770 11387 35771
rect 11387 35770 11399 35771
rect 11438 35770 11456 35771
rect 11456 35770 11472 35771
rect 11511 35770 11525 35771
rect 11525 35770 11545 35771
rect 11584 35770 11594 35771
rect 11594 35770 11618 35771
rect 11657 35770 11663 35771
rect 11663 35770 11691 35771
rect 11730 35770 11732 35771
rect 11732 35770 11764 35771
rect 11803 35770 11836 35771
rect 11836 35770 11837 35771
rect 11876 35770 11905 35771
rect 11905 35770 11910 35771
rect 11949 35770 11974 35771
rect 11974 35770 11983 35771
rect 12022 35770 12043 35771
rect 12043 35770 12056 35771
rect 12095 35770 12112 35771
rect 12112 35770 12129 35771
rect 12168 35770 12181 35771
rect 12181 35770 12202 35771
rect 12241 35770 12250 35771
rect 12250 35770 12275 35771
rect 12314 35770 12319 35771
rect 12319 35770 12348 35771
rect 12387 35770 12388 35771
rect 12388 35770 12421 35771
rect 12460 35770 12494 35771
rect 12533 35770 12567 35771
rect 12606 35770 12640 35771
rect 12679 35770 12713 35771
rect 12752 35770 12786 35771
rect 12825 35770 12859 35771
rect 12898 35770 12932 35771
rect 12971 35770 13005 35771
rect 13044 35770 13078 35771
rect 13117 35770 13151 35771
rect 13190 35770 13224 35771
rect 13263 35770 13297 35771
rect 13336 35770 13370 35771
rect 13409 35770 13443 35771
rect 13482 35770 13516 35771
rect 13555 35770 13589 35771
rect 13628 35770 13662 35771
rect 13701 35770 13735 35771
rect 13774 35770 13808 35771
rect 13846 35770 13880 35771
rect 13918 35770 13952 35771
rect 13990 35770 14024 35771
rect 14062 35770 14096 35771
rect 14134 35770 14168 35771
rect 14206 35770 14240 35771
rect 14278 35770 14312 35771
rect 14350 35770 14384 35771
rect 10927 35737 10961 35770
rect 11000 35737 11034 35770
rect 11073 35737 11107 35770
rect 11146 35737 11180 35770
rect 11219 35737 11253 35770
rect 11292 35737 11326 35770
rect 11365 35737 11399 35770
rect 11438 35737 11472 35770
rect 11511 35737 11545 35770
rect 11584 35737 11618 35770
rect 11657 35737 11691 35770
rect 11730 35737 11764 35770
rect 11803 35737 11837 35770
rect 11876 35737 11910 35770
rect 11949 35737 11983 35770
rect 12022 35737 12056 35770
rect 12095 35737 12129 35770
rect 12168 35737 12202 35770
rect 12241 35737 12275 35770
rect 12314 35737 12348 35770
rect 12387 35737 12421 35770
rect 12460 35737 12494 35770
rect 12533 35737 12567 35770
rect 12606 35737 12640 35770
rect 12679 35737 12713 35770
rect 12752 35737 12786 35770
rect 12825 35737 12859 35770
rect 12898 35737 12932 35770
rect 12971 35737 13005 35770
rect 13044 35737 13078 35770
rect 13117 35737 13151 35770
rect 13190 35737 13224 35770
rect 13263 35737 13297 35770
rect 13336 35737 13370 35770
rect 13409 35737 13443 35770
rect 13482 35737 13516 35770
rect 13555 35737 13589 35770
rect 13628 35737 13662 35770
rect 13701 35737 13735 35770
rect 13774 35737 13808 35770
rect 13846 35737 13880 35770
rect 13918 35737 13952 35770
rect 13990 35737 14024 35770
rect 14062 35737 14096 35770
rect 14134 35737 14168 35770
rect 14206 35737 14240 35770
rect 14278 35737 14312 35770
rect 14350 35737 14384 35770
rect 13216 35663 13250 35697
rect 13289 35663 13323 35697
rect 13362 35663 13396 35697
rect 13435 35663 13469 35697
rect 13508 35663 13542 35697
rect 13581 35663 13615 35697
rect 13654 35663 13688 35697
rect 13727 35663 13761 35697
rect 13800 35663 13834 35697
rect 13873 35663 13907 35697
rect 13946 35663 13980 35697
rect 14019 35663 14053 35697
rect 14092 35663 14126 35697
rect 14165 35663 14199 35697
rect 14238 35663 14272 35697
rect 14311 35663 14345 35697
rect 14384 35663 14392 35697
rect 14392 35663 14418 35697
rect 13216 35599 13250 35625
rect 13289 35599 13323 35625
rect 13362 35599 13396 35625
rect 13435 35599 13469 35625
rect 13508 35599 13542 35625
rect 13581 35599 13615 35625
rect 13654 35599 13688 35625
rect 13727 35599 13761 35625
rect 13800 35599 13834 35625
rect 13873 35599 13907 35625
rect 13946 35599 13980 35625
rect 14019 35599 14053 35625
rect 14092 35599 14126 35625
rect 14165 35599 14199 35625
rect 14238 35599 14272 35625
rect 14311 35599 14345 35625
rect 14384 35599 14392 35625
rect 14392 35599 14418 35625
rect 13216 35591 13250 35599
rect 13289 35591 13323 35599
rect 13362 35591 13396 35599
rect 13435 35591 13469 35599
rect 13508 35591 13542 35599
rect 13581 35591 13615 35599
rect 13654 35591 13688 35599
rect 13727 35591 13761 35599
rect 13800 35591 13834 35599
rect 13873 35591 13907 35599
rect 13946 35591 13980 35599
rect 14019 35591 14053 35599
rect 14092 35591 14126 35599
rect 14165 35591 14199 35599
rect 14238 35591 14272 35599
rect 14311 35591 14345 35599
rect 14384 35591 14418 35599
rect 13216 35530 13236 35553
rect 13236 35530 13250 35553
rect 13289 35530 13304 35553
rect 13304 35530 13323 35553
rect 13362 35530 13372 35553
rect 13372 35530 13396 35553
rect 13435 35530 13440 35553
rect 13440 35530 13469 35553
rect 13216 35519 13250 35530
rect 13289 35519 13323 35530
rect 13362 35519 13396 35530
rect 13435 35519 13469 35530
rect 13508 35519 13542 35553
rect 13581 35530 13610 35553
rect 13610 35530 13615 35553
rect 13654 35530 13678 35553
rect 13678 35530 13688 35553
rect 13727 35530 13746 35553
rect 13746 35530 13761 35553
rect 13800 35530 13814 35553
rect 13814 35530 13834 35553
rect 13873 35530 13882 35553
rect 13882 35530 13907 35553
rect 13946 35530 13950 35553
rect 13950 35530 13980 35553
rect 14019 35530 14052 35553
rect 14052 35530 14053 35553
rect 14092 35530 14120 35553
rect 14120 35530 14126 35553
rect 14165 35530 14188 35553
rect 14188 35530 14199 35553
rect 14238 35530 14256 35553
rect 14256 35530 14272 35553
rect 14311 35530 14324 35553
rect 14324 35530 14345 35553
rect 14384 35530 14392 35553
rect 14392 35530 14418 35553
rect 13581 35519 13615 35530
rect 13654 35519 13688 35530
rect 13727 35519 13761 35530
rect 13800 35519 13834 35530
rect 13873 35519 13907 35530
rect 13946 35519 13980 35530
rect 14019 35519 14053 35530
rect 14092 35519 14126 35530
rect 14165 35519 14199 35530
rect 14238 35519 14272 35530
rect 14311 35519 14345 35530
rect 14384 35519 14418 35530
rect 13216 35461 13236 35481
rect 13236 35461 13250 35481
rect 13289 35461 13304 35481
rect 13304 35461 13323 35481
rect 13362 35461 13372 35481
rect 13372 35461 13396 35481
rect 13435 35461 13440 35481
rect 13440 35461 13469 35481
rect 13216 35447 13250 35461
rect 13289 35447 13323 35461
rect 13362 35447 13396 35461
rect 13435 35447 13469 35461
rect 13508 35447 13542 35481
rect 13581 35461 13610 35481
rect 13610 35461 13615 35481
rect 13654 35461 13678 35481
rect 13678 35461 13688 35481
rect 13727 35461 13746 35481
rect 13746 35461 13761 35481
rect 13800 35461 13814 35481
rect 13814 35461 13834 35481
rect 13873 35461 13882 35481
rect 13882 35461 13907 35481
rect 13946 35461 13950 35481
rect 13950 35461 13980 35481
rect 14019 35461 14052 35481
rect 14052 35461 14053 35481
rect 14092 35461 14120 35481
rect 14120 35461 14126 35481
rect 14165 35461 14188 35481
rect 14188 35461 14199 35481
rect 14238 35461 14256 35481
rect 14256 35461 14272 35481
rect 14311 35461 14324 35481
rect 14324 35461 14345 35481
rect 14384 35461 14392 35481
rect 14392 35461 14418 35481
rect 13581 35447 13615 35461
rect 13654 35447 13688 35461
rect 13727 35447 13761 35461
rect 13800 35447 13834 35461
rect 13873 35447 13907 35461
rect 13946 35447 13980 35461
rect 14019 35447 14053 35461
rect 14092 35447 14126 35461
rect 14165 35447 14199 35461
rect 14238 35447 14272 35461
rect 14311 35447 14345 35461
rect 14384 35447 14418 35461
rect 13216 35392 13236 35409
rect 13236 35392 13250 35409
rect 13289 35392 13304 35409
rect 13304 35392 13323 35409
rect 13362 35392 13372 35409
rect 13372 35392 13396 35409
rect 13435 35392 13440 35409
rect 13440 35392 13469 35409
rect 13216 35375 13250 35392
rect 13289 35375 13323 35392
rect 13362 35375 13396 35392
rect 13435 35375 13469 35392
rect 13508 35375 13542 35409
rect 13581 35392 13610 35409
rect 13610 35392 13615 35409
rect 13654 35392 13678 35409
rect 13678 35392 13688 35409
rect 13727 35392 13746 35409
rect 13746 35392 13761 35409
rect 13800 35392 13814 35409
rect 13814 35392 13834 35409
rect 13873 35392 13882 35409
rect 13882 35392 13907 35409
rect 13946 35392 13950 35409
rect 13950 35392 13980 35409
rect 14019 35392 14052 35409
rect 14052 35392 14053 35409
rect 14092 35392 14120 35409
rect 14120 35392 14126 35409
rect 14165 35392 14188 35409
rect 14188 35392 14199 35409
rect 14238 35392 14256 35409
rect 14256 35392 14272 35409
rect 14311 35392 14324 35409
rect 14324 35392 14345 35409
rect 14384 35392 14392 35409
rect 14392 35392 14418 35409
rect 13581 35375 13615 35392
rect 13654 35375 13688 35392
rect 13727 35375 13761 35392
rect 13800 35375 13834 35392
rect 13873 35375 13907 35392
rect 13946 35375 13980 35392
rect 14019 35375 14053 35392
rect 14092 35375 14126 35392
rect 14165 35375 14199 35392
rect 14238 35375 14272 35392
rect 14311 35375 14345 35392
rect 14384 35375 14418 35392
rect 13216 35323 13236 35337
rect 13236 35323 13250 35337
rect 13289 35323 13304 35337
rect 13304 35323 13323 35337
rect 13362 35323 13372 35337
rect 13372 35323 13396 35337
rect 13435 35323 13440 35337
rect 13440 35323 13469 35337
rect 13216 35303 13250 35323
rect 13289 35303 13323 35323
rect 13362 35303 13396 35323
rect 13435 35303 13469 35323
rect 13508 35303 13542 35337
rect 13581 35323 13610 35337
rect 13610 35323 13615 35337
rect 13654 35323 13678 35337
rect 13678 35323 13688 35337
rect 13727 35323 13746 35337
rect 13746 35323 13761 35337
rect 13800 35323 13814 35337
rect 13814 35323 13834 35337
rect 13873 35323 13882 35337
rect 13882 35323 13907 35337
rect 13946 35323 13950 35337
rect 13950 35323 13980 35337
rect 14019 35323 14052 35337
rect 14052 35323 14053 35337
rect 14092 35323 14120 35337
rect 14120 35323 14126 35337
rect 14165 35323 14188 35337
rect 14188 35323 14199 35337
rect 14238 35323 14256 35337
rect 14256 35323 14272 35337
rect 14311 35323 14324 35337
rect 14324 35323 14345 35337
rect 14384 35323 14392 35337
rect 14392 35323 14418 35337
rect 13581 35303 13615 35323
rect 13654 35303 13688 35323
rect 13727 35303 13761 35323
rect 13800 35303 13834 35323
rect 13873 35303 13907 35323
rect 13946 35303 13980 35323
rect 14019 35303 14053 35323
rect 14092 35303 14126 35323
rect 14165 35303 14199 35323
rect 14238 35303 14272 35323
rect 14311 35303 14345 35323
rect 14384 35303 14418 35323
rect 13216 35254 13236 35265
rect 13236 35254 13250 35265
rect 13289 35254 13304 35265
rect 13304 35254 13323 35265
rect 13362 35254 13372 35265
rect 13372 35254 13396 35265
rect 13435 35254 13440 35265
rect 13440 35254 13469 35265
rect 13216 35231 13250 35254
rect 13289 35231 13323 35254
rect 13362 35231 13396 35254
rect 13435 35231 13469 35254
rect 13508 35231 13542 35265
rect 13581 35254 13610 35265
rect 13610 35254 13615 35265
rect 13654 35254 13678 35265
rect 13678 35254 13688 35265
rect 13727 35254 13746 35265
rect 13746 35254 13761 35265
rect 13800 35254 13814 35265
rect 13814 35254 13834 35265
rect 13873 35254 13882 35265
rect 13882 35254 13907 35265
rect 13946 35254 13950 35265
rect 13950 35254 13980 35265
rect 14019 35254 14052 35265
rect 14052 35254 14053 35265
rect 14092 35254 14120 35265
rect 14120 35254 14126 35265
rect 14165 35254 14188 35265
rect 14188 35254 14199 35265
rect 14238 35254 14256 35265
rect 14256 35254 14272 35265
rect 14311 35254 14324 35265
rect 14324 35254 14345 35265
rect 14384 35254 14392 35265
rect 14392 35254 14418 35265
rect 13581 35231 13615 35254
rect 13654 35231 13688 35254
rect 13727 35231 13761 35254
rect 13800 35231 13834 35254
rect 13873 35231 13907 35254
rect 13946 35231 13980 35254
rect 14019 35231 14053 35254
rect 14092 35231 14126 35254
rect 14165 35231 14199 35254
rect 14238 35231 14272 35254
rect 14311 35231 14345 35254
rect 14384 35231 14418 35254
rect 13216 35185 13236 35193
rect 13236 35185 13250 35193
rect 13289 35185 13304 35193
rect 13304 35185 13323 35193
rect 13362 35185 13372 35193
rect 13372 35185 13396 35193
rect 13435 35185 13440 35193
rect 13440 35185 13469 35193
rect 13216 35159 13250 35185
rect 13289 35159 13323 35185
rect 13362 35159 13396 35185
rect 13435 35159 13469 35185
rect 13508 35159 13542 35193
rect 13581 35185 13610 35193
rect 13610 35185 13615 35193
rect 13654 35185 13678 35193
rect 13678 35185 13688 35193
rect 13727 35185 13746 35193
rect 13746 35185 13761 35193
rect 13800 35185 13814 35193
rect 13814 35185 13834 35193
rect 13873 35185 13882 35193
rect 13882 35185 13907 35193
rect 13946 35185 13950 35193
rect 13950 35185 13980 35193
rect 14019 35185 14052 35193
rect 14052 35185 14053 35193
rect 14092 35185 14120 35193
rect 14120 35185 14126 35193
rect 14165 35185 14188 35193
rect 14188 35185 14199 35193
rect 14238 35185 14256 35193
rect 14256 35185 14272 35193
rect 14311 35185 14324 35193
rect 14324 35185 14345 35193
rect 14384 35185 14392 35193
rect 14392 35185 14418 35193
rect 13581 35159 13615 35185
rect 13654 35159 13688 35185
rect 13727 35159 13761 35185
rect 13800 35159 13834 35185
rect 13873 35159 13907 35185
rect 13946 35159 13980 35185
rect 14019 35159 14053 35185
rect 14092 35159 14126 35185
rect 14165 35159 14199 35185
rect 14238 35159 14272 35185
rect 14311 35159 14345 35185
rect 14384 35159 14418 35185
rect 13216 35116 13236 35121
rect 13236 35116 13250 35121
rect 13289 35116 13304 35121
rect 13304 35116 13323 35121
rect 13362 35116 13372 35121
rect 13372 35116 13396 35121
rect 13435 35116 13440 35121
rect 13440 35116 13469 35121
rect 13216 35087 13250 35116
rect 13289 35087 13323 35116
rect 13362 35087 13396 35116
rect 13435 35087 13469 35116
rect 13508 35087 13542 35121
rect 13581 35116 13610 35121
rect 13610 35116 13615 35121
rect 13654 35116 13678 35121
rect 13678 35116 13688 35121
rect 13727 35116 13746 35121
rect 13746 35116 13761 35121
rect 13800 35116 13814 35121
rect 13814 35116 13834 35121
rect 13873 35116 13882 35121
rect 13882 35116 13907 35121
rect 13946 35116 13950 35121
rect 13950 35116 13980 35121
rect 14019 35116 14052 35121
rect 14052 35116 14053 35121
rect 14092 35116 14120 35121
rect 14120 35116 14126 35121
rect 14165 35116 14188 35121
rect 14188 35116 14199 35121
rect 14238 35116 14256 35121
rect 14256 35116 14272 35121
rect 14311 35116 14324 35121
rect 14324 35116 14345 35121
rect 14384 35116 14392 35121
rect 14392 35116 14418 35121
rect 13581 35087 13615 35116
rect 13654 35087 13688 35116
rect 13727 35087 13761 35116
rect 13800 35087 13834 35116
rect 13873 35087 13907 35116
rect 13946 35087 13980 35116
rect 14019 35087 14053 35116
rect 14092 35087 14126 35116
rect 14165 35087 14199 35116
rect 14238 35087 14272 35116
rect 14311 35087 14345 35116
rect 14384 35087 14418 35116
rect 13216 35047 13236 35049
rect 13236 35047 13250 35049
rect 13289 35047 13304 35049
rect 13304 35047 13323 35049
rect 13362 35047 13372 35049
rect 13372 35047 13396 35049
rect 13435 35047 13440 35049
rect 13440 35047 13469 35049
rect 13216 35015 13250 35047
rect 13289 35015 13323 35047
rect 13362 35015 13396 35047
rect 13435 35015 13469 35047
rect 13508 35015 13542 35049
rect 13581 35047 13610 35049
rect 13610 35047 13615 35049
rect 13654 35047 13678 35049
rect 13678 35047 13688 35049
rect 13727 35047 13746 35049
rect 13746 35047 13761 35049
rect 13800 35047 13814 35049
rect 13814 35047 13834 35049
rect 13873 35047 13882 35049
rect 13882 35047 13907 35049
rect 13946 35047 13950 35049
rect 13950 35047 13980 35049
rect 14019 35047 14052 35049
rect 14052 35047 14053 35049
rect 14092 35047 14120 35049
rect 14120 35047 14126 35049
rect 14165 35047 14188 35049
rect 14188 35047 14199 35049
rect 14238 35047 14256 35049
rect 14256 35047 14272 35049
rect 14311 35047 14324 35049
rect 14324 35047 14345 35049
rect 14384 35047 14392 35049
rect 14392 35047 14418 35049
rect 13581 35015 13615 35047
rect 13654 35015 13688 35047
rect 13727 35015 13761 35047
rect 13800 35015 13834 35047
rect 13873 35015 13907 35047
rect 13946 35015 13980 35047
rect 14019 35015 14053 35047
rect 14092 35015 14126 35047
rect 14165 35015 14199 35047
rect 14238 35015 14272 35047
rect 14311 35015 14345 35047
rect 14384 35015 14418 35047
rect 13216 34943 13250 34977
rect 13289 34943 13323 34977
rect 13362 34943 13396 34977
rect 13435 34943 13469 34977
rect 13508 34943 13542 34977
rect 13581 34943 13615 34977
rect 13654 34943 13688 34977
rect 13727 34943 13761 34977
rect 13800 34943 13834 34977
rect 13873 34943 13907 34977
rect 13946 34943 13980 34977
rect 14019 34943 14053 34977
rect 14092 34943 14126 34977
rect 14165 34943 14199 34977
rect 14238 34943 14272 34977
rect 14311 34943 14345 34977
rect 14384 34943 14418 34977
rect 13216 34874 13250 34905
rect 13289 34874 13323 34905
rect 13362 34874 13396 34905
rect 13435 34874 13469 34905
rect 13216 34871 13236 34874
rect 13236 34871 13250 34874
rect 13289 34871 13304 34874
rect 13304 34871 13323 34874
rect 13362 34871 13372 34874
rect 13372 34871 13396 34874
rect 13435 34871 13440 34874
rect 13440 34871 13469 34874
rect 13508 34871 13542 34905
rect 13581 34874 13615 34905
rect 13654 34874 13688 34905
rect 13727 34874 13761 34905
rect 13800 34874 13834 34905
rect 13873 34874 13907 34905
rect 13946 34874 13980 34905
rect 14019 34874 14053 34905
rect 14092 34874 14126 34905
rect 14165 34874 14199 34905
rect 14238 34874 14272 34905
rect 14311 34874 14345 34905
rect 14384 34874 14418 34905
rect 13581 34871 13610 34874
rect 13610 34871 13615 34874
rect 13654 34871 13678 34874
rect 13678 34871 13688 34874
rect 13727 34871 13746 34874
rect 13746 34871 13761 34874
rect 13800 34871 13814 34874
rect 13814 34871 13834 34874
rect 13873 34871 13882 34874
rect 13882 34871 13907 34874
rect 13946 34871 13950 34874
rect 13950 34871 13980 34874
rect 14019 34871 14052 34874
rect 14052 34871 14053 34874
rect 14092 34871 14120 34874
rect 14120 34871 14126 34874
rect 14165 34871 14188 34874
rect 14188 34871 14199 34874
rect 14238 34871 14256 34874
rect 14256 34871 14272 34874
rect 14311 34871 14324 34874
rect 14324 34871 14345 34874
rect 14384 34871 14392 34874
rect 14392 34871 14418 34874
rect 13216 34805 13250 34833
rect 13289 34805 13323 34833
rect 13362 34805 13396 34833
rect 13435 34805 13469 34833
rect 13216 34799 13236 34805
rect 13236 34799 13250 34805
rect 13289 34799 13304 34805
rect 13304 34799 13323 34805
rect 13362 34799 13372 34805
rect 13372 34799 13396 34805
rect 13435 34799 13440 34805
rect 13440 34799 13469 34805
rect 13508 34799 13542 34833
rect 13581 34805 13615 34833
rect 13654 34805 13688 34833
rect 13727 34805 13761 34833
rect 13800 34805 13834 34833
rect 13873 34805 13907 34833
rect 13946 34805 13980 34833
rect 14019 34805 14053 34833
rect 14092 34805 14126 34833
rect 14165 34805 14199 34833
rect 14238 34805 14272 34833
rect 14311 34805 14345 34833
rect 14384 34805 14418 34833
rect 13581 34799 13610 34805
rect 13610 34799 13615 34805
rect 13654 34799 13678 34805
rect 13678 34799 13688 34805
rect 13727 34799 13746 34805
rect 13746 34799 13761 34805
rect 13800 34799 13814 34805
rect 13814 34799 13834 34805
rect 13873 34799 13882 34805
rect 13882 34799 13907 34805
rect 13946 34799 13950 34805
rect 13950 34799 13980 34805
rect 14019 34799 14052 34805
rect 14052 34799 14053 34805
rect 14092 34799 14120 34805
rect 14120 34799 14126 34805
rect 14165 34799 14188 34805
rect 14188 34799 14199 34805
rect 14238 34799 14256 34805
rect 14256 34799 14272 34805
rect 14311 34799 14324 34805
rect 14324 34799 14345 34805
rect 14384 34799 14392 34805
rect 14392 34799 14418 34805
rect 13216 34736 13250 34760
rect 13289 34736 13323 34760
rect 13362 34736 13396 34760
rect 13435 34736 13469 34760
rect 13216 34726 13236 34736
rect 13236 34726 13250 34736
rect 13289 34726 13304 34736
rect 13304 34726 13323 34736
rect 13362 34726 13372 34736
rect 13372 34726 13396 34736
rect 13435 34726 13440 34736
rect 13440 34726 13469 34736
rect 13508 34726 13542 34760
rect 13581 34736 13615 34760
rect 13654 34736 13688 34760
rect 13727 34736 13761 34760
rect 13800 34736 13834 34760
rect 13873 34736 13907 34760
rect 13946 34736 13980 34760
rect 14019 34736 14053 34760
rect 14092 34736 14126 34760
rect 14165 34736 14199 34760
rect 14238 34736 14272 34760
rect 14311 34736 14345 34760
rect 14384 34736 14418 34760
rect 13581 34726 13610 34736
rect 13610 34726 13615 34736
rect 13654 34726 13678 34736
rect 13678 34726 13688 34736
rect 13727 34726 13746 34736
rect 13746 34726 13761 34736
rect 13800 34726 13814 34736
rect 13814 34726 13834 34736
rect 13873 34726 13882 34736
rect 13882 34726 13907 34736
rect 13946 34726 13950 34736
rect 13950 34726 13980 34736
rect 14019 34726 14052 34736
rect 14052 34726 14053 34736
rect 14092 34726 14120 34736
rect 14120 34726 14126 34736
rect 14165 34726 14188 34736
rect 14188 34726 14199 34736
rect 14238 34726 14256 34736
rect 14256 34726 14272 34736
rect 14311 34726 14324 34736
rect 14324 34726 14345 34736
rect 14384 34726 14392 34736
rect 14392 34726 14418 34736
rect 13216 34667 13250 34687
rect 13289 34667 13323 34687
rect 13362 34667 13396 34687
rect 13435 34667 13469 34687
rect 13216 34653 13236 34667
rect 13236 34653 13250 34667
rect 13289 34653 13304 34667
rect 13304 34653 13323 34667
rect 13362 34653 13372 34667
rect 13372 34653 13396 34667
rect 13435 34653 13440 34667
rect 13440 34653 13469 34667
rect 13508 34653 13542 34687
rect 13581 34667 13615 34687
rect 13654 34667 13688 34687
rect 13727 34667 13761 34687
rect 13800 34667 13834 34687
rect 13873 34667 13907 34687
rect 13946 34667 13980 34687
rect 14019 34667 14053 34687
rect 14092 34667 14126 34687
rect 14165 34667 14199 34687
rect 14238 34667 14272 34687
rect 14311 34667 14345 34687
rect 14384 34667 14418 34687
rect 13581 34653 13610 34667
rect 13610 34653 13615 34667
rect 13654 34653 13678 34667
rect 13678 34653 13688 34667
rect 13727 34653 13746 34667
rect 13746 34653 13761 34667
rect 13800 34653 13814 34667
rect 13814 34653 13834 34667
rect 13873 34653 13882 34667
rect 13882 34653 13907 34667
rect 13946 34653 13950 34667
rect 13950 34653 13980 34667
rect 14019 34653 14052 34667
rect 14052 34653 14053 34667
rect 14092 34653 14120 34667
rect 14120 34653 14126 34667
rect 14165 34653 14188 34667
rect 14188 34653 14199 34667
rect 14238 34653 14256 34667
rect 14256 34653 14272 34667
rect 14311 34653 14324 34667
rect 14324 34653 14345 34667
rect 14384 34653 14392 34667
rect 14392 34653 14418 34667
rect 13216 34598 13250 34614
rect 13289 34598 13323 34614
rect 13362 34598 13396 34614
rect 13435 34598 13469 34614
rect 13216 34580 13236 34598
rect 13236 34580 13250 34598
rect 13289 34580 13304 34598
rect 13304 34580 13323 34598
rect 13362 34580 13372 34598
rect 13372 34580 13396 34598
rect 13435 34580 13440 34598
rect 13440 34580 13469 34598
rect 13508 34580 13542 34614
rect 13581 34598 13615 34614
rect 13654 34598 13688 34614
rect 13727 34598 13761 34614
rect 13800 34598 13834 34614
rect 13873 34598 13907 34614
rect 13946 34598 13980 34614
rect 14019 34598 14053 34614
rect 14092 34598 14126 34614
rect 14165 34598 14199 34614
rect 14238 34598 14272 34614
rect 14311 34598 14345 34614
rect 14384 34598 14418 34614
rect 13581 34580 13610 34598
rect 13610 34580 13615 34598
rect 13654 34580 13678 34598
rect 13678 34580 13688 34598
rect 13727 34580 13746 34598
rect 13746 34580 13761 34598
rect 13800 34580 13814 34598
rect 13814 34580 13834 34598
rect 13873 34580 13882 34598
rect 13882 34580 13907 34598
rect 13946 34580 13950 34598
rect 13950 34580 13980 34598
rect 14019 34580 14052 34598
rect 14052 34580 14053 34598
rect 14092 34580 14120 34598
rect 14120 34580 14126 34598
rect 14165 34580 14188 34598
rect 14188 34580 14199 34598
rect 14238 34580 14256 34598
rect 14256 34580 14272 34598
rect 14311 34580 14324 34598
rect 14324 34580 14345 34598
rect 14384 34580 14392 34598
rect 14392 34580 14418 34598
rect 13216 34529 13250 34541
rect 13289 34529 13323 34541
rect 13362 34529 13396 34541
rect 13435 34529 13469 34541
rect 13216 34507 13236 34529
rect 13236 34507 13250 34529
rect 13289 34507 13304 34529
rect 13304 34507 13323 34529
rect 13362 34507 13372 34529
rect 13372 34507 13396 34529
rect 13435 34507 13440 34529
rect 13440 34507 13469 34529
rect 13508 34507 13542 34541
rect 13581 34529 13615 34541
rect 13654 34529 13688 34541
rect 13727 34529 13761 34541
rect 13800 34529 13834 34541
rect 13873 34529 13907 34541
rect 13946 34529 13980 34541
rect 14019 34529 14053 34541
rect 14092 34529 14126 34541
rect 14165 34529 14199 34541
rect 14238 34529 14272 34541
rect 14311 34529 14345 34541
rect 14384 34529 14418 34541
rect 13581 34507 13610 34529
rect 13610 34507 13615 34529
rect 13654 34507 13678 34529
rect 13678 34507 13688 34529
rect 13727 34507 13746 34529
rect 13746 34507 13761 34529
rect 13800 34507 13814 34529
rect 13814 34507 13834 34529
rect 13873 34507 13882 34529
rect 13882 34507 13907 34529
rect 13946 34507 13950 34529
rect 13950 34507 13980 34529
rect 14019 34507 14052 34529
rect 14052 34507 14053 34529
rect 14092 34507 14120 34529
rect 14120 34507 14126 34529
rect 14165 34507 14188 34529
rect 14188 34507 14199 34529
rect 14238 34507 14256 34529
rect 14256 34507 14272 34529
rect 14311 34507 14324 34529
rect 14324 34507 14345 34529
rect 14384 34507 14392 34529
rect 14392 34507 14418 34529
rect 13216 34460 13250 34468
rect 13289 34460 13323 34468
rect 13362 34460 13396 34468
rect 13435 34460 13469 34468
rect 13216 34434 13236 34460
rect 13236 34434 13250 34460
rect 13289 34434 13304 34460
rect 13304 34434 13323 34460
rect 13362 34434 13372 34460
rect 13372 34434 13396 34460
rect 13435 34434 13440 34460
rect 13440 34434 13469 34460
rect 13508 34434 13542 34468
rect 13581 34460 13615 34468
rect 13654 34460 13688 34468
rect 13727 34460 13761 34468
rect 13800 34460 13834 34468
rect 13873 34460 13907 34468
rect 13946 34460 13980 34468
rect 14019 34460 14053 34468
rect 14092 34460 14126 34468
rect 14165 34460 14199 34468
rect 14238 34460 14272 34468
rect 14311 34460 14345 34468
rect 14384 34460 14418 34468
rect 13581 34434 13610 34460
rect 13610 34434 13615 34460
rect 13654 34434 13678 34460
rect 13678 34434 13688 34460
rect 13727 34434 13746 34460
rect 13746 34434 13761 34460
rect 13800 34434 13814 34460
rect 13814 34434 13834 34460
rect 13873 34434 13882 34460
rect 13882 34434 13907 34460
rect 13946 34434 13950 34460
rect 13950 34434 13980 34460
rect 14019 34434 14052 34460
rect 14052 34434 14053 34460
rect 14092 34434 14120 34460
rect 14120 34434 14126 34460
rect 14165 34434 14188 34460
rect 14188 34434 14199 34460
rect 14238 34434 14256 34460
rect 14256 34434 14272 34460
rect 14311 34434 14324 34460
rect 14324 34434 14345 34460
rect 14384 34434 14392 34460
rect 14392 34434 14418 34460
rect 13216 34391 13250 34395
rect 13289 34391 13323 34395
rect 13362 34391 13396 34395
rect 13435 34391 13469 34395
rect 13216 34361 13236 34391
rect 13236 34361 13250 34391
rect 13289 34361 13304 34391
rect 13304 34361 13323 34391
rect 13362 34361 13372 34391
rect 13372 34361 13396 34391
rect 13435 34361 13440 34391
rect 13440 34361 13469 34391
rect 13508 34361 13542 34395
rect 13581 34391 13615 34395
rect 13654 34391 13688 34395
rect 13727 34391 13761 34395
rect 13800 34391 13834 34395
rect 13873 34391 13907 34395
rect 13946 34391 13980 34395
rect 14019 34391 14053 34395
rect 14092 34391 14126 34395
rect 14165 34391 14199 34395
rect 14238 34391 14272 34395
rect 14311 34391 14345 34395
rect 14384 34391 14418 34395
rect 13581 34361 13610 34391
rect 13610 34361 13615 34391
rect 13654 34361 13678 34391
rect 13678 34361 13688 34391
rect 13727 34361 13746 34391
rect 13746 34361 13761 34391
rect 13800 34361 13814 34391
rect 13814 34361 13834 34391
rect 13873 34361 13882 34391
rect 13882 34361 13907 34391
rect 13946 34361 13950 34391
rect 13950 34361 13980 34391
rect 14019 34361 14052 34391
rect 14052 34361 14053 34391
rect 14092 34361 14120 34391
rect 14120 34361 14126 34391
rect 14165 34361 14188 34391
rect 14188 34361 14199 34391
rect 14238 34361 14256 34391
rect 14256 34361 14272 34391
rect 14311 34361 14324 34391
rect 14324 34361 14345 34391
rect 14384 34361 14392 34391
rect 14392 34361 14418 34391
rect 13216 34288 13236 34322
rect 13236 34288 13250 34322
rect 13289 34288 13304 34322
rect 13304 34288 13323 34322
rect 13362 34288 13372 34322
rect 13372 34288 13396 34322
rect 13435 34288 13440 34322
rect 13440 34288 13469 34322
rect 13508 34288 13542 34322
rect 13581 34288 13610 34322
rect 13610 34288 13615 34322
rect 13654 34288 13678 34322
rect 13678 34288 13688 34322
rect 13727 34288 13746 34322
rect 13746 34288 13761 34322
rect 13800 34288 13814 34322
rect 13814 34288 13834 34322
rect 13873 34288 13882 34322
rect 13882 34288 13907 34322
rect 13946 34288 13950 34322
rect 13950 34288 13980 34322
rect 14019 34288 14052 34322
rect 14052 34288 14053 34322
rect 14092 34288 14120 34322
rect 14120 34288 14126 34322
rect 14165 34288 14188 34322
rect 14188 34288 14199 34322
rect 14238 34288 14256 34322
rect 14256 34288 14272 34322
rect 14311 34288 14324 34322
rect 14324 34288 14345 34322
rect 14384 34288 14392 34322
rect 14392 34288 14418 34322
rect 13216 34219 13236 34249
rect 13236 34219 13250 34249
rect 13289 34219 13304 34249
rect 13304 34219 13323 34249
rect 13362 34219 13372 34249
rect 13372 34219 13396 34249
rect 13435 34219 13440 34249
rect 13440 34219 13469 34249
rect 13216 34215 13250 34219
rect 13289 34215 13323 34219
rect 13362 34215 13396 34219
rect 13435 34215 13469 34219
rect 13508 34215 13542 34249
rect 13581 34219 13610 34249
rect 13610 34219 13615 34249
rect 13654 34219 13678 34249
rect 13678 34219 13688 34249
rect 13727 34219 13746 34249
rect 13746 34219 13761 34249
rect 13800 34219 13814 34249
rect 13814 34219 13834 34249
rect 13873 34219 13882 34249
rect 13882 34219 13907 34249
rect 13946 34219 13950 34249
rect 13950 34219 13980 34249
rect 14019 34219 14052 34249
rect 14052 34219 14053 34249
rect 14092 34219 14120 34249
rect 14120 34219 14126 34249
rect 14165 34219 14188 34249
rect 14188 34219 14199 34249
rect 14238 34219 14256 34249
rect 14256 34219 14272 34249
rect 14311 34219 14324 34249
rect 14324 34219 14345 34249
rect 14384 34219 14392 34249
rect 14392 34219 14418 34249
rect 13581 34215 13615 34219
rect 13654 34215 13688 34219
rect 13727 34215 13761 34219
rect 13800 34215 13834 34219
rect 13873 34215 13907 34219
rect 13946 34215 13980 34219
rect 14019 34215 14053 34219
rect 14092 34215 14126 34219
rect 14165 34215 14199 34219
rect 14238 34215 14272 34219
rect 14311 34215 14345 34219
rect 14384 34215 14418 34219
rect 13216 34150 13236 34176
rect 13236 34150 13250 34176
rect 13289 34150 13304 34176
rect 13304 34150 13323 34176
rect 13362 34150 13372 34176
rect 13372 34150 13396 34176
rect 13435 34150 13440 34176
rect 13440 34150 13469 34176
rect 13216 34142 13250 34150
rect 13289 34142 13323 34150
rect 13362 34142 13396 34150
rect 13435 34142 13469 34150
rect 13508 34142 13542 34176
rect 13581 34150 13610 34176
rect 13610 34150 13615 34176
rect 13654 34150 13678 34176
rect 13678 34150 13688 34176
rect 13727 34150 13746 34176
rect 13746 34150 13761 34176
rect 13800 34150 13814 34176
rect 13814 34150 13834 34176
rect 13873 34150 13882 34176
rect 13882 34150 13907 34176
rect 13946 34150 13950 34176
rect 13950 34150 13980 34176
rect 14019 34150 14052 34176
rect 14052 34150 14053 34176
rect 14092 34150 14120 34176
rect 14120 34150 14126 34176
rect 14165 34150 14188 34176
rect 14188 34150 14199 34176
rect 14238 34150 14256 34176
rect 14256 34150 14272 34176
rect 14311 34150 14324 34176
rect 14324 34150 14345 34176
rect 14384 34150 14392 34176
rect 14392 34150 14418 34176
rect 13581 34142 13615 34150
rect 13654 34142 13688 34150
rect 13727 34142 13761 34150
rect 13800 34142 13834 34150
rect 13873 34142 13907 34150
rect 13946 34142 13980 34150
rect 14019 34142 14053 34150
rect 14092 34142 14126 34150
rect 14165 34142 14199 34150
rect 14238 34142 14272 34150
rect 14311 34142 14345 34150
rect 14384 34142 14418 34150
rect 13216 34081 13236 34103
rect 13236 34081 13250 34103
rect 13289 34081 13304 34103
rect 13304 34081 13323 34103
rect 13362 34081 13372 34103
rect 13372 34081 13396 34103
rect 13435 34081 13440 34103
rect 13440 34081 13469 34103
rect 13216 34069 13250 34081
rect 13289 34069 13323 34081
rect 13362 34069 13396 34081
rect 13435 34069 13469 34081
rect 13508 34069 13542 34103
rect 13581 34081 13610 34103
rect 13610 34081 13615 34103
rect 13654 34081 13678 34103
rect 13678 34081 13688 34103
rect 13727 34081 13746 34103
rect 13746 34081 13761 34103
rect 13800 34081 13814 34103
rect 13814 34081 13834 34103
rect 13873 34081 13882 34103
rect 13882 34081 13907 34103
rect 13946 34081 13950 34103
rect 13950 34081 13980 34103
rect 14019 34081 14052 34103
rect 14052 34081 14053 34103
rect 14092 34081 14120 34103
rect 14120 34081 14126 34103
rect 14165 34081 14188 34103
rect 14188 34081 14199 34103
rect 14238 34081 14256 34103
rect 14256 34081 14272 34103
rect 14311 34081 14324 34103
rect 14324 34081 14345 34103
rect 14384 34081 14392 34103
rect 14392 34081 14418 34103
rect 13581 34069 13615 34081
rect 13654 34069 13688 34081
rect 13727 34069 13761 34081
rect 13800 34069 13834 34081
rect 13873 34069 13907 34081
rect 13946 34069 13980 34081
rect 14019 34069 14053 34081
rect 14092 34069 14126 34081
rect 14165 34069 14199 34081
rect 14238 34069 14272 34081
rect 14311 34069 14345 34081
rect 14384 34069 14418 34081
rect 13216 34012 13236 34030
rect 13236 34012 13250 34030
rect 13289 34012 13304 34030
rect 13304 34012 13323 34030
rect 13362 34012 13372 34030
rect 13372 34012 13396 34030
rect 13435 34012 13440 34030
rect 13440 34012 13469 34030
rect 13216 33996 13250 34012
rect 13289 33996 13323 34012
rect 13362 33996 13396 34012
rect 13435 33996 13469 34012
rect 13508 33996 13542 34030
rect 13581 34012 13610 34030
rect 13610 34012 13615 34030
rect 13654 34012 13678 34030
rect 13678 34012 13688 34030
rect 13727 34012 13746 34030
rect 13746 34012 13761 34030
rect 13800 34012 13814 34030
rect 13814 34012 13834 34030
rect 13873 34012 13882 34030
rect 13882 34012 13907 34030
rect 13946 34012 13950 34030
rect 13950 34012 13980 34030
rect 14019 34012 14052 34030
rect 14052 34012 14053 34030
rect 14092 34012 14120 34030
rect 14120 34012 14126 34030
rect 14165 34012 14188 34030
rect 14188 34012 14199 34030
rect 14238 34012 14256 34030
rect 14256 34012 14272 34030
rect 14311 34012 14324 34030
rect 14324 34012 14345 34030
rect 14384 34012 14392 34030
rect 14392 34012 14418 34030
rect 13581 33996 13615 34012
rect 13654 33996 13688 34012
rect 13727 33996 13761 34012
rect 13800 33996 13834 34012
rect 13873 33996 13907 34012
rect 13946 33996 13980 34012
rect 14019 33996 14053 34012
rect 14092 33996 14126 34012
rect 14165 33996 14199 34012
rect 14238 33996 14272 34012
rect 14311 33996 14345 34012
rect 14384 33996 14418 34012
rect 13216 33943 13236 33957
rect 13236 33943 13250 33957
rect 13289 33943 13304 33957
rect 13304 33943 13323 33957
rect 13362 33943 13372 33957
rect 13372 33943 13396 33957
rect 13435 33943 13440 33957
rect 13440 33943 13469 33957
rect 13216 33923 13250 33943
rect 13289 33923 13323 33943
rect 13362 33923 13396 33943
rect 13435 33923 13469 33943
rect 13508 33923 13542 33957
rect 13581 33943 13610 33957
rect 13610 33943 13615 33957
rect 13654 33943 13678 33957
rect 13678 33943 13688 33957
rect 13727 33943 13746 33957
rect 13746 33943 13761 33957
rect 13800 33943 13814 33957
rect 13814 33943 13834 33957
rect 13873 33943 13882 33957
rect 13882 33943 13907 33957
rect 13946 33943 13950 33957
rect 13950 33943 13980 33957
rect 14019 33943 14052 33957
rect 14052 33943 14053 33957
rect 14092 33943 14120 33957
rect 14120 33943 14126 33957
rect 14165 33943 14188 33957
rect 14188 33943 14199 33957
rect 14238 33943 14256 33957
rect 14256 33943 14272 33957
rect 14311 33943 14324 33957
rect 14324 33943 14345 33957
rect 14384 33943 14392 33957
rect 14392 33943 14418 33957
rect 13581 33923 13615 33943
rect 13654 33923 13688 33943
rect 13727 33923 13761 33943
rect 13800 33923 13834 33943
rect 13873 33923 13907 33943
rect 13946 33923 13980 33943
rect 14019 33923 14053 33943
rect 14092 33923 14126 33943
rect 14165 33923 14199 33943
rect 14238 33923 14272 33943
rect 14311 33923 14345 33943
rect 14384 33923 14418 33943
rect 13216 33874 13236 33884
rect 13236 33874 13250 33884
rect 13289 33874 13304 33884
rect 13304 33874 13323 33884
rect 13362 33874 13372 33884
rect 13372 33874 13396 33884
rect 13435 33874 13440 33884
rect 13440 33874 13469 33884
rect 13216 33850 13250 33874
rect 13289 33850 13323 33874
rect 13362 33850 13396 33874
rect 13435 33850 13469 33874
rect 13508 33850 13542 33884
rect 13581 33874 13610 33884
rect 13610 33874 13615 33884
rect 13654 33874 13678 33884
rect 13678 33874 13688 33884
rect 13727 33874 13746 33884
rect 13746 33874 13761 33884
rect 13800 33874 13814 33884
rect 13814 33874 13834 33884
rect 13873 33874 13882 33884
rect 13882 33874 13907 33884
rect 13946 33874 13950 33884
rect 13950 33874 13980 33884
rect 14019 33874 14052 33884
rect 14052 33874 14053 33884
rect 14092 33874 14120 33884
rect 14120 33874 14126 33884
rect 14165 33874 14188 33884
rect 14188 33874 14199 33884
rect 14238 33874 14256 33884
rect 14256 33874 14272 33884
rect 14311 33874 14324 33884
rect 14324 33874 14345 33884
rect 14384 33874 14392 33884
rect 14392 33874 14418 33884
rect 13581 33850 13615 33874
rect 13654 33850 13688 33874
rect 13727 33850 13761 33874
rect 13800 33850 13834 33874
rect 13873 33850 13907 33874
rect 13946 33850 13980 33874
rect 14019 33850 14053 33874
rect 14092 33850 14126 33874
rect 14165 33850 14199 33874
rect 14238 33850 14272 33874
rect 14311 33850 14345 33874
rect 14384 33850 14418 33874
rect 13216 33805 13236 33811
rect 13236 33805 13250 33811
rect 13289 33805 13304 33811
rect 13304 33805 13323 33811
rect 13362 33805 13372 33811
rect 13372 33805 13396 33811
rect 13435 33805 13440 33811
rect 13440 33805 13469 33811
rect 13216 33777 13250 33805
rect 13289 33777 13323 33805
rect 13362 33777 13396 33805
rect 13435 33777 13469 33805
rect 13508 33777 13542 33811
rect 13581 33805 13610 33811
rect 13610 33805 13615 33811
rect 13654 33805 13678 33811
rect 13678 33805 13688 33811
rect 13727 33805 13746 33811
rect 13746 33805 13761 33811
rect 13800 33805 13814 33811
rect 13814 33805 13834 33811
rect 13873 33805 13882 33811
rect 13882 33805 13907 33811
rect 13946 33805 13950 33811
rect 13950 33805 13980 33811
rect 14019 33805 14052 33811
rect 14052 33805 14053 33811
rect 14092 33805 14120 33811
rect 14120 33805 14126 33811
rect 14165 33805 14188 33811
rect 14188 33805 14199 33811
rect 14238 33805 14256 33811
rect 14256 33805 14272 33811
rect 14311 33805 14324 33811
rect 14324 33805 14345 33811
rect 14384 33805 14392 33811
rect 14392 33805 14418 33811
rect 13581 33777 13615 33805
rect 13654 33777 13688 33805
rect 13727 33777 13761 33805
rect 13800 33777 13834 33805
rect 13873 33777 13907 33805
rect 13946 33777 13980 33805
rect 14019 33777 14053 33805
rect 14092 33777 14126 33805
rect 14165 33777 14199 33805
rect 14238 33777 14272 33805
rect 14311 33777 14345 33805
rect 14384 33777 14418 33805
rect 13216 33736 13236 33738
rect 13236 33736 13250 33738
rect 13289 33736 13304 33738
rect 13304 33736 13323 33738
rect 13362 33736 13372 33738
rect 13372 33736 13396 33738
rect 13435 33736 13440 33738
rect 13440 33736 13469 33738
rect 13216 33704 13250 33736
rect 13289 33704 13323 33736
rect 13362 33704 13396 33736
rect 13435 33704 13469 33736
rect 13508 33704 13542 33738
rect 13581 33736 13610 33738
rect 13610 33736 13615 33738
rect 13654 33736 13678 33738
rect 13678 33736 13688 33738
rect 13727 33736 13746 33738
rect 13746 33736 13761 33738
rect 13800 33736 13814 33738
rect 13814 33736 13834 33738
rect 13873 33736 13882 33738
rect 13882 33736 13907 33738
rect 13946 33736 13950 33738
rect 13950 33736 13980 33738
rect 14019 33736 14052 33738
rect 14052 33736 14053 33738
rect 14092 33736 14120 33738
rect 14120 33736 14126 33738
rect 14165 33736 14188 33738
rect 14188 33736 14199 33738
rect 14238 33736 14256 33738
rect 14256 33736 14272 33738
rect 14311 33736 14324 33738
rect 14324 33736 14345 33738
rect 14384 33736 14392 33738
rect 14392 33736 14418 33738
rect 13581 33704 13615 33736
rect 13654 33704 13688 33736
rect 13727 33704 13761 33736
rect 13800 33704 13834 33736
rect 13873 33704 13907 33736
rect 13946 33704 13980 33736
rect 14019 33704 14053 33736
rect 14092 33704 14126 33736
rect 14165 33704 14199 33736
rect 14238 33704 14272 33736
rect 14311 33704 14345 33736
rect 14384 33704 14418 33736
rect 13216 33632 13250 33665
rect 13289 33632 13323 33665
rect 13362 33632 13396 33665
rect 13435 33632 13469 33665
rect 13216 33631 13236 33632
rect 13236 33631 13250 33632
rect 13289 33631 13304 33632
rect 13304 33631 13323 33632
rect 13362 33631 13372 33632
rect 13372 33631 13396 33632
rect 13435 33631 13440 33632
rect 13440 33631 13469 33632
rect 13508 33631 13542 33665
rect 13581 33632 13615 33665
rect 13654 33632 13688 33665
rect 13727 33632 13761 33665
rect 13800 33632 13834 33665
rect 13873 33632 13907 33665
rect 13946 33632 13980 33665
rect 14019 33632 14053 33665
rect 14092 33632 14126 33665
rect 14165 33632 14199 33665
rect 14238 33632 14272 33665
rect 14311 33632 14345 33665
rect 14384 33632 14418 33665
rect 13581 33631 13610 33632
rect 13610 33631 13615 33632
rect 13654 33631 13678 33632
rect 13678 33631 13688 33632
rect 13727 33631 13746 33632
rect 13746 33631 13761 33632
rect 13800 33631 13814 33632
rect 13814 33631 13834 33632
rect 13873 33631 13882 33632
rect 13882 33631 13907 33632
rect 13946 33631 13950 33632
rect 13950 33631 13980 33632
rect 14019 33631 14052 33632
rect 14052 33631 14053 33632
rect 14092 33631 14120 33632
rect 14120 33631 14126 33632
rect 14165 33631 14188 33632
rect 14188 33631 14199 33632
rect 14238 33631 14256 33632
rect 14256 33631 14272 33632
rect 14311 33631 14324 33632
rect 14324 33631 14345 33632
rect 14384 33631 14392 33632
rect 14392 33631 14418 33632
rect 13216 33563 13250 33592
rect 13289 33563 13323 33592
rect 13362 33563 13396 33592
rect 13435 33563 13469 33592
rect 13216 33558 13236 33563
rect 13236 33558 13250 33563
rect 13289 33558 13304 33563
rect 13304 33558 13323 33563
rect 13362 33558 13372 33563
rect 13372 33558 13396 33563
rect 13435 33558 13440 33563
rect 13440 33558 13469 33563
rect 13508 33558 13542 33592
rect 13581 33563 13615 33592
rect 13654 33563 13688 33592
rect 13727 33563 13761 33592
rect 13800 33563 13834 33592
rect 13873 33563 13907 33592
rect 13946 33563 13980 33592
rect 14019 33563 14053 33592
rect 14092 33563 14126 33592
rect 14165 33563 14199 33592
rect 14238 33563 14272 33592
rect 14311 33563 14345 33592
rect 14384 33563 14418 33592
rect 13581 33558 13610 33563
rect 13610 33558 13615 33563
rect 13654 33558 13678 33563
rect 13678 33558 13688 33563
rect 13727 33558 13746 33563
rect 13746 33558 13761 33563
rect 13800 33558 13814 33563
rect 13814 33558 13834 33563
rect 13873 33558 13882 33563
rect 13882 33558 13907 33563
rect 13946 33558 13950 33563
rect 13950 33558 13980 33563
rect 14019 33558 14052 33563
rect 14052 33558 14053 33563
rect 14092 33558 14120 33563
rect 14120 33558 14126 33563
rect 14165 33558 14188 33563
rect 14188 33558 14199 33563
rect 14238 33558 14256 33563
rect 14256 33558 14272 33563
rect 14311 33558 14324 33563
rect 14324 33558 14345 33563
rect 14384 33558 14392 33563
rect 14392 33558 14418 33563
rect 13216 33494 13250 33519
rect 13289 33494 13323 33519
rect 13362 33494 13396 33519
rect 13435 33494 13469 33519
rect 13216 33485 13236 33494
rect 13236 33485 13250 33494
rect 13289 33485 13304 33494
rect 13304 33485 13323 33494
rect 13362 33485 13372 33494
rect 13372 33485 13396 33494
rect 13435 33485 13440 33494
rect 13440 33485 13469 33494
rect 13508 33485 13542 33519
rect 13581 33494 13615 33519
rect 13654 33494 13688 33519
rect 13727 33494 13761 33519
rect 13800 33494 13834 33519
rect 13873 33494 13907 33519
rect 13946 33494 13980 33519
rect 14019 33494 14053 33519
rect 14092 33494 14126 33519
rect 14165 33494 14199 33519
rect 14238 33494 14272 33519
rect 14311 33494 14345 33519
rect 14384 33494 14418 33519
rect 13581 33485 13610 33494
rect 13610 33485 13615 33494
rect 13654 33485 13678 33494
rect 13678 33485 13688 33494
rect 13727 33485 13746 33494
rect 13746 33485 13761 33494
rect 13800 33485 13814 33494
rect 13814 33485 13834 33494
rect 13873 33485 13882 33494
rect 13882 33485 13907 33494
rect 13946 33485 13950 33494
rect 13950 33485 13980 33494
rect 14019 33485 14052 33494
rect 14052 33485 14053 33494
rect 14092 33485 14120 33494
rect 14120 33485 14126 33494
rect 14165 33485 14188 33494
rect 14188 33485 14199 33494
rect 14238 33485 14256 33494
rect 14256 33485 14272 33494
rect 14311 33485 14324 33494
rect 14324 33485 14345 33494
rect 14384 33485 14392 33494
rect 14392 33485 14418 33494
rect 13216 33425 13250 33446
rect 13289 33425 13323 33446
rect 13362 33425 13396 33446
rect 13435 33425 13469 33446
rect 13216 33412 13236 33425
rect 13236 33412 13250 33425
rect 13289 33412 13304 33425
rect 13304 33412 13323 33425
rect 13362 33412 13372 33425
rect 13372 33412 13396 33425
rect 13435 33412 13440 33425
rect 13440 33412 13469 33425
rect 13508 33412 13542 33446
rect 13581 33425 13615 33446
rect 13654 33425 13688 33446
rect 13727 33425 13761 33446
rect 13800 33425 13834 33446
rect 13873 33425 13907 33446
rect 13946 33425 13980 33446
rect 14019 33425 14053 33446
rect 14092 33425 14126 33446
rect 14165 33425 14199 33446
rect 14238 33425 14272 33446
rect 14311 33425 14345 33446
rect 14384 33425 14418 33446
rect 13581 33412 13610 33425
rect 13610 33412 13615 33425
rect 13654 33412 13678 33425
rect 13678 33412 13688 33425
rect 13727 33412 13746 33425
rect 13746 33412 13761 33425
rect 13800 33412 13814 33425
rect 13814 33412 13834 33425
rect 13873 33412 13882 33425
rect 13882 33412 13907 33425
rect 13946 33412 13950 33425
rect 13950 33412 13980 33425
rect 14019 33412 14052 33425
rect 14052 33412 14053 33425
rect 14092 33412 14120 33425
rect 14120 33412 14126 33425
rect 14165 33412 14188 33425
rect 14188 33412 14199 33425
rect 14238 33412 14256 33425
rect 14256 33412 14272 33425
rect 14311 33412 14324 33425
rect 14324 33412 14345 33425
rect 14384 33412 14392 33425
rect 14392 33412 14418 33425
rect 13216 33356 13250 33373
rect 13289 33356 13323 33373
rect 13362 33356 13396 33373
rect 13435 33356 13469 33373
rect 13216 33339 13236 33356
rect 13236 33339 13250 33356
rect 13289 33339 13304 33356
rect 13304 33339 13323 33356
rect 13362 33339 13372 33356
rect 13372 33339 13396 33356
rect 13435 33339 13440 33356
rect 13440 33339 13469 33356
rect 13508 33339 13542 33373
rect 13581 33356 13615 33373
rect 13654 33356 13688 33373
rect 13727 33356 13761 33373
rect 13800 33356 13834 33373
rect 13873 33356 13907 33373
rect 13946 33356 13980 33373
rect 14019 33356 14053 33373
rect 14092 33356 14126 33373
rect 14165 33356 14199 33373
rect 14238 33356 14272 33373
rect 14311 33356 14345 33373
rect 14384 33356 14418 33373
rect 13581 33339 13610 33356
rect 13610 33339 13615 33356
rect 13654 33339 13678 33356
rect 13678 33339 13688 33356
rect 13727 33339 13746 33356
rect 13746 33339 13761 33356
rect 13800 33339 13814 33356
rect 13814 33339 13834 33356
rect 13873 33339 13882 33356
rect 13882 33339 13907 33356
rect 13946 33339 13950 33356
rect 13950 33339 13980 33356
rect 14019 33339 14052 33356
rect 14052 33339 14053 33356
rect 14092 33339 14120 33356
rect 14120 33339 14126 33356
rect 14165 33339 14188 33356
rect 14188 33339 14199 33356
rect 14238 33339 14256 33356
rect 14256 33339 14272 33356
rect 14311 33339 14324 33356
rect 14324 33339 14345 33356
rect 14384 33339 14392 33356
rect 14392 33339 14418 33356
rect 13216 33287 13250 33300
rect 13289 33287 13323 33300
rect 13362 33287 13396 33300
rect 13435 33287 13469 33300
rect 13216 33266 13236 33287
rect 13236 33266 13250 33287
rect 13289 33266 13304 33287
rect 13304 33266 13323 33287
rect 13362 33266 13372 33287
rect 13372 33266 13396 33287
rect 13435 33266 13440 33287
rect 13440 33266 13469 33287
rect 13508 33266 13542 33300
rect 13581 33287 13615 33300
rect 13654 33287 13688 33300
rect 13727 33287 13761 33300
rect 13800 33287 13834 33300
rect 13873 33287 13907 33300
rect 13946 33287 13980 33300
rect 14019 33287 14053 33300
rect 14092 33287 14126 33300
rect 14165 33287 14199 33300
rect 14238 33287 14272 33300
rect 14311 33287 14345 33300
rect 14384 33287 14418 33300
rect 13581 33266 13610 33287
rect 13610 33266 13615 33287
rect 13654 33266 13678 33287
rect 13678 33266 13688 33287
rect 13727 33266 13746 33287
rect 13746 33266 13761 33287
rect 13800 33266 13814 33287
rect 13814 33266 13834 33287
rect 13873 33266 13882 33287
rect 13882 33266 13907 33287
rect 13946 33266 13950 33287
rect 13950 33266 13980 33287
rect 14019 33266 14052 33287
rect 14052 33266 14053 33287
rect 14092 33266 14120 33287
rect 14120 33266 14126 33287
rect 14165 33266 14188 33287
rect 14188 33266 14199 33287
rect 14238 33266 14256 33287
rect 14256 33266 14272 33287
rect 14311 33266 14324 33287
rect 14324 33266 14345 33287
rect 14384 33266 14392 33287
rect 14392 33266 14418 33287
rect 13216 33218 13250 33227
rect 13289 33218 13323 33227
rect 13362 33218 13396 33227
rect 13435 33218 13469 33227
rect 13216 33193 13236 33218
rect 13236 33193 13250 33218
rect 13289 33193 13304 33218
rect 13304 33193 13323 33218
rect 13362 33193 13372 33218
rect 13372 33193 13396 33218
rect 13435 33193 13440 33218
rect 13440 33193 13469 33218
rect 13508 33193 13542 33227
rect 13581 33218 13615 33227
rect 13654 33218 13688 33227
rect 13727 33218 13761 33227
rect 13800 33218 13834 33227
rect 13873 33218 13907 33227
rect 13946 33218 13980 33227
rect 14019 33218 14053 33227
rect 14092 33218 14126 33227
rect 14165 33218 14199 33227
rect 14238 33218 14272 33227
rect 14311 33218 14345 33227
rect 14384 33218 14418 33227
rect 13581 33193 13610 33218
rect 13610 33193 13615 33218
rect 13654 33193 13678 33218
rect 13678 33193 13688 33218
rect 13727 33193 13746 33218
rect 13746 33193 13761 33218
rect 13800 33193 13814 33218
rect 13814 33193 13834 33218
rect 13873 33193 13882 33218
rect 13882 33193 13907 33218
rect 13946 33193 13950 33218
rect 13950 33193 13980 33218
rect 14019 33193 14052 33218
rect 14052 33193 14053 33218
rect 14092 33193 14120 33218
rect 14120 33193 14126 33218
rect 14165 33193 14188 33218
rect 14188 33193 14199 33218
rect 14238 33193 14256 33218
rect 14256 33193 14272 33218
rect 14311 33193 14324 33218
rect 14324 33193 14345 33218
rect 14384 33193 14392 33218
rect 14392 33193 14418 33218
rect 13216 33149 13250 33154
rect 13289 33149 13323 33154
rect 13362 33149 13396 33154
rect 13435 33149 13469 33154
rect 13216 33120 13236 33149
rect 13236 33120 13250 33149
rect 13289 33120 13304 33149
rect 13304 33120 13323 33149
rect 13362 33120 13372 33149
rect 13372 33120 13396 33149
rect 13435 33120 13440 33149
rect 13440 33120 13469 33149
rect 13508 33120 13542 33154
rect 13581 33149 13615 33154
rect 13654 33149 13688 33154
rect 13727 33149 13761 33154
rect 13800 33149 13834 33154
rect 13873 33149 13907 33154
rect 13946 33149 13980 33154
rect 14019 33149 14053 33154
rect 14092 33149 14126 33154
rect 14165 33149 14199 33154
rect 14238 33149 14272 33154
rect 14311 33149 14345 33154
rect 14384 33149 14418 33154
rect 13581 33120 13610 33149
rect 13610 33120 13615 33149
rect 13654 33120 13678 33149
rect 13678 33120 13688 33149
rect 13727 33120 13746 33149
rect 13746 33120 13761 33149
rect 13800 33120 13814 33149
rect 13814 33120 13834 33149
rect 13873 33120 13882 33149
rect 13882 33120 13907 33149
rect 13946 33120 13950 33149
rect 13950 33120 13980 33149
rect 14019 33120 14052 33149
rect 14052 33120 14053 33149
rect 14092 33120 14120 33149
rect 14120 33120 14126 33149
rect 14165 33120 14188 33149
rect 14188 33120 14199 33149
rect 14238 33120 14256 33149
rect 14256 33120 14272 33149
rect 14311 33120 14324 33149
rect 14324 33120 14345 33149
rect 14384 33120 14392 33149
rect 14392 33120 14418 33149
rect 13216 33080 13250 33081
rect 13289 33080 13323 33081
rect 13362 33080 13396 33081
rect 13435 33080 13469 33081
rect 13216 33047 13236 33080
rect 13236 33047 13250 33080
rect 13289 33047 13304 33080
rect 13304 33047 13323 33080
rect 13362 33047 13372 33080
rect 13372 33047 13396 33080
rect 13435 33047 13440 33080
rect 13440 33047 13469 33080
rect 13508 33047 13542 33081
rect 13581 33080 13615 33081
rect 13654 33080 13688 33081
rect 13727 33080 13761 33081
rect 13800 33080 13834 33081
rect 13873 33080 13907 33081
rect 13946 33080 13980 33081
rect 14019 33080 14053 33081
rect 14092 33080 14126 33081
rect 14165 33080 14199 33081
rect 14238 33080 14272 33081
rect 14311 33080 14345 33081
rect 14384 33080 14418 33081
rect 13581 33047 13610 33080
rect 13610 33047 13615 33080
rect 13654 33047 13678 33080
rect 13678 33047 13688 33080
rect 13727 33047 13746 33080
rect 13746 33047 13761 33080
rect 13800 33047 13814 33080
rect 13814 33047 13834 33080
rect 13873 33047 13882 33080
rect 13882 33047 13907 33080
rect 13946 33047 13950 33080
rect 13950 33047 13980 33080
rect 14019 33047 14052 33080
rect 14052 33047 14053 33080
rect 14092 33047 14120 33080
rect 14120 33047 14126 33080
rect 14165 33047 14188 33080
rect 14188 33047 14199 33080
rect 14238 33047 14256 33080
rect 14256 33047 14272 33080
rect 14311 33047 14324 33080
rect 14324 33047 14345 33080
rect 14384 33047 14392 33080
rect 14392 33047 14418 33080
rect 13216 32977 13236 33008
rect 13236 32977 13250 33008
rect 13289 32977 13304 33008
rect 13304 32977 13323 33008
rect 13362 32977 13372 33008
rect 13372 32977 13396 33008
rect 13435 32977 13440 33008
rect 13440 32977 13469 33008
rect 13216 32974 13250 32977
rect 13289 32974 13323 32977
rect 13362 32974 13396 32977
rect 13435 32974 13469 32977
rect 13508 32974 13542 33008
rect 13581 32977 13610 33008
rect 13610 32977 13615 33008
rect 13654 32977 13678 33008
rect 13678 32977 13688 33008
rect 13727 32977 13746 33008
rect 13746 32977 13761 33008
rect 13800 32977 13814 33008
rect 13814 32977 13834 33008
rect 13873 32977 13882 33008
rect 13882 32977 13907 33008
rect 13946 32977 13950 33008
rect 13950 32977 13980 33008
rect 14019 32977 14052 33008
rect 14052 32977 14053 33008
rect 14092 32977 14120 33008
rect 14120 32977 14126 33008
rect 14165 32977 14188 33008
rect 14188 32977 14199 33008
rect 14238 32977 14256 33008
rect 14256 32977 14272 33008
rect 14311 32977 14324 33008
rect 14324 32977 14345 33008
rect 14384 32977 14392 33008
rect 14392 32977 14418 33008
rect 13581 32974 13615 32977
rect 13654 32974 13688 32977
rect 13727 32974 13761 32977
rect 13800 32974 13834 32977
rect 13873 32974 13907 32977
rect 13946 32974 13980 32977
rect 14019 32974 14053 32977
rect 14092 32974 14126 32977
rect 14165 32974 14199 32977
rect 14238 32974 14272 32977
rect 14311 32974 14345 32977
rect 14384 32974 14418 32977
rect 13216 32908 13236 32935
rect 13236 32908 13250 32935
rect 13289 32908 13304 32935
rect 13304 32908 13323 32935
rect 13362 32908 13372 32935
rect 13372 32908 13396 32935
rect 13435 32908 13440 32935
rect 13440 32908 13469 32935
rect 13216 32901 13250 32908
rect 13289 32901 13323 32908
rect 13362 32901 13396 32908
rect 13435 32901 13469 32908
rect 13508 32901 13542 32935
rect 13581 32908 13610 32935
rect 13610 32908 13615 32935
rect 13654 32908 13678 32935
rect 13678 32908 13688 32935
rect 13727 32908 13746 32935
rect 13746 32908 13761 32935
rect 13800 32908 13814 32935
rect 13814 32908 13834 32935
rect 13873 32908 13882 32935
rect 13882 32908 13907 32935
rect 13946 32908 13950 32935
rect 13950 32908 13980 32935
rect 14019 32908 14052 32935
rect 14052 32908 14053 32935
rect 14092 32908 14120 32935
rect 14120 32908 14126 32935
rect 14165 32908 14188 32935
rect 14188 32908 14199 32935
rect 14238 32908 14256 32935
rect 14256 32908 14272 32935
rect 14311 32908 14324 32935
rect 14324 32908 14345 32935
rect 14384 32908 14392 32935
rect 14392 32908 14418 32935
rect 13581 32901 13615 32908
rect 13654 32901 13688 32908
rect 13727 32901 13761 32908
rect 13800 32901 13834 32908
rect 13873 32901 13907 32908
rect 13946 32901 13980 32908
rect 14019 32901 14053 32908
rect 14092 32901 14126 32908
rect 14165 32901 14199 32908
rect 14238 32901 14272 32908
rect 14311 32901 14345 32908
rect 14384 32901 14418 32908
rect 13216 32839 13236 32862
rect 13236 32839 13250 32862
rect 13289 32839 13304 32862
rect 13304 32839 13323 32862
rect 13362 32839 13372 32862
rect 13372 32839 13396 32862
rect 13435 32839 13440 32862
rect 13440 32839 13469 32862
rect 13216 32828 13250 32839
rect 13289 32828 13323 32839
rect 13362 32828 13396 32839
rect 13435 32828 13469 32839
rect 13508 32828 13542 32862
rect 13581 32839 13610 32862
rect 13610 32839 13615 32862
rect 13654 32839 13678 32862
rect 13678 32839 13688 32862
rect 13727 32839 13746 32862
rect 13746 32839 13761 32862
rect 13800 32839 13814 32862
rect 13814 32839 13834 32862
rect 13873 32839 13882 32862
rect 13882 32839 13907 32862
rect 13946 32839 13950 32862
rect 13950 32839 13980 32862
rect 14019 32839 14052 32862
rect 14052 32839 14053 32862
rect 14092 32839 14120 32862
rect 14120 32839 14126 32862
rect 14165 32839 14188 32862
rect 14188 32839 14199 32862
rect 14238 32839 14256 32862
rect 14256 32839 14272 32862
rect 14311 32839 14324 32862
rect 14324 32839 14345 32862
rect 14384 32839 14392 32862
rect 14392 32839 14418 32862
rect 13581 32828 13615 32839
rect 13654 32828 13688 32839
rect 13727 32828 13761 32839
rect 13800 32828 13834 32839
rect 13873 32828 13907 32839
rect 13946 32828 13980 32839
rect 14019 32828 14053 32839
rect 14092 32828 14126 32839
rect 14165 32828 14199 32839
rect 14238 32828 14272 32839
rect 14311 32828 14345 32839
rect 14384 32828 14418 32839
rect 13216 32770 13236 32789
rect 13236 32770 13250 32789
rect 13289 32770 13304 32789
rect 13304 32770 13323 32789
rect 13362 32770 13372 32789
rect 13372 32770 13396 32789
rect 13435 32770 13440 32789
rect 13440 32770 13469 32789
rect 13216 32755 13250 32770
rect 13289 32755 13323 32770
rect 13362 32755 13396 32770
rect 13435 32755 13469 32770
rect 13508 32755 13542 32789
rect 13581 32770 13610 32789
rect 13610 32770 13615 32789
rect 13654 32770 13678 32789
rect 13678 32770 13688 32789
rect 13727 32770 13746 32789
rect 13746 32770 13761 32789
rect 13800 32770 13814 32789
rect 13814 32770 13834 32789
rect 13873 32770 13882 32789
rect 13882 32770 13907 32789
rect 13946 32770 13950 32789
rect 13950 32770 13980 32789
rect 14019 32770 14052 32789
rect 14052 32770 14053 32789
rect 14092 32770 14120 32789
rect 14120 32770 14126 32789
rect 14165 32770 14188 32789
rect 14188 32770 14199 32789
rect 14238 32770 14256 32789
rect 14256 32770 14272 32789
rect 14311 32770 14324 32789
rect 14324 32770 14345 32789
rect 14384 32770 14392 32789
rect 14392 32770 14418 32789
rect 13581 32755 13615 32770
rect 13654 32755 13688 32770
rect 13727 32755 13761 32770
rect 13800 32755 13834 32770
rect 13873 32755 13907 32770
rect 13946 32755 13980 32770
rect 14019 32755 14053 32770
rect 14092 32755 14126 32770
rect 14165 32755 14199 32770
rect 14238 32755 14272 32770
rect 14311 32755 14345 32770
rect 14384 32755 14418 32770
rect 13216 32701 13236 32716
rect 13236 32701 13250 32716
rect 13289 32701 13304 32716
rect 13304 32701 13323 32716
rect 13362 32701 13372 32716
rect 13372 32701 13396 32716
rect 13435 32701 13440 32716
rect 13440 32701 13469 32716
rect 13216 32682 13250 32701
rect 13289 32682 13323 32701
rect 13362 32682 13396 32701
rect 13435 32682 13469 32701
rect 13508 32682 13542 32716
rect 13581 32701 13610 32716
rect 13610 32701 13615 32716
rect 13654 32701 13678 32716
rect 13678 32701 13688 32716
rect 13727 32701 13746 32716
rect 13746 32701 13761 32716
rect 13800 32701 13814 32716
rect 13814 32701 13834 32716
rect 13873 32701 13882 32716
rect 13882 32701 13907 32716
rect 13946 32701 13950 32716
rect 13950 32701 13980 32716
rect 14019 32701 14052 32716
rect 14052 32701 14053 32716
rect 14092 32701 14120 32716
rect 14120 32701 14126 32716
rect 14165 32701 14188 32716
rect 14188 32701 14199 32716
rect 14238 32701 14256 32716
rect 14256 32701 14272 32716
rect 14311 32701 14324 32716
rect 14324 32701 14345 32716
rect 14384 32701 14392 32716
rect 14392 32701 14418 32716
rect 13581 32682 13615 32701
rect 13654 32682 13688 32701
rect 13727 32682 13761 32701
rect 13800 32682 13834 32701
rect 13873 32682 13907 32701
rect 13946 32682 13980 32701
rect 14019 32682 14053 32701
rect 14092 32682 14126 32701
rect 14165 32682 14199 32701
rect 14238 32682 14272 32701
rect 14311 32682 14345 32701
rect 14384 32682 14418 32701
rect 13216 32632 13236 32643
rect 13236 32632 13250 32643
rect 13289 32632 13304 32643
rect 13304 32632 13323 32643
rect 13362 32632 13372 32643
rect 13372 32632 13396 32643
rect 13435 32632 13440 32643
rect 13440 32632 13469 32643
rect 13216 32609 13250 32632
rect 13289 32609 13323 32632
rect 13362 32609 13396 32632
rect 13435 32609 13469 32632
rect 13508 32609 13542 32643
rect 13581 32632 13610 32643
rect 13610 32632 13615 32643
rect 13654 32632 13678 32643
rect 13678 32632 13688 32643
rect 13727 32632 13746 32643
rect 13746 32632 13761 32643
rect 13800 32632 13814 32643
rect 13814 32632 13834 32643
rect 13873 32632 13882 32643
rect 13882 32632 13907 32643
rect 13946 32632 13950 32643
rect 13950 32632 13980 32643
rect 14019 32632 14052 32643
rect 14052 32632 14053 32643
rect 14092 32632 14120 32643
rect 14120 32632 14126 32643
rect 14165 32632 14188 32643
rect 14188 32632 14199 32643
rect 14238 32632 14256 32643
rect 14256 32632 14272 32643
rect 14311 32632 14324 32643
rect 14324 32632 14345 32643
rect 14384 32632 14392 32643
rect 14392 32632 14418 32643
rect 13581 32609 13615 32632
rect 13654 32609 13688 32632
rect 13727 32609 13761 32632
rect 13800 32609 13834 32632
rect 13873 32609 13907 32632
rect 13946 32609 13980 32632
rect 14019 32609 14053 32632
rect 14092 32609 14126 32632
rect 14165 32609 14199 32632
rect 14238 32609 14272 32632
rect 14311 32609 14345 32632
rect 14384 32609 14418 32632
rect 13216 32563 13236 32570
rect 13236 32563 13250 32570
rect 13289 32563 13304 32570
rect 13304 32563 13323 32570
rect 13362 32563 13372 32570
rect 13372 32563 13396 32570
rect 13435 32563 13440 32570
rect 13440 32563 13469 32570
rect 13216 32536 13250 32563
rect 13289 32536 13323 32563
rect 13362 32536 13396 32563
rect 13435 32536 13469 32563
rect 13508 32536 13542 32570
rect 13581 32563 13610 32570
rect 13610 32563 13615 32570
rect 13654 32563 13678 32570
rect 13678 32563 13688 32570
rect 13727 32563 13746 32570
rect 13746 32563 13761 32570
rect 13800 32563 13814 32570
rect 13814 32563 13834 32570
rect 13873 32563 13882 32570
rect 13882 32563 13907 32570
rect 13946 32563 13950 32570
rect 13950 32563 13980 32570
rect 14019 32563 14052 32570
rect 14052 32563 14053 32570
rect 14092 32563 14120 32570
rect 14120 32563 14126 32570
rect 14165 32563 14188 32570
rect 14188 32563 14199 32570
rect 14238 32563 14256 32570
rect 14256 32563 14272 32570
rect 14311 32563 14324 32570
rect 14324 32563 14345 32570
rect 14384 32563 14392 32570
rect 14392 32563 14418 32570
rect 13581 32536 13615 32563
rect 13654 32536 13688 32563
rect 13727 32536 13761 32563
rect 13800 32536 13834 32563
rect 13873 32536 13907 32563
rect 13946 32536 13980 32563
rect 14019 32536 14053 32563
rect 14092 32536 14126 32563
rect 14165 32536 14199 32563
rect 14238 32536 14272 32563
rect 14311 32536 14345 32563
rect 14384 32536 14418 32563
rect 13216 32494 13236 32497
rect 13236 32494 13250 32497
rect 13289 32494 13304 32497
rect 13304 32494 13323 32497
rect 13362 32494 13372 32497
rect 13372 32494 13396 32497
rect 13435 32494 13440 32497
rect 13440 32494 13469 32497
rect 13216 32463 13250 32494
rect 13289 32463 13323 32494
rect 13362 32463 13396 32494
rect 13435 32463 13469 32494
rect 13508 32463 13542 32497
rect 13581 32494 13610 32497
rect 13610 32494 13615 32497
rect 13654 32494 13678 32497
rect 13678 32494 13688 32497
rect 13727 32494 13746 32497
rect 13746 32494 13761 32497
rect 13800 32494 13814 32497
rect 13814 32494 13834 32497
rect 13873 32494 13882 32497
rect 13882 32494 13907 32497
rect 13946 32494 13950 32497
rect 13950 32494 13980 32497
rect 14019 32494 14052 32497
rect 14052 32494 14053 32497
rect 14092 32494 14120 32497
rect 14120 32494 14126 32497
rect 14165 32494 14188 32497
rect 14188 32494 14199 32497
rect 14238 32494 14256 32497
rect 14256 32494 14272 32497
rect 14311 32494 14324 32497
rect 14324 32494 14345 32497
rect 14384 32494 14392 32497
rect 14392 32494 14418 32497
rect 13581 32463 13615 32494
rect 13654 32463 13688 32494
rect 13727 32463 13761 32494
rect 13800 32463 13834 32494
rect 13873 32463 13907 32494
rect 13946 32463 13980 32494
rect 14019 32463 14053 32494
rect 14092 32463 14126 32494
rect 14165 32463 14199 32494
rect 14238 32463 14272 32494
rect 14311 32463 14345 32494
rect 14384 32463 14418 32494
rect 13216 32390 13250 32424
rect 13289 32390 13323 32424
rect 13362 32390 13396 32424
rect 13435 32390 13469 32424
rect 13508 32390 13542 32424
rect 13581 32390 13615 32424
rect 13654 32390 13688 32424
rect 13727 32390 13761 32424
rect 13800 32390 13834 32424
rect 13873 32390 13907 32424
rect 13946 32390 13980 32424
rect 14019 32390 14053 32424
rect 14092 32390 14126 32424
rect 14165 32390 14199 32424
rect 14238 32390 14272 32424
rect 14311 32390 14345 32424
rect 14384 32390 14418 32424
rect 13216 32321 13250 32351
rect 13289 32321 13323 32351
rect 13362 32321 13396 32351
rect 13435 32321 13469 32351
rect 13216 32317 13236 32321
rect 13236 32317 13250 32321
rect 13289 32317 13304 32321
rect 13304 32317 13323 32321
rect 13362 32317 13372 32321
rect 13372 32317 13396 32321
rect 13435 32317 13440 32321
rect 13440 32317 13469 32321
rect 13508 32317 13542 32351
rect 13581 32321 13615 32351
rect 13654 32321 13688 32351
rect 13727 32321 13761 32351
rect 13800 32321 13834 32351
rect 13873 32321 13907 32351
rect 13946 32321 13980 32351
rect 14019 32321 14053 32351
rect 14092 32321 14126 32351
rect 14165 32321 14199 32351
rect 14238 32321 14272 32351
rect 14311 32321 14345 32351
rect 14384 32321 14418 32351
rect 13581 32317 13610 32321
rect 13610 32317 13615 32321
rect 13654 32317 13678 32321
rect 13678 32317 13688 32321
rect 13727 32317 13746 32321
rect 13746 32317 13761 32321
rect 13800 32317 13814 32321
rect 13814 32317 13834 32321
rect 13873 32317 13882 32321
rect 13882 32317 13907 32321
rect 13946 32317 13950 32321
rect 13950 32317 13980 32321
rect 14019 32317 14052 32321
rect 14052 32317 14053 32321
rect 14092 32317 14120 32321
rect 14120 32317 14126 32321
rect 14165 32317 14188 32321
rect 14188 32317 14199 32321
rect 14238 32317 14256 32321
rect 14256 32317 14272 32321
rect 14311 32317 14324 32321
rect 14324 32317 14345 32321
rect 14384 32317 14392 32321
rect 14392 32317 14418 32321
rect 13216 32252 13250 32278
rect 13289 32252 13323 32278
rect 13362 32252 13396 32278
rect 13435 32252 13469 32278
rect 13216 32244 13236 32252
rect 13236 32244 13250 32252
rect 13289 32244 13304 32252
rect 13304 32244 13323 32252
rect 13362 32244 13372 32252
rect 13372 32244 13396 32252
rect 13435 32244 13440 32252
rect 13440 32244 13469 32252
rect 13508 32244 13542 32278
rect 13581 32252 13615 32278
rect 13654 32252 13688 32278
rect 13727 32252 13761 32278
rect 13800 32252 13834 32278
rect 13873 32252 13907 32278
rect 13946 32252 13980 32278
rect 14019 32252 14053 32278
rect 14092 32252 14126 32278
rect 14165 32252 14199 32278
rect 14238 32252 14272 32278
rect 14311 32252 14345 32278
rect 14384 32252 14418 32278
rect 13581 32244 13610 32252
rect 13610 32244 13615 32252
rect 13654 32244 13678 32252
rect 13678 32244 13688 32252
rect 13727 32244 13746 32252
rect 13746 32244 13761 32252
rect 13800 32244 13814 32252
rect 13814 32244 13834 32252
rect 13873 32244 13882 32252
rect 13882 32244 13907 32252
rect 13946 32244 13950 32252
rect 13950 32244 13980 32252
rect 14019 32244 14052 32252
rect 14052 32244 14053 32252
rect 14092 32244 14120 32252
rect 14120 32244 14126 32252
rect 14165 32244 14188 32252
rect 14188 32244 14199 32252
rect 14238 32244 14256 32252
rect 14256 32244 14272 32252
rect 14311 32244 14324 32252
rect 14324 32244 14345 32252
rect 14384 32244 14392 32252
rect 14392 32244 14418 32252
rect 13216 32183 13250 32205
rect 13289 32183 13323 32205
rect 13362 32183 13396 32205
rect 13435 32183 13469 32205
rect 13216 32171 13236 32183
rect 13236 32171 13250 32183
rect 13289 32171 13304 32183
rect 13304 32171 13323 32183
rect 13362 32171 13372 32183
rect 13372 32171 13396 32183
rect 13435 32171 13440 32183
rect 13440 32171 13469 32183
rect 13508 32171 13542 32205
rect 13581 32183 13615 32205
rect 13654 32183 13688 32205
rect 13727 32183 13761 32205
rect 13800 32183 13834 32205
rect 13873 32183 13907 32205
rect 13946 32183 13980 32205
rect 14019 32183 14053 32205
rect 14092 32183 14126 32205
rect 14165 32183 14199 32205
rect 14238 32183 14272 32205
rect 14311 32183 14345 32205
rect 14384 32183 14418 32205
rect 13581 32171 13610 32183
rect 13610 32171 13615 32183
rect 13654 32171 13678 32183
rect 13678 32171 13688 32183
rect 13727 32171 13746 32183
rect 13746 32171 13761 32183
rect 13800 32171 13814 32183
rect 13814 32171 13834 32183
rect 13873 32171 13882 32183
rect 13882 32171 13907 32183
rect 13946 32171 13950 32183
rect 13950 32171 13980 32183
rect 14019 32171 14052 32183
rect 14052 32171 14053 32183
rect 14092 32171 14120 32183
rect 14120 32171 14126 32183
rect 14165 32171 14188 32183
rect 14188 32171 14199 32183
rect 14238 32171 14256 32183
rect 14256 32171 14272 32183
rect 14311 32171 14324 32183
rect 14324 32171 14345 32183
rect 14384 32171 14392 32183
rect 14392 32171 14418 32183
rect 13216 32114 13250 32132
rect 13289 32114 13323 32132
rect 13362 32114 13396 32132
rect 13435 32114 13469 32132
rect 13216 32098 13236 32114
rect 13236 32098 13250 32114
rect 13289 32098 13304 32114
rect 13304 32098 13323 32114
rect 13362 32098 13372 32114
rect 13372 32098 13396 32114
rect 13435 32098 13440 32114
rect 13440 32098 13469 32114
rect 13508 32098 13542 32132
rect 13581 32114 13615 32132
rect 13654 32114 13688 32132
rect 13727 32114 13761 32132
rect 13800 32114 13834 32132
rect 13873 32114 13907 32132
rect 13946 32114 13980 32132
rect 14019 32114 14053 32132
rect 14092 32114 14126 32132
rect 14165 32114 14199 32132
rect 14238 32114 14272 32132
rect 14311 32114 14345 32132
rect 14384 32114 14418 32132
rect 13581 32098 13610 32114
rect 13610 32098 13615 32114
rect 13654 32098 13678 32114
rect 13678 32098 13688 32114
rect 13727 32098 13746 32114
rect 13746 32098 13761 32114
rect 13800 32098 13814 32114
rect 13814 32098 13834 32114
rect 13873 32098 13882 32114
rect 13882 32098 13907 32114
rect 13946 32098 13950 32114
rect 13950 32098 13980 32114
rect 14019 32098 14052 32114
rect 14052 32098 14053 32114
rect 14092 32098 14120 32114
rect 14120 32098 14126 32114
rect 14165 32098 14188 32114
rect 14188 32098 14199 32114
rect 14238 32098 14256 32114
rect 14256 32098 14272 32114
rect 14311 32098 14324 32114
rect 14324 32098 14345 32114
rect 14384 32098 14392 32114
rect 14392 32098 14418 32114
rect 13216 32045 13250 32059
rect 13289 32045 13323 32059
rect 13362 32045 13396 32059
rect 13435 32045 13469 32059
rect 13216 32025 13236 32045
rect 13236 32025 13250 32045
rect 13289 32025 13304 32045
rect 13304 32025 13323 32045
rect 13362 32025 13372 32045
rect 13372 32025 13396 32045
rect 13435 32025 13440 32045
rect 13440 32025 13469 32045
rect 13508 32025 13542 32059
rect 13581 32045 13615 32059
rect 13654 32045 13688 32059
rect 13727 32045 13761 32059
rect 13800 32045 13834 32059
rect 13873 32045 13907 32059
rect 13946 32045 13980 32059
rect 14019 32045 14053 32059
rect 14092 32045 14126 32059
rect 14165 32045 14199 32059
rect 14238 32045 14272 32059
rect 14311 32045 14345 32059
rect 14384 32045 14418 32059
rect 13581 32025 13610 32045
rect 13610 32025 13615 32045
rect 13654 32025 13678 32045
rect 13678 32025 13688 32045
rect 13727 32025 13746 32045
rect 13746 32025 13761 32045
rect 13800 32025 13814 32045
rect 13814 32025 13834 32045
rect 13873 32025 13882 32045
rect 13882 32025 13907 32045
rect 13946 32025 13950 32045
rect 13950 32025 13980 32045
rect 14019 32025 14052 32045
rect 14052 32025 14053 32045
rect 14092 32025 14120 32045
rect 14120 32025 14126 32045
rect 14165 32025 14188 32045
rect 14188 32025 14199 32045
rect 14238 32025 14256 32045
rect 14256 32025 14272 32045
rect 14311 32025 14324 32045
rect 14324 32025 14345 32045
rect 14384 32025 14392 32045
rect 14392 32025 14418 32045
rect 13216 31976 13250 31986
rect 13289 31976 13323 31986
rect 13362 31976 13396 31986
rect 13435 31976 13469 31986
rect 13216 31952 13236 31976
rect 13236 31952 13250 31976
rect 13289 31952 13304 31976
rect 13304 31952 13323 31976
rect 13362 31952 13372 31976
rect 13372 31952 13396 31976
rect 13435 31952 13440 31976
rect 13440 31952 13469 31976
rect 13508 31952 13542 31986
rect 13581 31976 13615 31986
rect 13654 31976 13688 31986
rect 13727 31976 13761 31986
rect 13800 31976 13834 31986
rect 13873 31976 13907 31986
rect 13946 31976 13980 31986
rect 14019 31976 14053 31986
rect 14092 31976 14126 31986
rect 14165 31976 14199 31986
rect 14238 31976 14272 31986
rect 14311 31976 14345 31986
rect 14384 31976 14418 31986
rect 13581 31952 13610 31976
rect 13610 31952 13615 31976
rect 13654 31952 13678 31976
rect 13678 31952 13688 31976
rect 13727 31952 13746 31976
rect 13746 31952 13761 31976
rect 13800 31952 13814 31976
rect 13814 31952 13834 31976
rect 13873 31952 13882 31976
rect 13882 31952 13907 31976
rect 13946 31952 13950 31976
rect 13950 31952 13980 31976
rect 14019 31952 14052 31976
rect 14052 31952 14053 31976
rect 14092 31952 14120 31976
rect 14120 31952 14126 31976
rect 14165 31952 14188 31976
rect 14188 31952 14199 31976
rect 14238 31952 14256 31976
rect 14256 31952 14272 31976
rect 14311 31952 14324 31976
rect 14324 31952 14345 31976
rect 14384 31952 14392 31976
rect 14392 31952 14418 31976
rect 13216 31907 13250 31913
rect 13289 31907 13323 31913
rect 13362 31907 13396 31913
rect 13435 31907 13469 31913
rect 13216 31879 13236 31907
rect 13236 31879 13250 31907
rect 13289 31879 13304 31907
rect 13304 31879 13323 31907
rect 13362 31879 13372 31907
rect 13372 31879 13396 31907
rect 13435 31879 13440 31907
rect 13440 31879 13469 31907
rect 13508 31879 13542 31913
rect 13581 31907 13615 31913
rect 13654 31907 13688 31913
rect 13727 31907 13761 31913
rect 13800 31907 13834 31913
rect 13873 31907 13907 31913
rect 13946 31907 13980 31913
rect 14019 31907 14053 31913
rect 14092 31907 14126 31913
rect 14165 31907 14199 31913
rect 14238 31907 14272 31913
rect 14311 31907 14345 31913
rect 14384 31907 14418 31913
rect 13581 31879 13610 31907
rect 13610 31879 13615 31907
rect 13654 31879 13678 31907
rect 13678 31879 13688 31907
rect 13727 31879 13746 31907
rect 13746 31879 13761 31907
rect 13800 31879 13814 31907
rect 13814 31879 13834 31907
rect 13873 31879 13882 31907
rect 13882 31879 13907 31907
rect 13946 31879 13950 31907
rect 13950 31879 13980 31907
rect 14019 31879 14052 31907
rect 14052 31879 14053 31907
rect 14092 31879 14120 31907
rect 14120 31879 14126 31907
rect 14165 31879 14188 31907
rect 14188 31879 14199 31907
rect 14238 31879 14256 31907
rect 14256 31879 14272 31907
rect 14311 31879 14324 31907
rect 14324 31879 14345 31907
rect 14384 31879 14392 31907
rect 14392 31879 14418 31907
rect 13216 31838 13250 31840
rect 13289 31838 13323 31840
rect 13362 31838 13396 31840
rect 13435 31838 13469 31840
rect 13216 31806 13236 31838
rect 13236 31806 13250 31838
rect 13289 31806 13304 31838
rect 13304 31806 13323 31838
rect 13362 31806 13372 31838
rect 13372 31806 13396 31838
rect 13435 31806 13440 31838
rect 13440 31806 13469 31838
rect 13508 31806 13542 31840
rect 13581 31838 13615 31840
rect 13654 31838 13688 31840
rect 13727 31838 13761 31840
rect 13800 31838 13834 31840
rect 13873 31838 13907 31840
rect 13946 31838 13980 31840
rect 14019 31838 14053 31840
rect 14092 31838 14126 31840
rect 14165 31838 14199 31840
rect 14238 31838 14272 31840
rect 14311 31838 14345 31840
rect 14384 31838 14418 31840
rect 13581 31806 13610 31838
rect 13610 31806 13615 31838
rect 13654 31806 13678 31838
rect 13678 31806 13688 31838
rect 13727 31806 13746 31838
rect 13746 31806 13761 31838
rect 13800 31806 13814 31838
rect 13814 31806 13834 31838
rect 13873 31806 13882 31838
rect 13882 31806 13907 31838
rect 13946 31806 13950 31838
rect 13950 31806 13980 31838
rect 14019 31806 14052 31838
rect 14052 31806 14053 31838
rect 14092 31806 14120 31838
rect 14120 31806 14126 31838
rect 14165 31806 14188 31838
rect 14188 31806 14199 31838
rect 14238 31806 14256 31838
rect 14256 31806 14272 31838
rect 14311 31806 14324 31838
rect 14324 31806 14345 31838
rect 14384 31806 14392 31838
rect 14392 31806 14418 31838
rect 13216 31735 13236 31767
rect 13236 31735 13250 31767
rect 13289 31735 13304 31767
rect 13304 31735 13323 31767
rect 13362 31735 13372 31767
rect 13372 31735 13396 31767
rect 13435 31735 13440 31767
rect 13440 31735 13469 31767
rect 13216 31733 13250 31735
rect 13289 31733 13323 31735
rect 13362 31733 13396 31735
rect 13435 31733 13469 31735
rect 13508 31733 13542 31767
rect 13581 31735 13610 31767
rect 13610 31735 13615 31767
rect 13654 31735 13678 31767
rect 13678 31735 13688 31767
rect 13727 31735 13746 31767
rect 13746 31735 13761 31767
rect 13800 31735 13814 31767
rect 13814 31735 13834 31767
rect 13873 31735 13882 31767
rect 13882 31735 13907 31767
rect 13946 31735 13950 31767
rect 13950 31735 13980 31767
rect 14019 31735 14052 31767
rect 14052 31735 14053 31767
rect 14092 31735 14120 31767
rect 14120 31735 14126 31767
rect 14165 31735 14188 31767
rect 14188 31735 14199 31767
rect 14238 31735 14256 31767
rect 14256 31735 14272 31767
rect 14311 31735 14324 31767
rect 14324 31735 14345 31767
rect 14384 31735 14392 31767
rect 14392 31735 14418 31767
rect 13581 31733 13615 31735
rect 13654 31733 13688 31735
rect 13727 31733 13761 31735
rect 13800 31733 13834 31735
rect 13873 31733 13907 31735
rect 13946 31733 13980 31735
rect 14019 31733 14053 31735
rect 14092 31733 14126 31735
rect 14165 31733 14199 31735
rect 14238 31733 14272 31735
rect 14311 31733 14345 31735
rect 14384 31733 14418 31735
rect 13216 31666 13236 31694
rect 13236 31666 13250 31694
rect 13289 31666 13304 31694
rect 13304 31666 13323 31694
rect 13362 31666 13372 31694
rect 13372 31666 13396 31694
rect 13435 31666 13440 31694
rect 13440 31666 13469 31694
rect 13216 31660 13250 31666
rect 13289 31660 13323 31666
rect 13362 31660 13396 31666
rect 13435 31660 13469 31666
rect 13508 31660 13542 31694
rect 13581 31666 13610 31694
rect 13610 31666 13615 31694
rect 13654 31666 13678 31694
rect 13678 31666 13688 31694
rect 13727 31666 13746 31694
rect 13746 31666 13761 31694
rect 13800 31666 13814 31694
rect 13814 31666 13834 31694
rect 13873 31666 13882 31694
rect 13882 31666 13907 31694
rect 13946 31666 13950 31694
rect 13950 31666 13980 31694
rect 14019 31666 14052 31694
rect 14052 31666 14053 31694
rect 14092 31666 14120 31694
rect 14120 31666 14126 31694
rect 14165 31666 14188 31694
rect 14188 31666 14199 31694
rect 14238 31666 14256 31694
rect 14256 31666 14272 31694
rect 14311 31666 14324 31694
rect 14324 31666 14345 31694
rect 14384 31666 14392 31694
rect 14392 31666 14418 31694
rect 13581 31660 13615 31666
rect 13654 31660 13688 31666
rect 13727 31660 13761 31666
rect 13800 31660 13834 31666
rect 13873 31660 13907 31666
rect 13946 31660 13980 31666
rect 14019 31660 14053 31666
rect 14092 31660 14126 31666
rect 14165 31660 14199 31666
rect 14238 31660 14272 31666
rect 14311 31660 14345 31666
rect 14384 31660 14418 31666
rect 13216 31597 13236 31621
rect 13236 31597 13250 31621
rect 13289 31597 13304 31621
rect 13304 31597 13323 31621
rect 13362 31597 13372 31621
rect 13372 31597 13396 31621
rect 13435 31597 13440 31621
rect 13440 31597 13469 31621
rect 13216 31587 13250 31597
rect 13289 31587 13323 31597
rect 13362 31587 13396 31597
rect 13435 31587 13469 31597
rect 13508 31587 13542 31621
rect 13581 31597 13610 31621
rect 13610 31597 13615 31621
rect 13654 31597 13678 31621
rect 13678 31597 13688 31621
rect 13727 31597 13746 31621
rect 13746 31597 13761 31621
rect 13800 31597 13814 31621
rect 13814 31597 13834 31621
rect 13873 31597 13882 31621
rect 13882 31597 13907 31621
rect 13946 31597 13950 31621
rect 13950 31597 13980 31621
rect 14019 31597 14052 31621
rect 14052 31597 14053 31621
rect 14092 31597 14120 31621
rect 14120 31597 14126 31621
rect 14165 31597 14188 31621
rect 14188 31597 14199 31621
rect 14238 31597 14256 31621
rect 14256 31597 14272 31621
rect 14311 31597 14324 31621
rect 14324 31597 14345 31621
rect 14384 31597 14392 31621
rect 14392 31597 14418 31621
rect 13581 31587 13615 31597
rect 13654 31587 13688 31597
rect 13727 31587 13761 31597
rect 13800 31587 13834 31597
rect 13873 31587 13907 31597
rect 13946 31587 13980 31597
rect 14019 31587 14053 31597
rect 14092 31587 14126 31597
rect 14165 31587 14199 31597
rect 14238 31587 14272 31597
rect 14311 31587 14345 31597
rect 14384 31587 14418 31597
rect 13216 31528 13236 31548
rect 13236 31528 13250 31548
rect 13289 31528 13304 31548
rect 13304 31528 13323 31548
rect 13362 31528 13372 31548
rect 13372 31528 13396 31548
rect 13435 31528 13440 31548
rect 13440 31528 13469 31548
rect 13216 31514 13250 31528
rect 13289 31514 13323 31528
rect 13362 31514 13396 31528
rect 13435 31514 13469 31528
rect 13508 31514 13542 31548
rect 13581 31528 13610 31548
rect 13610 31528 13615 31548
rect 13654 31528 13678 31548
rect 13678 31528 13688 31548
rect 13727 31528 13746 31548
rect 13746 31528 13761 31548
rect 13800 31528 13814 31548
rect 13814 31528 13834 31548
rect 13873 31528 13882 31548
rect 13882 31528 13907 31548
rect 13946 31528 13950 31548
rect 13950 31528 13980 31548
rect 14019 31528 14052 31548
rect 14052 31528 14053 31548
rect 14092 31528 14120 31548
rect 14120 31528 14126 31548
rect 14165 31528 14188 31548
rect 14188 31528 14199 31548
rect 14238 31528 14256 31548
rect 14256 31528 14272 31548
rect 14311 31528 14324 31548
rect 14324 31528 14345 31548
rect 14384 31528 14392 31548
rect 14392 31528 14418 31548
rect 13581 31514 13615 31528
rect 13654 31514 13688 31528
rect 13727 31514 13761 31528
rect 13800 31514 13834 31528
rect 13873 31514 13907 31528
rect 13946 31514 13980 31528
rect 14019 31514 14053 31528
rect 14092 31514 14126 31528
rect 14165 31514 14199 31528
rect 14238 31514 14272 31528
rect 14311 31514 14345 31528
rect 14384 31514 14418 31528
rect 13216 31459 13236 31475
rect 13236 31459 13250 31475
rect 13289 31459 13304 31475
rect 13304 31459 13323 31475
rect 13362 31459 13372 31475
rect 13372 31459 13396 31475
rect 13435 31459 13440 31475
rect 13440 31459 13469 31475
rect 13216 31441 13250 31459
rect 13289 31441 13323 31459
rect 13362 31441 13396 31459
rect 13435 31441 13469 31459
rect 13508 31441 13542 31475
rect 13581 31459 13610 31475
rect 13610 31459 13615 31475
rect 13654 31459 13678 31475
rect 13678 31459 13688 31475
rect 13727 31459 13746 31475
rect 13746 31459 13761 31475
rect 13800 31459 13814 31475
rect 13814 31459 13834 31475
rect 13873 31459 13882 31475
rect 13882 31459 13907 31475
rect 13946 31459 13950 31475
rect 13950 31459 13980 31475
rect 14019 31459 14052 31475
rect 14052 31459 14053 31475
rect 14092 31459 14120 31475
rect 14120 31459 14126 31475
rect 14165 31459 14188 31475
rect 14188 31459 14199 31475
rect 14238 31459 14256 31475
rect 14256 31459 14272 31475
rect 14311 31459 14324 31475
rect 14324 31459 14345 31475
rect 14384 31459 14392 31475
rect 14392 31459 14418 31475
rect 13581 31441 13615 31459
rect 13654 31441 13688 31459
rect 13727 31441 13761 31459
rect 13800 31441 13834 31459
rect 13873 31441 13907 31459
rect 13946 31441 13980 31459
rect 14019 31441 14053 31459
rect 14092 31441 14126 31459
rect 14165 31441 14199 31459
rect 14238 31441 14272 31459
rect 14311 31441 14345 31459
rect 14384 31441 14418 31459
rect 13216 31390 13236 31402
rect 13236 31390 13250 31402
rect 13289 31390 13304 31402
rect 13304 31390 13323 31402
rect 13362 31390 13372 31402
rect 13372 31390 13396 31402
rect 13435 31390 13440 31402
rect 13440 31390 13469 31402
rect 13216 31368 13250 31390
rect 13289 31368 13323 31390
rect 13362 31368 13396 31390
rect 13435 31368 13469 31390
rect 13508 31368 13542 31402
rect 13581 31390 13610 31402
rect 13610 31390 13615 31402
rect 13654 31390 13678 31402
rect 13678 31390 13688 31402
rect 13727 31390 13746 31402
rect 13746 31390 13761 31402
rect 13800 31390 13814 31402
rect 13814 31390 13834 31402
rect 13873 31390 13882 31402
rect 13882 31390 13907 31402
rect 13946 31390 13950 31402
rect 13950 31390 13980 31402
rect 14019 31390 14052 31402
rect 14052 31390 14053 31402
rect 14092 31390 14120 31402
rect 14120 31390 14126 31402
rect 14165 31390 14188 31402
rect 14188 31390 14199 31402
rect 14238 31390 14256 31402
rect 14256 31390 14272 31402
rect 14311 31390 14324 31402
rect 14324 31390 14345 31402
rect 14384 31390 14392 31402
rect 14392 31390 14418 31402
rect 13581 31368 13615 31390
rect 13654 31368 13688 31390
rect 13727 31368 13761 31390
rect 13800 31368 13834 31390
rect 13873 31368 13907 31390
rect 13946 31368 13980 31390
rect 14019 31368 14053 31390
rect 14092 31368 14126 31390
rect 14165 31368 14199 31390
rect 14238 31368 14272 31390
rect 14311 31368 14345 31390
rect 14384 31368 14418 31390
rect 13216 31321 13236 31329
rect 13236 31321 13250 31329
rect 13289 31321 13304 31329
rect 13304 31321 13323 31329
rect 13362 31321 13372 31329
rect 13372 31321 13396 31329
rect 13435 31321 13440 31329
rect 13440 31321 13469 31329
rect 13216 31295 13250 31321
rect 13289 31295 13323 31321
rect 13362 31295 13396 31321
rect 13435 31295 13469 31321
rect 13508 31295 13542 31329
rect 13581 31321 13610 31329
rect 13610 31321 13615 31329
rect 13654 31321 13678 31329
rect 13678 31321 13688 31329
rect 13727 31321 13746 31329
rect 13746 31321 13761 31329
rect 13800 31321 13814 31329
rect 13814 31321 13834 31329
rect 13873 31321 13882 31329
rect 13882 31321 13907 31329
rect 13946 31321 13950 31329
rect 13950 31321 13980 31329
rect 14019 31321 14052 31329
rect 14052 31321 14053 31329
rect 14092 31321 14120 31329
rect 14120 31321 14126 31329
rect 14165 31321 14188 31329
rect 14188 31321 14199 31329
rect 14238 31321 14256 31329
rect 14256 31321 14272 31329
rect 14311 31321 14324 31329
rect 14324 31321 14345 31329
rect 14384 31321 14392 31329
rect 14392 31321 14418 31329
rect 13581 31295 13615 31321
rect 13654 31295 13688 31321
rect 13727 31295 13761 31321
rect 13800 31295 13834 31321
rect 13873 31295 13907 31321
rect 13946 31295 13980 31321
rect 14019 31295 14053 31321
rect 14092 31295 14126 31321
rect 14165 31295 14199 31321
rect 14238 31295 14272 31321
rect 14311 31295 14345 31321
rect 14384 31295 14418 31321
rect 13216 31252 13236 31256
rect 13236 31252 13250 31256
rect 13289 31252 13304 31256
rect 13304 31252 13323 31256
rect 13362 31252 13372 31256
rect 13372 31252 13396 31256
rect 13435 31252 13440 31256
rect 13440 31252 13469 31256
rect 13216 31222 13250 31252
rect 13289 31222 13323 31252
rect 13362 31222 13396 31252
rect 13435 31222 13469 31252
rect 13508 31222 13542 31256
rect 13581 31252 13610 31256
rect 13610 31252 13615 31256
rect 13654 31252 13678 31256
rect 13678 31252 13688 31256
rect 13727 31252 13746 31256
rect 13746 31252 13761 31256
rect 13800 31252 13814 31256
rect 13814 31252 13834 31256
rect 13873 31252 13882 31256
rect 13882 31252 13907 31256
rect 13946 31252 13950 31256
rect 13950 31252 13980 31256
rect 14019 31252 14052 31256
rect 14052 31252 14053 31256
rect 14092 31252 14120 31256
rect 14120 31252 14126 31256
rect 14165 31252 14188 31256
rect 14188 31252 14199 31256
rect 14238 31252 14256 31256
rect 14256 31252 14272 31256
rect 14311 31252 14324 31256
rect 14324 31252 14345 31256
rect 14384 31252 14392 31256
rect 14392 31252 14418 31256
rect 13581 31222 13615 31252
rect 13654 31222 13688 31252
rect 13727 31222 13761 31252
rect 13800 31222 13834 31252
rect 13873 31222 13907 31252
rect 13946 31222 13980 31252
rect 14019 31222 14053 31252
rect 14092 31222 14126 31252
rect 14165 31222 14199 31252
rect 14238 31222 14272 31252
rect 14311 31222 14345 31252
rect 14384 31222 14418 31252
rect 13216 31149 13250 31183
rect 13289 31149 13323 31183
rect 13362 31149 13396 31183
rect 13435 31149 13469 31183
rect 13508 31149 13542 31183
rect 13581 31149 13615 31183
rect 13654 31149 13688 31183
rect 13727 31149 13761 31183
rect 13800 31149 13834 31183
rect 13873 31149 13907 31183
rect 13946 31149 13980 31183
rect 14019 31149 14053 31183
rect 14092 31149 14126 31183
rect 14165 31149 14199 31183
rect 14238 31149 14272 31183
rect 14311 31149 14345 31183
rect 14384 31149 14418 31183
rect 13051 30957 13078 30991
rect 13078 30957 13085 30991
rect 13124 30957 13158 30991
rect 13197 30957 13231 30991
rect 13270 30957 13304 30991
rect 13344 30957 13378 30991
rect 13418 30957 13452 30991
rect 13492 30957 13526 30991
rect 13566 30957 13600 30991
rect 13640 30957 13674 30991
rect 13714 30957 13748 30991
rect 13788 30957 13822 30991
rect 13862 30957 13896 30991
rect 13936 30957 13970 30991
rect 14010 30957 14044 30991
rect 14084 30957 14118 30991
rect 14158 30957 14192 30991
rect 14230 30889 14233 30919
rect 14233 30889 14264 30919
rect 14230 30885 14264 30889
rect 13051 30829 13077 30863
rect 13077 30829 13085 30863
rect 13126 30829 13160 30863
rect 13201 30829 13235 30863
rect 13276 30829 13310 30863
rect 13351 30829 13385 30863
rect 13426 30829 13460 30863
rect 13501 30829 13535 30863
rect 13576 30829 13610 30863
rect 13651 30829 13685 30863
rect 13726 30829 13760 30863
rect 13801 30829 13835 30863
rect 13876 30829 13910 30863
rect 13951 30829 13985 30863
rect 14026 30829 14060 30863
rect 14102 30829 14131 30863
rect 14131 30829 14136 30863
rect 14230 30813 14264 30847
rect 14102 30788 14136 30791
rect 10246 30636 10280 30664
rect 10320 30636 10354 30664
rect 10394 30636 10428 30664
rect 10467 30636 10501 30664
rect 10246 30630 10258 30636
rect 10258 30630 10280 30636
rect 10320 30630 10327 30636
rect 10327 30630 10354 30636
rect 10394 30630 10396 30636
rect 10396 30630 10428 30636
rect 10467 30630 10499 30636
rect 10499 30630 10501 30636
rect 10540 30630 10574 30664
rect 10613 30635 10647 30664
rect 10686 30635 10720 30664
rect 10759 30635 10793 30664
rect 10832 30635 10866 30664
rect 10905 30635 10939 30664
rect 10978 30635 11012 30664
rect 11051 30635 11085 30664
rect 11124 30635 11158 30664
rect 11197 30635 11231 30664
rect 11270 30635 11304 30664
rect 11343 30635 11377 30664
rect 11416 30635 11450 30664
rect 11489 30635 11523 30664
rect 11562 30635 11596 30664
rect 11635 30635 11669 30664
rect 11708 30635 11742 30664
rect 11781 30635 11815 30664
rect 11854 30635 11888 30664
rect 11927 30635 11961 30664
rect 12000 30635 12034 30664
rect 10613 30630 10644 30635
rect 10644 30630 10647 30635
rect 10686 30630 10713 30635
rect 10713 30630 10720 30635
rect 10759 30630 10781 30635
rect 10781 30630 10793 30635
rect 10832 30630 10849 30635
rect 10849 30630 10866 30635
rect 10905 30630 10917 30635
rect 10917 30630 10939 30635
rect 10978 30630 10985 30635
rect 10985 30630 11012 30635
rect 11051 30630 11053 30635
rect 11053 30630 11085 30635
rect 11124 30630 11155 30635
rect 11155 30630 11158 30635
rect 11197 30630 11223 30635
rect 11223 30630 11231 30635
rect 11270 30630 11291 30635
rect 11291 30630 11304 30635
rect 11343 30630 11359 30635
rect 11359 30630 11377 30635
rect 11416 30630 11427 30635
rect 11427 30630 11450 30635
rect 11489 30630 11495 30635
rect 11495 30630 11523 30635
rect 11562 30630 11563 30635
rect 11563 30630 11596 30635
rect 11635 30630 11665 30635
rect 11665 30630 11669 30635
rect 11708 30630 11733 30635
rect 11733 30630 11742 30635
rect 11781 30630 11801 30635
rect 11801 30630 11815 30635
rect 11854 30630 11869 30635
rect 11869 30630 11888 30635
rect 11927 30630 11937 30635
rect 11937 30630 11961 30635
rect 12000 30630 12005 30635
rect 12005 30630 12034 30635
rect 12073 30630 12107 30664
rect 12146 30635 12180 30664
rect 12219 30635 12253 30664
rect 12292 30635 12326 30664
rect 12365 30635 12399 30664
rect 12438 30635 12472 30664
rect 12511 30635 12545 30664
rect 12584 30635 12618 30664
rect 12657 30635 12691 30664
rect 12730 30635 12764 30664
rect 12803 30635 12837 30664
rect 12876 30635 12910 30664
rect 12949 30635 12983 30664
rect 13022 30635 13056 30664
rect 13095 30635 13129 30664
rect 13168 30635 13202 30664
rect 13241 30635 13275 30664
rect 13314 30635 13348 30664
rect 13387 30635 13421 30664
rect 13460 30635 13494 30664
rect 13533 30635 13567 30664
rect 13606 30635 13640 30664
rect 13679 30635 13713 30664
rect 13752 30635 13786 30664
rect 13825 30635 13859 30664
rect 13898 30635 13932 30664
rect 12146 30630 12175 30635
rect 12175 30630 12180 30635
rect 12219 30630 12243 30635
rect 12243 30630 12253 30635
rect 12292 30630 12311 30635
rect 12311 30630 12326 30635
rect 12365 30630 12379 30635
rect 12379 30630 12399 30635
rect 12438 30630 12447 30635
rect 12447 30630 12472 30635
rect 12511 30630 12515 30635
rect 12515 30630 12545 30635
rect 12584 30630 12617 30635
rect 12617 30630 12618 30635
rect 12657 30630 12685 30635
rect 12685 30630 12691 30635
rect 12730 30630 12753 30635
rect 12753 30630 12764 30635
rect 12803 30630 12821 30635
rect 12821 30630 12837 30635
rect 12876 30630 12889 30635
rect 12889 30630 12910 30635
rect 12949 30630 12957 30635
rect 12957 30630 12983 30635
rect 13022 30630 13025 30635
rect 13025 30630 13056 30635
rect 13095 30630 13127 30635
rect 13127 30630 13129 30635
rect 13168 30630 13195 30635
rect 13195 30630 13202 30635
rect 13241 30630 13263 30635
rect 13263 30630 13275 30635
rect 13314 30630 13331 30635
rect 13331 30630 13348 30635
rect 13387 30630 13399 30635
rect 13399 30630 13421 30635
rect 13460 30630 13467 30635
rect 13467 30630 13494 30635
rect 13533 30630 13535 30635
rect 13535 30630 13567 30635
rect 13606 30630 13637 30635
rect 13637 30630 13640 30635
rect 13679 30630 13705 30635
rect 13705 30630 13713 30635
rect 13752 30630 13773 30635
rect 13773 30630 13786 30635
rect 13825 30630 13841 30635
rect 13841 30630 13859 30635
rect 13898 30630 13909 30635
rect 13909 30630 13932 30635
rect 10246 30534 10258 30557
rect 10258 30534 10280 30557
rect 10320 30534 10327 30557
rect 10327 30534 10354 30557
rect 10394 30534 10396 30557
rect 10396 30534 10428 30557
rect 10467 30534 10499 30557
rect 10499 30534 10501 30557
rect 10246 30523 10280 30534
rect 10320 30523 10354 30534
rect 10394 30523 10428 30534
rect 10467 30523 10501 30534
rect 10540 30523 10574 30557
rect 10613 30526 10644 30557
rect 10644 30526 10647 30557
rect 10686 30526 10713 30557
rect 10713 30526 10720 30557
rect 10759 30526 10781 30557
rect 10781 30526 10793 30557
rect 10832 30526 10849 30557
rect 10849 30526 10866 30557
rect 10905 30526 10917 30557
rect 10917 30526 10939 30557
rect 10978 30526 10985 30557
rect 10985 30526 11012 30557
rect 11051 30526 11053 30557
rect 11053 30526 11085 30557
rect 11124 30526 11155 30557
rect 11155 30526 11158 30557
rect 11197 30526 11223 30557
rect 11223 30526 11231 30557
rect 11270 30526 11291 30557
rect 11291 30526 11304 30557
rect 11343 30526 11359 30557
rect 11359 30526 11377 30557
rect 11416 30526 11427 30557
rect 11427 30526 11450 30557
rect 11489 30526 11495 30557
rect 11495 30526 11523 30557
rect 11562 30526 11563 30557
rect 11563 30526 11596 30557
rect 11635 30526 11665 30557
rect 11665 30526 11669 30557
rect 11708 30526 11733 30557
rect 11733 30526 11742 30557
rect 11781 30526 11801 30557
rect 11801 30526 11815 30557
rect 11854 30526 11869 30557
rect 11869 30526 11888 30557
rect 11927 30526 11937 30557
rect 11937 30526 11961 30557
rect 12000 30526 12005 30557
rect 12005 30526 12034 30557
rect 10613 30523 10647 30526
rect 10686 30523 10720 30526
rect 10759 30523 10793 30526
rect 10832 30523 10866 30526
rect 10905 30523 10939 30526
rect 10978 30523 11012 30526
rect 11051 30523 11085 30526
rect 11124 30523 11158 30526
rect 11197 30523 11231 30526
rect 11270 30523 11304 30526
rect 11343 30523 11377 30526
rect 11416 30523 11450 30526
rect 11489 30523 11523 30526
rect 11562 30523 11596 30526
rect 11635 30523 11669 30526
rect 11708 30523 11742 30526
rect 11781 30523 11815 30526
rect 11854 30523 11888 30526
rect 11927 30523 11961 30526
rect 12000 30523 12034 30526
rect 12073 30523 12107 30557
rect 12146 30526 12175 30557
rect 12175 30526 12180 30557
rect 12219 30526 12243 30557
rect 12243 30526 12253 30557
rect 12292 30526 12311 30557
rect 12311 30526 12326 30557
rect 12365 30526 12379 30557
rect 12379 30526 12399 30557
rect 12438 30526 12447 30557
rect 12447 30526 12472 30557
rect 12511 30526 12515 30557
rect 12515 30526 12545 30557
rect 12584 30526 12617 30557
rect 12617 30526 12618 30557
rect 12657 30526 12685 30557
rect 12685 30526 12691 30557
rect 12730 30526 12753 30557
rect 12753 30526 12764 30557
rect 12803 30526 12821 30557
rect 12821 30526 12837 30557
rect 12876 30526 12889 30557
rect 12889 30526 12910 30557
rect 12949 30526 12957 30557
rect 12957 30526 12983 30557
rect 13022 30526 13025 30557
rect 13025 30526 13056 30557
rect 13095 30526 13127 30557
rect 13127 30526 13129 30557
rect 13168 30526 13195 30557
rect 13195 30526 13202 30557
rect 13241 30526 13263 30557
rect 13263 30526 13275 30557
rect 13314 30526 13331 30557
rect 13331 30526 13348 30557
rect 13387 30526 13399 30557
rect 13399 30526 13421 30557
rect 13460 30526 13467 30557
rect 13467 30526 13494 30557
rect 13533 30526 13535 30557
rect 13535 30526 13567 30557
rect 13606 30526 13637 30557
rect 13637 30526 13640 30557
rect 13679 30526 13705 30557
rect 13705 30526 13713 30557
rect 13752 30526 13773 30557
rect 13773 30526 13786 30557
rect 13825 30526 13841 30557
rect 13841 30526 13859 30557
rect 13898 30526 13909 30557
rect 13909 30526 13932 30557
rect 12146 30523 12180 30526
rect 12219 30523 12253 30526
rect 12292 30523 12326 30526
rect 12365 30523 12399 30526
rect 12438 30523 12472 30526
rect 12511 30523 12545 30526
rect 12584 30523 12618 30526
rect 12657 30523 12691 30526
rect 12730 30523 12764 30526
rect 12803 30523 12837 30526
rect 12876 30523 12910 30526
rect 12949 30523 12983 30526
rect 13022 30523 13056 30526
rect 13095 30523 13129 30526
rect 13168 30523 13202 30526
rect 13241 30523 13275 30526
rect 13314 30523 13348 30526
rect 13387 30523 13421 30526
rect 13460 30523 13494 30526
rect 13533 30523 13567 30526
rect 13606 30523 13640 30526
rect 13679 30523 13713 30526
rect 13752 30523 13786 30526
rect 13825 30523 13859 30526
rect 13898 30523 13932 30526
rect 10246 30432 10280 30450
rect 10320 30432 10354 30450
rect 10394 30432 10428 30450
rect 10467 30432 10501 30450
rect 10246 30416 10258 30432
rect 10258 30416 10280 30432
rect 10320 30416 10327 30432
rect 10327 30416 10354 30432
rect 10394 30416 10396 30432
rect 10396 30416 10428 30432
rect 10467 30416 10499 30432
rect 10499 30416 10501 30432
rect 10540 30416 10574 30450
rect 10613 30416 10647 30450
rect 10686 30416 10720 30450
rect 10759 30416 10793 30450
rect 10832 30416 10866 30450
rect 10905 30416 10939 30450
rect 10978 30416 11012 30450
rect 11051 30416 11085 30450
rect 11124 30416 11158 30450
rect 11197 30416 11231 30450
rect 11270 30416 11304 30450
rect 11343 30416 11377 30450
rect 11416 30416 11450 30450
rect 11489 30416 11523 30450
rect 11562 30416 11596 30450
rect 11635 30416 11669 30450
rect 11708 30416 11742 30450
rect 11781 30416 11815 30450
rect 11854 30416 11888 30450
rect 11927 30416 11961 30450
rect 12000 30416 12034 30450
rect 12073 30416 12107 30450
rect 12146 30416 12180 30450
rect 12219 30416 12253 30450
rect 12292 30416 12326 30450
rect 12365 30416 12399 30450
rect 12438 30416 12472 30450
rect 12511 30416 12545 30450
rect 12584 30416 12618 30450
rect 12657 30416 12691 30450
rect 12730 30416 12764 30450
rect 12803 30416 12837 30450
rect 12876 30416 12910 30450
rect 12949 30416 12983 30450
rect 13022 30416 13056 30450
rect 13095 30416 13129 30450
rect 13168 30416 13202 30450
rect 13241 30416 13275 30450
rect 13314 30416 13348 30450
rect 13387 30416 13421 30450
rect 13460 30416 13494 30450
rect 13533 30416 13567 30450
rect 13606 30416 13640 30450
rect 13679 30416 13713 30450
rect 13752 30416 13786 30450
rect 13825 30416 13859 30450
rect 13898 30416 13932 30450
rect 10248 29174 10258 29175
rect 10258 29174 10282 29175
rect 13705 30340 13738 30374
rect 13738 30340 13739 30374
rect 13807 30340 13841 30374
rect 13909 30340 13943 30374
rect 13705 30267 13738 30301
rect 13738 30267 13739 30301
rect 13807 30266 13841 30300
rect 13909 30267 13943 30301
rect 13705 30194 13738 30228
rect 13738 30194 13739 30228
rect 13807 30192 13841 30226
rect 13909 30194 13943 30228
rect 13705 30121 13738 30155
rect 13738 30121 13739 30155
rect 13807 30118 13841 30152
rect 13909 30121 13943 30155
rect 13705 30048 13738 30082
rect 13738 30048 13739 30082
rect 13807 30045 13841 30079
rect 13909 30048 13943 30082
rect 13705 29975 13738 30009
rect 13738 29975 13739 30009
rect 13807 29972 13841 30006
rect 13909 29975 13943 30009
rect 13705 29902 13738 29936
rect 13738 29902 13739 29936
rect 13807 29899 13841 29933
rect 13909 29902 13943 29936
rect 13705 29829 13738 29863
rect 13738 29829 13739 29863
rect 13807 29826 13841 29860
rect 13909 29829 13943 29863
rect 13705 29756 13738 29790
rect 13738 29756 13739 29790
rect 13807 29753 13841 29787
rect 13909 29756 13943 29790
rect 13705 29683 13738 29717
rect 13738 29683 13739 29717
rect 13807 29680 13841 29714
rect 13909 29683 13943 29717
rect 13705 29610 13738 29644
rect 13738 29610 13739 29644
rect 13807 29607 13841 29641
rect 13909 29610 13943 29644
rect 13705 29537 13738 29571
rect 13738 29537 13739 29571
rect 13807 29534 13841 29568
rect 13909 29538 13943 29572
rect 13705 29464 13738 29498
rect 13738 29464 13739 29498
rect 13807 29461 13841 29495
rect 13909 29466 13943 29500
rect 13705 29391 13738 29425
rect 13738 29391 13739 29425
rect 13807 29388 13841 29422
rect 13909 29394 13943 29428
rect 13705 29318 13738 29352
rect 13738 29318 13739 29352
rect 13807 29315 13841 29349
rect 13909 29322 13943 29356
rect 13705 29245 13738 29279
rect 13738 29245 13739 29279
rect 13807 29242 13841 29276
rect 13909 29250 13943 29284
rect 10331 29174 10361 29175
rect 10361 29174 10365 29175
rect 10414 29174 10430 29175
rect 10430 29174 10448 29175
rect 10497 29174 10499 29175
rect 10499 29174 10531 29175
rect 10248 29141 10282 29174
rect 10331 29141 10365 29174
rect 10414 29141 10448 29174
rect 10497 29141 10531 29174
rect 10580 29141 10614 29175
rect 10248 29072 10282 29102
rect 10331 29072 10365 29102
rect 10414 29072 10448 29102
rect 10497 29072 10531 29102
rect 10248 29068 10258 29072
rect 10258 29068 10282 29072
rect 10331 29068 10361 29072
rect 10361 29068 10365 29072
rect 10414 29068 10430 29072
rect 10430 29068 10448 29072
rect 10497 29068 10499 29072
rect 10499 29068 10531 29072
rect 10580 29068 10614 29102
rect 10248 29004 10282 29029
rect 10331 29004 10365 29029
rect 10414 29004 10448 29029
rect 10497 29004 10531 29029
rect 10248 28995 10258 29004
rect 10258 28995 10282 29004
rect 10331 28995 10361 29004
rect 10361 28995 10365 29004
rect 10414 28995 10430 29004
rect 10430 28995 10448 29004
rect 10497 28995 10499 29004
rect 10499 28995 10531 29004
rect 10580 28995 10614 29029
rect 10248 28936 10282 28956
rect 10331 28936 10365 28956
rect 10414 28936 10448 28956
rect 10497 28936 10531 28956
rect 10248 28922 10258 28936
rect 10258 28922 10282 28936
rect 10331 28922 10361 28936
rect 10361 28922 10365 28936
rect 10414 28922 10430 28936
rect 10430 28922 10448 28936
rect 10497 28922 10499 28936
rect 10499 28922 10531 28936
rect 10580 28922 10614 28956
rect 10248 28868 10282 28883
rect 10331 28868 10365 28883
rect 10414 28868 10448 28883
rect 10497 28868 10531 28883
rect 10248 28849 10258 28868
rect 10258 28849 10282 28868
rect 10331 28849 10361 28868
rect 10361 28849 10365 28868
rect 10414 28849 10430 28868
rect 10430 28849 10448 28868
rect 10497 28849 10499 28868
rect 10499 28849 10531 28868
rect 10580 28849 10614 28883
rect 10248 28800 10282 28810
rect 10331 28800 10365 28810
rect 10414 28800 10448 28810
rect 10497 28800 10531 28810
rect 10248 28776 10258 28800
rect 10258 28776 10282 28800
rect 10331 28776 10361 28800
rect 10361 28776 10365 28800
rect 10414 28776 10430 28800
rect 10430 28776 10448 28800
rect 10497 28776 10499 28800
rect 10499 28776 10531 28800
rect 10580 28776 10614 28810
rect 10248 28732 10282 28737
rect 10331 28732 10365 28737
rect 10414 28732 10448 28737
rect 10497 28732 10531 28737
rect 10248 28703 10258 28732
rect 10258 28703 10282 28732
rect 10331 28703 10361 28732
rect 10361 28703 10365 28732
rect 10414 28703 10430 28732
rect 10430 28703 10448 28732
rect 10497 28703 10499 28732
rect 10499 28703 10531 28732
rect 10580 28703 10614 28737
rect 10248 28630 10258 28664
rect 10258 28630 10282 28664
rect 10331 28630 10361 28664
rect 10361 28630 10365 28664
rect 10414 28630 10430 28664
rect 10430 28630 10448 28664
rect 10497 28630 10499 28664
rect 10499 28630 10531 28664
rect 10580 28630 10614 28664
rect 10248 28562 10258 28591
rect 10258 28562 10282 28591
rect 10331 28562 10361 28591
rect 10361 28562 10365 28591
rect 10414 28562 10430 28591
rect 10430 28562 10448 28591
rect 10497 28562 10499 28591
rect 10499 28562 10531 28591
rect 10248 28557 10282 28562
rect 10331 28557 10365 28562
rect 10414 28557 10448 28562
rect 10497 28557 10531 28562
rect 10580 28557 10614 28591
rect 10248 28494 10258 28518
rect 10258 28494 10282 28518
rect 10331 28494 10361 28518
rect 10361 28494 10365 28518
rect 10414 28494 10430 28518
rect 10430 28494 10448 28518
rect 10497 28494 10499 28518
rect 10499 28494 10531 28518
rect 10248 28484 10282 28494
rect 10331 28484 10365 28494
rect 10414 28484 10448 28494
rect 10497 28484 10531 28494
rect 10580 28484 10614 28518
rect 10248 28426 10258 28445
rect 10258 28426 10282 28445
rect 10331 28426 10361 28445
rect 10361 28426 10365 28445
rect 10414 28426 10430 28445
rect 10430 28426 10448 28445
rect 10497 28426 10499 28445
rect 10499 28426 10531 28445
rect 10248 28411 10282 28426
rect 10331 28411 10365 28426
rect 10414 28411 10448 28426
rect 10497 28411 10531 28426
rect 10580 28411 10614 28445
rect 10248 28358 10258 28372
rect 10258 28358 10282 28372
rect 10331 28358 10361 28372
rect 10361 28358 10365 28372
rect 10414 28358 10430 28372
rect 10430 28358 10448 28372
rect 10497 28358 10499 28372
rect 10499 28358 10531 28372
rect 10248 28338 10282 28358
rect 10331 28338 10365 28358
rect 10414 28338 10448 28358
rect 10497 28338 10531 28358
rect 10580 28338 10614 28372
rect 10248 28290 10258 28299
rect 10258 28290 10282 28299
rect 10331 28290 10361 28299
rect 10361 28290 10365 28299
rect 10414 28290 10430 28299
rect 10430 28290 10448 28299
rect 10497 28290 10499 28299
rect 10499 28290 10531 28299
rect 10248 28265 10282 28290
rect 10331 28265 10365 28290
rect 10414 28265 10448 28290
rect 10497 28265 10531 28290
rect 10580 28265 10614 28299
rect 10248 28222 10258 28226
rect 10258 28222 10282 28226
rect 10331 28222 10361 28226
rect 10361 28222 10365 28226
rect 10414 28222 10430 28226
rect 10430 28222 10448 28226
rect 10497 28222 10499 28226
rect 10499 28222 10531 28226
rect 10248 28192 10282 28222
rect 10331 28192 10365 28222
rect 10414 28192 10448 28222
rect 10497 28192 10531 28222
rect 10580 28192 10614 28226
rect 10248 28120 10282 28153
rect 10331 28120 10365 28153
rect 10414 28120 10448 28153
rect 10497 28120 10531 28153
rect 10248 28119 10258 28120
rect 10258 28119 10282 28120
rect 10331 28119 10361 28120
rect 10361 28119 10365 28120
rect 10414 28119 10430 28120
rect 10430 28119 10448 28120
rect 10497 28119 10499 28120
rect 10499 28119 10531 28120
rect 10580 28119 10614 28153
rect 10248 28052 10282 28080
rect 10331 28052 10365 28080
rect 10414 28052 10448 28080
rect 10497 28052 10531 28080
rect 10248 28046 10258 28052
rect 10258 28046 10282 28052
rect 10331 28046 10361 28052
rect 10361 28046 10365 28052
rect 10414 28046 10430 28052
rect 10430 28046 10448 28052
rect 10497 28046 10499 28052
rect 10499 28046 10531 28052
rect 10580 28046 10614 28080
rect 10248 27983 10282 28007
rect 10331 27983 10365 28007
rect 10414 27983 10448 28007
rect 10497 27983 10531 28007
rect 10248 27973 10258 27983
rect 10258 27973 10282 27983
rect 10331 27973 10361 27983
rect 10361 27973 10365 27983
rect 10414 27973 10430 27983
rect 10430 27973 10448 27983
rect 10497 27973 10499 27983
rect 10499 27973 10531 27983
rect 10580 27973 10614 28007
rect 10248 27914 10282 27934
rect 10331 27914 10365 27934
rect 10414 27914 10448 27934
rect 10497 27914 10531 27934
rect 10248 27900 10258 27914
rect 10258 27900 10282 27914
rect 10331 27900 10361 27914
rect 10361 27900 10365 27914
rect 10414 27900 10430 27914
rect 10430 27900 10448 27914
rect 10497 27900 10499 27914
rect 10499 27900 10531 27914
rect 10580 27900 10614 27934
rect 10248 27845 10282 27861
rect 10331 27845 10365 27861
rect 10414 27845 10448 27861
rect 10497 27845 10531 27861
rect 10248 27827 10258 27845
rect 10258 27827 10282 27845
rect 10331 27827 10361 27845
rect 10361 27827 10365 27845
rect 10414 27827 10430 27845
rect 10430 27827 10448 27845
rect 10497 27827 10499 27845
rect 10499 27827 10531 27845
rect 10580 27827 10614 27861
rect 10248 27776 10282 27788
rect 10331 27776 10365 27788
rect 10414 27776 10448 27788
rect 10497 27776 10531 27788
rect 10248 27754 10258 27776
rect 10258 27754 10282 27776
rect 10331 27754 10361 27776
rect 10361 27754 10365 27776
rect 10414 27754 10430 27776
rect 10430 27754 10448 27776
rect 10497 27754 10499 27776
rect 10499 27754 10531 27776
rect 10580 27754 10614 27788
rect 10248 27707 10282 27715
rect 10331 27707 10365 27715
rect 10414 27707 10448 27715
rect 10497 27707 10531 27715
rect 10248 27681 10258 27707
rect 10258 27681 10282 27707
rect 10331 27681 10361 27707
rect 10361 27681 10365 27707
rect 10414 27681 10430 27707
rect 10430 27681 10448 27707
rect 10497 27681 10499 27707
rect 10499 27681 10531 27707
rect 10580 27681 10614 27715
rect 10248 27638 10282 27642
rect 10331 27638 10365 27642
rect 10414 27638 10448 27642
rect 10497 27638 10531 27642
rect 10248 27608 10258 27638
rect 10258 27608 10282 27638
rect 10331 27608 10361 27638
rect 10361 27608 10365 27638
rect 10414 27608 10430 27638
rect 10430 27608 10448 27638
rect 10497 27608 10499 27638
rect 10499 27608 10531 27638
rect 10580 27608 10614 27642
rect 10248 27535 10258 27568
rect 10258 27535 10282 27568
rect 10331 27535 10361 27568
rect 10361 27535 10365 27568
rect 10414 27535 10430 27568
rect 10430 27535 10448 27568
rect 10497 27535 10499 27568
rect 10499 27535 10531 27568
rect 10248 27534 10282 27535
rect 10331 27534 10365 27535
rect 10414 27534 10448 27535
rect 10497 27534 10531 27535
rect 10580 27534 10614 27568
rect 10248 27466 10258 27494
rect 10258 27466 10282 27494
rect 10331 27466 10361 27494
rect 10361 27466 10365 27494
rect 10414 27466 10430 27494
rect 10430 27466 10448 27494
rect 10497 27466 10499 27494
rect 10499 27466 10531 27494
rect 10248 27460 10282 27466
rect 10331 27460 10365 27466
rect 10414 27460 10448 27466
rect 10497 27460 10531 27466
rect 10580 27460 10614 27494
rect 10248 27397 10258 27420
rect 10258 27397 10282 27420
rect 10331 27397 10361 27420
rect 10361 27397 10365 27420
rect 10414 27397 10430 27420
rect 10430 27397 10448 27420
rect 10497 27397 10499 27420
rect 10499 27397 10531 27420
rect 10248 27386 10282 27397
rect 10331 27386 10365 27397
rect 10414 27386 10448 27397
rect 10497 27386 10531 27397
rect 10580 27386 10614 27420
rect 10248 27328 10258 27346
rect 10258 27328 10282 27346
rect 10331 27328 10361 27346
rect 10361 27328 10365 27346
rect 10414 27328 10430 27346
rect 10430 27328 10448 27346
rect 10497 27328 10499 27346
rect 10499 27328 10531 27346
rect 10248 27312 10282 27328
rect 10331 27312 10365 27328
rect 10414 27312 10448 27328
rect 10497 27312 10531 27328
rect 10580 27312 10614 27346
rect 10248 27259 10258 27272
rect 10258 27259 10282 27272
rect 10331 27259 10361 27272
rect 10361 27259 10365 27272
rect 10414 27259 10430 27272
rect 10430 27259 10448 27272
rect 10497 27259 10499 27272
rect 10499 27259 10531 27272
rect 10248 27238 10282 27259
rect 10331 27238 10365 27259
rect 10414 27238 10448 27259
rect 10497 27238 10531 27259
rect 10580 27238 10614 27272
rect 10248 27190 10258 27198
rect 10258 27190 10282 27198
rect 10331 27190 10361 27198
rect 10361 27190 10365 27198
rect 10414 27190 10430 27198
rect 10430 27190 10448 27198
rect 10497 27190 10499 27198
rect 10499 27190 10531 27198
rect 10248 27164 10282 27190
rect 10331 27164 10365 27190
rect 10414 27164 10448 27190
rect 10497 27164 10531 27190
rect 10580 27164 10614 27198
rect 10248 27121 10258 27124
rect 10258 27121 10282 27124
rect 10331 27121 10361 27124
rect 10361 27121 10365 27124
rect 10414 27121 10430 27124
rect 10430 27121 10448 27124
rect 10497 27121 10499 27124
rect 10499 27121 10531 27124
rect 10248 27090 10282 27121
rect 10331 27090 10365 27121
rect 10414 27090 10448 27121
rect 10497 27090 10531 27121
rect 10580 27090 10614 27124
rect 10248 27016 10282 27050
rect 10331 27016 10365 27050
rect 10414 27016 10448 27050
rect 10497 27016 10531 27050
rect 10580 27016 10614 27050
rect 10248 26942 10282 26976
rect 10331 26942 10365 26976
rect 10414 26942 10448 26976
rect 10497 26942 10531 26976
rect 10580 26942 10614 26976
rect 13705 29172 13738 29206
rect 13738 29172 13739 29206
rect 13807 29169 13841 29203
rect 13909 29178 13943 29212
rect 13705 29099 13738 29133
rect 13738 29099 13739 29133
rect 13807 29096 13841 29130
rect 13909 29106 13943 29140
rect 13705 29026 13738 29060
rect 13738 29026 13739 29060
rect 13807 29023 13841 29057
rect 13909 29034 13943 29068
rect 13705 28972 13739 28987
rect 13807 28972 13841 28984
rect 13705 28953 13738 28972
rect 13738 28953 13739 28972
rect 13807 28950 13840 28972
rect 13840 28950 13841 28972
rect 13909 28962 13943 28996
rect 13705 28903 13739 28914
rect 13807 28903 13841 28911
rect 13705 28880 13738 28903
rect 13738 28880 13739 28903
rect 13807 28877 13840 28903
rect 13840 28877 13841 28903
rect 13909 28890 13943 28924
rect 13705 28834 13739 28841
rect 13807 28834 13841 28838
rect 13705 28807 13738 28834
rect 13738 28807 13739 28834
rect 13807 28804 13840 28834
rect 13840 28804 13841 28834
rect 13909 28818 13943 28852
rect 13705 28765 13739 28769
rect 13705 28735 13738 28765
rect 13738 28735 13739 28765
rect 13807 28731 13840 28765
rect 13840 28731 13841 28765
rect 13909 28746 13943 28780
rect 13705 28696 13739 28697
rect 13705 28663 13738 28696
rect 13738 28663 13739 28696
rect 13807 28662 13840 28692
rect 13840 28662 13841 28692
rect 13909 28674 13943 28708
rect 13807 28658 13841 28662
rect 13705 28593 13738 28625
rect 13738 28593 13739 28625
rect 13807 28593 13840 28619
rect 13840 28593 13841 28619
rect 13909 28602 13943 28636
rect 13705 28591 13739 28593
rect 13807 28585 13841 28593
rect 13705 28524 13738 28553
rect 13738 28524 13739 28553
rect 13807 28524 13840 28546
rect 13840 28524 13841 28546
rect 13909 28530 13943 28564
rect 13705 28519 13739 28524
rect 13807 28512 13841 28524
rect 13705 28455 13738 28481
rect 13738 28455 13739 28481
rect 13807 28455 13840 28473
rect 13840 28455 13841 28473
rect 13909 28458 13943 28492
rect 13705 28447 13739 28455
rect 13807 28439 13841 28455
rect 13705 28386 13738 28409
rect 13738 28386 13739 28409
rect 13807 28386 13840 28400
rect 13840 28386 13841 28400
rect 13909 28386 13943 28420
rect 13705 28375 13739 28386
rect 13807 28366 13841 28386
rect 13705 28317 13738 28337
rect 13738 28317 13739 28337
rect 13807 28317 13840 28327
rect 13840 28317 13841 28327
rect 13705 28303 13739 28317
rect 13807 28293 13841 28317
rect 13909 28314 13943 28348
rect 13705 28248 13738 28265
rect 13738 28248 13739 28265
rect 13807 28248 13840 28254
rect 13840 28248 13841 28254
rect 13705 28231 13739 28248
rect 13807 28220 13841 28248
rect 13909 28242 13943 28276
rect 13705 28179 13738 28193
rect 13738 28179 13739 28193
rect 13807 28179 13840 28181
rect 13840 28179 13841 28181
rect 13705 28159 13739 28179
rect 13807 28147 13841 28179
rect 13909 28170 13943 28204
rect 13705 28110 13738 28121
rect 13738 28110 13739 28121
rect 13705 28087 13739 28110
rect 13807 28075 13841 28108
rect 13909 28098 13943 28132
rect 13705 28041 13738 28049
rect 13738 28041 13739 28049
rect 13807 28074 13840 28075
rect 13840 28074 13841 28075
rect 13705 28015 13739 28041
rect 13807 28006 13841 28035
rect 13909 28026 13943 28060
rect 13705 27972 13738 27977
rect 13738 27972 13739 27977
rect 13807 28001 13840 28006
rect 13840 28001 13841 28006
rect 13705 27943 13739 27972
rect 13807 27937 13841 27962
rect 13909 27954 13943 27988
rect 13705 27903 13738 27905
rect 13738 27903 13739 27905
rect 13807 27928 13840 27937
rect 13840 27928 13841 27937
rect 13705 27871 13739 27903
rect 13807 27868 13841 27889
rect 13909 27882 13943 27916
rect 13807 27855 13840 27868
rect 13840 27855 13841 27868
rect 13705 27799 13739 27833
rect 13807 27799 13841 27816
rect 13909 27810 13943 27844
rect 13807 27782 13840 27799
rect 13840 27782 13841 27799
rect 13705 27730 13739 27761
rect 13807 27730 13841 27743
rect 13909 27738 13943 27772
rect 13705 27727 13738 27730
rect 13738 27727 13739 27730
rect 13807 27709 13840 27730
rect 13840 27709 13841 27730
rect 13705 27661 13739 27689
rect 13807 27661 13841 27670
rect 13909 27666 13943 27700
rect 13705 27655 13738 27661
rect 13738 27655 13739 27661
rect 13807 27636 13840 27661
rect 13840 27636 13841 27661
rect 13705 27592 13739 27617
rect 13807 27592 13841 27597
rect 13909 27594 13943 27628
rect 13705 27583 13738 27592
rect 13738 27583 13739 27592
rect 13807 27563 13840 27592
rect 13840 27563 13841 27592
rect 13705 27523 13739 27545
rect 13807 27523 13841 27524
rect 13705 27511 13738 27523
rect 13738 27511 13739 27523
rect 13807 27490 13840 27523
rect 13840 27490 13841 27523
rect 13909 27522 13943 27556
rect 13705 27454 13739 27473
rect 13705 27439 13738 27454
rect 13738 27439 13739 27454
rect 13807 27420 13840 27451
rect 13840 27420 13841 27451
rect 13909 27450 13943 27484
rect 13807 27417 13841 27420
rect 13705 27385 13739 27401
rect 13705 27367 13738 27385
rect 13738 27367 13739 27385
rect 13807 27351 13840 27378
rect 13840 27351 13841 27378
rect 13909 27378 13943 27412
rect 13807 27344 13841 27351
rect 13705 27316 13739 27329
rect 13705 27295 13738 27316
rect 13738 27295 13739 27316
rect 13807 27282 13840 27305
rect 13840 27282 13841 27305
rect 13909 27306 13943 27340
rect 13807 27271 13841 27282
rect 13705 27247 13739 27257
rect 13705 27223 13738 27247
rect 13738 27223 13739 27247
rect 13807 27213 13840 27232
rect 13840 27213 13841 27232
rect 13909 27234 13943 27268
rect 13807 27198 13841 27213
rect 13705 27178 13739 27185
rect 13705 27151 13738 27178
rect 13738 27151 13739 27178
rect 13807 27144 13840 27159
rect 13840 27144 13841 27159
rect 13909 27162 13943 27196
rect 13807 27125 13841 27144
rect 13705 27109 13739 27113
rect 13705 27079 13738 27109
rect 13738 27079 13739 27109
rect 13807 27075 13840 27086
rect 13840 27075 13841 27086
rect 13909 27090 13943 27124
rect 13807 27052 13841 27075
rect 13705 27040 13739 27041
rect 13705 27007 13738 27040
rect 13738 27007 13739 27040
rect 13807 27006 13840 27013
rect 13840 27006 13841 27013
rect 13909 27018 13943 27052
rect 13807 26979 13841 27006
rect 10659 26938 10693 26969
rect 10731 26938 10765 26969
rect 10803 26938 10837 26969
rect 10875 26938 10909 26969
rect 10947 26938 10981 26969
rect 11019 26938 11053 26969
rect 11091 26938 11125 26969
rect 11163 26938 11197 26969
rect 11235 26938 11269 26969
rect 11307 26938 11341 26969
rect 11379 26938 11413 26969
rect 11451 26938 11485 26969
rect 11523 26938 11557 26969
rect 11595 26938 11629 26969
rect 11667 26938 11701 26969
rect 11739 26938 11773 26969
rect 11811 26938 11845 26969
rect 11883 26938 11917 26969
rect 11955 26938 11989 26969
rect 12027 26938 12061 26969
rect 12099 26938 12133 26969
rect 12172 26938 12206 26969
rect 12245 26938 12279 26969
rect 12318 26938 12352 26969
rect 12391 26938 12425 26969
rect 12464 26938 12498 26969
rect 12537 26938 12571 26969
rect 12610 26938 12644 26969
rect 12683 26938 12717 26969
rect 12756 26938 12790 26969
rect 12829 26938 12863 26969
rect 12902 26938 12936 26969
rect 12975 26938 13009 26969
rect 13048 26938 13082 26969
rect 13121 26938 13155 26969
rect 13194 26938 13228 26969
rect 13267 26938 13301 26969
rect 13340 26938 13374 26969
rect 13413 26938 13447 26969
rect 13486 26938 13520 26969
rect 13559 26938 13593 26969
rect 13632 26938 13666 26969
rect 10659 26935 10670 26938
rect 10670 26935 10693 26938
rect 10731 26935 10739 26938
rect 10739 26935 10765 26938
rect 10803 26935 10808 26938
rect 10808 26935 10837 26938
rect 10875 26935 10877 26938
rect 10877 26935 10909 26938
rect 10947 26935 10980 26938
rect 10980 26935 10981 26938
rect 11019 26935 11049 26938
rect 11049 26935 11053 26938
rect 11091 26935 11118 26938
rect 11118 26935 11125 26938
rect 11163 26935 11187 26938
rect 11187 26935 11197 26938
rect 11235 26935 11256 26938
rect 11256 26935 11269 26938
rect 11307 26935 11325 26938
rect 11325 26935 11341 26938
rect 11379 26935 11393 26938
rect 11393 26935 11413 26938
rect 11451 26935 11461 26938
rect 11461 26935 11485 26938
rect 11523 26935 11529 26938
rect 11529 26935 11557 26938
rect 11595 26935 11597 26938
rect 11597 26935 11629 26938
rect 11667 26935 11699 26938
rect 11699 26935 11701 26938
rect 11739 26935 11767 26938
rect 11767 26935 11773 26938
rect 11811 26935 11835 26938
rect 11835 26935 11845 26938
rect 11883 26935 11903 26938
rect 11903 26935 11917 26938
rect 11955 26935 11971 26938
rect 11971 26935 11989 26938
rect 12027 26935 12039 26938
rect 12039 26935 12061 26938
rect 12099 26935 12107 26938
rect 12107 26935 12133 26938
rect 12172 26935 12175 26938
rect 12175 26935 12206 26938
rect 12245 26935 12277 26938
rect 12277 26935 12279 26938
rect 12318 26935 12345 26938
rect 12345 26935 12352 26938
rect 12391 26935 12413 26938
rect 12413 26935 12425 26938
rect 12464 26935 12481 26938
rect 12481 26935 12498 26938
rect 12537 26935 12549 26938
rect 12549 26935 12571 26938
rect 12610 26935 12617 26938
rect 12617 26935 12644 26938
rect 12683 26935 12685 26938
rect 12685 26935 12717 26938
rect 12756 26935 12787 26938
rect 12787 26935 12790 26938
rect 12829 26935 12855 26938
rect 12855 26935 12863 26938
rect 12902 26935 12923 26938
rect 12923 26935 12936 26938
rect 12975 26935 12991 26938
rect 12991 26935 13009 26938
rect 13048 26935 13059 26938
rect 13059 26935 13082 26938
rect 13121 26935 13127 26938
rect 13127 26935 13155 26938
rect 13194 26935 13195 26938
rect 13195 26935 13228 26938
rect 13267 26935 13297 26938
rect 13297 26935 13301 26938
rect 13340 26935 13365 26938
rect 13365 26935 13374 26938
rect 13413 26935 13433 26938
rect 13433 26935 13447 26938
rect 13486 26935 13501 26938
rect 13501 26935 13520 26938
rect 13559 26935 13569 26938
rect 13569 26935 13593 26938
rect 13632 26935 13637 26938
rect 13637 26935 13666 26938
rect 13705 26935 13739 26969
rect 13909 26946 13943 26980
rect 13807 26938 13841 26940
rect 13807 26906 13841 26938
rect 10248 26868 10282 26902
rect 10331 26868 10365 26902
rect 10414 26868 10448 26902
rect 10497 26868 10531 26902
rect 10580 26868 10614 26902
rect 13909 26874 13943 26908
rect 10659 26866 10693 26867
rect 10732 26866 10766 26867
rect 10805 26866 10839 26867
rect 10878 26866 10912 26867
rect 10951 26866 10985 26867
rect 11024 26866 11058 26867
rect 11097 26866 11131 26867
rect 11170 26866 11204 26867
rect 11243 26866 11277 26867
rect 11316 26866 11350 26867
rect 11389 26866 11423 26867
rect 11462 26866 11496 26867
rect 11535 26866 11569 26867
rect 11608 26866 11642 26867
rect 11681 26866 11715 26867
rect 11754 26866 11788 26867
rect 11827 26866 11861 26867
rect 11900 26866 11934 26867
rect 11973 26866 12007 26867
rect 12046 26866 12080 26867
rect 12119 26866 12153 26867
rect 12192 26866 12226 26867
rect 12265 26866 12299 26867
rect 12338 26866 12372 26867
rect 12411 26866 12445 26867
rect 12484 26866 12518 26867
rect 12557 26866 12591 26867
rect 12630 26866 12664 26867
rect 12703 26866 12737 26867
rect 12776 26866 12810 26867
rect 12849 26866 12883 26867
rect 12922 26866 12956 26867
rect 12995 26866 13029 26867
rect 13068 26866 13102 26867
rect 13141 26866 13175 26867
rect 13215 26866 13249 26867
rect 13289 26866 13323 26867
rect 13363 26866 13397 26867
rect 13437 26866 13471 26867
rect 13511 26866 13545 26867
rect 13585 26866 13619 26867
rect 13659 26866 13693 26867
rect 13733 26866 13767 26867
rect 13807 26866 13841 26867
rect 10659 26833 10670 26866
rect 10670 26833 10693 26866
rect 10732 26833 10739 26866
rect 10739 26833 10766 26866
rect 10805 26833 10808 26866
rect 10808 26833 10839 26866
rect 10878 26833 10911 26866
rect 10911 26833 10912 26866
rect 10951 26833 10980 26866
rect 10980 26833 10985 26866
rect 11024 26833 11049 26866
rect 11049 26833 11058 26866
rect 11097 26833 11118 26866
rect 11118 26833 11131 26866
rect 11170 26833 11187 26866
rect 11187 26833 11204 26866
rect 11243 26833 11256 26866
rect 11256 26833 11277 26866
rect 11316 26833 11325 26866
rect 11325 26833 11350 26866
rect 11389 26833 11393 26866
rect 11393 26833 11423 26866
rect 11462 26833 11495 26866
rect 11495 26833 11496 26866
rect 11535 26833 11563 26866
rect 11563 26833 11569 26866
rect 11608 26833 11631 26866
rect 11631 26833 11642 26866
rect 11681 26833 11699 26866
rect 11699 26833 11715 26866
rect 11754 26833 11767 26866
rect 11767 26833 11788 26866
rect 11827 26833 11835 26866
rect 11835 26833 11861 26866
rect 11900 26833 11903 26866
rect 11903 26833 11934 26866
rect 11973 26833 12005 26866
rect 12005 26833 12007 26866
rect 12046 26833 12073 26866
rect 12073 26833 12080 26866
rect 12119 26833 12141 26866
rect 12141 26833 12153 26866
rect 12192 26833 12209 26866
rect 12209 26833 12226 26866
rect 12265 26833 12277 26866
rect 12277 26833 12299 26866
rect 12338 26833 12345 26866
rect 12345 26833 12372 26866
rect 12411 26833 12413 26866
rect 12413 26833 12445 26866
rect 12484 26833 12515 26866
rect 12515 26833 12518 26866
rect 12557 26833 12583 26866
rect 12583 26833 12591 26866
rect 12630 26833 12651 26866
rect 12651 26833 12664 26866
rect 12703 26833 12719 26866
rect 12719 26833 12737 26866
rect 12776 26833 12787 26866
rect 12787 26833 12810 26866
rect 12849 26833 12855 26866
rect 12855 26833 12883 26866
rect 12922 26833 12923 26866
rect 12923 26833 12956 26866
rect 12995 26833 13025 26866
rect 13025 26833 13029 26866
rect 13068 26833 13093 26866
rect 13093 26833 13102 26866
rect 13141 26833 13161 26866
rect 13161 26833 13175 26866
rect 13215 26833 13229 26866
rect 13229 26833 13249 26866
rect 13289 26833 13297 26866
rect 13297 26833 13323 26866
rect 13363 26833 13365 26866
rect 13365 26833 13397 26866
rect 13437 26833 13467 26866
rect 13467 26833 13471 26866
rect 13511 26833 13535 26866
rect 13535 26833 13545 26866
rect 13585 26833 13603 26866
rect 13603 26833 13619 26866
rect 13659 26833 13671 26866
rect 13671 26833 13693 26866
rect 13733 26833 13739 26866
rect 13739 26833 13767 26866
rect 13807 26833 13841 26866
rect 10248 26794 10282 26828
rect 10331 26794 10365 26828
rect 10414 26794 10448 26828
rect 10497 26794 10531 26828
rect 10580 26794 10614 26828
rect 13909 26802 13943 26836
rect 10659 26760 10670 26765
rect 10670 26760 10693 26765
rect 10731 26760 10739 26765
rect 10739 26760 10765 26765
rect 10803 26760 10808 26765
rect 10808 26760 10837 26765
rect 10875 26760 10877 26765
rect 10877 26760 10909 26765
rect 10947 26760 10980 26765
rect 10980 26760 10981 26765
rect 11019 26760 11049 26765
rect 11049 26760 11053 26765
rect 11091 26760 11118 26765
rect 11118 26760 11125 26765
rect 11163 26760 11187 26765
rect 11187 26760 11197 26765
rect 11235 26760 11256 26765
rect 11256 26760 11269 26765
rect 11307 26760 11325 26765
rect 11325 26760 11341 26765
rect 11379 26760 11393 26765
rect 11393 26760 11413 26765
rect 11451 26760 11461 26765
rect 11461 26760 11485 26765
rect 11523 26760 11529 26765
rect 11529 26760 11557 26765
rect 11595 26760 11597 26765
rect 11597 26760 11629 26765
rect 11667 26760 11699 26765
rect 11699 26760 11701 26765
rect 11739 26760 11767 26765
rect 11767 26760 11773 26765
rect 11811 26760 11835 26765
rect 11835 26760 11845 26765
rect 11883 26760 11903 26765
rect 11903 26760 11917 26765
rect 11955 26760 11971 26765
rect 11971 26760 11989 26765
rect 12027 26760 12039 26765
rect 12039 26760 12061 26765
rect 12099 26760 12107 26765
rect 12107 26760 12133 26765
rect 12171 26760 12175 26765
rect 12175 26760 12205 26765
rect 12243 26760 12277 26765
rect 12315 26760 12345 26765
rect 12345 26760 12349 26765
rect 12387 26760 12413 26765
rect 12413 26760 12421 26765
rect 12459 26760 12481 26765
rect 12481 26760 12493 26765
rect 12531 26760 12549 26765
rect 12549 26760 12565 26765
rect 12603 26760 12617 26765
rect 12617 26760 12637 26765
rect 12675 26760 12685 26765
rect 12685 26760 12709 26765
rect 12747 26760 12753 26765
rect 12753 26760 12781 26765
rect 12819 26760 12821 26765
rect 12821 26760 12853 26765
rect 12891 26760 12923 26765
rect 12923 26760 12925 26765
rect 12963 26760 12991 26765
rect 12991 26760 12997 26765
rect 13035 26760 13059 26765
rect 13059 26760 13069 26765
rect 13108 26760 13127 26765
rect 13127 26760 13142 26765
rect 13181 26760 13195 26765
rect 13195 26760 13215 26765
rect 13254 26760 13263 26765
rect 13263 26760 13288 26765
rect 13327 26760 13331 26765
rect 13331 26760 13361 26765
rect 13400 26760 13433 26765
rect 13433 26760 13434 26765
rect 13473 26760 13501 26765
rect 13501 26760 13507 26765
rect 13546 26760 13569 26765
rect 13569 26760 13580 26765
rect 13619 26760 13637 26765
rect 13637 26760 13653 26765
rect 13692 26760 13705 26765
rect 13705 26760 13726 26765
rect 13765 26760 13773 26765
rect 13773 26760 13799 26765
rect 13838 26760 13841 26765
rect 13841 26760 13872 26765
rect 10248 26720 10282 26754
rect 10331 26720 10365 26754
rect 10414 26720 10448 26754
rect 10497 26720 10531 26754
rect 10580 26720 10614 26754
rect 10659 26731 10693 26760
rect 10731 26731 10765 26760
rect 10803 26731 10837 26760
rect 10875 26731 10909 26760
rect 10947 26731 10981 26760
rect 11019 26731 11053 26760
rect 11091 26731 11125 26760
rect 11163 26731 11197 26760
rect 11235 26731 11269 26760
rect 11307 26731 11341 26760
rect 11379 26731 11413 26760
rect 11451 26731 11485 26760
rect 11523 26731 11557 26760
rect 11595 26731 11629 26760
rect 11667 26731 11701 26760
rect 11739 26731 11773 26760
rect 11811 26731 11845 26760
rect 11883 26731 11917 26760
rect 11955 26731 11989 26760
rect 12027 26731 12061 26760
rect 12099 26731 12133 26760
rect 12171 26731 12205 26760
rect 12243 26731 12277 26760
rect 12315 26731 12349 26760
rect 12387 26731 12421 26760
rect 12459 26731 12493 26760
rect 12531 26731 12565 26760
rect 12603 26731 12637 26760
rect 12675 26731 12709 26760
rect 12747 26731 12781 26760
rect 12819 26731 12853 26760
rect 12891 26731 12925 26760
rect 12963 26731 12997 26760
rect 13035 26731 13069 26760
rect 13108 26731 13142 26760
rect 13181 26731 13215 26760
rect 13254 26731 13288 26760
rect 13327 26731 13361 26760
rect 13400 26731 13434 26760
rect 13473 26731 13507 26760
rect 13546 26731 13580 26760
rect 13619 26731 13653 26760
rect 13692 26731 13726 26760
rect 13765 26731 13799 26760
rect 13838 26731 13872 26760
rect 14102 30757 14136 30788
rect 14230 30741 14264 30775
rect 14102 30685 14136 30719
rect 14230 30669 14264 30703
rect 14102 30613 14136 30647
rect 14230 30597 14264 30631
rect 14102 30541 14136 30575
rect 14230 30525 14264 30559
rect 14102 30469 14136 30503
rect 14230 30453 14264 30487
rect 14102 30397 14136 30431
rect 14230 30381 14264 30415
rect 14102 30325 14136 30359
rect 14230 30309 14264 30343
rect 14102 30253 14136 30287
rect 14230 30237 14264 30271
rect 14102 30181 14136 30215
rect 14230 30165 14264 30199
rect 14102 30109 14136 30143
rect 14230 30093 14264 30127
rect 14102 30037 14136 30071
rect 14230 30021 14264 30055
rect 14102 29965 14136 29999
rect 14230 29949 14264 29983
rect 14102 29892 14136 29926
rect 14230 29877 14264 29911
rect 14102 29819 14136 29853
rect 14230 29805 14264 29839
rect 14102 29746 14136 29780
rect 14230 29733 14264 29767
rect 14102 29673 14136 29707
rect 14230 29661 14264 29695
rect 14102 29600 14136 29634
rect 14230 29589 14264 29623
rect 14102 29527 14136 29561
rect 14230 29517 14264 29551
rect 14102 29454 14136 29488
rect 14230 29445 14264 29479
rect 14102 29381 14136 29415
rect 14230 29373 14264 29407
rect 14102 29308 14136 29342
rect 14230 29301 14264 29335
rect 14102 29235 14136 29269
rect 14230 29229 14264 29263
rect 14102 29162 14136 29196
rect 14230 29157 14264 29191
rect 14102 29089 14136 29123
rect 14230 29085 14264 29119
rect 14102 29016 14136 29050
rect 14230 29013 14264 29047
rect 14102 28943 14136 28977
rect 14230 28941 14264 28975
rect 14102 28870 14136 28904
rect 14230 28869 14264 28903
rect 14102 28797 14136 28831
rect 14230 28797 14264 28831
rect 14102 28724 14136 28758
rect 14230 28725 14264 28759
rect 14102 28651 14136 28685
rect 14230 28653 14264 28687
rect 14102 28578 14136 28612
rect 14230 28581 14264 28615
rect 14102 28505 14136 28539
rect 14230 28509 14264 28543
rect 14102 28432 14136 28466
rect 14230 28437 14264 28471
rect 14102 28359 14136 28393
rect 14230 28365 14264 28399
rect 14102 28286 14136 28320
rect 14230 28293 14264 28327
rect 14102 28213 14136 28247
rect 14230 28221 14264 28255
rect 14102 28140 14136 28174
rect 14230 28149 14264 28183
rect 14102 28067 14136 28101
rect 14230 28077 14264 28111
rect 14102 27994 14136 28028
rect 14230 28005 14264 28039
rect 14102 27921 14136 27955
rect 14230 27933 14264 27967
rect 14102 27848 14136 27882
rect 14230 27861 14264 27895
rect 14102 27775 14136 27809
rect 14230 27789 14264 27823
rect 14102 27702 14136 27736
rect 14230 27717 14264 27751
rect 14102 27629 14136 27663
rect 14230 27645 14264 27679
rect 14102 27556 14136 27590
rect 14230 27573 14264 27607
rect 14102 27483 14136 27517
rect 14230 27500 14264 27534
rect 14102 27410 14136 27444
rect 14230 27427 14264 27461
rect 14102 27337 14136 27371
rect 14230 27354 14264 27388
rect 14102 27264 14136 27298
rect 14230 27281 14264 27315
rect 14102 27191 14136 27225
rect 14230 27208 14264 27242
rect 14102 27118 14136 27152
rect 14230 27135 14264 27169
rect 14102 27045 14136 27079
rect 14230 27062 14264 27096
rect 14102 26972 14136 27006
rect 14230 26989 14264 27023
rect 14102 26899 14136 26933
rect 14230 26916 14264 26950
rect 14102 26826 14136 26860
rect 14230 26843 14264 26877
rect 14102 26753 14136 26787
rect 14230 26770 14264 26804
rect 14102 26680 14136 26714
rect 14230 26697 14264 26731
rect 14102 26607 14136 26641
rect 14230 26624 14264 26658
rect 9765 26534 9799 26568
rect 9838 26534 9872 26568
rect 9911 26534 9945 26568
rect 9984 26534 10018 26568
rect 10057 26534 10091 26568
rect 10130 26534 10164 26568
rect 10203 26534 10237 26568
rect 10276 26534 10310 26568
rect 10349 26534 10383 26568
rect 10422 26534 10456 26568
rect 10495 26534 10529 26568
rect 10568 26534 10602 26568
rect 10641 26534 10675 26568
rect 10714 26534 10748 26568
rect 10787 26534 10821 26568
rect 10860 26534 10894 26568
rect 10933 26534 10967 26568
rect 11006 26534 11040 26568
rect 11078 26534 11112 26568
rect 11150 26534 11184 26568
rect 11222 26534 11256 26568
rect 11294 26534 11328 26568
rect 11366 26534 11400 26568
rect 11438 26534 11472 26568
rect 11510 26534 11544 26568
rect 11582 26534 11616 26568
rect 11654 26534 11688 26568
rect 11726 26534 11760 26568
rect 11798 26534 11832 26568
rect 11870 26534 11904 26568
rect 11942 26534 11976 26568
rect 12014 26534 12048 26568
rect 12086 26534 12120 26568
rect 12158 26534 12192 26568
rect 12230 26534 12264 26568
rect 12302 26534 12336 26568
rect 12374 26534 12408 26568
rect 12446 26534 12480 26568
rect 12518 26534 12552 26568
rect 12590 26534 12624 26568
rect 12662 26534 12696 26568
rect 12734 26534 12768 26568
rect 12806 26534 12840 26568
rect 12878 26534 12912 26568
rect 12950 26534 12984 26568
rect 13022 26534 13056 26568
rect 13094 26534 13128 26568
rect 13166 26534 13200 26568
rect 13238 26534 13272 26568
rect 13310 26534 13344 26568
rect 13382 26534 13416 26568
rect 13454 26534 13488 26568
rect 13526 26534 13560 26568
rect 13598 26534 13632 26568
rect 13670 26534 13704 26568
rect 13742 26534 13776 26568
rect 13814 26534 13848 26568
rect 13886 26534 13920 26568
rect 13958 26534 13992 26568
rect 14030 26534 14064 26568
rect 14102 26538 14136 26568
rect 14230 26551 14264 26585
rect 14102 26534 14136 26538
rect 14230 26478 14264 26512
rect 9765 26406 9799 26440
rect 9838 26406 9872 26440
rect 9910 26406 9944 26440
rect 9982 26406 10016 26440
rect 10054 26406 10088 26440
rect 10126 26406 10160 26440
rect 10198 26406 10232 26440
rect 10270 26406 10304 26440
rect 10342 26406 10376 26440
rect 10414 26406 10448 26440
rect 10486 26406 10520 26440
rect 10558 26406 10592 26440
rect 10630 26406 10664 26440
rect 10702 26406 10736 26440
rect 10774 26406 10808 26440
rect 10846 26406 10880 26440
rect 10918 26406 10952 26440
rect 10990 26406 11024 26440
rect 11062 26406 11096 26440
rect 11134 26406 11168 26440
rect 11206 26406 11240 26440
rect 11278 26406 11312 26440
rect 11350 26406 11384 26440
rect 11422 26406 11456 26440
rect 11494 26406 11528 26440
rect 11566 26406 11600 26440
rect 11638 26406 11672 26440
rect 11710 26406 11744 26440
rect 11782 26406 11816 26440
rect 11854 26406 11888 26440
rect 11926 26406 11960 26440
rect 11998 26406 12032 26440
rect 12070 26406 12104 26440
rect 12142 26406 12176 26440
rect 12214 26406 12248 26440
rect 12286 26406 12320 26440
rect 12358 26406 12392 26440
rect 12430 26406 12464 26440
rect 12502 26406 12536 26440
rect 12574 26406 12608 26440
rect 12646 26406 12680 26440
rect 12718 26406 12752 26440
rect 12790 26406 12824 26440
rect 12862 26406 12896 26440
rect 12934 26406 12968 26440
rect 13006 26406 13040 26440
rect 13078 26406 13112 26440
rect 13150 26406 13184 26440
rect 13222 26406 13256 26440
rect 13294 26406 13328 26440
rect 13366 26406 13400 26440
rect 13438 26406 13472 26440
rect 13510 26406 13544 26440
rect 13582 26406 13616 26440
rect 13654 26406 13688 26440
rect 13726 26406 13760 26440
rect 13798 26406 13832 26440
rect 13870 26406 13904 26440
rect 13942 26406 13976 26440
rect 14014 26406 14048 26440
rect 14086 26436 14120 26440
rect 14086 26406 14111 26436
rect 14111 26406 14120 26436
rect 14158 26406 14192 26440
rect 9909 26214 9943 26248
rect 9981 26214 10015 26248
rect 10053 26214 10087 26248
rect 10125 26214 10159 26248
rect 10197 26214 10231 26248
rect 10269 26214 10303 26248
rect 10341 26214 10375 26248
rect 10413 26214 10447 26248
rect 10485 26214 10519 26248
rect 10557 26214 10591 26248
rect 10629 26214 10663 26248
rect 10701 26214 10735 26248
rect 10773 26214 10807 26248
rect 10845 26214 10879 26248
rect 10917 26214 10951 26248
rect 10989 26214 11023 26248
rect 11061 26214 11095 26248
rect 11133 26214 11167 26248
rect 11205 26214 11239 26248
rect 11277 26214 11311 26248
rect 11349 26214 11383 26248
rect 11421 26214 11455 26248
rect 11493 26214 11527 26248
rect 11565 26214 11599 26248
rect 11637 26214 11671 26248
rect 11709 26214 11743 26248
rect 11781 26214 11815 26248
rect 11853 26214 11887 26248
rect 11925 26214 11959 26248
rect 11997 26214 12031 26248
rect 12069 26214 12103 26248
rect 12141 26214 12175 26248
rect 12213 26214 12247 26248
rect 12285 26214 12319 26248
rect 12357 26214 12391 26248
rect 12429 26214 12463 26248
rect 12501 26214 12535 26248
rect 12573 26214 12607 26248
rect 12645 26214 12679 26248
rect 12717 26214 12751 26248
rect 12789 26214 12823 26248
rect 12861 26214 12895 26248
rect 12933 26214 12967 26248
rect 13005 26214 13039 26248
rect 13077 26214 13111 26248
rect 13149 26214 13183 26248
rect 13221 26214 13255 26248
rect 13293 26214 13327 26248
rect 13365 26214 13399 26248
rect 13437 26214 13471 26248
rect 13509 26214 13543 26248
rect 13581 26214 13615 26248
rect 13653 26214 13687 26248
rect 13756 26214 13790 26248
rect 13828 26214 13862 26248
rect 13900 26214 13934 26248
rect 13972 26214 14006 26248
rect 14044 26214 14078 26248
rect 14116 26214 14150 26248
rect 9909 26165 9911 26174
rect 9911 26165 9943 26174
rect 9981 26165 10014 26174
rect 10014 26165 10015 26174
rect 10053 26165 10083 26174
rect 10083 26165 10087 26174
rect 10125 26165 10152 26174
rect 10152 26165 10159 26174
rect 10197 26165 10221 26174
rect 10221 26165 10231 26174
rect 10269 26165 10290 26174
rect 10290 26165 10303 26174
rect 10341 26165 10359 26174
rect 10359 26165 10375 26174
rect 10413 26165 10428 26174
rect 10428 26165 10447 26174
rect 10485 26165 10497 26174
rect 10497 26165 10519 26174
rect 10557 26165 10566 26174
rect 10566 26165 10591 26174
rect 10629 26165 10635 26174
rect 10635 26165 10663 26174
rect 10701 26165 10704 26174
rect 10704 26165 10735 26174
rect 9909 26140 9943 26165
rect 9981 26140 10015 26165
rect 10053 26140 10087 26165
rect 10125 26140 10159 26165
rect 10197 26140 10231 26165
rect 10269 26140 10303 26165
rect 10341 26140 10375 26165
rect 10413 26140 10447 26165
rect 10485 26140 10519 26165
rect 10557 26140 10591 26165
rect 10629 26140 10663 26165
rect 10701 26140 10735 26165
rect 10773 26140 10807 26174
rect 10845 26165 10875 26174
rect 10875 26165 10879 26174
rect 10917 26165 10943 26174
rect 10943 26165 10951 26174
rect 10989 26165 11011 26174
rect 11011 26165 11023 26174
rect 11061 26165 11079 26174
rect 11079 26165 11095 26174
rect 11133 26165 11147 26174
rect 11147 26165 11167 26174
rect 11205 26165 11215 26174
rect 11215 26165 11239 26174
rect 11277 26165 11283 26174
rect 11283 26165 11311 26174
rect 11349 26165 11351 26174
rect 11351 26165 11383 26174
rect 11421 26165 11453 26174
rect 11453 26165 11455 26174
rect 11493 26165 11521 26174
rect 11521 26165 11527 26174
rect 11565 26165 11589 26174
rect 11589 26165 11599 26174
rect 11637 26165 11657 26174
rect 11657 26165 11671 26174
rect 11709 26165 11725 26174
rect 11725 26165 11743 26174
rect 11781 26165 11793 26174
rect 11793 26165 11815 26174
rect 11853 26165 11861 26174
rect 11861 26165 11887 26174
rect 11925 26165 11929 26174
rect 11929 26165 11959 26174
rect 10845 26140 10879 26165
rect 10917 26140 10951 26165
rect 10989 26140 11023 26165
rect 11061 26140 11095 26165
rect 11133 26140 11167 26165
rect 11205 26140 11239 26165
rect 11277 26140 11311 26165
rect 11349 26140 11383 26165
rect 11421 26140 11455 26165
rect 11493 26140 11527 26165
rect 11565 26140 11599 26165
rect 11637 26140 11671 26165
rect 11709 26140 11743 26165
rect 11781 26140 11815 26165
rect 11853 26140 11887 26165
rect 11925 26140 11959 26165
rect 11997 26140 12031 26174
rect 12069 26165 12099 26174
rect 12099 26165 12103 26174
rect 12141 26165 12167 26174
rect 12167 26165 12175 26174
rect 12213 26165 12235 26174
rect 12235 26165 12247 26174
rect 12285 26165 12303 26174
rect 12303 26165 12319 26174
rect 12357 26165 12371 26174
rect 12371 26165 12391 26174
rect 12429 26165 12439 26174
rect 12439 26165 12463 26174
rect 12501 26165 12507 26174
rect 12507 26165 12535 26174
rect 12573 26165 12575 26174
rect 12575 26165 12607 26174
rect 12645 26165 12677 26174
rect 12677 26165 12679 26174
rect 12717 26165 12745 26174
rect 12745 26165 12751 26174
rect 12789 26165 12813 26174
rect 12813 26165 12823 26174
rect 12861 26165 12881 26174
rect 12881 26165 12895 26174
rect 12933 26165 12949 26174
rect 12949 26165 12967 26174
rect 13005 26165 13017 26174
rect 13017 26165 13039 26174
rect 13077 26165 13085 26174
rect 13085 26165 13111 26174
rect 13149 26165 13153 26174
rect 13153 26165 13183 26174
rect 12069 26140 12103 26165
rect 12141 26140 12175 26165
rect 12213 26140 12247 26165
rect 12285 26140 12319 26165
rect 12357 26140 12391 26165
rect 12429 26140 12463 26165
rect 12501 26140 12535 26165
rect 12573 26140 12607 26165
rect 12645 26140 12679 26165
rect 12717 26140 12751 26165
rect 12789 26140 12823 26165
rect 12861 26140 12895 26165
rect 12933 26140 12967 26165
rect 13005 26140 13039 26165
rect 13077 26140 13111 26165
rect 13149 26140 13183 26165
rect 13221 26140 13255 26174
rect 13293 26165 13323 26174
rect 13323 26165 13327 26174
rect 13365 26165 13391 26174
rect 13391 26165 13399 26174
rect 13437 26165 13459 26174
rect 13459 26165 13471 26174
rect 13509 26165 13527 26174
rect 13527 26165 13543 26174
rect 13581 26165 13595 26174
rect 13595 26165 13615 26174
rect 13653 26165 13663 26174
rect 13663 26165 13687 26174
rect 13756 26165 13765 26175
rect 13765 26165 13790 26175
rect 13828 26165 13833 26175
rect 13833 26165 13862 26175
rect 13900 26165 13901 26175
rect 13901 26165 13934 26175
rect 13972 26165 14003 26175
rect 14003 26165 14006 26175
rect 14044 26165 14071 26175
rect 14071 26165 14078 26175
rect 14116 26165 14139 26175
rect 14139 26165 14150 26175
rect 13293 26140 13327 26165
rect 13365 26140 13399 26165
rect 13437 26140 13471 26165
rect 13509 26140 13543 26165
rect 13581 26140 13615 26165
rect 13653 26140 13687 26165
rect 13756 26141 13790 26165
rect 13828 26141 13862 26165
rect 13900 26141 13934 26165
rect 13972 26141 14006 26165
rect 14044 26141 14078 26165
rect 14116 26141 14150 26165
rect 9909 26095 9911 26100
rect 9911 26095 9943 26100
rect 9981 26095 10014 26100
rect 10014 26095 10015 26100
rect 10053 26095 10083 26100
rect 10083 26095 10087 26100
rect 10125 26095 10152 26100
rect 10152 26095 10159 26100
rect 10197 26095 10221 26100
rect 10221 26095 10231 26100
rect 10269 26095 10290 26100
rect 10290 26095 10303 26100
rect 10341 26095 10359 26100
rect 10359 26095 10375 26100
rect 10413 26095 10428 26100
rect 10428 26095 10447 26100
rect 10485 26095 10497 26100
rect 10497 26095 10519 26100
rect 10557 26095 10566 26100
rect 10566 26095 10591 26100
rect 10629 26095 10635 26100
rect 10635 26095 10663 26100
rect 10701 26095 10704 26100
rect 10704 26095 10735 26100
rect 9909 26066 9943 26095
rect 9981 26066 10015 26095
rect 10053 26066 10087 26095
rect 10125 26066 10159 26095
rect 10197 26066 10231 26095
rect 10269 26066 10303 26095
rect 10341 26066 10375 26095
rect 10413 26066 10447 26095
rect 10485 26066 10519 26095
rect 10557 26066 10591 26095
rect 10629 26066 10663 26095
rect 10701 26066 10735 26095
rect 10773 26066 10807 26100
rect 10845 26095 10875 26100
rect 10875 26095 10879 26100
rect 10917 26095 10943 26100
rect 10943 26095 10951 26100
rect 10989 26095 11011 26100
rect 11011 26095 11023 26100
rect 11061 26095 11079 26100
rect 11079 26095 11095 26100
rect 11133 26095 11147 26100
rect 11147 26095 11167 26100
rect 11205 26095 11215 26100
rect 11215 26095 11239 26100
rect 11277 26095 11283 26100
rect 11283 26095 11311 26100
rect 11349 26095 11351 26100
rect 11351 26095 11383 26100
rect 11421 26095 11453 26100
rect 11453 26095 11455 26100
rect 11493 26095 11521 26100
rect 11521 26095 11527 26100
rect 11565 26095 11589 26100
rect 11589 26095 11599 26100
rect 11637 26095 11657 26100
rect 11657 26095 11671 26100
rect 11709 26095 11725 26100
rect 11725 26095 11743 26100
rect 11781 26095 11793 26100
rect 11793 26095 11815 26100
rect 11853 26095 11861 26100
rect 11861 26095 11887 26100
rect 11925 26095 11929 26100
rect 11929 26095 11959 26100
rect 10845 26066 10879 26095
rect 10917 26066 10951 26095
rect 10989 26066 11023 26095
rect 11061 26066 11095 26095
rect 11133 26066 11167 26095
rect 11205 26066 11239 26095
rect 11277 26066 11311 26095
rect 11349 26066 11383 26095
rect 11421 26066 11455 26095
rect 11493 26066 11527 26095
rect 11565 26066 11599 26095
rect 11637 26066 11671 26095
rect 11709 26066 11743 26095
rect 11781 26066 11815 26095
rect 11853 26066 11887 26095
rect 11925 26066 11959 26095
rect 11997 26066 12031 26100
rect 12069 26095 12099 26100
rect 12099 26095 12103 26100
rect 12141 26095 12167 26100
rect 12167 26095 12175 26100
rect 12213 26095 12235 26100
rect 12235 26095 12247 26100
rect 12285 26095 12303 26100
rect 12303 26095 12319 26100
rect 12357 26095 12371 26100
rect 12371 26095 12391 26100
rect 12429 26095 12439 26100
rect 12439 26095 12463 26100
rect 12501 26095 12507 26100
rect 12507 26095 12535 26100
rect 12573 26095 12575 26100
rect 12575 26095 12607 26100
rect 12645 26095 12677 26100
rect 12677 26095 12679 26100
rect 12717 26095 12745 26100
rect 12745 26095 12751 26100
rect 12789 26095 12813 26100
rect 12813 26095 12823 26100
rect 12861 26095 12881 26100
rect 12881 26095 12895 26100
rect 12933 26095 12949 26100
rect 12949 26095 12967 26100
rect 13005 26095 13017 26100
rect 13017 26095 13039 26100
rect 13077 26095 13085 26100
rect 13085 26095 13111 26100
rect 13149 26095 13153 26100
rect 13153 26095 13183 26100
rect 12069 26066 12103 26095
rect 12141 26066 12175 26095
rect 12213 26066 12247 26095
rect 12285 26066 12319 26095
rect 12357 26066 12391 26095
rect 12429 26066 12463 26095
rect 12501 26066 12535 26095
rect 12573 26066 12607 26095
rect 12645 26066 12679 26095
rect 12717 26066 12751 26095
rect 12789 26066 12823 26095
rect 12861 26066 12895 26095
rect 12933 26066 12967 26095
rect 13005 26066 13039 26095
rect 13077 26066 13111 26095
rect 13149 26066 13183 26095
rect 13221 26066 13255 26100
rect 13293 26095 13323 26100
rect 13323 26095 13327 26100
rect 13365 26095 13391 26100
rect 13391 26095 13399 26100
rect 13437 26095 13459 26100
rect 13459 26095 13471 26100
rect 13509 26095 13527 26100
rect 13527 26095 13543 26100
rect 13581 26095 13595 26100
rect 13595 26095 13615 26100
rect 13653 26095 13663 26100
rect 13663 26095 13687 26100
rect 13756 26095 13765 26102
rect 13765 26095 13790 26102
rect 13828 26095 13833 26102
rect 13833 26095 13862 26102
rect 13900 26095 13901 26102
rect 13901 26095 13934 26102
rect 13972 26095 14003 26102
rect 14003 26095 14006 26102
rect 14044 26095 14071 26102
rect 14071 26095 14078 26102
rect 14116 26095 14139 26102
rect 14139 26095 14150 26102
rect 13293 26066 13327 26095
rect 13365 26066 13399 26095
rect 13437 26066 13471 26095
rect 13509 26066 13543 26095
rect 13581 26066 13615 26095
rect 13653 26066 13687 26095
rect 13756 26068 13790 26095
rect 13828 26068 13862 26095
rect 13900 26068 13934 26095
rect 13972 26068 14006 26095
rect 14044 26068 14078 26095
rect 14116 26068 14150 26095
rect 9909 26025 9911 26026
rect 9911 26025 9943 26026
rect 9981 26025 10014 26026
rect 10014 26025 10015 26026
rect 10053 26025 10083 26026
rect 10083 26025 10087 26026
rect 10125 26025 10152 26026
rect 10152 26025 10159 26026
rect 10197 26025 10221 26026
rect 10221 26025 10231 26026
rect 10269 26025 10290 26026
rect 10290 26025 10303 26026
rect 10341 26025 10359 26026
rect 10359 26025 10375 26026
rect 10413 26025 10428 26026
rect 10428 26025 10447 26026
rect 10485 26025 10497 26026
rect 10497 26025 10519 26026
rect 10557 26025 10566 26026
rect 10566 26025 10591 26026
rect 10629 26025 10635 26026
rect 10635 26025 10663 26026
rect 10701 26025 10704 26026
rect 10704 26025 10735 26026
rect 9909 25992 9943 26025
rect 9981 25992 10015 26025
rect 10053 25992 10087 26025
rect 10125 25992 10159 26025
rect 10197 25992 10231 26025
rect 10269 25992 10303 26025
rect 10341 25992 10375 26025
rect 10413 25992 10447 26025
rect 10485 25992 10519 26025
rect 10557 25992 10591 26025
rect 10629 25992 10663 26025
rect 10701 25992 10735 26025
rect 10773 25992 10807 26026
rect 10845 26025 10875 26026
rect 10875 26025 10879 26026
rect 10917 26025 10943 26026
rect 10943 26025 10951 26026
rect 10989 26025 11011 26026
rect 11011 26025 11023 26026
rect 11061 26025 11079 26026
rect 11079 26025 11095 26026
rect 11133 26025 11147 26026
rect 11147 26025 11167 26026
rect 11205 26025 11215 26026
rect 11215 26025 11239 26026
rect 11277 26025 11283 26026
rect 11283 26025 11311 26026
rect 11349 26025 11351 26026
rect 11351 26025 11383 26026
rect 11421 26025 11453 26026
rect 11453 26025 11455 26026
rect 11493 26025 11521 26026
rect 11521 26025 11527 26026
rect 11565 26025 11589 26026
rect 11589 26025 11599 26026
rect 11637 26025 11657 26026
rect 11657 26025 11671 26026
rect 11709 26025 11725 26026
rect 11725 26025 11743 26026
rect 11781 26025 11793 26026
rect 11793 26025 11815 26026
rect 11853 26025 11861 26026
rect 11861 26025 11887 26026
rect 11925 26025 11929 26026
rect 11929 26025 11959 26026
rect 10845 25992 10879 26025
rect 10917 25992 10951 26025
rect 10989 25992 11023 26025
rect 11061 25992 11095 26025
rect 11133 25992 11167 26025
rect 11205 25992 11239 26025
rect 11277 25992 11311 26025
rect 11349 25992 11383 26025
rect 11421 25992 11455 26025
rect 11493 25992 11527 26025
rect 11565 25992 11599 26025
rect 11637 25992 11671 26025
rect 11709 25992 11743 26025
rect 11781 25992 11815 26025
rect 11853 25992 11887 26025
rect 11925 25992 11959 26025
rect 11997 25992 12031 26026
rect 12069 26025 12099 26026
rect 12099 26025 12103 26026
rect 12141 26025 12167 26026
rect 12167 26025 12175 26026
rect 12213 26025 12235 26026
rect 12235 26025 12247 26026
rect 12285 26025 12303 26026
rect 12303 26025 12319 26026
rect 12357 26025 12371 26026
rect 12371 26025 12391 26026
rect 12429 26025 12439 26026
rect 12439 26025 12463 26026
rect 12501 26025 12507 26026
rect 12507 26025 12535 26026
rect 12573 26025 12575 26026
rect 12575 26025 12607 26026
rect 12645 26025 12677 26026
rect 12677 26025 12679 26026
rect 12717 26025 12745 26026
rect 12745 26025 12751 26026
rect 12789 26025 12813 26026
rect 12813 26025 12823 26026
rect 12861 26025 12881 26026
rect 12881 26025 12895 26026
rect 12933 26025 12949 26026
rect 12949 26025 12967 26026
rect 13005 26025 13017 26026
rect 13017 26025 13039 26026
rect 13077 26025 13085 26026
rect 13085 26025 13111 26026
rect 13149 26025 13153 26026
rect 13153 26025 13183 26026
rect 12069 25992 12103 26025
rect 12141 25992 12175 26025
rect 12213 25992 12247 26025
rect 12285 25992 12319 26025
rect 12357 25992 12391 26025
rect 12429 25992 12463 26025
rect 12501 25992 12535 26025
rect 12573 25992 12607 26025
rect 12645 25992 12679 26025
rect 12717 25992 12751 26025
rect 12789 25992 12823 26025
rect 12861 25992 12895 26025
rect 12933 25992 12967 26025
rect 13005 25992 13039 26025
rect 13077 25992 13111 26025
rect 13149 25992 13183 26025
rect 13221 25992 13255 26026
rect 13293 26025 13323 26026
rect 13323 26025 13327 26026
rect 13365 26025 13391 26026
rect 13391 26025 13399 26026
rect 13437 26025 13459 26026
rect 13459 26025 13471 26026
rect 13509 26025 13527 26026
rect 13527 26025 13543 26026
rect 13581 26025 13595 26026
rect 13595 26025 13615 26026
rect 13653 26025 13663 26026
rect 13663 26025 13687 26026
rect 13756 26025 13765 26029
rect 13765 26025 13790 26029
rect 13828 26025 13833 26029
rect 13833 26025 13862 26029
rect 13900 26025 13901 26029
rect 13901 26025 13934 26029
rect 13972 26025 14003 26029
rect 14003 26025 14006 26029
rect 14044 26025 14071 26029
rect 14071 26025 14078 26029
rect 14116 26025 14139 26029
rect 14139 26025 14150 26029
rect 13293 25992 13327 26025
rect 13365 25992 13399 26025
rect 13437 25992 13471 26025
rect 13509 25992 13543 26025
rect 13581 25992 13615 26025
rect 13653 25992 13687 26025
rect 13756 25995 13790 26025
rect 13828 25995 13862 26025
rect 13900 25995 13934 26025
rect 13972 25995 14006 26025
rect 14044 25995 14078 26025
rect 14116 25995 14150 26025
rect 9909 25919 9943 25953
rect 9981 25919 10015 25953
rect 10053 25919 10087 25953
rect 10125 25919 10159 25953
rect 10197 25919 10231 25953
rect 10269 25919 10303 25953
rect 10341 25919 10375 25953
rect 10413 25919 10447 25953
rect 10485 25919 10519 25953
rect 10557 25919 10591 25953
rect 10629 25919 10663 25953
rect 10701 25919 10735 25953
rect 10773 25919 10807 25953
rect 10845 25919 10879 25953
rect 10917 25919 10951 25953
rect 10989 25919 11023 25953
rect 11061 25919 11095 25953
rect 11133 25919 11167 25953
rect 11205 25919 11239 25953
rect 11277 25919 11311 25953
rect 11349 25919 11383 25953
rect 11421 25919 11455 25953
rect 11493 25919 11527 25953
rect 11565 25919 11599 25953
rect 11637 25919 11671 25953
rect 11709 25919 11743 25953
rect 11781 25919 11815 25953
rect 11853 25919 11887 25953
rect 11925 25919 11959 25953
rect 11997 25919 12031 25953
rect 12069 25919 12103 25953
rect 12141 25919 12175 25953
rect 12213 25919 12247 25953
rect 12285 25919 12319 25953
rect 12357 25919 12391 25953
rect 12429 25919 12463 25953
rect 12501 25919 12535 25953
rect 12573 25919 12607 25953
rect 12645 25919 12679 25953
rect 12717 25919 12751 25953
rect 12789 25919 12823 25953
rect 12861 25919 12895 25953
rect 12933 25919 12967 25953
rect 13005 25919 13039 25953
rect 13077 25919 13111 25953
rect 13149 25919 13183 25953
rect 13221 25919 13255 25953
rect 13293 25919 13327 25953
rect 13365 25919 13399 25953
rect 13437 25919 13471 25953
rect 13509 25919 13543 25953
rect 13581 25919 13615 25953
rect 13653 25919 13687 25953
rect 13756 25921 13790 25955
rect 13828 25921 13862 25955
rect 13900 25921 13934 25955
rect 13972 25921 14006 25955
rect 14044 25921 14078 25955
rect 14116 25921 14150 25955
rect 9909 25849 9943 25880
rect 9981 25849 10015 25880
rect 10053 25849 10087 25880
rect 10125 25849 10159 25880
rect 10197 25849 10231 25880
rect 10269 25849 10303 25880
rect 10341 25849 10375 25880
rect 10413 25849 10447 25880
rect 10485 25849 10519 25880
rect 10557 25849 10591 25880
rect 10629 25849 10663 25880
rect 10701 25849 10735 25880
rect 9909 25846 9911 25849
rect 9911 25846 9943 25849
rect 9981 25846 10014 25849
rect 10014 25846 10015 25849
rect 10053 25846 10083 25849
rect 10083 25846 10087 25849
rect 10125 25846 10152 25849
rect 10152 25846 10159 25849
rect 10197 25846 10221 25849
rect 10221 25846 10231 25849
rect 10269 25846 10290 25849
rect 10290 25846 10303 25849
rect 10341 25846 10359 25849
rect 10359 25846 10375 25849
rect 10413 25846 10428 25849
rect 10428 25846 10447 25849
rect 10485 25846 10497 25849
rect 10497 25846 10519 25849
rect 10557 25846 10566 25849
rect 10566 25846 10591 25849
rect 10629 25846 10635 25849
rect 10635 25846 10663 25849
rect 10701 25846 10704 25849
rect 10704 25846 10735 25849
rect 10773 25846 10807 25880
rect 10845 25849 10879 25880
rect 10917 25849 10951 25880
rect 10989 25849 11023 25880
rect 11061 25849 11095 25880
rect 11133 25849 11167 25880
rect 11205 25849 11239 25880
rect 11277 25849 11311 25880
rect 11349 25849 11383 25880
rect 11421 25849 11455 25880
rect 11493 25849 11527 25880
rect 11565 25849 11599 25880
rect 11637 25849 11671 25880
rect 11709 25849 11743 25880
rect 11781 25849 11815 25880
rect 11853 25849 11887 25880
rect 11925 25849 11959 25880
rect 10845 25846 10875 25849
rect 10875 25846 10879 25849
rect 10917 25846 10943 25849
rect 10943 25846 10951 25849
rect 10989 25846 11011 25849
rect 11011 25846 11023 25849
rect 11061 25846 11079 25849
rect 11079 25846 11095 25849
rect 11133 25846 11147 25849
rect 11147 25846 11167 25849
rect 11205 25846 11215 25849
rect 11215 25846 11239 25849
rect 11277 25846 11283 25849
rect 11283 25846 11311 25849
rect 11349 25846 11351 25849
rect 11351 25846 11383 25849
rect 11421 25846 11453 25849
rect 11453 25846 11455 25849
rect 11493 25846 11521 25849
rect 11521 25846 11527 25849
rect 11565 25846 11589 25849
rect 11589 25846 11599 25849
rect 11637 25846 11657 25849
rect 11657 25846 11671 25849
rect 11709 25846 11725 25849
rect 11725 25846 11743 25849
rect 11781 25846 11793 25849
rect 11793 25846 11815 25849
rect 11853 25846 11861 25849
rect 11861 25846 11887 25849
rect 11925 25846 11929 25849
rect 11929 25846 11959 25849
rect 11997 25846 12031 25880
rect 12069 25849 12103 25880
rect 12141 25849 12175 25880
rect 12213 25849 12247 25880
rect 12285 25849 12319 25880
rect 12357 25849 12391 25880
rect 12429 25849 12463 25880
rect 12501 25849 12535 25880
rect 12573 25849 12607 25880
rect 12645 25849 12679 25880
rect 12717 25849 12751 25880
rect 12789 25849 12823 25880
rect 12861 25849 12895 25880
rect 12933 25849 12967 25880
rect 13005 25849 13039 25880
rect 13077 25849 13111 25880
rect 13149 25849 13183 25880
rect 12069 25846 12099 25849
rect 12099 25846 12103 25849
rect 12141 25846 12167 25849
rect 12167 25846 12175 25849
rect 12213 25846 12235 25849
rect 12235 25846 12247 25849
rect 12285 25846 12303 25849
rect 12303 25846 12319 25849
rect 12357 25846 12371 25849
rect 12371 25846 12391 25849
rect 12429 25846 12439 25849
rect 12439 25846 12463 25849
rect 12501 25846 12507 25849
rect 12507 25846 12535 25849
rect 12573 25846 12575 25849
rect 12575 25846 12607 25849
rect 12645 25846 12677 25849
rect 12677 25846 12679 25849
rect 12717 25846 12745 25849
rect 12745 25846 12751 25849
rect 12789 25846 12813 25849
rect 12813 25846 12823 25849
rect 12861 25846 12881 25849
rect 12881 25846 12895 25849
rect 12933 25846 12949 25849
rect 12949 25846 12967 25849
rect 13005 25846 13017 25849
rect 13017 25846 13039 25849
rect 13077 25846 13085 25849
rect 13085 25846 13111 25849
rect 13149 25846 13153 25849
rect 13153 25846 13183 25849
rect 13221 25846 13255 25880
rect 13293 25849 13327 25880
rect 13365 25849 13399 25880
rect 13437 25849 13471 25880
rect 13509 25849 13543 25880
rect 13581 25849 13615 25880
rect 13653 25849 13687 25880
rect 13756 25849 13790 25881
rect 13828 25849 13862 25881
rect 13900 25849 13934 25881
rect 13972 25849 14006 25881
rect 14044 25849 14078 25881
rect 14116 25849 14150 25881
rect 13293 25846 13323 25849
rect 13323 25846 13327 25849
rect 13365 25846 13391 25849
rect 13391 25846 13399 25849
rect 13437 25846 13459 25849
rect 13459 25846 13471 25849
rect 13509 25846 13527 25849
rect 13527 25846 13543 25849
rect 13581 25846 13595 25849
rect 13595 25846 13615 25849
rect 13653 25846 13663 25849
rect 13663 25846 13687 25849
rect 13756 25847 13765 25849
rect 13765 25847 13790 25849
rect 13828 25847 13833 25849
rect 13833 25847 13862 25849
rect 13900 25847 13901 25849
rect 13901 25847 13934 25849
rect 13972 25847 14003 25849
rect 14003 25847 14006 25849
rect 14044 25847 14071 25849
rect 14071 25847 14078 25849
rect 14116 25847 14139 25849
rect 14139 25847 14150 25849
rect 9909 25779 9943 25807
rect 9981 25779 10015 25807
rect 10053 25779 10087 25807
rect 10125 25779 10159 25807
rect 10197 25779 10231 25807
rect 10269 25779 10303 25807
rect 10341 25779 10375 25807
rect 10413 25779 10447 25807
rect 10485 25779 10519 25807
rect 10557 25779 10591 25807
rect 10629 25779 10663 25807
rect 10701 25779 10735 25807
rect 9909 25773 9911 25779
rect 9911 25773 9943 25779
rect 9981 25773 10014 25779
rect 10014 25773 10015 25779
rect 10053 25773 10083 25779
rect 10083 25773 10087 25779
rect 10125 25773 10152 25779
rect 10152 25773 10159 25779
rect 10197 25773 10221 25779
rect 10221 25773 10231 25779
rect 10269 25773 10290 25779
rect 10290 25773 10303 25779
rect 10341 25773 10359 25779
rect 10359 25773 10375 25779
rect 10413 25773 10428 25779
rect 10428 25773 10447 25779
rect 10485 25773 10497 25779
rect 10497 25773 10519 25779
rect 10557 25773 10566 25779
rect 10566 25773 10591 25779
rect 10629 25773 10635 25779
rect 10635 25773 10663 25779
rect 10701 25773 10704 25779
rect 10704 25773 10735 25779
rect 10773 25773 10807 25807
rect 10845 25779 10879 25807
rect 10917 25779 10951 25807
rect 10989 25779 11023 25807
rect 11061 25779 11095 25807
rect 11133 25779 11167 25807
rect 11205 25779 11239 25807
rect 11277 25779 11311 25807
rect 11349 25779 11383 25807
rect 11421 25779 11455 25807
rect 11493 25779 11527 25807
rect 11565 25779 11599 25807
rect 11637 25779 11671 25807
rect 11709 25779 11743 25807
rect 11781 25779 11815 25807
rect 11853 25779 11887 25807
rect 11925 25779 11959 25807
rect 10845 25773 10875 25779
rect 10875 25773 10879 25779
rect 10917 25773 10943 25779
rect 10943 25773 10951 25779
rect 10989 25773 11011 25779
rect 11011 25773 11023 25779
rect 11061 25773 11079 25779
rect 11079 25773 11095 25779
rect 11133 25773 11147 25779
rect 11147 25773 11167 25779
rect 11205 25773 11215 25779
rect 11215 25773 11239 25779
rect 11277 25773 11283 25779
rect 11283 25773 11311 25779
rect 11349 25773 11351 25779
rect 11351 25773 11383 25779
rect 11421 25773 11453 25779
rect 11453 25773 11455 25779
rect 11493 25773 11521 25779
rect 11521 25773 11527 25779
rect 11565 25773 11589 25779
rect 11589 25773 11599 25779
rect 11637 25773 11657 25779
rect 11657 25773 11671 25779
rect 11709 25773 11725 25779
rect 11725 25773 11743 25779
rect 11781 25773 11793 25779
rect 11793 25773 11815 25779
rect 11853 25773 11861 25779
rect 11861 25773 11887 25779
rect 11925 25773 11929 25779
rect 11929 25773 11959 25779
rect 11997 25773 12031 25807
rect 12069 25779 12103 25807
rect 12141 25779 12175 25807
rect 12213 25779 12247 25807
rect 12285 25779 12319 25807
rect 12357 25779 12391 25807
rect 12429 25779 12463 25807
rect 12501 25779 12535 25807
rect 12573 25779 12607 25807
rect 12645 25779 12679 25807
rect 12717 25779 12751 25807
rect 12789 25779 12823 25807
rect 12861 25779 12895 25807
rect 12933 25779 12967 25807
rect 13005 25779 13039 25807
rect 13077 25779 13111 25807
rect 13149 25779 13183 25807
rect 12069 25773 12099 25779
rect 12099 25773 12103 25779
rect 12141 25773 12167 25779
rect 12167 25773 12175 25779
rect 12213 25773 12235 25779
rect 12235 25773 12247 25779
rect 12285 25773 12303 25779
rect 12303 25773 12319 25779
rect 12357 25773 12371 25779
rect 12371 25773 12391 25779
rect 12429 25773 12439 25779
rect 12439 25773 12463 25779
rect 12501 25773 12507 25779
rect 12507 25773 12535 25779
rect 12573 25773 12575 25779
rect 12575 25773 12607 25779
rect 12645 25773 12677 25779
rect 12677 25773 12679 25779
rect 12717 25773 12745 25779
rect 12745 25773 12751 25779
rect 12789 25773 12813 25779
rect 12813 25773 12823 25779
rect 12861 25773 12881 25779
rect 12881 25773 12895 25779
rect 12933 25773 12949 25779
rect 12949 25773 12967 25779
rect 13005 25773 13017 25779
rect 13017 25773 13039 25779
rect 13077 25773 13085 25779
rect 13085 25773 13111 25779
rect 13149 25773 13153 25779
rect 13153 25773 13183 25779
rect 13221 25773 13255 25807
rect 13293 25779 13327 25807
rect 13365 25779 13399 25807
rect 13437 25779 13471 25807
rect 13509 25779 13543 25807
rect 13581 25779 13615 25807
rect 13653 25779 13687 25807
rect 13756 25779 13790 25807
rect 13828 25779 13862 25807
rect 13900 25779 13934 25807
rect 13972 25779 14006 25807
rect 14044 25779 14078 25807
rect 14116 25779 14150 25807
rect 13293 25773 13323 25779
rect 13323 25773 13327 25779
rect 13365 25773 13391 25779
rect 13391 25773 13399 25779
rect 13437 25773 13459 25779
rect 13459 25773 13471 25779
rect 13509 25773 13527 25779
rect 13527 25773 13543 25779
rect 13581 25773 13595 25779
rect 13595 25773 13615 25779
rect 13653 25773 13663 25779
rect 13663 25773 13687 25779
rect 13756 25773 13765 25779
rect 13765 25773 13790 25779
rect 13828 25773 13833 25779
rect 13833 25773 13862 25779
rect 13900 25773 13901 25779
rect 13901 25773 13934 25779
rect 13972 25773 14003 25779
rect 14003 25773 14006 25779
rect 14044 25773 14071 25779
rect 14071 25773 14078 25779
rect 14116 25773 14139 25779
rect 14139 25773 14150 25779
rect 9909 25709 9943 25734
rect 9981 25709 10015 25734
rect 10053 25709 10087 25734
rect 10125 25709 10159 25734
rect 10197 25709 10231 25734
rect 10269 25709 10303 25734
rect 10341 25709 10375 25734
rect 10413 25709 10447 25734
rect 10485 25709 10519 25734
rect 10557 25709 10591 25734
rect 10629 25709 10663 25734
rect 10701 25709 10735 25734
rect 9909 25700 9911 25709
rect 9911 25700 9943 25709
rect 9981 25700 10014 25709
rect 10014 25700 10015 25709
rect 10053 25700 10083 25709
rect 10083 25700 10087 25709
rect 10125 25700 10152 25709
rect 10152 25700 10159 25709
rect 10197 25700 10221 25709
rect 10221 25700 10231 25709
rect 10269 25700 10290 25709
rect 10290 25700 10303 25709
rect 10341 25700 10359 25709
rect 10359 25700 10375 25709
rect 10413 25700 10428 25709
rect 10428 25700 10447 25709
rect 10485 25700 10497 25709
rect 10497 25700 10519 25709
rect 10557 25700 10566 25709
rect 10566 25700 10591 25709
rect 10629 25700 10635 25709
rect 10635 25700 10663 25709
rect 10701 25700 10704 25709
rect 10704 25700 10735 25709
rect 10773 25700 10807 25734
rect 10845 25709 10879 25734
rect 10917 25709 10951 25734
rect 10989 25709 11023 25734
rect 11061 25709 11095 25734
rect 11133 25709 11167 25734
rect 11205 25709 11239 25734
rect 11277 25709 11311 25734
rect 11349 25709 11383 25734
rect 11421 25709 11455 25734
rect 11493 25709 11527 25734
rect 11565 25709 11599 25734
rect 11637 25709 11671 25734
rect 11709 25709 11743 25734
rect 11781 25709 11815 25734
rect 11853 25709 11887 25734
rect 11925 25709 11959 25734
rect 10845 25700 10875 25709
rect 10875 25700 10879 25709
rect 10917 25700 10943 25709
rect 10943 25700 10951 25709
rect 10989 25700 11011 25709
rect 11011 25700 11023 25709
rect 11061 25700 11079 25709
rect 11079 25700 11095 25709
rect 11133 25700 11147 25709
rect 11147 25700 11167 25709
rect 11205 25700 11215 25709
rect 11215 25700 11239 25709
rect 11277 25700 11283 25709
rect 11283 25700 11311 25709
rect 11349 25700 11351 25709
rect 11351 25700 11383 25709
rect 11421 25700 11453 25709
rect 11453 25700 11455 25709
rect 11493 25700 11521 25709
rect 11521 25700 11527 25709
rect 11565 25700 11589 25709
rect 11589 25700 11599 25709
rect 11637 25700 11657 25709
rect 11657 25700 11671 25709
rect 11709 25700 11725 25709
rect 11725 25700 11743 25709
rect 11781 25700 11793 25709
rect 11793 25700 11815 25709
rect 11853 25700 11861 25709
rect 11861 25700 11887 25709
rect 11925 25700 11929 25709
rect 11929 25700 11959 25709
rect 11997 25700 12031 25734
rect 12069 25709 12103 25734
rect 12141 25709 12175 25734
rect 12213 25709 12247 25734
rect 12285 25709 12319 25734
rect 12357 25709 12391 25734
rect 12429 25709 12463 25734
rect 12501 25709 12535 25734
rect 12573 25709 12607 25734
rect 12645 25709 12679 25734
rect 12717 25709 12751 25734
rect 12789 25709 12823 25734
rect 12861 25709 12895 25734
rect 12933 25709 12967 25734
rect 13005 25709 13039 25734
rect 13077 25709 13111 25734
rect 13149 25709 13183 25734
rect 12069 25700 12099 25709
rect 12099 25700 12103 25709
rect 12141 25700 12167 25709
rect 12167 25700 12175 25709
rect 12213 25700 12235 25709
rect 12235 25700 12247 25709
rect 12285 25700 12303 25709
rect 12303 25700 12319 25709
rect 12357 25700 12371 25709
rect 12371 25700 12391 25709
rect 12429 25700 12439 25709
rect 12439 25700 12463 25709
rect 12501 25700 12507 25709
rect 12507 25700 12535 25709
rect 12573 25700 12575 25709
rect 12575 25700 12607 25709
rect 12645 25700 12677 25709
rect 12677 25700 12679 25709
rect 12717 25700 12745 25709
rect 12745 25700 12751 25709
rect 12789 25700 12813 25709
rect 12813 25700 12823 25709
rect 12861 25700 12881 25709
rect 12881 25700 12895 25709
rect 12933 25700 12949 25709
rect 12949 25700 12967 25709
rect 13005 25700 13017 25709
rect 13017 25700 13039 25709
rect 13077 25700 13085 25709
rect 13085 25700 13111 25709
rect 13149 25700 13153 25709
rect 13153 25700 13183 25709
rect 13221 25700 13255 25734
rect 13293 25709 13327 25734
rect 13365 25709 13399 25734
rect 13437 25709 13471 25734
rect 13509 25709 13543 25734
rect 13581 25709 13615 25734
rect 13653 25709 13687 25734
rect 13756 25709 13790 25733
rect 13828 25709 13862 25733
rect 13900 25709 13934 25733
rect 13972 25709 14006 25733
rect 14044 25709 14078 25733
rect 14116 25709 14150 25733
rect 13293 25700 13323 25709
rect 13323 25700 13327 25709
rect 13365 25700 13391 25709
rect 13391 25700 13399 25709
rect 13437 25700 13459 25709
rect 13459 25700 13471 25709
rect 13509 25700 13527 25709
rect 13527 25700 13543 25709
rect 13581 25700 13595 25709
rect 13595 25700 13615 25709
rect 13653 25700 13663 25709
rect 13663 25700 13687 25709
rect 13756 25699 13765 25709
rect 13765 25699 13790 25709
rect 13828 25699 13833 25709
rect 13833 25699 13862 25709
rect 13900 25699 13901 25709
rect 13901 25699 13934 25709
rect 13972 25699 14003 25709
rect 14003 25699 14006 25709
rect 14044 25699 14071 25709
rect 14071 25699 14078 25709
rect 14116 25699 14139 25709
rect 14139 25699 14150 25709
rect 9909 25639 9943 25661
rect 9981 25639 10015 25661
rect 10053 25639 10087 25661
rect 10125 25639 10159 25661
rect 10197 25639 10231 25661
rect 10269 25639 10303 25661
rect 10341 25639 10375 25661
rect 10413 25639 10447 25661
rect 10485 25639 10519 25661
rect 10557 25639 10591 25661
rect 10629 25639 10663 25661
rect 10701 25639 10735 25661
rect 9909 25627 9911 25639
rect 9911 25627 9943 25639
rect 9981 25627 10014 25639
rect 10014 25627 10015 25639
rect 10053 25627 10083 25639
rect 10083 25627 10087 25639
rect 10125 25627 10152 25639
rect 10152 25627 10159 25639
rect 10197 25627 10221 25639
rect 10221 25627 10231 25639
rect 10269 25627 10290 25639
rect 10290 25627 10303 25639
rect 10341 25627 10359 25639
rect 10359 25627 10375 25639
rect 10413 25627 10428 25639
rect 10428 25627 10447 25639
rect 10485 25627 10497 25639
rect 10497 25627 10519 25639
rect 10557 25627 10566 25639
rect 10566 25627 10591 25639
rect 10629 25627 10635 25639
rect 10635 25627 10663 25639
rect 10701 25627 10704 25639
rect 10704 25627 10735 25639
rect 10773 25627 10807 25661
rect 10845 25639 10879 25661
rect 10917 25639 10951 25661
rect 10989 25639 11023 25661
rect 11061 25639 11095 25661
rect 11133 25639 11167 25661
rect 11205 25639 11239 25661
rect 11277 25639 11311 25661
rect 11349 25639 11383 25661
rect 11421 25639 11455 25661
rect 11493 25639 11527 25661
rect 11565 25639 11599 25661
rect 11637 25639 11671 25661
rect 11709 25639 11743 25661
rect 11781 25639 11815 25661
rect 11853 25639 11887 25661
rect 11925 25639 11959 25661
rect 10845 25627 10875 25639
rect 10875 25627 10879 25639
rect 10917 25627 10943 25639
rect 10943 25627 10951 25639
rect 10989 25627 11011 25639
rect 11011 25627 11023 25639
rect 11061 25627 11079 25639
rect 11079 25627 11095 25639
rect 11133 25627 11147 25639
rect 11147 25627 11167 25639
rect 11205 25627 11215 25639
rect 11215 25627 11239 25639
rect 11277 25627 11283 25639
rect 11283 25627 11311 25639
rect 11349 25627 11351 25639
rect 11351 25627 11383 25639
rect 11421 25627 11453 25639
rect 11453 25627 11455 25639
rect 11493 25627 11521 25639
rect 11521 25627 11527 25639
rect 11565 25627 11589 25639
rect 11589 25627 11599 25639
rect 11637 25627 11657 25639
rect 11657 25627 11671 25639
rect 11709 25627 11725 25639
rect 11725 25627 11743 25639
rect 11781 25627 11793 25639
rect 11793 25627 11815 25639
rect 11853 25627 11861 25639
rect 11861 25627 11887 25639
rect 11925 25627 11929 25639
rect 11929 25627 11959 25639
rect 11997 25627 12031 25661
rect 12069 25639 12103 25661
rect 12141 25639 12175 25661
rect 12213 25639 12247 25661
rect 12285 25639 12319 25661
rect 12357 25639 12391 25661
rect 12429 25639 12463 25661
rect 12501 25639 12535 25661
rect 12573 25639 12607 25661
rect 12645 25639 12679 25661
rect 12717 25639 12751 25661
rect 12789 25639 12823 25661
rect 12861 25639 12895 25661
rect 12933 25639 12967 25661
rect 13005 25639 13039 25661
rect 13077 25639 13111 25661
rect 13149 25639 13183 25661
rect 12069 25627 12099 25639
rect 12099 25627 12103 25639
rect 12141 25627 12167 25639
rect 12167 25627 12175 25639
rect 12213 25627 12235 25639
rect 12235 25627 12247 25639
rect 12285 25627 12303 25639
rect 12303 25627 12319 25639
rect 12357 25627 12371 25639
rect 12371 25627 12391 25639
rect 12429 25627 12439 25639
rect 12439 25627 12463 25639
rect 12501 25627 12507 25639
rect 12507 25627 12535 25639
rect 12573 25627 12575 25639
rect 12575 25627 12607 25639
rect 12645 25627 12677 25639
rect 12677 25627 12679 25639
rect 12717 25627 12745 25639
rect 12745 25627 12751 25639
rect 12789 25627 12813 25639
rect 12813 25627 12823 25639
rect 12861 25627 12881 25639
rect 12881 25627 12895 25639
rect 12933 25627 12949 25639
rect 12949 25627 12967 25639
rect 13005 25627 13017 25639
rect 13017 25627 13039 25639
rect 13077 25627 13085 25639
rect 13085 25627 13111 25639
rect 13149 25627 13153 25639
rect 13153 25627 13183 25639
rect 13221 25627 13255 25661
rect 13293 25639 13327 25661
rect 13365 25639 13399 25661
rect 13437 25639 13471 25661
rect 13509 25639 13543 25661
rect 13581 25639 13615 25661
rect 13653 25639 13687 25661
rect 13756 25639 13790 25659
rect 13828 25639 13862 25659
rect 13900 25639 13934 25659
rect 13972 25639 14006 25659
rect 14044 25639 14078 25659
rect 14116 25639 14150 25659
rect 13293 25627 13323 25639
rect 13323 25627 13327 25639
rect 13365 25627 13391 25639
rect 13391 25627 13399 25639
rect 13437 25627 13459 25639
rect 13459 25627 13471 25639
rect 13509 25627 13527 25639
rect 13527 25627 13543 25639
rect 13581 25627 13595 25639
rect 13595 25627 13615 25639
rect 13653 25627 13663 25639
rect 13663 25627 13687 25639
rect 13756 25625 13765 25639
rect 13765 25625 13790 25639
rect 13828 25625 13833 25639
rect 13833 25625 13862 25639
rect 13900 25625 13901 25639
rect 13901 25625 13934 25639
rect 13972 25625 14003 25639
rect 14003 25625 14006 25639
rect 14044 25625 14071 25639
rect 14071 25625 14078 25639
rect 14116 25625 14139 25639
rect 14139 25625 14150 25639
rect 9909 25569 9943 25588
rect 9981 25569 10015 25588
rect 10053 25569 10087 25588
rect 10125 25569 10159 25588
rect 10197 25569 10231 25588
rect 10269 25569 10303 25588
rect 10341 25569 10375 25588
rect 10413 25569 10447 25588
rect 10485 25569 10519 25588
rect 10557 25569 10591 25588
rect 10629 25569 10663 25588
rect 10701 25569 10735 25588
rect 9909 25554 9911 25569
rect 9911 25554 9943 25569
rect 9981 25554 10014 25569
rect 10014 25554 10015 25569
rect 10053 25554 10083 25569
rect 10083 25554 10087 25569
rect 10125 25554 10152 25569
rect 10152 25554 10159 25569
rect 10197 25554 10221 25569
rect 10221 25554 10231 25569
rect 10269 25554 10290 25569
rect 10290 25554 10303 25569
rect 10341 25554 10359 25569
rect 10359 25554 10375 25569
rect 10413 25554 10428 25569
rect 10428 25554 10447 25569
rect 10485 25554 10497 25569
rect 10497 25554 10519 25569
rect 10557 25554 10566 25569
rect 10566 25554 10591 25569
rect 10629 25554 10635 25569
rect 10635 25554 10663 25569
rect 10701 25554 10704 25569
rect 10704 25554 10735 25569
rect 10773 25554 10807 25588
rect 10845 25569 10879 25588
rect 10917 25569 10951 25588
rect 10989 25569 11023 25588
rect 11061 25569 11095 25588
rect 11133 25569 11167 25588
rect 11205 25569 11239 25588
rect 11277 25569 11311 25588
rect 11349 25569 11383 25588
rect 11421 25569 11455 25588
rect 11493 25569 11527 25588
rect 11565 25569 11599 25588
rect 11637 25569 11671 25588
rect 11709 25569 11743 25588
rect 11781 25569 11815 25588
rect 11853 25569 11887 25588
rect 11925 25569 11959 25588
rect 10845 25554 10875 25569
rect 10875 25554 10879 25569
rect 10917 25554 10943 25569
rect 10943 25554 10951 25569
rect 10989 25554 11011 25569
rect 11011 25554 11023 25569
rect 11061 25554 11079 25569
rect 11079 25554 11095 25569
rect 11133 25554 11147 25569
rect 11147 25554 11167 25569
rect 11205 25554 11215 25569
rect 11215 25554 11239 25569
rect 11277 25554 11283 25569
rect 11283 25554 11311 25569
rect 11349 25554 11351 25569
rect 11351 25554 11383 25569
rect 11421 25554 11453 25569
rect 11453 25554 11455 25569
rect 11493 25554 11521 25569
rect 11521 25554 11527 25569
rect 11565 25554 11589 25569
rect 11589 25554 11599 25569
rect 11637 25554 11657 25569
rect 11657 25554 11671 25569
rect 11709 25554 11725 25569
rect 11725 25554 11743 25569
rect 11781 25554 11793 25569
rect 11793 25554 11815 25569
rect 11853 25554 11861 25569
rect 11861 25554 11887 25569
rect 11925 25554 11929 25569
rect 11929 25554 11959 25569
rect 11997 25554 12031 25588
rect 12069 25569 12103 25588
rect 12141 25569 12175 25588
rect 12213 25569 12247 25588
rect 12285 25569 12319 25588
rect 12357 25569 12391 25588
rect 12429 25569 12463 25588
rect 12501 25569 12535 25588
rect 12573 25569 12607 25588
rect 12645 25569 12679 25588
rect 12717 25569 12751 25588
rect 12789 25569 12823 25588
rect 12861 25569 12895 25588
rect 12933 25569 12967 25588
rect 13005 25569 13039 25588
rect 13077 25569 13111 25588
rect 13149 25569 13183 25588
rect 12069 25554 12099 25569
rect 12099 25554 12103 25569
rect 12141 25554 12167 25569
rect 12167 25554 12175 25569
rect 12213 25554 12235 25569
rect 12235 25554 12247 25569
rect 12285 25554 12303 25569
rect 12303 25554 12319 25569
rect 12357 25554 12371 25569
rect 12371 25554 12391 25569
rect 12429 25554 12439 25569
rect 12439 25554 12463 25569
rect 12501 25554 12507 25569
rect 12507 25554 12535 25569
rect 12573 25554 12575 25569
rect 12575 25554 12607 25569
rect 12645 25554 12677 25569
rect 12677 25554 12679 25569
rect 12717 25554 12745 25569
rect 12745 25554 12751 25569
rect 12789 25554 12813 25569
rect 12813 25554 12823 25569
rect 12861 25554 12881 25569
rect 12881 25554 12895 25569
rect 12933 25554 12949 25569
rect 12949 25554 12967 25569
rect 13005 25554 13017 25569
rect 13017 25554 13039 25569
rect 13077 25554 13085 25569
rect 13085 25554 13111 25569
rect 13149 25554 13153 25569
rect 13153 25554 13183 25569
rect 13221 25554 13255 25588
rect 13293 25569 13327 25588
rect 13365 25569 13399 25588
rect 13437 25569 13471 25588
rect 13509 25569 13543 25588
rect 13581 25569 13615 25588
rect 13653 25569 13687 25588
rect 13756 25569 13790 25585
rect 13828 25569 13862 25585
rect 13900 25569 13934 25585
rect 13972 25569 14006 25585
rect 14044 25569 14078 25585
rect 14116 25569 14150 25585
rect 13293 25554 13323 25569
rect 13323 25554 13327 25569
rect 13365 25554 13391 25569
rect 13391 25554 13399 25569
rect 13437 25554 13459 25569
rect 13459 25554 13471 25569
rect 13509 25554 13527 25569
rect 13527 25554 13543 25569
rect 13581 25554 13595 25569
rect 13595 25554 13615 25569
rect 13653 25554 13663 25569
rect 13663 25554 13687 25569
rect 13756 25551 13765 25569
rect 13765 25551 13790 25569
rect 13828 25551 13833 25569
rect 13833 25551 13862 25569
rect 13900 25551 13901 25569
rect 13901 25551 13934 25569
rect 13972 25551 14003 25569
rect 14003 25551 14006 25569
rect 14044 25551 14071 25569
rect 14071 25551 14078 25569
rect 14116 25551 14139 25569
rect 14139 25551 14150 25569
rect 9909 25499 9943 25515
rect 9981 25499 10015 25515
rect 10053 25499 10087 25515
rect 10125 25499 10159 25515
rect 10197 25499 10231 25515
rect 10269 25499 10303 25515
rect 10341 25499 10375 25515
rect 10413 25499 10447 25515
rect 10485 25499 10519 25515
rect 10557 25499 10591 25515
rect 10629 25499 10663 25515
rect 10701 25499 10735 25515
rect 9909 25481 9911 25499
rect 9911 25481 9943 25499
rect 9981 25481 10014 25499
rect 10014 25481 10015 25499
rect 10053 25481 10083 25499
rect 10083 25481 10087 25499
rect 10125 25481 10152 25499
rect 10152 25481 10159 25499
rect 10197 25481 10221 25499
rect 10221 25481 10231 25499
rect 10269 25481 10290 25499
rect 10290 25481 10303 25499
rect 10341 25481 10359 25499
rect 10359 25481 10375 25499
rect 10413 25481 10428 25499
rect 10428 25481 10447 25499
rect 10485 25481 10497 25499
rect 10497 25481 10519 25499
rect 10557 25481 10566 25499
rect 10566 25481 10591 25499
rect 10629 25481 10635 25499
rect 10635 25481 10663 25499
rect 10701 25481 10704 25499
rect 10704 25481 10735 25499
rect 10773 25481 10807 25515
rect 10845 25499 10879 25515
rect 10917 25499 10951 25515
rect 10989 25499 11023 25515
rect 11061 25499 11095 25515
rect 11133 25499 11167 25515
rect 11205 25499 11239 25515
rect 11277 25499 11311 25515
rect 11349 25499 11383 25515
rect 11421 25499 11455 25515
rect 11493 25499 11527 25515
rect 11565 25499 11599 25515
rect 11637 25499 11671 25515
rect 11709 25499 11743 25515
rect 11781 25499 11815 25515
rect 11853 25499 11887 25515
rect 11925 25499 11959 25515
rect 10845 25481 10875 25499
rect 10875 25481 10879 25499
rect 10917 25481 10943 25499
rect 10943 25481 10951 25499
rect 10989 25481 11011 25499
rect 11011 25481 11023 25499
rect 11061 25481 11079 25499
rect 11079 25481 11095 25499
rect 11133 25481 11147 25499
rect 11147 25481 11167 25499
rect 11205 25481 11215 25499
rect 11215 25481 11239 25499
rect 11277 25481 11283 25499
rect 11283 25481 11311 25499
rect 11349 25481 11351 25499
rect 11351 25481 11383 25499
rect 11421 25481 11453 25499
rect 11453 25481 11455 25499
rect 11493 25481 11521 25499
rect 11521 25481 11527 25499
rect 11565 25481 11589 25499
rect 11589 25481 11599 25499
rect 11637 25481 11657 25499
rect 11657 25481 11671 25499
rect 11709 25481 11725 25499
rect 11725 25481 11743 25499
rect 11781 25481 11793 25499
rect 11793 25481 11815 25499
rect 11853 25481 11861 25499
rect 11861 25481 11887 25499
rect 11925 25481 11929 25499
rect 11929 25481 11959 25499
rect 11997 25481 12031 25515
rect 12069 25499 12103 25515
rect 12141 25499 12175 25515
rect 12213 25499 12247 25515
rect 12285 25499 12319 25515
rect 12357 25499 12391 25515
rect 12429 25499 12463 25515
rect 12501 25499 12535 25515
rect 12573 25499 12607 25515
rect 12645 25499 12679 25515
rect 12717 25499 12751 25515
rect 12789 25499 12823 25515
rect 12861 25499 12895 25515
rect 12933 25499 12967 25515
rect 13005 25499 13039 25515
rect 13077 25499 13111 25515
rect 13149 25499 13183 25515
rect 12069 25481 12099 25499
rect 12099 25481 12103 25499
rect 12141 25481 12167 25499
rect 12167 25481 12175 25499
rect 12213 25481 12235 25499
rect 12235 25481 12247 25499
rect 12285 25481 12303 25499
rect 12303 25481 12319 25499
rect 12357 25481 12371 25499
rect 12371 25481 12391 25499
rect 12429 25481 12439 25499
rect 12439 25481 12463 25499
rect 12501 25481 12507 25499
rect 12507 25481 12535 25499
rect 12573 25481 12575 25499
rect 12575 25481 12607 25499
rect 12645 25481 12677 25499
rect 12677 25481 12679 25499
rect 12717 25481 12745 25499
rect 12745 25481 12751 25499
rect 12789 25481 12813 25499
rect 12813 25481 12823 25499
rect 12861 25481 12881 25499
rect 12881 25481 12895 25499
rect 12933 25481 12949 25499
rect 12949 25481 12967 25499
rect 13005 25481 13017 25499
rect 13017 25481 13039 25499
rect 13077 25481 13085 25499
rect 13085 25481 13111 25499
rect 13149 25481 13153 25499
rect 13153 25481 13183 25499
rect 13221 25481 13255 25515
rect 13293 25499 13327 25515
rect 13365 25499 13399 25515
rect 13437 25499 13471 25515
rect 13509 25499 13543 25515
rect 13581 25499 13615 25515
rect 13653 25499 13687 25515
rect 13756 25499 13790 25511
rect 13828 25499 13862 25511
rect 13900 25499 13934 25511
rect 13972 25499 14006 25511
rect 14044 25499 14078 25511
rect 14116 25499 14150 25511
rect 13293 25481 13323 25499
rect 13323 25481 13327 25499
rect 13365 25481 13391 25499
rect 13391 25481 13399 25499
rect 13437 25481 13459 25499
rect 13459 25481 13471 25499
rect 13509 25481 13527 25499
rect 13527 25481 13543 25499
rect 13581 25481 13595 25499
rect 13595 25481 13615 25499
rect 13653 25481 13663 25499
rect 13663 25481 13687 25499
rect 13756 25477 13765 25499
rect 13765 25477 13790 25499
rect 13828 25477 13833 25499
rect 13833 25477 13862 25499
rect 13900 25477 13901 25499
rect 13901 25477 13934 25499
rect 13972 25477 14003 25499
rect 14003 25477 14006 25499
rect 14044 25477 14071 25499
rect 14071 25477 14078 25499
rect 14116 25477 14139 25499
rect 14139 25477 14150 25499
rect 9909 25429 9943 25442
rect 9981 25429 10015 25442
rect 10053 25429 10087 25442
rect 10125 25429 10159 25442
rect 10197 25429 10231 25442
rect 10269 25429 10303 25442
rect 10341 25429 10375 25442
rect 10413 25429 10447 25442
rect 10485 25429 10519 25442
rect 10557 25429 10591 25442
rect 10629 25429 10663 25442
rect 10701 25429 10735 25442
rect 9909 25408 9911 25429
rect 9911 25408 9943 25429
rect 9981 25408 10014 25429
rect 10014 25408 10015 25429
rect 10053 25408 10083 25429
rect 10083 25408 10087 25429
rect 10125 25408 10152 25429
rect 10152 25408 10159 25429
rect 10197 25408 10221 25429
rect 10221 25408 10231 25429
rect 10269 25408 10290 25429
rect 10290 25408 10303 25429
rect 10341 25408 10359 25429
rect 10359 25408 10375 25429
rect 10413 25408 10428 25429
rect 10428 25408 10447 25429
rect 10485 25408 10497 25429
rect 10497 25408 10519 25429
rect 10557 25408 10566 25429
rect 10566 25408 10591 25429
rect 10629 25408 10635 25429
rect 10635 25408 10663 25429
rect 10701 25408 10704 25429
rect 10704 25408 10735 25429
rect 10773 25408 10807 25442
rect 10845 25429 10879 25442
rect 10917 25429 10951 25442
rect 10989 25429 11023 25442
rect 11061 25429 11095 25442
rect 11133 25429 11167 25442
rect 11205 25429 11239 25442
rect 11277 25429 11311 25442
rect 11349 25429 11383 25442
rect 11421 25429 11455 25442
rect 11493 25429 11527 25442
rect 11565 25429 11599 25442
rect 11637 25429 11671 25442
rect 11709 25429 11743 25442
rect 11781 25429 11815 25442
rect 11853 25429 11887 25442
rect 11925 25429 11959 25442
rect 10845 25408 10875 25429
rect 10875 25408 10879 25429
rect 10917 25408 10943 25429
rect 10943 25408 10951 25429
rect 10989 25408 11011 25429
rect 11011 25408 11023 25429
rect 11061 25408 11079 25429
rect 11079 25408 11095 25429
rect 11133 25408 11147 25429
rect 11147 25408 11167 25429
rect 11205 25408 11215 25429
rect 11215 25408 11239 25429
rect 11277 25408 11283 25429
rect 11283 25408 11311 25429
rect 11349 25408 11351 25429
rect 11351 25408 11383 25429
rect 11421 25408 11453 25429
rect 11453 25408 11455 25429
rect 11493 25408 11521 25429
rect 11521 25408 11527 25429
rect 11565 25408 11589 25429
rect 11589 25408 11599 25429
rect 11637 25408 11657 25429
rect 11657 25408 11671 25429
rect 11709 25408 11725 25429
rect 11725 25408 11743 25429
rect 11781 25408 11793 25429
rect 11793 25408 11815 25429
rect 11853 25408 11861 25429
rect 11861 25408 11887 25429
rect 11925 25408 11929 25429
rect 11929 25408 11959 25429
rect 11997 25408 12031 25442
rect 12069 25429 12103 25442
rect 12141 25429 12175 25442
rect 12213 25429 12247 25442
rect 12285 25429 12319 25442
rect 12357 25429 12391 25442
rect 12429 25429 12463 25442
rect 12501 25429 12535 25442
rect 12573 25429 12607 25442
rect 12645 25429 12679 25442
rect 12717 25429 12751 25442
rect 12789 25429 12823 25442
rect 12861 25429 12895 25442
rect 12933 25429 12967 25442
rect 13005 25429 13039 25442
rect 13077 25429 13111 25442
rect 13149 25429 13183 25442
rect 12069 25408 12099 25429
rect 12099 25408 12103 25429
rect 12141 25408 12167 25429
rect 12167 25408 12175 25429
rect 12213 25408 12235 25429
rect 12235 25408 12247 25429
rect 12285 25408 12303 25429
rect 12303 25408 12319 25429
rect 12357 25408 12371 25429
rect 12371 25408 12391 25429
rect 12429 25408 12439 25429
rect 12439 25408 12463 25429
rect 12501 25408 12507 25429
rect 12507 25408 12535 25429
rect 12573 25408 12575 25429
rect 12575 25408 12607 25429
rect 12645 25408 12677 25429
rect 12677 25408 12679 25429
rect 12717 25408 12745 25429
rect 12745 25408 12751 25429
rect 12789 25408 12813 25429
rect 12813 25408 12823 25429
rect 12861 25408 12881 25429
rect 12881 25408 12895 25429
rect 12933 25408 12949 25429
rect 12949 25408 12967 25429
rect 13005 25408 13017 25429
rect 13017 25408 13039 25429
rect 13077 25408 13085 25429
rect 13085 25408 13111 25429
rect 13149 25408 13153 25429
rect 13153 25408 13183 25429
rect 13221 25408 13255 25442
rect 13293 25429 13327 25442
rect 13365 25429 13399 25442
rect 13437 25429 13471 25442
rect 13509 25429 13543 25442
rect 13581 25429 13615 25442
rect 13653 25429 13687 25442
rect 13756 25429 13790 25437
rect 13828 25429 13862 25437
rect 13900 25429 13934 25437
rect 13972 25429 14006 25437
rect 14044 25429 14078 25437
rect 14116 25429 14150 25437
rect 13293 25408 13323 25429
rect 13323 25408 13327 25429
rect 13365 25408 13391 25429
rect 13391 25408 13399 25429
rect 13437 25408 13459 25429
rect 13459 25408 13471 25429
rect 13509 25408 13527 25429
rect 13527 25408 13543 25429
rect 13581 25408 13595 25429
rect 13595 25408 13615 25429
rect 13653 25408 13663 25429
rect 13663 25408 13687 25429
rect 13756 25403 13765 25429
rect 13765 25403 13790 25429
rect 13828 25403 13833 25429
rect 13833 25403 13862 25429
rect 13900 25403 13901 25429
rect 13901 25403 13934 25429
rect 13972 25403 14003 25429
rect 14003 25403 14006 25429
rect 14044 25403 14071 25429
rect 14071 25403 14078 25429
rect 14116 25403 14139 25429
rect 14139 25403 14150 25429
rect 9909 25359 9943 25369
rect 9981 25359 10015 25369
rect 10053 25359 10087 25369
rect 10125 25359 10159 25369
rect 10197 25359 10231 25369
rect 10269 25359 10303 25369
rect 10341 25359 10375 25369
rect 10413 25359 10447 25369
rect 10485 25359 10519 25369
rect 10557 25359 10591 25369
rect 10629 25359 10663 25369
rect 10701 25359 10735 25369
rect 9909 25335 9911 25359
rect 9911 25335 9943 25359
rect 9981 25335 10014 25359
rect 10014 25335 10015 25359
rect 10053 25335 10083 25359
rect 10083 25335 10087 25359
rect 10125 25335 10152 25359
rect 10152 25335 10159 25359
rect 10197 25335 10221 25359
rect 10221 25335 10231 25359
rect 10269 25335 10290 25359
rect 10290 25335 10303 25359
rect 10341 25335 10359 25359
rect 10359 25335 10375 25359
rect 10413 25335 10428 25359
rect 10428 25335 10447 25359
rect 10485 25335 10497 25359
rect 10497 25335 10519 25359
rect 10557 25335 10566 25359
rect 10566 25335 10591 25359
rect 10629 25335 10635 25359
rect 10635 25335 10663 25359
rect 10701 25335 10704 25359
rect 10704 25335 10735 25359
rect 10773 25335 10807 25369
rect 10845 25359 10879 25369
rect 10917 25359 10951 25369
rect 10989 25359 11023 25369
rect 11061 25359 11095 25369
rect 11133 25359 11167 25369
rect 11205 25359 11239 25369
rect 11277 25359 11311 25369
rect 11349 25359 11383 25369
rect 11421 25359 11455 25369
rect 11493 25359 11527 25369
rect 11565 25359 11599 25369
rect 11637 25359 11671 25369
rect 11709 25359 11743 25369
rect 11781 25359 11815 25369
rect 11853 25359 11887 25369
rect 11925 25359 11959 25369
rect 10845 25335 10875 25359
rect 10875 25335 10879 25359
rect 10917 25335 10943 25359
rect 10943 25335 10951 25359
rect 10989 25335 11011 25359
rect 11011 25335 11023 25359
rect 11061 25335 11079 25359
rect 11079 25335 11095 25359
rect 11133 25335 11147 25359
rect 11147 25335 11167 25359
rect 11205 25335 11215 25359
rect 11215 25335 11239 25359
rect 11277 25335 11283 25359
rect 11283 25335 11311 25359
rect 11349 25335 11351 25359
rect 11351 25335 11383 25359
rect 11421 25335 11453 25359
rect 11453 25335 11455 25359
rect 11493 25335 11521 25359
rect 11521 25335 11527 25359
rect 11565 25335 11589 25359
rect 11589 25335 11599 25359
rect 11637 25335 11657 25359
rect 11657 25335 11671 25359
rect 11709 25335 11725 25359
rect 11725 25335 11743 25359
rect 11781 25335 11793 25359
rect 11793 25335 11815 25359
rect 11853 25335 11861 25359
rect 11861 25335 11887 25359
rect 11925 25335 11929 25359
rect 11929 25335 11959 25359
rect 11997 25335 12031 25369
rect 12069 25359 12103 25369
rect 12141 25359 12175 25369
rect 12213 25359 12247 25369
rect 12285 25359 12319 25369
rect 12357 25359 12391 25369
rect 12429 25359 12463 25369
rect 12501 25359 12535 25369
rect 12573 25359 12607 25369
rect 12645 25359 12679 25369
rect 12717 25359 12751 25369
rect 12789 25359 12823 25369
rect 12861 25359 12895 25369
rect 12933 25359 12967 25369
rect 13005 25359 13039 25369
rect 13077 25359 13111 25369
rect 13149 25359 13183 25369
rect 12069 25335 12099 25359
rect 12099 25335 12103 25359
rect 12141 25335 12167 25359
rect 12167 25335 12175 25359
rect 12213 25335 12235 25359
rect 12235 25335 12247 25359
rect 12285 25335 12303 25359
rect 12303 25335 12319 25359
rect 12357 25335 12371 25359
rect 12371 25335 12391 25359
rect 12429 25335 12439 25359
rect 12439 25335 12463 25359
rect 12501 25335 12507 25359
rect 12507 25335 12535 25359
rect 12573 25335 12575 25359
rect 12575 25335 12607 25359
rect 12645 25335 12677 25359
rect 12677 25335 12679 25359
rect 12717 25335 12745 25359
rect 12745 25335 12751 25359
rect 12789 25335 12813 25359
rect 12813 25335 12823 25359
rect 12861 25335 12881 25359
rect 12881 25335 12895 25359
rect 12933 25335 12949 25359
rect 12949 25335 12967 25359
rect 13005 25335 13017 25359
rect 13017 25335 13039 25359
rect 13077 25335 13085 25359
rect 13085 25335 13111 25359
rect 13149 25335 13153 25359
rect 13153 25335 13183 25359
rect 13221 25335 13255 25369
rect 13293 25359 13327 25369
rect 13365 25359 13399 25369
rect 13437 25359 13471 25369
rect 13509 25359 13543 25369
rect 13581 25359 13615 25369
rect 13653 25359 13687 25369
rect 13756 25359 13790 25363
rect 13828 25359 13862 25363
rect 13900 25359 13934 25363
rect 13972 25359 14006 25363
rect 14044 25359 14078 25363
rect 14116 25359 14150 25363
rect 13293 25335 13323 25359
rect 13323 25335 13327 25359
rect 13365 25335 13391 25359
rect 13391 25335 13399 25359
rect 13437 25335 13459 25359
rect 13459 25335 13471 25359
rect 13509 25335 13527 25359
rect 13527 25335 13543 25359
rect 13581 25335 13595 25359
rect 13595 25335 13615 25359
rect 13653 25335 13663 25359
rect 13663 25335 13687 25359
rect 13756 25329 13765 25359
rect 13765 25329 13790 25359
rect 13828 25329 13833 25359
rect 13833 25329 13862 25359
rect 13900 25329 13901 25359
rect 13901 25329 13934 25359
rect 13972 25329 14003 25359
rect 14003 25329 14006 25359
rect 14044 25329 14071 25359
rect 14071 25329 14078 25359
rect 14116 25329 14139 25359
rect 14139 25329 14150 25359
rect 9909 25289 9943 25296
rect 9981 25289 10015 25296
rect 10053 25289 10087 25296
rect 10125 25289 10159 25296
rect 10197 25289 10231 25296
rect 10269 25289 10303 25296
rect 10341 25289 10375 25296
rect 10413 25289 10447 25296
rect 10485 25289 10519 25296
rect 10557 25289 10591 25296
rect 10629 25289 10663 25296
rect 10701 25289 10735 25296
rect 9909 25262 9911 25289
rect 9911 25262 9943 25289
rect 9981 25262 10014 25289
rect 10014 25262 10015 25289
rect 10053 25262 10083 25289
rect 10083 25262 10087 25289
rect 10125 25262 10152 25289
rect 10152 25262 10159 25289
rect 10197 25262 10221 25289
rect 10221 25262 10231 25289
rect 10269 25262 10290 25289
rect 10290 25262 10303 25289
rect 10341 25262 10359 25289
rect 10359 25262 10375 25289
rect 10413 25262 10428 25289
rect 10428 25262 10447 25289
rect 10485 25262 10497 25289
rect 10497 25262 10519 25289
rect 10557 25262 10566 25289
rect 10566 25262 10591 25289
rect 10629 25262 10635 25289
rect 10635 25262 10663 25289
rect 10701 25262 10704 25289
rect 10704 25262 10735 25289
rect 10773 25262 10807 25296
rect 10845 25289 10879 25296
rect 10917 25289 10951 25296
rect 10989 25289 11023 25296
rect 11061 25289 11095 25296
rect 11133 25289 11167 25296
rect 11205 25289 11239 25296
rect 11277 25289 11311 25296
rect 11349 25289 11383 25296
rect 11421 25289 11455 25296
rect 11493 25289 11527 25296
rect 11565 25289 11599 25296
rect 11637 25289 11671 25296
rect 11709 25289 11743 25296
rect 11781 25289 11815 25296
rect 11853 25289 11887 25296
rect 11925 25289 11959 25296
rect 10845 25262 10875 25289
rect 10875 25262 10879 25289
rect 10917 25262 10943 25289
rect 10943 25262 10951 25289
rect 10989 25262 11011 25289
rect 11011 25262 11023 25289
rect 11061 25262 11079 25289
rect 11079 25262 11095 25289
rect 11133 25262 11147 25289
rect 11147 25262 11167 25289
rect 11205 25262 11215 25289
rect 11215 25262 11239 25289
rect 11277 25262 11283 25289
rect 11283 25262 11311 25289
rect 11349 25262 11351 25289
rect 11351 25262 11383 25289
rect 11421 25262 11453 25289
rect 11453 25262 11455 25289
rect 11493 25262 11521 25289
rect 11521 25262 11527 25289
rect 11565 25262 11589 25289
rect 11589 25262 11599 25289
rect 11637 25262 11657 25289
rect 11657 25262 11671 25289
rect 11709 25262 11725 25289
rect 11725 25262 11743 25289
rect 11781 25262 11793 25289
rect 11793 25262 11815 25289
rect 11853 25262 11861 25289
rect 11861 25262 11887 25289
rect 11925 25262 11929 25289
rect 11929 25262 11959 25289
rect 11997 25262 12031 25296
rect 12069 25289 12103 25296
rect 12141 25289 12175 25296
rect 12213 25289 12247 25296
rect 12285 25289 12319 25296
rect 12357 25289 12391 25296
rect 12429 25289 12463 25296
rect 12501 25289 12535 25296
rect 12573 25289 12607 25296
rect 12645 25289 12679 25296
rect 12717 25289 12751 25296
rect 12789 25289 12823 25296
rect 12861 25289 12895 25296
rect 12933 25289 12967 25296
rect 13005 25289 13039 25296
rect 13077 25289 13111 25296
rect 13149 25289 13183 25296
rect 12069 25262 12099 25289
rect 12099 25262 12103 25289
rect 12141 25262 12167 25289
rect 12167 25262 12175 25289
rect 12213 25262 12235 25289
rect 12235 25262 12247 25289
rect 12285 25262 12303 25289
rect 12303 25262 12319 25289
rect 12357 25262 12371 25289
rect 12371 25262 12391 25289
rect 12429 25262 12439 25289
rect 12439 25262 12463 25289
rect 12501 25262 12507 25289
rect 12507 25262 12535 25289
rect 12573 25262 12575 25289
rect 12575 25262 12607 25289
rect 12645 25262 12677 25289
rect 12677 25262 12679 25289
rect 12717 25262 12745 25289
rect 12745 25262 12751 25289
rect 12789 25262 12813 25289
rect 12813 25262 12823 25289
rect 12861 25262 12881 25289
rect 12881 25262 12895 25289
rect 12933 25262 12949 25289
rect 12949 25262 12967 25289
rect 13005 25262 13017 25289
rect 13017 25262 13039 25289
rect 13077 25262 13085 25289
rect 13085 25262 13111 25289
rect 13149 25262 13153 25289
rect 13153 25262 13183 25289
rect 13221 25262 13255 25296
rect 13293 25289 13327 25296
rect 13365 25289 13399 25296
rect 13437 25289 13471 25296
rect 13509 25289 13543 25296
rect 13581 25289 13615 25296
rect 13653 25289 13687 25296
rect 13293 25262 13323 25289
rect 13323 25262 13327 25289
rect 13365 25262 13391 25289
rect 13391 25262 13399 25289
rect 13437 25262 13459 25289
rect 13459 25262 13471 25289
rect 13509 25262 13527 25289
rect 13527 25262 13543 25289
rect 13581 25262 13595 25289
rect 13595 25262 13615 25289
rect 13653 25262 13663 25289
rect 13663 25262 13687 25289
rect 13756 25255 13765 25289
rect 13765 25255 13790 25289
rect 13828 25255 13833 25289
rect 13833 25255 13862 25289
rect 13900 25255 13901 25289
rect 13901 25255 13934 25289
rect 13972 25255 14003 25289
rect 14003 25255 14006 25289
rect 14044 25255 14071 25289
rect 14071 25255 14078 25289
rect 14116 25255 14139 25289
rect 14139 25255 14150 25289
rect 9909 25219 9943 25223
rect 9981 25219 10015 25223
rect 10053 25219 10087 25223
rect 10125 25219 10159 25223
rect 10197 25219 10231 25223
rect 10269 25219 10303 25223
rect 10341 25219 10375 25223
rect 10413 25219 10447 25223
rect 10485 25219 10519 25223
rect 10557 25219 10591 25223
rect 10629 25219 10663 25223
rect 10701 25219 10735 25223
rect 9909 25189 9911 25219
rect 9911 25189 9943 25219
rect 9981 25189 10014 25219
rect 10014 25189 10015 25219
rect 10053 25189 10083 25219
rect 10083 25189 10087 25219
rect 10125 25189 10152 25219
rect 10152 25189 10159 25219
rect 10197 25189 10221 25219
rect 10221 25189 10231 25219
rect 10269 25189 10290 25219
rect 10290 25189 10303 25219
rect 10341 25189 10359 25219
rect 10359 25189 10375 25219
rect 10413 25189 10428 25219
rect 10428 25189 10447 25219
rect 10485 25189 10497 25219
rect 10497 25189 10519 25219
rect 10557 25189 10566 25219
rect 10566 25189 10591 25219
rect 10629 25189 10635 25219
rect 10635 25189 10663 25219
rect 10701 25189 10704 25219
rect 10704 25189 10735 25219
rect 10773 25189 10807 25223
rect 10845 25219 10879 25223
rect 10917 25219 10951 25223
rect 10989 25219 11023 25223
rect 11061 25219 11095 25223
rect 11133 25219 11167 25223
rect 11205 25219 11239 25223
rect 11277 25219 11311 25223
rect 11349 25219 11383 25223
rect 11421 25219 11455 25223
rect 11493 25219 11527 25223
rect 11565 25219 11599 25223
rect 11637 25219 11671 25223
rect 11709 25219 11743 25223
rect 11781 25219 11815 25223
rect 11853 25219 11887 25223
rect 11925 25219 11959 25223
rect 10845 25189 10875 25219
rect 10875 25189 10879 25219
rect 10917 25189 10943 25219
rect 10943 25189 10951 25219
rect 10989 25189 11011 25219
rect 11011 25189 11023 25219
rect 11061 25189 11079 25219
rect 11079 25189 11095 25219
rect 11133 25189 11147 25219
rect 11147 25189 11167 25219
rect 11205 25189 11215 25219
rect 11215 25189 11239 25219
rect 11277 25189 11283 25219
rect 11283 25189 11311 25219
rect 11349 25189 11351 25219
rect 11351 25189 11383 25219
rect 11421 25189 11453 25219
rect 11453 25189 11455 25219
rect 11493 25189 11521 25219
rect 11521 25189 11527 25219
rect 11565 25189 11589 25219
rect 11589 25189 11599 25219
rect 11637 25189 11657 25219
rect 11657 25189 11671 25219
rect 11709 25189 11725 25219
rect 11725 25189 11743 25219
rect 11781 25189 11793 25219
rect 11793 25189 11815 25219
rect 11853 25189 11861 25219
rect 11861 25189 11887 25219
rect 11925 25189 11929 25219
rect 11929 25189 11959 25219
rect 11997 25189 12031 25223
rect 12069 25219 12103 25223
rect 12141 25219 12175 25223
rect 12213 25219 12247 25223
rect 12285 25219 12319 25223
rect 12357 25219 12391 25223
rect 12429 25219 12463 25223
rect 12501 25219 12535 25223
rect 12573 25219 12607 25223
rect 12645 25219 12679 25223
rect 12717 25219 12751 25223
rect 12789 25219 12823 25223
rect 12861 25219 12895 25223
rect 12933 25219 12967 25223
rect 13005 25219 13039 25223
rect 13077 25219 13111 25223
rect 13149 25219 13183 25223
rect 12069 25189 12099 25219
rect 12099 25189 12103 25219
rect 12141 25189 12167 25219
rect 12167 25189 12175 25219
rect 12213 25189 12235 25219
rect 12235 25189 12247 25219
rect 12285 25189 12303 25219
rect 12303 25189 12319 25219
rect 12357 25189 12371 25219
rect 12371 25189 12391 25219
rect 12429 25189 12439 25219
rect 12439 25189 12463 25219
rect 12501 25189 12507 25219
rect 12507 25189 12535 25219
rect 12573 25189 12575 25219
rect 12575 25189 12607 25219
rect 12645 25189 12677 25219
rect 12677 25189 12679 25219
rect 12717 25189 12745 25219
rect 12745 25189 12751 25219
rect 12789 25189 12813 25219
rect 12813 25189 12823 25219
rect 12861 25189 12881 25219
rect 12881 25189 12895 25219
rect 12933 25189 12949 25219
rect 12949 25189 12967 25219
rect 13005 25189 13017 25219
rect 13017 25189 13039 25219
rect 13077 25189 13085 25219
rect 13085 25189 13111 25219
rect 13149 25189 13153 25219
rect 13153 25189 13183 25219
rect 13221 25189 13255 25223
rect 13293 25219 13327 25223
rect 13365 25219 13399 25223
rect 13437 25219 13471 25223
rect 13509 25219 13543 25223
rect 13581 25219 13615 25223
rect 13653 25219 13687 25223
rect 13293 25189 13323 25219
rect 13323 25189 13327 25219
rect 13365 25189 13391 25219
rect 13391 25189 13399 25219
rect 13437 25189 13459 25219
rect 13459 25189 13471 25219
rect 13509 25189 13527 25219
rect 13527 25189 13543 25219
rect 13581 25189 13595 25219
rect 13595 25189 13615 25219
rect 13653 25189 13663 25219
rect 13663 25189 13687 25219
rect 13756 25185 13765 25215
rect 13765 25185 13790 25215
rect 13828 25185 13833 25215
rect 13833 25185 13862 25215
rect 13900 25185 13901 25215
rect 13901 25185 13934 25215
rect 13972 25185 14003 25215
rect 14003 25185 14006 25215
rect 14044 25185 14071 25215
rect 14071 25185 14078 25215
rect 14116 25185 14139 25215
rect 14139 25185 14150 25215
rect 14252 25207 14286 25241
rect 14324 25207 14358 25241
rect 13756 25181 13790 25185
rect 13828 25181 13862 25185
rect 13900 25181 13934 25185
rect 13972 25181 14006 25185
rect 14044 25181 14078 25185
rect 14116 25181 14150 25185
rect 9909 25149 9943 25150
rect 9981 25149 10015 25150
rect 10053 25149 10087 25150
rect 10125 25149 10159 25150
rect 10197 25149 10231 25150
rect 10269 25149 10303 25150
rect 10341 25149 10375 25150
rect 10413 25149 10447 25150
rect 10485 25149 10519 25150
rect 10557 25149 10591 25150
rect 10629 25149 10663 25150
rect 10701 25149 10735 25150
rect 9909 25116 9911 25149
rect 9911 25116 9943 25149
rect 9981 25116 10014 25149
rect 10014 25116 10015 25149
rect 10053 25116 10083 25149
rect 10083 25116 10087 25149
rect 10125 25116 10152 25149
rect 10152 25116 10159 25149
rect 10197 25116 10221 25149
rect 10221 25116 10231 25149
rect 10269 25116 10290 25149
rect 10290 25116 10303 25149
rect 10341 25116 10359 25149
rect 10359 25116 10375 25149
rect 10413 25116 10428 25149
rect 10428 25116 10447 25149
rect 10485 25116 10497 25149
rect 10497 25116 10519 25149
rect 10557 25116 10566 25149
rect 10566 25116 10591 25149
rect 10629 25116 10635 25149
rect 10635 25116 10663 25149
rect 10701 25116 10704 25149
rect 10704 25116 10735 25149
rect 10773 25116 10807 25150
rect 10845 25149 10879 25150
rect 10917 25149 10951 25150
rect 10989 25149 11023 25150
rect 11061 25149 11095 25150
rect 11133 25149 11167 25150
rect 11205 25149 11239 25150
rect 11277 25149 11311 25150
rect 11349 25149 11383 25150
rect 11421 25149 11455 25150
rect 11493 25149 11527 25150
rect 11565 25149 11599 25150
rect 11637 25149 11671 25150
rect 11709 25149 11743 25150
rect 11781 25149 11815 25150
rect 11853 25149 11887 25150
rect 11925 25149 11959 25150
rect 10845 25116 10875 25149
rect 10875 25116 10879 25149
rect 10917 25116 10943 25149
rect 10943 25116 10951 25149
rect 10989 25116 11011 25149
rect 11011 25116 11023 25149
rect 11061 25116 11079 25149
rect 11079 25116 11095 25149
rect 11133 25116 11147 25149
rect 11147 25116 11167 25149
rect 11205 25116 11215 25149
rect 11215 25116 11239 25149
rect 11277 25116 11283 25149
rect 11283 25116 11311 25149
rect 11349 25116 11351 25149
rect 11351 25116 11383 25149
rect 11421 25116 11453 25149
rect 11453 25116 11455 25149
rect 11493 25116 11521 25149
rect 11521 25116 11527 25149
rect 11565 25116 11589 25149
rect 11589 25116 11599 25149
rect 11637 25116 11657 25149
rect 11657 25116 11671 25149
rect 11709 25116 11725 25149
rect 11725 25116 11743 25149
rect 11781 25116 11793 25149
rect 11793 25116 11815 25149
rect 11853 25116 11861 25149
rect 11861 25116 11887 25149
rect 11925 25116 11929 25149
rect 11929 25116 11959 25149
rect 11997 25116 12031 25150
rect 12069 25149 12103 25150
rect 12141 25149 12175 25150
rect 12213 25149 12247 25150
rect 12285 25149 12319 25150
rect 12357 25149 12391 25150
rect 12429 25149 12463 25150
rect 12501 25149 12535 25150
rect 12573 25149 12607 25150
rect 12645 25149 12679 25150
rect 12717 25149 12751 25150
rect 12789 25149 12823 25150
rect 12861 25149 12895 25150
rect 12933 25149 12967 25150
rect 13005 25149 13039 25150
rect 13077 25149 13111 25150
rect 13149 25149 13183 25150
rect 12069 25116 12099 25149
rect 12099 25116 12103 25149
rect 12141 25116 12167 25149
rect 12167 25116 12175 25149
rect 12213 25116 12235 25149
rect 12235 25116 12247 25149
rect 12285 25116 12303 25149
rect 12303 25116 12319 25149
rect 12357 25116 12371 25149
rect 12371 25116 12391 25149
rect 12429 25116 12439 25149
rect 12439 25116 12463 25149
rect 12501 25116 12507 25149
rect 12507 25116 12535 25149
rect 12573 25116 12575 25149
rect 12575 25116 12607 25149
rect 12645 25116 12677 25149
rect 12677 25116 12679 25149
rect 12717 25116 12745 25149
rect 12745 25116 12751 25149
rect 12789 25116 12813 25149
rect 12813 25116 12823 25149
rect 12861 25116 12881 25149
rect 12881 25116 12895 25149
rect 12933 25116 12949 25149
rect 12949 25116 12967 25149
rect 13005 25116 13017 25149
rect 13017 25116 13039 25149
rect 13077 25116 13085 25149
rect 13085 25116 13111 25149
rect 13149 25116 13153 25149
rect 13153 25116 13183 25149
rect 13221 25116 13255 25150
rect 13293 25149 13327 25150
rect 13365 25149 13399 25150
rect 13437 25149 13471 25150
rect 13509 25149 13543 25150
rect 13581 25149 13615 25150
rect 13653 25149 13687 25150
rect 13293 25116 13323 25149
rect 13323 25116 13327 25149
rect 13365 25116 13391 25149
rect 13391 25116 13399 25149
rect 13437 25116 13459 25149
rect 13459 25116 13471 25149
rect 13509 25116 13527 25149
rect 13527 25116 13543 25149
rect 13581 25116 13595 25149
rect 13595 25116 13615 25149
rect 13653 25116 13663 25149
rect 13663 25116 13687 25149
rect 13756 25115 13765 25141
rect 13765 25115 13790 25141
rect 13828 25115 13833 25141
rect 13833 25115 13862 25141
rect 13900 25115 13901 25141
rect 13901 25115 13934 25141
rect 13972 25115 14003 25141
rect 14003 25115 14006 25141
rect 14044 25115 14071 25141
rect 14071 25115 14078 25141
rect 14116 25115 14139 25141
rect 14139 25115 14150 25141
rect 14252 25134 14286 25168
rect 14324 25134 14358 25168
rect 13756 25107 13790 25115
rect 13828 25107 13862 25115
rect 13900 25107 13934 25115
rect 13972 25107 14006 25115
rect 14044 25107 14078 25115
rect 14116 25107 14150 25115
rect 13756 25045 13765 25067
rect 13765 25045 13790 25067
rect 13828 25045 13833 25067
rect 13833 25045 13862 25067
rect 13900 25045 13901 25067
rect 13901 25045 13934 25067
rect 13972 25045 14003 25067
rect 14003 25045 14006 25067
rect 14044 25045 14071 25067
rect 14071 25045 14078 25067
rect 14116 25045 14139 25067
rect 14139 25045 14150 25067
rect 14252 25061 14286 25095
rect 14324 25061 14358 25095
rect 13756 25033 13790 25045
rect 13828 25033 13862 25045
rect 13900 25033 13934 25045
rect 13972 25033 14006 25045
rect 14044 25033 14078 25045
rect 14116 25033 14150 25045
rect 14252 24988 14286 25022
rect 14324 24988 14358 25022
rect 14252 24915 14286 24949
rect 14324 24915 14358 24949
rect 14252 24842 14286 24876
rect 14324 24842 14358 24876
rect 9914 24549 9948 24562
rect 9990 24549 10024 24562
rect 10066 24549 10100 24562
rect 10142 24549 10176 24562
rect 10218 24549 10252 24562
rect 10294 24549 10328 24562
rect 10369 24549 10403 24562
rect 10444 24549 10478 24562
rect 10519 24549 10553 24562
rect 10594 24549 10628 24562
rect 10669 24549 10703 24562
rect 10744 24549 10778 24562
rect 10819 24549 10853 24562
rect 10894 24549 10928 24562
rect 10969 24549 11003 24562
rect 11044 24549 11078 24562
rect 11119 24549 11153 24562
rect 11194 24549 11228 24562
rect 9914 24528 9945 24549
rect 9945 24528 9948 24549
rect 9990 24528 10015 24549
rect 10015 24528 10024 24549
rect 10066 24528 10085 24549
rect 10085 24528 10100 24549
rect 10142 24528 10155 24549
rect 10155 24528 10176 24549
rect 10218 24528 10225 24549
rect 10225 24528 10252 24549
rect 10294 24528 10295 24549
rect 10295 24528 10328 24549
rect 10369 24528 10401 24549
rect 10401 24528 10403 24549
rect 10444 24528 10471 24549
rect 10471 24528 10478 24549
rect 10519 24528 10541 24549
rect 10541 24528 10553 24549
rect 10594 24528 10611 24549
rect 10611 24528 10628 24549
rect 10669 24528 10681 24549
rect 10681 24528 10703 24549
rect 10744 24528 10750 24549
rect 10750 24528 10778 24549
rect 10819 24528 10853 24549
rect 10894 24528 10922 24549
rect 10922 24528 10928 24549
rect 10969 24528 10991 24549
rect 10991 24528 11003 24549
rect 11044 24528 11060 24549
rect 11060 24528 11078 24549
rect 11119 24528 11129 24549
rect 11129 24528 11153 24549
rect 11194 24528 11198 24549
rect 11198 24528 11228 24549
rect 9914 24481 9948 24490
rect 9990 24481 10024 24490
rect 10066 24481 10100 24490
rect 10142 24481 10176 24490
rect 10218 24481 10252 24490
rect 10294 24481 10328 24490
rect 10369 24481 10403 24490
rect 10444 24481 10478 24490
rect 10519 24481 10553 24490
rect 10594 24481 10628 24490
rect 10669 24481 10703 24490
rect 10744 24481 10778 24490
rect 10819 24481 10853 24490
rect 10894 24481 10928 24490
rect 10969 24481 11003 24490
rect 11044 24481 11078 24490
rect 11119 24481 11153 24490
rect 11194 24481 11228 24490
rect 9914 24456 9945 24481
rect 9945 24456 9948 24481
rect 9990 24456 10015 24481
rect 10015 24456 10024 24481
rect 10066 24456 10085 24481
rect 10085 24456 10100 24481
rect 10142 24456 10155 24481
rect 10155 24456 10176 24481
rect 10218 24456 10225 24481
rect 10225 24456 10252 24481
rect 10294 24456 10295 24481
rect 10295 24456 10328 24481
rect 10369 24456 10401 24481
rect 10401 24456 10403 24481
rect 10444 24456 10471 24481
rect 10471 24456 10478 24481
rect 10519 24456 10541 24481
rect 10541 24456 10553 24481
rect 10594 24456 10611 24481
rect 10611 24456 10628 24481
rect 10669 24456 10681 24481
rect 10681 24456 10703 24481
rect 10744 24456 10750 24481
rect 10750 24456 10778 24481
rect 10819 24456 10853 24481
rect 10894 24456 10922 24481
rect 10922 24456 10928 24481
rect 10969 24456 10991 24481
rect 10991 24456 11003 24481
rect 11044 24456 11060 24481
rect 11060 24456 11078 24481
rect 11119 24456 11129 24481
rect 11129 24456 11153 24481
rect 11194 24456 11198 24481
rect 11198 24456 11228 24481
rect 9914 24413 9948 24418
rect 9990 24413 10024 24418
rect 10066 24413 10100 24418
rect 10142 24413 10176 24418
rect 10218 24413 10252 24418
rect 10294 24413 10328 24418
rect 10369 24413 10403 24418
rect 10444 24413 10478 24418
rect 10519 24413 10553 24418
rect 10594 24413 10628 24418
rect 10669 24413 10703 24418
rect 10744 24413 10778 24418
rect 10819 24413 10853 24418
rect 10894 24413 10928 24418
rect 10969 24413 11003 24418
rect 11044 24413 11078 24418
rect 11119 24413 11153 24418
rect 11194 24413 11228 24418
rect 9914 24384 9945 24413
rect 9945 24384 9948 24413
rect 9990 24384 10015 24413
rect 10015 24384 10024 24413
rect 10066 24384 10085 24413
rect 10085 24384 10100 24413
rect 10142 24384 10155 24413
rect 10155 24384 10176 24413
rect 10218 24384 10225 24413
rect 10225 24384 10252 24413
rect 10294 24384 10295 24413
rect 10295 24384 10328 24413
rect 10369 24384 10401 24413
rect 10401 24384 10403 24413
rect 10444 24384 10471 24413
rect 10471 24384 10478 24413
rect 10519 24384 10541 24413
rect 10541 24384 10553 24413
rect 10594 24384 10611 24413
rect 10611 24384 10628 24413
rect 10669 24384 10681 24413
rect 10681 24384 10703 24413
rect 10744 24384 10750 24413
rect 10750 24384 10778 24413
rect 10819 24384 10853 24413
rect 10894 24384 10922 24413
rect 10922 24384 10928 24413
rect 10969 24384 10991 24413
rect 10991 24384 11003 24413
rect 11044 24384 11060 24413
rect 11060 24384 11078 24413
rect 11119 24384 11129 24413
rect 11129 24384 11153 24413
rect 11194 24384 11198 24413
rect 11198 24384 11228 24413
rect 9914 24345 9948 24346
rect 9990 24345 10024 24346
rect 10066 24345 10100 24346
rect 10142 24345 10176 24346
rect 10218 24345 10252 24346
rect 10294 24345 10328 24346
rect 10369 24345 10403 24346
rect 10444 24345 10478 24346
rect 10519 24345 10553 24346
rect 10594 24345 10628 24346
rect 10669 24345 10703 24346
rect 10744 24345 10778 24346
rect 10819 24345 10853 24346
rect 10894 24345 10928 24346
rect 10969 24345 11003 24346
rect 11044 24345 11078 24346
rect 11119 24345 11153 24346
rect 11194 24345 11228 24346
rect 9914 24312 9945 24345
rect 9945 24312 9948 24345
rect 9990 24312 10015 24345
rect 10015 24312 10024 24345
rect 10066 24312 10085 24345
rect 10085 24312 10100 24345
rect 10142 24312 10155 24345
rect 10155 24312 10176 24345
rect 10218 24312 10225 24345
rect 10225 24312 10252 24345
rect 10294 24312 10295 24345
rect 10295 24312 10328 24345
rect 10369 24312 10401 24345
rect 10401 24312 10403 24345
rect 10444 24312 10471 24345
rect 10471 24312 10478 24345
rect 10519 24312 10541 24345
rect 10541 24312 10553 24345
rect 10594 24312 10611 24345
rect 10611 24312 10628 24345
rect 10669 24312 10681 24345
rect 10681 24312 10703 24345
rect 10744 24312 10750 24345
rect 10750 24312 10778 24345
rect 10819 24312 10853 24345
rect 10894 24312 10922 24345
rect 10922 24312 10928 24345
rect 10969 24312 10991 24345
rect 10991 24312 11003 24345
rect 11044 24312 11060 24345
rect 11060 24312 11078 24345
rect 11119 24312 11129 24345
rect 11129 24312 11153 24345
rect 11194 24312 11198 24345
rect 11198 24312 11228 24345
rect 9914 24243 9945 24274
rect 9945 24243 9948 24274
rect 9990 24243 10015 24274
rect 10015 24243 10024 24274
rect 10066 24243 10085 24274
rect 10085 24243 10100 24274
rect 10142 24243 10155 24274
rect 10155 24243 10176 24274
rect 10218 24243 10225 24274
rect 10225 24243 10252 24274
rect 10294 24243 10295 24274
rect 10295 24243 10328 24274
rect 10369 24243 10401 24274
rect 10401 24243 10403 24274
rect 10444 24243 10471 24274
rect 10471 24243 10478 24274
rect 10519 24243 10541 24274
rect 10541 24243 10553 24274
rect 10594 24243 10611 24274
rect 10611 24243 10628 24274
rect 10669 24243 10681 24274
rect 10681 24243 10703 24274
rect 10744 24243 10750 24274
rect 10750 24243 10778 24274
rect 10819 24243 10853 24274
rect 10894 24243 10922 24274
rect 10922 24243 10928 24274
rect 10969 24243 10991 24274
rect 10991 24243 11003 24274
rect 11044 24243 11060 24274
rect 11060 24243 11078 24274
rect 11119 24243 11129 24274
rect 11129 24243 11153 24274
rect 11194 24243 11198 24274
rect 11198 24243 11228 24274
rect 9914 24240 9948 24243
rect 9990 24240 10024 24243
rect 10066 24240 10100 24243
rect 10142 24240 10176 24243
rect 10218 24240 10252 24243
rect 10294 24240 10328 24243
rect 10369 24240 10403 24243
rect 10444 24240 10478 24243
rect 10519 24240 10553 24243
rect 10594 24240 10628 24243
rect 10669 24240 10703 24243
rect 10744 24240 10778 24243
rect 10819 24240 10853 24243
rect 10894 24240 10928 24243
rect 10969 24240 11003 24243
rect 11044 24240 11078 24243
rect 11119 24240 11153 24243
rect 11194 24240 11228 24243
rect 9905 24142 9914 24171
rect 9914 24142 9939 24171
rect 9981 24142 9984 24171
rect 9984 24142 10015 24171
rect 10057 24142 10088 24171
rect 10088 24142 10091 24171
rect 10133 24142 10158 24171
rect 10158 24142 10167 24171
rect 10209 24142 10228 24171
rect 10228 24142 10243 24171
rect 10285 24142 10298 24171
rect 10298 24142 10319 24171
rect 10361 24142 10368 24171
rect 10368 24142 10395 24171
rect 10437 24142 10438 24171
rect 10438 24142 10471 24171
rect 10513 24142 10544 24171
rect 10544 24142 10547 24171
rect 10589 24142 10614 24171
rect 10614 24142 10623 24171
rect 10665 24142 10684 24171
rect 10684 24142 10699 24171
rect 9905 24137 9939 24142
rect 9981 24137 10015 24142
rect 10057 24137 10091 24142
rect 10133 24137 10167 24142
rect 10209 24137 10243 24142
rect 10285 24137 10319 24142
rect 10361 24137 10395 24142
rect 10437 24137 10471 24142
rect 10513 24137 10547 24142
rect 10589 24137 10623 24142
rect 10665 24137 10699 24142
rect 9905 24074 9914 24097
rect 9914 24074 9939 24097
rect 9981 24074 9984 24097
rect 9984 24074 10015 24097
rect 10057 24074 10088 24097
rect 10088 24074 10091 24097
rect 10133 24074 10158 24097
rect 10158 24074 10167 24097
rect 10209 24074 10228 24097
rect 10228 24074 10243 24097
rect 10285 24074 10298 24097
rect 10298 24074 10319 24097
rect 10361 24074 10368 24097
rect 10368 24074 10395 24097
rect 10437 24074 10438 24097
rect 10438 24074 10471 24097
rect 10513 24074 10544 24097
rect 10544 24074 10547 24097
rect 10589 24074 10614 24097
rect 10614 24074 10623 24097
rect 10665 24074 10684 24097
rect 10684 24074 10699 24097
rect 9905 24063 9939 24074
rect 9981 24063 10015 24074
rect 10057 24063 10091 24074
rect 10133 24063 10167 24074
rect 10209 24063 10243 24074
rect 10285 24063 10319 24074
rect 10361 24063 10395 24074
rect 10437 24063 10471 24074
rect 10513 24063 10547 24074
rect 10589 24063 10623 24074
rect 10665 24063 10699 24074
rect 9905 24006 9914 24023
rect 9914 24006 9939 24023
rect 9981 24006 9984 24023
rect 9984 24006 10015 24023
rect 10057 24006 10088 24023
rect 10088 24006 10091 24023
rect 10133 24006 10158 24023
rect 10158 24006 10167 24023
rect 10209 24006 10228 24023
rect 10228 24006 10243 24023
rect 10285 24006 10298 24023
rect 10298 24006 10319 24023
rect 10361 24006 10368 24023
rect 10368 24006 10395 24023
rect 10437 24006 10438 24023
rect 10438 24006 10471 24023
rect 10513 24006 10544 24023
rect 10544 24006 10547 24023
rect 10589 24006 10614 24023
rect 10614 24006 10623 24023
rect 10665 24006 10684 24023
rect 10684 24006 10699 24023
rect 9905 23989 9939 24006
rect 9981 23989 10015 24006
rect 10057 23989 10091 24006
rect 10133 23989 10167 24006
rect 10209 23989 10243 24006
rect 10285 23989 10319 24006
rect 10361 23989 10395 24006
rect 10437 23989 10471 24006
rect 10513 23989 10547 24006
rect 10589 23989 10623 24006
rect 10665 23989 10699 24006
rect 9905 23937 9914 23949
rect 9914 23937 9939 23949
rect 9981 23937 9984 23949
rect 9984 23937 10015 23949
rect 10057 23937 10088 23949
rect 10088 23937 10091 23949
rect 10133 23937 10158 23949
rect 10158 23937 10167 23949
rect 10209 23937 10228 23949
rect 10228 23937 10243 23949
rect 10285 23937 10298 23949
rect 10298 23937 10319 23949
rect 10361 23937 10368 23949
rect 10368 23937 10395 23949
rect 10437 23937 10438 23949
rect 10438 23937 10471 23949
rect 10513 23937 10544 23949
rect 10544 23937 10547 23949
rect 10589 23937 10614 23949
rect 10614 23937 10623 23949
rect 10665 23937 10684 23949
rect 10684 23937 10699 23949
rect 9905 23915 9939 23937
rect 9981 23915 10015 23937
rect 10057 23915 10091 23937
rect 10133 23915 10167 23937
rect 10209 23915 10243 23937
rect 10285 23915 10319 23937
rect 10361 23915 10395 23937
rect 10437 23915 10471 23937
rect 10513 23915 10547 23937
rect 10589 23915 10623 23937
rect 10665 23915 10699 23937
rect 9905 23868 9914 23875
rect 9914 23868 9939 23875
rect 9981 23868 9984 23875
rect 9984 23868 10015 23875
rect 10057 23868 10088 23875
rect 10088 23868 10091 23875
rect 10133 23868 10158 23875
rect 10158 23868 10167 23875
rect 10209 23868 10228 23875
rect 10228 23868 10243 23875
rect 10285 23868 10298 23875
rect 10298 23868 10319 23875
rect 10361 23868 10368 23875
rect 10368 23868 10395 23875
rect 10437 23868 10438 23875
rect 10438 23868 10471 23875
rect 10513 23868 10544 23875
rect 10544 23868 10547 23875
rect 10589 23868 10614 23875
rect 10614 23868 10623 23875
rect 10665 23868 10684 23875
rect 10684 23868 10699 23875
rect 9905 23841 9939 23868
rect 9981 23841 10015 23868
rect 10057 23841 10091 23868
rect 10133 23841 10167 23868
rect 10209 23841 10243 23868
rect 10285 23841 10319 23868
rect 10361 23841 10395 23868
rect 10437 23841 10471 23868
rect 10513 23841 10547 23868
rect 10589 23841 10623 23868
rect 10665 23841 10699 23868
rect 9905 23799 9914 23801
rect 9914 23799 9939 23801
rect 9981 23799 9984 23801
rect 9984 23799 10015 23801
rect 10057 23799 10088 23801
rect 10088 23799 10091 23801
rect 10133 23799 10158 23801
rect 10158 23799 10167 23801
rect 10209 23799 10228 23801
rect 10228 23799 10243 23801
rect 10285 23799 10298 23801
rect 10298 23799 10319 23801
rect 10361 23799 10368 23801
rect 10368 23799 10395 23801
rect 10437 23799 10438 23801
rect 10438 23799 10471 23801
rect 10513 23799 10544 23801
rect 10544 23799 10547 23801
rect 10589 23799 10614 23801
rect 10614 23799 10623 23801
rect 10665 23799 10684 23801
rect 10684 23799 10699 23801
rect 9905 23767 9939 23799
rect 9981 23767 10015 23799
rect 10057 23767 10091 23799
rect 10133 23767 10167 23799
rect 10209 23767 10243 23799
rect 10285 23767 10319 23799
rect 10361 23767 10395 23799
rect 10437 23767 10471 23799
rect 10513 23767 10547 23799
rect 10589 23767 10623 23799
rect 10665 23767 10699 23799
rect 9905 23695 9939 23727
rect 9981 23695 10015 23727
rect 10057 23695 10091 23727
rect 10133 23695 10167 23727
rect 10209 23695 10243 23727
rect 10285 23695 10319 23727
rect 10361 23695 10395 23727
rect 10437 23695 10471 23727
rect 10513 23695 10547 23727
rect 10589 23695 10623 23727
rect 10665 23695 10699 23727
rect 9905 23693 9914 23695
rect 9914 23693 9939 23695
rect 9981 23693 9984 23695
rect 9984 23693 10015 23695
rect 10057 23693 10088 23695
rect 10088 23693 10091 23695
rect 10133 23693 10158 23695
rect 10158 23693 10167 23695
rect 10209 23693 10228 23695
rect 10228 23693 10243 23695
rect 10285 23693 10298 23695
rect 10298 23693 10319 23695
rect 10361 23693 10368 23695
rect 10368 23693 10395 23695
rect 10437 23693 10438 23695
rect 10438 23693 10471 23695
rect 10513 23693 10544 23695
rect 10544 23693 10547 23695
rect 10589 23693 10614 23695
rect 10614 23693 10623 23695
rect 10665 23693 10684 23695
rect 10684 23693 10699 23695
rect 9905 23626 9939 23653
rect 9981 23626 10015 23653
rect 10057 23626 10091 23653
rect 10133 23626 10167 23653
rect 10209 23626 10243 23653
rect 10285 23626 10319 23653
rect 10361 23626 10395 23653
rect 10437 23626 10471 23653
rect 10513 23626 10547 23653
rect 10589 23626 10623 23653
rect 10665 23626 10699 23653
rect 9905 23619 9914 23626
rect 9914 23619 9939 23626
rect 9981 23619 9984 23626
rect 9984 23619 10015 23626
rect 10057 23619 10088 23626
rect 10088 23619 10091 23626
rect 10133 23619 10158 23626
rect 10158 23619 10167 23626
rect 10209 23619 10228 23626
rect 10228 23619 10243 23626
rect 10285 23619 10298 23626
rect 10298 23619 10319 23626
rect 10361 23619 10368 23626
rect 10368 23619 10395 23626
rect 10437 23619 10438 23626
rect 10438 23619 10471 23626
rect 10513 23619 10544 23626
rect 10544 23619 10547 23626
rect 10589 23619 10614 23626
rect 10614 23619 10623 23626
rect 10665 23619 10684 23626
rect 10684 23619 10699 23626
rect 9905 23557 9939 23579
rect 9981 23557 10015 23579
rect 10057 23557 10091 23579
rect 10133 23557 10167 23579
rect 10209 23557 10243 23579
rect 10285 23557 10319 23579
rect 10361 23557 10395 23579
rect 10437 23557 10471 23579
rect 10513 23557 10547 23579
rect 10589 23557 10623 23579
rect 10665 23557 10699 23579
rect 9905 23545 9914 23557
rect 9914 23545 9939 23557
rect 9981 23545 9984 23557
rect 9984 23545 10015 23557
rect 10057 23545 10088 23557
rect 10088 23545 10091 23557
rect 10133 23545 10158 23557
rect 10158 23545 10167 23557
rect 10209 23545 10228 23557
rect 10228 23545 10243 23557
rect 10285 23545 10298 23557
rect 10298 23545 10319 23557
rect 10361 23545 10368 23557
rect 10368 23545 10395 23557
rect 10437 23545 10438 23557
rect 10438 23545 10471 23557
rect 10513 23545 10544 23557
rect 10544 23545 10547 23557
rect 10589 23545 10614 23557
rect 10614 23545 10623 23557
rect 10665 23545 10684 23557
rect 10684 23545 10699 23557
rect 9905 23488 9939 23505
rect 9981 23488 10015 23505
rect 10057 23488 10091 23505
rect 10133 23488 10167 23505
rect 10209 23488 10243 23505
rect 10285 23488 10319 23505
rect 10361 23488 10395 23505
rect 10437 23488 10471 23505
rect 10513 23488 10547 23505
rect 10589 23488 10623 23505
rect 10665 23488 10699 23505
rect 9905 23471 9914 23488
rect 9914 23471 9939 23488
rect 9981 23471 9984 23488
rect 9984 23471 10015 23488
rect 10057 23471 10088 23488
rect 10088 23471 10091 23488
rect 10133 23471 10158 23488
rect 10158 23471 10167 23488
rect 10209 23471 10228 23488
rect 10228 23471 10243 23488
rect 10285 23471 10298 23488
rect 10298 23471 10319 23488
rect 10361 23471 10368 23488
rect 10368 23471 10395 23488
rect 10437 23471 10438 23488
rect 10438 23471 10471 23488
rect 10513 23471 10544 23488
rect 10544 23471 10547 23488
rect 10589 23471 10614 23488
rect 10614 23471 10623 23488
rect 10665 23471 10684 23488
rect 10684 23471 10699 23488
rect 9905 23419 9939 23431
rect 9981 23419 10015 23431
rect 10057 23419 10091 23431
rect 10133 23419 10167 23431
rect 10209 23419 10243 23431
rect 10285 23419 10319 23431
rect 10361 23419 10395 23431
rect 10437 23419 10471 23431
rect 10513 23419 10547 23431
rect 10589 23419 10623 23431
rect 10665 23419 10699 23431
rect 9905 23397 9914 23419
rect 9914 23397 9939 23419
rect 9981 23397 9984 23419
rect 9984 23397 10015 23419
rect 10057 23397 10088 23419
rect 10088 23397 10091 23419
rect 10133 23397 10158 23419
rect 10158 23397 10167 23419
rect 10209 23397 10228 23419
rect 10228 23397 10243 23419
rect 10285 23397 10298 23419
rect 10298 23397 10319 23419
rect 10361 23397 10368 23419
rect 10368 23397 10395 23419
rect 10437 23397 10438 23419
rect 10438 23397 10471 23419
rect 10513 23397 10544 23419
rect 10544 23397 10547 23419
rect 10589 23397 10614 23419
rect 10614 23397 10623 23419
rect 10665 23397 10684 23419
rect 10684 23397 10699 23419
rect 9905 23350 9939 23357
rect 9981 23350 10015 23357
rect 10057 23350 10091 23357
rect 10133 23350 10167 23357
rect 10209 23350 10243 23357
rect 10285 23350 10319 23357
rect 10361 23350 10395 23357
rect 10437 23350 10471 23357
rect 10513 23350 10547 23357
rect 10589 23350 10623 23357
rect 10665 23350 10699 23357
rect 9905 23323 9914 23350
rect 9914 23323 9939 23350
rect 9981 23323 9984 23350
rect 9984 23323 10015 23350
rect 10057 23323 10088 23350
rect 10088 23323 10091 23350
rect 10133 23323 10158 23350
rect 10158 23323 10167 23350
rect 10209 23323 10228 23350
rect 10228 23323 10243 23350
rect 10285 23323 10298 23350
rect 10298 23323 10319 23350
rect 10361 23323 10368 23350
rect 10368 23323 10395 23350
rect 10437 23323 10438 23350
rect 10438 23323 10471 23350
rect 10513 23323 10544 23350
rect 10544 23323 10547 23350
rect 10589 23323 10614 23350
rect 10614 23323 10623 23350
rect 10665 23323 10684 23350
rect 10684 23323 10699 23350
rect 9905 23281 9939 23283
rect 9981 23281 10015 23283
rect 10057 23281 10091 23283
rect 10133 23281 10167 23283
rect 10209 23281 10243 23283
rect 10285 23281 10319 23283
rect 10361 23281 10395 23283
rect 10437 23281 10471 23283
rect 10513 23281 10547 23283
rect 10589 23281 10623 23283
rect 10665 23281 10699 23283
rect 9905 23249 9914 23281
rect 9914 23249 9939 23281
rect 9981 23249 9984 23281
rect 9984 23249 10015 23281
rect 10057 23249 10088 23281
rect 10088 23249 10091 23281
rect 10133 23249 10158 23281
rect 10158 23249 10167 23281
rect 10209 23249 10228 23281
rect 10228 23249 10243 23281
rect 10285 23249 10298 23281
rect 10298 23249 10319 23281
rect 10361 23249 10368 23281
rect 10368 23249 10395 23281
rect 10437 23249 10438 23281
rect 10438 23249 10471 23281
rect 10513 23249 10544 23281
rect 10544 23249 10547 23281
rect 10589 23249 10614 23281
rect 10614 23249 10623 23281
rect 10665 23249 10684 23281
rect 10684 23249 10699 23281
rect 9905 23178 9914 23209
rect 9914 23178 9939 23209
rect 9981 23178 9984 23209
rect 9984 23178 10015 23209
rect 10057 23178 10088 23209
rect 10088 23178 10091 23209
rect 10133 23178 10158 23209
rect 10158 23178 10167 23209
rect 10209 23178 10228 23209
rect 10228 23178 10243 23209
rect 10285 23178 10298 23209
rect 10298 23178 10319 23209
rect 10361 23178 10368 23209
rect 10368 23178 10395 23209
rect 10437 23178 10438 23209
rect 10438 23178 10471 23209
rect 10513 23178 10544 23209
rect 10544 23178 10547 23209
rect 10589 23178 10614 23209
rect 10614 23178 10623 23209
rect 10665 23178 10684 23209
rect 10684 23178 10699 23209
rect 9905 23175 9939 23178
rect 9981 23175 10015 23178
rect 10057 23175 10091 23178
rect 10133 23175 10167 23178
rect 10209 23175 10243 23178
rect 10285 23175 10319 23178
rect 10361 23175 10395 23178
rect 10437 23175 10471 23178
rect 10513 23175 10547 23178
rect 10589 23175 10623 23178
rect 10665 23175 10699 23178
rect 9905 23109 9914 23135
rect 9914 23109 9939 23135
rect 9981 23109 9984 23135
rect 9984 23109 10015 23135
rect 10057 23109 10088 23135
rect 10088 23109 10091 23135
rect 10133 23109 10158 23135
rect 10158 23109 10167 23135
rect 10209 23109 10228 23135
rect 10228 23109 10243 23135
rect 10285 23109 10298 23135
rect 10298 23109 10319 23135
rect 10361 23109 10368 23135
rect 10368 23109 10395 23135
rect 10437 23109 10438 23135
rect 10438 23109 10471 23135
rect 10513 23109 10544 23135
rect 10544 23109 10547 23135
rect 10589 23109 10614 23135
rect 10614 23109 10623 23135
rect 10665 23109 10684 23135
rect 10684 23109 10699 23135
rect 9905 23101 9939 23109
rect 9981 23101 10015 23109
rect 10057 23101 10091 23109
rect 10133 23101 10167 23109
rect 10209 23101 10243 23109
rect 10285 23101 10319 23109
rect 10361 23101 10395 23109
rect 10437 23101 10471 23109
rect 10513 23101 10547 23109
rect 10589 23101 10623 23109
rect 10665 23101 10699 23109
rect 9905 23040 9914 23061
rect 9914 23040 9939 23061
rect 9981 23040 9984 23061
rect 9984 23040 10015 23061
rect 10057 23040 10088 23061
rect 10088 23040 10091 23061
rect 10133 23040 10158 23061
rect 10158 23040 10167 23061
rect 10209 23040 10228 23061
rect 10228 23040 10243 23061
rect 10285 23040 10298 23061
rect 10298 23040 10319 23061
rect 10361 23040 10368 23061
rect 10368 23040 10395 23061
rect 10437 23040 10438 23061
rect 10438 23040 10471 23061
rect 10513 23040 10544 23061
rect 10544 23040 10547 23061
rect 10589 23040 10614 23061
rect 10614 23040 10623 23061
rect 10665 23040 10684 23061
rect 10684 23040 10699 23061
rect 14252 24769 14286 24803
rect 14324 24769 14358 24803
rect 14252 24696 14286 24730
rect 14324 24696 14358 24730
rect 14252 24623 14286 24657
rect 14324 24623 14358 24657
rect 14252 24550 14286 24584
rect 14324 24550 14358 24584
rect 14252 24477 14286 24511
rect 14324 24477 14358 24511
rect 14252 24404 14286 24438
rect 14324 24404 14358 24438
rect 14252 24331 14286 24365
rect 14324 24331 14358 24365
rect 14252 24258 14286 24292
rect 14324 24258 14358 24292
rect 14252 24185 14286 24219
rect 14324 24185 14358 24219
rect 14252 24115 14286 24146
rect 14324 24115 14358 24146
rect 14252 24112 14267 24115
rect 14267 24112 14286 24115
rect 14324 24112 14335 24115
rect 14335 24112 14358 24115
rect 14252 24046 14286 24073
rect 14324 24046 14358 24073
rect 14252 24039 14267 24046
rect 14267 24039 14286 24046
rect 14324 24039 14335 24046
rect 14335 24039 14358 24046
rect 14252 23977 14286 24000
rect 14324 23977 14358 24000
rect 14252 23966 14267 23977
rect 14267 23966 14286 23977
rect 14324 23966 14335 23977
rect 14335 23966 14358 23977
rect 14252 23908 14286 23927
rect 14324 23908 14358 23927
rect 14252 23893 14267 23908
rect 14267 23893 14286 23908
rect 14324 23893 14335 23908
rect 14335 23893 14358 23908
rect 14252 23839 14286 23854
rect 14324 23839 14358 23854
rect 14252 23820 14267 23839
rect 14267 23820 14286 23839
rect 14324 23820 14335 23839
rect 14335 23820 14358 23839
rect 14252 23770 14286 23781
rect 14324 23770 14358 23781
rect 14252 23747 14267 23770
rect 14267 23747 14286 23770
rect 14324 23747 14335 23770
rect 14335 23747 14358 23770
rect 14252 23701 14286 23708
rect 14324 23701 14358 23708
rect 14252 23674 14267 23701
rect 14267 23674 14286 23701
rect 14324 23674 14335 23701
rect 14335 23674 14358 23701
rect 14252 23632 14286 23635
rect 14324 23632 14358 23635
rect 14252 23601 14267 23632
rect 14267 23601 14286 23632
rect 14324 23601 14335 23632
rect 14335 23601 14358 23632
rect 14252 23529 14267 23562
rect 14267 23529 14286 23562
rect 14324 23529 14335 23562
rect 14335 23529 14358 23562
rect 14252 23528 14286 23529
rect 14324 23528 14358 23529
rect 14252 23460 14267 23489
rect 14267 23460 14286 23489
rect 14324 23460 14335 23489
rect 14335 23460 14358 23489
rect 14252 23455 14286 23460
rect 14324 23455 14358 23460
rect 14252 23391 14267 23416
rect 14267 23391 14286 23416
rect 14324 23391 14335 23416
rect 14335 23391 14358 23416
rect 14252 23382 14286 23391
rect 14324 23382 14358 23391
rect 14252 23322 14267 23343
rect 14267 23322 14286 23343
rect 14324 23322 14335 23343
rect 14335 23322 14358 23343
rect 14252 23309 14286 23322
rect 14324 23309 14358 23322
rect 14252 23253 14267 23270
rect 14267 23253 14286 23270
rect 14324 23253 14335 23270
rect 14335 23253 14358 23270
rect 14252 23236 14286 23253
rect 14324 23236 14358 23253
rect 14252 23184 14267 23197
rect 14267 23184 14286 23197
rect 14324 23184 14335 23197
rect 14335 23184 14358 23197
rect 14252 23163 14286 23184
rect 14324 23163 14358 23184
rect 14252 23115 14267 23124
rect 14267 23115 14286 23124
rect 14324 23115 14335 23124
rect 14335 23115 14358 23124
rect 14252 23090 14286 23115
rect 14324 23090 14358 23115
rect 14252 23046 14267 23051
rect 14267 23046 14286 23051
rect 14324 23046 14335 23051
rect 14335 23046 14358 23051
rect 9905 23027 9939 23040
rect 9981 23027 10015 23040
rect 10057 23027 10091 23040
rect 10133 23027 10167 23040
rect 10209 23027 10243 23040
rect 10285 23027 10319 23040
rect 10361 23027 10395 23040
rect 10437 23027 10471 23040
rect 10513 23027 10547 23040
rect 10589 23027 10623 23040
rect 10665 23027 10699 23040
rect 14252 23017 14286 23046
rect 14324 23017 14358 23046
rect 9905 22971 9914 22987
rect 9914 22971 9939 22987
rect 9981 22971 9984 22987
rect 9984 22971 10015 22987
rect 10057 22971 10088 22987
rect 10088 22971 10091 22987
rect 10133 22971 10158 22987
rect 10158 22971 10167 22987
rect 10209 22971 10228 22987
rect 10228 22971 10243 22987
rect 10285 22971 10298 22987
rect 10298 22971 10319 22987
rect 10361 22971 10368 22987
rect 10368 22971 10395 22987
rect 10437 22971 10438 22987
rect 10438 22971 10471 22987
rect 10513 22971 10544 22987
rect 10544 22971 10547 22987
rect 10589 22971 10614 22987
rect 10614 22971 10623 22987
rect 10665 22971 10684 22987
rect 10684 22971 10699 22987
rect 10759 22971 10788 23000
rect 10788 22971 10793 23000
rect 9905 22953 9939 22971
rect 9981 22953 10015 22971
rect 10057 22953 10091 22971
rect 10133 22953 10167 22971
rect 10209 22953 10243 22971
rect 10285 22953 10319 22971
rect 10361 22953 10395 22971
rect 10437 22953 10471 22971
rect 10513 22953 10547 22971
rect 10589 22953 10623 22971
rect 10665 22953 10699 22971
rect 10759 22966 10793 22971
rect 10832 22969 10859 23000
rect 10859 22969 10866 23000
rect 10905 22969 10928 23000
rect 10928 22969 10939 23000
rect 10978 22969 10997 23000
rect 10997 22969 11012 23000
rect 11051 22969 11066 23000
rect 11066 22969 11085 23000
rect 11124 22969 11135 23000
rect 11135 22969 11158 23000
rect 11197 22969 11204 23000
rect 11204 22969 11231 23000
rect 11270 22969 11273 23000
rect 11273 22969 11304 23000
rect 11343 22969 11376 23000
rect 11376 22969 11377 23000
rect 11416 22969 11445 23000
rect 11445 22969 11450 23000
rect 11489 22969 11514 23000
rect 11514 22969 11523 23000
rect 11562 22969 11583 23000
rect 11583 22969 11596 23000
rect 11635 22969 11652 23000
rect 11652 22969 11669 23000
rect 11707 22969 11721 23000
rect 11721 22969 11741 23000
rect 11779 22969 11790 23000
rect 11790 22969 11813 23000
rect 11851 22969 11859 23000
rect 11859 22969 11885 23000
rect 11923 22969 11928 23000
rect 11928 22969 11957 23000
rect 11995 22969 11997 23000
rect 11997 22969 12029 23000
rect 12067 22969 12099 23000
rect 12099 22969 12101 23000
rect 12139 22969 12167 23000
rect 12167 22969 12173 23000
rect 12211 22969 12235 23000
rect 12235 22969 12245 23000
rect 12476 22969 12507 22984
rect 12507 22969 12510 22984
rect 12550 22969 12575 22984
rect 12575 22969 12584 22984
rect 12624 22969 12643 22984
rect 12643 22969 12658 22984
rect 12698 22969 12711 22984
rect 12711 22969 12732 22984
rect 12772 22969 12779 22984
rect 12779 22969 12806 22984
rect 12846 22969 12847 22984
rect 12847 22969 12880 22984
rect 12920 22969 12949 22984
rect 12949 22969 12954 22984
rect 12994 22969 13017 22984
rect 13017 22969 13028 22984
rect 13068 22969 13085 22984
rect 13085 22969 13102 22984
rect 13141 22969 13153 22984
rect 13153 22969 13175 22984
rect 13214 22969 13221 22984
rect 13221 22969 13248 22984
rect 13287 22969 13289 22984
rect 13289 22969 13321 22984
rect 13360 22969 13391 22984
rect 13391 22969 13394 22984
rect 13433 22969 13459 22984
rect 13459 22969 13467 22984
rect 13506 22969 13527 22984
rect 13527 22969 13540 22984
rect 13579 22969 13595 22984
rect 13595 22969 13613 22984
rect 13652 22969 13663 22984
rect 13663 22969 13686 22984
rect 13756 22969 13765 22999
rect 13765 22969 13790 22999
rect 13828 22969 13833 22999
rect 13833 22969 13862 22999
rect 13900 22969 13901 22999
rect 13901 22969 13934 22999
rect 10832 22966 10866 22969
rect 10905 22966 10939 22969
rect 10978 22966 11012 22969
rect 11051 22966 11085 22969
rect 11124 22966 11158 22969
rect 11197 22966 11231 22969
rect 11270 22966 11304 22969
rect 11343 22966 11377 22969
rect 11416 22966 11450 22969
rect 11489 22966 11523 22969
rect 11562 22966 11596 22969
rect 11635 22966 11669 22969
rect 11707 22966 11741 22969
rect 11779 22966 11813 22969
rect 11851 22966 11885 22969
rect 11923 22966 11957 22969
rect 11995 22966 12029 22969
rect 12067 22966 12101 22969
rect 12139 22966 12173 22969
rect 12211 22966 12245 22969
rect 12476 22950 12510 22969
rect 12550 22950 12584 22969
rect 12624 22950 12658 22969
rect 12698 22950 12732 22969
rect 12772 22950 12806 22969
rect 12846 22950 12880 22969
rect 12920 22950 12954 22969
rect 12994 22950 13028 22969
rect 13068 22950 13102 22969
rect 13141 22950 13175 22969
rect 13214 22950 13248 22969
rect 13287 22950 13321 22969
rect 13360 22950 13394 22969
rect 13433 22950 13467 22969
rect 13506 22950 13540 22969
rect 13579 22950 13613 22969
rect 13652 22950 13686 22969
rect 13756 22965 13790 22969
rect 13828 22965 13862 22969
rect 13900 22965 13934 22969
rect 13972 22998 14006 22999
rect 14044 22998 14078 22999
rect 14116 22998 14150 22999
rect 13972 22965 13978 22998
rect 13978 22965 14006 22998
rect 14044 22965 14048 22998
rect 14048 22965 14078 22998
rect 14116 22965 14118 22998
rect 14118 22965 14150 22998
rect 14252 22977 14267 22978
rect 14267 22977 14286 22978
rect 14324 22977 14335 22978
rect 14335 22977 14358 22978
rect 14252 22944 14286 22977
rect 14324 22944 14358 22977
rect 9905 22901 9935 22913
rect 9935 22901 9939 22913
rect 9981 22901 10005 22913
rect 10005 22901 10015 22913
rect 10057 22901 10075 22913
rect 10075 22901 10091 22913
rect 10133 22901 10145 22913
rect 10145 22901 10167 22913
rect 10209 22901 10215 22913
rect 10215 22901 10243 22913
rect 9905 22879 9939 22901
rect 9981 22879 10015 22901
rect 10057 22879 10091 22901
rect 10133 22879 10167 22901
rect 10209 22879 10243 22901
rect 10285 22879 10319 22913
rect 10361 22901 10391 22913
rect 10391 22901 10395 22913
rect 10437 22901 10461 22913
rect 10461 22901 10471 22913
rect 10513 22901 10530 22913
rect 10530 22901 10547 22913
rect 10589 22901 10599 22913
rect 10599 22901 10623 22913
rect 10665 22901 10668 22913
rect 10668 22901 10699 22913
rect 10759 22901 10771 22914
rect 10771 22901 10793 22914
rect 10832 22901 10840 22914
rect 10840 22901 10866 22914
rect 10905 22901 10909 22914
rect 10909 22901 10939 22914
rect 10361 22879 10395 22901
rect 10437 22879 10471 22901
rect 10513 22879 10547 22901
rect 10589 22879 10623 22901
rect 10665 22879 10699 22901
rect 10759 22880 10793 22901
rect 10832 22880 10866 22901
rect 10905 22880 10939 22901
rect 10978 22880 11012 22914
rect 11051 22901 11082 22914
rect 11082 22901 11085 22914
rect 11124 22901 11151 22914
rect 11151 22901 11158 22914
rect 11197 22901 11220 22914
rect 11220 22901 11231 22914
rect 11270 22901 11289 22914
rect 11289 22901 11304 22914
rect 11343 22901 11358 22914
rect 11358 22901 11377 22914
rect 11416 22901 11427 22914
rect 11427 22901 11450 22914
rect 11489 22901 11496 22914
rect 11496 22901 11523 22914
rect 11562 22901 11565 22914
rect 11565 22901 11596 22914
rect 11635 22901 11668 22914
rect 11668 22901 11669 22914
rect 11707 22901 11737 22914
rect 11737 22901 11741 22914
rect 11779 22901 11806 22914
rect 11806 22901 11813 22914
rect 11851 22901 11875 22914
rect 11875 22901 11885 22914
rect 11923 22901 11944 22914
rect 11944 22901 11957 22914
rect 11995 22901 12013 22914
rect 12013 22901 12029 22914
rect 12067 22901 12082 22914
rect 12082 22901 12101 22914
rect 12139 22901 12151 22914
rect 12151 22901 12173 22914
rect 12211 22901 12220 22914
rect 12220 22901 12245 22914
rect 11051 22880 11085 22901
rect 11124 22880 11158 22901
rect 11197 22880 11231 22901
rect 11270 22880 11304 22901
rect 11343 22880 11377 22901
rect 11416 22880 11450 22901
rect 11489 22880 11523 22901
rect 11562 22880 11596 22901
rect 11635 22880 11669 22901
rect 11707 22880 11741 22901
rect 11779 22880 11813 22901
rect 11851 22880 11885 22901
rect 11923 22880 11957 22901
rect 11995 22880 12029 22901
rect 12067 22880 12101 22901
rect 12139 22880 12173 22901
rect 12211 22880 12245 22901
rect 9905 22831 9935 22839
rect 9935 22831 9939 22839
rect 9981 22831 10005 22839
rect 10005 22831 10015 22839
rect 10057 22831 10075 22839
rect 10075 22831 10091 22839
rect 10133 22831 10145 22839
rect 10145 22831 10167 22839
rect 10209 22831 10215 22839
rect 10215 22831 10243 22839
rect 9905 22805 9939 22831
rect 9981 22805 10015 22831
rect 10057 22805 10091 22831
rect 10133 22805 10167 22831
rect 10209 22805 10243 22831
rect 10285 22805 10319 22839
rect 10361 22831 10391 22839
rect 10391 22831 10395 22839
rect 10437 22831 10461 22839
rect 10461 22831 10471 22839
rect 10513 22831 10530 22839
rect 10530 22831 10547 22839
rect 10589 22831 10599 22839
rect 10599 22831 10623 22839
rect 10665 22831 10668 22839
rect 10668 22831 10699 22839
rect 10361 22805 10395 22831
rect 10437 22805 10471 22831
rect 10513 22805 10547 22831
rect 10589 22805 10623 22831
rect 10665 22805 10699 22831
rect 10759 22795 10793 22828
rect 10832 22795 10866 22828
rect 10905 22795 10939 22828
rect 9905 22761 9935 22765
rect 9935 22761 9939 22765
rect 9981 22761 10005 22765
rect 10005 22761 10015 22765
rect 10057 22761 10075 22765
rect 10075 22761 10091 22765
rect 10133 22761 10145 22765
rect 10145 22761 10167 22765
rect 10209 22761 10215 22765
rect 10215 22761 10243 22765
rect 9905 22731 9939 22761
rect 9981 22731 10015 22761
rect 10057 22731 10091 22761
rect 10133 22731 10167 22761
rect 10209 22731 10243 22761
rect 10285 22731 10319 22765
rect 10361 22761 10391 22765
rect 10391 22761 10395 22765
rect 10437 22761 10461 22765
rect 10461 22761 10471 22765
rect 10513 22761 10530 22765
rect 10530 22761 10547 22765
rect 10589 22761 10599 22765
rect 10599 22761 10623 22765
rect 10665 22761 10668 22765
rect 10668 22761 10699 22765
rect 10759 22794 10771 22795
rect 10771 22794 10793 22795
rect 10832 22794 10840 22795
rect 10840 22794 10866 22795
rect 10905 22794 10909 22795
rect 10909 22794 10939 22795
rect 10978 22794 11012 22828
rect 11051 22795 11085 22828
rect 11124 22795 11158 22828
rect 11197 22795 11231 22828
rect 11270 22795 11304 22828
rect 11343 22795 11377 22828
rect 11416 22795 11450 22828
rect 11489 22795 11523 22828
rect 11562 22795 11596 22828
rect 11635 22795 11669 22828
rect 11707 22795 11741 22828
rect 11779 22795 11813 22828
rect 11851 22795 11885 22828
rect 11923 22795 11957 22828
rect 11995 22795 12029 22828
rect 12067 22795 12101 22828
rect 12139 22795 12173 22828
rect 12211 22795 12245 22828
rect 11051 22794 11082 22795
rect 11082 22794 11085 22795
rect 11124 22794 11151 22795
rect 11151 22794 11158 22795
rect 11197 22794 11220 22795
rect 11220 22794 11231 22795
rect 11270 22794 11289 22795
rect 11289 22794 11304 22795
rect 11343 22794 11358 22795
rect 11358 22794 11377 22795
rect 11416 22794 11427 22795
rect 11427 22794 11450 22795
rect 11489 22794 11496 22795
rect 11496 22794 11523 22795
rect 11562 22794 11565 22795
rect 11565 22794 11596 22795
rect 11635 22794 11668 22795
rect 11668 22794 11669 22795
rect 11707 22794 11737 22795
rect 11737 22794 11741 22795
rect 11779 22794 11806 22795
rect 11806 22794 11813 22795
rect 11851 22794 11875 22795
rect 11875 22794 11885 22795
rect 11923 22794 11944 22795
rect 11944 22794 11957 22795
rect 11995 22794 12013 22795
rect 12013 22794 12029 22795
rect 12067 22794 12082 22795
rect 12082 22794 12101 22795
rect 12139 22794 12151 22795
rect 12151 22794 12173 22795
rect 12211 22794 12220 22795
rect 12220 22794 12245 22795
rect 10361 22731 10395 22761
rect 10437 22731 10471 22761
rect 10513 22731 10547 22761
rect 10589 22731 10623 22761
rect 10665 22731 10699 22761
rect 10759 22725 10793 22742
rect 10832 22725 10866 22742
rect 10905 22725 10939 22742
rect 10759 22708 10771 22725
rect 10771 22708 10793 22725
rect 10832 22708 10840 22725
rect 10840 22708 10866 22725
rect 10905 22708 10909 22725
rect 10909 22708 10939 22725
rect 10978 22708 11012 22742
rect 11051 22725 11085 22742
rect 11124 22725 11158 22742
rect 11197 22725 11231 22742
rect 11270 22725 11304 22742
rect 11343 22725 11377 22742
rect 11416 22725 11450 22742
rect 11489 22725 11523 22742
rect 11562 22725 11596 22742
rect 11635 22725 11669 22742
rect 11707 22725 11741 22742
rect 11779 22725 11813 22742
rect 11851 22725 11885 22742
rect 11923 22725 11957 22742
rect 11995 22725 12029 22742
rect 12067 22725 12101 22742
rect 12139 22725 12173 22742
rect 12211 22725 12245 22742
rect 11051 22708 11082 22725
rect 11082 22708 11085 22725
rect 11124 22708 11151 22725
rect 11151 22708 11158 22725
rect 11197 22708 11220 22725
rect 11220 22708 11231 22725
rect 11270 22708 11289 22725
rect 11289 22708 11304 22725
rect 11343 22708 11358 22725
rect 11358 22708 11377 22725
rect 11416 22708 11427 22725
rect 11427 22708 11450 22725
rect 11489 22708 11496 22725
rect 11496 22708 11523 22725
rect 11562 22708 11565 22725
rect 11565 22708 11596 22725
rect 11635 22708 11668 22725
rect 11668 22708 11669 22725
rect 11707 22708 11737 22725
rect 11737 22708 11741 22725
rect 11779 22708 11806 22725
rect 11806 22708 11813 22725
rect 11851 22708 11875 22725
rect 11875 22708 11885 22725
rect 11923 22708 11944 22725
rect 11944 22708 11957 22725
rect 11995 22708 12013 22725
rect 12013 22708 12029 22725
rect 12067 22708 12082 22725
rect 12082 22708 12101 22725
rect 12139 22708 12151 22725
rect 12151 22708 12173 22725
rect 12211 22708 12220 22725
rect 12220 22708 12245 22725
rect 9905 22657 9939 22691
rect 9981 22657 10015 22691
rect 10057 22657 10091 22691
rect 10133 22657 10167 22691
rect 10209 22657 10243 22691
rect 10285 22657 10319 22691
rect 10361 22657 10395 22691
rect 10437 22657 10471 22691
rect 10513 22657 10547 22691
rect 10589 22657 10623 22691
rect 10665 22657 10699 22691
rect 10759 22655 10793 22656
rect 10832 22655 10866 22656
rect 10905 22655 10939 22656
rect 10759 22622 10771 22655
rect 10771 22622 10793 22655
rect 10832 22622 10840 22655
rect 10840 22622 10866 22655
rect 10905 22622 10909 22655
rect 10909 22622 10939 22655
rect 10978 22622 11012 22656
rect 11051 22655 11085 22656
rect 11124 22655 11158 22656
rect 11197 22655 11231 22656
rect 11270 22655 11304 22656
rect 11343 22655 11377 22656
rect 11416 22655 11450 22656
rect 11489 22655 11523 22656
rect 11562 22655 11596 22656
rect 11635 22655 11669 22656
rect 11707 22655 11741 22656
rect 11779 22655 11813 22656
rect 11851 22655 11885 22656
rect 11923 22655 11957 22656
rect 11995 22655 12029 22656
rect 12067 22655 12101 22656
rect 12139 22655 12173 22656
rect 12211 22655 12245 22656
rect 11051 22622 11082 22655
rect 11082 22622 11085 22655
rect 11124 22622 11151 22655
rect 11151 22622 11158 22655
rect 11197 22622 11220 22655
rect 11220 22622 11231 22655
rect 11270 22622 11289 22655
rect 11289 22622 11304 22655
rect 11343 22622 11358 22655
rect 11358 22622 11377 22655
rect 11416 22622 11427 22655
rect 11427 22622 11450 22655
rect 11489 22622 11496 22655
rect 11496 22622 11523 22655
rect 11562 22622 11565 22655
rect 11565 22622 11596 22655
rect 11635 22622 11668 22655
rect 11668 22622 11669 22655
rect 11707 22622 11737 22655
rect 11737 22622 11741 22655
rect 11779 22622 11806 22655
rect 11806 22622 11813 22655
rect 11851 22622 11875 22655
rect 11875 22622 11885 22655
rect 11923 22622 11944 22655
rect 11944 22622 11957 22655
rect 11995 22622 12013 22655
rect 12013 22622 12029 22655
rect 12067 22622 12082 22655
rect 12082 22622 12101 22655
rect 12139 22622 12151 22655
rect 12151 22622 12173 22655
rect 12211 22622 12220 22655
rect 12220 22622 12245 22655
rect 9905 22585 9939 22617
rect 9981 22585 10015 22617
rect 10057 22585 10091 22617
rect 10133 22585 10167 22617
rect 10209 22585 10243 22617
rect 9905 22583 9935 22585
rect 9935 22583 9939 22585
rect 9981 22583 10005 22585
rect 10005 22583 10015 22585
rect 10057 22583 10075 22585
rect 10075 22583 10091 22585
rect 10133 22583 10145 22585
rect 10145 22583 10167 22585
rect 10209 22583 10215 22585
rect 10215 22583 10243 22585
rect 10285 22583 10319 22617
rect 10361 22585 10395 22617
rect 10437 22585 10471 22617
rect 10513 22585 10547 22617
rect 10589 22585 10623 22617
rect 10665 22585 10699 22617
rect 10361 22583 10391 22585
rect 10391 22583 10395 22585
rect 10437 22583 10461 22585
rect 10461 22583 10471 22585
rect 10513 22583 10530 22585
rect 10530 22583 10547 22585
rect 10589 22583 10599 22585
rect 10599 22583 10623 22585
rect 10665 22583 10668 22585
rect 10668 22583 10699 22585
rect 13756 22891 13790 22925
rect 13828 22903 13862 22925
rect 13900 22903 13934 22925
rect 13972 22903 14006 22925
rect 14044 22903 14078 22925
rect 13828 22891 13830 22903
rect 13830 22891 13862 22903
rect 13900 22891 13932 22903
rect 13932 22891 13934 22903
rect 13972 22891 14000 22903
rect 14000 22891 14006 22903
rect 14044 22891 14068 22903
rect 14068 22891 14078 22903
rect 14116 22891 14150 22925
rect 14252 22873 14286 22905
rect 14324 22873 14358 22905
rect 14252 22871 14267 22873
rect 14267 22871 14286 22873
rect 14324 22871 14335 22873
rect 14335 22871 14358 22873
rect 13756 22817 13790 22851
rect 13828 22833 13862 22851
rect 13900 22833 13934 22851
rect 13972 22833 14006 22851
rect 14044 22833 14078 22851
rect 13828 22817 13830 22833
rect 13830 22817 13862 22833
rect 13900 22817 13932 22833
rect 13932 22817 13934 22833
rect 13972 22817 14000 22833
rect 14000 22817 14006 22833
rect 14044 22817 14068 22833
rect 14068 22817 14078 22833
rect 14116 22817 14150 22851
rect 14252 22804 14286 22832
rect 14324 22804 14358 22832
rect 14252 22798 14267 22804
rect 14267 22798 14286 22804
rect 14324 22798 14335 22804
rect 14335 22798 14358 22804
rect 13756 22743 13790 22777
rect 13828 22763 13862 22777
rect 13900 22763 13934 22777
rect 13972 22763 14006 22777
rect 14044 22763 14078 22777
rect 13828 22743 13830 22763
rect 13830 22743 13862 22763
rect 13900 22743 13932 22763
rect 13932 22743 13934 22763
rect 13972 22743 14000 22763
rect 14000 22743 14006 22763
rect 14044 22743 14068 22763
rect 14068 22743 14078 22763
rect 14116 22743 14150 22777
rect 14252 22735 14286 22759
rect 14324 22735 14358 22759
rect 14252 22725 14267 22735
rect 14267 22725 14286 22735
rect 14324 22725 14335 22735
rect 14335 22725 14358 22735
rect 13756 22669 13790 22703
rect 13828 22693 13862 22703
rect 13900 22693 13934 22703
rect 13972 22693 14006 22703
rect 14044 22693 14078 22703
rect 13828 22669 13830 22693
rect 13830 22669 13862 22693
rect 13900 22669 13932 22693
rect 13932 22669 13934 22693
rect 13972 22669 14000 22693
rect 14000 22669 14006 22693
rect 14044 22669 14068 22693
rect 14068 22669 14078 22693
rect 14116 22669 14150 22703
rect 14252 22666 14286 22686
rect 14324 22666 14358 22686
rect 14252 22652 14267 22666
rect 14267 22652 14286 22666
rect 14324 22652 14335 22666
rect 14335 22652 14358 22666
rect 13756 22595 13790 22629
rect 13828 22623 13862 22629
rect 13900 22623 13934 22629
rect 13972 22623 14006 22629
rect 14044 22623 14078 22629
rect 13828 22595 13830 22623
rect 13830 22595 13862 22623
rect 13900 22595 13932 22623
rect 13932 22595 13934 22623
rect 13972 22595 14000 22623
rect 14000 22595 14006 22623
rect 14044 22595 14068 22623
rect 14068 22595 14078 22623
rect 14116 22595 14150 22629
rect 14252 22597 14286 22613
rect 14324 22597 14358 22613
rect 14252 22579 14267 22597
rect 14267 22579 14286 22597
rect 14324 22579 14335 22597
rect 14335 22579 14358 22597
rect 13756 22521 13790 22555
rect 13828 22553 13862 22555
rect 13900 22553 13934 22555
rect 13972 22553 14006 22555
rect 14044 22553 14078 22555
rect 13828 22521 13830 22553
rect 13830 22521 13862 22553
rect 13900 22521 13932 22553
rect 13932 22521 13934 22553
rect 13972 22521 14000 22553
rect 14000 22521 14006 22553
rect 14044 22521 14068 22553
rect 14068 22521 14078 22553
rect 14116 22521 14150 22555
rect 14252 22528 14286 22540
rect 14324 22528 14358 22540
rect 14252 22506 14267 22528
rect 14267 22506 14286 22528
rect 14324 22506 14335 22528
rect 14335 22506 14358 22528
rect 13756 22447 13790 22481
rect 13828 22449 13830 22481
rect 13830 22449 13862 22481
rect 13900 22449 13932 22481
rect 13932 22449 13934 22481
rect 13972 22449 14000 22481
rect 14000 22449 14006 22481
rect 14044 22449 14068 22481
rect 14068 22449 14078 22481
rect 13828 22447 13862 22449
rect 13900 22447 13934 22449
rect 13972 22447 14006 22449
rect 14044 22447 14078 22449
rect 14116 22447 14150 22481
rect 14252 22459 14286 22467
rect 14324 22459 14358 22467
rect 14252 22433 14267 22459
rect 14267 22433 14286 22459
rect 14324 22433 14335 22459
rect 14335 22433 14358 22459
rect 13756 22373 13790 22407
rect 13828 22379 13830 22407
rect 13830 22379 13862 22407
rect 13900 22379 13932 22407
rect 13932 22379 13934 22407
rect 13972 22379 14000 22407
rect 14000 22379 14006 22407
rect 14044 22379 14068 22407
rect 14068 22379 14078 22407
rect 13828 22373 13862 22379
rect 13900 22373 13934 22379
rect 13972 22373 14006 22379
rect 14044 22373 14078 22379
rect 14116 22373 14150 22407
rect 14252 22390 14286 22394
rect 14324 22390 14358 22394
rect 14252 22360 14267 22390
rect 14267 22360 14286 22390
rect 14324 22360 14335 22390
rect 14335 22360 14358 22390
rect 13756 22299 13790 22333
rect 13828 22309 13830 22333
rect 13830 22309 13862 22333
rect 13900 22309 13932 22333
rect 13932 22309 13934 22333
rect 13972 22309 14000 22333
rect 14000 22309 14006 22333
rect 14044 22309 14068 22333
rect 14068 22309 14078 22333
rect 13828 22299 13862 22309
rect 13900 22299 13934 22309
rect 13972 22299 14006 22309
rect 14044 22299 14078 22309
rect 14116 22299 14150 22333
rect 14252 22287 14267 22321
rect 14267 22287 14286 22321
rect 14324 22287 14335 22321
rect 14335 22287 14358 22321
rect 13756 22225 13790 22259
rect 13828 22239 13830 22259
rect 13830 22239 13862 22259
rect 13900 22239 13932 22259
rect 13932 22239 13934 22259
rect 13972 22239 14000 22259
rect 14000 22239 14006 22259
rect 14044 22239 14068 22259
rect 14068 22239 14078 22259
rect 13828 22225 13862 22239
rect 13900 22225 13934 22239
rect 13972 22225 14006 22239
rect 14044 22225 14078 22239
rect 14116 22225 14150 22259
rect 14252 22218 14267 22248
rect 14267 22218 14286 22248
rect 14324 22218 14335 22248
rect 14335 22218 14358 22248
rect 14252 22214 14286 22218
rect 14324 22214 14358 22218
rect 13756 22151 13790 22185
rect 13828 22169 13830 22185
rect 13830 22169 13862 22185
rect 13900 22169 13932 22185
rect 13932 22169 13934 22185
rect 13972 22169 14000 22185
rect 14000 22169 14006 22185
rect 14044 22169 14068 22185
rect 14068 22169 14078 22185
rect 13828 22151 13862 22169
rect 13900 22151 13934 22169
rect 13972 22151 14006 22169
rect 14044 22151 14078 22169
rect 14116 22151 14150 22185
rect 14252 22149 14267 22175
rect 14267 22149 14286 22175
rect 14324 22149 14335 22175
rect 14335 22149 14358 22175
rect 14252 22141 14286 22149
rect 14324 22141 14358 22149
rect 13756 22077 13790 22111
rect 13828 22099 13830 22111
rect 13830 22099 13862 22111
rect 13900 22099 13932 22111
rect 13932 22099 13934 22111
rect 13972 22099 14000 22111
rect 14000 22099 14006 22111
rect 14044 22099 14068 22111
rect 14068 22099 14078 22111
rect 13828 22077 13862 22099
rect 13900 22077 13934 22099
rect 13972 22077 14006 22099
rect 14044 22077 14078 22099
rect 14116 22077 14150 22111
rect 14252 22080 14267 22102
rect 14267 22080 14286 22102
rect 14324 22080 14335 22102
rect 14335 22080 14358 22102
rect 14252 22068 14286 22080
rect 14324 22068 14358 22080
rect 13756 22003 13790 22037
rect 13828 22029 13830 22037
rect 13830 22029 13862 22037
rect 13900 22029 13932 22037
rect 13932 22029 13934 22037
rect 13972 22029 14000 22037
rect 14000 22029 14006 22037
rect 14044 22029 14068 22037
rect 14068 22029 14078 22037
rect 13828 22003 13862 22029
rect 13900 22003 13934 22029
rect 13972 22003 14006 22029
rect 14044 22003 14078 22029
rect 14116 22003 14150 22037
rect 14252 22011 14267 22029
rect 14267 22011 14286 22029
rect 14324 22011 14335 22029
rect 14335 22011 14358 22029
rect 14252 21995 14286 22011
rect 14324 21995 14358 22011
rect 13756 21929 13790 21963
rect 13828 21959 13830 21963
rect 13830 21959 13862 21963
rect 13900 21959 13932 21963
rect 13932 21959 13934 21963
rect 13972 21959 14000 21963
rect 14000 21959 14006 21963
rect 14044 21959 14068 21963
rect 14068 21959 14078 21963
rect 13828 21929 13862 21959
rect 13900 21929 13934 21959
rect 13972 21929 14006 21959
rect 14044 21929 14078 21959
rect 14116 21929 14150 21963
rect 14252 21942 14267 21956
rect 14267 21942 14286 21956
rect 14324 21942 14335 21956
rect 14335 21942 14358 21956
rect 14252 21922 14286 21942
rect 14324 21922 14358 21942
rect 13756 21855 13790 21889
rect 13828 21855 13862 21889
rect 13900 21855 13934 21889
rect 13972 21855 14006 21889
rect 14044 21855 14078 21889
rect 14116 21855 14150 21889
rect 14252 21873 14267 21883
rect 14267 21873 14286 21883
rect 14324 21873 14335 21883
rect 14335 21873 14358 21883
rect 14252 21849 14286 21873
rect 14324 21849 14358 21873
rect 13756 21781 13790 21815
rect 13828 21783 13862 21815
rect 13900 21783 13934 21815
rect 13972 21783 14006 21815
rect 14044 21783 14078 21815
rect 13828 21781 13830 21783
rect 13830 21781 13862 21783
rect 13900 21781 13932 21783
rect 13932 21781 13934 21783
rect 13972 21781 14000 21783
rect 14000 21781 14006 21783
rect 14044 21781 14068 21783
rect 14068 21781 14078 21783
rect 14116 21781 14150 21815
rect 14252 21804 14267 21810
rect 14267 21804 14286 21810
rect 14324 21804 14335 21810
rect 14335 21804 14358 21810
rect 14252 21776 14286 21804
rect 14324 21776 14358 21804
rect 13756 21707 13790 21741
rect 13828 21713 13862 21741
rect 13900 21713 13934 21741
rect 13972 21713 14006 21741
rect 14044 21713 14078 21741
rect 13828 21707 13830 21713
rect 13830 21707 13862 21713
rect 13900 21707 13932 21713
rect 13932 21707 13934 21713
rect 13972 21707 14000 21713
rect 14000 21707 14006 21713
rect 14044 21707 14068 21713
rect 14068 21707 14078 21713
rect 14116 21707 14150 21741
rect 14252 21735 14267 21737
rect 14267 21735 14286 21737
rect 14324 21735 14335 21737
rect 14335 21735 14358 21737
rect 14252 21703 14286 21735
rect 14324 21703 14358 21735
rect 13756 21632 13790 21666
rect 13828 21643 13862 21666
rect 13900 21643 13934 21666
rect 13972 21643 14006 21666
rect 14044 21643 14078 21666
rect 13828 21632 13830 21643
rect 13830 21632 13862 21643
rect 13900 21632 13932 21643
rect 13932 21632 13934 21643
rect 13972 21632 14000 21643
rect 14000 21632 14006 21643
rect 14044 21632 14068 21643
rect 14068 21632 14078 21643
rect 14116 21632 14150 21666
rect 14252 21631 14286 21664
rect 14324 21631 14358 21664
rect 14252 21630 14267 21631
rect 14267 21630 14286 21631
rect 14324 21630 14335 21631
rect 14335 21630 14358 21631
rect 13756 21557 13790 21591
rect 13828 21573 13862 21591
rect 13900 21573 13934 21591
rect 13972 21573 14006 21591
rect 14044 21573 14078 21591
rect 13828 21557 13830 21573
rect 13830 21557 13862 21573
rect 13900 21557 13932 21573
rect 13932 21557 13934 21573
rect 13972 21557 14000 21573
rect 14000 21557 14006 21573
rect 14044 21557 14068 21573
rect 14068 21557 14078 21573
rect 14116 21557 14150 21591
rect 14252 21562 14286 21591
rect 14324 21562 14358 21591
rect 14252 21557 14267 21562
rect 14267 21557 14286 21562
rect 14324 21557 14335 21562
rect 14335 21557 14358 21562
rect 13756 21482 13790 21516
rect 13828 21503 13862 21516
rect 13900 21503 13934 21516
rect 13972 21503 14006 21516
rect 14044 21503 14078 21516
rect 13828 21482 13830 21503
rect 13830 21482 13862 21503
rect 13900 21482 13932 21503
rect 13932 21482 13934 21503
rect 13972 21482 14000 21503
rect 14000 21482 14006 21503
rect 14044 21482 14068 21503
rect 14068 21482 14078 21503
rect 14116 21482 14150 21516
rect 14252 21493 14286 21518
rect 14324 21493 14358 21518
rect 14252 21484 14267 21493
rect 14267 21484 14286 21493
rect 14324 21484 14335 21493
rect 14335 21484 14358 21493
rect 13756 21407 13790 21441
rect 13828 21433 13862 21441
rect 13900 21433 13934 21441
rect 13972 21433 14006 21441
rect 14044 21433 14078 21441
rect 13828 21407 13830 21433
rect 13830 21407 13862 21433
rect 13900 21407 13932 21433
rect 13932 21407 13934 21433
rect 13972 21407 14000 21433
rect 14000 21407 14006 21433
rect 14044 21407 14068 21433
rect 14068 21407 14078 21433
rect 14116 21407 14150 21441
rect 14252 21424 14286 21445
rect 14324 21424 14358 21445
rect 14252 21411 14267 21424
rect 14267 21411 14286 21424
rect 14324 21411 14335 21424
rect 14335 21411 14358 21424
rect 13756 21332 13790 21366
rect 13828 21363 13862 21366
rect 13900 21363 13934 21366
rect 13972 21363 14006 21366
rect 14044 21363 14078 21366
rect 13828 21332 13830 21363
rect 13830 21332 13862 21363
rect 13900 21332 13932 21363
rect 13932 21332 13934 21363
rect 13972 21332 14000 21363
rect 14000 21332 14006 21363
rect 14044 21332 14068 21363
rect 14068 21332 14078 21363
rect 14116 21332 14150 21366
rect 14252 21355 14286 21371
rect 14324 21355 14358 21371
rect 14252 21337 14267 21355
rect 14267 21337 14286 21355
rect 14324 21337 14335 21355
rect 14335 21337 14358 21355
rect 13756 21257 13790 21291
rect 13828 21259 13830 21291
rect 13830 21259 13862 21291
rect 13900 21259 13932 21291
rect 13932 21259 13934 21291
rect 13972 21259 14000 21291
rect 14000 21259 14006 21291
rect 14044 21259 14068 21291
rect 14068 21259 14078 21291
rect 13828 21257 13862 21259
rect 13900 21257 13934 21259
rect 13972 21257 14006 21259
rect 14044 21257 14078 21259
rect 14116 21257 14150 21291
rect 14252 21286 14286 21297
rect 14324 21286 14358 21297
rect 14252 21263 14267 21286
rect 14267 21263 14286 21286
rect 14324 21263 14335 21286
rect 14335 21263 14358 21286
rect 13756 21182 13790 21216
rect 13828 21189 13830 21216
rect 13830 21189 13862 21216
rect 14252 21217 14286 21223
rect 14324 21217 14358 21223
rect 13900 21189 13932 21216
rect 13932 21189 13934 21216
rect 13972 21189 14000 21216
rect 14000 21189 14006 21216
rect 14044 21189 14068 21216
rect 14068 21189 14078 21216
rect 13828 21182 13862 21189
rect 13900 21182 13934 21189
rect 13972 21182 14006 21189
rect 14044 21182 14078 21189
rect 14116 21182 14150 21216
rect 14252 21189 14267 21217
rect 14267 21189 14286 21217
rect 14324 21189 14335 21217
rect 14335 21189 14358 21217
rect 13756 21107 13790 21141
rect 13828 21119 13830 21141
rect 13830 21119 13862 21141
rect 14252 21148 14286 21149
rect 14324 21148 14358 21149
rect 13900 21119 13932 21141
rect 13932 21119 13934 21141
rect 13972 21119 14000 21141
rect 14000 21119 14006 21141
rect 14044 21119 14068 21141
rect 14068 21119 14078 21141
rect 13828 21107 13862 21119
rect 13900 21107 13934 21119
rect 13972 21107 14006 21119
rect 14044 21107 14078 21119
rect 14116 21107 14150 21141
rect 14252 21115 14267 21148
rect 14267 21115 14286 21148
rect 14324 21115 14335 21148
rect 14335 21115 14358 21148
rect 13756 21032 13790 21066
rect 13828 21049 13830 21066
rect 13830 21049 13862 21066
rect 13900 21049 13932 21066
rect 13932 21049 13934 21066
rect 13972 21049 14000 21066
rect 14000 21049 14006 21066
rect 14044 21049 14068 21066
rect 14068 21049 14078 21066
rect 13828 21032 13862 21049
rect 13900 21032 13934 21049
rect 13972 21032 14006 21049
rect 14044 21032 14078 21049
rect 14116 21032 14150 21066
rect 14252 21045 14267 21075
rect 14267 21045 14286 21075
rect 14324 21045 14335 21075
rect 14335 21045 14358 21075
rect 14252 21041 14286 21045
rect 14324 21041 14358 21045
rect 10911 17325 10945 17359
rect 10911 17253 10945 17287
rect 1807 10981 1841 11015
rect 1807 10909 1841 10943
rect 1807 10837 1841 10871
rect 1807 10765 1841 10799
rect 1923 10981 1957 11015
rect 1923 10909 1957 10943
rect 1923 10837 1957 10871
rect 1923 10765 1957 10799
rect 846 5349 880 5383
rect 926 5349 960 5383
rect 1005 5349 1039 5383
rect 1084 5349 1118 5383
rect 1163 5349 1197 5383
rect 1242 5349 1276 5383
rect 1321 5349 1355 5383
rect 1400 5349 1434 5383
rect 1479 5349 1513 5383
rect 1558 5349 1592 5383
rect 951 3271 985 3305
rect 951 3199 985 3233
rect 1807 3298 1841 3332
rect 1807 3226 1841 3260
rect 1807 3154 1841 3188
rect 1807 3082 1841 3116
rect 1923 3298 1957 3332
rect 1923 3226 1957 3260
rect 1923 3154 1957 3188
rect 1923 3082 1957 3116
rect 11365 1468 11399 1486
rect 11365 1452 11399 1468
rect 11437 1458 11471 1492
rect 11509 1458 11543 1492
rect 11581 1458 11615 1492
rect 11653 1458 11687 1492
rect 11725 1458 11759 1492
rect 11797 1458 11831 1492
rect 11869 1458 11903 1492
rect 11941 1458 11975 1492
rect 12013 1458 12047 1492
rect 12085 1458 12119 1492
rect 12157 1458 12191 1492
rect 12229 1458 12263 1492
rect 12301 1458 12335 1492
rect 12373 1458 12407 1492
rect 12445 1458 12479 1492
rect 12517 1458 12551 1492
rect 12589 1458 12623 1492
rect 12661 1458 12695 1492
rect 12733 1458 12767 1492
rect 12805 1458 12839 1492
rect 12877 1458 12911 1492
rect 12949 1458 12983 1492
rect 13021 1458 13055 1492
rect 13093 1458 13127 1492
rect 13165 1458 13199 1492
rect 13237 1458 13271 1492
rect 13309 1458 13343 1492
rect 13381 1468 13415 1486
rect 11365 1393 11399 1406
rect 11365 1372 11399 1393
rect 13381 1452 13415 1468
rect 13381 1393 13415 1406
rect 11365 1318 11399 1325
rect 11365 1291 11399 1318
rect 11365 1243 11399 1244
rect 11365 1210 11399 1243
rect 13381 1372 13415 1393
rect 13381 1318 13415 1325
rect 13381 1291 13415 1318
rect 13381 1243 13415 1244
rect 11365 1134 11399 1163
rect 11365 1129 11399 1134
rect 11365 1058 11399 1082
rect 11365 1048 11399 1058
rect 11481 1192 11515 1226
rect 11481 1120 11515 1154
rect 11481 1048 11515 1082
rect 11737 1192 11771 1226
rect 11737 1120 11771 1154
rect 11737 1048 11771 1082
rect 11861 1192 11895 1226
rect 11861 1120 11895 1154
rect 11861 1048 11895 1082
rect 12117 1192 12151 1226
rect 12117 1120 12151 1154
rect 12243 1192 12277 1226
rect 12243 1120 12277 1154
rect 12373 1192 12407 1226
rect 12373 1120 12407 1154
rect 12503 1192 12537 1226
rect 12503 1120 12537 1154
rect 12629 1192 12663 1226
rect 12629 1120 12663 1154
rect 12117 1048 12151 1082
rect 12373 1048 12407 1082
rect 12629 1048 12663 1082
rect 12885 1192 12919 1226
rect 12885 1120 12919 1154
rect 12885 1048 12919 1082
rect 13009 1192 13043 1226
rect 13009 1120 13043 1154
rect 13009 1048 13043 1082
rect 13265 1192 13299 1226
rect 13265 1120 13299 1154
rect 13265 1048 13299 1082
rect 13381 1210 13415 1243
rect 13381 1134 13415 1163
rect 13381 1129 13415 1134
rect 13381 1058 13415 1082
rect 13381 1048 13415 1058
rect 11365 798 11399 814
rect 11365 780 11399 798
rect 11365 714 11399 719
rect 11365 685 11399 714
rect 11481 780 11515 814
rect 11481 708 11515 742
rect 11481 636 11515 670
rect 11737 780 11771 814
rect 11737 708 11771 742
rect 11737 636 11771 670
rect 11993 780 12027 814
rect 11993 708 12027 742
rect 12753 780 12787 814
rect 12753 708 12787 742
rect 11993 636 12027 670
rect 12093 624 12127 658
rect 12165 624 12199 658
rect 12237 624 12271 658
rect 12369 644 12403 678
rect 11365 596 11399 624
rect 11365 590 11399 596
rect 12509 624 12543 658
rect 12581 624 12615 658
rect 12653 624 12687 658
rect 12753 636 12787 670
rect 13009 780 13043 814
rect 13009 708 13043 742
rect 13009 636 13043 670
rect 13265 780 13299 814
rect 13265 708 13299 742
rect 13265 636 13299 670
rect 13381 798 13415 814
rect 13381 780 13415 798
rect 13381 714 13415 719
rect 13381 685 13415 714
rect 12369 560 12403 594
rect 13381 596 13415 624
rect 13381 590 13415 596
rect 11365 512 11399 528
rect 11365 494 11399 512
rect 11437 488 11471 522
rect 11509 488 11543 522
rect 11581 488 11615 522
rect 11653 488 11687 522
rect 11725 488 11759 522
rect 11797 488 11831 522
rect 11869 488 11903 522
rect 11941 488 11975 522
rect 12013 488 12047 522
rect 12085 488 12119 522
rect 12157 488 12191 522
rect 12229 488 12263 522
rect 12301 488 12335 522
rect 12373 488 12407 522
rect 12445 488 12479 522
rect 12517 488 12551 522
rect 12589 488 12623 522
rect 12661 488 12695 522
rect 12733 488 12767 522
rect 12805 488 12839 522
rect 12877 488 12911 522
rect 12949 488 12983 522
rect 13021 488 13055 522
rect 13093 488 13127 522
rect 13165 488 13199 522
rect 13237 488 13271 522
rect 13309 488 13343 522
rect 13381 512 13415 528
rect 13381 494 13415 512
<< metal1 >>
rect 9877 36379 14429 36388
rect 9877 36351 10927 36379
rect 9877 36317 9915 36351
rect 9949 36317 9987 36351
rect 10021 36317 10059 36351
rect 10093 36317 10131 36351
rect 10165 36317 10203 36351
rect 10237 36317 10275 36351
rect 10309 36317 10347 36351
rect 10381 36317 10419 36351
rect 10453 36317 10491 36351
rect 10525 36317 10563 36351
rect 10597 36317 10635 36351
rect 10669 36317 10707 36351
rect 10741 36317 10779 36351
rect 10813 36317 10851 36351
rect 10885 36345 10927 36351
rect 10961 36345 11000 36379
rect 11034 36345 11073 36379
rect 11107 36345 11146 36379
rect 11180 36345 11219 36379
rect 11253 36345 11292 36379
rect 11326 36345 11365 36379
rect 11399 36345 11438 36379
rect 11472 36345 11511 36379
rect 11545 36345 11584 36379
rect 11618 36345 11657 36379
rect 11691 36345 11730 36379
rect 11764 36345 11803 36379
rect 11837 36345 11876 36379
rect 11910 36345 11949 36379
rect 11983 36345 12022 36379
rect 12056 36345 12095 36379
rect 12129 36345 12168 36379
rect 12202 36345 12241 36379
rect 12275 36345 12314 36379
rect 12348 36345 12387 36379
rect 12421 36345 12460 36379
rect 12494 36345 12533 36379
rect 12567 36345 12606 36379
rect 12640 36345 12679 36379
rect 12713 36345 12752 36379
rect 12786 36345 12825 36379
rect 12859 36345 12898 36379
rect 12932 36345 12971 36379
rect 13005 36345 13044 36379
rect 13078 36345 13117 36379
rect 13151 36345 13190 36379
rect 13224 36345 13263 36379
rect 13297 36345 13336 36379
rect 13370 36345 13409 36379
rect 13443 36345 13482 36379
rect 13516 36345 13555 36379
rect 13589 36345 13628 36379
rect 13662 36345 13701 36379
rect 13735 36345 13774 36379
rect 13808 36345 13846 36379
rect 13880 36345 13918 36379
rect 13952 36345 13990 36379
rect 14024 36345 14062 36379
rect 14096 36345 14134 36379
rect 14168 36345 14206 36379
rect 14240 36345 14278 36379
rect 14312 36345 14350 36379
rect 14384 36345 14429 36379
rect 10885 36317 14429 36345
rect 9877 36303 14429 36317
rect 9877 36273 10927 36303
rect 9877 36239 9915 36273
rect 9949 36239 9987 36273
rect 10021 36239 10059 36273
rect 10093 36239 10131 36273
rect 10165 36239 10203 36273
rect 10237 36239 10275 36273
rect 10309 36239 10347 36273
rect 10381 36239 10419 36273
rect 10453 36239 10491 36273
rect 10525 36239 10563 36273
rect 10597 36239 10635 36273
rect 10669 36239 10707 36273
rect 10741 36239 10779 36273
rect 10813 36239 10851 36273
rect 10885 36269 10927 36273
rect 10961 36269 11000 36303
rect 11034 36269 11073 36303
rect 11107 36269 11146 36303
rect 11180 36269 11219 36303
rect 11253 36269 11292 36303
rect 11326 36269 11365 36303
rect 11399 36269 11438 36303
rect 11472 36269 11511 36303
rect 11545 36269 11584 36303
rect 11618 36269 11657 36303
rect 11691 36269 11730 36303
rect 11764 36269 11803 36303
rect 11837 36269 11876 36303
rect 11910 36269 11949 36303
rect 11983 36269 12022 36303
rect 12056 36269 12095 36303
rect 12129 36269 12168 36303
rect 12202 36269 12241 36303
rect 12275 36269 12314 36303
rect 12348 36269 12387 36303
rect 12421 36269 12460 36303
rect 12494 36269 12533 36303
rect 12567 36269 12606 36303
rect 12640 36269 12679 36303
rect 12713 36269 12752 36303
rect 12786 36269 12825 36303
rect 12859 36269 12898 36303
rect 12932 36269 12971 36303
rect 13005 36269 13044 36303
rect 13078 36269 13117 36303
rect 13151 36269 13190 36303
rect 13224 36269 13263 36303
rect 13297 36269 13336 36303
rect 13370 36269 13409 36303
rect 13443 36269 13482 36303
rect 13516 36269 13555 36303
rect 13589 36269 13628 36303
rect 13662 36269 13701 36303
rect 13735 36269 13774 36303
rect 13808 36269 13846 36303
rect 13880 36269 13918 36303
rect 13952 36269 13990 36303
rect 14024 36269 14062 36303
rect 14096 36269 14134 36303
rect 14168 36269 14206 36303
rect 14240 36269 14278 36303
rect 14312 36269 14350 36303
rect 14384 36269 14429 36303
rect 10885 36239 14429 36269
rect 9877 36227 14429 36239
rect 9877 36195 10927 36227
rect 9877 36161 9915 36195
rect 9949 36161 9987 36195
rect 10021 36161 10059 36195
rect 10093 36161 10131 36195
rect 10165 36161 10203 36195
rect 10237 36161 10275 36195
rect 10309 36161 10347 36195
rect 10381 36161 10419 36195
rect 10453 36161 10491 36195
rect 10525 36161 10563 36195
rect 10597 36161 10635 36195
rect 10669 36161 10707 36195
rect 10741 36161 10779 36195
rect 10813 36161 10851 36195
rect 10885 36193 10927 36195
rect 10961 36193 11000 36227
rect 11034 36193 11073 36227
rect 11107 36193 11146 36227
rect 11180 36193 11219 36227
rect 11253 36193 11292 36227
rect 11326 36193 11365 36227
rect 11399 36193 11438 36227
rect 11472 36193 11511 36227
rect 11545 36193 11584 36227
rect 11618 36193 11657 36227
rect 11691 36193 11730 36227
rect 11764 36193 11803 36227
rect 11837 36193 11876 36227
rect 11910 36193 11949 36227
rect 11983 36193 12022 36227
rect 12056 36193 12095 36227
rect 12129 36193 12168 36227
rect 12202 36193 12241 36227
rect 12275 36193 12314 36227
rect 12348 36193 12387 36227
rect 12421 36193 12460 36227
rect 12494 36193 12533 36227
rect 12567 36193 12606 36227
rect 12640 36193 12679 36227
rect 12713 36193 12752 36227
rect 12786 36193 12825 36227
rect 12859 36193 12898 36227
rect 12932 36193 12971 36227
rect 13005 36193 13044 36227
rect 13078 36193 13117 36227
rect 13151 36193 13190 36227
rect 13224 36193 13263 36227
rect 13297 36193 13336 36227
rect 13370 36193 13409 36227
rect 13443 36193 13482 36227
rect 13516 36193 13555 36227
rect 13589 36193 13628 36227
rect 13662 36193 13701 36227
rect 13735 36193 13774 36227
rect 13808 36193 13846 36227
rect 13880 36193 13918 36227
rect 13952 36193 13990 36227
rect 14024 36193 14062 36227
rect 14096 36193 14134 36227
rect 14168 36193 14206 36227
rect 14240 36193 14278 36227
rect 14312 36193 14350 36227
rect 14384 36193 14429 36227
rect 10885 36161 14429 36193
rect 9877 36151 14429 36161
rect 9877 36117 10927 36151
rect 10961 36117 11000 36151
rect 11034 36117 11073 36151
rect 11107 36117 11146 36151
rect 11180 36117 11219 36151
rect 11253 36117 11292 36151
rect 11326 36117 11365 36151
rect 11399 36117 11438 36151
rect 11472 36117 11511 36151
rect 11545 36117 11584 36151
rect 11618 36117 11657 36151
rect 11691 36117 11730 36151
rect 11764 36117 11803 36151
rect 11837 36117 11876 36151
rect 11910 36117 11949 36151
rect 11983 36117 12022 36151
rect 12056 36117 12095 36151
rect 12129 36117 12168 36151
rect 12202 36117 12241 36151
rect 12275 36117 12314 36151
rect 12348 36117 12387 36151
rect 12421 36117 12460 36151
rect 12494 36117 12533 36151
rect 12567 36117 12606 36151
rect 12640 36117 12679 36151
rect 12713 36117 12752 36151
rect 12786 36117 12825 36151
rect 12859 36117 12898 36151
rect 12932 36117 12971 36151
rect 13005 36117 13044 36151
rect 13078 36117 13117 36151
rect 13151 36117 13190 36151
rect 13224 36117 13263 36151
rect 13297 36117 13336 36151
rect 13370 36117 13409 36151
rect 13443 36117 13482 36151
rect 13516 36117 13555 36151
rect 13589 36117 13628 36151
rect 13662 36117 13701 36151
rect 13735 36117 13774 36151
rect 13808 36117 13846 36151
rect 13880 36117 13918 36151
rect 13952 36117 13990 36151
rect 14024 36117 14062 36151
rect 14096 36117 14134 36151
rect 14168 36117 14206 36151
rect 14240 36117 14278 36151
rect 14312 36117 14350 36151
rect 14384 36117 14429 36151
rect 9877 36116 14429 36117
rect 9877 36082 9915 36116
rect 9949 36082 9987 36116
rect 10021 36082 10059 36116
rect 10093 36082 10131 36116
rect 10165 36082 10203 36116
rect 10237 36082 10275 36116
rect 10309 36082 10347 36116
rect 10381 36082 10419 36116
rect 10453 36082 10491 36116
rect 10525 36082 10563 36116
rect 10597 36082 10635 36116
rect 10669 36082 10707 36116
rect 10741 36082 10779 36116
rect 10813 36082 10851 36116
rect 10885 36082 14429 36116
rect 9877 36075 14429 36082
rect 9877 36041 10927 36075
rect 10961 36041 11000 36075
rect 11034 36041 11073 36075
rect 11107 36041 11146 36075
rect 11180 36041 11219 36075
rect 11253 36041 11292 36075
rect 11326 36041 11365 36075
rect 11399 36041 11438 36075
rect 11472 36041 11511 36075
rect 11545 36041 11584 36075
rect 11618 36041 11657 36075
rect 11691 36041 11730 36075
rect 11764 36041 11803 36075
rect 11837 36041 11876 36075
rect 11910 36041 11949 36075
rect 11983 36041 12022 36075
rect 12056 36041 12095 36075
rect 12129 36041 12168 36075
rect 12202 36041 12241 36075
rect 12275 36041 12314 36075
rect 12348 36041 12387 36075
rect 12421 36041 12460 36075
rect 12494 36041 12533 36075
rect 12567 36041 12606 36075
rect 12640 36041 12679 36075
rect 12713 36041 12752 36075
rect 12786 36041 12825 36075
rect 12859 36041 12898 36075
rect 12932 36041 12971 36075
rect 13005 36041 13044 36075
rect 13078 36041 13117 36075
rect 13151 36041 13190 36075
rect 13224 36041 13263 36075
rect 13297 36041 13336 36075
rect 13370 36041 13409 36075
rect 13443 36041 13482 36075
rect 13516 36041 13555 36075
rect 13589 36041 13628 36075
rect 13662 36041 13701 36075
rect 13735 36041 13774 36075
rect 13808 36041 13846 36075
rect 13880 36041 13918 36075
rect 13952 36041 13990 36075
rect 14024 36041 14062 36075
rect 14096 36041 14134 36075
rect 14168 36041 14206 36075
rect 14240 36041 14278 36075
rect 14312 36041 14350 36075
rect 14384 36041 14429 36075
rect 9877 36037 14429 36041
rect 9877 36003 9915 36037
rect 9949 36003 9987 36037
rect 10021 36003 10059 36037
rect 10093 36003 10131 36037
rect 10165 36003 10203 36037
rect 10237 36003 10275 36037
rect 10309 36003 10347 36037
rect 10381 36003 10419 36037
rect 10453 36003 10491 36037
rect 10525 36003 10563 36037
rect 10597 36003 10635 36037
rect 10669 36003 10707 36037
rect 10741 36003 10779 36037
rect 10813 36003 10851 36037
rect 10885 36003 14429 36037
rect 9877 35999 14429 36003
rect 9877 35965 10927 35999
rect 10961 35965 11000 35999
rect 11034 35965 11073 35999
rect 11107 35965 11146 35999
rect 11180 35965 11219 35999
rect 11253 35965 11292 35999
rect 11326 35965 11365 35999
rect 11399 35965 11438 35999
rect 11472 35965 11511 35999
rect 11545 35965 11584 35999
rect 11618 35965 11657 35999
rect 11691 35965 11730 35999
rect 11764 35965 11803 35999
rect 11837 35965 11876 35999
rect 11910 35965 11949 35999
rect 11983 35965 12022 35999
rect 12056 35965 12095 35999
rect 12129 35965 12168 35999
rect 12202 35965 12241 35999
rect 12275 35965 12314 35999
rect 12348 35965 12387 35999
rect 12421 35965 12460 35999
rect 12494 35965 12533 35999
rect 12567 35965 12606 35999
rect 12640 35965 12679 35999
rect 12713 35965 12752 35999
rect 12786 35965 12825 35999
rect 12859 35965 12898 35999
rect 12932 35965 12971 35999
rect 13005 35965 13044 35999
rect 13078 35965 13117 35999
rect 13151 35965 13190 35999
rect 13224 35965 13263 35999
rect 13297 35965 13336 35999
rect 13370 35965 13409 35999
rect 13443 35965 13482 35999
rect 13516 35965 13555 35999
rect 13589 35965 13628 35999
rect 13662 35965 13701 35999
rect 13735 35965 13774 35999
rect 13808 35965 13846 35999
rect 13880 35965 13918 35999
rect 13952 35965 13990 35999
rect 14024 35965 14062 35999
rect 14096 35965 14134 35999
rect 14168 35965 14206 35999
rect 14240 35965 14278 35999
rect 14312 35965 14350 35999
rect 14384 35965 14429 35999
rect 9877 35958 14429 35965
rect 9877 35924 9915 35958
rect 9949 35924 9987 35958
rect 10021 35924 10059 35958
rect 10093 35924 10131 35958
rect 10165 35924 10203 35958
rect 10237 35924 10275 35958
rect 10309 35924 10347 35958
rect 10381 35924 10419 35958
rect 10453 35924 10491 35958
rect 10525 35924 10563 35958
rect 10597 35924 10635 35958
rect 10669 35924 10707 35958
rect 10741 35924 10779 35958
rect 10813 35924 10851 35958
rect 10885 35924 14429 35958
rect 9877 35923 14429 35924
rect 9877 35889 10927 35923
rect 10961 35889 11000 35923
rect 11034 35889 11073 35923
rect 11107 35889 11146 35923
rect 11180 35889 11219 35923
rect 11253 35889 11292 35923
rect 11326 35889 11365 35923
rect 11399 35889 11438 35923
rect 11472 35889 11511 35923
rect 11545 35889 11584 35923
rect 11618 35889 11657 35923
rect 11691 35889 11730 35923
rect 11764 35889 11803 35923
rect 11837 35889 11876 35923
rect 11910 35889 11949 35923
rect 11983 35889 12022 35923
rect 12056 35889 12095 35923
rect 12129 35889 12168 35923
rect 12202 35889 12241 35923
rect 12275 35889 12314 35923
rect 12348 35889 12387 35923
rect 12421 35889 12460 35923
rect 12494 35889 12533 35923
rect 12567 35889 12606 35923
rect 12640 35889 12679 35923
rect 12713 35889 12752 35923
rect 12786 35889 12825 35923
rect 12859 35889 12898 35923
rect 12932 35889 12971 35923
rect 13005 35889 13044 35923
rect 13078 35889 13117 35923
rect 13151 35889 13190 35923
rect 13224 35889 13263 35923
rect 13297 35889 13336 35923
rect 13370 35889 13409 35923
rect 13443 35889 13482 35923
rect 13516 35889 13555 35923
rect 13589 35889 13628 35923
rect 13662 35889 13701 35923
rect 13735 35889 13774 35923
rect 13808 35889 13846 35923
rect 13880 35889 13918 35923
rect 13952 35889 13990 35923
rect 14024 35889 14062 35923
rect 14096 35889 14134 35923
rect 14168 35889 14206 35923
rect 14240 35889 14278 35923
rect 14312 35889 14350 35923
rect 14384 35889 14429 35923
rect 9877 35879 14429 35889
rect 9877 35845 9915 35879
rect 9949 35845 9987 35879
rect 10021 35845 10059 35879
rect 10093 35845 10131 35879
rect 10165 35845 10203 35879
rect 10237 35845 10275 35879
rect 10309 35845 10347 35879
rect 10381 35845 10419 35879
rect 10453 35845 10491 35879
rect 10525 35845 10563 35879
rect 10597 35845 10635 35879
rect 10669 35845 10707 35879
rect 10741 35845 10779 35879
rect 10813 35845 10851 35879
rect 10885 35847 14429 35879
rect 10885 35845 10927 35847
rect 9877 35813 10927 35845
rect 10961 35813 11000 35847
rect 11034 35813 11073 35847
rect 11107 35813 11146 35847
rect 11180 35813 11219 35847
rect 11253 35813 11292 35847
rect 11326 35813 11365 35847
rect 11399 35813 11438 35847
rect 11472 35813 11511 35847
rect 11545 35813 11584 35847
rect 11618 35813 11657 35847
rect 11691 35813 11730 35847
rect 11764 35813 11803 35847
rect 11837 35813 11876 35847
rect 11910 35813 11949 35847
rect 11983 35813 12022 35847
rect 12056 35813 12095 35847
rect 12129 35813 12168 35847
rect 12202 35813 12241 35847
rect 12275 35813 12314 35847
rect 12348 35813 12387 35847
rect 12421 35813 12460 35847
rect 12494 35813 12533 35847
rect 12567 35813 12606 35847
rect 12640 35813 12679 35847
rect 12713 35813 12752 35847
rect 12786 35813 12825 35847
rect 12859 35813 12898 35847
rect 12932 35813 12971 35847
rect 13005 35813 13044 35847
rect 13078 35813 13117 35847
rect 13151 35813 13190 35847
rect 13224 35813 13263 35847
rect 13297 35813 13336 35847
rect 13370 35813 13409 35847
rect 13443 35813 13482 35847
rect 13516 35813 13555 35847
rect 13589 35813 13628 35847
rect 13662 35813 13701 35847
rect 13735 35813 13774 35847
rect 13808 35813 13846 35847
rect 13880 35813 13918 35847
rect 13952 35813 13990 35847
rect 14024 35813 14062 35847
rect 14096 35813 14134 35847
rect 14168 35813 14206 35847
rect 14240 35813 14278 35847
rect 14312 35813 14350 35847
rect 14384 35813 14429 35847
rect 9877 35800 14429 35813
rect 9877 35766 9915 35800
rect 9949 35766 9987 35800
rect 10021 35766 10059 35800
rect 10093 35766 10131 35800
rect 10165 35766 10203 35800
rect 10237 35766 10275 35800
rect 10309 35766 10347 35800
rect 10381 35766 10419 35800
rect 10453 35766 10491 35800
rect 10525 35766 10563 35800
rect 10597 35766 10635 35800
rect 10669 35766 10707 35800
rect 10741 35766 10779 35800
rect 10813 35766 10851 35800
rect 10885 35771 14429 35800
rect 10885 35766 10927 35771
rect 9877 35737 10927 35766
rect 10961 35737 11000 35771
rect 11034 35737 11073 35771
rect 11107 35737 11146 35771
rect 11180 35737 11219 35771
rect 11253 35737 11292 35771
rect 11326 35737 11365 35771
rect 11399 35737 11438 35771
rect 11472 35737 11511 35771
rect 11545 35737 11584 35771
rect 11618 35737 11657 35771
rect 11691 35737 11730 35771
rect 11764 35737 11803 35771
rect 11837 35737 11876 35771
rect 11910 35737 11949 35771
rect 11983 35737 12022 35771
rect 12056 35737 12095 35771
rect 12129 35737 12168 35771
rect 12202 35737 12241 35771
rect 12275 35737 12314 35771
rect 12348 35737 12387 35771
rect 12421 35737 12460 35771
rect 12494 35737 12533 35771
rect 12567 35737 12606 35771
rect 12640 35737 12679 35771
rect 12713 35737 12752 35771
rect 12786 35737 12825 35771
rect 12859 35737 12898 35771
rect 12932 35737 12971 35771
rect 13005 35737 13044 35771
rect 13078 35737 13117 35771
rect 13151 35737 13190 35771
rect 13224 35737 13263 35771
rect 13297 35737 13336 35771
rect 13370 35737 13409 35771
rect 13443 35737 13482 35771
rect 13516 35737 13555 35771
rect 13589 35737 13628 35771
rect 13662 35737 13701 35771
rect 13735 35737 13774 35771
rect 13808 35737 13846 35771
rect 13880 35737 13918 35771
rect 13952 35737 13990 35771
rect 14024 35737 14062 35771
rect 14096 35737 14134 35771
rect 14168 35737 14206 35771
rect 14240 35737 14278 35771
rect 14312 35737 14350 35771
rect 14384 35737 14429 35771
rect 9877 35697 14429 35737
rect 9877 35687 13216 35697
tri 12949 35663 12973 35687 ne
rect 12973 35663 13216 35687
rect 13250 35663 13289 35697
rect 13323 35663 13362 35697
rect 13396 35663 13435 35697
rect 13469 35663 13508 35697
rect 13542 35663 13581 35697
rect 13615 35663 13654 35697
rect 13688 35663 13727 35697
rect 13761 35663 13800 35697
rect 13834 35663 13873 35697
rect 13907 35663 13946 35697
rect 13980 35663 14019 35697
rect 14053 35663 14092 35697
rect 14126 35663 14165 35697
rect 14199 35663 14238 35697
rect 14272 35663 14311 35697
rect 14345 35663 14384 35697
rect 14418 35663 14429 35697
tri 12973 35625 13011 35663 ne
rect 13011 35625 14429 35663
tri 13011 35591 13045 35625 ne
rect 13045 35591 13216 35625
rect 13250 35591 13289 35625
rect 13323 35591 13362 35625
rect 13396 35591 13435 35625
rect 13469 35591 13508 35625
rect 13542 35591 13581 35625
rect 13615 35591 13654 35625
rect 13688 35591 13727 35625
rect 13761 35591 13800 35625
rect 13834 35591 13873 35625
rect 13907 35591 13946 35625
rect 13980 35591 14019 35625
rect 14053 35591 14092 35625
rect 14126 35591 14165 35625
rect 14199 35591 14238 35625
rect 14272 35591 14311 35625
rect 14345 35591 14384 35625
rect 14418 35591 14429 35625
tri 13045 35553 13083 35591 ne
rect 13083 35553 14429 35591
tri 13083 35519 13117 35553 ne
rect 13117 35519 13216 35553
rect 13250 35519 13289 35553
rect 13323 35519 13362 35553
rect 13396 35519 13435 35553
rect 13469 35519 13508 35553
rect 13542 35519 13581 35553
rect 13615 35519 13654 35553
rect 13688 35519 13727 35553
rect 13761 35519 13800 35553
rect 13834 35519 13873 35553
rect 13907 35519 13946 35553
rect 13980 35519 14019 35553
rect 14053 35519 14092 35553
rect 14126 35519 14165 35553
rect 14199 35519 14238 35553
rect 14272 35519 14311 35553
rect 14345 35519 14384 35553
rect 14418 35519 14429 35553
tri 13117 35481 13155 35519 ne
rect 13155 35481 14429 35519
tri 13155 35461 13175 35481 ne
rect 13175 35447 13216 35481
rect 13250 35447 13289 35481
rect 13323 35447 13362 35481
rect 13396 35447 13435 35481
rect 13469 35447 13508 35481
rect 13542 35447 13581 35481
rect 13615 35447 13654 35481
rect 13688 35447 13727 35481
rect 13761 35447 13800 35481
rect 13834 35447 13873 35481
rect 13907 35447 13946 35481
rect 13980 35447 14019 35481
rect 14053 35447 14092 35481
rect 14126 35447 14165 35481
rect 14199 35447 14238 35481
rect 14272 35447 14311 35481
rect 14345 35447 14384 35481
rect 14418 35447 14429 35481
rect 13175 35409 14429 35447
rect 13175 35375 13216 35409
rect 13250 35375 13289 35409
rect 13323 35375 13362 35409
rect 13396 35375 13435 35409
rect 13469 35375 13508 35409
rect 13542 35375 13581 35409
rect 13615 35375 13654 35409
rect 13688 35375 13727 35409
rect 13761 35375 13800 35409
rect 13834 35375 13873 35409
rect 13907 35375 13946 35409
rect 13980 35375 14019 35409
rect 14053 35375 14092 35409
rect 14126 35375 14165 35409
rect 14199 35375 14238 35409
rect 14272 35375 14311 35409
rect 14345 35375 14384 35409
rect 14418 35375 14429 35409
rect 13175 35337 14429 35375
rect 13175 35303 13216 35337
rect 13250 35303 13289 35337
rect 13323 35303 13362 35337
rect 13396 35303 13435 35337
rect 13469 35303 13508 35337
rect 13542 35303 13581 35337
rect 13615 35303 13654 35337
rect 13688 35303 13727 35337
rect 13761 35303 13800 35337
rect 13834 35303 13873 35337
rect 13907 35303 13946 35337
rect 13980 35303 14019 35337
rect 14053 35303 14092 35337
rect 14126 35303 14165 35337
rect 14199 35303 14238 35337
rect 14272 35303 14311 35337
rect 14345 35303 14384 35337
rect 14418 35303 14429 35337
rect 13175 35265 14429 35303
rect 13175 35231 13216 35265
rect 13250 35231 13289 35265
rect 13323 35231 13362 35265
rect 13396 35231 13435 35265
rect 13469 35231 13508 35265
rect 13542 35231 13581 35265
rect 13615 35231 13654 35265
rect 13688 35231 13727 35265
rect 13761 35231 13800 35265
rect 13834 35231 13873 35265
rect 13907 35231 13946 35265
rect 13980 35231 14019 35265
rect 14053 35231 14092 35265
rect 14126 35231 14165 35265
rect 14199 35231 14238 35265
rect 14272 35231 14311 35265
rect 14345 35231 14384 35265
rect 14418 35231 14429 35265
rect 13175 35193 14429 35231
rect 13175 35159 13216 35193
rect 13250 35159 13289 35193
rect 13323 35159 13362 35193
rect 13396 35159 13435 35193
rect 13469 35159 13508 35193
rect 13542 35159 13581 35193
rect 13615 35159 13654 35193
rect 13688 35159 13727 35193
rect 13761 35159 13800 35193
rect 13834 35159 13873 35193
rect 13907 35159 13946 35193
rect 13980 35159 14019 35193
rect 14053 35159 14092 35193
rect 14126 35159 14165 35193
rect 14199 35159 14238 35193
rect 14272 35159 14311 35193
rect 14345 35159 14384 35193
rect 14418 35159 14429 35193
rect 13175 35121 14429 35159
rect 13175 35087 13216 35121
rect 13250 35087 13289 35121
rect 13323 35087 13362 35121
rect 13396 35087 13435 35121
rect 13469 35087 13508 35121
rect 13542 35087 13581 35121
rect 13615 35087 13654 35121
rect 13688 35087 13727 35121
rect 13761 35087 13800 35121
rect 13834 35087 13873 35121
rect 13907 35087 13946 35121
rect 13980 35087 14019 35121
rect 14053 35087 14092 35121
rect 14126 35087 14165 35121
rect 14199 35087 14238 35121
rect 14272 35087 14311 35121
rect 14345 35087 14384 35121
rect 14418 35087 14429 35121
rect 13175 35049 14429 35087
rect 13175 35015 13216 35049
rect 13250 35015 13289 35049
rect 13323 35015 13362 35049
rect 13396 35015 13435 35049
rect 13469 35015 13508 35049
rect 13542 35015 13581 35049
rect 13615 35015 13654 35049
rect 13688 35015 13727 35049
rect 13761 35015 13800 35049
rect 13834 35015 13873 35049
rect 13907 35015 13946 35049
rect 13980 35015 14019 35049
rect 14053 35015 14092 35049
rect 14126 35015 14165 35049
rect 14199 35015 14238 35049
rect 14272 35015 14311 35049
rect 14345 35015 14384 35049
rect 14418 35015 14429 35049
rect 13175 34977 14429 35015
rect 13175 34943 13216 34977
rect 13250 34943 13289 34977
rect 13323 34943 13362 34977
rect 13396 34943 13435 34977
rect 13469 34943 13508 34977
rect 13542 34943 13581 34977
rect 13615 34943 13654 34977
rect 13688 34943 13727 34977
rect 13761 34943 13800 34977
rect 13834 34943 13873 34977
rect 13907 34943 13946 34977
rect 13980 34943 14019 34977
rect 14053 34943 14092 34977
rect 14126 34943 14165 34977
rect 14199 34943 14238 34977
rect 14272 34943 14311 34977
rect 14345 34943 14384 34977
rect 14418 34943 14429 34977
rect 13175 34905 14429 34943
rect 13175 34871 13216 34905
rect 13250 34871 13289 34905
rect 13323 34871 13362 34905
rect 13396 34871 13435 34905
rect 13469 34871 13508 34905
rect 13542 34871 13581 34905
rect 13615 34871 13654 34905
rect 13688 34871 13727 34905
rect 13761 34871 13800 34905
rect 13834 34871 13873 34905
rect 13907 34871 13946 34905
rect 13980 34871 14019 34905
rect 14053 34871 14092 34905
rect 14126 34871 14165 34905
rect 14199 34871 14238 34905
rect 14272 34871 14311 34905
rect 14345 34871 14384 34905
rect 14418 34871 14429 34905
rect 13175 34833 14429 34871
rect 13175 34799 13216 34833
rect 13250 34799 13289 34833
rect 13323 34799 13362 34833
rect 13396 34799 13435 34833
rect 13469 34799 13508 34833
rect 13542 34799 13581 34833
rect 13615 34799 13654 34833
rect 13688 34799 13727 34833
rect 13761 34799 13800 34833
rect 13834 34799 13873 34833
rect 13907 34799 13946 34833
rect 13980 34799 14019 34833
rect 14053 34799 14092 34833
rect 14126 34799 14165 34833
rect 14199 34799 14238 34833
rect 14272 34799 14311 34833
rect 14345 34799 14384 34833
rect 14418 34799 14429 34833
rect 13175 34760 14429 34799
rect 13175 34726 13216 34760
rect 13250 34726 13289 34760
rect 13323 34726 13362 34760
rect 13396 34726 13435 34760
rect 13469 34726 13508 34760
rect 13542 34726 13581 34760
rect 13615 34726 13654 34760
rect 13688 34726 13727 34760
rect 13761 34726 13800 34760
rect 13834 34726 13873 34760
rect 13907 34726 13946 34760
rect 13980 34726 14019 34760
rect 14053 34726 14092 34760
rect 14126 34726 14165 34760
rect 14199 34726 14238 34760
rect 14272 34726 14311 34760
rect 14345 34726 14384 34760
rect 14418 34726 14429 34760
rect 13175 34687 14429 34726
rect 13175 34653 13216 34687
rect 13250 34653 13289 34687
rect 13323 34653 13362 34687
rect 13396 34653 13435 34687
rect 13469 34653 13508 34687
rect 13542 34653 13581 34687
rect 13615 34653 13654 34687
rect 13688 34653 13727 34687
rect 13761 34653 13800 34687
rect 13834 34653 13873 34687
rect 13907 34653 13946 34687
rect 13980 34653 14019 34687
rect 14053 34653 14092 34687
rect 14126 34653 14165 34687
rect 14199 34653 14238 34687
rect 14272 34653 14311 34687
rect 14345 34653 14384 34687
rect 14418 34653 14429 34687
rect 13175 34614 14429 34653
rect 13175 34580 13216 34614
rect 13250 34580 13289 34614
rect 13323 34580 13362 34614
rect 13396 34580 13435 34614
rect 13469 34580 13508 34614
rect 13542 34580 13581 34614
rect 13615 34580 13654 34614
rect 13688 34580 13727 34614
rect 13761 34580 13800 34614
rect 13834 34580 13873 34614
rect 13907 34580 13946 34614
rect 13980 34580 14019 34614
rect 14053 34580 14092 34614
rect 14126 34580 14165 34614
rect 14199 34580 14238 34614
rect 14272 34580 14311 34614
rect 14345 34580 14384 34614
rect 14418 34580 14429 34614
rect 13175 34541 14429 34580
rect 13175 34507 13216 34541
rect 13250 34507 13289 34541
rect 13323 34507 13362 34541
rect 13396 34507 13435 34541
rect 13469 34507 13508 34541
rect 13542 34507 13581 34541
rect 13615 34507 13654 34541
rect 13688 34507 13727 34541
rect 13761 34507 13800 34541
rect 13834 34507 13873 34541
rect 13907 34507 13946 34541
rect 13980 34507 14019 34541
rect 14053 34507 14092 34541
rect 14126 34507 14165 34541
rect 14199 34507 14238 34541
rect 14272 34507 14311 34541
rect 14345 34507 14384 34541
rect 14418 34507 14429 34541
rect 13175 34468 14429 34507
rect 13175 34434 13216 34468
rect 13250 34434 13289 34468
rect 13323 34434 13362 34468
rect 13396 34434 13435 34468
rect 13469 34434 13508 34468
rect 13542 34434 13581 34468
rect 13615 34434 13654 34468
rect 13688 34434 13727 34468
rect 13761 34434 13800 34468
rect 13834 34434 13873 34468
rect 13907 34434 13946 34468
rect 13980 34434 14019 34468
rect 14053 34434 14092 34468
rect 14126 34434 14165 34468
rect 14199 34434 14238 34468
rect 14272 34434 14311 34468
rect 14345 34434 14384 34468
rect 14418 34434 14429 34468
rect 13175 34395 14429 34434
rect 13175 34361 13216 34395
rect 13250 34361 13289 34395
rect 13323 34361 13362 34395
rect 13396 34361 13435 34395
rect 13469 34361 13508 34395
rect 13542 34361 13581 34395
rect 13615 34361 13654 34395
rect 13688 34361 13727 34395
rect 13761 34361 13800 34395
rect 13834 34361 13873 34395
rect 13907 34361 13946 34395
rect 13980 34361 14019 34395
rect 14053 34361 14092 34395
rect 14126 34361 14165 34395
rect 14199 34361 14238 34395
rect 14272 34361 14311 34395
rect 14345 34361 14384 34395
rect 14418 34361 14429 34395
rect 13175 34322 14429 34361
rect 13175 34288 13216 34322
rect 13250 34288 13289 34322
rect 13323 34288 13362 34322
rect 13396 34288 13435 34322
rect 13469 34288 13508 34322
rect 13542 34288 13581 34322
rect 13615 34288 13654 34322
rect 13688 34288 13727 34322
rect 13761 34288 13800 34322
rect 13834 34288 13873 34322
rect 13907 34288 13946 34322
rect 13980 34288 14019 34322
rect 14053 34288 14092 34322
rect 14126 34288 14165 34322
rect 14199 34288 14238 34322
rect 14272 34288 14311 34322
rect 14345 34288 14384 34322
rect 14418 34288 14429 34322
rect 13175 34249 14429 34288
rect 13175 34215 13216 34249
rect 13250 34215 13289 34249
rect 13323 34215 13362 34249
rect 13396 34215 13435 34249
rect 13469 34215 13508 34249
rect 13542 34215 13581 34249
rect 13615 34215 13654 34249
rect 13688 34215 13727 34249
rect 13761 34215 13800 34249
rect 13834 34215 13873 34249
rect 13907 34215 13946 34249
rect 13980 34215 14019 34249
rect 14053 34215 14092 34249
rect 14126 34215 14165 34249
rect 14199 34215 14238 34249
rect 14272 34215 14311 34249
rect 14345 34215 14384 34249
rect 14418 34215 14429 34249
rect 13175 34176 14429 34215
rect 13175 34142 13216 34176
rect 13250 34142 13289 34176
rect 13323 34142 13362 34176
rect 13396 34142 13435 34176
rect 13469 34142 13508 34176
rect 13542 34142 13581 34176
rect 13615 34142 13654 34176
rect 13688 34142 13727 34176
rect 13761 34142 13800 34176
rect 13834 34142 13873 34176
rect 13907 34142 13946 34176
rect 13980 34142 14019 34176
rect 14053 34142 14092 34176
rect 14126 34142 14165 34176
rect 14199 34142 14238 34176
rect 14272 34142 14311 34176
rect 14345 34142 14384 34176
rect 14418 34142 14429 34176
rect 13175 34103 14429 34142
rect 13175 34069 13216 34103
rect 13250 34069 13289 34103
rect 13323 34069 13362 34103
rect 13396 34069 13435 34103
rect 13469 34069 13508 34103
rect 13542 34069 13581 34103
rect 13615 34069 13654 34103
rect 13688 34069 13727 34103
rect 13761 34069 13800 34103
rect 13834 34069 13873 34103
rect 13907 34069 13946 34103
rect 13980 34069 14019 34103
rect 14053 34069 14092 34103
rect 14126 34069 14165 34103
rect 14199 34069 14238 34103
rect 14272 34069 14311 34103
rect 14345 34069 14384 34103
rect 14418 34069 14429 34103
rect 13175 34030 14429 34069
rect 13175 33996 13216 34030
rect 13250 33996 13289 34030
rect 13323 33996 13362 34030
rect 13396 33996 13435 34030
rect 13469 33996 13508 34030
rect 13542 33996 13581 34030
rect 13615 33996 13654 34030
rect 13688 33996 13727 34030
rect 13761 33996 13800 34030
rect 13834 33996 13873 34030
rect 13907 33996 13946 34030
rect 13980 33996 14019 34030
rect 14053 33996 14092 34030
rect 14126 33996 14165 34030
rect 14199 33996 14238 34030
rect 14272 33996 14311 34030
rect 14345 33996 14384 34030
rect 14418 33996 14429 34030
rect 13175 33957 14429 33996
rect 13175 33923 13216 33957
rect 13250 33923 13289 33957
rect 13323 33923 13362 33957
rect 13396 33923 13435 33957
rect 13469 33923 13508 33957
rect 13542 33923 13581 33957
rect 13615 33923 13654 33957
rect 13688 33923 13727 33957
rect 13761 33923 13800 33957
rect 13834 33923 13873 33957
rect 13907 33923 13946 33957
rect 13980 33923 14019 33957
rect 14053 33923 14092 33957
rect 14126 33923 14165 33957
rect 14199 33923 14238 33957
rect 14272 33923 14311 33957
rect 14345 33923 14384 33957
rect 14418 33923 14429 33957
rect 13175 33884 14429 33923
rect 13175 33850 13216 33884
rect 13250 33850 13289 33884
rect 13323 33850 13362 33884
rect 13396 33850 13435 33884
rect 13469 33850 13508 33884
rect 13542 33850 13581 33884
rect 13615 33850 13654 33884
rect 13688 33850 13727 33884
rect 13761 33850 13800 33884
rect 13834 33850 13873 33884
rect 13907 33850 13946 33884
rect 13980 33850 14019 33884
rect 14053 33850 14092 33884
rect 14126 33850 14165 33884
rect 14199 33850 14238 33884
rect 14272 33850 14311 33884
rect 14345 33850 14384 33884
rect 14418 33850 14429 33884
rect 13175 33811 14429 33850
rect 13175 33777 13216 33811
rect 13250 33777 13289 33811
rect 13323 33777 13362 33811
rect 13396 33777 13435 33811
rect 13469 33777 13508 33811
rect 13542 33777 13581 33811
rect 13615 33777 13654 33811
rect 13688 33777 13727 33811
rect 13761 33777 13800 33811
rect 13834 33777 13873 33811
rect 13907 33777 13946 33811
rect 13980 33777 14019 33811
rect 14053 33777 14092 33811
rect 14126 33777 14165 33811
rect 14199 33777 14238 33811
rect 14272 33777 14311 33811
rect 14345 33777 14384 33811
rect 14418 33777 14429 33811
rect 13175 33738 14429 33777
rect 13175 33704 13216 33738
rect 13250 33704 13289 33738
rect 13323 33704 13362 33738
rect 13396 33704 13435 33738
rect 13469 33704 13508 33738
rect 13542 33704 13581 33738
rect 13615 33704 13654 33738
rect 13688 33704 13727 33738
rect 13761 33704 13800 33738
rect 13834 33704 13873 33738
rect 13907 33704 13946 33738
rect 13980 33704 14019 33738
rect 14053 33704 14092 33738
rect 14126 33704 14165 33738
rect 14199 33704 14238 33738
rect 14272 33704 14311 33738
rect 14345 33704 14384 33738
rect 14418 33704 14429 33738
rect 13175 33665 14429 33704
rect 13175 33631 13216 33665
rect 13250 33631 13289 33665
rect 13323 33631 13362 33665
rect 13396 33631 13435 33665
rect 13469 33631 13508 33665
rect 13542 33631 13581 33665
rect 13615 33631 13654 33665
rect 13688 33631 13727 33665
rect 13761 33631 13800 33665
rect 13834 33631 13873 33665
rect 13907 33631 13946 33665
rect 13980 33631 14019 33665
rect 14053 33631 14092 33665
rect 14126 33631 14165 33665
rect 14199 33631 14238 33665
rect 14272 33631 14311 33665
rect 14345 33631 14384 33665
rect 14418 33631 14429 33665
rect 13175 33592 14429 33631
rect 13175 33558 13216 33592
rect 13250 33558 13289 33592
rect 13323 33558 13362 33592
rect 13396 33558 13435 33592
rect 13469 33558 13508 33592
rect 13542 33558 13581 33592
rect 13615 33558 13654 33592
rect 13688 33558 13727 33592
rect 13761 33558 13800 33592
rect 13834 33558 13873 33592
rect 13907 33558 13946 33592
rect 13980 33558 14019 33592
rect 14053 33558 14092 33592
rect 14126 33558 14165 33592
rect 14199 33558 14238 33592
rect 14272 33558 14311 33592
rect 14345 33558 14384 33592
rect 14418 33558 14429 33592
rect 13175 33519 14429 33558
rect 13175 33485 13216 33519
rect 13250 33485 13289 33519
rect 13323 33485 13362 33519
rect 13396 33485 13435 33519
rect 13469 33485 13508 33519
rect 13542 33485 13581 33519
rect 13615 33485 13654 33519
rect 13688 33485 13727 33519
rect 13761 33485 13800 33519
rect 13834 33485 13873 33519
rect 13907 33485 13946 33519
rect 13980 33485 14019 33519
rect 14053 33485 14092 33519
rect 14126 33485 14165 33519
rect 14199 33485 14238 33519
rect 14272 33485 14311 33519
rect 14345 33485 14384 33519
rect 14418 33485 14429 33519
rect 13175 33446 14429 33485
rect 13175 33412 13216 33446
rect 13250 33412 13289 33446
rect 13323 33412 13362 33446
rect 13396 33412 13435 33446
rect 13469 33412 13508 33446
rect 13542 33412 13581 33446
rect 13615 33412 13654 33446
rect 13688 33412 13727 33446
rect 13761 33412 13800 33446
rect 13834 33412 13873 33446
rect 13907 33412 13946 33446
rect 13980 33412 14019 33446
rect 14053 33412 14092 33446
rect 14126 33412 14165 33446
rect 14199 33412 14238 33446
rect 14272 33412 14311 33446
rect 14345 33412 14384 33446
rect 14418 33412 14429 33446
rect 13175 33373 14429 33412
rect 13175 33339 13216 33373
rect 13250 33339 13289 33373
rect 13323 33339 13362 33373
rect 13396 33339 13435 33373
rect 13469 33339 13508 33373
rect 13542 33339 13581 33373
rect 13615 33339 13654 33373
rect 13688 33339 13727 33373
rect 13761 33339 13800 33373
rect 13834 33339 13873 33373
rect 13907 33339 13946 33373
rect 13980 33339 14019 33373
rect 14053 33339 14092 33373
rect 14126 33339 14165 33373
rect 14199 33339 14238 33373
rect 14272 33339 14311 33373
rect 14345 33339 14384 33373
rect 14418 33339 14429 33373
rect 13175 33300 14429 33339
rect 13175 33266 13216 33300
rect 13250 33266 13289 33300
rect 13323 33266 13362 33300
rect 13396 33266 13435 33300
rect 13469 33266 13508 33300
rect 13542 33266 13581 33300
rect 13615 33266 13654 33300
rect 13688 33266 13727 33300
rect 13761 33266 13800 33300
rect 13834 33266 13873 33300
rect 13907 33266 13946 33300
rect 13980 33266 14019 33300
rect 14053 33266 14092 33300
rect 14126 33266 14165 33300
rect 14199 33266 14238 33300
rect 14272 33266 14311 33300
rect 14345 33266 14384 33300
rect 14418 33266 14429 33300
rect 13175 33227 14429 33266
rect 13175 33193 13216 33227
rect 13250 33193 13289 33227
rect 13323 33193 13362 33227
rect 13396 33193 13435 33227
rect 13469 33193 13508 33227
rect 13542 33193 13581 33227
rect 13615 33193 13654 33227
rect 13688 33193 13727 33227
rect 13761 33193 13800 33227
rect 13834 33193 13873 33227
rect 13907 33193 13946 33227
rect 13980 33193 14019 33227
rect 14053 33193 14092 33227
rect 14126 33193 14165 33227
rect 14199 33193 14238 33227
rect 14272 33193 14311 33227
rect 14345 33193 14384 33227
rect 14418 33193 14429 33227
rect 13175 33154 14429 33193
rect 13175 33120 13216 33154
rect 13250 33120 13289 33154
rect 13323 33120 13362 33154
rect 13396 33120 13435 33154
rect 13469 33120 13508 33154
rect 13542 33120 13581 33154
rect 13615 33120 13654 33154
rect 13688 33120 13727 33154
rect 13761 33120 13800 33154
rect 13834 33120 13873 33154
rect 13907 33120 13946 33154
rect 13980 33120 14019 33154
rect 14053 33120 14092 33154
rect 14126 33120 14165 33154
rect 14199 33120 14238 33154
rect 14272 33120 14311 33154
rect 14345 33120 14384 33154
rect 14418 33120 14429 33154
rect 13175 33081 14429 33120
rect 13175 33047 13216 33081
rect 13250 33047 13289 33081
rect 13323 33047 13362 33081
rect 13396 33047 13435 33081
rect 13469 33047 13508 33081
rect 13542 33047 13581 33081
rect 13615 33047 13654 33081
rect 13688 33047 13727 33081
rect 13761 33047 13800 33081
rect 13834 33047 13873 33081
rect 13907 33047 13946 33081
rect 13980 33047 14019 33081
rect 14053 33047 14092 33081
rect 14126 33047 14165 33081
rect 14199 33047 14238 33081
rect 14272 33047 14311 33081
rect 14345 33047 14384 33081
rect 14418 33047 14429 33081
rect 13175 33008 14429 33047
rect 13175 32974 13216 33008
rect 13250 32974 13289 33008
rect 13323 32974 13362 33008
rect 13396 32974 13435 33008
rect 13469 32974 13508 33008
rect 13542 32974 13581 33008
rect 13615 32974 13654 33008
rect 13688 32974 13727 33008
rect 13761 32974 13800 33008
rect 13834 32974 13873 33008
rect 13907 32974 13946 33008
rect 13980 32974 14019 33008
rect 14053 32974 14092 33008
rect 14126 32974 14165 33008
rect 14199 32974 14238 33008
rect 14272 32974 14311 33008
rect 14345 32974 14384 33008
rect 14418 32974 14429 33008
rect 13175 32935 14429 32974
rect 13175 32901 13216 32935
rect 13250 32901 13289 32935
rect 13323 32901 13362 32935
rect 13396 32901 13435 32935
rect 13469 32901 13508 32935
rect 13542 32901 13581 32935
rect 13615 32901 13654 32935
rect 13688 32901 13727 32935
rect 13761 32901 13800 32935
rect 13834 32901 13873 32935
rect 13907 32901 13946 32935
rect 13980 32901 14019 32935
rect 14053 32901 14092 32935
rect 14126 32901 14165 32935
rect 14199 32901 14238 32935
rect 14272 32901 14311 32935
rect 14345 32901 14384 32935
rect 14418 32901 14429 32935
rect 13175 32862 14429 32901
rect 13175 32828 13216 32862
rect 13250 32828 13289 32862
rect 13323 32828 13362 32862
rect 13396 32828 13435 32862
rect 13469 32828 13508 32862
rect 13542 32828 13581 32862
rect 13615 32828 13654 32862
rect 13688 32828 13727 32862
rect 13761 32828 13800 32862
rect 13834 32828 13873 32862
rect 13907 32828 13946 32862
rect 13980 32828 14019 32862
rect 14053 32828 14092 32862
rect 14126 32828 14165 32862
rect 14199 32828 14238 32862
rect 14272 32828 14311 32862
rect 14345 32828 14384 32862
rect 14418 32828 14429 32862
rect 13175 32789 14429 32828
rect 13175 32755 13216 32789
rect 13250 32755 13289 32789
rect 13323 32755 13362 32789
rect 13396 32755 13435 32789
rect 13469 32755 13508 32789
rect 13542 32755 13581 32789
rect 13615 32755 13654 32789
rect 13688 32755 13727 32789
rect 13761 32755 13800 32789
rect 13834 32755 13873 32789
rect 13907 32755 13946 32789
rect 13980 32755 14019 32789
rect 14053 32755 14092 32789
rect 14126 32755 14165 32789
rect 14199 32755 14238 32789
rect 14272 32755 14311 32789
rect 14345 32755 14384 32789
rect 14418 32755 14429 32789
rect 13175 32716 14429 32755
rect 13175 32682 13216 32716
rect 13250 32682 13289 32716
rect 13323 32682 13362 32716
rect 13396 32682 13435 32716
rect 13469 32682 13508 32716
rect 13542 32682 13581 32716
rect 13615 32682 13654 32716
rect 13688 32682 13727 32716
rect 13761 32682 13800 32716
rect 13834 32682 13873 32716
rect 13907 32682 13946 32716
rect 13980 32682 14019 32716
rect 14053 32682 14092 32716
rect 14126 32682 14165 32716
rect 14199 32682 14238 32716
rect 14272 32682 14311 32716
rect 14345 32682 14384 32716
rect 14418 32682 14429 32716
rect 13175 32643 14429 32682
rect 13175 32609 13216 32643
rect 13250 32609 13289 32643
rect 13323 32609 13362 32643
rect 13396 32609 13435 32643
rect 13469 32609 13508 32643
rect 13542 32609 13581 32643
rect 13615 32609 13654 32643
rect 13688 32609 13727 32643
rect 13761 32609 13800 32643
rect 13834 32609 13873 32643
rect 13907 32609 13946 32643
rect 13980 32609 14019 32643
rect 14053 32609 14092 32643
rect 14126 32609 14165 32643
rect 14199 32609 14238 32643
rect 14272 32609 14311 32643
rect 14345 32609 14384 32643
rect 14418 32609 14429 32643
rect 13175 32570 14429 32609
rect 13175 32536 13216 32570
rect 13250 32536 13289 32570
rect 13323 32536 13362 32570
rect 13396 32536 13435 32570
rect 13469 32536 13508 32570
rect 13542 32536 13581 32570
rect 13615 32536 13654 32570
rect 13688 32536 13727 32570
rect 13761 32536 13800 32570
rect 13834 32536 13873 32570
rect 13907 32536 13946 32570
rect 13980 32536 14019 32570
rect 14053 32536 14092 32570
rect 14126 32536 14165 32570
rect 14199 32536 14238 32570
rect 14272 32536 14311 32570
rect 14345 32536 14384 32570
rect 14418 32536 14429 32570
rect 13175 32497 14429 32536
rect 13175 32463 13216 32497
rect 13250 32463 13289 32497
rect 13323 32463 13362 32497
rect 13396 32463 13435 32497
rect 13469 32463 13508 32497
rect 13542 32463 13581 32497
rect 13615 32463 13654 32497
rect 13688 32463 13727 32497
rect 13761 32463 13800 32497
rect 13834 32463 13873 32497
rect 13907 32463 13946 32497
rect 13980 32463 14019 32497
rect 14053 32463 14092 32497
rect 14126 32463 14165 32497
rect 14199 32463 14238 32497
rect 14272 32463 14311 32497
rect 14345 32463 14384 32497
rect 14418 32463 14429 32497
rect 13175 32424 14429 32463
rect 13175 32390 13216 32424
rect 13250 32390 13289 32424
rect 13323 32390 13362 32424
rect 13396 32390 13435 32424
rect 13469 32390 13508 32424
rect 13542 32390 13581 32424
rect 13615 32390 13654 32424
rect 13688 32390 13727 32424
rect 13761 32390 13800 32424
rect 13834 32390 13873 32424
rect 13907 32390 13946 32424
rect 13980 32390 14019 32424
rect 14053 32390 14092 32424
rect 14126 32390 14165 32424
rect 14199 32390 14238 32424
rect 14272 32390 14311 32424
rect 14345 32390 14384 32424
rect 14418 32390 14429 32424
rect 13175 32351 14429 32390
rect 13175 32317 13216 32351
rect 13250 32317 13289 32351
rect 13323 32317 13362 32351
rect 13396 32317 13435 32351
rect 13469 32317 13508 32351
rect 13542 32317 13581 32351
rect 13615 32317 13654 32351
rect 13688 32317 13727 32351
rect 13761 32317 13800 32351
rect 13834 32317 13873 32351
rect 13907 32317 13946 32351
rect 13980 32317 14019 32351
rect 14053 32317 14092 32351
rect 14126 32317 14165 32351
rect 14199 32317 14238 32351
rect 14272 32317 14311 32351
rect 14345 32317 14384 32351
rect 14418 32317 14429 32351
rect 13175 32278 14429 32317
rect 13175 32244 13216 32278
rect 13250 32244 13289 32278
rect 13323 32244 13362 32278
rect 13396 32244 13435 32278
rect 13469 32244 13508 32278
rect 13542 32244 13581 32278
rect 13615 32244 13654 32278
rect 13688 32244 13727 32278
rect 13761 32244 13800 32278
rect 13834 32244 13873 32278
rect 13907 32244 13946 32278
rect 13980 32244 14019 32278
rect 14053 32244 14092 32278
rect 14126 32244 14165 32278
rect 14199 32244 14238 32278
rect 14272 32244 14311 32278
rect 14345 32244 14384 32278
rect 14418 32244 14429 32278
rect 13175 32205 14429 32244
rect 13175 32171 13216 32205
rect 13250 32171 13289 32205
rect 13323 32171 13362 32205
rect 13396 32171 13435 32205
rect 13469 32171 13508 32205
rect 13542 32171 13581 32205
rect 13615 32171 13654 32205
rect 13688 32171 13727 32205
rect 13761 32171 13800 32205
rect 13834 32171 13873 32205
rect 13907 32171 13946 32205
rect 13980 32171 14019 32205
rect 14053 32171 14092 32205
rect 14126 32171 14165 32205
rect 14199 32171 14238 32205
rect 14272 32171 14311 32205
rect 14345 32171 14384 32205
rect 14418 32171 14429 32205
rect 13175 32132 14429 32171
rect 13175 32098 13216 32132
rect 13250 32098 13289 32132
rect 13323 32098 13362 32132
rect 13396 32098 13435 32132
rect 13469 32098 13508 32132
rect 13542 32098 13581 32132
rect 13615 32098 13654 32132
rect 13688 32098 13727 32132
rect 13761 32098 13800 32132
rect 13834 32098 13873 32132
rect 13907 32098 13946 32132
rect 13980 32098 14019 32132
rect 14053 32098 14092 32132
rect 14126 32098 14165 32132
rect 14199 32098 14238 32132
rect 14272 32098 14311 32132
rect 14345 32098 14384 32132
rect 14418 32098 14429 32132
rect 13175 32059 14429 32098
rect 13175 32025 13216 32059
rect 13250 32025 13289 32059
rect 13323 32025 13362 32059
rect 13396 32025 13435 32059
rect 13469 32025 13508 32059
rect 13542 32025 13581 32059
rect 13615 32025 13654 32059
rect 13688 32025 13727 32059
rect 13761 32025 13800 32059
rect 13834 32025 13873 32059
rect 13907 32025 13946 32059
rect 13980 32025 14019 32059
rect 14053 32025 14092 32059
rect 14126 32025 14165 32059
rect 14199 32025 14238 32059
rect 14272 32025 14311 32059
rect 14345 32025 14384 32059
rect 14418 32025 14429 32059
rect 13175 31986 14429 32025
rect 13175 31952 13216 31986
rect 13250 31952 13289 31986
rect 13323 31952 13362 31986
rect 13396 31952 13435 31986
rect 13469 31952 13508 31986
rect 13542 31952 13581 31986
rect 13615 31952 13654 31986
rect 13688 31952 13727 31986
rect 13761 31952 13800 31986
rect 13834 31952 13873 31986
rect 13907 31952 13946 31986
rect 13980 31952 14019 31986
rect 14053 31952 14092 31986
rect 14126 31952 14165 31986
rect 14199 31952 14238 31986
rect 14272 31952 14311 31986
rect 14345 31952 14384 31986
rect 14418 31952 14429 31986
rect 13175 31913 14429 31952
rect 13175 31879 13216 31913
rect 13250 31879 13289 31913
rect 13323 31879 13362 31913
rect 13396 31879 13435 31913
rect 13469 31879 13508 31913
rect 13542 31879 13581 31913
rect 13615 31879 13654 31913
rect 13688 31879 13727 31913
rect 13761 31879 13800 31913
rect 13834 31879 13873 31913
rect 13907 31879 13946 31913
rect 13980 31879 14019 31913
rect 14053 31879 14092 31913
rect 14126 31879 14165 31913
rect 14199 31879 14238 31913
rect 14272 31879 14311 31913
rect 14345 31879 14384 31913
rect 14418 31879 14429 31913
rect 13175 31840 14429 31879
rect 13175 31806 13216 31840
rect 13250 31806 13289 31840
rect 13323 31806 13362 31840
rect 13396 31806 13435 31840
rect 13469 31806 13508 31840
rect 13542 31806 13581 31840
rect 13615 31806 13654 31840
rect 13688 31806 13727 31840
rect 13761 31806 13800 31840
rect 13834 31806 13873 31840
rect 13907 31806 13946 31840
rect 13980 31806 14019 31840
rect 14053 31806 14092 31840
rect 14126 31806 14165 31840
rect 14199 31806 14238 31840
rect 14272 31806 14311 31840
rect 14345 31806 14384 31840
rect 14418 31806 14429 31840
rect 13175 31767 14429 31806
rect 13175 31733 13216 31767
rect 13250 31733 13289 31767
rect 13323 31733 13362 31767
rect 13396 31733 13435 31767
rect 13469 31733 13508 31767
rect 13542 31733 13581 31767
rect 13615 31733 13654 31767
rect 13688 31733 13727 31767
rect 13761 31733 13800 31767
rect 13834 31733 13873 31767
rect 13907 31733 13946 31767
rect 13980 31733 14019 31767
rect 14053 31733 14092 31767
rect 14126 31733 14165 31767
rect 14199 31733 14238 31767
rect 14272 31733 14311 31767
rect 14345 31733 14384 31767
rect 14418 31733 14429 31767
rect 13175 31694 14429 31733
rect 13175 31660 13216 31694
rect 13250 31660 13289 31694
rect 13323 31660 13362 31694
rect 13396 31660 13435 31694
rect 13469 31660 13508 31694
rect 13542 31660 13581 31694
rect 13615 31660 13654 31694
rect 13688 31660 13727 31694
rect 13761 31660 13800 31694
rect 13834 31660 13873 31694
rect 13907 31660 13946 31694
rect 13980 31660 14019 31694
rect 14053 31660 14092 31694
rect 14126 31660 14165 31694
rect 14199 31660 14238 31694
rect 14272 31660 14311 31694
rect 14345 31660 14384 31694
rect 14418 31660 14429 31694
rect 13175 31621 14429 31660
rect 13175 31587 13216 31621
rect 13250 31587 13289 31621
rect 13323 31587 13362 31621
rect 13396 31587 13435 31621
rect 13469 31587 13508 31621
rect 13542 31587 13581 31621
rect 13615 31587 13654 31621
rect 13688 31587 13727 31621
rect 13761 31587 13800 31621
rect 13834 31587 13873 31621
rect 13907 31587 13946 31621
rect 13980 31587 14019 31621
rect 14053 31587 14092 31621
rect 14126 31587 14165 31621
rect 14199 31587 14238 31621
rect 14272 31587 14311 31621
rect 14345 31587 14384 31621
rect 14418 31587 14429 31621
rect 13175 31548 14429 31587
rect 13175 31514 13216 31548
rect 13250 31514 13289 31548
rect 13323 31514 13362 31548
rect 13396 31514 13435 31548
rect 13469 31514 13508 31548
rect 13542 31514 13581 31548
rect 13615 31514 13654 31548
rect 13688 31514 13727 31548
rect 13761 31514 13800 31548
rect 13834 31514 13873 31548
rect 13907 31514 13946 31548
rect 13980 31514 14019 31548
rect 14053 31514 14092 31548
rect 14126 31514 14165 31548
rect 14199 31514 14238 31548
rect 14272 31514 14311 31548
rect 14345 31514 14384 31548
rect 14418 31514 14429 31548
rect 13175 31475 14429 31514
rect 13175 31441 13216 31475
rect 13250 31441 13289 31475
rect 13323 31441 13362 31475
rect 13396 31441 13435 31475
rect 13469 31441 13508 31475
rect 13542 31441 13581 31475
rect 13615 31441 13654 31475
rect 13688 31441 13727 31475
rect 13761 31441 13800 31475
rect 13834 31441 13873 31475
rect 13907 31441 13946 31475
rect 13980 31441 14019 31475
rect 14053 31441 14092 31475
rect 14126 31441 14165 31475
rect 14199 31441 14238 31475
rect 14272 31441 14311 31475
rect 14345 31441 14384 31475
rect 14418 31441 14429 31475
rect 13175 31402 14429 31441
rect 13175 31368 13216 31402
rect 13250 31368 13289 31402
rect 13323 31368 13362 31402
rect 13396 31368 13435 31402
rect 13469 31368 13508 31402
rect 13542 31368 13581 31402
rect 13615 31368 13654 31402
rect 13688 31368 13727 31402
rect 13761 31368 13800 31402
rect 13834 31368 13873 31402
rect 13907 31368 13946 31402
rect 13980 31368 14019 31402
rect 14053 31368 14092 31402
rect 14126 31368 14165 31402
rect 14199 31368 14238 31402
rect 14272 31368 14311 31402
rect 14345 31368 14384 31402
rect 14418 31368 14429 31402
rect 13175 31329 14429 31368
rect 13175 31295 13216 31329
rect 13250 31295 13289 31329
rect 13323 31295 13362 31329
rect 13396 31295 13435 31329
rect 13469 31295 13508 31329
rect 13542 31295 13581 31329
rect 13615 31295 13654 31329
rect 13688 31295 13727 31329
rect 13761 31295 13800 31329
rect 13834 31295 13873 31329
rect 13907 31295 13946 31329
rect 13980 31295 14019 31329
rect 14053 31295 14092 31329
rect 14126 31295 14165 31329
rect 14199 31295 14238 31329
rect 14272 31295 14311 31329
rect 14345 31295 14384 31329
rect 14418 31295 14429 31329
rect 13175 31256 14429 31295
rect 13175 31222 13216 31256
rect 13250 31222 13289 31256
rect 13323 31222 13362 31256
rect 13396 31222 13435 31256
rect 13469 31222 13508 31256
rect 13542 31222 13581 31256
rect 13615 31222 13654 31256
rect 13688 31222 13727 31256
rect 13761 31222 13800 31256
rect 13834 31222 13873 31256
rect 13907 31222 13946 31256
rect 13980 31222 14019 31256
rect 14053 31222 14092 31256
rect 14126 31222 14165 31256
rect 14199 31222 14238 31256
rect 14272 31222 14311 31256
rect 14345 31222 14384 31256
rect 14418 31222 14429 31256
rect 13175 31183 14429 31222
rect 13175 31149 13216 31183
rect 13250 31149 13289 31183
rect 13323 31149 13362 31183
rect 13396 31149 13435 31183
rect 13469 31149 13508 31183
rect 13542 31149 13581 31183
rect 13615 31149 13654 31183
rect 13688 31149 13727 31183
rect 13761 31149 13800 31183
rect 13834 31149 13873 31183
rect 13907 31149 13946 31183
rect 13980 31149 14019 31183
rect 14053 31149 14092 31183
rect 14126 31149 14165 31183
rect 14199 31149 14238 31183
rect 14272 31149 14311 31183
rect 14345 31149 14384 31183
rect 14418 31149 14429 31183
rect 13175 31137 14429 31149
tri 13012 30997 13050 31035 sw
rect 13012 30991 14270 30997
rect 13012 30957 13051 30991
rect 13085 30957 13124 30991
rect 13158 30957 13197 30991
rect 13231 30957 13270 30991
rect 13304 30957 13344 30991
rect 13378 30957 13418 30991
rect 13452 30957 13492 30991
rect 13526 30957 13566 30991
rect 13600 30957 13640 30991
rect 13674 30957 13714 30991
rect 13748 30957 13788 30991
rect 13822 30957 13862 30991
rect 13896 30957 13936 30991
rect 13970 30957 14010 30991
rect 14044 30957 14084 30991
rect 14118 30957 14158 30991
rect 14192 30957 14270 30991
rect 13012 30919 14270 30957
rect 13012 30885 14230 30919
rect 14264 30885 14270 30919
rect 13012 30863 14270 30885
rect 13012 30829 13051 30863
rect 13085 30829 13126 30863
rect 13160 30829 13201 30863
rect 13235 30829 13276 30863
rect 13310 30829 13351 30863
rect 13385 30829 13426 30863
rect 13460 30829 13501 30863
rect 13535 30829 13576 30863
rect 13610 30829 13651 30863
rect 13685 30829 13726 30863
rect 13760 30829 13801 30863
rect 13835 30829 13876 30863
rect 13910 30829 13951 30863
rect 13985 30829 14026 30863
rect 14060 30829 14102 30863
rect 14136 30847 14270 30863
rect 14136 30829 14230 30847
rect 13012 30823 14230 30829
rect 9699 30813 9854 30823
tri 9854 30813 9864 30823 nw
tri 13931 30813 13941 30823 ne
rect 13941 30813 14230 30823
rect 14264 30813 14270 30847
rect 9699 30791 9832 30813
tri 9832 30791 9854 30813 nw
tri 13941 30791 13963 30813 ne
rect 13963 30791 14270 30813
rect 9699 30757 9798 30791
tri 9798 30757 9832 30791 nw
tri 13963 30757 13997 30791 ne
rect 13997 30757 14102 30791
rect 14136 30775 14270 30791
rect 14136 30757 14230 30775
rect 9699 30741 9782 30757
tri 9782 30741 9798 30757 nw
tri 13997 30741 14013 30757 ne
rect 14013 30741 14230 30757
rect 14264 30741 14270 30775
rect 9699 30719 9760 30741
tri 9760 30719 9782 30741 nw
tri 14013 30719 14035 30741 ne
rect 14035 30719 14270 30741
rect 9699 30685 9726 30719
tri 9726 30685 9760 30719 nw
tri 14035 30685 14069 30719 ne
rect 14069 30685 14102 30719
rect 14136 30703 14270 30719
rect 14136 30685 14230 30703
rect 9699 30670 9711 30685
tri 9711 30670 9726 30685 nw
tri 14069 30670 14084 30685 ne
rect 14084 30670 14230 30685
rect 9699 30669 9710 30670
tri 9710 30669 9711 30670 nw
rect 9699 30664 9705 30669
tri 9705 30664 9710 30669 nw
rect 9901 30664 13950 30670
tri 14084 30669 14085 30670 ne
rect 14085 30669 14230 30670
rect 14264 30669 14270 30703
tri 9699 30658 9705 30664 nw
rect 9901 30630 10246 30664
rect 10280 30630 10320 30664
rect 10354 30630 10394 30664
rect 10428 30630 10467 30664
rect 10501 30630 10540 30664
rect 10574 30630 10613 30664
rect 10647 30630 10686 30664
rect 10720 30630 10759 30664
rect 10793 30630 10832 30664
rect 10866 30630 10905 30664
rect 10939 30630 10978 30664
rect 11012 30630 11051 30664
rect 11085 30630 11124 30664
rect 11158 30630 11197 30664
rect 11231 30630 11270 30664
rect 11304 30630 11343 30664
rect 11377 30630 11416 30664
rect 11450 30630 11489 30664
rect 11523 30630 11562 30664
rect 11596 30630 11635 30664
rect 11669 30630 11708 30664
rect 11742 30630 11781 30664
rect 11815 30630 11854 30664
rect 11888 30630 11927 30664
rect 11961 30630 12000 30664
rect 12034 30630 12073 30664
rect 12107 30630 12146 30664
rect 12180 30630 12219 30664
rect 12253 30630 12292 30664
rect 12326 30630 12365 30664
rect 12399 30630 12438 30664
rect 12472 30630 12511 30664
rect 12545 30630 12584 30664
rect 12618 30630 12657 30664
rect 12691 30630 12730 30664
rect 12764 30630 12803 30664
rect 12837 30630 12876 30664
rect 12910 30630 12949 30664
rect 12983 30630 13022 30664
rect 13056 30630 13095 30664
rect 13129 30630 13168 30664
rect 13202 30630 13241 30664
rect 13275 30630 13314 30664
rect 13348 30630 13387 30664
rect 13421 30630 13460 30664
rect 13494 30630 13533 30664
rect 13567 30630 13606 30664
rect 13640 30630 13679 30664
rect 13713 30630 13752 30664
rect 13786 30630 13825 30664
rect 13859 30630 13898 30664
rect 13932 30630 13950 30664
tri 14085 30658 14096 30669 ne
rect 9901 30557 13950 30630
rect 9901 30523 10246 30557
rect 10280 30523 10320 30557
rect 10354 30523 10394 30557
rect 10428 30523 10467 30557
rect 10501 30523 10540 30557
rect 10574 30523 10613 30557
rect 10647 30523 10686 30557
rect 10720 30523 10759 30557
rect 10793 30523 10832 30557
rect 10866 30523 10905 30557
rect 10939 30523 10978 30557
rect 11012 30523 11051 30557
rect 11085 30523 11124 30557
rect 11158 30523 11197 30557
rect 11231 30523 11270 30557
rect 11304 30523 11343 30557
rect 11377 30523 11416 30557
rect 11450 30523 11489 30557
rect 11523 30523 11562 30557
rect 11596 30523 11635 30557
rect 11669 30523 11708 30557
rect 11742 30523 11781 30557
rect 11815 30523 11854 30557
rect 11888 30523 11927 30557
rect 11961 30523 12000 30557
rect 12034 30523 12073 30557
rect 12107 30523 12146 30557
rect 12180 30523 12219 30557
rect 12253 30523 12292 30557
rect 12326 30523 12365 30557
rect 12399 30523 12438 30557
rect 12472 30523 12511 30557
rect 12545 30523 12584 30557
rect 12618 30523 12657 30557
rect 12691 30523 12730 30557
rect 12764 30523 12803 30557
rect 12837 30523 12876 30557
rect 12910 30523 12949 30557
rect 12983 30523 13022 30557
rect 13056 30523 13095 30557
rect 13129 30523 13168 30557
rect 13202 30523 13241 30557
rect 13275 30523 13314 30557
rect 13348 30523 13387 30557
rect 13421 30523 13460 30557
rect 13494 30523 13533 30557
rect 13567 30523 13606 30557
rect 13640 30523 13679 30557
rect 13713 30523 13752 30557
rect 13786 30523 13825 30557
rect 13859 30523 13898 30557
rect 13932 30523 13950 30557
rect 9901 30450 13950 30523
rect 9901 30416 10246 30450
rect 10280 30416 10320 30450
rect 10354 30416 10394 30450
rect 10428 30416 10467 30450
rect 10501 30416 10540 30450
rect 10574 30416 10613 30450
rect 10647 30416 10686 30450
rect 10720 30416 10759 30450
rect 10793 30416 10832 30450
rect 10866 30416 10905 30450
rect 10939 30416 10978 30450
rect 11012 30416 11051 30450
rect 11085 30416 11124 30450
rect 11158 30416 11197 30450
rect 11231 30416 11270 30450
rect 11304 30416 11343 30450
rect 11377 30416 11416 30450
rect 11450 30416 11489 30450
rect 11523 30416 11562 30450
rect 11596 30416 11635 30450
rect 11669 30416 11708 30450
rect 11742 30416 11781 30450
rect 11815 30416 11854 30450
rect 11888 30416 11927 30450
rect 11961 30416 12000 30450
rect 12034 30416 12073 30450
rect 12107 30416 12146 30450
rect 12180 30416 12219 30450
rect 12253 30416 12292 30450
rect 12326 30416 12365 30450
rect 12399 30416 12438 30450
rect 12472 30416 12511 30450
rect 12545 30416 12584 30450
rect 12618 30416 12657 30450
rect 12691 30416 12730 30450
rect 12764 30416 12803 30450
rect 12837 30416 12876 30450
rect 12910 30416 12949 30450
rect 12983 30416 13022 30450
rect 13056 30416 13095 30450
rect 13129 30416 13168 30450
rect 13202 30416 13241 30450
rect 13275 30416 13314 30450
rect 13348 30416 13387 30450
rect 13421 30416 13460 30450
rect 13494 30416 13533 30450
rect 13567 30416 13606 30450
rect 13640 30416 13679 30450
rect 13713 30416 13752 30450
rect 13786 30416 13825 30450
rect 13859 30416 13898 30450
rect 13932 30416 13950 30450
rect 9901 30410 13950 30416
rect 9901 30397 10400 30410
tri 10400 30397 10413 30410 nw
tri 13456 30397 13469 30410 ne
rect 13469 30397 13950 30410
rect 9901 30386 10389 30397
tri 10389 30386 10400 30397 nw
tri 13469 30386 13480 30397 ne
rect 13480 30386 13950 30397
rect 9901 30381 10384 30386
tri 10384 30381 10389 30386 nw
tri 13480 30381 13485 30386 ne
rect 13485 30381 13950 30386
rect 9901 30374 10377 30381
tri 10377 30374 10384 30381 nw
tri 13485 30374 13492 30381 ne
rect 13492 30374 13950 30381
rect 9901 30340 10343 30374
tri 10343 30340 10377 30374 nw
tri 13492 30340 13526 30374 ne
rect 13526 30340 13705 30374
rect 13739 30340 13807 30374
rect 13841 30340 13909 30374
rect 13943 30340 13950 30374
rect 9901 30325 10328 30340
tri 10328 30325 10343 30340 nw
tri 13526 30325 13541 30340 ne
rect 13541 30325 13950 30340
rect 9901 30309 10312 30325
tri 10312 30309 10328 30325 nw
tri 13541 30309 13557 30325 ne
rect 13557 30309 13950 30325
rect 9901 30301 10304 30309
tri 10304 30301 10312 30309 nw
tri 13557 30301 13565 30309 ne
rect 13565 30301 13950 30309
rect 9901 30267 10270 30301
tri 10270 30267 10304 30301 nw
tri 13565 30267 13599 30301 ne
rect 13599 30267 13705 30301
rect 13739 30300 13909 30301
rect 13739 30267 13807 30300
rect 9901 30266 10269 30267
tri 10269 30266 10270 30267 nw
tri 13599 30266 13600 30267 ne
rect 13600 30266 13807 30267
rect 13841 30267 13909 30300
rect 13943 30267 13950 30301
rect 13841 30266 13950 30267
rect 9901 30253 10256 30266
tri 10256 30253 10269 30266 nw
tri 13600 30253 13613 30266 ne
rect 13613 30253 13950 30266
rect 9901 30237 10240 30253
tri 10240 30237 10256 30253 nw
tri 13613 30237 13629 30253 ne
rect 13629 30237 13950 30253
rect 9901 30228 10231 30237
tri 10231 30228 10240 30237 nw
tri 13629 30228 13638 30237 ne
rect 13638 30228 13950 30237
rect -12267 29874 -11883 29955
rect -10936 29951 -10744 30003
rect -10112 29907 -9920 29940
tri 5506 29907 5519 29920 sw
rect 5506 29902 5519 29907
tri 5519 29902 5524 29907 sw
rect 5506 29899 5524 29902
tri 5524 29899 5527 29902 sw
rect 5506 29895 5527 29899
tri 5527 29895 5531 29899 sw
rect 4679 29857 4795 29863
rect -16902 29735 -16786 29787
rect -16515 29705 -16414 29772
rect -16009 29699 -15957 29734
rect -15929 29699 -15877 29734
rect -10716 29727 -10348 29823
rect -9779 29727 -9032 29781
rect -8541 29755 -7795 29809
rect -7622 29727 -5887 29781
rect -5656 29755 -4910 29809
rect -4418 29755 -3672 29809
rect -3493 29727 -1757 29781
rect -1534 29755 -787 29809
rect -296 29755 450 29809
rect 4731 29805 4743 29857
rect 4679 29799 4795 29805
rect 5097 29857 5213 29863
rect 5149 29805 5161 29857
rect 5097 29799 5213 29805
rect 5243 29857 5359 29863
rect 5295 29805 5307 29857
rect 5243 29799 5359 29805
rect 639 29727 1600 29781
rect 5388 29767 8391 29895
tri 8838 29572 8848 29582 se
rect 8848 29572 8900 29815
rect 8928 29733 8980 29844
rect 8928 29669 8980 29681
rect 8928 29611 8980 29617
rect 9008 29733 9060 29842
rect 9008 29669 9060 29681
rect 9008 29611 9060 29617
tri 9078 29589 9088 29599 se
rect 9088 29589 9140 29815
tri 9061 29572 9078 29589 se
rect 9078 29577 9140 29589
rect 9078 29572 9135 29577
tri 9135 29572 9140 29577 nw
tri 8837 29571 8838 29572 se
rect 8838 29571 8900 29572
tri 9060 29571 9061 29572 se
rect 9061 29571 9134 29572
tri 9134 29571 9135 29572 nw
tri 8823 29557 8837 29571 se
rect 8837 29557 8900 29571
tri 2076 29541 2092 29557 se
rect 2092 29541 2098 29557
rect 1664 29537 1733 29541
tri 1733 29537 1737 29541 sw
tri 2072 29537 2076 29541 se
rect 2076 29537 2098 29541
rect 1664 29535 1737 29537
rect 1664 29489 1680 29535
tri 1664 29477 1676 29489 ne
rect 1676 29483 1680 29489
rect 1732 29534 1737 29535
tri 1737 29534 1740 29537 sw
tri 2069 29534 2072 29537 se
rect 2072 29534 2098 29537
rect 1732 29529 1740 29534
tri 1740 29529 1745 29534 sw
tri 2064 29529 2069 29534 se
rect 2069 29529 2098 29534
rect 1732 29527 1745 29529
tri 1745 29527 1747 29529 sw
rect 1732 29517 1747 29527
tri 1747 29517 1757 29527 sw
rect 2034 29523 2098 29529
rect 1732 29510 1757 29517
tri 1757 29510 1764 29517 sw
rect 1732 29500 1764 29510
tri 1764 29500 1774 29510 sw
rect 1732 29498 1774 29500
tri 1774 29498 1776 29500 sw
rect 1732 29483 1776 29498
tri 1776 29483 1791 29498 sw
rect 1676 29478 1791 29483
rect 1676 29477 1733 29478
tri 1676 29465 1688 29477 ne
rect 1688 29465 1733 29477
tri 1688 29464 1689 29465 ne
rect 1689 29464 1733 29465
tri 1689 29461 1692 29464 ne
rect 1692 29461 1733 29464
tri 1692 29454 1699 29461 ne
rect 1699 29454 1733 29461
tri 1699 29445 1708 29454 ne
rect 1708 29445 1733 29454
tri 1708 29428 1725 29445 ne
rect 1725 29428 1733 29445
tri 1725 29426 1727 29428 ne
rect 1727 29426 1733 29428
rect 1785 29426 1791 29478
rect 2086 29505 2098 29523
rect 2150 29505 7564 29557
rect 7616 29505 7628 29557
rect 7680 29505 7686 29557
rect 7998 29505 8004 29557
rect 8056 29505 8068 29557
rect 8120 29554 8900 29557
rect 8120 29537 8883 29554
tri 8883 29537 8900 29554 nw
tri 9026 29537 9060 29571 se
rect 9060 29537 9100 29571
tri 9100 29537 9134 29571 nw
rect 8120 29534 8880 29537
tri 8880 29534 8883 29537 nw
tri 9023 29534 9026 29537 se
rect 9026 29534 9097 29537
tri 9097 29534 9100 29537 nw
rect 8120 29527 8873 29534
tri 8873 29527 8880 29534 nw
tri 9016 29527 9023 29534 se
rect 9023 29527 9090 29534
tri 9090 29527 9097 29534 nw
rect 8120 29517 8863 29527
tri 8863 29517 8873 29527 nw
tri 9014 29525 9016 29527 se
rect 9016 29525 9088 29527
tri 9088 29525 9090 29527 nw
tri 9006 29517 9014 29525 se
rect 9014 29517 9080 29525
tri 9080 29517 9088 29525 nw
rect 8120 29505 8851 29517
tri 8851 29505 8863 29517 nw
tri 8994 29505 9006 29517 se
rect 9006 29505 9063 29517
rect 2086 29500 2141 29505
tri 2141 29500 2146 29505 nw
tri 8989 29500 8994 29505 se
rect 8994 29500 9063 29505
tri 9063 29500 9080 29517 nw
rect 2086 29498 2139 29500
tri 2139 29498 2141 29500 nw
tri 8987 29498 8989 29500 se
rect 8989 29498 9061 29500
tri 9061 29498 9063 29500 nw
rect 2086 29471 2109 29498
rect 2034 29468 2109 29471
tri 2109 29468 2139 29498 nw
tri 8957 29468 8987 29498 se
rect 8987 29468 9031 29498
tri 9031 29468 9061 29498 nw
rect 2034 29465 2106 29468
tri 2106 29465 2109 29468 nw
tri 2147 29465 2150 29468 se
rect 2150 29465 7564 29468
tri 2146 29464 2147 29465 se
rect 2147 29464 7564 29465
tri 2143 29461 2146 29464 se
rect 2146 29461 7564 29464
tri 2136 29454 2143 29461 se
rect 2143 29454 7564 29461
tri 2127 29445 2136 29454 se
rect 2136 29445 7564 29454
tri 2110 29428 2127 29445 se
rect 2127 29428 7564 29445
tri 2108 29426 2110 29428 se
rect 2110 29426 7564 29428
tri 2107 29425 2108 29426 se
rect 2108 29425 7564 29426
tri 2098 29416 2107 29425 se
rect 2107 29416 7564 29425
rect 7616 29416 7628 29468
rect 7680 29416 7686 29468
rect 7998 29416 8004 29468
rect 8056 29416 8068 29468
rect 8120 29464 9027 29468
tri 9027 29464 9031 29468 nw
rect 8120 29461 9024 29464
tri 9024 29461 9027 29464 nw
rect 8120 29454 9017 29461
tri 9017 29454 9024 29461 nw
rect 8120 29445 9008 29454
tri 9008 29445 9017 29454 nw
rect 8120 29428 8991 29445
tri 8991 29428 9008 29445 nw
rect 8120 29425 8988 29428
tri 8988 29425 8991 29428 nw
rect 8120 29416 8979 29425
tri 8979 29416 8988 29425 nw
rect 2098 29410 2200 29416
rect 1680 29392 1736 29398
rect 1732 29391 1736 29392
tri 1736 29391 1743 29398 sw
rect 1732 29388 1743 29391
tri 1743 29388 1746 29391 sw
rect 1732 29381 1746 29388
tri 1746 29381 1753 29388 sw
rect 1732 29373 1753 29381
tri 1753 29373 1761 29381 sw
rect 1732 29371 1761 29373
tri 1761 29371 1763 29373 sw
rect 1732 29356 1763 29371
tri 1763 29356 1778 29371 sw
rect 2150 29391 2200 29410
tri 2200 29391 2225 29416 nw
rect 9901 29391 10230 30228
tri 10230 30227 10231 30228 nw
tri 13638 30227 13639 30228 ne
rect 13639 30227 13705 30228
tri 13639 30194 13672 30227 ne
rect 13672 30194 13705 30227
rect 13739 30226 13909 30228
rect 13739 30194 13807 30226
tri 13672 30192 13674 30194 ne
rect 13674 30192 13807 30194
rect 13841 30194 13909 30226
rect 13943 30194 13950 30228
rect 13841 30192 13950 30194
tri 13674 30181 13685 30192 ne
rect 13685 30181 13950 30192
tri 13685 30168 13698 30181 ne
rect 13698 30155 13950 30181
rect 13698 30121 13705 30155
rect 13739 30152 13909 30155
rect 13739 30121 13807 30152
rect 13698 30118 13807 30121
rect 13841 30121 13909 30152
rect 13943 30121 13950 30155
rect 13841 30118 13950 30121
rect 13698 30082 13950 30118
rect 13698 30048 13705 30082
rect 13739 30079 13909 30082
rect 13739 30048 13807 30079
rect 13698 30045 13807 30048
rect 13841 30048 13909 30079
rect 13943 30048 13950 30082
rect 13841 30045 13950 30048
rect 13698 30009 13950 30045
rect 13698 29975 13705 30009
rect 13739 30006 13909 30009
rect 13739 29975 13807 30006
rect 13698 29972 13807 29975
rect 13841 29975 13909 30006
rect 13943 29975 13950 30009
rect 13841 29972 13950 29975
rect 13698 29936 13950 29972
rect 13698 29902 13705 29936
rect 13739 29933 13909 29936
rect 13739 29902 13807 29933
rect 13698 29899 13807 29902
rect 13841 29902 13909 29933
rect 13943 29902 13950 29936
rect 13841 29899 13950 29902
rect 13698 29863 13950 29899
rect 13698 29829 13705 29863
rect 13739 29860 13909 29863
rect 13739 29829 13807 29860
rect 13698 29826 13807 29829
rect 13841 29829 13909 29860
rect 13943 29829 13950 29863
rect 13841 29826 13950 29829
rect 13698 29790 13950 29826
rect 13698 29756 13705 29790
rect 13739 29787 13909 29790
rect 13739 29756 13807 29787
rect 13698 29753 13807 29756
rect 13841 29756 13909 29787
rect 13943 29756 13950 29790
rect 13841 29753 13950 29756
rect 13698 29717 13950 29753
rect 13698 29683 13705 29717
rect 13739 29714 13909 29717
rect 13739 29683 13807 29714
rect 13698 29680 13807 29683
rect 13841 29683 13909 29714
rect 13943 29683 13950 29717
rect 13841 29680 13950 29683
rect 13698 29644 13950 29680
rect 13698 29610 13705 29644
rect 13739 29641 13909 29644
rect 13739 29610 13807 29641
rect 13698 29607 13807 29610
rect 13841 29610 13909 29641
rect 13943 29610 13950 29644
rect 13841 29607 13950 29610
rect 13698 29572 13950 29607
rect 13698 29571 13909 29572
rect 13698 29537 13705 29571
rect 13739 29568 13909 29571
rect 13739 29537 13807 29568
rect 13698 29534 13807 29537
rect 13841 29538 13909 29568
rect 13943 29538 13950 29572
rect 13841 29534 13950 29538
rect 13698 29500 13950 29534
rect 13698 29498 13909 29500
rect 13698 29464 13705 29498
rect 13739 29495 13909 29498
rect 13739 29464 13807 29495
rect 13698 29461 13807 29464
rect 13841 29466 13909 29495
rect 13943 29466 13950 29500
rect 13841 29461 13950 29466
rect 13698 29428 13950 29461
rect 13698 29425 13909 29428
tri 10230 29391 10231 29392 sw
rect 13698 29391 13705 29425
rect 13739 29422 13909 29425
rect 13739 29391 13807 29422
rect 2150 29388 2197 29391
tri 2197 29388 2200 29391 nw
rect 9901 29388 10231 29391
tri 10231 29388 10234 29391 sw
rect 13698 29388 13807 29391
rect 13841 29394 13909 29422
rect 13943 29394 13950 29428
rect 13841 29388 13950 29394
rect 2150 29381 2190 29388
tri 2190 29381 2197 29388 nw
rect 9901 29381 10234 29388
tri 10234 29381 10241 29388 sw
rect 2150 29373 2182 29381
tri 2182 29373 2190 29381 nw
rect 9901 29373 10241 29381
tri 10241 29373 10249 29381 sw
rect 2150 29358 2165 29373
rect 2098 29356 2165 29358
tri 2165 29356 2182 29373 nw
rect 9901 29356 10249 29373
tri 10249 29356 10266 29373 sw
rect 13698 29356 13950 29388
rect 1732 29352 1778 29356
tri 1778 29352 1782 29356 sw
rect 2098 29352 2161 29356
tri 2161 29352 2165 29356 nw
rect 9901 29352 10266 29356
tri 10266 29352 10270 29356 sw
rect 13698 29352 13909 29356
rect 1732 29342 1782 29352
tri 1782 29342 1792 29352 sw
rect 1732 29340 1792 29342
rect 1680 29337 1792 29340
rect 1680 29333 1734 29337
tri 1680 29326 1687 29333 ne
rect 1687 29326 1734 29333
tri 1687 29318 1695 29326 ne
rect 1695 29318 1734 29326
tri 1695 29315 1698 29318 ne
rect 1698 29315 1734 29318
tri 1698 29308 1705 29315 ne
rect 1705 29308 1734 29315
tri 1705 29301 1712 29308 ne
rect 1712 29301 1734 29308
tri 1712 29285 1728 29301 ne
rect 1728 29285 1734 29301
rect 1786 29285 1792 29337
rect 2098 29346 2150 29352
tri 2150 29341 2161 29352 nw
rect 2098 29288 2150 29294
rect 9901 29318 10270 29352
tri 10270 29318 10304 29352 sw
rect 13698 29318 13705 29352
rect 13739 29349 13909 29352
rect 13739 29318 13807 29349
rect 9901 29315 10304 29318
tri 10304 29315 10307 29318 sw
rect 13698 29315 13807 29318
rect 13841 29322 13909 29349
rect 13943 29322 13950 29356
rect 13841 29315 13950 29322
rect 9901 29308 10307 29315
tri 10307 29308 10314 29315 sw
rect 9901 29301 10314 29308
tri 10314 29301 10321 29308 sw
rect 9901 29288 10321 29301
tri 10321 29288 10334 29301 sw
rect 9901 29285 10334 29288
tri 10334 29285 10337 29288 sw
rect 9901 29284 10337 29285
tri 10337 29284 10338 29285 sw
rect 13698 29284 13950 29315
rect 9901 29279 10338 29284
tri 10338 29279 10343 29284 sw
rect 13698 29279 13909 29284
rect 9901 29245 10343 29279
tri 10343 29245 10377 29279 sw
rect 13698 29245 13705 29279
rect 13739 29276 13909 29279
rect 13739 29245 13807 29276
rect 9901 29242 10377 29245
tri 10377 29242 10380 29245 sw
rect 13698 29242 13807 29245
rect 13841 29250 13909 29276
rect 13943 29250 13950 29284
rect 13841 29242 13950 29250
rect 9901 29235 10380 29242
tri 10380 29235 10387 29242 sw
rect 9901 29229 10387 29235
tri 10387 29229 10393 29235 sw
rect 9901 29212 10393 29229
tri 10393 29212 10410 29229 sw
rect 13698 29212 13950 29242
rect 9901 29206 10410 29212
tri 10410 29206 10416 29212 sw
rect 13698 29206 13909 29212
rect 9901 29187 10416 29206
tri 10416 29187 10435 29206 sw
rect 9901 29175 10621 29187
rect 9901 29141 10248 29175
rect 10282 29141 10331 29175
rect 10365 29141 10414 29175
rect 10448 29141 10497 29175
rect 10531 29141 10580 29175
rect 10614 29141 10621 29175
rect 9901 29102 10621 29141
rect 9901 29068 10248 29102
rect 10282 29068 10331 29102
rect 10365 29068 10414 29102
rect 10448 29068 10497 29102
rect 10531 29068 10580 29102
rect 10614 29068 10621 29102
rect 9901 29029 10621 29068
rect 9901 28995 10248 29029
rect 10282 28995 10331 29029
rect 10365 28995 10414 29029
rect 10448 28995 10497 29029
rect 10531 28995 10580 29029
rect 10614 28995 10621 29029
rect 9901 28956 10621 28995
rect 9901 28922 10248 28956
rect 10282 28922 10331 28956
rect 10365 28922 10414 28956
rect 10448 28922 10497 28956
rect 10531 28922 10580 28956
rect 10614 28922 10621 28956
rect 9901 28883 10621 28922
rect 9901 28849 10248 28883
rect 10282 28849 10331 28883
rect 10365 28849 10414 28883
rect 10448 28849 10497 28883
rect 10531 28849 10580 28883
rect 10614 28849 10621 28883
rect 9901 28810 10621 28849
rect 9901 28776 10248 28810
rect 10282 28776 10331 28810
rect 10365 28776 10414 28810
rect 10448 28776 10497 28810
rect 10531 28776 10580 28810
rect 10614 28776 10621 28810
rect 9901 28737 10621 28776
rect 9901 28703 10248 28737
rect 10282 28703 10331 28737
rect 10365 28703 10414 28737
rect 10448 28703 10497 28737
rect 10531 28703 10580 28737
rect 10614 28703 10621 28737
rect 9901 28664 10621 28703
rect 9901 28630 10248 28664
rect 10282 28630 10331 28664
rect 10365 28630 10414 28664
rect 10448 28630 10497 28664
rect 10531 28630 10580 28664
rect 10614 28630 10621 28664
rect 9901 28591 10621 28630
rect 9901 28557 10248 28591
rect 10282 28557 10331 28591
rect 10365 28557 10414 28591
rect 10448 28557 10497 28591
rect 10531 28557 10580 28591
rect 10614 28557 10621 28591
rect 9901 28518 10621 28557
rect 9901 28484 10248 28518
rect 10282 28484 10331 28518
rect 10365 28484 10414 28518
rect 10448 28484 10497 28518
rect 10531 28484 10580 28518
rect 10614 28484 10621 28518
rect 9901 28445 10621 28484
rect 9901 28411 10248 28445
rect 10282 28411 10331 28445
rect 10365 28411 10414 28445
rect 10448 28411 10497 28445
rect 10531 28411 10580 28445
rect 10614 28411 10621 28445
rect 9901 28372 10621 28411
rect 9901 28338 10248 28372
rect 10282 28338 10331 28372
rect 10365 28338 10414 28372
rect 10448 28338 10497 28372
rect 10531 28338 10580 28372
rect 10614 28338 10621 28372
rect 9901 28299 10621 28338
rect 9901 28265 10248 28299
rect 10282 28265 10331 28299
rect 10365 28265 10414 28299
rect 10448 28265 10497 28299
rect 10531 28265 10580 28299
rect 10614 28265 10621 28299
rect 9901 28226 10621 28265
rect 9901 28192 10248 28226
rect 10282 28192 10331 28226
rect 10365 28192 10414 28226
rect 10448 28192 10497 28226
rect 10531 28192 10580 28226
rect 10614 28192 10621 28226
rect 9901 28153 10621 28192
rect 9901 28119 10248 28153
rect 10282 28119 10331 28153
rect 10365 28119 10414 28153
rect 10448 28119 10497 28153
rect 10531 28119 10580 28153
rect 10614 28119 10621 28153
rect 9901 28080 10621 28119
rect 9901 28046 10248 28080
rect 10282 28046 10331 28080
rect 10365 28046 10414 28080
rect 10448 28046 10497 28080
rect 10531 28046 10580 28080
rect 10614 28046 10621 28080
rect 9901 28007 10621 28046
rect 9901 27973 10248 28007
rect 10282 27973 10331 28007
rect 10365 27973 10414 28007
rect 10448 27973 10497 28007
rect 10531 27973 10580 28007
rect 10614 27973 10621 28007
rect 9901 27934 10621 27973
rect 9901 27900 10248 27934
rect 10282 27900 10331 27934
rect 10365 27900 10414 27934
rect 10448 27900 10497 27934
rect 10531 27900 10580 27934
rect 10614 27900 10621 27934
rect 9901 27861 10621 27900
rect 9901 27827 10248 27861
rect 10282 27827 10331 27861
rect 10365 27827 10414 27861
rect 10448 27827 10497 27861
rect 10531 27827 10580 27861
rect 10614 27827 10621 27861
rect 9901 27788 10621 27827
rect 9901 27754 10248 27788
rect 10282 27754 10331 27788
rect 10365 27754 10414 27788
rect 10448 27754 10497 27788
rect 10531 27754 10580 27788
rect 10614 27754 10621 27788
rect 9901 27715 10621 27754
rect 9901 27681 10248 27715
rect 10282 27681 10331 27715
rect 10365 27681 10414 27715
rect 10448 27681 10497 27715
rect 10531 27681 10580 27715
rect 10614 27681 10621 27715
rect 9901 27642 10621 27681
rect 9901 27608 10248 27642
rect 10282 27608 10331 27642
rect 10365 27608 10414 27642
rect 10448 27608 10497 27642
rect 10531 27608 10580 27642
rect 10614 27608 10621 27642
rect 9901 27568 10621 27608
rect 9901 27534 10248 27568
rect 10282 27534 10331 27568
rect 10365 27534 10414 27568
rect 10448 27534 10497 27568
rect 10531 27534 10580 27568
rect 10614 27534 10621 27568
rect 9901 27494 10621 27534
rect 9901 27460 10248 27494
rect 10282 27460 10331 27494
rect 10365 27460 10414 27494
rect 10448 27460 10497 27494
rect 10531 27460 10580 27494
rect 10614 27460 10621 27494
rect 9901 27420 10621 27460
rect 9901 27386 10248 27420
rect 10282 27386 10331 27420
rect 10365 27386 10414 27420
rect 10448 27386 10497 27420
rect 10531 27386 10580 27420
rect 10614 27386 10621 27420
rect 9901 27346 10621 27386
rect 9901 27312 10248 27346
rect 10282 27312 10331 27346
rect 10365 27312 10414 27346
rect 10448 27312 10497 27346
rect 10531 27312 10580 27346
rect 10614 27312 10621 27346
rect 9901 27272 10621 27312
rect 9901 27238 10248 27272
rect 10282 27238 10331 27272
rect 10365 27238 10414 27272
rect 10448 27238 10497 27272
rect 10531 27238 10580 27272
rect 10614 27238 10621 27272
rect 9901 27198 10621 27238
rect 13698 29172 13705 29206
rect 13739 29203 13909 29206
rect 13739 29172 13807 29203
rect 13698 29169 13807 29172
rect 13841 29178 13909 29203
rect 13943 29178 13950 29212
rect 13841 29169 13950 29178
rect 13698 29140 13950 29169
rect 13698 29133 13909 29140
rect 13698 29099 13705 29133
rect 13739 29130 13909 29133
rect 13739 29099 13807 29130
rect 13698 29096 13807 29099
rect 13841 29106 13909 29130
rect 13943 29106 13950 29140
rect 13841 29096 13950 29106
rect 13698 29068 13950 29096
rect 13698 29060 13909 29068
rect 13698 29026 13705 29060
rect 13739 29057 13909 29060
rect 13739 29026 13807 29057
rect 13698 29023 13807 29026
rect 13841 29034 13909 29057
rect 13943 29034 13950 29068
rect 13841 29023 13950 29034
rect 13698 28996 13950 29023
rect 13698 28987 13909 28996
rect 13698 28953 13705 28987
rect 13739 28984 13909 28987
rect 13739 28953 13807 28984
rect 13698 28950 13807 28953
rect 13841 28962 13909 28984
rect 13943 28962 13950 28996
rect 13841 28950 13950 28962
rect 13698 28924 13950 28950
rect 13698 28914 13909 28924
rect 13698 28880 13705 28914
rect 13739 28911 13909 28914
rect 13739 28880 13807 28911
rect 13698 28877 13807 28880
rect 13841 28890 13909 28911
rect 13943 28890 13950 28924
rect 13841 28877 13950 28890
rect 13698 28852 13950 28877
rect 13698 28841 13909 28852
rect 13698 28807 13705 28841
rect 13739 28838 13909 28841
rect 13739 28807 13807 28838
rect 13698 28804 13807 28807
rect 13841 28818 13909 28838
rect 13943 28818 13950 28852
rect 13841 28804 13950 28818
rect 13698 28780 13950 28804
rect 13698 28769 13909 28780
rect 13698 28735 13705 28769
rect 13739 28765 13909 28769
rect 13739 28735 13807 28765
rect 13698 28731 13807 28735
rect 13841 28746 13909 28765
rect 13943 28746 13950 28780
rect 13841 28731 13950 28746
rect 13698 28708 13950 28731
rect 13698 28697 13909 28708
rect 13698 28663 13705 28697
rect 13739 28692 13909 28697
rect 13739 28663 13807 28692
rect 13698 28658 13807 28663
rect 13841 28674 13909 28692
rect 13943 28674 13950 28708
rect 13841 28658 13950 28674
rect 13698 28636 13950 28658
rect 13698 28625 13909 28636
rect 13698 28591 13705 28625
rect 13739 28619 13909 28625
rect 13739 28591 13807 28619
rect 13698 28585 13807 28591
rect 13841 28602 13909 28619
rect 13943 28602 13950 28636
rect 13841 28585 13950 28602
rect 13698 28564 13950 28585
rect 13698 28553 13909 28564
rect 13698 28519 13705 28553
rect 13739 28546 13909 28553
rect 13739 28519 13807 28546
rect 13698 28512 13807 28519
rect 13841 28530 13909 28546
rect 13943 28530 13950 28564
rect 13841 28512 13950 28530
rect 13698 28492 13950 28512
rect 13698 28481 13909 28492
rect 13698 28447 13705 28481
rect 13739 28473 13909 28481
rect 13739 28447 13807 28473
rect 13698 28439 13807 28447
rect 13841 28458 13909 28473
rect 13943 28458 13950 28492
rect 13841 28439 13950 28458
rect 13698 28420 13950 28439
rect 13698 28409 13909 28420
rect 13698 28375 13705 28409
rect 13739 28400 13909 28409
rect 13739 28375 13807 28400
rect 13698 28366 13807 28375
rect 13841 28386 13909 28400
rect 13943 28386 13950 28420
rect 13841 28366 13950 28386
rect 13698 28348 13950 28366
rect 13698 28337 13909 28348
rect 13698 28303 13705 28337
rect 13739 28327 13909 28337
rect 13739 28303 13807 28327
rect 13698 28293 13807 28303
rect 13841 28314 13909 28327
rect 13943 28314 13950 28348
rect 13841 28293 13950 28314
rect 13698 28276 13950 28293
rect 13698 28265 13909 28276
rect 13698 28231 13705 28265
rect 13739 28254 13909 28265
rect 13739 28231 13807 28254
rect 13698 28220 13807 28231
rect 13841 28242 13909 28254
rect 13943 28242 13950 28276
rect 13841 28220 13950 28242
rect 13698 28204 13950 28220
rect 13698 28193 13909 28204
rect 13698 28159 13705 28193
rect 13739 28181 13909 28193
rect 13739 28159 13807 28181
rect 13698 28147 13807 28159
rect 13841 28170 13909 28181
rect 13943 28170 13950 28204
rect 13841 28147 13950 28170
rect 13698 28132 13950 28147
rect 13698 28121 13909 28132
rect 13698 28087 13705 28121
rect 13739 28108 13909 28121
rect 13739 28087 13807 28108
rect 13698 28074 13807 28087
rect 13841 28098 13909 28108
rect 13943 28098 13950 28132
rect 13841 28074 13950 28098
rect 13698 28060 13950 28074
rect 13698 28049 13909 28060
rect 13698 28015 13705 28049
rect 13739 28035 13909 28049
rect 13739 28015 13807 28035
rect 13698 28001 13807 28015
rect 13841 28026 13909 28035
rect 13943 28026 13950 28060
rect 13841 28001 13950 28026
rect 13698 27988 13950 28001
rect 13698 27977 13909 27988
rect 13698 27943 13705 27977
rect 13739 27962 13909 27977
rect 13739 27943 13807 27962
rect 13698 27928 13807 27943
rect 13841 27954 13909 27962
rect 13943 27954 13950 27988
rect 13841 27928 13950 27954
rect 13698 27916 13950 27928
rect 13698 27905 13909 27916
rect 13698 27871 13705 27905
rect 13739 27889 13909 27905
rect 13739 27871 13807 27889
rect 13698 27855 13807 27871
rect 13841 27882 13909 27889
rect 13943 27882 13950 27916
rect 13841 27855 13950 27882
rect 13698 27844 13950 27855
rect 13698 27833 13909 27844
rect 13698 27799 13705 27833
rect 13739 27816 13909 27833
rect 13739 27799 13807 27816
rect 13698 27782 13807 27799
rect 13841 27810 13909 27816
rect 13943 27810 13950 27844
rect 13841 27782 13950 27810
rect 13698 27772 13950 27782
rect 13698 27761 13909 27772
rect 13698 27727 13705 27761
rect 13739 27743 13909 27761
rect 13739 27727 13807 27743
rect 13698 27709 13807 27727
rect 13841 27738 13909 27743
rect 13943 27738 13950 27772
rect 13841 27709 13950 27738
rect 13698 27700 13950 27709
rect 13698 27689 13909 27700
rect 13698 27655 13705 27689
rect 13739 27670 13909 27689
rect 13739 27655 13807 27670
rect 13698 27636 13807 27655
rect 13841 27666 13909 27670
rect 13943 27666 13950 27700
rect 13841 27636 13950 27666
rect 13698 27628 13950 27636
rect 13698 27617 13909 27628
rect 13698 27583 13705 27617
rect 13739 27597 13909 27617
rect 13739 27583 13807 27597
rect 13698 27563 13807 27583
rect 13841 27594 13909 27597
rect 13943 27594 13950 27628
rect 13841 27563 13950 27594
rect 13698 27556 13950 27563
rect 13698 27545 13909 27556
rect 13698 27511 13705 27545
rect 13739 27524 13909 27545
rect 13739 27511 13807 27524
rect 13698 27490 13807 27511
rect 13841 27522 13909 27524
rect 13943 27522 13950 27556
rect 13841 27490 13950 27522
rect 13698 27484 13950 27490
rect 13698 27473 13909 27484
rect 13698 27439 13705 27473
rect 13739 27451 13909 27473
rect 13739 27439 13807 27451
rect 13698 27417 13807 27439
rect 13841 27450 13909 27451
rect 13943 27450 13950 27484
rect 13841 27417 13950 27450
rect 13698 27412 13950 27417
rect 13698 27401 13909 27412
rect 13698 27367 13705 27401
rect 13739 27378 13909 27401
rect 13943 27378 13950 27412
rect 13739 27367 13807 27378
rect 13698 27344 13807 27367
rect 13841 27344 13950 27378
rect 13698 27340 13950 27344
rect 13698 27329 13909 27340
rect 13698 27295 13705 27329
rect 13739 27306 13909 27329
rect 13943 27306 13950 27340
rect 13739 27305 13950 27306
rect 13739 27295 13807 27305
rect 13698 27271 13807 27295
rect 13841 27271 13950 27305
rect 13698 27268 13950 27271
rect 13698 27257 13909 27268
rect 13698 27223 13705 27257
rect 13739 27234 13909 27257
rect 13943 27234 13950 27268
rect 13739 27232 13950 27234
rect 13739 27223 13807 27232
tri 13682 27198 13698 27214 se
rect 13698 27198 13807 27223
rect 13841 27198 13950 27232
rect 9901 27164 10248 27198
rect 10282 27164 10331 27198
rect 10365 27164 10414 27198
rect 10448 27164 10497 27198
rect 10531 27164 10580 27198
rect 10614 27164 10621 27198
tri 13680 27196 13682 27198 se
rect 13682 27196 13950 27198
tri 13669 27185 13680 27196 se
rect 13680 27185 13909 27196
rect 9901 27125 10621 27164
tri 13635 27151 13669 27185 se
rect 13669 27151 13705 27185
rect 13739 27162 13909 27185
rect 13943 27162 13950 27196
rect 13739 27159 13950 27162
rect 13739 27151 13807 27159
tri 13631 27147 13635 27151 se
rect 13635 27147 13807 27151
tri 10621 27125 10643 27147 sw
tri 13609 27125 13631 27147 se
rect 13631 27125 13807 27147
rect 13841 27125 13950 27159
rect 9901 27124 10643 27125
tri 10643 27124 10644 27125 sw
tri 13608 27124 13609 27125 se
rect 13609 27124 13950 27125
rect 9901 27090 10248 27124
rect 10282 27090 10331 27124
rect 10365 27090 10414 27124
rect 10448 27090 10497 27124
rect 10531 27090 10580 27124
rect 10614 27113 10644 27124
tri 10644 27113 10655 27124 sw
tri 13597 27113 13608 27124 se
rect 13608 27113 13909 27124
rect 10614 27090 10655 27113
rect 9901 27079 10655 27090
tri 10655 27079 10689 27113 sw
tri 13563 27079 13597 27113 se
rect 13597 27079 13705 27113
rect 13739 27090 13909 27113
rect 13943 27090 13950 27124
rect 13739 27086 13950 27090
rect 13739 27079 13807 27086
rect 9901 27052 10689 27079
tri 10689 27052 10716 27079 sw
tri 13536 27052 13563 27079 se
rect 13563 27052 13807 27079
rect 13841 27052 13950 27086
rect 9901 27050 10716 27052
rect 9901 27016 10248 27050
rect 10282 27016 10331 27050
rect 10365 27016 10414 27050
rect 10448 27016 10497 27050
rect 10531 27016 10580 27050
rect 10614 27041 10716 27050
tri 10716 27041 10727 27052 sw
tri 13525 27041 13536 27052 se
rect 13536 27041 13909 27052
rect 10614 27016 10727 27041
rect 9901 27007 10727 27016
tri 10727 27007 10761 27041 sw
tri 13491 27007 13525 27041 se
rect 13525 27007 13705 27041
rect 13739 27018 13909 27041
rect 13943 27018 13950 27052
rect 13739 27013 13950 27018
rect 13739 27007 13807 27013
rect 9901 26979 10761 27007
tri 10761 26979 10789 27007 sw
tri 13463 26979 13491 27007 se
rect 13491 26979 13807 27007
rect 13841 26980 13950 27013
rect 13841 26979 13909 26980
rect 9901 26976 10789 26979
tri 10789 26976 10792 26979 sw
tri 13460 26976 13463 26979 se
rect 13463 26976 13909 26979
rect 9901 26942 10248 26976
rect 10282 26942 10331 26976
rect 10365 26942 10414 26976
rect 10448 26942 10497 26976
rect 10531 26942 10580 26976
rect 10614 26973 13909 26976
rect 10614 26969 13024 26973
rect 13076 26969 13093 26973
rect 13145 26969 13162 26973
rect 13214 26969 13231 26973
rect 13283 26969 13300 26973
rect 13352 26969 13369 26973
rect 13421 26969 13439 26973
rect 13491 26969 13509 26973
rect 13561 26969 13579 26973
rect 13631 26969 13649 26973
rect 13701 26969 13909 26973
rect 10614 26942 10659 26969
rect 9901 26935 10659 26942
rect 10693 26935 10731 26969
rect 10765 26935 10803 26969
rect 10837 26935 10875 26969
rect 10909 26935 10947 26969
rect 10981 26935 11019 26969
rect 11053 26935 11091 26969
rect 11125 26935 11163 26969
rect 11197 26935 11235 26969
rect 11269 26935 11307 26969
rect 11341 26935 11379 26969
rect 11413 26935 11451 26969
rect 11485 26935 11523 26969
rect 11557 26935 11595 26969
rect 11629 26935 11667 26969
rect 11701 26935 11739 26969
rect 11773 26935 11811 26969
rect 11845 26935 11883 26969
rect 11917 26935 11955 26969
rect 11989 26935 12027 26969
rect 12061 26935 12099 26969
rect 12133 26935 12172 26969
rect 12206 26935 12245 26969
rect 12279 26935 12318 26969
rect 12352 26935 12391 26969
rect 12425 26935 12464 26969
rect 12498 26935 12537 26969
rect 12571 26935 12610 26969
rect 12644 26935 12683 26969
rect 12717 26935 12756 26969
rect 12790 26935 12829 26969
rect 12863 26935 12902 26969
rect 12936 26935 12975 26969
rect 13009 26935 13024 26969
rect 13082 26935 13093 26969
rect 13155 26935 13162 26969
rect 13228 26935 13231 26969
rect 13631 26935 13632 26969
rect 13701 26935 13705 26969
rect 13739 26946 13909 26969
rect 13943 26946 13950 26980
rect 13739 26940 13950 26946
rect 13739 26935 13807 26940
rect 9901 26921 13024 26935
rect 13076 26921 13093 26935
rect 13145 26921 13162 26935
rect 13214 26921 13231 26935
rect 13283 26921 13300 26935
rect 13352 26921 13369 26935
rect 13421 26921 13439 26935
rect 13491 26921 13509 26935
rect 13561 26921 13579 26935
rect 13631 26921 13649 26935
rect 13701 26921 13807 26935
rect 9901 26909 13807 26921
rect 9901 26902 13024 26909
rect 9901 26868 10248 26902
rect 10282 26868 10331 26902
rect 10365 26868 10414 26902
rect 10448 26868 10497 26902
rect 10531 26868 10580 26902
rect 10614 26868 13024 26902
rect 9901 26867 13024 26868
rect 13076 26867 13093 26909
rect 13145 26867 13162 26909
rect 13214 26867 13231 26909
rect 13283 26867 13300 26909
rect 13352 26867 13369 26909
rect 13421 26867 13439 26909
rect 9901 26833 10659 26867
rect 10693 26833 10732 26867
rect 10766 26833 10805 26867
rect 10839 26833 10878 26867
rect 10912 26833 10951 26867
rect 10985 26833 11024 26867
rect 11058 26833 11097 26867
rect 11131 26833 11170 26867
rect 11204 26833 11243 26867
rect 11277 26833 11316 26867
rect 11350 26833 11389 26867
rect 11423 26833 11462 26867
rect 11496 26833 11535 26867
rect 11569 26833 11608 26867
rect 11642 26833 11681 26867
rect 11715 26833 11754 26867
rect 11788 26833 11827 26867
rect 11861 26833 11900 26867
rect 11934 26833 11973 26867
rect 12007 26833 12046 26867
rect 12080 26833 12119 26867
rect 12153 26833 12192 26867
rect 12226 26833 12265 26867
rect 12299 26833 12338 26867
rect 12372 26833 12411 26867
rect 12445 26833 12484 26867
rect 12518 26833 12557 26867
rect 12591 26833 12630 26867
rect 12664 26833 12703 26867
rect 12737 26833 12776 26867
rect 12810 26833 12849 26867
rect 12883 26833 12922 26867
rect 12956 26833 12995 26867
rect 13214 26857 13215 26867
rect 13283 26857 13289 26867
rect 13352 26857 13363 26867
rect 13421 26857 13437 26867
rect 13491 26857 13509 26909
rect 13561 26857 13579 26909
rect 13631 26857 13649 26909
rect 13701 26906 13807 26909
rect 13841 26908 13950 26940
rect 13841 26906 13909 26908
rect 13701 26874 13909 26906
rect 13943 26874 13950 26908
rect 13701 26867 13950 26874
rect 13701 26857 13733 26867
rect 13029 26845 13068 26857
rect 13102 26845 13141 26857
rect 13175 26845 13215 26857
rect 13249 26845 13289 26857
rect 13323 26845 13363 26857
rect 13397 26845 13437 26857
rect 13471 26845 13511 26857
rect 13545 26845 13585 26857
rect 13619 26845 13659 26857
rect 13693 26845 13733 26857
rect 13214 26833 13215 26845
rect 13283 26833 13289 26845
rect 13352 26833 13363 26845
rect 13421 26833 13437 26845
rect 9901 26828 13024 26833
rect 9901 26794 10248 26828
rect 10282 26794 10331 26828
rect 10365 26794 10414 26828
rect 10448 26794 10497 26828
rect 10531 26794 10580 26828
rect 10614 26794 13024 26828
rect 9901 26793 13024 26794
rect 13076 26793 13093 26833
rect 13145 26793 13162 26833
rect 13214 26793 13231 26833
rect 13283 26793 13300 26833
rect 13352 26793 13369 26833
rect 13421 26793 13439 26833
rect 13491 26793 13509 26845
rect 13561 26793 13579 26845
rect 13631 26793 13649 26845
rect 13701 26833 13733 26845
rect 13767 26833 13807 26867
rect 13841 26836 13950 26867
rect 13841 26833 13909 26836
rect 13701 26802 13909 26833
rect 13943 26802 13950 26836
rect 13701 26793 13950 26802
rect 9901 26781 13950 26793
rect 9901 26765 13024 26781
rect 9901 26754 10659 26765
rect 9901 26720 10248 26754
rect 10282 26720 10331 26754
rect 10365 26720 10414 26754
rect 10448 26720 10497 26754
rect 10531 26720 10580 26754
rect 10614 26731 10659 26754
rect 10693 26731 10731 26765
rect 10765 26731 10803 26765
rect 10837 26731 10875 26765
rect 10909 26731 10947 26765
rect 10981 26731 11019 26765
rect 11053 26731 11091 26765
rect 11125 26731 11163 26765
rect 11197 26731 11235 26765
rect 11269 26731 11307 26765
rect 11341 26731 11379 26765
rect 11413 26731 11451 26765
rect 11485 26731 11523 26765
rect 11557 26731 11595 26765
rect 11629 26731 11667 26765
rect 11701 26731 11739 26765
rect 11773 26731 11811 26765
rect 11845 26731 11883 26765
rect 11917 26731 11955 26765
rect 11989 26731 12027 26765
rect 12061 26731 12099 26765
rect 12133 26731 12171 26765
rect 12205 26731 12243 26765
rect 12277 26731 12315 26765
rect 12349 26731 12387 26765
rect 12421 26731 12459 26765
rect 12493 26731 12531 26765
rect 12565 26731 12603 26765
rect 12637 26731 12675 26765
rect 12709 26731 12747 26765
rect 12781 26731 12819 26765
rect 12853 26731 12891 26765
rect 12925 26731 12963 26765
rect 12997 26731 13024 26765
rect 10614 26729 13024 26731
rect 13076 26729 13093 26781
rect 13145 26729 13162 26781
rect 13214 26765 13231 26781
rect 13283 26765 13300 26781
rect 13352 26765 13369 26781
rect 13421 26765 13439 26781
rect 13491 26765 13509 26781
rect 13561 26765 13579 26781
rect 13631 26765 13649 26781
rect 13701 26765 13950 26781
rect 13215 26731 13231 26765
rect 13288 26731 13300 26765
rect 13361 26731 13369 26765
rect 13434 26731 13439 26765
rect 13507 26731 13509 26765
rect 13726 26731 13765 26765
rect 13799 26731 13838 26765
rect 13872 26731 13950 26765
rect 14096 30647 14270 30669
rect 14096 30613 14102 30647
rect 14136 30631 14270 30647
rect 14136 30613 14230 30631
rect 14096 30597 14230 30613
rect 14264 30597 14270 30631
rect 14096 30575 14270 30597
rect 14096 30541 14102 30575
rect 14136 30559 14270 30575
rect 14136 30541 14230 30559
rect 14096 30525 14230 30541
rect 14264 30525 14270 30559
rect 14096 30503 14270 30525
rect 14096 30469 14102 30503
rect 14136 30487 14270 30503
rect 14136 30469 14230 30487
rect 14096 30453 14230 30469
rect 14264 30453 14270 30487
rect 14096 30431 14270 30453
rect 14096 30397 14102 30431
rect 14136 30415 14270 30431
rect 14136 30397 14230 30415
rect 14096 30381 14230 30397
rect 14264 30381 14270 30415
rect 14096 30359 14270 30381
rect 14096 30325 14102 30359
rect 14136 30343 14270 30359
rect 14136 30325 14230 30343
rect 14096 30309 14230 30325
rect 14264 30309 14270 30343
rect 14096 30287 14270 30309
rect 14096 30253 14102 30287
rect 14136 30271 14270 30287
rect 14136 30253 14230 30271
rect 14096 30237 14230 30253
rect 14264 30237 14270 30271
rect 14096 30215 14270 30237
rect 14096 30181 14102 30215
rect 14136 30199 14270 30215
rect 14136 30181 14230 30199
rect 14096 30165 14230 30181
rect 14264 30165 14270 30199
rect 14096 30143 14270 30165
rect 14096 30109 14102 30143
rect 14136 30127 14270 30143
rect 14136 30109 14230 30127
rect 14096 30093 14230 30109
rect 14264 30093 14270 30127
rect 14096 30071 14270 30093
rect 14096 30037 14102 30071
rect 14136 30055 14270 30071
rect 14136 30037 14230 30055
rect 14096 30021 14230 30037
rect 14264 30021 14270 30055
rect 14096 29999 14270 30021
rect 14096 29965 14102 29999
rect 14136 29983 14270 29999
rect 14136 29965 14230 29983
rect 14096 29949 14230 29965
rect 14264 29949 14270 29983
rect 14096 29926 14270 29949
rect 14096 29892 14102 29926
rect 14136 29911 14270 29926
rect 14136 29892 14230 29911
rect 14096 29877 14230 29892
rect 14264 29877 14270 29911
rect 14096 29853 14270 29877
rect 14096 29819 14102 29853
rect 14136 29839 14270 29853
rect 14136 29819 14230 29839
rect 14096 29805 14230 29819
rect 14264 29805 14270 29839
rect 14096 29780 14270 29805
rect 14096 29746 14102 29780
rect 14136 29767 14270 29780
rect 14136 29746 14230 29767
rect 14096 29733 14230 29746
rect 14264 29733 14270 29767
rect 14096 29707 14270 29733
rect 14096 29673 14102 29707
rect 14136 29695 14270 29707
rect 14136 29673 14230 29695
rect 14096 29661 14230 29673
rect 14264 29661 14270 29695
rect 14096 29634 14270 29661
rect 14096 29600 14102 29634
rect 14136 29623 14270 29634
rect 14136 29600 14230 29623
rect 14096 29589 14230 29600
rect 14264 29589 14270 29623
rect 14096 29561 14270 29589
rect 14096 29527 14102 29561
rect 14136 29551 14270 29561
rect 14136 29527 14230 29551
rect 14096 29517 14230 29527
rect 14264 29517 14270 29551
rect 14096 29488 14270 29517
rect 14096 29454 14102 29488
rect 14136 29479 14270 29488
rect 14136 29454 14230 29479
rect 14096 29445 14230 29454
rect 14264 29445 14270 29479
rect 14096 29415 14270 29445
rect 14096 29381 14102 29415
rect 14136 29407 14270 29415
rect 14136 29381 14230 29407
rect 14096 29373 14230 29381
rect 14264 29373 14270 29407
rect 14096 29342 14270 29373
rect 14096 29308 14102 29342
rect 14136 29335 14270 29342
rect 14136 29308 14230 29335
rect 14096 29301 14230 29308
rect 14264 29301 14270 29335
rect 14096 29269 14270 29301
rect 14096 29235 14102 29269
rect 14136 29263 14270 29269
rect 14136 29235 14230 29263
rect 14096 29229 14230 29235
rect 14264 29229 14270 29263
rect 14096 29196 14270 29229
rect 14096 29162 14102 29196
rect 14136 29191 14270 29196
rect 14136 29162 14230 29191
rect 14096 29157 14230 29162
rect 14264 29157 14270 29191
rect 14096 29123 14270 29157
rect 14096 29089 14102 29123
rect 14136 29119 14270 29123
rect 14136 29089 14230 29119
rect 14096 29085 14230 29089
rect 14264 29085 14270 29119
rect 14096 29050 14270 29085
rect 14096 29016 14102 29050
rect 14136 29047 14270 29050
rect 14136 29016 14230 29047
rect 14096 29013 14230 29016
rect 14264 29013 14270 29047
rect 14096 28977 14270 29013
rect 14096 28943 14102 28977
rect 14136 28975 14270 28977
rect 14136 28943 14230 28975
rect 14096 28941 14230 28943
rect 14264 28941 14270 28975
rect 14096 28904 14270 28941
rect 14096 28870 14102 28904
rect 14136 28903 14270 28904
rect 14136 28870 14230 28903
rect 14096 28869 14230 28870
rect 14264 28869 14270 28903
rect 14096 28831 14270 28869
rect 14096 28797 14102 28831
rect 14136 28797 14230 28831
rect 14264 28797 14270 28831
rect 14096 28759 14270 28797
rect 14096 28758 14230 28759
rect 14096 28724 14102 28758
rect 14136 28725 14230 28758
rect 14264 28725 14270 28759
rect 14136 28724 14270 28725
rect 14096 28687 14270 28724
rect 14096 28685 14230 28687
rect 14096 28651 14102 28685
rect 14136 28653 14230 28685
rect 14264 28653 14270 28687
rect 14136 28651 14270 28653
rect 14096 28615 14270 28651
rect 14096 28612 14230 28615
rect 14096 28578 14102 28612
rect 14136 28581 14230 28612
rect 14264 28581 14270 28615
rect 14136 28578 14270 28581
rect 14096 28543 14270 28578
rect 14096 28539 14230 28543
rect 14096 28505 14102 28539
rect 14136 28509 14230 28539
rect 14264 28509 14270 28543
rect 14136 28505 14270 28509
rect 14096 28471 14270 28505
rect 14096 28466 14230 28471
rect 14096 28432 14102 28466
rect 14136 28437 14230 28466
rect 14264 28437 14270 28471
rect 14136 28432 14270 28437
rect 14096 28399 14270 28432
rect 14096 28393 14230 28399
rect 14096 28359 14102 28393
rect 14136 28365 14230 28393
rect 14264 28365 14270 28399
rect 14136 28359 14270 28365
rect 14096 28327 14270 28359
rect 14096 28320 14230 28327
rect 14096 28286 14102 28320
rect 14136 28293 14230 28320
rect 14264 28293 14270 28327
rect 14136 28286 14270 28293
rect 14096 28255 14270 28286
rect 14096 28247 14230 28255
rect 14096 28213 14102 28247
rect 14136 28221 14230 28247
rect 14264 28221 14270 28255
rect 14136 28213 14270 28221
rect 14096 28183 14270 28213
rect 14096 28174 14230 28183
rect 14096 28140 14102 28174
rect 14136 28149 14230 28174
rect 14264 28149 14270 28183
rect 14136 28140 14270 28149
rect 14096 28111 14270 28140
rect 14096 28101 14230 28111
rect 14096 28067 14102 28101
rect 14136 28077 14230 28101
rect 14264 28077 14270 28111
rect 14136 28067 14270 28077
rect 14096 28039 14270 28067
rect 14096 28028 14230 28039
rect 14096 27994 14102 28028
rect 14136 28005 14230 28028
rect 14264 28005 14270 28039
rect 14136 27994 14270 28005
rect 14096 27967 14270 27994
rect 14096 27955 14230 27967
rect 14096 27921 14102 27955
rect 14136 27933 14230 27955
rect 14264 27933 14270 27967
rect 14136 27921 14270 27933
rect 14096 27895 14270 27921
rect 14096 27882 14230 27895
rect 14096 27848 14102 27882
rect 14136 27861 14230 27882
rect 14264 27861 14270 27895
rect 14136 27848 14270 27861
rect 14096 27823 14270 27848
rect 14096 27809 14230 27823
rect 14096 27775 14102 27809
rect 14136 27789 14230 27809
rect 14264 27789 14270 27823
rect 14136 27775 14270 27789
rect 14096 27751 14270 27775
rect 14096 27736 14230 27751
rect 14096 27702 14102 27736
rect 14136 27717 14230 27736
rect 14264 27717 14270 27751
rect 14136 27702 14270 27717
rect 14096 27679 14270 27702
rect 14096 27663 14230 27679
rect 14096 27629 14102 27663
rect 14136 27645 14230 27663
rect 14264 27645 14270 27679
rect 14136 27629 14270 27645
rect 14096 27607 14270 27629
rect 14096 27590 14230 27607
rect 14096 27556 14102 27590
rect 14136 27573 14230 27590
rect 14264 27573 14270 27607
rect 14136 27556 14270 27573
rect 14096 27534 14270 27556
rect 14096 27517 14230 27534
rect 14096 27483 14102 27517
rect 14136 27500 14230 27517
rect 14264 27500 14270 27534
rect 14136 27483 14270 27500
rect 14096 27461 14270 27483
rect 14096 27444 14230 27461
rect 14096 27410 14102 27444
rect 14136 27427 14230 27444
rect 14264 27427 14270 27461
rect 14136 27410 14270 27427
rect 14096 27388 14270 27410
rect 14096 27371 14230 27388
rect 14096 27337 14102 27371
rect 14136 27354 14230 27371
rect 14264 27354 14270 27388
rect 14136 27337 14270 27354
rect 14096 27315 14270 27337
rect 14096 27298 14230 27315
rect 14096 27264 14102 27298
rect 14136 27281 14230 27298
rect 14264 27281 14270 27315
rect 14136 27264 14270 27281
rect 14096 27242 14270 27264
rect 14096 27225 14230 27242
rect 14096 27191 14102 27225
rect 14136 27208 14230 27225
rect 14264 27208 14270 27242
rect 14136 27191 14270 27208
rect 14096 27169 14270 27191
rect 14096 27152 14230 27169
rect 14096 27118 14102 27152
rect 14136 27135 14230 27152
rect 14264 27135 14270 27169
rect 14136 27118 14270 27135
rect 14096 27096 14270 27118
rect 14096 27079 14230 27096
rect 14096 27045 14102 27079
rect 14136 27062 14230 27079
rect 14264 27062 14270 27096
rect 14136 27045 14270 27062
rect 14096 27023 14270 27045
rect 14096 27006 14230 27023
rect 14096 26972 14102 27006
rect 14136 26989 14230 27006
rect 14264 26989 14270 27023
rect 14136 26972 14270 26989
rect 14096 26950 14270 26972
rect 14096 26933 14230 26950
rect 14096 26899 14102 26933
rect 14136 26916 14230 26933
rect 14264 26916 14270 26950
rect 14818 27556 15258 27562
rect 14818 26992 14820 27556
rect 15256 26992 15258 27556
rect 14818 26979 15258 26992
rect 14818 26927 14820 26979
rect 14872 26927 14884 26979
rect 14936 26927 14948 26979
rect 15000 26927 15012 26979
rect 15064 26927 15076 26979
rect 15128 26927 15140 26979
rect 15192 26927 15204 26979
rect 15256 26927 15258 26979
rect 14818 26921 15258 26927
rect 14136 26899 14270 26916
rect 14096 26877 14270 26899
rect 14096 26860 14230 26877
rect 14096 26826 14102 26860
rect 14136 26843 14230 26860
rect 14264 26843 14270 26877
rect 14136 26826 14270 26843
rect 14096 26804 14270 26826
rect 14096 26787 14230 26804
rect 14096 26753 14102 26787
rect 14136 26770 14230 26787
rect 14264 26770 14270 26804
rect 14136 26753 14270 26770
tri 14090 26731 14096 26737 se
rect 14096 26731 14270 26753
rect 13214 26729 13231 26731
rect 13283 26729 13300 26731
rect 13352 26729 13369 26731
rect 13421 26729 13439 26731
rect 13491 26729 13509 26731
rect 13561 26729 13579 26731
rect 13631 26729 13649 26731
rect 13701 26729 13950 26731
rect 10614 26724 13950 26729
tri 14083 26724 14090 26731 se
rect 14090 26724 14230 26731
rect 10614 26720 10653 26724
rect 9901 26714 10653 26720
tri 10653 26714 10663 26724 nw
tri 14073 26714 14083 26724 se
rect 14083 26714 14230 26724
rect 9901 26708 10647 26714
tri 10647 26708 10653 26714 nw
tri 14067 26708 14073 26714 se
rect 14073 26708 14102 26714
tri 14065 26706 14067 26708 se
rect 14067 26706 14102 26708
tri 9726 26680 9752 26706 sw
tri 14039 26680 14065 26706 se
rect 14065 26680 14102 26706
rect 14136 26697 14230 26714
rect 14264 26697 14270 26731
rect 14136 26680 14270 26697
rect 9726 26658 9752 26680
tri 9752 26658 9774 26680 sw
tri 14017 26658 14039 26680 se
rect 14039 26658 14270 26680
rect 9726 26641 9774 26658
tri 9774 26641 9791 26658 sw
tri 14000 26641 14017 26658 se
rect 14017 26641 14230 26658
rect 9726 26607 9791 26641
tri 9791 26607 9825 26641 sw
tri 13966 26607 14000 26641 se
rect 14000 26607 14102 26641
rect 14136 26624 14230 26641
rect 14264 26624 14270 26658
rect 14136 26607 14270 26624
rect 9726 26585 9825 26607
tri 9825 26585 9847 26607 sw
tri 13944 26585 13966 26607 se
rect 13966 26585 14270 26607
rect 9726 26574 9847 26585
tri 9847 26574 9858 26585 sw
tri 13933 26574 13944 26585 se
rect 13944 26574 14230 26585
rect 9726 26568 14230 26574
rect 9726 26534 9765 26568
rect 9799 26534 9838 26568
rect 9872 26534 9911 26568
rect 9945 26534 9984 26568
rect 10018 26534 10057 26568
rect 10091 26534 10130 26568
rect 10164 26534 10203 26568
rect 10237 26534 10276 26568
rect 10310 26534 10349 26568
rect 10383 26534 10422 26568
rect 10456 26534 10495 26568
rect 10529 26534 10568 26568
rect 10602 26534 10641 26568
rect 10675 26534 10714 26568
rect 10748 26534 10787 26568
rect 10821 26534 10860 26568
rect 10894 26534 10933 26568
rect 10967 26534 11006 26568
rect 11040 26534 11078 26568
rect 11112 26534 11150 26568
rect 11184 26534 11222 26568
rect 11256 26534 11294 26568
rect 11328 26534 11366 26568
rect 11400 26534 11438 26568
rect 11472 26534 11510 26568
rect 11544 26534 11582 26568
rect 11616 26534 11654 26568
rect 11688 26534 11726 26568
rect 11760 26534 11798 26568
rect 11832 26534 11870 26568
rect 11904 26534 11942 26568
rect 11976 26534 12014 26568
rect 12048 26534 12086 26568
rect 12120 26534 12158 26568
rect 12192 26534 12230 26568
rect 12264 26534 12302 26568
rect 12336 26534 12374 26568
rect 12408 26534 12446 26568
rect 12480 26534 12518 26568
rect 12552 26534 12590 26568
rect 12624 26534 12662 26568
rect 12696 26534 12734 26568
rect 12768 26534 12806 26568
rect 12840 26534 12878 26568
rect 12912 26534 12950 26568
rect 12984 26534 13022 26568
rect 13056 26534 13094 26568
rect 13128 26534 13166 26568
rect 13200 26534 13238 26568
rect 13272 26534 13310 26568
rect 13344 26534 13382 26568
rect 13416 26534 13454 26568
rect 13488 26534 13526 26568
rect 13560 26534 13598 26568
rect 13632 26534 13670 26568
rect 13704 26534 13742 26568
rect 13776 26534 13814 26568
rect 13848 26534 13886 26568
rect 13920 26534 13958 26568
rect 13992 26534 14030 26568
rect 14064 26534 14102 26568
rect 14136 26551 14230 26568
rect 14264 26551 14270 26585
rect 14136 26534 14270 26551
rect 9726 26512 14270 26534
rect 9726 26478 14230 26512
rect 14264 26478 14270 26512
rect 9726 26440 14270 26478
rect 9726 26406 9765 26440
rect 9799 26406 9838 26440
rect 9872 26406 9910 26440
rect 9944 26406 9982 26440
rect 10016 26406 10054 26440
rect 10088 26406 10126 26440
rect 10160 26406 10198 26440
rect 10232 26406 10270 26440
rect 10304 26406 10342 26440
rect 10376 26406 10414 26440
rect 10448 26406 10486 26440
rect 10520 26406 10558 26440
rect 10592 26406 10630 26440
rect 10664 26406 10702 26440
rect 10736 26406 10774 26440
rect 10808 26406 10846 26440
rect 10880 26406 10918 26440
rect 10952 26406 10990 26440
rect 11024 26406 11062 26440
rect 11096 26406 11134 26440
rect 11168 26406 11206 26440
rect 11240 26406 11278 26440
rect 11312 26406 11350 26440
rect 11384 26406 11422 26440
rect 11456 26406 11494 26440
rect 11528 26406 11566 26440
rect 11600 26406 11638 26440
rect 11672 26406 11710 26440
rect 11744 26406 11782 26440
rect 11816 26406 11854 26440
rect 11888 26406 11926 26440
rect 11960 26406 11998 26440
rect 12032 26406 12070 26440
rect 12104 26406 12142 26440
rect 12176 26406 12214 26440
rect 12248 26406 12286 26440
rect 12320 26406 12358 26440
rect 12392 26406 12430 26440
rect 12464 26406 12502 26440
rect 12536 26406 12574 26440
rect 12608 26406 12646 26440
rect 12680 26406 12718 26440
rect 12752 26406 12790 26440
rect 12824 26406 12862 26440
rect 12896 26406 12934 26440
rect 12968 26406 13006 26440
rect 13040 26406 13078 26440
rect 13112 26406 13150 26440
rect 13184 26406 13222 26440
rect 13256 26406 13294 26440
rect 13328 26406 13366 26440
rect 13400 26406 13438 26440
rect 13472 26406 13510 26440
rect 13544 26406 13582 26440
rect 13616 26406 13654 26440
rect 13688 26406 13726 26440
rect 13760 26406 13798 26440
rect 13832 26406 13870 26440
rect 13904 26406 13942 26440
rect 13976 26406 14014 26440
rect 14048 26406 14086 26440
rect 14120 26406 14158 26440
rect 14192 26406 14270 26440
rect 9726 26400 14270 26406
tri 9726 26268 9858 26400 nw
rect 9901 26253 14194 26260
rect 9901 26248 13022 26253
rect 13074 26248 13092 26253
rect 13144 26248 13162 26253
rect 13214 26248 13232 26253
rect 13284 26248 13302 26253
rect 13354 26248 13372 26253
rect 13424 26248 13442 26253
rect 13494 26248 13512 26253
rect 13564 26248 13582 26253
rect 9901 26214 9909 26248
rect 9943 26214 9981 26248
rect 10015 26214 10053 26248
rect 10087 26214 10125 26248
rect 10159 26214 10197 26248
rect 10231 26214 10269 26248
rect 10303 26214 10341 26248
rect 10375 26214 10413 26248
rect 10447 26214 10485 26248
rect 10519 26214 10557 26248
rect 10591 26214 10629 26248
rect 10663 26214 10701 26248
rect 10735 26214 10773 26248
rect 10807 26214 10845 26248
rect 10879 26214 10917 26248
rect 10951 26214 10989 26248
rect 11023 26214 11061 26248
rect 11095 26214 11133 26248
rect 11167 26214 11205 26248
rect 11239 26214 11277 26248
rect 11311 26214 11349 26248
rect 11383 26214 11421 26248
rect 11455 26214 11493 26248
rect 11527 26214 11565 26248
rect 11599 26214 11637 26248
rect 11671 26214 11709 26248
rect 11743 26214 11781 26248
rect 11815 26214 11853 26248
rect 11887 26214 11925 26248
rect 11959 26214 11997 26248
rect 12031 26214 12069 26248
rect 12103 26214 12141 26248
rect 12175 26214 12213 26248
rect 12247 26214 12285 26248
rect 12319 26214 12357 26248
rect 12391 26214 12429 26248
rect 12463 26214 12501 26248
rect 12535 26214 12573 26248
rect 12607 26214 12645 26248
rect 12679 26214 12717 26248
rect 12751 26214 12789 26248
rect 12823 26214 12861 26248
rect 12895 26214 12933 26248
rect 12967 26214 13005 26248
rect 13074 26214 13077 26248
rect 13144 26214 13149 26248
rect 13214 26214 13221 26248
rect 13284 26214 13293 26248
rect 13354 26214 13365 26248
rect 13424 26214 13437 26248
rect 13494 26214 13509 26248
rect 13564 26214 13581 26248
rect 9901 26201 13022 26214
rect 13074 26201 13092 26214
rect 13144 26201 13162 26214
rect 13214 26201 13232 26214
rect 13284 26201 13302 26214
rect 13354 26201 13372 26214
rect 13424 26201 13442 26214
rect 13494 26201 13512 26214
rect 13564 26201 13582 26214
rect 13634 26201 13652 26253
rect 13704 26248 14194 26253
rect 13704 26214 13756 26248
rect 13790 26214 13828 26248
rect 13862 26214 13900 26248
rect 13934 26214 13972 26248
rect 14006 26214 14044 26248
rect 14078 26214 14116 26248
rect 14150 26214 14194 26248
rect 13704 26201 14194 26214
rect 9901 26186 14194 26201
rect 9901 26174 13022 26186
rect 13074 26174 13092 26186
rect 13144 26174 13162 26186
rect 13214 26174 13232 26186
rect 13284 26174 13302 26186
rect 13354 26174 13372 26186
rect 13424 26174 13442 26186
rect 13494 26174 13512 26186
rect 13564 26174 13582 26186
rect 9901 26140 9909 26174
rect 9943 26140 9981 26174
rect 10015 26140 10053 26174
rect 10087 26140 10125 26174
rect 10159 26140 10197 26174
rect 10231 26140 10269 26174
rect 10303 26140 10341 26174
rect 10375 26140 10413 26174
rect 10447 26140 10485 26174
rect 10519 26140 10557 26174
rect 10591 26140 10629 26174
rect 10663 26140 10701 26174
rect 10735 26140 10773 26174
rect 10807 26140 10845 26174
rect 10879 26140 10917 26174
rect 10951 26140 10989 26174
rect 11023 26140 11061 26174
rect 11095 26140 11133 26174
rect 11167 26140 11205 26174
rect 11239 26140 11277 26174
rect 11311 26140 11349 26174
rect 11383 26140 11421 26174
rect 11455 26140 11493 26174
rect 11527 26140 11565 26174
rect 11599 26140 11637 26174
rect 11671 26140 11709 26174
rect 11743 26140 11781 26174
rect 11815 26140 11853 26174
rect 11887 26140 11925 26174
rect 11959 26140 11997 26174
rect 12031 26140 12069 26174
rect 12103 26140 12141 26174
rect 12175 26140 12213 26174
rect 12247 26140 12285 26174
rect 12319 26140 12357 26174
rect 12391 26140 12429 26174
rect 12463 26140 12501 26174
rect 12535 26140 12573 26174
rect 12607 26140 12645 26174
rect 12679 26140 12717 26174
rect 12751 26140 12789 26174
rect 12823 26140 12861 26174
rect 12895 26140 12933 26174
rect 12967 26140 13005 26174
rect 13074 26140 13077 26174
rect 13144 26140 13149 26174
rect 13214 26140 13221 26174
rect 13284 26140 13293 26174
rect 13354 26140 13365 26174
rect 13424 26140 13437 26174
rect 13494 26140 13509 26174
rect 13564 26140 13581 26174
rect 9901 26134 13022 26140
rect 13074 26134 13092 26140
rect 13144 26134 13162 26140
rect 13214 26134 13232 26140
rect 13284 26134 13302 26140
rect 13354 26134 13372 26140
rect 13424 26134 13442 26140
rect 13494 26134 13512 26140
rect 13564 26134 13582 26140
rect 13634 26134 13652 26186
rect 13704 26175 14194 26186
rect 13704 26141 13756 26175
rect 13790 26141 13828 26175
rect 13862 26141 13900 26175
rect 13934 26141 13972 26175
rect 14006 26141 14044 26175
rect 14078 26141 14116 26175
rect 14150 26141 14194 26175
rect 13704 26134 14194 26141
rect 9901 26119 14194 26134
rect 9901 26100 13022 26119
rect 13074 26100 13092 26119
rect 13144 26100 13162 26119
rect 13214 26100 13232 26119
rect 13284 26100 13302 26119
rect 13354 26100 13372 26119
rect 13424 26100 13442 26119
rect 13494 26100 13512 26119
rect 13564 26100 13582 26119
rect 9901 26066 9909 26100
rect 9943 26066 9981 26100
rect 10015 26066 10053 26100
rect 10087 26066 10125 26100
rect 10159 26066 10197 26100
rect 10231 26066 10269 26100
rect 10303 26066 10341 26100
rect 10375 26066 10413 26100
rect 10447 26066 10485 26100
rect 10519 26066 10557 26100
rect 10591 26066 10629 26100
rect 10663 26066 10701 26100
rect 10735 26066 10773 26100
rect 10807 26066 10845 26100
rect 10879 26066 10917 26100
rect 10951 26066 10989 26100
rect 11023 26066 11061 26100
rect 11095 26066 11133 26100
rect 11167 26066 11205 26100
rect 11239 26066 11277 26100
rect 11311 26066 11349 26100
rect 11383 26066 11421 26100
rect 11455 26066 11493 26100
rect 11527 26066 11565 26100
rect 11599 26066 11637 26100
rect 11671 26066 11709 26100
rect 11743 26066 11781 26100
rect 11815 26066 11853 26100
rect 11887 26066 11925 26100
rect 11959 26066 11997 26100
rect 12031 26066 12069 26100
rect 12103 26066 12141 26100
rect 12175 26066 12213 26100
rect 12247 26066 12285 26100
rect 12319 26066 12357 26100
rect 12391 26066 12429 26100
rect 12463 26066 12501 26100
rect 12535 26066 12573 26100
rect 12607 26066 12645 26100
rect 12679 26066 12717 26100
rect 12751 26066 12789 26100
rect 12823 26066 12861 26100
rect 12895 26066 12933 26100
rect 12967 26066 13005 26100
rect 13074 26067 13077 26100
rect 13144 26067 13149 26100
rect 13214 26067 13221 26100
rect 13284 26067 13293 26100
rect 13354 26067 13365 26100
rect 13424 26067 13437 26100
rect 13494 26067 13509 26100
rect 13564 26067 13581 26100
rect 13634 26067 13652 26119
rect 13704 26102 14194 26119
rect 13704 26068 13756 26102
rect 13790 26068 13828 26102
rect 13862 26068 13900 26102
rect 13934 26068 13972 26102
rect 14006 26068 14044 26102
rect 14078 26068 14116 26102
rect 14150 26068 14194 26102
rect 13704 26067 14194 26068
rect 13039 26066 13077 26067
rect 13111 26066 13149 26067
rect 13183 26066 13221 26067
rect 13255 26066 13293 26067
rect 13327 26066 13365 26067
rect 13399 26066 13437 26067
rect 13471 26066 13509 26067
rect 13543 26066 13581 26067
rect 13615 26066 13653 26067
rect 13687 26066 14194 26067
rect 9901 26052 14194 26066
rect 9901 26026 13022 26052
rect 13074 26026 13092 26052
rect 13144 26026 13162 26052
rect 13214 26026 13232 26052
rect 13284 26026 13302 26052
rect 13354 26026 13372 26052
rect 13424 26026 13442 26052
rect 13494 26026 13512 26052
rect 13564 26026 13582 26052
rect 9901 25992 9909 26026
rect 9943 25992 9981 26026
rect 10015 25992 10053 26026
rect 10087 25992 10125 26026
rect 10159 25992 10197 26026
rect 10231 25992 10269 26026
rect 10303 25992 10341 26026
rect 10375 25992 10413 26026
rect 10447 25992 10485 26026
rect 10519 25992 10557 26026
rect 10591 25992 10629 26026
rect 10663 25992 10701 26026
rect 10735 25992 10773 26026
rect 10807 25992 10845 26026
rect 10879 25992 10917 26026
rect 10951 25992 10989 26026
rect 11023 25992 11061 26026
rect 11095 25992 11133 26026
rect 11167 25992 11205 26026
rect 11239 25992 11277 26026
rect 11311 25992 11349 26026
rect 11383 25992 11421 26026
rect 11455 25992 11493 26026
rect 11527 25992 11565 26026
rect 11599 25992 11637 26026
rect 11671 25992 11709 26026
rect 11743 25992 11781 26026
rect 11815 25992 11853 26026
rect 11887 25992 11925 26026
rect 11959 25992 11997 26026
rect 12031 25992 12069 26026
rect 12103 25992 12141 26026
rect 12175 25992 12213 26026
rect 12247 25992 12285 26026
rect 12319 25992 12357 26026
rect 12391 25992 12429 26026
rect 12463 25992 12501 26026
rect 12535 25992 12573 26026
rect 12607 25992 12645 26026
rect 12679 25992 12717 26026
rect 12751 25992 12789 26026
rect 12823 25992 12861 26026
rect 12895 25992 12933 26026
rect 12967 25992 13005 26026
rect 13074 26000 13077 26026
rect 13144 26000 13149 26026
rect 13214 26000 13221 26026
rect 13284 26000 13293 26026
rect 13354 26000 13365 26026
rect 13424 26000 13437 26026
rect 13494 26000 13509 26026
rect 13564 26000 13581 26026
rect 13634 26000 13652 26052
rect 13704 26029 14194 26052
rect 13704 26000 13756 26029
rect 13039 25992 13077 26000
rect 13111 25992 13149 26000
rect 13183 25992 13221 26000
rect 13255 25992 13293 26000
rect 13327 25992 13365 26000
rect 13399 25992 13437 26000
rect 13471 25992 13509 26000
rect 13543 25992 13581 26000
rect 13615 25992 13653 26000
rect 13687 25995 13756 26000
rect 13790 25995 13828 26029
rect 13862 25995 13900 26029
rect 13934 25995 13972 26029
rect 14006 25995 14044 26029
rect 14078 25995 14116 26029
rect 14150 25995 14194 26029
rect 13687 25992 14194 25995
rect 9901 25985 14194 25992
rect 9901 25953 13022 25985
rect 13074 25953 13092 25985
rect 13144 25953 13162 25985
rect 13214 25953 13232 25985
rect 13284 25953 13302 25985
rect 13354 25953 13372 25985
rect 13424 25953 13442 25985
rect 13494 25953 13512 25985
rect 13564 25953 13582 25985
rect 9901 25919 9909 25953
rect 9943 25919 9981 25953
rect 10015 25919 10053 25953
rect 10087 25919 10125 25953
rect 10159 25919 10197 25953
rect 10231 25919 10269 25953
rect 10303 25919 10341 25953
rect 10375 25919 10413 25953
rect 10447 25919 10485 25953
rect 10519 25919 10557 25953
rect 10591 25919 10629 25953
rect 10663 25919 10701 25953
rect 10735 25919 10773 25953
rect 10807 25919 10845 25953
rect 10879 25919 10917 25953
rect 10951 25919 10989 25953
rect 11023 25919 11061 25953
rect 11095 25919 11133 25953
rect 11167 25919 11205 25953
rect 11239 25919 11277 25953
rect 11311 25919 11349 25953
rect 11383 25919 11421 25953
rect 11455 25919 11493 25953
rect 11527 25919 11565 25953
rect 11599 25919 11637 25953
rect 11671 25919 11709 25953
rect 11743 25919 11781 25953
rect 11815 25919 11853 25953
rect 11887 25919 11925 25953
rect 11959 25919 11997 25953
rect 12031 25919 12069 25953
rect 12103 25919 12141 25953
rect 12175 25919 12213 25953
rect 12247 25919 12285 25953
rect 12319 25919 12357 25953
rect 12391 25919 12429 25953
rect 12463 25919 12501 25953
rect 12535 25919 12573 25953
rect 12607 25919 12645 25953
rect 12679 25919 12717 25953
rect 12751 25919 12789 25953
rect 12823 25919 12861 25953
rect 12895 25919 12933 25953
rect 12967 25919 13005 25953
rect 13074 25933 13077 25953
rect 13144 25933 13149 25953
rect 13214 25933 13221 25953
rect 13284 25933 13293 25953
rect 13354 25933 13365 25953
rect 13424 25933 13437 25953
rect 13494 25933 13509 25953
rect 13564 25933 13581 25953
rect 13634 25933 13652 25985
rect 13704 25955 14194 25985
rect 13704 25933 13756 25955
rect 13039 25919 13077 25933
rect 13111 25919 13149 25933
rect 13183 25919 13221 25933
rect 13255 25919 13293 25933
rect 13327 25919 13365 25933
rect 13399 25919 13437 25933
rect 13471 25919 13509 25933
rect 13543 25919 13581 25933
rect 13615 25919 13653 25933
rect 13687 25921 13756 25933
rect 13790 25921 13828 25955
rect 13862 25921 13900 25955
rect 13934 25921 13972 25955
rect 14006 25921 14044 25955
rect 14078 25921 14116 25955
rect 14150 25921 14194 25955
rect 13687 25919 14194 25921
rect 9901 25918 14194 25919
rect 9901 25880 13022 25918
rect 13074 25880 13092 25918
rect 13144 25880 13162 25918
rect 13214 25880 13232 25918
rect 13284 25880 13302 25918
rect 13354 25880 13372 25918
rect 13424 25880 13442 25918
rect 13494 25880 13512 25918
rect 13564 25880 13582 25918
rect 9901 25846 9909 25880
rect 9943 25846 9981 25880
rect 10015 25846 10053 25880
rect 10087 25846 10125 25880
rect 10159 25846 10197 25880
rect 10231 25846 10269 25880
rect 10303 25846 10341 25880
rect 10375 25846 10413 25880
rect 10447 25846 10485 25880
rect 10519 25846 10557 25880
rect 10591 25846 10629 25880
rect 10663 25846 10701 25880
rect 10735 25846 10773 25880
rect 10807 25846 10845 25880
rect 10879 25846 10917 25880
rect 10951 25846 10989 25880
rect 11023 25846 11061 25880
rect 11095 25846 11133 25880
rect 11167 25846 11205 25880
rect 11239 25846 11277 25880
rect 11311 25846 11349 25880
rect 11383 25846 11421 25880
rect 11455 25846 11493 25880
rect 11527 25846 11565 25880
rect 11599 25846 11637 25880
rect 11671 25846 11709 25880
rect 11743 25846 11781 25880
rect 11815 25846 11853 25880
rect 11887 25846 11925 25880
rect 11959 25846 11997 25880
rect 12031 25846 12069 25880
rect 12103 25846 12141 25880
rect 12175 25846 12213 25880
rect 12247 25846 12285 25880
rect 12319 25846 12357 25880
rect 12391 25846 12429 25880
rect 12463 25846 12501 25880
rect 12535 25846 12573 25880
rect 12607 25846 12645 25880
rect 12679 25846 12717 25880
rect 12751 25846 12789 25880
rect 12823 25846 12861 25880
rect 12895 25846 12933 25880
rect 12967 25846 13005 25880
rect 13074 25866 13077 25880
rect 13144 25866 13149 25880
rect 13214 25866 13221 25880
rect 13284 25866 13293 25880
rect 13354 25866 13365 25880
rect 13424 25866 13437 25880
rect 13494 25866 13509 25880
rect 13564 25866 13581 25880
rect 13634 25866 13652 25918
rect 13704 25881 14194 25918
rect 13704 25866 13756 25881
rect 13039 25851 13077 25866
rect 13111 25851 13149 25866
rect 13183 25851 13221 25866
rect 13255 25851 13293 25866
rect 13327 25851 13365 25866
rect 13399 25851 13437 25866
rect 13471 25851 13509 25866
rect 13543 25851 13581 25866
rect 13615 25851 13653 25866
rect 13687 25851 13756 25866
rect 13074 25846 13077 25851
rect 13144 25846 13149 25851
rect 13214 25846 13221 25851
rect 13284 25846 13293 25851
rect 13354 25846 13365 25851
rect 13424 25846 13437 25851
rect 13494 25846 13509 25851
rect 13564 25846 13581 25851
rect 9901 25807 13022 25846
rect 13074 25807 13092 25846
rect 13144 25807 13162 25846
rect 13214 25807 13232 25846
rect 13284 25807 13302 25846
rect 13354 25807 13372 25846
rect 13424 25807 13442 25846
rect 13494 25807 13512 25846
rect 13564 25807 13582 25846
rect 9901 25773 9909 25807
rect 9943 25773 9981 25807
rect 10015 25773 10053 25807
rect 10087 25773 10125 25807
rect 10159 25773 10197 25807
rect 10231 25773 10269 25807
rect 10303 25773 10341 25807
rect 10375 25773 10413 25807
rect 10447 25773 10485 25807
rect 10519 25773 10557 25807
rect 10591 25773 10629 25807
rect 10663 25773 10701 25807
rect 10735 25773 10773 25807
rect 10807 25773 10845 25807
rect 10879 25773 10917 25807
rect 10951 25773 10989 25807
rect 11023 25773 11061 25807
rect 11095 25773 11133 25807
rect 11167 25773 11205 25807
rect 11239 25773 11277 25807
rect 11311 25773 11349 25807
rect 11383 25773 11421 25807
rect 11455 25773 11493 25807
rect 11527 25773 11565 25807
rect 11599 25773 11637 25807
rect 11671 25773 11709 25807
rect 11743 25773 11781 25807
rect 11815 25773 11853 25807
rect 11887 25773 11925 25807
rect 11959 25773 11997 25807
rect 12031 25773 12069 25807
rect 12103 25773 12141 25807
rect 12175 25773 12213 25807
rect 12247 25773 12285 25807
rect 12319 25773 12357 25807
rect 12391 25773 12429 25807
rect 12463 25773 12501 25807
rect 12535 25773 12573 25807
rect 12607 25773 12645 25807
rect 12679 25773 12717 25807
rect 12751 25773 12789 25807
rect 12823 25773 12861 25807
rect 12895 25773 12933 25807
rect 12967 25773 13005 25807
rect 13074 25799 13077 25807
rect 13144 25799 13149 25807
rect 13214 25799 13221 25807
rect 13284 25799 13293 25807
rect 13354 25799 13365 25807
rect 13424 25799 13437 25807
rect 13494 25799 13509 25807
rect 13564 25799 13581 25807
rect 13634 25799 13652 25851
rect 13704 25847 13756 25851
rect 13790 25847 13828 25881
rect 13862 25847 13900 25881
rect 13934 25847 13972 25881
rect 14006 25847 14044 25881
rect 14078 25847 14116 25881
rect 14150 25847 14194 25881
rect 13704 25807 14194 25847
rect 13704 25799 13756 25807
rect 13039 25784 13077 25799
rect 13111 25784 13149 25799
rect 13183 25784 13221 25799
rect 13255 25784 13293 25799
rect 13327 25784 13365 25799
rect 13399 25784 13437 25799
rect 13471 25784 13509 25799
rect 13543 25784 13581 25799
rect 13615 25784 13653 25799
rect 13687 25784 13756 25799
rect 13074 25773 13077 25784
rect 13144 25773 13149 25784
rect 13214 25773 13221 25784
rect 13284 25773 13293 25784
rect 13354 25773 13365 25784
rect 13424 25773 13437 25784
rect 13494 25773 13509 25784
rect 13564 25773 13581 25784
rect 9901 25734 13022 25773
rect 13074 25734 13092 25773
rect 13144 25734 13162 25773
rect 13214 25734 13232 25773
rect 13284 25734 13302 25773
rect 13354 25734 13372 25773
rect 13424 25734 13442 25773
rect 13494 25734 13512 25773
rect 13564 25734 13582 25773
rect 9901 25700 9909 25734
rect 9943 25700 9981 25734
rect 10015 25700 10053 25734
rect 10087 25700 10125 25734
rect 10159 25700 10197 25734
rect 10231 25700 10269 25734
rect 10303 25700 10341 25734
rect 10375 25700 10413 25734
rect 10447 25700 10485 25734
rect 10519 25700 10557 25734
rect 10591 25700 10629 25734
rect 10663 25700 10701 25734
rect 10735 25700 10773 25734
rect 10807 25700 10845 25734
rect 10879 25700 10917 25734
rect 10951 25700 10989 25734
rect 11023 25700 11061 25734
rect 11095 25700 11133 25734
rect 11167 25700 11205 25734
rect 11239 25700 11277 25734
rect 11311 25700 11349 25734
rect 11383 25700 11421 25734
rect 11455 25700 11493 25734
rect 11527 25700 11565 25734
rect 11599 25700 11637 25734
rect 11671 25700 11709 25734
rect 11743 25700 11781 25734
rect 11815 25700 11853 25734
rect 11887 25700 11925 25734
rect 11959 25700 11997 25734
rect 12031 25700 12069 25734
rect 12103 25700 12141 25734
rect 12175 25700 12213 25734
rect 12247 25700 12285 25734
rect 12319 25700 12357 25734
rect 12391 25700 12429 25734
rect 12463 25700 12501 25734
rect 12535 25700 12573 25734
rect 12607 25700 12645 25734
rect 12679 25700 12717 25734
rect 12751 25700 12789 25734
rect 12823 25700 12861 25734
rect 12895 25700 12933 25734
rect 12967 25700 13005 25734
rect 13074 25732 13077 25734
rect 13144 25732 13149 25734
rect 13214 25732 13221 25734
rect 13284 25732 13293 25734
rect 13354 25732 13365 25734
rect 13424 25732 13437 25734
rect 13494 25732 13509 25734
rect 13564 25732 13581 25734
rect 13634 25732 13652 25784
rect 13704 25773 13756 25784
rect 13790 25773 13828 25807
rect 13862 25773 13900 25807
rect 13934 25773 13972 25807
rect 14006 25773 14044 25807
rect 14078 25773 14116 25807
rect 14150 25773 14194 25807
rect 13704 25733 14194 25773
rect 13704 25732 13756 25733
rect 13039 25717 13077 25732
rect 13111 25717 13149 25732
rect 13183 25717 13221 25732
rect 13255 25717 13293 25732
rect 13327 25717 13365 25732
rect 13399 25717 13437 25732
rect 13471 25717 13509 25732
rect 13543 25717 13581 25732
rect 13615 25717 13653 25732
rect 13687 25717 13756 25732
rect 13074 25700 13077 25717
rect 13144 25700 13149 25717
rect 13214 25700 13221 25717
rect 13284 25700 13293 25717
rect 13354 25700 13365 25717
rect 13424 25700 13437 25717
rect 13494 25700 13509 25717
rect 13564 25700 13581 25717
rect 9901 25665 13022 25700
rect 13074 25665 13092 25700
rect 13144 25665 13162 25700
rect 13214 25665 13232 25700
rect 13284 25665 13302 25700
rect 13354 25665 13372 25700
rect 13424 25665 13442 25700
rect 13494 25665 13512 25700
rect 13564 25665 13582 25700
rect 13634 25665 13652 25717
rect 13704 25699 13756 25717
rect 13790 25699 13828 25733
rect 13862 25699 13900 25733
rect 13934 25699 13972 25733
rect 14006 25699 14044 25733
rect 14078 25699 14116 25733
rect 14150 25699 14194 25733
rect 13704 25665 14194 25699
rect 9901 25661 14194 25665
rect 9901 25627 9909 25661
rect 9943 25627 9981 25661
rect 10015 25627 10053 25661
rect 10087 25627 10125 25661
rect 10159 25627 10197 25661
rect 10231 25627 10269 25661
rect 10303 25627 10341 25661
rect 10375 25627 10413 25661
rect 10447 25627 10485 25661
rect 10519 25627 10557 25661
rect 10591 25627 10629 25661
rect 10663 25627 10701 25661
rect 10735 25627 10773 25661
rect 10807 25627 10845 25661
rect 10879 25627 10917 25661
rect 10951 25627 10989 25661
rect 11023 25627 11061 25661
rect 11095 25627 11133 25661
rect 11167 25627 11205 25661
rect 11239 25627 11277 25661
rect 11311 25627 11349 25661
rect 11383 25627 11421 25661
rect 11455 25627 11493 25661
rect 11527 25627 11565 25661
rect 11599 25627 11637 25661
rect 11671 25627 11709 25661
rect 11743 25627 11781 25661
rect 11815 25627 11853 25661
rect 11887 25627 11925 25661
rect 11959 25627 11997 25661
rect 12031 25627 12069 25661
rect 12103 25627 12141 25661
rect 12175 25627 12213 25661
rect 12247 25627 12285 25661
rect 12319 25627 12357 25661
rect 12391 25627 12429 25661
rect 12463 25627 12501 25661
rect 12535 25627 12573 25661
rect 12607 25627 12645 25661
rect 12679 25627 12717 25661
rect 12751 25627 12789 25661
rect 12823 25627 12861 25661
rect 12895 25627 12933 25661
rect 12967 25627 13005 25661
rect 13039 25650 13077 25661
rect 13111 25650 13149 25661
rect 13183 25650 13221 25661
rect 13255 25650 13293 25661
rect 13327 25650 13365 25661
rect 13399 25650 13437 25661
rect 13471 25650 13509 25661
rect 13543 25650 13581 25661
rect 13615 25650 13653 25661
rect 13687 25659 14194 25661
rect 13687 25650 13756 25659
rect 13074 25627 13077 25650
rect 13144 25627 13149 25650
rect 13214 25627 13221 25650
rect 13284 25627 13293 25650
rect 13354 25627 13365 25650
rect 13424 25627 13437 25650
rect 13494 25627 13509 25650
rect 13564 25627 13581 25650
rect 9901 25598 13022 25627
rect 13074 25598 13092 25627
rect 13144 25598 13162 25627
rect 13214 25598 13232 25627
rect 13284 25598 13302 25627
rect 13354 25598 13372 25627
rect 13424 25598 13442 25627
rect 13494 25598 13512 25627
rect 13564 25598 13582 25627
rect 13634 25598 13652 25650
rect 13704 25625 13756 25650
rect 13790 25625 13828 25659
rect 13862 25625 13900 25659
rect 13934 25625 13972 25659
rect 14006 25625 14044 25659
rect 14078 25625 14116 25659
rect 14150 25625 14194 25659
rect 13704 25598 14194 25625
rect 9901 25588 14194 25598
rect 9901 25554 9909 25588
rect 9943 25554 9981 25588
rect 10015 25554 10053 25588
rect 10087 25554 10125 25588
rect 10159 25554 10197 25588
rect 10231 25554 10269 25588
rect 10303 25554 10341 25588
rect 10375 25554 10413 25588
rect 10447 25554 10485 25588
rect 10519 25554 10557 25588
rect 10591 25554 10629 25588
rect 10663 25554 10701 25588
rect 10735 25554 10773 25588
rect 10807 25554 10845 25588
rect 10879 25554 10917 25588
rect 10951 25554 10989 25588
rect 11023 25554 11061 25588
rect 11095 25554 11133 25588
rect 11167 25554 11205 25588
rect 11239 25554 11277 25588
rect 11311 25554 11349 25588
rect 11383 25554 11421 25588
rect 11455 25554 11493 25588
rect 11527 25554 11565 25588
rect 11599 25554 11637 25588
rect 11671 25554 11709 25588
rect 11743 25554 11781 25588
rect 11815 25554 11853 25588
rect 11887 25554 11925 25588
rect 11959 25554 11997 25588
rect 12031 25554 12069 25588
rect 12103 25554 12141 25588
rect 12175 25554 12213 25588
rect 12247 25554 12285 25588
rect 12319 25554 12357 25588
rect 12391 25554 12429 25588
rect 12463 25554 12501 25588
rect 12535 25554 12573 25588
rect 12607 25554 12645 25588
rect 12679 25554 12717 25588
rect 12751 25554 12789 25588
rect 12823 25554 12861 25588
rect 12895 25554 12933 25588
rect 12967 25554 13005 25588
rect 13039 25582 13077 25588
rect 13111 25582 13149 25588
rect 13183 25582 13221 25588
rect 13255 25582 13293 25588
rect 13327 25582 13365 25588
rect 13399 25582 13437 25588
rect 13471 25582 13509 25588
rect 13543 25582 13581 25588
rect 13615 25582 13653 25588
rect 13687 25585 14194 25588
rect 13687 25582 13756 25585
rect 13074 25554 13077 25582
rect 13144 25554 13149 25582
rect 13214 25554 13221 25582
rect 13284 25554 13293 25582
rect 13354 25554 13365 25582
rect 13424 25554 13437 25582
rect 13494 25554 13509 25582
rect 13564 25554 13581 25582
rect 9901 25530 13022 25554
rect 13074 25530 13092 25554
rect 13144 25530 13162 25554
rect 13214 25530 13232 25554
rect 13284 25530 13302 25554
rect 13354 25530 13372 25554
rect 13424 25530 13442 25554
rect 13494 25530 13512 25554
rect 13564 25530 13582 25554
rect 13634 25530 13652 25582
rect 13704 25551 13756 25582
rect 13790 25551 13828 25585
rect 13862 25551 13900 25585
rect 13934 25551 13972 25585
rect 14006 25551 14044 25585
rect 14078 25551 14116 25585
rect 14150 25551 14194 25585
rect 13704 25530 14194 25551
rect 9901 25515 14194 25530
rect 9901 25481 9909 25515
rect 9943 25481 9981 25515
rect 10015 25481 10053 25515
rect 10087 25481 10125 25515
rect 10159 25481 10197 25515
rect 10231 25481 10269 25515
rect 10303 25481 10341 25515
rect 10375 25481 10413 25515
rect 10447 25481 10485 25515
rect 10519 25481 10557 25515
rect 10591 25481 10629 25515
rect 10663 25481 10701 25515
rect 10735 25481 10773 25515
rect 10807 25481 10845 25515
rect 10879 25481 10917 25515
rect 10951 25481 10989 25515
rect 11023 25481 11061 25515
rect 11095 25481 11133 25515
rect 11167 25481 11205 25515
rect 11239 25481 11277 25515
rect 11311 25481 11349 25515
rect 11383 25481 11421 25515
rect 11455 25481 11493 25515
rect 11527 25481 11565 25515
rect 11599 25481 11637 25515
rect 11671 25481 11709 25515
rect 11743 25481 11781 25515
rect 11815 25481 11853 25515
rect 11887 25481 11925 25515
rect 11959 25481 11997 25515
rect 12031 25481 12069 25515
rect 12103 25481 12141 25515
rect 12175 25481 12213 25515
rect 12247 25481 12285 25515
rect 12319 25481 12357 25515
rect 12391 25481 12429 25515
rect 12463 25481 12501 25515
rect 12535 25481 12573 25515
rect 12607 25481 12645 25515
rect 12679 25481 12717 25515
rect 12751 25481 12789 25515
rect 12823 25481 12861 25515
rect 12895 25481 12933 25515
rect 12967 25481 13005 25515
rect 13039 25514 13077 25515
rect 13111 25514 13149 25515
rect 13183 25514 13221 25515
rect 13255 25514 13293 25515
rect 13327 25514 13365 25515
rect 13399 25514 13437 25515
rect 13471 25514 13509 25515
rect 13543 25514 13581 25515
rect 13615 25514 13653 25515
rect 13687 25514 14194 25515
rect 13074 25481 13077 25514
rect 13144 25481 13149 25514
rect 13214 25481 13221 25514
rect 13284 25481 13293 25514
rect 13354 25481 13365 25514
rect 13424 25481 13437 25514
rect 13494 25481 13509 25514
rect 13564 25481 13581 25514
rect 9901 25462 13022 25481
rect 13074 25462 13092 25481
rect 13144 25462 13162 25481
rect 13214 25462 13232 25481
rect 13284 25462 13302 25481
rect 13354 25462 13372 25481
rect 13424 25462 13442 25481
rect 13494 25462 13512 25481
rect 13564 25462 13582 25481
rect 13634 25462 13652 25514
rect 13704 25511 14194 25514
rect 13704 25477 13756 25511
rect 13790 25477 13828 25511
rect 13862 25477 13900 25511
rect 13934 25477 13972 25511
rect 14006 25477 14044 25511
rect 14078 25477 14116 25511
rect 14150 25477 14194 25511
rect 13704 25462 14194 25477
rect 9901 25446 14194 25462
rect 9901 25442 13022 25446
rect 13074 25442 13092 25446
rect 13144 25442 13162 25446
rect 13214 25442 13232 25446
rect 13284 25442 13302 25446
rect 13354 25442 13372 25446
rect 13424 25442 13442 25446
rect 13494 25442 13512 25446
rect 13564 25442 13582 25446
rect 9901 25408 9909 25442
rect 9943 25408 9981 25442
rect 10015 25408 10053 25442
rect 10087 25408 10125 25442
rect 10159 25408 10197 25442
rect 10231 25408 10269 25442
rect 10303 25408 10341 25442
rect 10375 25408 10413 25442
rect 10447 25408 10485 25442
rect 10519 25408 10557 25442
rect 10591 25408 10629 25442
rect 10663 25408 10701 25442
rect 10735 25408 10773 25442
rect 10807 25408 10845 25442
rect 10879 25408 10917 25442
rect 10951 25408 10989 25442
rect 11023 25408 11061 25442
rect 11095 25408 11133 25442
rect 11167 25408 11205 25442
rect 11239 25408 11277 25442
rect 11311 25408 11349 25442
rect 11383 25408 11421 25442
rect 11455 25408 11493 25442
rect 11527 25408 11565 25442
rect 11599 25408 11637 25442
rect 11671 25408 11709 25442
rect 11743 25408 11781 25442
rect 11815 25408 11853 25442
rect 11887 25408 11925 25442
rect 11959 25408 11997 25442
rect 12031 25408 12069 25442
rect 12103 25408 12141 25442
rect 12175 25408 12213 25442
rect 12247 25408 12285 25442
rect 12319 25408 12357 25442
rect 12391 25408 12429 25442
rect 12463 25408 12501 25442
rect 12535 25408 12573 25442
rect 12607 25408 12645 25442
rect 12679 25408 12717 25442
rect 12751 25408 12789 25442
rect 12823 25408 12861 25442
rect 12895 25408 12933 25442
rect 12967 25408 13005 25442
rect 13074 25408 13077 25442
rect 13144 25408 13149 25442
rect 13214 25408 13221 25442
rect 13284 25408 13293 25442
rect 13354 25408 13365 25442
rect 13424 25408 13437 25442
rect 13494 25408 13509 25442
rect 13564 25408 13581 25442
rect 9901 25394 13022 25408
rect 13074 25394 13092 25408
rect 13144 25394 13162 25408
rect 13214 25394 13232 25408
rect 13284 25394 13302 25408
rect 13354 25394 13372 25408
rect 13424 25394 13442 25408
rect 13494 25394 13512 25408
rect 13564 25394 13582 25408
rect 13634 25394 13652 25446
rect 13704 25437 14194 25446
rect 13704 25403 13756 25437
rect 13790 25403 13828 25437
rect 13862 25403 13900 25437
rect 13934 25403 13972 25437
rect 14006 25403 14044 25437
rect 14078 25403 14116 25437
rect 14150 25403 14194 25437
rect 13704 25394 14194 25403
rect 9901 25378 14194 25394
rect 9901 25369 13022 25378
rect 13074 25369 13092 25378
rect 13144 25369 13162 25378
rect 13214 25369 13232 25378
rect 13284 25369 13302 25378
rect 13354 25369 13372 25378
rect 13424 25369 13442 25378
rect 13494 25369 13512 25378
rect 13564 25369 13582 25378
rect 9901 25335 9909 25369
rect 9943 25335 9981 25369
rect 10015 25335 10053 25369
rect 10087 25335 10125 25369
rect 10159 25335 10197 25369
rect 10231 25335 10269 25369
rect 10303 25335 10341 25369
rect 10375 25335 10413 25369
rect 10447 25335 10485 25369
rect 10519 25335 10557 25369
rect 10591 25335 10629 25369
rect 10663 25335 10701 25369
rect 10735 25335 10773 25369
rect 10807 25335 10845 25369
rect 10879 25335 10917 25369
rect 10951 25335 10989 25369
rect 11023 25335 11061 25369
rect 11095 25335 11133 25369
rect 11167 25335 11205 25369
rect 11239 25335 11277 25369
rect 11311 25335 11349 25369
rect 11383 25335 11421 25369
rect 11455 25335 11493 25369
rect 11527 25335 11565 25369
rect 11599 25335 11637 25369
rect 11671 25335 11709 25369
rect 11743 25335 11781 25369
rect 11815 25335 11853 25369
rect 11887 25335 11925 25369
rect 11959 25335 11997 25369
rect 12031 25335 12069 25369
rect 12103 25335 12141 25369
rect 12175 25335 12213 25369
rect 12247 25335 12285 25369
rect 12319 25335 12357 25369
rect 12391 25335 12429 25369
rect 12463 25335 12501 25369
rect 12535 25335 12573 25369
rect 12607 25335 12645 25369
rect 12679 25335 12717 25369
rect 12751 25335 12789 25369
rect 12823 25335 12861 25369
rect 12895 25335 12933 25369
rect 12967 25335 13005 25369
rect 13074 25335 13077 25369
rect 13144 25335 13149 25369
rect 13214 25335 13221 25369
rect 13284 25335 13293 25369
rect 13354 25335 13365 25369
rect 13424 25335 13437 25369
rect 13494 25335 13509 25369
rect 13564 25335 13581 25369
rect 9901 25326 13022 25335
rect 13074 25326 13092 25335
rect 13144 25326 13162 25335
rect 13214 25326 13232 25335
rect 13284 25326 13302 25335
rect 13354 25326 13372 25335
rect 13424 25326 13442 25335
rect 13494 25326 13512 25335
rect 13564 25326 13582 25335
rect 13634 25326 13652 25378
rect 13704 25363 14194 25378
rect 13704 25329 13756 25363
rect 13790 25329 13828 25363
rect 13862 25329 13900 25363
rect 13934 25329 13972 25363
rect 14006 25329 14044 25363
rect 14078 25329 14116 25363
rect 14150 25329 14194 25363
rect 13704 25326 14194 25329
rect 9901 25310 14194 25326
rect 9901 25296 13022 25310
rect 13074 25296 13092 25310
rect 13144 25296 13162 25310
rect 13214 25296 13232 25310
rect 13284 25296 13302 25310
rect 13354 25296 13372 25310
rect 13424 25296 13442 25310
rect 13494 25296 13512 25310
rect 13564 25296 13582 25310
rect 9901 25262 9909 25296
rect 9943 25262 9981 25296
rect 10015 25262 10053 25296
rect 10087 25262 10125 25296
rect 10159 25262 10197 25296
rect 10231 25262 10269 25296
rect 10303 25262 10341 25296
rect 10375 25262 10413 25296
rect 10447 25262 10485 25296
rect 10519 25262 10557 25296
rect 10591 25262 10629 25296
rect 10663 25262 10701 25296
rect 10735 25262 10773 25296
rect 10807 25262 10845 25296
rect 10879 25262 10917 25296
rect 10951 25262 10989 25296
rect 11023 25262 11061 25296
rect 11095 25262 11133 25296
rect 11167 25262 11205 25296
rect 11239 25262 11277 25296
rect 11311 25262 11349 25296
rect 11383 25262 11421 25296
rect 11455 25262 11493 25296
rect 11527 25262 11565 25296
rect 11599 25262 11637 25296
rect 11671 25262 11709 25296
rect 11743 25262 11781 25296
rect 11815 25262 11853 25296
rect 11887 25262 11925 25296
rect 11959 25262 11997 25296
rect 12031 25262 12069 25296
rect 12103 25262 12141 25296
rect 12175 25262 12213 25296
rect 12247 25262 12285 25296
rect 12319 25262 12357 25296
rect 12391 25262 12429 25296
rect 12463 25262 12501 25296
rect 12535 25262 12573 25296
rect 12607 25262 12645 25296
rect 12679 25262 12717 25296
rect 12751 25262 12789 25296
rect 12823 25262 12861 25296
rect 12895 25262 12933 25296
rect 12967 25262 13005 25296
rect 13074 25262 13077 25296
rect 13144 25262 13149 25296
rect 13214 25262 13221 25296
rect 13284 25262 13293 25296
rect 13354 25262 13365 25296
rect 13424 25262 13437 25296
rect 13494 25262 13509 25296
rect 13564 25262 13581 25296
rect 9901 25258 13022 25262
rect 13074 25258 13092 25262
rect 13144 25258 13162 25262
rect 13214 25258 13232 25262
rect 13284 25258 13302 25262
rect 13354 25258 13372 25262
rect 13424 25258 13442 25262
rect 13494 25258 13512 25262
rect 13564 25258 13582 25262
rect 13634 25258 13652 25310
rect 13704 25289 14194 25310
rect 13704 25258 13756 25289
rect 9901 25255 13756 25258
rect 13790 25255 13828 25289
rect 13862 25255 13900 25289
rect 13934 25255 13972 25289
rect 14006 25255 14044 25289
rect 14078 25255 14116 25289
rect 14150 25255 14194 25289
rect 9901 25253 14194 25255
tri 14194 25253 14403 25462 sw
rect 9901 25242 14403 25253
rect 9901 25223 13022 25242
rect 13074 25223 13092 25242
rect 13144 25223 13162 25242
rect 13214 25223 13232 25242
rect 13284 25223 13302 25242
rect 13354 25223 13372 25242
rect 13424 25223 13442 25242
rect 13494 25223 13512 25242
rect 13564 25223 13582 25242
rect 9901 25189 9909 25223
rect 9943 25189 9981 25223
rect 10015 25189 10053 25223
rect 10087 25189 10125 25223
rect 10159 25189 10197 25223
rect 10231 25189 10269 25223
rect 10303 25189 10341 25223
rect 10375 25189 10413 25223
rect 10447 25189 10485 25223
rect 10519 25189 10557 25223
rect 10591 25189 10629 25223
rect 10663 25189 10701 25223
rect 10735 25189 10773 25223
rect 10807 25189 10845 25223
rect 10879 25189 10917 25223
rect 10951 25189 10989 25223
rect 11023 25189 11061 25223
rect 11095 25189 11133 25223
rect 11167 25189 11205 25223
rect 11239 25189 11277 25223
rect 11311 25189 11349 25223
rect 11383 25189 11421 25223
rect 11455 25189 11493 25223
rect 11527 25189 11565 25223
rect 11599 25189 11637 25223
rect 11671 25189 11709 25223
rect 11743 25189 11781 25223
rect 11815 25189 11853 25223
rect 11887 25189 11925 25223
rect 11959 25189 11997 25223
rect 12031 25189 12069 25223
rect 12103 25189 12141 25223
rect 12175 25189 12213 25223
rect 12247 25189 12285 25223
rect 12319 25189 12357 25223
rect 12391 25189 12429 25223
rect 12463 25189 12501 25223
rect 12535 25189 12573 25223
rect 12607 25189 12645 25223
rect 12679 25189 12717 25223
rect 12751 25189 12789 25223
rect 12823 25189 12861 25223
rect 12895 25189 12933 25223
rect 12967 25189 13005 25223
rect 13074 25190 13077 25223
rect 13144 25190 13149 25223
rect 13214 25190 13221 25223
rect 13284 25190 13293 25223
rect 13354 25190 13365 25223
rect 13424 25190 13437 25223
rect 13494 25190 13509 25223
rect 13564 25190 13581 25223
rect 13634 25190 13652 25242
rect 13704 25241 14403 25242
rect 13704 25215 14252 25241
rect 13704 25190 13756 25215
rect 13039 25189 13077 25190
rect 13111 25189 13149 25190
rect 13183 25189 13221 25190
rect 13255 25189 13293 25190
rect 13327 25189 13365 25190
rect 13399 25189 13437 25190
rect 13471 25189 13509 25190
rect 13543 25189 13581 25190
rect 13615 25189 13653 25190
rect 13687 25189 13756 25190
rect 9901 25181 13756 25189
rect 13790 25181 13828 25215
rect 13862 25181 13900 25215
rect 13934 25181 13972 25215
rect 14006 25181 14044 25215
rect 14078 25181 14116 25215
rect 14150 25207 14252 25215
rect 14286 25207 14324 25241
rect 14358 25207 14403 25241
rect 14150 25181 14403 25207
rect 9901 25174 14403 25181
rect 9901 25150 13022 25174
rect 13074 25150 13092 25174
rect 13144 25150 13162 25174
rect 13214 25150 13232 25174
rect 13284 25150 13302 25174
rect 13354 25150 13372 25174
rect 13424 25150 13442 25174
rect 13494 25150 13512 25174
rect 13564 25150 13582 25174
rect 6814 25017 7070 25135
rect 9901 25116 9909 25150
rect 9943 25116 9981 25150
rect 10015 25116 10053 25150
rect 10087 25116 10125 25150
rect 10159 25116 10197 25150
rect 10231 25116 10269 25150
rect 10303 25116 10341 25150
rect 10375 25116 10413 25150
rect 10447 25116 10485 25150
rect 10519 25116 10557 25150
rect 10591 25116 10629 25150
rect 10663 25116 10701 25150
rect 10735 25116 10773 25150
rect 10807 25116 10845 25150
rect 10879 25116 10917 25150
rect 10951 25116 10989 25150
rect 11023 25116 11061 25150
rect 11095 25116 11133 25150
rect 11167 25116 11205 25150
rect 11239 25116 11277 25150
rect 11311 25116 11349 25150
rect 11383 25116 11421 25150
rect 11455 25116 11493 25150
rect 11527 25116 11565 25150
rect 11599 25116 11637 25150
rect 11671 25116 11709 25150
rect 11743 25116 11781 25150
rect 11815 25116 11853 25150
rect 11887 25116 11925 25150
rect 11959 25116 11997 25150
rect 12031 25116 12069 25150
rect 12103 25116 12141 25150
rect 12175 25116 12213 25150
rect 12247 25116 12285 25150
rect 12319 25116 12357 25150
rect 12391 25116 12429 25150
rect 12463 25116 12501 25150
rect 12535 25116 12573 25150
rect 12607 25116 12645 25150
rect 12679 25116 12717 25150
rect 12751 25116 12789 25150
rect 12823 25116 12861 25150
rect 12895 25116 12933 25150
rect 12967 25116 13005 25150
rect 13074 25122 13077 25150
rect 13144 25122 13149 25150
rect 13214 25122 13221 25150
rect 13284 25122 13293 25150
rect 13354 25122 13365 25150
rect 13424 25122 13437 25150
rect 13494 25122 13509 25150
rect 13564 25122 13581 25150
rect 13634 25122 13652 25174
rect 13704 25168 14403 25174
rect 13704 25141 14252 25168
rect 13704 25122 13756 25141
rect 13039 25116 13077 25122
rect 13111 25116 13149 25122
rect 13183 25116 13221 25122
rect 13255 25116 13293 25122
rect 13327 25116 13365 25122
rect 13399 25116 13437 25122
rect 13471 25116 13509 25122
rect 13543 25116 13581 25122
rect 13615 25116 13653 25122
rect 13687 25116 13756 25122
rect 9901 25107 13756 25116
rect 13790 25107 13828 25141
rect 13862 25107 13900 25141
rect 13934 25107 13972 25141
rect 14006 25107 14044 25141
rect 14078 25107 14116 25141
rect 14150 25134 14252 25141
rect 14286 25134 14324 25168
rect 14358 25134 14403 25168
rect 14150 25107 14403 25134
rect 9901 25103 14403 25107
tri 8474 25067 8481 25074 se
rect 8481 25067 8497 25074
tri 8440 25033 8474 25067 se
rect 8474 25033 8497 25067
tri 8429 25022 8440 25033 se
rect 8440 25022 8497 25033
rect 8549 25022 8561 25074
rect 8613 25022 8619 25074
tri 8424 25017 8429 25022 se
rect 8429 25019 8619 25022
rect 8429 25017 8610 25019
tri 8417 25010 8424 25017 se
rect 8424 25010 8610 25017
tri 8610 25010 8619 25019 nw
tri 8396 24989 8417 25010 se
rect 8417 24989 8433 25010
rect 5800 24937 5806 24989
rect 5858 24937 5870 24989
rect 5922 24958 8433 24989
rect 8485 24958 8497 25010
rect 8549 24988 8588 25010
tri 8588 24988 8610 25010 nw
rect 8549 24958 8558 24988
tri 8558 24958 8588 24988 nw
rect 5922 24949 8549 24958
tri 8549 24949 8558 24958 nw
rect 5922 24937 8537 24949
tri 8537 24937 8549 24949 nw
rect 5947 24857 5953 24909
rect 6005 24857 6017 24909
rect 6069 24857 8497 24909
rect 8549 24857 8561 24909
rect 8613 24857 8619 24909
rect 9901 24562 11240 25103
tri 13642 25095 13650 25103 ne
rect 13650 25095 14403 25103
tri 13650 25067 13678 25095 ne
rect 13678 25067 14252 25095
tri 13678 25033 13712 25067 ne
rect 13712 25033 13756 25067
rect 13790 25033 13828 25067
rect 13862 25033 13900 25067
rect 13934 25033 13972 25067
rect 14006 25033 14044 25067
rect 14078 25033 14116 25067
rect 14150 25061 14252 25067
rect 14286 25061 14324 25095
rect 14358 25061 14403 25095
rect 14150 25033 14403 25061
tri 13712 25022 13723 25033 ne
rect 13723 25022 14403 25033
tri 13723 25021 13724 25022 ne
rect 13724 25021 14252 25022
tri 13724 24988 13757 25021 ne
rect 13757 24988 14252 25021
rect 14286 24988 14324 25022
rect 14358 24988 14403 25022
tri 13757 24949 13796 24988 ne
rect 13796 24949 14403 24988
tri 13796 24915 13830 24949 ne
rect 13830 24915 14252 24949
rect 14286 24915 14324 24949
rect 14358 24915 14403 24949
tri 13830 24876 13869 24915 ne
rect 13869 24876 14403 24915
tri 13869 24842 13903 24876 ne
rect 13903 24842 14252 24876
rect 14286 24842 14324 24876
rect 14358 24842 14403 24876
tri 13903 24803 13942 24842 ne
rect 13942 24803 14403 24842
tri 13942 24769 13976 24803 ne
rect 13976 24769 14252 24803
rect 14286 24769 14324 24803
rect 14358 24769 14403 24803
tri 13976 24730 14015 24769 ne
rect 14015 24730 14403 24769
tri 14015 24696 14049 24730 ne
rect 14049 24696 14252 24730
rect 14286 24696 14324 24730
rect 14358 24696 14403 24730
tri 14049 24692 14053 24696 ne
rect 9901 24528 9914 24562
rect 9948 24528 9990 24562
rect 10024 24528 10066 24562
rect 10100 24528 10142 24562
rect 10176 24528 10218 24562
rect 10252 24528 10294 24562
rect 10328 24528 10369 24562
rect 10403 24528 10444 24562
rect 10478 24528 10519 24562
rect 10553 24528 10594 24562
rect 10628 24528 10669 24562
rect 10703 24528 10744 24562
rect 10778 24528 10819 24562
rect 10853 24528 10894 24562
rect 10928 24528 10969 24562
rect 11003 24528 11044 24562
rect 11078 24528 11119 24562
rect 11153 24528 11194 24562
rect 11228 24528 11240 24562
rect 9901 24490 11240 24528
rect 9901 24456 9914 24490
rect 9948 24456 9990 24490
rect 10024 24456 10066 24490
rect 10100 24456 10142 24490
rect 10176 24456 10218 24490
rect 10252 24456 10294 24490
rect 10328 24456 10369 24490
rect 10403 24456 10444 24490
rect 10478 24456 10519 24490
rect 10553 24456 10594 24490
rect 10628 24456 10669 24490
rect 10703 24456 10744 24490
rect 10778 24456 10819 24490
rect 10853 24456 10894 24490
rect 10928 24456 10969 24490
rect 11003 24456 11044 24490
rect 11078 24456 11119 24490
rect 11153 24456 11194 24490
rect 11228 24456 11240 24490
rect 9901 24418 11240 24456
rect 9901 24384 9914 24418
rect 9948 24384 9990 24418
rect 10024 24384 10066 24418
rect 10100 24384 10142 24418
rect 10176 24384 10218 24418
rect 10252 24384 10294 24418
rect 10328 24384 10369 24418
rect 10403 24384 10444 24418
rect 10478 24384 10519 24418
rect 10553 24384 10594 24418
rect 10628 24384 10669 24418
rect 10703 24384 10744 24418
rect 10778 24384 10819 24418
rect 10853 24384 10894 24418
rect 10928 24384 10969 24418
rect 11003 24384 11044 24418
rect 11078 24384 11119 24418
rect 11153 24384 11194 24418
rect 11228 24384 11240 24418
rect 9901 24346 11240 24384
rect 9901 24312 9914 24346
rect 9948 24312 9990 24346
rect 10024 24312 10066 24346
rect 10100 24312 10142 24346
rect 10176 24312 10218 24346
rect 10252 24312 10294 24346
rect 10328 24312 10369 24346
rect 10403 24312 10444 24346
rect 10478 24312 10519 24346
rect 10553 24312 10594 24346
rect 10628 24312 10669 24346
rect 10703 24312 10744 24346
rect 10778 24312 10819 24346
rect 10853 24312 10894 24346
rect 10928 24312 10969 24346
rect 11003 24312 11044 24346
rect 11078 24312 11119 24346
rect 11153 24312 11194 24346
rect 11228 24312 11240 24346
rect 9901 24274 11240 24312
rect 9901 24240 9914 24274
rect 9948 24240 9990 24274
rect 10024 24240 10066 24274
rect 10100 24240 10142 24274
rect 10176 24240 10218 24274
rect 10252 24240 10294 24274
rect 10328 24240 10369 24274
rect 10403 24240 10444 24274
rect 10478 24240 10519 24274
rect 10553 24240 10594 24274
rect 10628 24240 10669 24274
rect 10703 24240 10744 24274
rect 10778 24240 10819 24274
rect 10853 24240 10894 24274
rect 10928 24240 10969 24274
rect 11003 24240 11044 24274
rect 11078 24240 11119 24274
rect 11153 24240 11194 24274
rect 11228 24240 11240 24274
tri 9899 24229 9901 24231 se
rect 9901 24229 11240 24240
rect 14053 24657 14403 24696
rect 14053 24623 14252 24657
rect 14286 24623 14324 24657
rect 14358 24623 14403 24657
rect 14053 24584 14403 24623
rect 14053 24550 14252 24584
rect 14286 24550 14324 24584
rect 14358 24550 14403 24584
rect 14053 24511 14403 24550
rect 14053 24477 14252 24511
rect 14286 24477 14324 24511
rect 14358 24477 14403 24511
rect 14053 24438 14403 24477
rect 14053 24404 14252 24438
rect 14286 24404 14324 24438
rect 14358 24404 14403 24438
rect 14053 24365 14403 24404
rect 14053 24331 14252 24365
rect 14286 24331 14324 24365
rect 14358 24331 14403 24365
rect 14053 24292 14403 24331
rect 14053 24258 14252 24292
rect 14286 24258 14324 24292
rect 14358 24258 14403 24292
tri 9896 24226 9899 24229 se
rect 9899 24226 11086 24229
tri 11086 24226 11089 24229 nw
rect 9896 24219 11079 24226
tri 11079 24219 11086 24226 nw
rect 14053 24219 14403 24258
rect 9896 24185 11045 24219
tri 11045 24185 11079 24219 nw
rect 14053 24185 14252 24219
rect 14286 24185 14324 24219
rect 14358 24185 14403 24219
rect 9896 24171 11006 24185
rect 9896 24137 9905 24171
rect 9939 24137 9981 24171
rect 10015 24137 10057 24171
rect 10091 24137 10133 24171
rect 10167 24137 10209 24171
rect 10243 24137 10285 24171
rect 10319 24137 10361 24171
rect 10395 24137 10437 24171
rect 10471 24137 10513 24171
rect 10547 24137 10589 24171
rect 10623 24137 10665 24171
rect 10699 24146 11006 24171
tri 11006 24146 11045 24185 nw
rect 14053 24146 14403 24185
rect 10699 24137 10972 24146
rect 9896 24112 10972 24137
tri 10972 24112 11006 24146 nw
rect 14053 24112 14252 24146
rect 14286 24112 14324 24146
rect 14358 24112 14403 24146
rect 9896 24097 10933 24112
rect 9896 24063 9905 24097
rect 9939 24063 9981 24097
rect 10015 24063 10057 24097
rect 10091 24063 10133 24097
rect 10167 24063 10209 24097
rect 10243 24063 10285 24097
rect 10319 24063 10361 24097
rect 10395 24063 10437 24097
rect 10471 24063 10513 24097
rect 10547 24063 10589 24097
rect 10623 24063 10665 24097
rect 10699 24073 10933 24097
tri 10933 24073 10972 24112 nw
rect 14053 24073 14403 24112
rect 10699 24063 10899 24073
rect 9896 24039 10899 24063
tri 10899 24039 10933 24073 nw
rect 14053 24039 14252 24073
rect 14286 24039 14324 24073
rect 14358 24039 14403 24073
rect 9896 24023 10860 24039
rect 9896 23989 9905 24023
rect 9939 23989 9981 24023
rect 10015 23989 10057 24023
rect 10091 23989 10133 24023
rect 10167 23989 10209 24023
rect 10243 23989 10285 24023
rect 10319 23989 10361 24023
rect 10395 23989 10437 24023
rect 10471 23989 10513 24023
rect 10547 23989 10589 24023
rect 10623 23989 10665 24023
rect 10699 24000 10860 24023
tri 10860 24000 10899 24039 nw
rect 14053 24000 14403 24039
rect 10699 23989 10826 24000
rect 9896 23966 10826 23989
tri 10826 23966 10860 24000 nw
rect 14053 23966 14252 24000
rect 14286 23966 14324 24000
rect 14358 23966 14403 24000
rect 9896 23949 10787 23966
rect 9896 23915 9905 23949
rect 9939 23915 9981 23949
rect 10015 23915 10057 23949
rect 10091 23915 10133 23949
rect 10167 23915 10209 23949
rect 10243 23915 10285 23949
rect 10319 23915 10361 23949
rect 10395 23915 10437 23949
rect 10471 23915 10513 23949
rect 10547 23915 10589 23949
rect 10623 23915 10665 23949
rect 10699 23927 10787 23949
tri 10787 23927 10826 23966 nw
rect 14053 23927 14403 23966
rect 10699 23915 10753 23927
rect 9896 23893 10753 23915
tri 10753 23893 10787 23927 nw
rect 14053 23893 14252 23927
rect 14286 23893 14324 23927
rect 14358 23893 14403 23927
rect 9896 23875 10714 23893
rect 9896 23841 9905 23875
rect 9939 23841 9981 23875
rect 10015 23841 10057 23875
rect 10091 23841 10133 23875
rect 10167 23841 10209 23875
rect 10243 23841 10285 23875
rect 10319 23841 10361 23875
rect 10395 23841 10437 23875
rect 10471 23841 10513 23875
rect 10547 23841 10589 23875
rect 10623 23841 10665 23875
rect 10699 23854 10714 23875
tri 10714 23854 10753 23893 nw
rect 14053 23886 14403 23893
tri 14053 23877 14062 23886 nw
rect 14062 23854 14403 23886
rect 10699 23841 10708 23854
tri 10708 23848 10714 23854 nw
rect 9896 23801 10708 23841
rect 9896 23767 9905 23801
rect 9939 23767 9981 23801
rect 10015 23767 10057 23801
rect 10091 23767 10133 23801
rect 10167 23767 10209 23801
rect 10243 23767 10285 23801
rect 10319 23767 10361 23801
rect 10395 23767 10437 23801
rect 10471 23767 10513 23801
rect 10547 23767 10589 23801
rect 10623 23767 10665 23801
rect 10699 23767 10708 23801
rect 9896 23727 10708 23767
rect 9896 23693 9905 23727
rect 9939 23693 9981 23727
rect 10015 23693 10057 23727
rect 10091 23693 10133 23727
rect 10167 23693 10209 23727
rect 10243 23693 10285 23727
rect 10319 23693 10361 23727
rect 10395 23693 10437 23727
rect 10471 23693 10513 23727
rect 10547 23693 10589 23727
rect 10623 23693 10665 23727
rect 10699 23693 10708 23727
rect 9896 23653 10708 23693
rect 9896 23619 9905 23653
rect 9939 23619 9981 23653
rect 10015 23619 10057 23653
rect 10091 23619 10133 23653
rect 10167 23619 10209 23653
rect 10243 23619 10285 23653
rect 10319 23619 10361 23653
rect 10395 23619 10437 23653
rect 10471 23619 10513 23653
rect 10547 23619 10589 23653
rect 10623 23619 10665 23653
rect 10699 23619 10708 23653
rect 9896 23579 10708 23619
rect 9896 23545 9905 23579
rect 9939 23545 9981 23579
rect 10015 23545 10057 23579
rect 10091 23545 10133 23579
rect 10167 23545 10209 23579
rect 10243 23545 10285 23579
rect 10319 23545 10361 23579
rect 10395 23545 10437 23579
rect 10471 23545 10513 23579
rect 10547 23545 10589 23579
rect 10623 23545 10665 23579
rect 10699 23545 10708 23579
rect 9896 23505 10708 23545
rect 9896 23471 9905 23505
rect 9939 23471 9981 23505
rect 10015 23471 10057 23505
rect 10091 23471 10133 23505
rect 10167 23471 10209 23505
rect 10243 23471 10285 23505
rect 10319 23471 10361 23505
rect 10395 23471 10437 23505
rect 10471 23471 10513 23505
rect 10547 23471 10589 23505
rect 10623 23471 10665 23505
rect 10699 23471 10708 23505
rect 9896 23431 10708 23471
rect 9896 23397 9905 23431
rect 9939 23397 9981 23431
rect 10015 23397 10057 23431
rect 10091 23397 10133 23431
rect 10167 23397 10209 23431
rect 10243 23397 10285 23431
rect 10319 23397 10361 23431
rect 10395 23397 10437 23431
rect 10471 23397 10513 23431
rect 10547 23397 10589 23431
rect 10623 23397 10665 23431
rect 10699 23397 10708 23431
rect 9896 23357 10708 23397
rect 9896 23323 9905 23357
rect 9939 23323 9981 23357
rect 10015 23323 10057 23357
rect 10091 23323 10133 23357
rect 10167 23323 10209 23357
rect 10243 23323 10285 23357
rect 10319 23323 10361 23357
rect 10395 23323 10437 23357
rect 10471 23323 10513 23357
rect 10547 23323 10589 23357
rect 10623 23323 10665 23357
rect 10699 23323 10708 23357
rect 9896 23283 10708 23323
rect 9896 23249 9905 23283
rect 9939 23249 9981 23283
rect 10015 23249 10057 23283
rect 10091 23249 10133 23283
rect 10167 23249 10209 23283
rect 10243 23249 10285 23283
rect 10319 23249 10361 23283
rect 10395 23249 10437 23283
rect 10471 23249 10513 23283
rect 10547 23249 10589 23283
rect 10623 23249 10665 23283
rect 10699 23249 10708 23283
rect 9896 23209 10708 23249
rect 14062 23820 14252 23854
rect 14286 23820 14324 23854
rect 14358 23820 14403 23854
rect 14062 23781 14403 23820
rect 14062 23747 14252 23781
rect 14286 23747 14324 23781
rect 14358 23747 14403 23781
rect 14062 23708 14403 23747
rect 14062 23674 14252 23708
rect 14286 23674 14324 23708
rect 14358 23674 14403 23708
rect 14062 23635 14403 23674
rect 14062 23601 14252 23635
rect 14286 23601 14324 23635
rect 14358 23601 14403 23635
rect 14062 23562 14403 23601
rect 14062 23528 14252 23562
rect 14286 23528 14324 23562
rect 14358 23528 14403 23562
rect 14062 23489 14403 23528
rect 14062 23455 14252 23489
rect 14286 23455 14324 23489
rect 14358 23455 14403 23489
rect 14062 23416 14403 23455
rect 14062 23382 14252 23416
rect 14286 23382 14324 23416
rect 14358 23382 14403 23416
rect 14062 23343 14403 23382
rect 14062 23309 14252 23343
rect 14286 23309 14324 23343
rect 14358 23309 14403 23343
rect 14062 23270 14403 23309
rect 14062 23236 14252 23270
rect 14286 23236 14324 23270
rect 14358 23236 14403 23270
rect 9896 23175 9905 23209
rect 9939 23175 9981 23209
rect 10015 23175 10057 23209
rect 10091 23175 10133 23209
rect 10167 23175 10209 23209
rect 10243 23175 10285 23209
rect 10319 23175 10361 23209
rect 10395 23175 10437 23209
rect 10471 23175 10513 23209
rect 10547 23175 10589 23209
rect 10623 23175 10665 23209
rect 10699 23197 10708 23209
tri 10708 23197 10743 23232 sw
rect 14062 23197 14403 23236
rect 10699 23175 10743 23197
rect 9896 23163 10743 23175
tri 10743 23163 10777 23197 sw
rect 14062 23163 14252 23197
rect 14286 23163 14324 23197
rect 14358 23163 14403 23197
rect 9896 23135 10777 23163
rect 9896 23101 9905 23135
rect 9939 23101 9981 23135
rect 10015 23101 10057 23135
rect 10091 23101 10133 23135
rect 10167 23101 10209 23135
rect 10243 23101 10285 23135
rect 10319 23101 10361 23135
rect 10395 23101 10437 23135
rect 10471 23101 10513 23135
rect 10547 23101 10589 23135
rect 10623 23101 10665 23135
rect 10699 23124 10777 23135
tri 10777 23124 10816 23163 sw
tri 14051 23124 14062 23135 se
rect 14062 23124 14403 23163
rect 10699 23101 10816 23124
rect 9896 23090 10816 23101
tri 10816 23090 10850 23124 sw
tri 14017 23090 14051 23124 se
rect 14051 23090 14252 23124
rect 14286 23090 14324 23124
rect 14358 23090 14403 23124
rect 9896 23061 10850 23090
rect 9896 23027 9905 23061
rect 9939 23027 9981 23061
rect 10015 23027 10057 23061
rect 10091 23027 10133 23061
rect 10167 23027 10209 23061
rect 10243 23027 10285 23061
rect 10319 23027 10361 23061
rect 10395 23027 10437 23061
rect 10471 23027 10513 23061
rect 10547 23027 10589 23061
rect 10623 23027 10665 23061
rect 10699 23051 10850 23061
tri 10850 23051 10889 23090 sw
tri 13978 23051 14017 23090 se
rect 14017 23051 14403 23090
rect 10699 23027 10889 23051
rect 9896 23017 10889 23027
tri 10889 23017 10923 23051 sw
tri 13944 23017 13978 23051 se
rect 13978 23017 14252 23051
rect 14286 23017 14324 23051
rect 14358 23017 14403 23051
rect 9896 23011 10923 23017
tri 10923 23011 10929 23017 sw
tri 13938 23011 13944 23017 se
rect 13944 23011 14403 23017
rect 9896 23000 14403 23011
rect 9896 22987 10759 23000
rect 9896 22953 9905 22987
rect 9939 22953 9981 22987
rect 10015 22953 10057 22987
rect 10091 22953 10133 22987
rect 10167 22953 10209 22987
rect 10243 22953 10285 22987
rect 10319 22953 10361 22987
rect 10395 22953 10437 22987
rect 10471 22953 10513 22987
rect 10547 22953 10589 22987
rect 10623 22953 10665 22987
rect 10699 22966 10759 22987
rect 10793 22966 10832 23000
rect 10866 22966 10905 23000
rect 10939 22966 10978 23000
rect 11012 22966 11051 23000
rect 11085 22966 11124 23000
rect 11158 22966 11197 23000
rect 11231 22966 11270 23000
rect 11304 22966 11343 23000
rect 11377 22966 11416 23000
rect 11450 22966 11489 23000
rect 11523 22966 11562 23000
rect 11596 22966 11635 23000
rect 11669 22966 11707 23000
rect 11741 22966 11779 23000
rect 11813 22966 11851 23000
rect 11885 22966 11923 23000
rect 11957 22966 11995 23000
rect 12029 22966 12067 23000
rect 12101 22966 12139 23000
rect 12173 22966 12211 23000
rect 12245 22999 14403 23000
rect 12245 22984 13756 22999
rect 12245 22966 12476 22984
rect 10699 22953 12476 22966
rect 9896 22950 12476 22953
rect 12510 22950 12550 22984
rect 12584 22950 12624 22984
rect 12658 22950 12698 22984
rect 12732 22950 12772 22984
rect 12806 22950 12846 22984
rect 12880 22950 12920 22984
rect 12954 22950 12994 22984
rect 13028 22950 13068 22984
rect 13102 22950 13141 22984
rect 13175 22950 13214 22984
rect 13248 22950 13287 22984
rect 13321 22950 13360 22984
rect 13394 22950 13433 22984
rect 13467 22950 13506 22984
rect 13540 22950 13579 22984
rect 13613 22950 13652 22984
rect 13686 22965 13756 22984
rect 13790 22965 13828 22999
rect 13862 22965 13900 22999
rect 13934 22965 13972 22999
rect 14006 22965 14044 22999
rect 14078 22965 14116 22999
rect 14150 22978 14403 22999
rect 14150 22965 14252 22978
rect 13686 22950 14252 22965
rect 9896 22944 14252 22950
rect 14286 22944 14324 22978
rect 14358 22944 14403 22978
rect 9896 22925 14403 22944
rect 9896 22923 13756 22925
rect 9896 22914 12322 22923
rect 9896 22913 10759 22914
rect 9896 22879 9905 22913
rect 9939 22879 9981 22913
rect 10015 22879 10057 22913
rect 10091 22879 10133 22913
rect 10167 22879 10209 22913
rect 10243 22879 10285 22913
rect 10319 22879 10361 22913
rect 10395 22879 10437 22913
rect 10471 22879 10513 22913
rect 10547 22879 10589 22913
rect 10623 22879 10665 22913
rect 10699 22880 10759 22913
rect 10793 22880 10832 22914
rect 10866 22880 10905 22914
rect 10939 22880 10978 22914
rect 11012 22880 11051 22914
rect 11085 22880 11124 22914
rect 11158 22880 11197 22914
rect 11231 22880 11270 22914
rect 11304 22880 11343 22914
rect 11377 22880 11416 22914
rect 11450 22880 11489 22914
rect 11523 22880 11562 22914
rect 11596 22880 11635 22914
rect 11669 22880 11707 22914
rect 11741 22880 11779 22914
rect 11813 22880 11851 22914
rect 11885 22880 11923 22914
rect 11957 22880 11995 22914
rect 12029 22880 12067 22914
rect 12101 22880 12139 22914
rect 12173 22880 12211 22914
rect 12245 22891 12322 22914
tri 12322 22891 12354 22923 nw
tri 13599 22891 13631 22923 ne
rect 13631 22891 13756 22923
rect 13790 22891 13828 22925
rect 13862 22891 13900 22925
rect 13934 22891 13972 22925
rect 14006 22891 14044 22925
rect 14078 22891 14116 22925
rect 14150 22905 14403 22925
rect 14150 22891 14252 22905
rect 12245 22880 12302 22891
rect 10699 22879 12302 22880
rect 9896 22871 12302 22879
tri 12302 22871 12322 22891 nw
tri 13631 22871 13651 22891 ne
rect 13651 22871 14252 22891
rect 14286 22871 14324 22905
rect 14358 22871 14403 22905
rect 9896 22851 12282 22871
tri 12282 22851 12302 22871 nw
tri 13651 22851 13671 22871 ne
rect 13671 22851 14403 22871
rect 9896 22839 12257 22851
rect 9896 22805 9905 22839
rect 9939 22805 9981 22839
rect 10015 22805 10057 22839
rect 10091 22805 10133 22839
rect 10167 22805 10209 22839
rect 10243 22805 10285 22839
rect 10319 22805 10361 22839
rect 10395 22805 10437 22839
rect 10471 22805 10513 22839
rect 10547 22805 10589 22839
rect 10623 22805 10665 22839
rect 10699 22828 12257 22839
rect 10699 22805 10759 22828
rect 9896 22794 10759 22805
rect 10793 22794 10832 22828
rect 10866 22794 10905 22828
rect 10939 22794 10978 22828
rect 11012 22794 11051 22828
rect 11085 22794 11124 22828
rect 11158 22794 11197 22828
rect 11231 22794 11270 22828
rect 11304 22794 11343 22828
rect 11377 22794 11416 22828
rect 11450 22794 11489 22828
rect 11523 22794 11562 22828
rect 11596 22794 11635 22828
rect 11669 22794 11707 22828
rect 11741 22794 11779 22828
rect 11813 22794 11851 22828
rect 11885 22794 11923 22828
rect 11957 22794 11995 22828
rect 12029 22794 12067 22828
rect 12101 22794 12139 22828
rect 12173 22794 12211 22828
rect 12245 22794 12257 22828
tri 12257 22826 12282 22851 nw
tri 13671 22826 13696 22851 ne
rect 13696 22826 13756 22851
tri 13696 22817 13705 22826 ne
rect 13705 22817 13756 22826
rect 13790 22817 13828 22851
rect 13862 22817 13900 22851
rect 13934 22817 13972 22851
rect 14006 22817 14044 22851
rect 14078 22817 14116 22851
rect 14150 22832 14403 22851
rect 14150 22817 14252 22832
tri 13705 22809 13713 22817 ne
rect 9896 22765 12257 22794
rect 9896 22731 9905 22765
rect 9939 22731 9981 22765
rect 10015 22731 10057 22765
rect 10091 22731 10133 22765
rect 10167 22731 10209 22765
rect 10243 22731 10285 22765
rect 10319 22731 10361 22765
rect 10395 22731 10437 22765
rect 10471 22731 10513 22765
rect 10547 22731 10589 22765
rect 10623 22731 10665 22765
rect 10699 22742 12257 22765
rect 10699 22731 10759 22742
rect 9896 22708 10759 22731
rect 10793 22708 10832 22742
rect 10866 22708 10905 22742
rect 10939 22708 10978 22742
rect 11012 22708 11051 22742
rect 11085 22708 11124 22742
rect 11158 22708 11197 22742
rect 11231 22708 11270 22742
rect 11304 22708 11343 22742
rect 11377 22708 11416 22742
rect 11450 22708 11489 22742
rect 11523 22708 11562 22742
rect 11596 22708 11635 22742
rect 11669 22708 11707 22742
rect 11741 22708 11779 22742
rect 11813 22708 11851 22742
rect 11885 22708 11923 22742
rect 11957 22708 11995 22742
rect 12029 22708 12067 22742
rect 12101 22708 12139 22742
rect 12173 22708 12211 22742
rect 12245 22708 12257 22742
rect 9896 22691 12257 22708
rect 9896 22657 9905 22691
rect 9939 22657 9981 22691
rect 10015 22657 10057 22691
rect 10091 22657 10133 22691
rect 10167 22657 10209 22691
rect 10243 22657 10285 22691
rect 10319 22657 10361 22691
rect 10395 22657 10437 22691
rect 10471 22657 10513 22691
rect 10547 22657 10589 22691
rect 10623 22657 10665 22691
rect 10699 22657 12257 22691
rect 9896 22656 12257 22657
rect 9896 22622 10759 22656
rect 10793 22622 10832 22656
rect 10866 22622 10905 22656
rect 10939 22622 10978 22656
rect 11012 22622 11051 22656
rect 11085 22622 11124 22656
rect 11158 22622 11197 22656
rect 11231 22622 11270 22656
rect 11304 22622 11343 22656
rect 11377 22622 11416 22656
rect 11450 22622 11489 22656
rect 11523 22622 11562 22656
rect 11596 22622 11635 22656
rect 11669 22622 11707 22656
rect 11741 22622 11779 22656
rect 11813 22622 11851 22656
rect 11885 22622 11923 22656
rect 11957 22622 11995 22656
rect 12029 22622 12067 22656
rect 12101 22622 12139 22656
rect 12173 22622 12211 22656
rect 12245 22622 12257 22656
rect 9896 22617 12257 22622
rect 9896 22583 9905 22617
rect 9939 22583 9981 22617
rect 10015 22583 10057 22617
rect 10091 22583 10133 22617
rect 10167 22583 10209 22617
rect 10243 22583 10285 22617
rect 10319 22583 10361 22617
rect 10395 22583 10437 22617
rect 10471 22583 10513 22617
rect 10547 22583 10589 22617
rect 10623 22583 10665 22617
rect 10699 22614 12257 22617
rect 13713 22798 14252 22817
rect 14286 22798 14324 22832
rect 14358 22798 14403 22832
rect 13713 22777 14403 22798
rect 13713 22743 13756 22777
rect 13790 22743 13828 22777
rect 13862 22743 13900 22777
rect 13934 22743 13972 22777
rect 14006 22743 14044 22777
rect 14078 22743 14116 22777
rect 14150 22759 14403 22777
rect 14150 22743 14252 22759
rect 13713 22725 14252 22743
rect 14286 22725 14324 22759
rect 14358 22725 14403 22759
rect 13713 22703 14403 22725
rect 13713 22669 13756 22703
rect 13790 22669 13828 22703
rect 13862 22669 13900 22703
rect 13934 22669 13972 22703
rect 14006 22669 14044 22703
rect 14078 22669 14116 22703
rect 14150 22686 14403 22703
rect 14150 22669 14252 22686
rect 13713 22652 14252 22669
rect 14286 22652 14324 22686
rect 14358 22652 14403 22686
rect 13713 22629 14403 22652
rect 10699 22595 10732 22614
tri 10732 22595 10751 22614 nw
rect 13713 22595 13756 22629
rect 13790 22595 13828 22629
rect 13862 22595 13900 22629
rect 13934 22595 13972 22629
rect 14006 22595 14044 22629
rect 14078 22595 14116 22629
rect 14150 22613 14403 22629
rect 14150 22595 14252 22613
rect 10699 22583 10716 22595
rect 9896 22579 10716 22583
tri 10716 22579 10732 22595 nw
rect 13713 22579 14252 22595
rect 14286 22579 14324 22613
rect 14358 22579 14403 22613
rect 9896 22571 10708 22579
tri 10708 22571 10716 22579 nw
rect 13713 22555 14403 22579
rect 13713 22521 13756 22555
rect 13790 22521 13828 22555
rect 13862 22521 13900 22555
rect 13934 22521 13972 22555
rect 14006 22521 14044 22555
rect 14078 22521 14116 22555
rect 14150 22540 14403 22555
rect 14150 22521 14252 22540
rect 13713 22506 14252 22521
rect 14286 22506 14324 22540
rect 14358 22506 14403 22540
rect 13713 22481 14403 22506
rect 13713 22447 13756 22481
rect 13790 22447 13828 22481
rect 13862 22447 13900 22481
rect 13934 22447 13972 22481
rect 14006 22447 14044 22481
rect 14078 22447 14116 22481
rect 14150 22467 14403 22481
rect 14150 22447 14252 22467
rect 13713 22433 14252 22447
rect 14286 22433 14324 22467
rect 14358 22433 14403 22467
rect 13713 22407 14403 22433
rect 13713 22373 13756 22407
rect 13790 22373 13828 22407
rect 13862 22373 13900 22407
rect 13934 22373 13972 22407
rect 14006 22373 14044 22407
rect 14078 22373 14116 22407
rect 14150 22394 14403 22407
rect 14150 22373 14252 22394
rect 13713 22360 14252 22373
rect 14286 22360 14324 22394
rect 14358 22360 14403 22394
rect 13713 22333 14403 22360
rect 13713 22299 13756 22333
rect 13790 22299 13828 22333
rect 13862 22299 13900 22333
rect 13934 22299 13972 22333
rect 14006 22299 14044 22333
rect 14078 22299 14116 22333
rect 14150 22321 14403 22333
rect 14150 22299 14252 22321
rect 13713 22287 14252 22299
rect 14286 22287 14324 22321
rect 14358 22287 14403 22321
rect 13713 22259 14403 22287
rect 13713 22225 13756 22259
rect 13790 22225 13828 22259
rect 13862 22225 13900 22259
rect 13934 22225 13972 22259
rect 14006 22225 14044 22259
rect 14078 22225 14116 22259
rect 14150 22248 14403 22259
rect 14150 22225 14252 22248
rect 13713 22214 14252 22225
rect 14286 22214 14324 22248
rect 14358 22214 14403 22248
rect 13713 22185 14403 22214
rect 13713 22151 13756 22185
rect 13790 22151 13828 22185
rect 13862 22151 13900 22185
rect 13934 22151 13972 22185
rect 14006 22151 14044 22185
rect 14078 22151 14116 22185
rect 14150 22175 14403 22185
rect 14150 22151 14252 22175
rect 13713 22141 14252 22151
rect 14286 22141 14324 22175
rect 14358 22141 14403 22175
rect 13713 22111 14403 22141
rect 5390 22104 7582 22110
rect 5506 21994 7582 22104
rect 7698 21994 7704 22110
rect 5506 21988 7704 21994
rect 5390 21982 7704 21988
rect 13713 22077 13756 22111
rect 13790 22077 13828 22111
rect 13862 22077 13900 22111
rect 13934 22077 13972 22111
rect 14006 22077 14044 22111
rect 14078 22077 14116 22111
rect 14150 22102 14403 22111
rect 14150 22077 14252 22102
rect 13713 22068 14252 22077
rect 14286 22068 14324 22102
rect 14358 22068 14403 22102
rect 13713 22037 14403 22068
rect 13713 22003 13756 22037
rect 13790 22003 13828 22037
rect 13862 22003 13900 22037
rect 13934 22003 13972 22037
rect 14006 22003 14044 22037
rect 14078 22003 14116 22037
rect 14150 22029 14403 22037
rect 14150 22003 14252 22029
rect 13713 21995 14252 22003
rect 14286 21995 14324 22029
rect 14358 21995 14403 22029
rect 13713 21963 14403 21995
rect 4973 21919 7940 21954
rect 4973 21916 7760 21919
rect 5089 21803 7760 21916
rect 5089 21800 7940 21803
rect 4973 21774 7940 21800
rect 13713 21929 13756 21963
rect 13790 21929 13828 21963
rect 13862 21929 13900 21963
rect 13934 21929 13972 21963
rect 14006 21929 14044 21963
rect 14078 21929 14116 21963
rect 14150 21956 14403 21963
rect 14150 21929 14252 21956
rect 13713 21922 14252 21929
rect 14286 21922 14324 21956
rect 14358 21922 14403 21956
rect 13713 21889 14403 21922
rect 13713 21855 13756 21889
rect 13790 21855 13828 21889
rect 13862 21855 13900 21889
rect 13934 21855 13972 21889
rect 14006 21855 14044 21889
rect 14078 21855 14116 21889
rect 14150 21883 14403 21889
rect 14150 21855 14252 21883
rect 13713 21849 14252 21855
rect 14286 21849 14324 21883
rect 14358 21849 14403 21883
rect 13713 21815 14403 21849
rect 13713 21781 13756 21815
rect 13790 21781 13828 21815
rect 13862 21781 13900 21815
rect 13934 21781 13972 21815
rect 14006 21781 14044 21815
rect 14078 21781 14116 21815
rect 14150 21810 14403 21815
rect 14150 21781 14252 21810
rect 13713 21776 14252 21781
rect 14286 21776 14324 21810
rect 14358 21776 14403 21810
rect 13713 21741 14403 21776
rect 6819 21711 7067 21717
rect 6819 21659 6821 21711
rect 6873 21659 6885 21711
rect 6937 21659 6949 21711
rect 7001 21659 7013 21711
rect 7065 21659 7067 21711
rect 6819 21645 7067 21659
rect 6819 21593 6821 21645
rect 6873 21593 6885 21645
rect 6937 21593 6949 21645
rect 7001 21593 7013 21645
rect 7065 21593 7067 21645
rect 6819 21579 7067 21593
rect 6819 21527 6821 21579
rect 6873 21527 6885 21579
rect 6937 21527 6949 21579
rect 7001 21527 7013 21579
rect 7065 21527 7067 21579
rect 6819 21513 7067 21527
rect 6819 21461 6821 21513
rect 6873 21461 6885 21513
rect 6937 21461 6949 21513
rect 7001 21461 7013 21513
rect 7065 21461 7067 21513
rect 6819 21447 7067 21461
rect 6819 21395 6821 21447
rect 6873 21395 6885 21447
rect 6937 21395 6949 21447
rect 7001 21395 7013 21447
rect 7065 21395 7067 21447
rect 6819 21389 7067 21395
rect 13713 21707 13756 21741
rect 13790 21707 13828 21741
rect 13862 21707 13900 21741
rect 13934 21707 13972 21741
rect 14006 21707 14044 21741
rect 14078 21707 14116 21741
rect 14150 21737 14403 21741
rect 14150 21707 14252 21737
rect 13713 21703 14252 21707
rect 14286 21703 14324 21737
rect 14358 21703 14403 21737
rect 13713 21666 14403 21703
rect 13713 21632 13756 21666
rect 13790 21632 13828 21666
rect 13862 21632 13900 21666
rect 13934 21632 13972 21666
rect 14006 21632 14044 21666
rect 14078 21632 14116 21666
rect 14150 21664 14403 21666
rect 14150 21632 14252 21664
rect 13713 21630 14252 21632
rect 14286 21630 14324 21664
rect 14358 21630 14403 21664
rect 13713 21591 14403 21630
rect 13713 21557 13756 21591
rect 13790 21557 13828 21591
rect 13862 21557 13900 21591
rect 13934 21557 13972 21591
rect 14006 21557 14044 21591
rect 14078 21557 14116 21591
rect 14150 21557 14252 21591
rect 14286 21557 14324 21591
rect 14358 21557 14403 21591
rect 13713 21518 14403 21557
rect 13713 21516 14252 21518
rect 13713 21482 13756 21516
rect 13790 21482 13828 21516
rect 13862 21482 13900 21516
rect 13934 21482 13972 21516
rect 14006 21482 14044 21516
rect 14078 21482 14116 21516
rect 14150 21484 14252 21516
rect 14286 21484 14324 21518
rect 14358 21484 14403 21518
rect 14150 21482 14403 21484
rect 13713 21445 14403 21482
rect 13713 21441 14252 21445
rect 13713 21407 13756 21441
rect 13790 21407 13828 21441
rect 13862 21407 13900 21441
rect 13934 21407 13972 21441
rect 14006 21407 14044 21441
rect 14078 21407 14116 21441
rect 14150 21411 14252 21441
rect 14286 21411 14324 21445
rect 14358 21411 14403 21445
rect 14150 21407 14403 21411
rect 13713 21371 14403 21407
rect 13713 21366 14252 21371
rect 13713 21332 13756 21366
rect 13790 21332 13828 21366
rect 13862 21332 13900 21366
rect 13934 21332 13972 21366
rect 14006 21332 14044 21366
rect 14078 21332 14116 21366
rect 14150 21337 14252 21366
rect 14286 21337 14324 21371
rect 14358 21337 14403 21371
rect 14150 21332 14403 21337
rect 13713 21297 14403 21332
rect 13713 21291 14252 21297
rect 13713 21257 13756 21291
rect 13790 21257 13828 21291
rect 13862 21257 13900 21291
rect 13934 21257 13972 21291
rect 14006 21257 14044 21291
rect 14078 21257 14116 21291
rect 14150 21263 14252 21291
rect 14286 21263 14324 21297
rect 14358 21263 14403 21297
rect 14150 21257 14403 21263
rect 13713 21223 14403 21257
rect 13713 21216 14252 21223
rect 13713 21182 13756 21216
rect 13790 21182 13828 21216
rect 13862 21182 13900 21216
rect 13934 21182 13972 21216
rect 14006 21182 14044 21216
rect 14078 21182 14116 21216
rect 14150 21189 14252 21216
rect 14286 21189 14324 21223
rect 14358 21189 14403 21223
rect 14150 21182 14403 21189
tri 13680 21149 13713 21182 se
rect 13713 21149 14403 21182
tri 13672 21141 13680 21149 se
rect 13680 21141 14252 21149
tri 13638 21107 13672 21141 se
rect 13672 21107 13756 21141
rect 13790 21107 13828 21141
rect 13862 21107 13900 21141
rect 13934 21107 13972 21141
rect 14006 21107 14044 21141
rect 14078 21107 14116 21141
rect 14150 21115 14252 21141
rect 14286 21115 14324 21149
rect 14358 21115 14403 21149
rect 14150 21107 14403 21115
tri 13606 21075 13638 21107 se
rect 13638 21075 14403 21107
tri 13597 21066 13606 21075 se
rect 13606 21066 14252 21075
tri 13563 21032 13597 21066 se
rect 13597 21032 13756 21066
rect 13790 21032 13828 21066
rect 13862 21032 13900 21066
rect 13934 21032 13972 21066
rect 14006 21032 14044 21066
rect 14078 21032 14116 21066
rect 14150 21041 14252 21066
rect 14286 21041 14324 21075
rect 14358 21041 14403 21075
rect 14150 21032 14403 21041
tri 13529 20998 13563 21032 se
rect 13563 20998 14403 21032
rect 13529 20952 14403 20998
tri 14285 20916 14321 20952 ne
rect 14321 20916 14367 20952
tri 14367 20916 14403 20952 nw
rect 3003 20732 3009 20848
rect 3189 20732 3195 20848
rect 4518 20732 4524 20848
rect 4640 20732 4646 20848
rect 729 19976 735 20028
rect 787 19976 799 20028
rect 851 19976 4884 20028
rect 4936 19976 4948 20028
rect 5000 19976 5006 20028
rect 729 19868 735 19920
rect 787 19868 799 19920
rect 851 19868 4884 19920
rect 4936 19868 4948 19920
rect 5000 19868 5006 19920
rect 9399 19423 9477 19429
rect 9399 19371 9412 19423
rect 9464 19371 9477 19423
rect 9399 19359 9477 19371
rect 9399 19307 9412 19359
rect 9464 19307 9477 19359
rect 9399 19295 9477 19307
rect 9399 19243 9412 19295
rect 9464 19243 9477 19295
rect 9399 19231 9477 19243
rect 9399 19179 9412 19231
rect 9464 19179 9477 19231
rect 9399 19167 9477 19179
rect 9399 19115 9412 19167
rect 9464 19115 9477 19167
rect 9399 19103 9477 19115
rect 9399 19051 9412 19103
rect 9464 19051 9477 19103
rect 9399 19039 9477 19051
rect 9399 18987 9412 19039
rect 9464 18987 9477 19039
rect 9399 18975 9477 18987
rect 9399 18923 9412 18975
rect 9464 18923 9477 18975
rect 9399 18911 9477 18923
rect 9399 18859 9412 18911
rect 9464 18859 9477 18911
rect 9399 18847 9477 18859
rect 9399 18795 9412 18847
rect 9464 18795 9477 18847
rect 9399 18783 9477 18795
rect 9399 18731 9412 18783
rect 9464 18731 9477 18783
rect 9399 18719 9477 18731
rect 9399 18667 9412 18719
rect 9464 18667 9477 18719
rect 9399 18655 9477 18667
rect 9399 18603 9412 18655
rect 9464 18603 9477 18655
rect 9399 18591 9477 18603
rect 6652 18500 6658 18552
rect 6710 18500 6716 18552
rect 6652 18488 6716 18500
rect 6652 18436 6658 18488
rect 6710 18436 6716 18488
rect 6652 18424 6716 18436
rect 6652 18372 6658 18424
rect 6710 18372 6716 18424
rect 6652 18360 6716 18372
rect 6652 18308 6658 18360
rect 6710 18308 6716 18360
rect 9399 18539 9412 18591
rect 9464 18539 9477 18591
rect 9399 18527 9477 18539
rect 9399 18475 9412 18527
rect 9464 18475 9477 18527
rect 9399 18463 9477 18475
rect 9399 18411 9412 18463
rect 9464 18411 9477 18463
rect 9706 19423 9902 19429
rect 9706 19371 9714 19423
rect 9766 19371 9778 19423
rect 9830 19371 9842 19423
rect 9894 19371 9902 19423
rect 9706 19358 9902 19371
rect 9706 19306 9714 19358
rect 9766 19306 9778 19358
rect 9830 19306 9842 19358
rect 9894 19306 9902 19358
rect 9706 19293 9902 19306
rect 9706 19241 9714 19293
rect 9766 19241 9778 19293
rect 9830 19241 9842 19293
rect 9894 19241 9902 19293
rect 9706 19228 9902 19241
rect 9706 19176 9714 19228
rect 9766 19176 9778 19228
rect 9830 19176 9842 19228
rect 9894 19176 9902 19228
rect 9706 19163 9902 19176
rect 9706 19111 9714 19163
rect 9766 19111 9778 19163
rect 9830 19111 9842 19163
rect 9894 19111 9902 19163
rect 9706 19098 9902 19111
rect 9706 19046 9714 19098
rect 9766 19046 9778 19098
rect 9830 19046 9842 19098
rect 9894 19046 9902 19098
rect 9706 19033 9902 19046
rect 9706 18981 9714 19033
rect 9766 18981 9778 19033
rect 9830 18981 9842 19033
rect 9894 18981 9902 19033
rect 9706 18968 9902 18981
rect 9706 18916 9714 18968
rect 9766 18916 9778 18968
rect 9830 18916 9842 18968
rect 9894 18916 9902 18968
rect 9706 18903 9902 18916
rect 9706 18851 9714 18903
rect 9766 18851 9778 18903
rect 9830 18851 9842 18903
rect 9894 18851 9902 18903
rect 9706 18837 9902 18851
rect 9706 18785 9714 18837
rect 9766 18785 9778 18837
rect 9830 18785 9842 18837
rect 9894 18785 9902 18837
rect 9706 18771 9902 18785
rect 9706 18719 9714 18771
rect 9766 18719 9778 18771
rect 9830 18719 9842 18771
rect 9894 18719 9902 18771
rect 9706 18705 9902 18719
rect 9706 18653 9714 18705
rect 9766 18653 9778 18705
rect 9830 18653 9842 18705
rect 9894 18653 9902 18705
rect 9706 18639 9902 18653
rect 9706 18587 9714 18639
rect 9766 18587 9778 18639
rect 9830 18587 9842 18639
rect 9894 18587 9902 18639
rect 9706 18573 9902 18587
rect 9706 18521 9714 18573
rect 9766 18521 9778 18573
rect 9830 18521 9842 18573
rect 9894 18521 9902 18573
rect 9706 18507 9902 18521
rect 9706 18455 9714 18507
rect 9766 18455 9778 18507
rect 9830 18455 9842 18507
rect 9894 18455 9902 18507
rect 9706 18449 9902 18455
rect 9399 18399 9477 18411
rect 9399 18347 9412 18399
rect 9464 18347 9477 18399
rect 9399 18334 9477 18347
rect 9399 18282 9412 18334
rect 9464 18282 9477 18334
rect 9399 18269 9477 18282
rect 9399 18217 9412 18269
rect 9464 18217 9477 18269
rect 9399 18204 9477 18217
rect 9399 18152 9412 18204
rect 9464 18152 9477 18204
rect 9399 18146 9477 18152
rect 3003 18024 3009 18140
rect 3189 18024 3195 18140
tri 14344 18107 14345 18108 se
rect 14345 18107 14388 18108
rect 5847 18088 5893 18107
tri 5893 18088 5912 18107 sw
tri 14325 18088 14344 18107 se
rect 14344 18088 14388 18107
rect 5847 18063 5912 18088
tri 5912 18063 5937 18088 sw
tri 13171 18063 13196 18088 se
rect 13196 18063 13242 18088
tri 13242 18063 13267 18088 sw
tri 14300 18063 14325 18088 se
rect 14325 18063 14388 18088
rect 5847 17939 14388 18063
rect 6652 17859 6658 17911
rect 6710 17859 6722 17911
rect 6774 17864 13697 17911
rect 6774 17859 6851 17864
tri 6851 17859 6856 17864 nw
tri 13686 17859 13691 17864 ne
rect 13691 17859 13697 17864
rect 13749 17859 13765 17911
rect 13817 17859 13823 17911
rect 14026 17864 14041 17911
tri 14026 17859 14031 17864 ne
rect 14031 17859 14041 17864
rect 14093 17859 14105 17911
rect 14157 17859 14170 17911
rect 6652 17851 6843 17859
tri 6843 17851 6851 17859 nw
tri 14031 17851 14039 17859 ne
rect 14039 17851 14170 17859
rect 5901 17784 5907 17836
rect 5959 17784 5971 17836
rect 6023 17823 6627 17836
tri 6627 17823 6640 17836 sw
tri 6859 17823 6872 17836 se
rect 6872 17823 13341 17836
rect 6023 17784 13341 17823
rect 13393 17784 13405 17836
rect 13457 17784 13463 17836
tri 5523 17756 5548 17781 se
tri 5666 17756 5691 17781 sw
rect 13691 17704 13697 17756
rect 13749 17704 13765 17756
rect 13817 17704 13823 17756
rect 10905 17359 10951 17371
rect 10905 17325 10911 17359
rect 10945 17325 10951 17359
rect 1789 17294 1919 17300
rect 1789 17242 1796 17294
rect 1848 17242 1860 17294
rect 1912 17242 1919 17294
rect 1789 17229 1919 17242
rect 10905 17287 10951 17325
rect 10905 17253 10911 17287
rect 10945 17253 10951 17287
rect 10905 17241 10951 17253
rect 1789 17177 1796 17229
rect 1848 17177 1860 17229
rect 1912 17177 1919 17229
rect 1789 17164 1919 17177
rect 1789 17112 1796 17164
rect 1848 17112 1860 17164
rect 1912 17112 1919 17164
rect 1789 17099 1919 17112
rect 1789 17047 1796 17099
rect 1848 17047 1860 17099
rect 1912 17047 1919 17099
rect 1789 17034 1919 17047
rect 1789 16982 1796 17034
rect 1848 16982 1860 17034
rect 1912 16982 1919 17034
rect 1789 16969 1919 16982
rect 1789 16917 1796 16969
rect 1848 16917 1860 16969
rect 1912 16917 1919 16969
rect 1789 16904 1919 16917
rect 1789 16852 1796 16904
rect 1848 16852 1860 16904
rect 1912 16852 1919 16904
rect 1789 16839 1919 16852
rect 1789 16787 1796 16839
rect 1848 16787 1860 16839
rect 1912 16787 1919 16839
rect 1789 16774 1919 16787
rect 1789 16722 1796 16774
rect 1848 16722 1860 16774
rect 1912 16722 1919 16774
rect 1789 16709 1919 16722
rect 1789 16657 1796 16709
rect 1848 16657 1860 16709
rect 1912 16657 1919 16709
rect 1789 16644 1919 16657
rect 1789 16592 1796 16644
rect 1848 16592 1860 16644
rect 1912 16592 1919 16644
rect 1789 16579 1919 16592
rect 1789 16527 1796 16579
rect 1848 16527 1860 16579
rect 1912 16527 1919 16579
rect 1789 16514 1919 16527
rect 1789 16462 1796 16514
rect 1848 16462 1860 16514
rect 1912 16462 1919 16514
rect 1789 16449 1919 16462
rect 1789 16397 1796 16449
rect 1848 16397 1860 16449
rect 1912 16397 1919 16449
rect 1789 16384 1919 16397
rect 1789 16332 1796 16384
rect 1848 16332 1860 16384
rect 1912 16332 1919 16384
rect 1789 16319 1919 16332
rect 1789 16267 1796 16319
rect 1848 16267 1860 16319
rect 1912 16267 1919 16319
rect 1789 16254 1919 16267
rect 1789 16202 1796 16254
rect 1848 16202 1860 16254
rect 1912 16202 1919 16254
rect 1789 16189 1919 16202
rect 1789 16137 1796 16189
rect 1848 16137 1860 16189
rect 1912 16137 1919 16189
rect 1789 16124 1919 16137
rect 1789 16072 1796 16124
rect 1848 16072 1860 16124
rect 1912 16072 1919 16124
rect 1789 16059 1919 16072
rect 1789 16007 1796 16059
rect 1848 16007 1860 16059
rect 1912 16007 1919 16059
rect 1789 15993 1919 16007
rect 1789 15941 1796 15993
rect 1848 15941 1860 15993
rect 1912 15941 1919 15993
rect 1789 15927 1919 15941
rect 1789 15875 1796 15927
rect 1848 15875 1860 15927
rect 1912 15875 1919 15927
rect 1789 15861 1919 15875
rect 1789 15809 1796 15861
rect 1848 15809 1860 15861
rect 1912 15809 1919 15861
rect 1789 15795 1919 15809
rect 1789 15743 1796 15795
rect 1848 15743 1860 15795
rect 1912 15743 1919 15795
rect 1789 15729 1919 15743
rect 1789 15677 1796 15729
rect 1848 15677 1860 15729
rect 1912 15677 1919 15729
rect 1789 15663 1919 15677
rect 1789 15611 1796 15663
rect 1848 15611 1860 15663
rect 1912 15611 1919 15663
rect 1789 15597 1919 15611
rect 1789 15545 1796 15597
rect 1848 15545 1860 15597
rect 1912 15545 1919 15597
rect 1789 15531 1919 15545
rect 1789 15479 1796 15531
rect 1848 15479 1860 15531
rect 1912 15479 1919 15531
rect 1789 15465 1919 15479
rect 1789 15413 1796 15465
rect 1848 15413 1860 15465
rect 1912 15413 1919 15465
rect 1789 15399 1919 15413
rect 1789 15347 1796 15399
rect 1848 15347 1860 15399
rect 1912 15347 1919 15399
rect 1789 15333 1919 15347
rect 1789 15281 1796 15333
rect 1848 15281 1860 15333
rect 1912 15281 1919 15333
rect 1789 15267 1919 15281
rect 1789 15215 1796 15267
rect 1848 15215 1860 15267
rect 1912 15215 1919 15267
rect 1789 15201 1919 15215
rect 1789 15149 1796 15201
rect 1848 15149 1860 15201
rect 1912 15149 1919 15201
rect 1789 15135 1919 15149
rect 1789 15083 1796 15135
rect 1848 15083 1860 15135
rect 1912 15083 1919 15135
rect 1789 15069 1919 15083
rect 1789 15017 1796 15069
rect 1848 15017 1860 15069
rect 1912 15017 1919 15069
rect 1789 15003 1919 15017
rect 1789 14951 1796 15003
rect 1848 14951 1860 15003
rect 1912 14951 1919 15003
rect 1789 14945 1919 14951
rect 9399 11961 9657 11987
rect 9399 11909 9405 11961
rect 9457 11909 9470 11961
rect 9522 11909 9535 11961
rect 9587 11909 9599 11961
rect 9651 11909 9657 11961
rect 9399 11883 9657 11909
rect 1798 11021 1850 11027
rect 1798 10957 1850 10969
rect 1798 10893 1850 10905
rect 1798 10837 1807 10841
rect 1841 10837 1850 10841
rect 1798 10829 1850 10837
rect 1798 10765 1807 10777
rect 1841 10765 1850 10777
rect 473 10641 523 10750
rect 1798 10707 1850 10713
rect 1914 11021 1966 11027
rect 1914 10957 1966 10969
rect 1914 10893 1966 10905
rect 1914 10837 1923 10841
rect 1957 10837 1966 10841
rect 1914 10829 1966 10837
rect 1914 10765 1923 10777
rect 1957 10765 1966 10777
rect 1914 10707 1966 10713
tri 523 10641 548 10666 sw
rect 473 10578 545 10641
rect 473 10577 547 10578
tri 547 10577 548 10578 nw
rect 473 10229 523 10577
tri 523 10552 548 10577 nw
tri 523 10229 548 10254 sw
rect 12029 10236 12157 10242
rect 473 10165 545 10229
rect 473 9717 523 10165
tri 523 10140 548 10165 nw
tri 523 9717 548 9742 sw
rect 473 9653 545 9717
rect 473 9276 523 9653
tri 523 9628 548 9653 nw
rect 1875 9523 1963 10229
rect 12029 10184 12035 10236
rect 12087 10184 12099 10236
rect 12151 10184 12157 10236
rect 12029 10163 12157 10184
rect 12029 10111 12035 10163
rect 12087 10111 12099 10163
rect 12151 10111 12157 10163
rect 12029 10090 12157 10111
rect 12029 10038 12035 10090
rect 12087 10038 12099 10090
rect 12151 10038 12157 10090
rect 12029 10017 12157 10038
rect 12029 9965 12035 10017
rect 12087 9965 12099 10017
rect 12151 9965 12157 10017
rect 12029 9944 12157 9965
rect 12029 9892 12035 9944
rect 12087 9892 12099 9944
rect 12151 9892 12157 9944
rect 12029 9870 12157 9892
rect 12029 9818 12035 9870
rect 12087 9818 12099 9870
rect 12151 9818 12157 9870
rect 12029 9812 12157 9818
rect 12029 9626 12157 9632
rect 12029 9574 12035 9626
rect 12087 9574 12099 9626
rect 12151 9574 12157 9626
rect 12029 9561 12157 9574
tri 1701 9307 1917 9523 ne
rect 12029 9509 12035 9561
rect 12087 9509 12099 9561
rect 12151 9509 12157 9561
rect 12029 9496 12157 9509
rect 12029 9444 12035 9496
rect 12087 9444 12099 9496
rect 12151 9444 12157 9496
rect 12029 9431 12157 9444
rect 12029 9379 12035 9431
rect 12087 9379 12099 9431
rect 12151 9379 12157 9431
rect 12029 9365 12157 9379
rect 12029 9313 12035 9365
rect 12087 9313 12099 9365
rect 12151 9313 12157 9365
tri 523 9276 548 9301 sw
rect 12029 9299 12157 9313
rect 473 9146 628 9276
rect 12029 9247 12035 9299
rect 12087 9247 12099 9299
rect 12151 9247 12157 9299
rect 12029 9233 12157 9247
rect 12029 9181 12035 9233
rect 12087 9181 12099 9233
rect 12151 9181 12157 9233
rect 12029 9175 12157 9181
rect 473 8773 523 9146
tri 523 9121 548 9146 nw
tri 523 8773 626 8876 sw
rect 3361 8767 3413 8773
rect 3361 8703 3413 8715
rect 3361 8645 3413 8651
rect 12029 8596 12157 8602
rect 12029 8544 12035 8596
rect 12087 8544 12099 8596
rect 12151 8544 12157 8596
rect 12029 8529 12157 8544
rect 12029 8477 12035 8529
rect 12087 8477 12099 8529
rect 12151 8477 12157 8529
rect 12029 8462 12157 8477
rect 12029 8410 12035 8462
rect 12087 8410 12099 8462
rect 12151 8410 12157 8462
rect 12029 8395 12157 8410
rect 12029 8343 12035 8395
rect 12087 8343 12099 8395
rect 12151 8343 12157 8395
rect 12029 8328 12157 8343
rect 12029 8276 12035 8328
rect 12087 8276 12099 8328
rect 12151 8276 12157 8328
rect 12029 8270 12157 8276
rect 12029 7336 12157 7342
rect 12029 7284 12035 7336
rect 12087 7284 12099 7336
rect 12151 7284 12157 7336
rect 12029 7269 12157 7284
rect 12029 7217 12035 7269
rect 12087 7217 12099 7269
rect 12151 7217 12157 7269
rect 12029 7202 12157 7217
rect 12029 7150 12035 7202
rect 12087 7150 12099 7202
rect 12151 7150 12157 7202
rect 12029 7135 12157 7150
rect 12029 7083 12035 7135
rect 12087 7083 12099 7135
rect 12151 7083 12157 7135
rect 12029 7068 12157 7083
rect 12029 7016 12035 7068
rect 12087 7016 12099 7068
rect 12151 7016 12157 7068
rect 12029 7010 12157 7016
rect 5489 6748 5495 6864
rect 5675 6748 5681 6864
rect 6670 6748 6676 6864
rect 6856 6748 6862 6864
rect 7192 6748 7198 6864
rect 7378 6748 7384 6864
rect 12029 6824 12157 6830
rect 12029 6772 12035 6824
rect 12087 6772 12099 6824
rect 12151 6772 12157 6824
rect 12029 6750 12157 6772
rect 12029 6698 12035 6750
rect 12087 6698 12099 6750
rect 12151 6698 12157 6750
rect 12029 6675 12157 6698
rect 12029 6623 12035 6675
rect 12087 6623 12099 6675
rect 12151 6623 12157 6675
rect 12029 6600 12157 6623
rect 12029 6548 12035 6600
rect 12087 6548 12099 6600
rect 12151 6548 12157 6600
rect 12029 6525 12157 6548
rect 12029 6473 12035 6525
rect 12087 6473 12099 6525
rect 12151 6473 12157 6525
rect 12029 6467 12157 6473
rect 12029 5578 12157 5584
rect 12029 5526 12035 5578
rect 12087 5526 12099 5578
rect 12151 5526 12157 5578
rect 12029 5505 12157 5526
rect 12029 5453 12035 5505
rect 12087 5453 12099 5505
rect 12151 5453 12157 5505
rect 12029 5432 12157 5453
tri 1604 5420 1615 5431 sw
tri 801 5383 834 5416 se
rect 834 5383 1615 5420
tri 767 5349 801 5383 se
rect 801 5349 846 5383
rect 880 5349 926 5383
rect 960 5349 1005 5383
rect 1039 5349 1084 5383
rect 1118 5349 1163 5383
rect 1197 5349 1242 5383
rect 1276 5349 1321 5383
rect 1355 5349 1400 5383
rect 1434 5349 1479 5383
rect 1513 5349 1558 5383
rect 1592 5349 1615 5383
tri 693 5275 767 5349 se
rect 767 5275 1615 5349
tri 1615 5275 1760 5420 sw
rect 12029 5380 12035 5432
rect 12087 5380 12099 5432
rect 12151 5380 12157 5432
rect 12029 5358 12157 5380
rect 12029 5306 12035 5358
rect 12087 5306 12099 5358
rect 12151 5306 12157 5358
rect 12029 5300 12157 5306
rect 473 5145 1604 5275
rect 3361 5267 3413 5273
rect 3361 5203 3413 5215
rect 3361 5145 3413 5151
rect 473 4770 523 5145
tri 523 5120 548 5145 nw
tri 523 4770 548 4795 sw
rect 473 4640 550 4770
rect 12029 4699 12157 4705
rect 473 4263 523 4640
tri 523 4615 548 4640 nw
tri 1701 4393 1917 4609 se
tri 523 4263 548 4288 sw
rect 473 4199 545 4263
rect 473 3751 523 4199
tri 523 4174 548 4199 nw
tri 523 3751 548 3776 sw
rect 473 3687 545 3751
rect 1875 3687 1963 4393
rect 12029 4391 12035 4699
rect 12151 4391 12157 4699
rect 12029 4378 12157 4391
rect 12029 4326 12035 4378
rect 12087 4326 12099 4378
rect 12151 4326 12157 4378
rect 12029 4313 12157 4326
rect 12029 4261 12035 4313
rect 12087 4261 12099 4313
rect 12151 4261 12157 4313
rect 12029 4255 12157 4261
rect 12029 4066 12157 4072
rect 12029 4014 12035 4066
rect 12087 4014 12099 4066
rect 12151 4014 12157 4066
rect 12029 4000 12157 4014
rect 12029 3948 12035 4000
rect 12087 3948 12099 4000
rect 12151 3948 12157 4000
rect 12029 3934 12157 3948
rect 12029 3882 12035 3934
rect 12087 3882 12099 3934
rect 12151 3882 12157 3934
rect 12029 3868 12157 3882
rect 12029 3816 12035 3868
rect 12087 3816 12099 3868
rect 12151 3816 12157 3868
rect 12029 3802 12157 3816
rect 12029 3750 12035 3802
rect 12087 3750 12099 3802
rect 12151 3750 12157 3802
rect 12029 3736 12157 3750
rect 473 3339 523 3687
tri 523 3662 548 3687 nw
rect 12029 3684 12035 3736
rect 12087 3684 12099 3736
rect 12151 3684 12157 3736
rect 12029 3678 12157 3684
rect 1798 3384 1850 3390
tri 523 3339 548 3364 sw
rect 473 3338 547 3339
tri 547 3338 548 3339 sw
rect 473 3166 545 3338
rect 773 3305 991 3339
rect 773 3271 951 3305
rect 985 3271 991 3305
rect 773 3233 991 3271
rect 773 3199 951 3233
rect 985 3199 991 3233
rect 773 3174 991 3199
rect 773 3166 803 3174
tri 803 3166 811 3174 nw
tri 881 3166 889 3174 ne
rect 889 3166 991 3174
rect 1798 3320 1807 3332
rect 1841 3320 1850 3332
rect 1798 3260 1850 3268
rect 1798 3256 1807 3260
rect 1841 3256 1850 3260
rect 1798 3192 1850 3204
rect 1798 3128 1850 3140
rect 1798 3070 1850 3076
rect 1914 3384 1966 3390
rect 1914 3320 1923 3332
rect 1957 3320 1966 3332
rect 1914 3260 1966 3268
rect 1914 3256 1923 3260
rect 1957 3256 1966 3260
rect 1914 3192 1966 3204
rect 1914 3128 1966 3140
rect 1914 3070 1966 3076
rect 4793 2462 4923 2463
rect 4793 2410 4799 2462
rect 4851 2410 4865 2462
rect 4917 2410 4923 2462
rect 4793 2398 4923 2410
rect 4793 2346 4799 2398
rect 4851 2346 4865 2398
rect 4917 2346 4923 2398
rect 4793 2345 4923 2346
rect 7996 2462 8189 2463
rect 7996 2410 8002 2462
rect 8054 2410 8067 2462
rect 7996 2398 8067 2410
rect 7996 2346 8002 2398
rect 8054 2346 8067 2398
rect 8183 2346 8189 2462
rect 7996 2345 8189 2346
tri 4048 2150 4054 2156 se
rect 4054 2150 4060 2156
rect 4048 2104 4060 2150
rect 4112 2104 4124 2156
rect 4176 2104 4188 2156
rect 4240 2150 4246 2156
tri 4246 2150 4252 2156 sw
rect 4240 2104 4252 2150
tri 5483 2150 5489 2156 se
rect 5489 2150 5495 2156
rect 5483 2104 5495 2150
rect 5547 2104 5559 2156
rect 5611 2104 5623 2156
rect 5675 2150 5681 2156
tri 5681 2150 5687 2156 sw
rect 5675 2104 5687 2150
tri 6664 2150 6670 2156 se
rect 6670 2150 6676 2156
rect 6664 2104 6676 2150
rect 6728 2104 6740 2156
rect 6792 2104 6804 2156
rect 6856 2150 6862 2156
tri 6862 2150 6868 2156 sw
rect 6856 2104 6868 2150
tri 7186 2150 7192 2156 se
rect 7192 2150 7198 2156
rect 7186 2104 7198 2150
rect 7250 2104 7262 2156
rect 7314 2104 7326 2156
rect 7378 2150 7384 2156
tri 7384 2150 7390 2156 sw
rect 7378 2104 7390 2150
tri 8311 2150 8317 2156 se
rect 8317 2150 8323 2156
rect 8311 2104 8323 2150
rect 8375 2104 8391 2156
rect 8443 2104 8458 2156
rect 8510 2104 8525 2156
rect 8577 2150 8583 2156
tri 8583 2150 8589 2156 sw
rect 8577 2104 8589 2150
rect -102 1819 -16 1871
rect 10096 1828 10282 1834
rect 10096 1776 10099 1828
rect 10151 1776 10163 1828
rect 10215 1776 10227 1828
rect 10279 1776 10282 1828
rect 10096 1763 10282 1776
rect -102 1705 -16 1757
rect 10096 1711 10099 1763
rect 10151 1711 10163 1763
rect 10215 1711 10227 1763
rect 10279 1711 10282 1763
rect 10096 1697 10282 1711
rect 10096 1645 10099 1697
rect 10151 1645 10163 1697
rect 10215 1645 10227 1697
rect 10279 1645 10282 1697
rect 10096 1639 10282 1645
rect -102 1580 -15 1632
rect 13859 1622 13975 1732
rect 11359 1492 11941 1504
rect 11993 1492 12020 1504
rect 12072 1492 12099 1504
rect 12151 1492 13421 1504
rect 11359 1486 11437 1492
rect 11359 1452 11365 1486
rect 11399 1458 11437 1486
rect 11471 1458 11509 1492
rect 11543 1458 11581 1492
rect 11615 1458 11653 1492
rect 11687 1458 11725 1492
rect 11759 1458 11797 1492
rect 11831 1458 11869 1492
rect 11903 1458 11941 1492
rect 11993 1458 12013 1492
rect 12072 1458 12085 1492
rect 12151 1458 12157 1492
rect 12191 1458 12229 1492
rect 12263 1458 12301 1492
rect 12335 1458 12373 1492
rect 12407 1458 12445 1492
rect 12479 1458 12517 1492
rect 12551 1458 12589 1492
rect 12623 1458 12661 1492
rect 12695 1458 12733 1492
rect 12767 1458 12805 1492
rect 12839 1458 12877 1492
rect 12911 1458 12949 1492
rect 12983 1458 13021 1492
rect 13055 1458 13093 1492
rect 13127 1458 13165 1492
rect 13199 1458 13237 1492
rect 13271 1458 13309 1492
rect 13343 1486 13421 1492
rect 13343 1458 13381 1486
rect 11399 1452 11941 1458
rect 11993 1452 12020 1458
rect 12072 1452 12099 1458
rect 12151 1452 13381 1458
rect 13415 1452 13421 1486
rect 11359 1412 11518 1452
tri 11518 1412 11558 1452 nw
tri 13223 1412 13263 1452 ne
rect 13263 1412 13421 1452
rect 11359 1406 11512 1412
tri 11512 1406 11518 1412 nw
tri 11589 1406 11595 1412 se
rect 11595 1406 13216 1412
tri 13216 1406 13222 1412 sw
tri 13263 1406 13269 1412 ne
rect 13269 1406 13421 1412
rect 11359 1372 11365 1406
rect 11399 1375 11481 1406
tri 11481 1375 11512 1406 nw
tri 11558 1375 11589 1406 se
rect 11589 1405 13222 1406
tri 13222 1405 13223 1406 sw
tri 13269 1405 13270 1406 ne
rect 13270 1405 13381 1406
rect 11589 1375 13223 1405
rect 11399 1372 11478 1375
tri 11478 1372 11481 1375 nw
tri 11555 1372 11558 1375 se
rect 11558 1372 13223 1375
tri 13223 1372 13256 1405 sw
tri 13270 1372 13303 1405 ne
rect 13303 1372 13381 1405
rect 13415 1372 13421 1406
rect 11359 1325 11431 1372
tri 11431 1325 11478 1372 nw
tri 11508 1325 11555 1372 se
rect 11555 1370 13256 1372
tri 13256 1370 13258 1372 sw
tri 13303 1370 13305 1372 ne
rect 13305 1370 13421 1372
rect 11555 1325 13258 1370
tri 13258 1325 13303 1370 sw
tri 13305 1325 13350 1370 ne
rect 13350 1325 13421 1370
rect 11359 1291 11365 1325
rect 11399 1323 11429 1325
tri 11429 1323 11431 1325 nw
tri 11506 1323 11508 1325 se
rect 11508 1323 13303 1325
tri 13303 1323 13305 1325 sw
rect 11399 1291 11405 1323
tri 11405 1299 11429 1323 nw
tri 11482 1299 11506 1323 se
rect 11506 1299 13305 1323
tri 13350 1300 13375 1325 ne
rect 11359 1244 11405 1291
rect 11359 1210 11365 1244
rect 11399 1210 11405 1244
rect 11359 1163 11405 1210
rect 11359 1129 11365 1163
rect 11399 1129 11405 1163
tri 9402 1082 9424 1104 se
tri 9398 1078 9402 1082 se
rect 9402 1078 9424 1082
rect 4056 1067 4242 1073
rect 4056 1015 4059 1067
rect 4111 1015 4123 1067
rect 4175 1015 4187 1067
rect 4239 1015 4242 1067
rect 4056 1001 4242 1015
rect 4056 949 4059 1001
rect 4111 949 4123 1001
rect 4175 949 4187 1001
rect 4239 949 4242 1001
rect 4056 935 4242 949
rect 4056 883 4059 935
rect 4111 883 4123 935
rect 4175 883 4187 935
rect 4239 883 4242 935
rect 4056 877 4242 883
rect 5491 1067 5677 1073
rect 5491 1015 5494 1067
rect 5546 1015 5558 1067
rect 5610 1015 5622 1067
rect 5674 1015 5677 1067
rect 5491 1001 5677 1015
rect 5491 949 5494 1001
rect 5546 949 5558 1001
rect 5610 949 5622 1001
rect 5674 949 5677 1001
rect 5491 935 5677 949
rect 5491 883 5494 935
rect 5546 883 5558 935
rect 5610 883 5622 935
rect 5674 883 5677 935
rect 5491 877 5677 883
rect 6672 1067 6858 1073
rect 6672 1015 6675 1067
rect 6727 1015 6739 1067
rect 6791 1015 6803 1067
rect 6855 1015 6858 1067
rect 6672 1001 6858 1015
rect 6672 949 6675 1001
rect 6727 949 6739 1001
rect 6791 949 6803 1001
rect 6855 949 6858 1001
rect 6672 935 6858 949
rect 6672 883 6675 935
rect 6727 883 6739 935
rect 6791 883 6803 935
rect 6855 883 6858 935
rect 6672 877 6858 883
rect 7194 1067 7380 1073
rect 7194 1015 7197 1067
rect 7249 1015 7261 1067
rect 7313 1015 7325 1067
rect 7377 1015 7380 1067
rect 7194 1001 7380 1015
rect 7194 949 7197 1001
rect 7249 949 7261 1001
rect 7313 949 7325 1001
rect 7377 949 7380 1001
rect 8321 1067 8579 1071
rect 8321 1015 8327 1067
rect 8379 1015 8392 1067
rect 8444 1015 8457 1067
rect 8321 1003 8457 1015
rect 8321 951 8327 1003
rect 8379 951 8392 1003
rect 8444 951 8457 1003
rect 8321 950 8457 951
rect 7194 935 7380 949
rect 7194 883 7197 935
rect 7249 883 7261 935
rect 7313 883 7325 935
rect 7377 883 7380 935
rect 7927 939 8457 950
rect 7927 922 8327 939
rect 8321 887 8327 922
rect 8379 887 8392 939
rect 8444 887 8457 939
rect 8573 950 8579 1067
rect 9383 950 9424 1078
rect 11359 1082 11405 1129
rect 11359 1048 11365 1082
rect 11399 1048 11405 1082
rect 11359 1036 11405 1048
tri 11475 1292 11482 1299 se
rect 11482 1292 13305 1299
rect 11475 1284 13305 1292
rect 11475 1226 11673 1284
tri 11673 1259 11698 1284 nw
tri 11830 1259 11855 1284 ne
rect 11475 1192 11481 1226
rect 11515 1192 11673 1226
rect 11475 1154 11673 1192
rect 11475 1120 11481 1154
rect 11515 1120 11673 1154
rect 11475 1082 11673 1120
rect 11475 1048 11481 1082
rect 11515 1048 11673 1082
tri 11450 986 11475 1011 se
rect 11475 986 11673 1048
rect 8573 922 9424 950
rect 8573 887 8579 922
rect 8321 883 8579 887
rect 10984 903 11673 986
rect 10984 883 11653 903
tri 11653 883 11673 903 nw
rect 11731 1226 11777 1238
rect 11731 1192 11737 1226
rect 11771 1192 11777 1226
rect 11731 1154 11777 1192
rect 11731 1120 11737 1154
rect 11771 1120 11777 1154
rect 11731 1082 11777 1120
rect 11731 1048 11737 1082
rect 11771 1048 11777 1082
rect 7194 877 7380 883
rect 10984 877 11647 883
tri 11647 877 11653 883 nw
rect 10984 870 11640 877
tri 11640 870 11647 877 nw
rect 11359 814 11521 826
rect 10096 785 10282 791
rect 10096 733 10099 785
rect 10151 733 10163 785
rect 10215 733 10227 785
rect 10279 733 10282 785
rect 10096 720 10282 733
rect 7996 710 8189 711
rect 7996 658 8002 710
rect 8054 658 8067 710
rect 7996 646 8067 658
rect -102 588 -35 640
rect 4787 593 4801 639
tri 4787 590 4790 593 ne
rect 4790 590 4801 593
tri 4790 588 4792 590 ne
rect 4792 588 4801 590
tri 4792 587 4793 588 ne
rect 4793 587 4801 588
rect 4853 587 4865 639
rect 4917 593 4929 639
rect 7996 594 8002 646
rect 8054 594 8067 646
rect 8183 594 8189 710
rect 10096 668 10099 720
rect 10151 668 10163 720
rect 10215 668 10227 720
rect 10279 668 10282 720
rect 10096 654 10282 668
rect 10096 602 10099 654
rect 10151 602 10163 654
rect 10215 602 10227 654
rect 10279 602 10282 654
rect 10096 596 10282 602
rect 11359 780 11365 814
rect 11399 780 11481 814
rect 11515 780 11521 814
rect 11359 742 11521 780
rect 11359 719 11481 742
rect 11359 685 11365 719
rect 11399 708 11481 719
rect 11515 708 11521 742
rect 11399 685 11521 708
rect 11359 670 11521 685
rect 11359 636 11481 670
rect 11515 636 11521 670
rect 11359 624 11521 636
rect 11731 814 11777 1048
rect 11855 1226 11901 1284
tri 11901 1259 11926 1284 nw
tri 12342 1259 12367 1284 ne
rect 11855 1192 11861 1226
rect 11895 1192 11901 1226
rect 11855 1154 11901 1192
rect 11855 1120 11861 1154
rect 11895 1120 11901 1154
rect 11855 1082 11901 1120
rect 11855 1048 11861 1082
rect 11895 1048 11901 1082
rect 11855 1036 11901 1048
rect 12081 1226 12157 1238
rect 12081 1192 12117 1226
rect 12151 1192 12157 1226
rect 12081 1154 12157 1192
rect 12081 1120 12117 1154
rect 12151 1120 12157 1154
rect 12081 1082 12157 1120
rect 12234 1232 12286 1238
rect 12234 1166 12286 1180
rect 12234 1108 12286 1114
rect 12367 1226 12413 1284
tri 12413 1259 12438 1284 nw
tri 12854 1259 12879 1284 ne
rect 12367 1192 12373 1226
rect 12407 1192 12413 1226
rect 12367 1154 12413 1192
rect 12367 1120 12373 1154
rect 12407 1120 12413 1154
rect 12081 1048 12117 1082
rect 12151 1048 12157 1082
rect 12081 1036 12157 1048
rect 12367 1082 12413 1120
rect 12494 1232 12546 1238
rect 12494 1166 12546 1180
rect 12494 1108 12546 1114
rect 12623 1226 12699 1238
rect 12623 1192 12629 1226
rect 12663 1192 12699 1226
rect 12623 1154 12699 1192
rect 12623 1120 12629 1154
rect 12663 1120 12699 1154
rect 12367 1048 12373 1082
rect 12407 1048 12413 1082
rect 12367 1036 12413 1048
rect 12623 1082 12699 1120
rect 12623 1048 12629 1082
rect 12663 1048 12699 1082
rect 12623 1036 12699 1048
rect 12879 1226 12925 1284
tri 12925 1259 12950 1284 nw
tri 13234 1259 13259 1284 ne
rect 12879 1192 12885 1226
rect 12919 1192 12925 1226
rect 12879 1154 12925 1192
rect 12879 1120 12885 1154
rect 12919 1120 12925 1154
rect 12879 1082 12925 1120
rect 12879 1048 12885 1082
rect 12919 1048 12925 1082
rect 12879 1036 12925 1048
rect 13003 1226 13049 1238
rect 13003 1192 13009 1226
rect 13043 1192 13049 1226
rect 13003 1154 13049 1192
rect 13003 1120 13009 1154
rect 13043 1120 13049 1154
rect 13003 1082 13049 1120
rect 13003 1048 13009 1082
rect 13043 1048 13049 1082
rect 11731 780 11737 814
rect 11771 780 11777 814
rect 11731 742 11777 780
rect 11731 708 11737 742
rect 11771 708 11777 742
rect 11731 670 11777 708
rect 11731 636 11737 670
rect 11771 636 11777 670
rect 11731 624 11777 636
rect 11987 814 12033 826
rect 11987 780 11993 814
rect 12027 780 12033 814
rect 11987 742 12033 780
rect 11987 708 11993 742
rect 12027 708 12033 742
rect 11987 670 12033 708
rect 11987 636 11993 670
rect 12027 636 12033 670
rect 7996 593 8189 594
rect 4917 590 4926 593
tri 4926 590 4929 593 nw
rect 11359 590 11365 624
rect 11399 596 11521 624
tri 11521 596 11534 609 sw
tri 11974 596 11987 609 se
rect 11987 596 12033 636
rect 12081 685 12127 1036
tri 12127 1006 12157 1036 nw
tri 12623 1006 12653 1036 ne
tri 12127 685 12131 689 sw
rect 12081 678 12131 685
tri 12131 678 12138 685 sw
rect 12363 678 12409 690
tri 12649 685 12653 689 se
rect 12653 685 12699 1036
rect 12081 664 12138 678
tri 12138 664 12152 678 sw
rect 12081 658 12283 664
rect 12081 624 12093 658
rect 12127 624 12165 658
rect 12199 624 12237 658
rect 12271 624 12283 658
rect 12081 618 12283 624
rect 12363 644 12369 678
rect 12403 644 12409 678
tri 12634 670 12649 685 se
rect 12649 670 12699 685
tri 12628 664 12634 670 se
rect 12634 664 12699 670
tri 12033 596 12046 609 sw
tri 12350 596 12363 609 se
rect 12363 596 12409 644
rect 12497 658 12699 664
rect 12497 624 12509 658
rect 12543 624 12581 658
rect 12615 624 12653 658
rect 12687 624 12699 658
rect 12497 618 12699 624
rect 12747 814 12793 826
rect 12747 780 12753 814
rect 12787 780 12793 814
rect 12747 742 12793 780
rect 12747 708 12753 742
rect 12787 708 12793 742
rect 12747 670 12793 708
rect 12747 636 12753 670
rect 12787 636 12793 670
tri 12409 596 12422 609 sw
tri 12734 596 12747 609 se
rect 12747 596 12793 636
rect 13003 814 13049 1048
rect 13259 1226 13305 1284
rect 13259 1192 13265 1226
rect 13299 1192 13305 1226
rect 13259 1154 13305 1192
rect 13259 1120 13265 1154
rect 13299 1120 13305 1154
rect 13259 1082 13305 1120
rect 13259 1048 13265 1082
rect 13299 1048 13305 1082
rect 13259 1036 13305 1048
rect 13375 1291 13381 1325
rect 13415 1291 13421 1325
rect 13375 1244 13421 1291
rect 13375 1210 13381 1244
rect 13415 1210 13421 1244
rect 13375 1163 13421 1210
rect 13375 1129 13381 1163
rect 13415 1129 13421 1163
rect 13375 1082 13421 1129
rect 13375 1048 13381 1082
rect 13415 1048 13421 1082
rect 13375 1036 13421 1048
tri 13506 826 13531 851 se
rect 13531 826 13693 1598
rect 13003 780 13009 814
rect 13043 780 13049 814
rect 13003 742 13049 780
rect 13003 708 13009 742
rect 13043 708 13049 742
rect 13003 670 13049 708
rect 13003 636 13009 670
rect 13043 636 13049 670
rect 13003 624 13049 636
rect 13259 814 13693 826
rect 13259 780 13265 814
rect 13299 780 13381 814
rect 13415 780 13693 814
rect 13259 742 13693 780
rect 13259 708 13265 742
rect 13299 719 13693 742
rect 13299 708 13381 719
rect 13259 685 13381 708
rect 13415 685 13693 719
rect 13259 670 13693 685
rect 13259 636 13265 670
rect 13299 636 13693 670
rect 13259 624 13693 636
tri 12793 596 12806 609 sw
tri 13246 596 13259 609 se
rect 13259 596 13381 624
rect 11399 594 11534 596
tri 11534 594 11536 596 sw
tri 11972 594 11974 596 se
rect 11974 594 12046 596
tri 12046 594 12048 596 sw
tri 12348 594 12350 596 se
rect 12350 594 12422 596
rect 11399 593 11536 594
tri 11536 593 11537 594 sw
tri 11971 593 11972 594 se
rect 11972 593 12048 594
tri 12048 593 12049 594 sw
tri 12347 593 12348 594 se
rect 12348 593 12369 594
rect 11399 590 11537 593
rect 4917 587 4923 590
tri 4923 587 4926 590 nw
rect 11359 587 11537 590
tri 11537 587 11543 593 sw
tri 11965 587 11971 593 se
rect 11971 587 12049 593
tri 12049 587 12055 593 sw
tri 12341 587 12347 593 se
rect 12347 587 12369 593
rect 11359 584 11543 587
tri 11543 584 11546 587 sw
tri 11962 584 11965 587 se
rect 11965 584 12055 587
tri 12055 584 12058 587 sw
tri 12338 584 12341 587 se
rect 12341 584 12369 587
rect 11359 560 12369 584
rect 12403 593 12422 594
tri 12422 593 12425 596 sw
tri 12731 593 12734 596 se
rect 12734 593 12806 596
tri 12806 593 12809 596 sw
tri 13243 593 13246 596 se
rect 13246 593 13381 596
rect 12403 590 12425 593
tri 12425 590 12428 593 sw
tri 12728 590 12731 593 se
rect 12731 590 12809 593
tri 12809 590 12812 593 sw
tri 13240 590 13243 593 se
rect 13243 590 13381 593
rect 13415 603 13693 624
tri 13693 603 13725 635 sw
rect 13415 590 13725 603
rect 12403 587 12428 590
tri 12428 587 12431 590 sw
tri 12725 587 12728 590 se
rect 12728 587 12812 590
tri 12812 587 12815 590 sw
tri 13237 587 13240 590 se
rect 13240 587 13725 590
rect 12403 584 12431 587
tri 12431 584 12434 587 sw
tri 12722 584 12725 587 se
rect 12725 584 12815 587
tri 12815 584 12818 587 sw
tri 13234 584 13237 587 se
rect 13237 584 13725 587
rect 12403 560 13725 584
rect -102 496 -33 548
rect -29 496 23 548
rect 24 497 25 547
rect 53 497 54 547
rect 55 521 107 548
rect 11359 528 13725 560
rect 13913 547 13975 1622
rect 13827 528 13975 547
rect 55 496 210 521
rect 80 471 210 496
rect 11359 494 11365 528
rect 11399 522 13381 528
rect 11399 494 11437 522
rect 11359 488 11437 494
rect 11471 488 11509 522
rect 11543 488 11581 522
rect 11615 488 11653 522
rect 11687 488 11725 522
rect 11759 488 11797 522
rect 11831 488 11869 522
rect 11903 488 11941 522
rect 11975 488 12013 522
rect 12047 488 12085 522
rect 12119 488 12157 522
rect 12191 488 12229 522
rect 12263 488 12301 522
rect 12335 488 12373 522
rect 12407 488 12445 522
rect 12479 488 12517 522
rect 12551 488 12589 522
rect 12623 488 12661 522
rect 12695 488 12733 522
rect 12767 488 12805 522
rect 12839 488 12877 522
rect 12911 488 12949 522
rect 12983 488 13021 522
rect 13055 488 13093 522
rect 13127 488 13165 522
rect 13199 488 13237 522
rect 13271 488 13309 522
rect 13343 494 13381 522
rect 13415 494 13725 528
rect 13343 488 13725 494
rect 11359 482 13725 488
rect 81 469 209 470
rect 80 435 210 469
rect 81 434 209 435
rect -102 356 -5 408
rect 80 381 210 433
rect -102 276 2 328
tri 1288 107 1294 113 se
rect 1294 107 1300 113
rect 1288 61 1300 107
rect 1352 61 1366 113
rect 1418 61 1432 113
rect 1484 61 1498 113
rect 1550 61 1564 113
rect 1616 61 1630 113
rect 1682 61 1696 113
rect 1748 61 1762 113
rect 1814 61 1827 113
rect 1879 61 1892 113
rect 1944 61 1957 113
rect 2009 61 2022 113
rect 2074 61 2087 113
rect 2139 61 2152 113
rect 2204 61 2217 113
rect 2269 61 2282 113
rect 2334 61 2347 113
rect 2399 107 2405 113
tri 2405 107 2411 113 sw
rect 2399 61 2411 107
tri 4048 107 4054 113 se
rect 4054 107 4060 113
rect 4048 61 4060 107
rect 4112 61 4124 113
rect 4176 61 4188 113
rect 4240 107 4246 113
tri 4246 107 4252 113 sw
rect 4240 61 4252 107
tri 5483 107 5489 113 se
rect 5489 107 5495 113
rect 5483 61 5495 107
rect 5547 61 5559 113
rect 5611 61 5623 113
rect 5675 107 5681 113
tri 5681 107 5687 113 sw
rect 5675 61 5687 107
tri 6664 107 6670 113 se
rect 6670 107 6676 113
rect 6664 61 6676 107
rect 6728 61 6740 113
rect 6792 61 6804 113
rect 6856 107 6862 113
tri 6862 107 6868 113 sw
rect 6856 61 6868 107
tri 7186 107 7192 113 se
rect 7192 107 7198 113
rect 7186 61 7198 107
rect 7250 61 7262 113
rect 7314 61 7326 113
rect 7378 107 7384 113
tri 7384 107 7390 113 sw
rect 7378 61 7390 107
tri 8311 107 8317 113 se
rect 8317 107 8323 113
rect 8311 61 8323 107
rect 8375 61 8391 113
rect 8443 61 8458 113
rect 8510 61 8525 113
rect 8577 107 8583 113
tri 8583 107 8589 113 sw
rect 8577 61 8589 107
tri 10739 107 10745 113 se
rect 10745 107 10751 113
rect 10739 61 10751 107
rect 10803 61 10819 113
rect 10871 61 10886 113
rect 10938 61 10953 113
rect 11005 107 11011 113
tri 11011 107 11017 113 sw
rect 11005 61 11017 107
<< rmetal1 >>
rect 23 547 25 548
rect 23 497 24 547
rect 23 496 25 497
rect 53 547 55 548
rect 54 497 55 547
rect 53 496 55 497
rect 80 470 210 471
rect 80 469 81 470
rect 209 469 210 470
rect 80 434 81 435
rect 209 434 210 435
rect 80 433 210 434
<< via1 >>
rect 4679 29805 4731 29857
rect 4743 29805 4795 29857
rect 5097 29805 5149 29857
rect 5161 29805 5213 29857
rect 5243 29805 5295 29857
rect 5307 29805 5359 29857
rect 8928 29681 8980 29733
rect 8928 29617 8980 29669
rect 9008 29681 9060 29733
rect 9008 29617 9060 29669
rect 1680 29483 1732 29535
rect 1733 29426 1785 29478
rect 2034 29471 2086 29523
rect 2098 29505 2150 29557
rect 7564 29505 7616 29557
rect 7628 29505 7680 29557
rect 8004 29505 8056 29557
rect 8068 29505 8120 29557
rect 7564 29416 7616 29468
rect 7628 29416 7680 29468
rect 8004 29416 8056 29468
rect 8068 29416 8120 29468
rect 1680 29340 1732 29392
rect 2098 29358 2150 29410
rect 1734 29285 1786 29337
rect 2098 29294 2150 29346
rect 13024 26969 13076 26973
rect 13093 26969 13145 26973
rect 13162 26969 13214 26973
rect 13231 26969 13283 26973
rect 13300 26969 13352 26973
rect 13369 26969 13421 26973
rect 13439 26969 13491 26973
rect 13509 26969 13561 26973
rect 13579 26969 13631 26973
rect 13649 26969 13701 26973
rect 13024 26935 13048 26969
rect 13048 26935 13076 26969
rect 13093 26935 13121 26969
rect 13121 26935 13145 26969
rect 13162 26935 13194 26969
rect 13194 26935 13214 26969
rect 13231 26935 13267 26969
rect 13267 26935 13283 26969
rect 13300 26935 13301 26969
rect 13301 26935 13340 26969
rect 13340 26935 13352 26969
rect 13369 26935 13374 26969
rect 13374 26935 13413 26969
rect 13413 26935 13421 26969
rect 13439 26935 13447 26969
rect 13447 26935 13486 26969
rect 13486 26935 13491 26969
rect 13509 26935 13520 26969
rect 13520 26935 13559 26969
rect 13559 26935 13561 26969
rect 13579 26935 13593 26969
rect 13593 26935 13631 26969
rect 13649 26935 13666 26969
rect 13666 26935 13701 26969
rect 13024 26921 13076 26935
rect 13093 26921 13145 26935
rect 13162 26921 13214 26935
rect 13231 26921 13283 26935
rect 13300 26921 13352 26935
rect 13369 26921 13421 26935
rect 13439 26921 13491 26935
rect 13509 26921 13561 26935
rect 13579 26921 13631 26935
rect 13649 26921 13701 26935
rect 13024 26867 13076 26909
rect 13093 26867 13145 26909
rect 13162 26867 13214 26909
rect 13231 26867 13283 26909
rect 13300 26867 13352 26909
rect 13369 26867 13421 26909
rect 13439 26867 13491 26909
rect 13024 26857 13029 26867
rect 13029 26857 13068 26867
rect 13068 26857 13076 26867
rect 13093 26857 13102 26867
rect 13102 26857 13141 26867
rect 13141 26857 13145 26867
rect 13162 26857 13175 26867
rect 13175 26857 13214 26867
rect 13231 26857 13249 26867
rect 13249 26857 13283 26867
rect 13300 26857 13323 26867
rect 13323 26857 13352 26867
rect 13369 26857 13397 26867
rect 13397 26857 13421 26867
rect 13439 26857 13471 26867
rect 13471 26857 13491 26867
rect 13509 26867 13561 26909
rect 13509 26857 13511 26867
rect 13511 26857 13545 26867
rect 13545 26857 13561 26867
rect 13579 26867 13631 26909
rect 13579 26857 13585 26867
rect 13585 26857 13619 26867
rect 13619 26857 13631 26867
rect 13649 26867 13701 26909
rect 13649 26857 13659 26867
rect 13659 26857 13693 26867
rect 13693 26857 13701 26867
rect 13024 26833 13029 26845
rect 13029 26833 13068 26845
rect 13068 26833 13076 26845
rect 13093 26833 13102 26845
rect 13102 26833 13141 26845
rect 13141 26833 13145 26845
rect 13162 26833 13175 26845
rect 13175 26833 13214 26845
rect 13231 26833 13249 26845
rect 13249 26833 13283 26845
rect 13300 26833 13323 26845
rect 13323 26833 13352 26845
rect 13369 26833 13397 26845
rect 13397 26833 13421 26845
rect 13439 26833 13471 26845
rect 13471 26833 13491 26845
rect 13024 26793 13076 26833
rect 13093 26793 13145 26833
rect 13162 26793 13214 26833
rect 13231 26793 13283 26833
rect 13300 26793 13352 26833
rect 13369 26793 13421 26833
rect 13439 26793 13491 26833
rect 13509 26833 13511 26845
rect 13511 26833 13545 26845
rect 13545 26833 13561 26845
rect 13509 26793 13561 26833
rect 13579 26833 13585 26845
rect 13585 26833 13619 26845
rect 13619 26833 13631 26845
rect 13579 26793 13631 26833
rect 13649 26833 13659 26845
rect 13659 26833 13693 26845
rect 13693 26833 13701 26845
rect 13649 26793 13701 26833
rect 13024 26765 13076 26781
rect 13024 26731 13035 26765
rect 13035 26731 13069 26765
rect 13069 26731 13076 26765
rect 13024 26729 13076 26731
rect 13093 26765 13145 26781
rect 13093 26731 13108 26765
rect 13108 26731 13142 26765
rect 13142 26731 13145 26765
rect 13093 26729 13145 26731
rect 13162 26765 13214 26781
rect 13231 26765 13283 26781
rect 13300 26765 13352 26781
rect 13369 26765 13421 26781
rect 13439 26765 13491 26781
rect 13509 26765 13561 26781
rect 13579 26765 13631 26781
rect 13649 26765 13701 26781
rect 13162 26731 13181 26765
rect 13181 26731 13214 26765
rect 13231 26731 13254 26765
rect 13254 26731 13283 26765
rect 13300 26731 13327 26765
rect 13327 26731 13352 26765
rect 13369 26731 13400 26765
rect 13400 26731 13421 26765
rect 13439 26731 13473 26765
rect 13473 26731 13491 26765
rect 13509 26731 13546 26765
rect 13546 26731 13561 26765
rect 13579 26731 13580 26765
rect 13580 26731 13619 26765
rect 13619 26731 13631 26765
rect 13649 26731 13653 26765
rect 13653 26731 13692 26765
rect 13692 26731 13701 26765
rect 14820 26992 15256 27556
rect 14820 26927 14872 26979
rect 14884 26927 14936 26979
rect 14948 26927 15000 26979
rect 15012 26927 15064 26979
rect 15076 26927 15128 26979
rect 15140 26927 15192 26979
rect 15204 26927 15256 26979
rect 13162 26729 13214 26731
rect 13231 26729 13283 26731
rect 13300 26729 13352 26731
rect 13369 26729 13421 26731
rect 13439 26729 13491 26731
rect 13509 26729 13561 26731
rect 13579 26729 13631 26731
rect 13649 26729 13701 26731
rect 13022 26248 13074 26253
rect 13092 26248 13144 26253
rect 13162 26248 13214 26253
rect 13232 26248 13284 26253
rect 13302 26248 13354 26253
rect 13372 26248 13424 26253
rect 13442 26248 13494 26253
rect 13512 26248 13564 26253
rect 13582 26248 13634 26253
rect 13022 26214 13039 26248
rect 13039 26214 13074 26248
rect 13092 26214 13111 26248
rect 13111 26214 13144 26248
rect 13162 26214 13183 26248
rect 13183 26214 13214 26248
rect 13232 26214 13255 26248
rect 13255 26214 13284 26248
rect 13302 26214 13327 26248
rect 13327 26214 13354 26248
rect 13372 26214 13399 26248
rect 13399 26214 13424 26248
rect 13442 26214 13471 26248
rect 13471 26214 13494 26248
rect 13512 26214 13543 26248
rect 13543 26214 13564 26248
rect 13582 26214 13615 26248
rect 13615 26214 13634 26248
rect 13022 26201 13074 26214
rect 13092 26201 13144 26214
rect 13162 26201 13214 26214
rect 13232 26201 13284 26214
rect 13302 26201 13354 26214
rect 13372 26201 13424 26214
rect 13442 26201 13494 26214
rect 13512 26201 13564 26214
rect 13582 26201 13634 26214
rect 13652 26248 13704 26253
rect 13652 26214 13653 26248
rect 13653 26214 13687 26248
rect 13687 26214 13704 26248
rect 13652 26201 13704 26214
rect 13022 26174 13074 26186
rect 13092 26174 13144 26186
rect 13162 26174 13214 26186
rect 13232 26174 13284 26186
rect 13302 26174 13354 26186
rect 13372 26174 13424 26186
rect 13442 26174 13494 26186
rect 13512 26174 13564 26186
rect 13582 26174 13634 26186
rect 13022 26140 13039 26174
rect 13039 26140 13074 26174
rect 13092 26140 13111 26174
rect 13111 26140 13144 26174
rect 13162 26140 13183 26174
rect 13183 26140 13214 26174
rect 13232 26140 13255 26174
rect 13255 26140 13284 26174
rect 13302 26140 13327 26174
rect 13327 26140 13354 26174
rect 13372 26140 13399 26174
rect 13399 26140 13424 26174
rect 13442 26140 13471 26174
rect 13471 26140 13494 26174
rect 13512 26140 13543 26174
rect 13543 26140 13564 26174
rect 13582 26140 13615 26174
rect 13615 26140 13634 26174
rect 13022 26134 13074 26140
rect 13092 26134 13144 26140
rect 13162 26134 13214 26140
rect 13232 26134 13284 26140
rect 13302 26134 13354 26140
rect 13372 26134 13424 26140
rect 13442 26134 13494 26140
rect 13512 26134 13564 26140
rect 13582 26134 13634 26140
rect 13652 26174 13704 26186
rect 13652 26140 13653 26174
rect 13653 26140 13687 26174
rect 13687 26140 13704 26174
rect 13652 26134 13704 26140
rect 13022 26100 13074 26119
rect 13092 26100 13144 26119
rect 13162 26100 13214 26119
rect 13232 26100 13284 26119
rect 13302 26100 13354 26119
rect 13372 26100 13424 26119
rect 13442 26100 13494 26119
rect 13512 26100 13564 26119
rect 13582 26100 13634 26119
rect 13022 26067 13039 26100
rect 13039 26067 13074 26100
rect 13092 26067 13111 26100
rect 13111 26067 13144 26100
rect 13162 26067 13183 26100
rect 13183 26067 13214 26100
rect 13232 26067 13255 26100
rect 13255 26067 13284 26100
rect 13302 26067 13327 26100
rect 13327 26067 13354 26100
rect 13372 26067 13399 26100
rect 13399 26067 13424 26100
rect 13442 26067 13471 26100
rect 13471 26067 13494 26100
rect 13512 26067 13543 26100
rect 13543 26067 13564 26100
rect 13582 26067 13615 26100
rect 13615 26067 13634 26100
rect 13652 26100 13704 26119
rect 13652 26067 13653 26100
rect 13653 26067 13687 26100
rect 13687 26067 13704 26100
rect 13022 26026 13074 26052
rect 13092 26026 13144 26052
rect 13162 26026 13214 26052
rect 13232 26026 13284 26052
rect 13302 26026 13354 26052
rect 13372 26026 13424 26052
rect 13442 26026 13494 26052
rect 13512 26026 13564 26052
rect 13582 26026 13634 26052
rect 13022 26000 13039 26026
rect 13039 26000 13074 26026
rect 13092 26000 13111 26026
rect 13111 26000 13144 26026
rect 13162 26000 13183 26026
rect 13183 26000 13214 26026
rect 13232 26000 13255 26026
rect 13255 26000 13284 26026
rect 13302 26000 13327 26026
rect 13327 26000 13354 26026
rect 13372 26000 13399 26026
rect 13399 26000 13424 26026
rect 13442 26000 13471 26026
rect 13471 26000 13494 26026
rect 13512 26000 13543 26026
rect 13543 26000 13564 26026
rect 13582 26000 13615 26026
rect 13615 26000 13634 26026
rect 13652 26026 13704 26052
rect 13652 26000 13653 26026
rect 13653 26000 13687 26026
rect 13687 26000 13704 26026
rect 13022 25953 13074 25985
rect 13092 25953 13144 25985
rect 13162 25953 13214 25985
rect 13232 25953 13284 25985
rect 13302 25953 13354 25985
rect 13372 25953 13424 25985
rect 13442 25953 13494 25985
rect 13512 25953 13564 25985
rect 13582 25953 13634 25985
rect 13022 25933 13039 25953
rect 13039 25933 13074 25953
rect 13092 25933 13111 25953
rect 13111 25933 13144 25953
rect 13162 25933 13183 25953
rect 13183 25933 13214 25953
rect 13232 25933 13255 25953
rect 13255 25933 13284 25953
rect 13302 25933 13327 25953
rect 13327 25933 13354 25953
rect 13372 25933 13399 25953
rect 13399 25933 13424 25953
rect 13442 25933 13471 25953
rect 13471 25933 13494 25953
rect 13512 25933 13543 25953
rect 13543 25933 13564 25953
rect 13582 25933 13615 25953
rect 13615 25933 13634 25953
rect 13652 25953 13704 25985
rect 13652 25933 13653 25953
rect 13653 25933 13687 25953
rect 13687 25933 13704 25953
rect 13022 25880 13074 25918
rect 13092 25880 13144 25918
rect 13162 25880 13214 25918
rect 13232 25880 13284 25918
rect 13302 25880 13354 25918
rect 13372 25880 13424 25918
rect 13442 25880 13494 25918
rect 13512 25880 13564 25918
rect 13582 25880 13634 25918
rect 13022 25866 13039 25880
rect 13039 25866 13074 25880
rect 13092 25866 13111 25880
rect 13111 25866 13144 25880
rect 13162 25866 13183 25880
rect 13183 25866 13214 25880
rect 13232 25866 13255 25880
rect 13255 25866 13284 25880
rect 13302 25866 13327 25880
rect 13327 25866 13354 25880
rect 13372 25866 13399 25880
rect 13399 25866 13424 25880
rect 13442 25866 13471 25880
rect 13471 25866 13494 25880
rect 13512 25866 13543 25880
rect 13543 25866 13564 25880
rect 13582 25866 13615 25880
rect 13615 25866 13634 25880
rect 13652 25880 13704 25918
rect 13652 25866 13653 25880
rect 13653 25866 13687 25880
rect 13687 25866 13704 25880
rect 13022 25846 13039 25851
rect 13039 25846 13074 25851
rect 13092 25846 13111 25851
rect 13111 25846 13144 25851
rect 13162 25846 13183 25851
rect 13183 25846 13214 25851
rect 13232 25846 13255 25851
rect 13255 25846 13284 25851
rect 13302 25846 13327 25851
rect 13327 25846 13354 25851
rect 13372 25846 13399 25851
rect 13399 25846 13424 25851
rect 13442 25846 13471 25851
rect 13471 25846 13494 25851
rect 13512 25846 13543 25851
rect 13543 25846 13564 25851
rect 13582 25846 13615 25851
rect 13615 25846 13634 25851
rect 13022 25807 13074 25846
rect 13092 25807 13144 25846
rect 13162 25807 13214 25846
rect 13232 25807 13284 25846
rect 13302 25807 13354 25846
rect 13372 25807 13424 25846
rect 13442 25807 13494 25846
rect 13512 25807 13564 25846
rect 13582 25807 13634 25846
rect 13022 25799 13039 25807
rect 13039 25799 13074 25807
rect 13092 25799 13111 25807
rect 13111 25799 13144 25807
rect 13162 25799 13183 25807
rect 13183 25799 13214 25807
rect 13232 25799 13255 25807
rect 13255 25799 13284 25807
rect 13302 25799 13327 25807
rect 13327 25799 13354 25807
rect 13372 25799 13399 25807
rect 13399 25799 13424 25807
rect 13442 25799 13471 25807
rect 13471 25799 13494 25807
rect 13512 25799 13543 25807
rect 13543 25799 13564 25807
rect 13582 25799 13615 25807
rect 13615 25799 13634 25807
rect 13652 25846 13653 25851
rect 13653 25846 13687 25851
rect 13687 25846 13704 25851
rect 13652 25807 13704 25846
rect 13652 25799 13653 25807
rect 13653 25799 13687 25807
rect 13687 25799 13704 25807
rect 13022 25773 13039 25784
rect 13039 25773 13074 25784
rect 13092 25773 13111 25784
rect 13111 25773 13144 25784
rect 13162 25773 13183 25784
rect 13183 25773 13214 25784
rect 13232 25773 13255 25784
rect 13255 25773 13284 25784
rect 13302 25773 13327 25784
rect 13327 25773 13354 25784
rect 13372 25773 13399 25784
rect 13399 25773 13424 25784
rect 13442 25773 13471 25784
rect 13471 25773 13494 25784
rect 13512 25773 13543 25784
rect 13543 25773 13564 25784
rect 13582 25773 13615 25784
rect 13615 25773 13634 25784
rect 13022 25734 13074 25773
rect 13092 25734 13144 25773
rect 13162 25734 13214 25773
rect 13232 25734 13284 25773
rect 13302 25734 13354 25773
rect 13372 25734 13424 25773
rect 13442 25734 13494 25773
rect 13512 25734 13564 25773
rect 13582 25734 13634 25773
rect 13022 25732 13039 25734
rect 13039 25732 13074 25734
rect 13092 25732 13111 25734
rect 13111 25732 13144 25734
rect 13162 25732 13183 25734
rect 13183 25732 13214 25734
rect 13232 25732 13255 25734
rect 13255 25732 13284 25734
rect 13302 25732 13327 25734
rect 13327 25732 13354 25734
rect 13372 25732 13399 25734
rect 13399 25732 13424 25734
rect 13442 25732 13471 25734
rect 13471 25732 13494 25734
rect 13512 25732 13543 25734
rect 13543 25732 13564 25734
rect 13582 25732 13615 25734
rect 13615 25732 13634 25734
rect 13652 25773 13653 25784
rect 13653 25773 13687 25784
rect 13687 25773 13704 25784
rect 13652 25734 13704 25773
rect 13652 25732 13653 25734
rect 13653 25732 13687 25734
rect 13687 25732 13704 25734
rect 13022 25700 13039 25717
rect 13039 25700 13074 25717
rect 13092 25700 13111 25717
rect 13111 25700 13144 25717
rect 13162 25700 13183 25717
rect 13183 25700 13214 25717
rect 13232 25700 13255 25717
rect 13255 25700 13284 25717
rect 13302 25700 13327 25717
rect 13327 25700 13354 25717
rect 13372 25700 13399 25717
rect 13399 25700 13424 25717
rect 13442 25700 13471 25717
rect 13471 25700 13494 25717
rect 13512 25700 13543 25717
rect 13543 25700 13564 25717
rect 13582 25700 13615 25717
rect 13615 25700 13634 25717
rect 13022 25665 13074 25700
rect 13092 25665 13144 25700
rect 13162 25665 13214 25700
rect 13232 25665 13284 25700
rect 13302 25665 13354 25700
rect 13372 25665 13424 25700
rect 13442 25665 13494 25700
rect 13512 25665 13564 25700
rect 13582 25665 13634 25700
rect 13652 25700 13653 25717
rect 13653 25700 13687 25717
rect 13687 25700 13704 25717
rect 13652 25665 13704 25700
rect 13022 25627 13039 25650
rect 13039 25627 13074 25650
rect 13092 25627 13111 25650
rect 13111 25627 13144 25650
rect 13162 25627 13183 25650
rect 13183 25627 13214 25650
rect 13232 25627 13255 25650
rect 13255 25627 13284 25650
rect 13302 25627 13327 25650
rect 13327 25627 13354 25650
rect 13372 25627 13399 25650
rect 13399 25627 13424 25650
rect 13442 25627 13471 25650
rect 13471 25627 13494 25650
rect 13512 25627 13543 25650
rect 13543 25627 13564 25650
rect 13582 25627 13615 25650
rect 13615 25627 13634 25650
rect 13022 25598 13074 25627
rect 13092 25598 13144 25627
rect 13162 25598 13214 25627
rect 13232 25598 13284 25627
rect 13302 25598 13354 25627
rect 13372 25598 13424 25627
rect 13442 25598 13494 25627
rect 13512 25598 13564 25627
rect 13582 25598 13634 25627
rect 13652 25627 13653 25650
rect 13653 25627 13687 25650
rect 13687 25627 13704 25650
rect 13652 25598 13704 25627
rect 13022 25554 13039 25582
rect 13039 25554 13074 25582
rect 13092 25554 13111 25582
rect 13111 25554 13144 25582
rect 13162 25554 13183 25582
rect 13183 25554 13214 25582
rect 13232 25554 13255 25582
rect 13255 25554 13284 25582
rect 13302 25554 13327 25582
rect 13327 25554 13354 25582
rect 13372 25554 13399 25582
rect 13399 25554 13424 25582
rect 13442 25554 13471 25582
rect 13471 25554 13494 25582
rect 13512 25554 13543 25582
rect 13543 25554 13564 25582
rect 13582 25554 13615 25582
rect 13615 25554 13634 25582
rect 13022 25530 13074 25554
rect 13092 25530 13144 25554
rect 13162 25530 13214 25554
rect 13232 25530 13284 25554
rect 13302 25530 13354 25554
rect 13372 25530 13424 25554
rect 13442 25530 13494 25554
rect 13512 25530 13564 25554
rect 13582 25530 13634 25554
rect 13652 25554 13653 25582
rect 13653 25554 13687 25582
rect 13687 25554 13704 25582
rect 13652 25530 13704 25554
rect 13022 25481 13039 25514
rect 13039 25481 13074 25514
rect 13092 25481 13111 25514
rect 13111 25481 13144 25514
rect 13162 25481 13183 25514
rect 13183 25481 13214 25514
rect 13232 25481 13255 25514
rect 13255 25481 13284 25514
rect 13302 25481 13327 25514
rect 13327 25481 13354 25514
rect 13372 25481 13399 25514
rect 13399 25481 13424 25514
rect 13442 25481 13471 25514
rect 13471 25481 13494 25514
rect 13512 25481 13543 25514
rect 13543 25481 13564 25514
rect 13582 25481 13615 25514
rect 13615 25481 13634 25514
rect 13022 25462 13074 25481
rect 13092 25462 13144 25481
rect 13162 25462 13214 25481
rect 13232 25462 13284 25481
rect 13302 25462 13354 25481
rect 13372 25462 13424 25481
rect 13442 25462 13494 25481
rect 13512 25462 13564 25481
rect 13582 25462 13634 25481
rect 13652 25481 13653 25514
rect 13653 25481 13687 25514
rect 13687 25481 13704 25514
rect 13652 25462 13704 25481
rect 13022 25442 13074 25446
rect 13092 25442 13144 25446
rect 13162 25442 13214 25446
rect 13232 25442 13284 25446
rect 13302 25442 13354 25446
rect 13372 25442 13424 25446
rect 13442 25442 13494 25446
rect 13512 25442 13564 25446
rect 13582 25442 13634 25446
rect 13022 25408 13039 25442
rect 13039 25408 13074 25442
rect 13092 25408 13111 25442
rect 13111 25408 13144 25442
rect 13162 25408 13183 25442
rect 13183 25408 13214 25442
rect 13232 25408 13255 25442
rect 13255 25408 13284 25442
rect 13302 25408 13327 25442
rect 13327 25408 13354 25442
rect 13372 25408 13399 25442
rect 13399 25408 13424 25442
rect 13442 25408 13471 25442
rect 13471 25408 13494 25442
rect 13512 25408 13543 25442
rect 13543 25408 13564 25442
rect 13582 25408 13615 25442
rect 13615 25408 13634 25442
rect 13022 25394 13074 25408
rect 13092 25394 13144 25408
rect 13162 25394 13214 25408
rect 13232 25394 13284 25408
rect 13302 25394 13354 25408
rect 13372 25394 13424 25408
rect 13442 25394 13494 25408
rect 13512 25394 13564 25408
rect 13582 25394 13634 25408
rect 13652 25442 13704 25446
rect 13652 25408 13653 25442
rect 13653 25408 13687 25442
rect 13687 25408 13704 25442
rect 13652 25394 13704 25408
rect 13022 25369 13074 25378
rect 13092 25369 13144 25378
rect 13162 25369 13214 25378
rect 13232 25369 13284 25378
rect 13302 25369 13354 25378
rect 13372 25369 13424 25378
rect 13442 25369 13494 25378
rect 13512 25369 13564 25378
rect 13582 25369 13634 25378
rect 13022 25335 13039 25369
rect 13039 25335 13074 25369
rect 13092 25335 13111 25369
rect 13111 25335 13144 25369
rect 13162 25335 13183 25369
rect 13183 25335 13214 25369
rect 13232 25335 13255 25369
rect 13255 25335 13284 25369
rect 13302 25335 13327 25369
rect 13327 25335 13354 25369
rect 13372 25335 13399 25369
rect 13399 25335 13424 25369
rect 13442 25335 13471 25369
rect 13471 25335 13494 25369
rect 13512 25335 13543 25369
rect 13543 25335 13564 25369
rect 13582 25335 13615 25369
rect 13615 25335 13634 25369
rect 13022 25326 13074 25335
rect 13092 25326 13144 25335
rect 13162 25326 13214 25335
rect 13232 25326 13284 25335
rect 13302 25326 13354 25335
rect 13372 25326 13424 25335
rect 13442 25326 13494 25335
rect 13512 25326 13564 25335
rect 13582 25326 13634 25335
rect 13652 25369 13704 25378
rect 13652 25335 13653 25369
rect 13653 25335 13687 25369
rect 13687 25335 13704 25369
rect 13652 25326 13704 25335
rect 13022 25296 13074 25310
rect 13092 25296 13144 25310
rect 13162 25296 13214 25310
rect 13232 25296 13284 25310
rect 13302 25296 13354 25310
rect 13372 25296 13424 25310
rect 13442 25296 13494 25310
rect 13512 25296 13564 25310
rect 13582 25296 13634 25310
rect 13022 25262 13039 25296
rect 13039 25262 13074 25296
rect 13092 25262 13111 25296
rect 13111 25262 13144 25296
rect 13162 25262 13183 25296
rect 13183 25262 13214 25296
rect 13232 25262 13255 25296
rect 13255 25262 13284 25296
rect 13302 25262 13327 25296
rect 13327 25262 13354 25296
rect 13372 25262 13399 25296
rect 13399 25262 13424 25296
rect 13442 25262 13471 25296
rect 13471 25262 13494 25296
rect 13512 25262 13543 25296
rect 13543 25262 13564 25296
rect 13582 25262 13615 25296
rect 13615 25262 13634 25296
rect 13022 25258 13074 25262
rect 13092 25258 13144 25262
rect 13162 25258 13214 25262
rect 13232 25258 13284 25262
rect 13302 25258 13354 25262
rect 13372 25258 13424 25262
rect 13442 25258 13494 25262
rect 13512 25258 13564 25262
rect 13582 25258 13634 25262
rect 13652 25296 13704 25310
rect 13652 25262 13653 25296
rect 13653 25262 13687 25296
rect 13687 25262 13704 25296
rect 13652 25258 13704 25262
rect 13022 25223 13074 25242
rect 13092 25223 13144 25242
rect 13162 25223 13214 25242
rect 13232 25223 13284 25242
rect 13302 25223 13354 25242
rect 13372 25223 13424 25242
rect 13442 25223 13494 25242
rect 13512 25223 13564 25242
rect 13582 25223 13634 25242
rect 13022 25190 13039 25223
rect 13039 25190 13074 25223
rect 13092 25190 13111 25223
rect 13111 25190 13144 25223
rect 13162 25190 13183 25223
rect 13183 25190 13214 25223
rect 13232 25190 13255 25223
rect 13255 25190 13284 25223
rect 13302 25190 13327 25223
rect 13327 25190 13354 25223
rect 13372 25190 13399 25223
rect 13399 25190 13424 25223
rect 13442 25190 13471 25223
rect 13471 25190 13494 25223
rect 13512 25190 13543 25223
rect 13543 25190 13564 25223
rect 13582 25190 13615 25223
rect 13615 25190 13634 25223
rect 13652 25223 13704 25242
rect 13652 25190 13653 25223
rect 13653 25190 13687 25223
rect 13687 25190 13704 25223
rect 13022 25150 13074 25174
rect 13092 25150 13144 25174
rect 13162 25150 13214 25174
rect 13232 25150 13284 25174
rect 13302 25150 13354 25174
rect 13372 25150 13424 25174
rect 13442 25150 13494 25174
rect 13512 25150 13564 25174
rect 13582 25150 13634 25174
rect 13022 25122 13039 25150
rect 13039 25122 13074 25150
rect 13092 25122 13111 25150
rect 13111 25122 13144 25150
rect 13162 25122 13183 25150
rect 13183 25122 13214 25150
rect 13232 25122 13255 25150
rect 13255 25122 13284 25150
rect 13302 25122 13327 25150
rect 13327 25122 13354 25150
rect 13372 25122 13399 25150
rect 13399 25122 13424 25150
rect 13442 25122 13471 25150
rect 13471 25122 13494 25150
rect 13512 25122 13543 25150
rect 13543 25122 13564 25150
rect 13582 25122 13615 25150
rect 13615 25122 13634 25150
rect 13652 25150 13704 25174
rect 13652 25122 13653 25150
rect 13653 25122 13687 25150
rect 13687 25122 13704 25150
rect 8497 25022 8549 25074
rect 8561 25022 8613 25074
rect 5806 24937 5858 24989
rect 5870 24937 5922 24989
rect 8433 24958 8485 25010
rect 8497 24958 8549 25010
rect 5953 24857 6005 24909
rect 6017 24857 6069 24909
rect 8497 24857 8549 24909
rect 8561 24857 8613 24909
rect 5390 21988 5506 22104
rect 7582 21994 7698 22110
rect 4973 21800 5089 21916
rect 7760 21803 7940 21919
rect 6821 21659 6873 21711
rect 6885 21659 6937 21711
rect 6949 21659 7001 21711
rect 7013 21659 7065 21711
rect 6821 21593 6873 21645
rect 6885 21593 6937 21645
rect 6949 21593 7001 21645
rect 7013 21593 7065 21645
rect 6821 21527 6873 21579
rect 6885 21527 6937 21579
rect 6949 21527 7001 21579
rect 7013 21527 7065 21579
rect 6821 21461 6873 21513
rect 6885 21461 6937 21513
rect 6949 21461 7001 21513
rect 7013 21461 7065 21513
rect 6821 21395 6873 21447
rect 6885 21395 6937 21447
rect 6949 21395 7001 21447
rect 7013 21395 7065 21447
rect 3009 20732 3189 20848
rect 4524 20732 4640 20848
rect 735 19976 787 20028
rect 799 19976 851 20028
rect 4884 19976 4936 20028
rect 4948 19976 5000 20028
rect 735 19868 787 19920
rect 799 19868 851 19920
rect 4884 19868 4936 19920
rect 4948 19868 5000 19920
rect 9412 19371 9464 19423
rect 9412 19307 9464 19359
rect 9412 19243 9464 19295
rect 9412 19179 9464 19231
rect 9412 19115 9464 19167
rect 9412 19051 9464 19103
rect 9412 18987 9464 19039
rect 9412 18923 9464 18975
rect 9412 18859 9464 18911
rect 9412 18795 9464 18847
rect 9412 18731 9464 18783
rect 9412 18667 9464 18719
rect 9412 18603 9464 18655
rect 6658 18500 6710 18552
rect 6658 18436 6710 18488
rect 6658 18372 6710 18424
rect 6658 18308 6710 18360
rect 9412 18539 9464 18591
rect 9412 18475 9464 18527
rect 9412 18411 9464 18463
rect 9714 19371 9766 19423
rect 9778 19371 9830 19423
rect 9842 19371 9894 19423
rect 9714 19306 9766 19358
rect 9778 19306 9830 19358
rect 9842 19306 9894 19358
rect 9714 19241 9766 19293
rect 9778 19241 9830 19293
rect 9842 19241 9894 19293
rect 9714 19176 9766 19228
rect 9778 19176 9830 19228
rect 9842 19176 9894 19228
rect 9714 19111 9766 19163
rect 9778 19111 9830 19163
rect 9842 19111 9894 19163
rect 9714 19046 9766 19098
rect 9778 19046 9830 19098
rect 9842 19046 9894 19098
rect 9714 18981 9766 19033
rect 9778 18981 9830 19033
rect 9842 18981 9894 19033
rect 9714 18916 9766 18968
rect 9778 18916 9830 18968
rect 9842 18916 9894 18968
rect 9714 18851 9766 18903
rect 9778 18851 9830 18903
rect 9842 18851 9894 18903
rect 9714 18785 9766 18837
rect 9778 18785 9830 18837
rect 9842 18785 9894 18837
rect 9714 18719 9766 18771
rect 9778 18719 9830 18771
rect 9842 18719 9894 18771
rect 9714 18653 9766 18705
rect 9778 18653 9830 18705
rect 9842 18653 9894 18705
rect 9714 18587 9766 18639
rect 9778 18587 9830 18639
rect 9842 18587 9894 18639
rect 9714 18521 9766 18573
rect 9778 18521 9830 18573
rect 9842 18521 9894 18573
rect 9714 18455 9766 18507
rect 9778 18455 9830 18507
rect 9842 18455 9894 18507
rect 9412 18347 9464 18399
rect 9412 18282 9464 18334
rect 9412 18217 9464 18269
rect 9412 18152 9464 18204
rect 3009 18024 3189 18140
rect 6658 17859 6710 17911
rect 6722 17859 6774 17911
rect 13697 17859 13749 17911
rect 13765 17859 13817 17911
rect 14041 17859 14093 17911
rect 14105 17859 14157 17911
rect 5907 17784 5959 17836
rect 5971 17784 6023 17836
rect 13341 17784 13393 17836
rect 13405 17784 13457 17836
rect 13697 17704 13749 17756
rect 13765 17704 13817 17756
rect 1796 17242 1848 17294
rect 1860 17242 1912 17294
rect 1796 17177 1848 17229
rect 1860 17177 1912 17229
rect 1796 17112 1848 17164
rect 1860 17112 1912 17164
rect 1796 17047 1848 17099
rect 1860 17047 1912 17099
rect 1796 16982 1848 17034
rect 1860 16982 1912 17034
rect 1796 16917 1848 16969
rect 1860 16917 1912 16969
rect 1796 16852 1848 16904
rect 1860 16852 1912 16904
rect 1796 16787 1848 16839
rect 1860 16787 1912 16839
rect 1796 16722 1848 16774
rect 1860 16722 1912 16774
rect 1796 16657 1848 16709
rect 1860 16657 1912 16709
rect 1796 16592 1848 16644
rect 1860 16592 1912 16644
rect 1796 16527 1848 16579
rect 1860 16527 1912 16579
rect 1796 16462 1848 16514
rect 1860 16462 1912 16514
rect 1796 16397 1848 16449
rect 1860 16397 1912 16449
rect 1796 16332 1848 16384
rect 1860 16332 1912 16384
rect 1796 16267 1848 16319
rect 1860 16267 1912 16319
rect 1796 16202 1848 16254
rect 1860 16202 1912 16254
rect 1796 16137 1848 16189
rect 1860 16137 1912 16189
rect 1796 16072 1848 16124
rect 1860 16072 1912 16124
rect 1796 16007 1848 16059
rect 1860 16007 1912 16059
rect 1796 15941 1848 15993
rect 1860 15941 1912 15993
rect 1796 15875 1848 15927
rect 1860 15875 1912 15927
rect 1796 15809 1848 15861
rect 1860 15809 1912 15861
rect 1796 15743 1848 15795
rect 1860 15743 1912 15795
rect 1796 15677 1848 15729
rect 1860 15677 1912 15729
rect 1796 15611 1848 15663
rect 1860 15611 1912 15663
rect 1796 15545 1848 15597
rect 1860 15545 1912 15597
rect 1796 15479 1848 15531
rect 1860 15479 1912 15531
rect 1796 15413 1848 15465
rect 1860 15413 1912 15465
rect 1796 15347 1848 15399
rect 1860 15347 1912 15399
rect 1796 15281 1848 15333
rect 1860 15281 1912 15333
rect 1796 15215 1848 15267
rect 1860 15215 1912 15267
rect 1796 15149 1848 15201
rect 1860 15149 1912 15201
rect 1796 15083 1848 15135
rect 1860 15083 1912 15135
rect 1796 15017 1848 15069
rect 1860 15017 1912 15069
rect 1796 14951 1848 15003
rect 1860 14951 1912 15003
rect 9405 11909 9457 11961
rect 9470 11909 9522 11961
rect 9535 11909 9587 11961
rect 9599 11909 9651 11961
rect 1798 11015 1850 11021
rect 1798 10981 1807 11015
rect 1807 10981 1841 11015
rect 1841 10981 1850 11015
rect 1798 10969 1850 10981
rect 1798 10943 1850 10957
rect 1798 10909 1807 10943
rect 1807 10909 1841 10943
rect 1841 10909 1850 10943
rect 1798 10905 1850 10909
rect 1798 10871 1850 10893
rect 1798 10841 1807 10871
rect 1807 10841 1841 10871
rect 1841 10841 1850 10871
rect 1798 10799 1850 10829
rect 1798 10777 1807 10799
rect 1807 10777 1841 10799
rect 1841 10777 1850 10799
rect 1798 10713 1850 10765
rect 1914 11015 1966 11021
rect 1914 10981 1923 11015
rect 1923 10981 1957 11015
rect 1957 10981 1966 11015
rect 1914 10969 1966 10981
rect 1914 10943 1966 10957
rect 1914 10909 1923 10943
rect 1923 10909 1957 10943
rect 1957 10909 1966 10943
rect 1914 10905 1966 10909
rect 1914 10871 1966 10893
rect 1914 10841 1923 10871
rect 1923 10841 1957 10871
rect 1957 10841 1966 10871
rect 1914 10799 1966 10829
rect 1914 10777 1923 10799
rect 1923 10777 1957 10799
rect 1957 10777 1966 10799
rect 1914 10713 1966 10765
rect 12035 10184 12087 10236
rect 12099 10184 12151 10236
rect 12035 10111 12087 10163
rect 12099 10111 12151 10163
rect 12035 10038 12087 10090
rect 12099 10038 12151 10090
rect 12035 9965 12087 10017
rect 12099 9965 12151 10017
rect 12035 9892 12087 9944
rect 12099 9892 12151 9944
rect 12035 9818 12087 9870
rect 12099 9818 12151 9870
rect 12035 9574 12087 9626
rect 12099 9574 12151 9626
rect 12035 9509 12087 9561
rect 12099 9509 12151 9561
rect 12035 9444 12087 9496
rect 12099 9444 12151 9496
rect 12035 9379 12087 9431
rect 12099 9379 12151 9431
rect 12035 9313 12087 9365
rect 12099 9313 12151 9365
rect 12035 9247 12087 9299
rect 12099 9247 12151 9299
rect 12035 9181 12087 9233
rect 12099 9181 12151 9233
rect 3361 8715 3413 8767
rect 3361 8651 3413 8703
rect 12035 8544 12087 8596
rect 12099 8544 12151 8596
rect 12035 8477 12087 8529
rect 12099 8477 12151 8529
rect 12035 8410 12087 8462
rect 12099 8410 12151 8462
rect 12035 8343 12087 8395
rect 12099 8343 12151 8395
rect 12035 8276 12087 8328
rect 12099 8276 12151 8328
rect 12035 7284 12087 7336
rect 12099 7284 12151 7336
rect 12035 7217 12087 7269
rect 12099 7217 12151 7269
rect 12035 7150 12087 7202
rect 12099 7150 12151 7202
rect 12035 7083 12087 7135
rect 12099 7083 12151 7135
rect 12035 7016 12087 7068
rect 12099 7016 12151 7068
rect 5495 6748 5675 6864
rect 6676 6748 6856 6864
rect 7198 6748 7378 6864
rect 12035 6772 12087 6824
rect 12099 6772 12151 6824
rect 12035 6698 12087 6750
rect 12099 6698 12151 6750
rect 12035 6623 12087 6675
rect 12099 6623 12151 6675
rect 12035 6548 12087 6600
rect 12099 6548 12151 6600
rect 12035 6473 12087 6525
rect 12099 6473 12151 6525
rect 12035 5526 12087 5578
rect 12099 5526 12151 5578
rect 12035 5453 12087 5505
rect 12099 5453 12151 5505
rect 12035 5380 12087 5432
rect 12099 5380 12151 5432
rect 12035 5306 12087 5358
rect 12099 5306 12151 5358
rect 3361 5215 3413 5267
rect 3361 5151 3413 5203
rect 12035 4391 12151 4699
rect 12035 4326 12087 4378
rect 12099 4326 12151 4378
rect 12035 4261 12087 4313
rect 12099 4261 12151 4313
rect 12035 4014 12087 4066
rect 12099 4014 12151 4066
rect 12035 3948 12087 4000
rect 12099 3948 12151 4000
rect 12035 3882 12087 3934
rect 12099 3882 12151 3934
rect 12035 3816 12087 3868
rect 12099 3816 12151 3868
rect 12035 3750 12087 3802
rect 12099 3750 12151 3802
rect 12035 3684 12087 3736
rect 12099 3684 12151 3736
rect 1798 3332 1850 3384
rect 1798 3298 1807 3320
rect 1807 3298 1841 3320
rect 1841 3298 1850 3320
rect 1798 3268 1850 3298
rect 1798 3226 1807 3256
rect 1807 3226 1841 3256
rect 1841 3226 1850 3256
rect 1798 3204 1850 3226
rect 1798 3188 1850 3192
rect 1798 3154 1807 3188
rect 1807 3154 1841 3188
rect 1841 3154 1850 3188
rect 1798 3140 1850 3154
rect 1798 3116 1850 3128
rect 1798 3082 1807 3116
rect 1807 3082 1841 3116
rect 1841 3082 1850 3116
rect 1798 3076 1850 3082
rect 1914 3332 1966 3384
rect 1914 3298 1923 3320
rect 1923 3298 1957 3320
rect 1957 3298 1966 3320
rect 1914 3268 1966 3298
rect 1914 3226 1923 3256
rect 1923 3226 1957 3256
rect 1957 3226 1966 3256
rect 1914 3204 1966 3226
rect 1914 3188 1966 3192
rect 1914 3154 1923 3188
rect 1923 3154 1957 3188
rect 1957 3154 1966 3188
rect 1914 3140 1966 3154
rect 1914 3116 1966 3128
rect 1914 3082 1923 3116
rect 1923 3082 1957 3116
rect 1957 3082 1966 3116
rect 1914 3076 1966 3082
rect 4799 2410 4851 2462
rect 4865 2410 4917 2462
rect 4799 2346 4851 2398
rect 4865 2346 4917 2398
rect 8002 2410 8054 2462
rect 8002 2346 8054 2398
rect 8067 2346 8183 2462
rect 4060 2104 4112 2156
rect 4124 2104 4176 2156
rect 4188 2104 4240 2156
rect 5495 2104 5547 2156
rect 5559 2104 5611 2156
rect 5623 2104 5675 2156
rect 6676 2104 6728 2156
rect 6740 2104 6792 2156
rect 6804 2104 6856 2156
rect 7198 2104 7250 2156
rect 7262 2104 7314 2156
rect 7326 2104 7378 2156
rect 8323 2104 8375 2156
rect 8391 2104 8443 2156
rect 8458 2104 8510 2156
rect 8525 2104 8577 2156
rect 10099 1776 10151 1828
rect 10163 1776 10215 1828
rect 10227 1776 10279 1828
rect 10099 1711 10151 1763
rect 10163 1711 10215 1763
rect 10227 1711 10279 1763
rect 10099 1645 10151 1697
rect 10163 1645 10215 1697
rect 10227 1645 10279 1697
rect 11941 1492 11993 1504
rect 12020 1492 12072 1504
rect 12099 1492 12151 1504
rect 11941 1458 11975 1492
rect 11975 1458 11993 1492
rect 12020 1458 12047 1492
rect 12047 1458 12072 1492
rect 12099 1458 12119 1492
rect 12119 1458 12151 1492
rect 11941 1452 11993 1458
rect 12020 1452 12072 1458
rect 12099 1452 12151 1458
rect 4059 1015 4111 1067
rect 4123 1015 4175 1067
rect 4187 1015 4239 1067
rect 4059 949 4111 1001
rect 4123 949 4175 1001
rect 4187 949 4239 1001
rect 4059 883 4111 935
rect 4123 883 4175 935
rect 4187 883 4239 935
rect 5494 1015 5546 1067
rect 5558 1015 5610 1067
rect 5622 1015 5674 1067
rect 5494 949 5546 1001
rect 5558 949 5610 1001
rect 5622 949 5674 1001
rect 5494 883 5546 935
rect 5558 883 5610 935
rect 5622 883 5674 935
rect 6675 1015 6727 1067
rect 6739 1015 6791 1067
rect 6803 1015 6855 1067
rect 6675 949 6727 1001
rect 6739 949 6791 1001
rect 6803 949 6855 1001
rect 6675 883 6727 935
rect 6739 883 6791 935
rect 6803 883 6855 935
rect 7197 1015 7249 1067
rect 7261 1015 7313 1067
rect 7325 1015 7377 1067
rect 7197 949 7249 1001
rect 7261 949 7313 1001
rect 7325 949 7377 1001
rect 8327 1015 8379 1067
rect 8392 1015 8444 1067
rect 8327 951 8379 1003
rect 8392 951 8444 1003
rect 7197 883 7249 935
rect 7261 883 7313 935
rect 7325 883 7377 935
rect 8327 887 8379 939
rect 8392 887 8444 939
rect 8457 887 8573 1067
rect 10099 733 10151 785
rect 10163 733 10215 785
rect 10227 733 10279 785
rect 8002 658 8054 710
rect 4801 587 4853 639
rect 4865 587 4917 639
rect 8002 594 8054 646
rect 8067 594 8183 710
rect 10099 668 10151 720
rect 10163 668 10215 720
rect 10227 668 10279 720
rect 10099 602 10151 654
rect 10163 602 10215 654
rect 10227 602 10279 654
rect 12234 1226 12286 1232
rect 12234 1192 12243 1226
rect 12243 1192 12277 1226
rect 12277 1192 12286 1226
rect 12234 1180 12286 1192
rect 12234 1154 12286 1166
rect 12234 1120 12243 1154
rect 12243 1120 12277 1154
rect 12277 1120 12286 1154
rect 12234 1114 12286 1120
rect 12494 1226 12546 1232
rect 12494 1192 12503 1226
rect 12503 1192 12537 1226
rect 12537 1192 12546 1226
rect 12494 1180 12546 1192
rect 12494 1154 12546 1166
rect 12494 1120 12503 1154
rect 12503 1120 12537 1154
rect 12537 1120 12546 1154
rect 12494 1114 12546 1120
rect 1300 61 1352 113
rect 1366 61 1418 113
rect 1432 61 1484 113
rect 1498 61 1550 113
rect 1564 61 1616 113
rect 1630 61 1682 113
rect 1696 61 1748 113
rect 1762 61 1814 113
rect 1827 61 1879 113
rect 1892 61 1944 113
rect 1957 61 2009 113
rect 2022 61 2074 113
rect 2087 61 2139 113
rect 2152 61 2204 113
rect 2217 61 2269 113
rect 2282 61 2334 113
rect 2347 61 2399 113
rect 4060 61 4112 113
rect 4124 61 4176 113
rect 4188 61 4240 113
rect 5495 61 5547 113
rect 5559 61 5611 113
rect 5623 61 5675 113
rect 6676 61 6728 113
rect 6740 61 6792 113
rect 6804 61 6856 113
rect 7198 61 7250 113
rect 7262 61 7314 113
rect 7326 61 7378 113
rect 8323 61 8375 113
rect 8391 61 8443 113
rect 8458 61 8510 113
rect 8525 61 8577 113
rect 10751 61 10803 113
rect 10819 61 10871 113
rect 10886 61 10938 113
rect 10953 61 11005 113
<< metal2 >>
rect 9307 29935 10256 30075
rect 8147 29863 10433 29895
tri 10433 29863 10465 29895 sw
rect 4678 29857 4796 29863
rect 4678 29805 4679 29857
rect 4731 29805 4743 29857
rect 4795 29805 4796 29857
tri 2076 29541 2092 29557 se
rect 2092 29541 2098 29557
rect 1680 29535 2098 29541
rect 1732 29523 2098 29535
rect 1732 29483 2034 29523
rect 1680 29478 2034 29483
rect 1680 29473 1733 29478
tri 1680 29426 1727 29473 ne
rect 1727 29426 1733 29473
rect 1785 29471 2034 29478
rect 2086 29505 2098 29523
rect 2150 29505 2156 29557
rect 2086 29471 2156 29505
rect 1785 29465 2156 29471
rect 1785 29426 1791 29465
tri 1791 29426 1830 29465 nw
tri 1815 29410 1821 29416 se
rect 1821 29410 2150 29416
tri 1803 29398 1815 29410 se
rect 1815 29398 2098 29410
rect 1680 29392 2098 29398
rect 1732 29366 2098 29392
rect 1732 29358 1865 29366
tri 1865 29358 1873 29366 nw
tri 2073 29358 2081 29366 ne
rect 2081 29358 2098 29366
rect 1732 29346 1853 29358
tri 1853 29346 1865 29358 nw
tri 2081 29346 2093 29358 ne
rect 2093 29346 2150 29358
rect 1732 29340 1844 29346
rect 1680 29337 1844 29340
tri 1844 29337 1853 29346 nw
tri 2093 29341 2098 29346 ne
rect 1680 29333 1734 29337
tri 1680 29285 1728 29333 ne
rect 1728 29285 1734 29333
rect 1786 29294 1801 29337
tri 1801 29294 1844 29337 nw
rect 1786 29288 1795 29294
tri 1795 29288 1801 29294 nw
rect 2098 29288 2150 29294
rect 1786 29285 1792 29288
tri 1792 29285 1795 29288 nw
rect -13399 29062 -12677 29204
tri 4663 21711 4678 21726 se
rect 4678 21711 4796 29805
rect 5097 29857 5213 29863
rect 5149 29805 5161 29857
tri 4611 21659 4663 21711 se
rect 4663 21678 4796 21711
rect 4663 21659 4777 21678
tri 4777 21659 4796 21678 nw
tri 4973 24370 5097 24494 se
rect 5097 24453 5213 29805
rect 5097 24370 5130 24453
tri 5130 24370 5213 24453 nw
rect 5243 29857 5359 29863
rect 5295 29805 5307 29857
rect 5243 24453 5359 29805
rect 8147 29767 10465 29863
tri 10372 29739 10400 29767 ne
rect 10400 29739 10465 29767
tri 10465 29739 10589 29863 sw
rect 8928 29733 8980 29739
rect 8928 29669 8980 29681
rect 7558 29505 7564 29557
rect 7616 29505 7628 29557
rect 7680 29505 8004 29557
rect 8056 29505 8068 29557
rect 8120 29505 8126 29557
rect 7558 29416 7564 29468
rect 7616 29416 7628 29468
rect 7680 29416 8004 29468
rect 8056 29416 8068 29468
rect 8120 29416 8126 29468
tri 8893 25135 8928 25170 se
rect 8928 25148 8980 29617
rect 8928 25135 8954 25148
rect 5799 24937 5806 24989
rect 5858 24937 5870 24989
rect 5922 24937 5928 24989
tri 5243 24370 5326 24453 ne
rect 5326 24370 5359 24453
rect 4973 24358 5118 24370
tri 5118 24358 5130 24370 nw
tri 5326 24358 5338 24370 ne
rect 5338 24358 5359 24370
tri 5359 24358 5506 24505 sw
rect 4973 24337 5097 24358
tri 5097 24337 5118 24358 nw
tri 5338 24337 5359 24358 ne
rect 5359 24337 5506 24358
rect 4973 21916 5089 24337
tri 5089 24329 5097 24337 nw
tri 5359 24329 5367 24337 ne
rect 5367 24329 5506 24337
tri 5367 24306 5390 24329 ne
rect 5390 22104 5506 24329
rect 5390 21982 5506 21988
tri 4597 21645 4611 21659 se
rect 4611 21645 4763 21659
tri 4763 21645 4777 21659 nw
tri 4545 21593 4597 21645 se
rect 4597 21593 4711 21645
tri 4711 21593 4763 21645 nw
tri 4531 21579 4545 21593 se
rect 4545 21579 4697 21593
tri 4697 21579 4711 21593 nw
tri 4518 21566 4531 21579 se
rect 4531 21566 4684 21579
tri 4684 21566 4697 21579 nw
rect 4518 20848 4646 21566
tri 4646 21528 4684 21566 nw
tri 4964 21513 4973 21522 se
rect 4973 21513 5089 21800
tri 5738 21711 5799 21772 se
rect 5799 21750 5851 24937
tri 5851 24912 5876 24937 nw
rect 5947 24857 5953 24909
rect 6005 24857 6017 24909
rect 6069 24857 6075 24909
tri 5998 24832 6023 24857 ne
rect 5799 21711 5812 21750
tri 5812 21711 5851 21750 nw
tri 5949 21717 6023 21791 se
rect 6023 21769 6075 24857
tri 6023 21717 6075 21769 nw
tri 5943 21711 5949 21717 se
rect 5949 21711 6017 21717
tri 6017 21711 6023 21717 nw
tri 5725 21698 5738 21711 se
rect 5738 21698 5799 21711
tri 5799 21698 5812 21711 nw
tri 5930 21698 5943 21711 se
rect 5943 21698 5996 21711
tri 5717 21690 5725 21698 se
rect 5725 21690 5791 21698
tri 5791 21690 5799 21698 nw
tri 5922 21690 5930 21698 se
rect 5930 21690 5996 21698
tri 5996 21690 6017 21711 nw
tri 5686 21659 5717 21690 se
rect 5717 21659 5760 21690
tri 5760 21659 5791 21690 nw
tri 5891 21659 5922 21690 se
rect 5922 21659 5965 21690
tri 5965 21659 5996 21690 nw
tri 6128 21659 6159 21690 se
rect 6159 21659 6419 24546
tri 5672 21645 5686 21659 se
rect 5686 21645 5746 21659
tri 5746 21645 5760 21659 nw
tri 5877 21645 5891 21659 se
rect 5891 21645 5951 21659
tri 5951 21645 5965 21659 nw
tri 6114 21645 6128 21659 se
rect 6128 21645 6419 21659
tri 5651 21624 5672 21645 se
rect 5672 21624 5725 21645
tri 5725 21624 5746 21645 nw
tri 5875 21643 5877 21645 se
rect 5877 21643 5949 21645
tri 5949 21643 5951 21645 nw
tri 6112 21643 6114 21645 se
rect 6114 21643 6419 21645
tri 5856 21624 5875 21643 se
rect 5875 21624 5899 21643
tri 5620 21593 5651 21624 se
rect 5651 21593 5694 21624
tri 5694 21593 5725 21624 nw
tri 5825 21593 5856 21624 se
rect 5856 21593 5899 21624
tri 5899 21593 5949 21643 nw
tri 6062 21593 6112 21643 se
rect 6112 21593 6419 21643
tri 5606 21579 5620 21593 se
rect 5620 21579 5680 21593
tri 5680 21579 5694 21593 nw
tri 5811 21579 5825 21593 se
rect 5825 21579 5885 21593
tri 5885 21579 5899 21593 nw
tri 6048 21579 6062 21593 se
rect 6062 21582 6419 21593
rect 6062 21579 6416 21582
tri 6416 21579 6419 21582 nw
rect 6814 21711 7070 25135
tri 8880 25122 8893 25135 se
rect 8893 25122 8954 25135
tri 8954 25122 8980 25148 nw
rect 9008 29733 9060 29739
tri 10400 29730 10409 29739 ne
rect 10409 29730 10589 29739
tri 10589 29730 10598 29739 sw
tri 10409 29706 10433 29730 ne
rect 10433 29706 10598 29730
rect 9008 29669 9060 29681
tri 10433 29669 10470 29706 ne
tri 8854 25096 8880 25122 se
rect 8880 25096 8928 25122
tri 8928 25096 8954 25122 nw
tri 8832 25074 8854 25096 se
rect 8854 25074 8906 25096
tri 8906 25074 8928 25096 nw
tri 9005 25074 9008 25077 se
rect 9008 25074 9060 29617
rect 10470 27776 10598 29706
tri 10470 27775 10471 27776 ne
rect 10471 27775 10598 27776
tri 10598 27775 10613 27790 sw
tri 10471 27648 10598 27775 ne
rect 10598 27648 10613 27775
tri 10598 27633 10613 27648 ne
tri 10613 27633 10755 27775 sw
tri 10613 27556 10690 27633 ne
rect 10690 27563 10755 27633
tri 10755 27563 10825 27633 sw
rect 10690 27556 10825 27563
tri 10825 27556 10832 27563 sw
rect 14800 27556 15258 27563
tri 10690 27491 10755 27556 ne
rect 10755 27491 10832 27556
tri 10832 27491 10897 27556 sw
rect 14800 27554 14820 27556
rect 15256 27554 15258 27556
rect 14800 27498 14801 27554
rect 15257 27498 15258 27554
tri 10755 27349 10897 27491 ne
tri 10897 27349 11039 27491 sw
tri 10897 27335 10911 27349 ne
tri 8439 25022 8491 25074 se
rect 8491 25022 8497 25074
rect 8549 25022 8561 25074
rect 8613 25022 8854 25074
tri 8854 25022 8906 25074 nw
tri 8953 25022 9005 25074 se
rect 9005 25055 9060 25074
rect 9005 25022 9008 25055
tri 8427 25010 8439 25022 se
rect 8439 25010 8607 25022
tri 8607 25010 8619 25022 nw
tri 8941 25010 8953 25022 se
rect 8953 25010 9008 25022
rect 8427 24958 8433 25010
rect 8485 24958 8497 25010
rect 8549 24958 8555 25010
tri 8555 24958 8607 25010 nw
tri 8934 25003 8941 25010 se
rect 8941 25003 9008 25010
tri 9008 25003 9060 25055 nw
tri 8889 24958 8934 25003 se
tri 8860 24929 8889 24958 se
rect 8889 24929 8934 24958
tri 8934 24929 9008 25003 nw
tri 8840 24909 8860 24929 se
rect 8860 24909 8914 24929
tri 8914 24909 8934 24929 nw
rect 8491 24857 8497 24909
rect 8549 24857 8561 24909
rect 8613 24857 8862 24909
tri 8862 24857 8914 24909 nw
rect 10911 23217 11039 27349
rect 14800 27411 14820 27498
rect 15256 27411 15258 27498
rect 14800 27355 14801 27411
rect 15257 27355 15258 27411
rect 14800 27268 14820 27355
rect 15256 27268 15258 27355
rect 14800 27212 14801 27268
rect 15257 27212 15258 27268
rect 14800 27125 14820 27212
rect 15256 27125 15258 27212
rect 14800 27069 14801 27125
rect 15257 27069 15258 27125
rect 14800 26992 14820 27069
rect 15256 26992 15258 27069
rect 14800 26981 15258 26992
rect 13017 26973 13709 26976
rect 13017 26921 13024 26973
rect 13076 26955 13093 26973
rect 13145 26955 13162 26973
rect 13214 26955 13231 26973
rect 13283 26955 13300 26973
rect 13085 26921 13093 26955
rect 13283 26921 13293 26955
rect 13352 26921 13369 26973
rect 13421 26955 13439 26973
rect 13491 26955 13509 26973
rect 13561 26955 13579 26973
rect 13631 26955 13649 26973
rect 13437 26921 13439 26955
rect 13631 26921 13645 26955
rect 13017 26909 13029 26921
rect 13085 26909 13117 26921
rect 13173 26909 13205 26921
rect 13261 26909 13293 26921
rect 13349 26909 13381 26921
rect 13437 26909 13469 26921
rect 13525 26909 13557 26921
rect 13613 26909 13645 26921
rect 13017 26857 13024 26909
rect 13085 26899 13093 26909
rect 13283 26899 13293 26909
rect 13076 26875 13093 26899
rect 13145 26875 13162 26899
rect 13214 26875 13231 26899
rect 13283 26875 13300 26899
rect 13085 26857 13093 26875
rect 13283 26857 13293 26875
rect 13352 26857 13369 26909
rect 13437 26899 13439 26909
rect 13631 26899 13645 26909
rect 13421 26875 13439 26899
rect 13491 26875 13509 26899
rect 13561 26875 13579 26899
rect 13631 26875 13649 26899
rect 13437 26857 13439 26875
rect 13631 26857 13645 26875
rect 13017 26845 13029 26857
rect 13085 26845 13117 26857
rect 13173 26845 13205 26857
rect 13261 26845 13293 26857
rect 13349 26845 13381 26857
rect 13437 26845 13469 26857
rect 13525 26845 13557 26857
rect 13613 26845 13645 26857
rect 13017 26793 13024 26845
rect 13085 26819 13093 26845
rect 13283 26819 13293 26845
rect 13076 26795 13093 26819
rect 13145 26795 13162 26819
rect 13214 26795 13231 26819
rect 13283 26795 13300 26819
rect 13085 26793 13093 26795
rect 13283 26793 13293 26795
rect 13352 26793 13369 26845
rect 13437 26819 13439 26845
rect 13631 26819 13645 26845
rect 13421 26795 13439 26819
rect 13491 26795 13509 26819
rect 13561 26795 13579 26819
rect 13631 26795 13649 26819
rect 13437 26793 13439 26795
rect 13631 26793 13645 26795
rect 13017 26781 13029 26793
rect 13085 26781 13117 26793
rect 13173 26781 13205 26793
rect 13261 26781 13293 26793
rect 13349 26781 13381 26793
rect 13437 26781 13469 26793
rect 13525 26781 13557 26793
rect 13613 26781 13645 26793
rect 13017 26729 13024 26781
rect 13085 26739 13093 26781
rect 13283 26739 13293 26781
rect 13076 26729 13093 26739
rect 13145 26729 13162 26739
rect 13214 26729 13231 26739
rect 13283 26729 13300 26739
rect 13352 26729 13369 26781
rect 13437 26739 13439 26781
rect 13631 26739 13645 26781
rect 13421 26729 13439 26739
rect 13491 26729 13509 26739
rect 13561 26729 13579 26739
rect 13631 26729 13649 26739
rect 13701 26729 13709 26973
rect 14800 26925 14801 26981
rect 14857 26979 14901 26981
rect 14957 26979 15001 26981
rect 15057 26979 15101 26981
rect 15157 26979 15201 26981
rect 14872 26927 14884 26979
rect 15000 26927 15001 26979
rect 15064 26927 15076 26979
rect 15192 26927 15201 26979
rect 14857 26925 14901 26927
rect 14957 26925 15001 26927
rect 15057 26925 15101 26927
rect 15157 26925 15201 26927
rect 15257 26925 15258 26981
rect 14800 26916 15258 26925
rect 13017 26715 13709 26729
rect 13017 26659 13029 26715
rect 13085 26659 13117 26715
rect 13173 26659 13205 26715
rect 13261 26659 13293 26715
rect 13349 26659 13381 26715
rect 13437 26659 13469 26715
rect 13525 26659 13557 26715
rect 13613 26659 13645 26715
rect 13701 26659 13709 26715
rect 13017 26635 13709 26659
rect 13017 26579 13029 26635
rect 13085 26579 13117 26635
rect 13173 26579 13205 26635
rect 13261 26579 13293 26635
rect 13349 26579 13381 26635
rect 13437 26579 13469 26635
rect 13525 26579 13557 26635
rect 13613 26579 13645 26635
rect 13701 26579 13709 26635
rect 13017 26555 13709 26579
rect 13017 26499 13029 26555
rect 13085 26499 13117 26555
rect 13173 26499 13205 26555
rect 13261 26499 13293 26555
rect 13349 26499 13381 26555
rect 13437 26499 13469 26555
rect 13525 26499 13557 26555
rect 13613 26499 13645 26555
rect 13701 26499 13709 26555
rect 13017 26475 13709 26499
rect 13017 26419 13029 26475
rect 13085 26419 13117 26475
rect 13173 26419 13205 26475
rect 13261 26419 13293 26475
rect 13349 26419 13381 26475
rect 13437 26419 13469 26475
rect 13525 26419 13557 26475
rect 13613 26419 13645 26475
rect 13701 26419 13709 26475
rect 13017 26395 13709 26419
rect 13017 26339 13029 26395
rect 13085 26339 13117 26395
rect 13173 26339 13205 26395
rect 13261 26339 13293 26395
rect 13349 26339 13381 26395
rect 13437 26339 13469 26395
rect 13525 26339 13557 26395
rect 13613 26339 13645 26395
rect 13701 26339 13709 26395
rect 13017 26315 13709 26339
rect 13017 26259 13029 26315
rect 13085 26259 13117 26315
rect 13173 26259 13205 26315
rect 13261 26259 13293 26315
rect 13349 26259 13381 26315
rect 13437 26259 13469 26315
rect 13525 26259 13557 26315
rect 13613 26259 13645 26315
rect 13701 26259 13709 26315
rect 13017 26253 13709 26259
rect 13017 26201 13022 26253
rect 13074 26235 13092 26253
rect 13144 26235 13162 26253
rect 13214 26235 13232 26253
rect 13284 26235 13302 26253
rect 13085 26201 13092 26235
rect 13284 26201 13293 26235
rect 13354 26201 13372 26253
rect 13424 26235 13442 26253
rect 13494 26235 13512 26253
rect 13564 26235 13582 26253
rect 13634 26235 13652 26253
rect 13437 26201 13442 26235
rect 13634 26201 13645 26235
rect 13704 26201 13709 26253
rect 13017 26186 13029 26201
rect 13085 26186 13117 26201
rect 13173 26186 13205 26201
rect 13261 26186 13293 26201
rect 13349 26186 13381 26201
rect 13437 26186 13469 26201
rect 13525 26186 13557 26201
rect 13613 26186 13645 26201
rect 13701 26186 13709 26201
rect 13017 26134 13022 26186
rect 13085 26179 13092 26186
rect 13284 26179 13293 26186
rect 13074 26155 13092 26179
rect 13144 26155 13162 26179
rect 13214 26155 13232 26179
rect 13284 26155 13302 26179
rect 13085 26134 13092 26155
rect 13284 26134 13293 26155
rect 13354 26134 13372 26186
rect 13437 26179 13442 26186
rect 13634 26179 13645 26186
rect 13424 26155 13442 26179
rect 13494 26155 13512 26179
rect 13564 26155 13582 26179
rect 13634 26155 13652 26179
rect 13437 26134 13442 26155
rect 13634 26134 13645 26155
rect 13704 26134 13709 26186
rect 13017 26119 13029 26134
rect 13085 26119 13117 26134
rect 13173 26119 13205 26134
rect 13261 26119 13293 26134
rect 13349 26119 13381 26134
rect 13437 26119 13469 26134
rect 13525 26119 13557 26134
rect 13613 26119 13645 26134
rect 13701 26119 13709 26134
rect 13017 26067 13022 26119
rect 13085 26099 13092 26119
rect 13284 26099 13293 26119
rect 13074 26075 13092 26099
rect 13144 26075 13162 26099
rect 13214 26075 13232 26099
rect 13284 26075 13302 26099
rect 13085 26067 13092 26075
rect 13284 26067 13293 26075
rect 13354 26067 13372 26119
rect 13437 26099 13442 26119
rect 13634 26099 13645 26119
rect 13424 26075 13442 26099
rect 13494 26075 13512 26099
rect 13564 26075 13582 26099
rect 13634 26075 13652 26099
rect 13437 26067 13442 26075
rect 13634 26067 13645 26075
rect 13704 26067 13709 26119
rect 13017 26052 13029 26067
rect 13085 26052 13117 26067
rect 13173 26052 13205 26067
rect 13261 26052 13293 26067
rect 13349 26052 13381 26067
rect 13437 26052 13469 26067
rect 13525 26052 13557 26067
rect 13613 26052 13645 26067
rect 13701 26052 13709 26067
rect 13017 26000 13022 26052
rect 13085 26019 13092 26052
rect 13284 26019 13293 26052
rect 13074 26000 13092 26019
rect 13144 26000 13162 26019
rect 13214 26000 13232 26019
rect 13284 26000 13302 26019
rect 13354 26000 13372 26052
rect 13437 26019 13442 26052
rect 13634 26019 13645 26052
rect 13424 26000 13442 26019
rect 13494 26000 13512 26019
rect 13564 26000 13582 26019
rect 13634 26000 13652 26019
rect 13704 26000 13709 26052
rect 13017 25995 13709 26000
rect 13017 25985 13029 25995
rect 13085 25985 13117 25995
rect 13173 25985 13205 25995
rect 13261 25985 13293 25995
rect 13349 25985 13381 25995
rect 13437 25985 13469 25995
rect 13525 25985 13557 25995
rect 13613 25985 13645 25995
rect 13701 25985 13709 25995
rect 13017 25933 13022 25985
rect 13085 25939 13092 25985
rect 13284 25939 13293 25985
rect 13074 25933 13092 25939
rect 13144 25933 13162 25939
rect 13214 25933 13232 25939
rect 13284 25933 13302 25939
rect 13354 25933 13372 25985
rect 13437 25939 13442 25985
rect 13634 25939 13645 25985
rect 13424 25933 13442 25939
rect 13494 25933 13512 25939
rect 13564 25933 13582 25939
rect 13634 25933 13652 25939
rect 13704 25933 13709 25985
rect 13017 25918 13709 25933
rect 13017 25866 13022 25918
rect 13074 25915 13092 25918
rect 13144 25915 13162 25918
rect 13214 25915 13232 25918
rect 13284 25915 13302 25918
rect 13085 25866 13092 25915
rect 13284 25866 13293 25915
rect 13354 25866 13372 25918
rect 13424 25915 13442 25918
rect 13494 25915 13512 25918
rect 13564 25915 13582 25918
rect 13634 25915 13652 25918
rect 13437 25866 13442 25915
rect 13634 25866 13645 25915
rect 13704 25866 13709 25918
rect 13017 25859 13029 25866
rect 13085 25859 13117 25866
rect 13173 25859 13205 25866
rect 13261 25859 13293 25866
rect 13349 25859 13381 25866
rect 13437 25859 13469 25866
rect 13525 25859 13557 25866
rect 13613 25859 13645 25866
rect 13701 25859 13709 25866
rect 13017 25851 13709 25859
rect 13017 25799 13022 25851
rect 13074 25835 13092 25851
rect 13144 25835 13162 25851
rect 13214 25835 13232 25851
rect 13284 25835 13302 25851
rect 13085 25799 13092 25835
rect 13284 25799 13293 25835
rect 13354 25799 13372 25851
rect 13424 25835 13442 25851
rect 13494 25835 13512 25851
rect 13564 25835 13582 25851
rect 13634 25835 13652 25851
rect 13437 25799 13442 25835
rect 13634 25799 13645 25835
rect 13704 25799 13709 25851
rect 13017 25784 13029 25799
rect 13085 25784 13117 25799
rect 13173 25784 13205 25799
rect 13261 25784 13293 25799
rect 13349 25784 13381 25799
rect 13437 25784 13469 25799
rect 13525 25784 13557 25799
rect 13613 25784 13645 25799
rect 13701 25784 13709 25799
rect 13017 25732 13022 25784
rect 13085 25779 13092 25784
rect 13284 25779 13293 25784
rect 13074 25754 13092 25779
rect 13144 25754 13162 25779
rect 13214 25754 13232 25779
rect 13284 25754 13302 25779
rect 13085 25732 13092 25754
rect 13284 25732 13293 25754
rect 13354 25732 13372 25784
rect 13437 25779 13442 25784
rect 13634 25779 13645 25784
rect 13424 25754 13442 25779
rect 13494 25754 13512 25779
rect 13564 25754 13582 25779
rect 13634 25754 13652 25779
rect 13437 25732 13442 25754
rect 13634 25732 13645 25754
rect 13704 25732 13709 25784
rect 13017 25717 13029 25732
rect 13085 25717 13117 25732
rect 13173 25717 13205 25732
rect 13261 25717 13293 25732
rect 13349 25717 13381 25732
rect 13437 25717 13469 25732
rect 13525 25717 13557 25732
rect 13613 25717 13645 25732
rect 13701 25717 13709 25732
rect 13017 25665 13022 25717
rect 13085 25698 13092 25717
rect 13284 25698 13293 25717
rect 13074 25665 13092 25698
rect 13144 25665 13162 25698
rect 13214 25665 13232 25698
rect 13284 25665 13302 25698
rect 13354 25665 13372 25717
rect 13437 25698 13442 25717
rect 13634 25698 13645 25717
rect 13424 25665 13442 25698
rect 13494 25665 13512 25698
rect 13564 25665 13582 25698
rect 13634 25665 13652 25698
rect 13704 25665 13709 25717
rect 13017 25650 13709 25665
rect 13017 25598 13022 25650
rect 13074 25598 13092 25650
rect 13144 25598 13162 25650
rect 13214 25598 13232 25650
rect 13284 25598 13302 25650
rect 13354 25598 13372 25650
rect 13424 25598 13442 25650
rect 13494 25598 13512 25650
rect 13564 25598 13582 25650
rect 13634 25598 13652 25650
rect 13704 25598 13709 25650
rect 13017 25582 13709 25598
rect 13017 25530 13022 25582
rect 13074 25530 13092 25582
rect 13144 25530 13162 25582
rect 13214 25530 13232 25582
rect 13284 25530 13302 25582
rect 13354 25530 13372 25582
rect 13424 25530 13442 25582
rect 13494 25530 13512 25582
rect 13564 25530 13582 25582
rect 13634 25530 13652 25582
rect 13704 25530 13709 25582
rect 13017 25514 13709 25530
rect 13017 25462 13022 25514
rect 13074 25462 13092 25514
rect 13144 25462 13162 25514
rect 13214 25462 13232 25514
rect 13284 25462 13302 25514
rect 13354 25462 13372 25514
rect 13424 25462 13442 25514
rect 13494 25462 13512 25514
rect 13564 25462 13582 25514
rect 13634 25462 13652 25514
rect 13704 25462 13709 25514
rect 13017 25446 13709 25462
rect 13017 25394 13022 25446
rect 13074 25394 13092 25446
rect 13144 25394 13162 25446
rect 13214 25394 13232 25446
rect 13284 25394 13302 25446
rect 13354 25394 13372 25446
rect 13424 25394 13442 25446
rect 13494 25394 13512 25446
rect 13564 25394 13582 25446
rect 13634 25394 13652 25446
rect 13704 25394 13709 25446
rect 13017 25378 13709 25394
rect 13017 25326 13022 25378
rect 13074 25326 13092 25378
rect 13144 25326 13162 25378
rect 13214 25326 13232 25378
rect 13284 25326 13302 25378
rect 13354 25326 13372 25378
rect 13424 25326 13442 25378
rect 13494 25326 13512 25378
rect 13564 25326 13582 25378
rect 13634 25326 13652 25378
rect 13704 25326 13709 25378
rect 13017 25310 13709 25326
rect 13017 25258 13022 25310
rect 13074 25258 13092 25310
rect 13144 25258 13162 25310
rect 13214 25258 13232 25310
rect 13284 25258 13302 25310
rect 13354 25258 13372 25310
rect 13424 25258 13442 25310
rect 13494 25258 13512 25310
rect 13564 25258 13582 25310
rect 13634 25258 13652 25310
rect 13704 25258 13709 25310
rect 13017 25242 13709 25258
rect 13017 25190 13022 25242
rect 13074 25190 13092 25242
rect 13144 25190 13162 25242
rect 13214 25190 13232 25242
rect 13284 25190 13302 25242
rect 13354 25190 13372 25242
rect 13424 25190 13442 25242
rect 13494 25190 13512 25242
rect 13564 25190 13582 25242
rect 13634 25190 13652 25242
rect 13704 25190 13709 25242
rect 13017 25174 13709 25190
rect 13017 25122 13022 25174
rect 13074 25122 13092 25174
rect 13144 25122 13162 25174
rect 13214 25122 13232 25174
rect 13284 25122 13302 25174
rect 13354 25122 13372 25174
rect 13424 25122 13442 25174
rect 13494 25122 13512 25174
rect 13564 25122 13582 25174
rect 13634 25122 13652 25174
rect 13704 25122 13709 25174
rect 13017 25116 13709 25122
tri 10911 23210 10918 23217 ne
rect 10918 23210 11039 23217
tri 11039 23210 11060 23231 sw
tri 10918 23089 11039 23210 ne
rect 11039 23089 11060 23210
tri 11039 23068 11060 23089 ne
tri 11060 23068 11202 23210 sw
tri 11060 22926 11202 23068 ne
tri 11202 22926 11344 23068 sw
tri 11202 22874 11254 22926 ne
rect 11254 22874 13503 22926
tri 13467 22851 13490 22874 ne
rect 13490 22851 13503 22874
tri 13503 22851 13578 22926 sw
tri 13490 22838 13503 22851 ne
rect 13503 22838 13578 22851
tri 13503 22815 13526 22838 ne
rect 6814 21659 6821 21711
rect 6873 21659 6885 21711
rect 6937 21659 6949 21711
rect 7001 21659 7013 21711
rect 7065 21659 7070 21711
rect 6814 21645 7070 21659
rect 6814 21593 6821 21645
rect 6873 21593 6885 21645
rect 6937 21593 6949 21645
rect 7001 21593 7013 21645
rect 7065 21593 7070 21645
rect 6814 21579 7070 21593
tri 5577 21550 5606 21579 se
rect 5606 21550 5651 21579
tri 5651 21550 5680 21579 nw
tri 5801 21569 5811 21579 se
rect 5811 21569 5875 21579
tri 5875 21569 5885 21579 nw
tri 6038 21569 6048 21579 se
rect 6048 21569 6364 21579
tri 5782 21550 5801 21569 se
rect 5801 21550 5833 21569
tri 5554 21527 5577 21550 se
rect 5577 21527 5628 21550
tri 5628 21527 5651 21550 nw
tri 5759 21527 5782 21550 se
rect 5782 21527 5833 21550
tri 5833 21527 5875 21569 nw
tri 5996 21527 6038 21569 se
rect 6038 21527 6364 21569
tri 6364 21527 6416 21579 nw
rect 6814 21527 6821 21579
rect 6873 21527 6885 21579
rect 6937 21527 6949 21579
rect 7001 21527 7013 21579
rect 7065 21527 7070 21579
tri 5540 21513 5554 21527 se
rect 5554 21513 5614 21527
tri 5614 21513 5628 21527 nw
tri 5745 21513 5759 21527 se
rect 5759 21513 5819 21527
tri 5819 21513 5833 21527 nw
tri 5982 21513 5996 21527 se
rect 5996 21513 6350 21527
tri 6350 21513 6364 21527 nw
rect 6814 21513 7070 21527
tri 4912 21461 4964 21513 se
rect 4964 21474 5089 21513
tri 5503 21476 5540 21513 se
rect 5540 21476 5577 21513
tri 5577 21476 5614 21513 nw
tri 5727 21495 5745 21513 se
rect 5745 21495 5801 21513
tri 5801 21495 5819 21513 nw
tri 5964 21495 5982 21513 se
rect 5982 21495 6298 21513
tri 5708 21476 5727 21495 se
rect 5727 21476 5767 21495
rect 4964 21461 5076 21474
tri 5076 21461 5089 21474 nw
tri 5488 21461 5503 21476 se
rect 5503 21461 5562 21476
tri 5562 21461 5577 21476 nw
tri 5693 21461 5708 21476 se
rect 5708 21461 5767 21476
tri 5767 21461 5801 21495 nw
tri 5930 21461 5964 21495 se
rect 5964 21461 6298 21495
tri 6298 21461 6350 21513 nw
rect 6814 21461 6821 21513
rect 6873 21461 6885 21513
rect 6937 21461 6949 21513
rect 7001 21461 7013 21513
rect 7065 21461 7070 21513
tri 4898 21447 4912 21461 se
rect 4912 21447 5062 21461
tri 5062 21447 5076 21461 nw
tri 5474 21447 5488 21461 se
rect 5488 21447 5548 21461
tri 5548 21447 5562 21461 nw
tri 5679 21447 5693 21461 se
rect 5693 21447 5753 21461
tri 5753 21447 5767 21461 nw
tri 5916 21447 5930 21461 se
rect 5930 21447 6284 21461
tri 6284 21447 6298 21461 nw
rect 6814 21447 7070 21461
tri 4846 21395 4898 21447 se
rect 4898 21395 5010 21447
tri 5010 21395 5062 21447 nw
tri 5429 21402 5474 21447 se
rect 5474 21402 5503 21447
tri 5503 21402 5548 21447 nw
tri 5653 21421 5679 21447 se
rect 5679 21421 5727 21447
tri 5727 21421 5753 21447 nw
tri 5890 21421 5916 21447 se
rect 5916 21421 6232 21447
tri 5634 21402 5653 21421 se
rect 5653 21402 5701 21421
tri 5422 21395 5429 21402 se
rect 5429 21395 5496 21402
tri 5496 21395 5503 21402 nw
tri 5627 21395 5634 21402 se
rect 5634 21395 5701 21402
tri 5701 21395 5727 21421 nw
tri 5864 21395 5890 21421 se
rect 5890 21395 6232 21421
tri 6232 21395 6284 21447 nw
rect 6814 21395 6821 21447
rect 6873 21395 6885 21447
rect 6937 21395 6949 21447
rect 7001 21395 7013 21447
rect 7065 21395 7070 21447
tri 4809 21358 4846 21395 se
rect 4846 21358 4973 21395
tri 4973 21358 5010 21395 nw
tri 5416 21389 5422 21395 se
rect 5422 21389 5490 21395
tri 5490 21389 5496 21395 nw
tri 5621 21389 5627 21395 se
rect 5627 21389 5695 21395
tri 5695 21389 5701 21395 nw
tri 5858 21389 5864 21395 se
rect 5864 21389 6226 21395
tri 6226 21389 6232 21395 nw
tri 5385 21358 5416 21389 se
rect 5416 21358 5459 21389
tri 5459 21358 5490 21389 nw
tri 5590 21358 5621 21389 se
rect 5621 21358 5664 21389
tri 5664 21358 5695 21389 nw
tri 5827 21358 5858 21389 se
rect 5858 21358 6159 21389
tri 4734 21283 4809 21358 se
rect 4809 21283 4898 21358
tri 4898 21283 4973 21358 nw
tri 5355 21328 5385 21358 se
rect 5385 21328 5429 21358
tri 5429 21328 5459 21358 nw
tri 5579 21347 5590 21358 se
rect 5590 21347 5653 21358
tri 5653 21347 5664 21358 nw
tri 5816 21347 5827 21358 se
rect 5827 21347 6159 21358
tri 5560 21328 5579 21347 se
rect 5579 21328 5628 21347
tri 5349 21322 5355 21328 se
rect 5355 21322 5423 21328
tri 5423 21322 5429 21328 nw
tri 5554 21322 5560 21328 se
rect 5560 21322 5628 21328
tri 5628 21322 5653 21347 nw
tri 5791 21322 5816 21347 se
rect 5816 21322 6159 21347
tri 6159 21322 6226 21389 nw
tri 5310 21283 5349 21322 se
rect 5349 21283 5384 21322
tri 5384 21283 5423 21322 nw
tri 5515 21283 5554 21322 se
rect 5554 21283 5589 21322
tri 5589 21283 5628 21322 nw
tri 5752 21283 5791 21322 se
rect 5791 21283 5845 21322
rect 4734 20900 4850 21283
tri 4850 21235 4898 21283 nw
tri 5281 21254 5310 21283 se
rect 5310 21254 5355 21283
tri 5355 21254 5384 21283 nw
tri 5505 21273 5515 21283 se
rect 5515 21273 5579 21283
tri 5579 21273 5589 21283 nw
tri 5742 21273 5752 21283 se
rect 5752 21273 5845 21283
tri 5486 21254 5505 21273 se
rect 5505 21254 5541 21273
tri 5262 21235 5281 21254 se
rect 5281 21235 5336 21254
tri 5336 21235 5355 21254 nw
tri 5467 21235 5486 21254 se
rect 5486 21235 5541 21254
tri 5541 21235 5579 21273 nw
tri 5704 21235 5742 21273 se
rect 5742 21235 5845 21273
tri 5207 21180 5262 21235 se
rect 5262 21180 5281 21235
tri 5281 21180 5336 21235 nw
tri 5431 21199 5467 21235 se
rect 5467 21199 5505 21235
tri 5505 21199 5541 21235 nw
tri 5668 21199 5704 21235 se
rect 5704 21199 5845 21235
tri 5412 21180 5431 21199 se
tri 5133 21106 5207 21180 se
tri 5207 21106 5281 21180 nw
tri 5357 21125 5412 21180 se
rect 5412 21125 5431 21180
tri 5431 21125 5505 21199 nw
tri 5594 21125 5668 21199 se
rect 5668 21125 5845 21199
tri 5338 21106 5357 21125 se
tri 5123 21096 5133 21106 se
rect 5133 21096 5197 21106
tri 5197 21096 5207 21106 nw
tri 5328 21096 5338 21106 se
rect 5338 21096 5357 21106
rect 3003 20732 3009 20848
rect 3189 20732 3202 20848
rect 4518 20732 4524 20848
rect 4640 20732 4646 20848
tri 479 19976 531 20028 se
rect 531 19976 735 20028
rect 787 19976 799 20028
rect 851 19976 857 20028
tri 457 19954 479 19976 se
rect 479 19954 531 19976
tri 531 19954 553 19976 nw
tri 423 19920 457 19954 se
rect 457 19920 497 19954
tri 497 19920 531 19954 nw
tri 383 19880 423 19920 se
rect 423 19880 457 19920
tri 457 19880 497 19920 nw
tri 611 19880 651 19920 se
rect 651 19880 735 19920
tri 371 19868 383 19880 se
rect 383 19868 445 19880
tri 445 19868 457 19880 nw
tri 599 19868 611 19880 se
rect 611 19868 735 19880
rect 787 19868 799 19920
rect 851 19868 857 19920
tri 349 19846 371 19868 se
rect 371 19846 423 19868
tri 423 19846 445 19868 nw
tri 577 19846 599 19868 se
rect 599 19846 651 19868
tri 651 19846 673 19868 nw
tri 309 19806 349 19846 se
rect 349 19806 383 19846
tri 383 19806 423 19846 nw
tri 537 19806 577 19846 se
tri 281 19778 309 19806 se
rect 309 19778 355 19806
tri 355 19778 383 19806 nw
tri 509 19778 537 19806 se
rect 537 19778 577 19806
rect 281 19772 349 19778
tri 349 19772 355 19778 nw
tri 503 19772 509 19778 se
rect 509 19772 577 19778
tri 577 19772 651 19846 nw
rect 281 17756 333 19772
tri 333 19756 349 19772 nw
tri 487 19756 503 19772 se
tri 429 19698 487 19756 se
rect 487 19698 503 19756
tri 503 19698 577 19772 nw
tri 373 19642 429 19698 se
rect 429 19642 447 19698
tri 447 19642 503 19698 nw
rect 373 17756 425 19642
tri 425 19620 447 19642 nw
rect 3003 18140 3202 20732
tri 5053 20028 5123 20098 se
rect 5123 20076 5175 21096
tri 5175 21074 5197 21096 nw
tri 5306 21074 5328 21096 se
rect 5328 21074 5357 21096
tri 5283 21051 5306 21074 se
rect 5306 21051 5357 21074
tri 5357 21051 5431 21125 nw
tri 5520 21051 5594 21125 se
rect 5594 21051 5845 21125
rect 5123 20028 5127 20076
tri 5127 20028 5175 20076 nw
tri 5253 21021 5283 21051 se
rect 5283 21021 5327 21051
tri 5327 21021 5357 21051 nw
tri 5490 21021 5520 21051 se
rect 5520 21021 5845 21051
rect 4878 19976 4884 20028
rect 4936 19976 4948 20028
rect 5000 19976 5075 20028
tri 5075 19976 5127 20028 nw
tri 5202 19976 5253 20027 se
rect 5253 20005 5305 21021
tri 5305 20999 5327 21021 nw
tri 5477 21008 5490 21021 se
rect 5490 21008 5845 21021
tri 5845 21008 6159 21322 nw
tri 5180 19954 5202 19976 se
rect 5202 19954 5253 19976
tri 5179 19953 5180 19954 se
rect 5180 19953 5253 19954
tri 5253 19953 5305 20005 nw
tri 5146 19920 5179 19953 se
rect 5179 19920 5220 19953
tri 5220 19920 5253 19953 nw
rect 4878 19868 4884 19920
rect 4936 19868 4948 19920
rect 5000 19868 5168 19920
tri 5168 19868 5220 19920 nw
tri 5473 18269 5477 18273 se
rect 5477 18269 5737 21008
tri 5737 20900 5845 21008 nw
tri 5421 18217 5473 18269 se
rect 5473 18217 5737 18269
tri 5408 18204 5421 18217 se
rect 5421 18204 5737 18217
tri 5356 18152 5408 18204 se
rect 5408 18152 5737 18204
tri 5344 18140 5356 18152 se
rect 5356 18140 5737 18152
rect 3003 18024 3009 18140
rect 3189 18024 3202 18140
tri 5333 18129 5344 18140 se
rect 5344 18129 5737 18140
tri 4795 18024 4900 18129 se
rect 4900 18091 5737 18129
rect 4900 18024 5602 18091
rect 3003 17911 3202 18024
tri 4727 17956 4795 18024 se
rect 4795 17956 5602 18024
tri 5602 17956 5737 18091 nw
rect 6652 18500 6658 18552
rect 6710 18500 6716 18552
rect 6652 18488 6716 18500
rect 6652 18436 6658 18488
rect 6710 18436 6716 18488
rect 6652 18424 6716 18436
rect 6652 18372 6658 18424
rect 6710 18372 6716 18424
rect 6652 18360 6716 18372
rect 6652 18308 6658 18360
rect 6710 18308 6716 18360
tri 3202 17911 3213 17922 sw
rect 4727 17911 5557 17956
tri 5557 17911 5602 17956 nw
rect 6652 17911 6716 18308
rect 6814 17939 7070 21395
rect 7574 21994 7582 22110
rect 7698 21994 7704 22110
tri 6716 17911 6741 17936 sw
rect 3003 17859 3213 17911
tri 3213 17859 3265 17911 sw
rect 4727 17872 5518 17911
tri 5518 17872 5557 17911 nw
rect 4727 17859 5116 17872
tri 5116 17859 5129 17872 nw
rect 6652 17859 6658 17911
rect 6710 17859 6722 17911
rect 6774 17859 6780 17911
rect 3003 17836 3265 17859
tri 3265 17836 3288 17859 sw
rect 4727 17836 5093 17859
tri 5093 17836 5116 17859 nw
tri 2999 17816 3003 17820 se
rect 3003 17816 3288 17836
tri 3288 17816 3308 17836 sw
tri 2967 17784 2999 17816 se
rect 2999 17784 3308 17816
tri 3308 17784 3340 17816 sw
rect 4727 17784 5041 17836
tri 5041 17784 5093 17836 nw
rect 5901 17784 5907 17836
rect 5959 17784 5971 17836
rect 6023 17784 6029 17836
tri 2939 17756 2967 17784 se
rect 2967 17756 3340 17784
tri 3340 17756 3368 17784 sw
rect 1783 17709 2109 17756
tri 2926 17743 2939 17756 se
rect 2939 17743 3368 17756
rect 2926 17697 3368 17743
rect 4727 17756 5013 17784
tri 5013 17756 5041 17784 nw
tri 5952 17759 5977 17784 ne
rect 5977 17756 6029 17784
rect 7574 17756 7704 21994
rect 7760 21919 7940 21954
rect 7760 17756 7940 21803
rect 9399 19423 9905 19429
rect 9399 19371 9412 19423
rect 9464 19371 9714 19423
rect 9766 19371 9778 19423
rect 9830 19371 9842 19423
rect 9894 19371 9905 19423
rect 9399 19359 9905 19371
rect 9399 19307 9412 19359
rect 9464 19358 9905 19359
rect 9464 19307 9714 19358
rect 9399 19306 9714 19307
rect 9766 19306 9778 19358
rect 9830 19306 9842 19358
rect 9894 19306 9905 19358
rect 9399 19295 9905 19306
rect 9399 19243 9412 19295
rect 9464 19293 9905 19295
rect 9464 19243 9714 19293
rect 9399 19241 9714 19243
rect 9766 19241 9778 19293
rect 9830 19241 9842 19293
rect 9894 19241 9905 19293
rect 9399 19231 9905 19241
rect 9399 19179 9412 19231
rect 9464 19228 9905 19231
rect 9464 19179 9714 19228
rect 9399 19176 9714 19179
rect 9766 19176 9778 19228
rect 9830 19176 9842 19228
rect 9894 19176 9905 19228
rect 9399 19167 9905 19176
rect 9399 19115 9412 19167
rect 9464 19163 9905 19167
rect 9464 19115 9714 19163
rect 9399 19111 9714 19115
rect 9766 19111 9778 19163
rect 9830 19111 9842 19163
rect 9894 19111 9905 19163
rect 9399 19103 9905 19111
rect 9399 19051 9412 19103
rect 9464 19098 9905 19103
rect 9464 19051 9714 19098
rect 9399 19046 9714 19051
rect 9766 19046 9778 19098
rect 9830 19046 9842 19098
rect 9894 19046 9905 19098
rect 9399 19039 9905 19046
rect 9399 18987 9412 19039
rect 9464 19033 9905 19039
rect 9464 18987 9714 19033
rect 9399 18981 9714 18987
rect 9766 18981 9778 19033
rect 9830 18981 9842 19033
rect 9894 18981 9905 19033
rect 9399 18975 9905 18981
rect 9399 18923 9412 18975
rect 9464 18968 9905 18975
rect 9464 18923 9714 18968
rect 9399 18916 9714 18923
rect 9766 18916 9778 18968
rect 9830 18916 9842 18968
rect 9894 18916 9905 18968
rect 9399 18911 9905 18916
rect 9399 18859 9412 18911
rect 9464 18903 9905 18911
rect 9464 18859 9714 18903
rect 9399 18851 9714 18859
rect 9766 18851 9778 18903
rect 9830 18851 9842 18903
rect 9894 18851 9905 18903
rect 9399 18847 9905 18851
rect 9399 18795 9412 18847
rect 9464 18837 9905 18847
rect 9464 18795 9714 18837
rect 9399 18785 9714 18795
rect 9766 18785 9778 18837
rect 9830 18785 9842 18837
rect 9894 18785 9905 18837
rect 9399 18783 9905 18785
rect 9399 18731 9412 18783
rect 9464 18771 9905 18783
rect 9464 18731 9714 18771
rect 9399 18719 9714 18731
rect 9766 18719 9778 18771
rect 9830 18719 9842 18771
rect 9894 18719 9905 18771
rect 9399 18667 9412 18719
rect 9464 18705 9905 18719
rect 9464 18667 9714 18705
rect 9399 18655 9714 18667
rect 9399 18603 9412 18655
rect 9464 18653 9714 18655
rect 9766 18653 9778 18705
rect 9830 18653 9842 18705
rect 9894 18653 9905 18705
rect 9464 18639 9905 18653
rect 9464 18603 9714 18639
rect 9399 18591 9714 18603
rect 9399 18539 9412 18591
rect 9464 18587 9714 18591
rect 9766 18587 9778 18639
rect 9830 18587 9842 18639
rect 9894 18587 9905 18639
rect 9464 18573 9905 18587
rect 9464 18539 9714 18573
rect 9399 18527 9714 18539
rect 9399 18475 9412 18527
rect 9464 18521 9714 18527
rect 9766 18521 9778 18573
rect 9830 18521 9842 18573
rect 9894 18521 9905 18573
rect 9464 18507 9905 18521
rect 9464 18475 9714 18507
rect 9399 18463 9714 18475
rect 9399 18411 9412 18463
rect 9464 18455 9714 18463
rect 9766 18455 9778 18507
rect 9830 18455 9842 18507
rect 9894 18455 9905 18507
rect 9464 18411 9905 18455
rect 9399 18399 9905 18411
rect 9399 18347 9412 18399
rect 9464 18354 9905 18399
rect 9464 18347 9859 18354
rect 9399 18334 9859 18347
tri 8733 18282 8768 18317 se
rect 8768 18282 9024 18317
tri 8720 18269 8733 18282 se
rect 8733 18269 9024 18282
tri 8668 18217 8720 18269 se
rect 8720 18217 9024 18269
tri 8655 18204 8668 18217 se
rect 8668 18204 9024 18217
tri 8603 18152 8655 18204 se
rect 8655 18198 9024 18204
rect 8655 18152 8978 18198
tri 8978 18152 9024 18198 nw
rect 9399 18282 9412 18334
rect 9464 18308 9859 18334
tri 9859 18308 9905 18354 nw
rect 9464 18282 9691 18308
rect 9399 18269 9691 18282
rect 9399 18217 9412 18269
rect 9464 18217 9691 18269
rect 9399 18204 9691 18217
rect 9399 18152 9412 18204
rect 9464 18152 9691 18204
tri 8393 17942 8603 18152 se
rect 8603 17942 8768 18152
tri 8768 17942 8978 18152 nw
rect 9399 18140 9691 18152
tri 9691 18140 9859 18308 nw
tri 8362 17911 8393 17942 se
rect 8393 17911 8737 17942
tri 8737 17911 8768 17942 nw
tri 8317 17866 8362 17911 se
rect 8362 17866 8692 17911
tri 8692 17866 8737 17911 nw
rect 8317 17859 8685 17866
tri 8685 17859 8692 17866 nw
rect 8317 17836 8662 17859
tri 8662 17836 8685 17859 nw
rect 8317 17784 8610 17836
tri 8610 17784 8662 17836 nw
rect 4727 17730 4987 17756
tri 4987 17730 5013 17756 nw
rect 5170 17710 5430 17756
rect 7996 17704 8189 17756
rect 8317 17710 8582 17784
tri 8582 17756 8610 17784 nw
rect 9399 17710 9657 18140
tri 9657 18106 9691 18140 nw
rect 10093 17710 10286 21170
rect 12346 18308 12453 18395
tri 12453 18308 12540 18395 sw
rect 12346 18140 12540 18308
tri 12540 18140 12708 18308 sw
rect 12346 18109 12708 18140
tri 12708 18109 12739 18140 sw
rect 12966 18136 13248 18370
tri 13519 18166 13526 18173 se
rect 13526 18166 13578 22838
rect 13519 18151 13578 18166
rect 12966 18109 13221 18136
tri 13221 18109 13248 18136 nw
rect 12346 18047 12739 18109
tri 12739 18047 12801 18109 sw
tri 12904 18047 12966 18109 se
rect 12966 18047 13159 18109
tri 13159 18047 13221 18109 nw
rect 13335 18091 13463 18143
tri 13335 18047 13379 18091 ne
rect 13379 18047 13463 18091
rect 12346 18024 13136 18047
tri 13136 18024 13159 18047 nw
tri 13379 18024 13402 18047 ne
rect 13402 18024 13463 18047
rect 12346 17989 13101 18024
tri 13101 17989 13136 18024 nw
tri 13402 18015 13411 18024 ne
tri 12346 17911 12424 17989 ne
rect 12424 17911 13023 17989
tri 13023 17911 13101 17989 nw
tri 12424 17859 12476 17911 ne
rect 12476 17859 12971 17911
tri 12971 17859 13023 17911 nw
tri 13409 17859 13411 17861 se
rect 13411 17859 13463 18024
tri 12476 17836 12499 17859 ne
rect 12499 17836 12948 17859
tri 12948 17836 12971 17859 nw
tri 13386 17836 13409 17859 se
rect 13409 17836 13463 17859
tri 12499 17784 12551 17836 ne
rect 12551 17784 12896 17836
tri 12896 17784 12948 17836 nw
rect 13335 17784 13341 17836
rect 13393 17784 13405 17836
rect 13457 17784 13463 17836
tri 12551 17756 12579 17784 ne
rect 12579 17756 12868 17784
tri 12868 17756 12896 17784 nw
rect 13519 17756 13571 18151
tri 13571 18144 13578 18151 nw
rect 13691 17859 13697 17911
rect 13749 17859 13765 17911
rect 13817 17859 13823 17911
rect 14026 17859 14041 17911
rect 14093 17859 14105 17911
rect 14157 17859 14170 17911
tri 13691 17836 13714 17859 ne
rect 13714 17836 13792 17859
tri 13792 17836 13815 17859 nw
tri 13714 17825 13725 17836 ne
tri 13719 17784 13725 17790 se
rect 13725 17784 13781 17836
tri 13781 17825 13792 17836 nw
tri 13781 17784 13787 17790 sw
tri 13691 17756 13719 17784 se
rect 13719 17756 13787 17784
tri 13787 17756 13815 17784 sw
rect 12801 17730 12842 17756
tri 12842 17730 12868 17756 nw
rect 12801 17704 12816 17730
tri 12816 17704 12842 17730 nw
rect 13691 17704 13697 17756
rect 13749 17704 13765 17756
rect 13817 17704 13823 17756
rect 12801 17697 12809 17704
tri 12809 17697 12816 17704 nw
tri 12801 17689 12809 17697 nw
rect 14026 17621 14170 17859
rect 14250 17616 14378 17756
rect 14436 17616 14564 17756
rect 1789 17294 1919 17300
rect 1789 17242 1796 17294
rect 1848 17242 1860 17294
rect 1912 17242 1919 17294
rect 1789 17229 1919 17242
rect 1789 17177 1796 17229
rect 1848 17177 1860 17229
rect 1912 17177 1919 17229
rect 1789 17164 1919 17177
rect 1789 17112 1796 17164
rect 1848 17112 1860 17164
rect 1912 17112 1919 17164
rect 1789 17099 1919 17112
rect 1789 17047 1796 17099
rect 1848 17047 1860 17099
rect 1912 17047 1919 17099
rect 1789 17034 1919 17047
rect 1789 16982 1796 17034
rect 1848 16982 1860 17034
rect 1912 16982 1919 17034
rect 1789 16969 1919 16982
rect 1789 16917 1796 16969
rect 1848 16917 1860 16969
rect 1912 16917 1919 16969
rect 1789 16904 1919 16917
rect 1789 16852 1796 16904
rect 1848 16852 1860 16904
rect 1912 16852 1919 16904
rect 1789 16839 1919 16852
rect 1789 16787 1796 16839
rect 1848 16787 1860 16839
rect 1912 16787 1919 16839
rect 1789 16774 1919 16787
rect 1789 16722 1796 16774
rect 1848 16722 1860 16774
rect 1912 16722 1919 16774
rect 1789 16709 1919 16722
rect 1789 16657 1796 16709
rect 1848 16657 1860 16709
rect 1912 16657 1919 16709
rect 1789 16644 1919 16657
rect 1789 16592 1796 16644
rect 1848 16592 1860 16644
rect 1912 16592 1919 16644
rect 1789 16579 1919 16592
rect 1789 16527 1796 16579
rect 1848 16527 1860 16579
rect 1912 16527 1919 16579
rect 1789 16514 1919 16527
rect 1789 16462 1796 16514
rect 1848 16462 1860 16514
rect 1912 16462 1919 16514
rect 1789 16449 1919 16462
rect 1789 16397 1796 16449
rect 1848 16397 1860 16449
rect 1912 16397 1919 16449
rect 1789 16384 1919 16397
rect 1789 16332 1796 16384
rect 1848 16332 1860 16384
rect 1912 16332 1919 16384
rect 1789 16319 1919 16332
rect 1789 16267 1796 16319
rect 1848 16267 1860 16319
rect 1912 16267 1919 16319
rect 1789 16254 1919 16267
rect 1789 16202 1796 16254
rect 1848 16202 1860 16254
rect 1912 16202 1919 16254
rect 1789 16189 1919 16202
rect 1789 16137 1796 16189
rect 1848 16137 1860 16189
rect 1912 16137 1919 16189
rect 1789 16124 1919 16137
rect 1789 16072 1796 16124
rect 1848 16072 1860 16124
rect 1912 16072 1919 16124
rect 1789 16059 1919 16072
rect 1789 16007 1796 16059
rect 1848 16007 1860 16059
rect 1912 16007 1919 16059
rect 1789 15993 1919 16007
rect 1789 15941 1796 15993
rect 1848 15941 1860 15993
rect 1912 15941 1919 15993
rect 1789 15927 1919 15941
rect 1789 15875 1796 15927
rect 1848 15875 1860 15927
rect 1912 15875 1919 15927
rect 1789 15861 1919 15875
rect 1789 15809 1796 15861
rect 1848 15809 1860 15861
rect 1912 15809 1919 15861
rect 1789 15795 1919 15809
rect 1789 15743 1796 15795
rect 1848 15743 1860 15795
rect 1912 15743 1919 15795
rect 1789 15729 1919 15743
rect 1789 15677 1796 15729
rect 1848 15677 1860 15729
rect 1912 15677 1919 15729
rect 1789 15663 1919 15677
rect 1789 15611 1796 15663
rect 1848 15611 1860 15663
rect 1912 15611 1919 15663
rect 1789 15597 1919 15611
rect 1789 15545 1796 15597
rect 1848 15545 1860 15597
rect 1912 15545 1919 15597
rect 1789 15531 1919 15545
rect 1789 15479 1796 15531
rect 1848 15479 1860 15531
rect 1912 15479 1919 15531
rect 1789 15465 1919 15479
rect 1789 15413 1796 15465
rect 1848 15413 1860 15465
rect 1912 15413 1919 15465
rect 1789 15399 1919 15413
rect 1789 15347 1796 15399
rect 1848 15347 1860 15399
rect 1912 15347 1919 15399
rect 1789 15333 1919 15347
rect 1789 15281 1796 15333
rect 1848 15281 1860 15333
rect 1912 15281 1919 15333
rect 1789 15267 1919 15281
rect 1789 15215 1796 15267
rect 1848 15215 1860 15267
rect 1912 15215 1919 15267
rect 1789 15201 1919 15215
rect 1789 15149 1796 15201
rect 1848 15149 1860 15201
rect 1912 15149 1919 15201
rect 1789 15135 1919 15149
rect 1789 15083 1796 15135
rect 1848 15083 1860 15135
rect 1912 15083 1919 15135
rect 1789 15069 1919 15083
rect 1789 15017 1796 15069
rect 1848 15017 1860 15069
rect 1912 15017 1919 15069
rect 1789 15003 1919 15017
rect 1789 14951 1796 15003
rect 1848 14951 1860 15003
rect 1912 14951 1919 15003
rect 1789 14945 1919 14951
rect 9399 11961 9657 11987
rect 9399 11909 9405 11961
rect 9457 11909 9470 11961
rect 9522 11909 9535 11961
rect 9587 11909 9599 11961
rect 9651 11909 9657 11961
rect 9399 11883 9657 11909
rect 1798 11021 1850 11027
rect 1798 10957 1850 10969
rect 1798 10893 1850 10905
rect 1798 10829 1850 10841
rect 1798 10765 1850 10777
rect 1798 10707 1850 10713
rect 1914 11021 1966 11027
rect 1914 10957 1966 10969
rect 1914 10893 1966 10905
rect 1914 10829 1966 10841
rect 1914 10765 1966 10777
rect 1914 10707 1966 10713
rect 12029 10236 12157 10242
rect 12029 10184 12035 10236
rect 12087 10184 12099 10236
rect 12151 10184 12157 10236
rect 12029 10163 12157 10184
rect 12029 10111 12035 10163
rect 12087 10111 12099 10163
rect 12151 10111 12157 10163
rect 12029 10090 12157 10111
rect 12029 10038 12035 10090
rect 12087 10038 12099 10090
rect 12151 10038 12157 10090
rect 12029 10017 12157 10038
rect 12029 9965 12035 10017
rect 12087 9965 12099 10017
rect 12151 9965 12157 10017
rect 12029 9944 12157 9965
rect 12029 9892 12035 9944
rect 12087 9892 12099 9944
rect 12151 9892 12157 9944
rect 12029 9870 12157 9892
rect 12029 9818 12035 9870
rect 12087 9818 12099 9870
rect 12151 9818 12157 9870
rect 12029 9812 12157 9818
rect 12029 9626 12157 9632
rect 12029 9574 12035 9626
rect 12087 9574 12099 9626
rect 12151 9574 12157 9626
rect 12029 9561 12157 9574
rect 12029 9509 12035 9561
rect 12087 9509 12099 9561
rect 12151 9509 12157 9561
rect 12029 9496 12157 9509
rect 12029 9444 12035 9496
rect 12087 9444 12099 9496
rect 12151 9444 12157 9496
rect 12029 9431 12157 9444
rect 12029 9379 12035 9431
rect 12087 9379 12099 9431
rect 12151 9379 12157 9431
rect 12029 9365 12157 9379
rect 12029 9313 12035 9365
rect 12087 9313 12099 9365
rect 12151 9313 12157 9365
rect 12029 9299 12157 9313
rect 12029 9247 12035 9299
rect 12087 9247 12099 9299
rect 12151 9247 12157 9299
rect 12029 9233 12157 9247
rect 7677 9068 7807 9198
rect 12029 9181 12035 9233
rect 12087 9181 12099 9233
rect 12151 9181 12157 9233
rect 12029 9175 12157 9181
rect 3361 8767 3413 8773
rect 3361 8703 3413 8715
rect -252 7199 68 7353
rect 3361 5267 3413 8651
rect 12029 8596 12157 8602
rect 12029 8544 12035 8596
rect 12087 8544 12099 8596
rect 12151 8544 12157 8596
rect 12029 8529 12157 8544
rect 12029 8477 12035 8529
rect 12087 8477 12099 8529
rect 12151 8477 12157 8529
rect 12029 8462 12157 8477
rect 12029 8410 12035 8462
rect 12087 8410 12099 8462
rect 12151 8410 12157 8462
rect 12029 8395 12157 8410
rect 12029 8343 12035 8395
rect 12087 8343 12099 8395
rect 12151 8343 12157 8395
rect 12029 8328 12157 8343
rect 12029 8276 12035 8328
rect 12087 8276 12099 8328
rect 12151 8276 12157 8328
rect 12029 8270 12157 8276
rect 5195 7294 5325 7346
rect 12029 7336 12157 7342
rect 12029 7284 12035 7336
rect 12087 7284 12099 7336
rect 12151 7284 12157 7336
rect 12029 7269 12157 7284
rect 12029 7217 12035 7269
rect 12087 7217 12099 7269
rect 12151 7217 12157 7269
rect 12029 7202 12157 7217
rect 12029 7150 12035 7202
rect 12087 7150 12099 7202
rect 12151 7150 12157 7202
rect 12029 7135 12157 7150
rect 12029 7083 12035 7135
rect 12087 7083 12099 7135
rect 12151 7083 12157 7135
rect 12029 7068 12157 7083
rect 12029 7016 12035 7068
rect 12087 7016 12099 7068
rect 12151 7016 12157 7068
rect 12029 7010 12157 7016
rect 5489 6748 5495 6864
rect 5675 6748 5681 6864
rect 6670 6748 6676 6864
rect 6856 6748 6862 6864
rect 7192 6748 7198 6864
rect 7378 6748 7384 6864
rect 12029 6824 12157 6830
rect 12029 6772 12035 6824
rect 12087 6772 12099 6824
rect 12151 6772 12157 6824
rect 12029 6750 12157 6772
rect 12029 6698 12035 6750
rect 12087 6698 12099 6750
rect 12151 6698 12157 6750
rect 12029 6675 12157 6698
rect 12029 6623 12035 6675
rect 12087 6623 12099 6675
rect 12151 6623 12157 6675
rect 12029 6600 12157 6623
rect 12029 6548 12035 6600
rect 12087 6548 12099 6600
rect 12151 6548 12157 6600
rect 12029 6525 12157 6548
rect 12029 6473 12035 6525
rect 12087 6473 12099 6525
rect 12151 6473 12157 6525
rect 12029 6467 12157 6473
rect 3361 5203 3413 5215
rect 3361 5145 3413 5151
rect 8008 6068 8176 6077
rect 8008 6012 8024 6068
rect 8080 6012 8104 6068
rect 8160 6012 8176 6068
rect 8008 5985 8176 6012
rect 8008 5929 8024 5985
rect 8080 5929 8104 5985
rect 8160 5929 8176 5985
rect 8008 5902 8176 5929
rect 8008 5846 8024 5902
rect 8080 5846 8104 5902
rect 8160 5846 8176 5902
rect 8008 5819 8176 5846
rect 8008 5763 8024 5819
rect 8080 5763 8104 5819
rect 8160 5763 8176 5819
rect 8008 5736 8176 5763
rect 8008 5680 8024 5736
rect 8080 5680 8104 5736
rect 8160 5680 8176 5736
rect 8008 5653 8176 5680
rect 8008 5597 8024 5653
rect 8080 5597 8104 5653
rect 8160 5597 8176 5653
rect 8008 5570 8176 5597
rect 8008 5514 8024 5570
rect 8080 5514 8104 5570
rect 8160 5514 8176 5570
rect 8008 5487 8176 5514
rect 8008 5431 8024 5487
rect 8080 5431 8104 5487
rect 8160 5431 8176 5487
rect 8008 5404 8176 5431
rect 8008 5348 8024 5404
rect 8080 5348 8104 5404
rect 8160 5348 8176 5404
rect 8008 5320 8176 5348
rect 8008 5264 8024 5320
rect 8080 5264 8104 5320
rect 8160 5264 8176 5320
rect 8008 5236 8176 5264
rect 8008 5180 8024 5236
rect 8080 5180 8104 5236
rect 8160 5180 8176 5236
rect 8008 5152 8176 5180
rect 8008 5096 8024 5152
rect 8080 5096 8104 5152
rect 8160 5096 8176 5152
rect 8008 5068 8176 5096
rect 8008 5012 8024 5068
rect 8080 5012 8104 5068
rect 8160 5012 8176 5068
rect 8008 4984 8176 5012
rect 8008 4928 8024 4984
rect 8080 4928 8104 4984
rect 8160 4928 8176 4984
rect 8008 4900 8176 4928
rect 8008 4844 8024 4900
rect 8080 4844 8104 4900
rect 8160 4844 8176 4900
rect 8008 4816 8176 4844
rect 8008 4760 8024 4816
rect 8080 4760 8104 4816
rect 8160 4760 8176 4816
rect 8008 4732 8176 4760
rect 8008 4676 8024 4732
rect 8080 4676 8104 4732
rect 8160 4676 8176 4732
rect 8008 4648 8176 4676
rect 8008 4592 8024 4648
rect 8080 4592 8104 4648
rect 8160 4592 8176 4648
rect 8008 4564 8176 4592
rect 8008 4508 8024 4564
rect 8080 4508 8104 4564
rect 8160 4508 8176 4564
rect 8008 4480 8176 4508
rect 8008 4424 8024 4480
rect 8080 4424 8104 4480
rect 8160 4424 8176 4480
rect 8008 4396 8176 4424
rect 8008 4340 8024 4396
rect 8080 4340 8104 4396
rect 8160 4340 8176 4396
rect 8008 4312 8176 4340
rect 8008 4256 8024 4312
rect 8080 4256 8104 4312
rect 8160 4256 8176 4312
rect 8008 4247 8176 4256
rect 10104 6068 10272 6077
rect 10104 6012 10120 6068
rect 10176 6012 10200 6068
rect 10256 6012 10272 6068
rect 10104 5985 10272 6012
rect 10104 5929 10120 5985
rect 10176 5929 10200 5985
rect 10256 5929 10272 5985
rect 10104 5902 10272 5929
rect 10104 5846 10120 5902
rect 10176 5846 10200 5902
rect 10256 5846 10272 5902
rect 10104 5819 10272 5846
rect 10104 5763 10120 5819
rect 10176 5763 10200 5819
rect 10256 5763 10272 5819
rect 10104 5736 10272 5763
rect 10104 5680 10120 5736
rect 10176 5680 10200 5736
rect 10256 5680 10272 5736
rect 10104 5653 10272 5680
rect 10104 5597 10120 5653
rect 10176 5597 10200 5653
rect 10256 5597 10272 5653
rect 10104 5570 10272 5597
rect 10104 5514 10120 5570
rect 10176 5514 10200 5570
rect 10256 5514 10272 5570
rect 10104 5487 10272 5514
rect 10104 5431 10120 5487
rect 10176 5431 10200 5487
rect 10256 5431 10272 5487
rect 10104 5404 10272 5431
rect 10104 5348 10120 5404
rect 10176 5348 10200 5404
rect 10256 5348 10272 5404
rect 10104 5320 10272 5348
rect 10104 5264 10120 5320
rect 10176 5264 10200 5320
rect 10256 5264 10272 5320
rect 10104 5236 10272 5264
rect 10104 5180 10120 5236
rect 10176 5180 10200 5236
rect 10256 5180 10272 5236
rect 10104 5152 10272 5180
rect 10104 5096 10120 5152
rect 10176 5096 10200 5152
rect 10256 5096 10272 5152
rect 10104 5068 10272 5096
rect 10104 5012 10120 5068
rect 10176 5012 10200 5068
rect 10256 5012 10272 5068
rect 10104 4984 10272 5012
rect 10104 4928 10120 4984
rect 10176 4928 10200 4984
rect 10256 4928 10272 4984
rect 10104 4900 10272 4928
rect 10104 4844 10120 4900
rect 10176 4844 10200 4900
rect 10256 4844 10272 4900
rect 10104 4816 10272 4844
rect 10104 4760 10120 4816
rect 10176 4760 10200 4816
rect 10256 4760 10272 4816
rect 10104 4732 10272 4760
rect 10104 4676 10120 4732
rect 10176 4676 10200 4732
rect 10256 4676 10272 4732
rect 10104 4648 10272 4676
rect 10104 4592 10120 4648
rect 10176 4592 10200 4648
rect 10256 4592 10272 4648
rect 10104 4564 10272 4592
rect 10104 4508 10120 4564
rect 10176 4508 10200 4564
rect 10256 4508 10272 4564
rect 10104 4480 10272 4508
rect 10104 4424 10120 4480
rect 10176 4424 10200 4480
rect 10256 4424 10272 4480
rect 10104 4396 10272 4424
rect 10104 4340 10120 4396
rect 10176 4340 10200 4396
rect 10256 4340 10272 4396
rect 10104 4312 10272 4340
rect 10104 4256 10120 4312
rect 10176 4256 10200 4312
rect 10256 4256 10272 4312
rect 10104 4247 10272 4256
rect 11472 6049 11856 6058
rect 11472 5993 11476 6049
rect 11532 5993 11556 6049
rect 11612 5993 11636 6049
rect 11692 5993 11716 6049
rect 11772 5993 11796 6049
rect 11852 5993 11856 6049
rect 11472 5967 11856 5993
rect 11472 5911 11476 5967
rect 11532 5911 11556 5967
rect 11612 5911 11636 5967
rect 11692 5911 11716 5967
rect 11772 5911 11796 5967
rect 11852 5911 11856 5967
rect 11472 5885 11856 5911
rect 11472 5829 11476 5885
rect 11532 5829 11556 5885
rect 11612 5829 11636 5885
rect 11692 5829 11716 5885
rect 11772 5829 11796 5885
rect 11852 5829 11856 5885
rect 11472 5803 11856 5829
rect 11472 5747 11476 5803
rect 11532 5747 11556 5803
rect 11612 5747 11636 5803
rect 11692 5747 11716 5803
rect 11772 5747 11796 5803
rect 11852 5747 11856 5803
rect 11472 5721 11856 5747
rect 11472 5665 11476 5721
rect 11532 5665 11556 5721
rect 11612 5665 11636 5721
rect 11692 5665 11716 5721
rect 11772 5665 11796 5721
rect 11852 5665 11856 5721
rect 11472 5639 11856 5665
rect 11472 5583 11476 5639
rect 11532 5583 11556 5639
rect 11612 5583 11636 5639
rect 11692 5583 11716 5639
rect 11772 5583 11796 5639
rect 11852 5583 11856 5639
rect 11472 5557 11856 5583
rect 11472 5501 11476 5557
rect 11532 5501 11556 5557
rect 11612 5501 11636 5557
rect 11692 5501 11716 5557
rect 11772 5501 11796 5557
rect 11852 5501 11856 5557
rect 11472 5475 11856 5501
rect 11472 5419 11476 5475
rect 11532 5419 11556 5475
rect 11612 5419 11636 5475
rect 11692 5419 11716 5475
rect 11772 5419 11796 5475
rect 11852 5419 11856 5475
rect 11472 5392 11856 5419
rect 11472 5336 11476 5392
rect 11532 5336 11556 5392
rect 11612 5336 11636 5392
rect 11692 5336 11716 5392
rect 11772 5336 11796 5392
rect 11852 5336 11856 5392
rect 11472 5309 11856 5336
rect 11472 5253 11476 5309
rect 11532 5253 11556 5309
rect 11612 5253 11636 5309
rect 11692 5253 11716 5309
rect 11772 5253 11796 5309
rect 11852 5253 11856 5309
rect 12029 5578 12157 5584
rect 12029 5526 12035 5578
rect 12087 5526 12099 5578
rect 12151 5526 12157 5578
rect 12029 5505 12157 5526
rect 12029 5453 12035 5505
rect 12087 5453 12099 5505
rect 12151 5453 12157 5505
rect 12029 5432 12157 5453
rect 12029 5380 12035 5432
rect 12087 5380 12099 5432
rect 12151 5380 12157 5432
rect 12029 5358 12157 5380
rect 12029 5306 12035 5358
rect 12087 5306 12099 5358
rect 12151 5306 12157 5358
rect 12029 5300 12157 5306
rect 11472 5226 11856 5253
rect 11472 5170 11476 5226
rect 11532 5170 11556 5226
rect 11612 5170 11636 5226
rect 11692 5170 11716 5226
rect 11772 5170 11796 5226
rect 11852 5170 11856 5226
rect 11472 5143 11856 5170
rect 11472 5087 11476 5143
rect 11532 5087 11556 5143
rect 11612 5087 11636 5143
rect 11692 5087 11716 5143
rect 11772 5087 11796 5143
rect 11852 5087 11856 5143
rect 11472 5060 11856 5087
rect 11472 5004 11476 5060
rect 11532 5004 11556 5060
rect 11612 5004 11636 5060
rect 11692 5004 11716 5060
rect 11772 5004 11796 5060
rect 11852 5004 11856 5060
rect 11472 4977 11856 5004
rect 11472 4921 11476 4977
rect 11532 4921 11556 4977
rect 11612 4921 11636 4977
rect 11692 4921 11716 4977
rect 11772 4921 11796 4977
rect 11852 4921 11856 4977
rect 11472 4894 11856 4921
rect 11472 4838 11476 4894
rect 11532 4838 11556 4894
rect 11612 4838 11636 4894
rect 11692 4838 11716 4894
rect 11772 4838 11796 4894
rect 11852 4838 11856 4894
rect 11472 4811 11856 4838
rect 11472 4755 11476 4811
rect 11532 4755 11556 4811
rect 11612 4755 11636 4811
rect 11692 4755 11716 4811
rect 11772 4755 11796 4811
rect 11852 4755 11856 4811
rect 11472 4728 11856 4755
rect 11472 4672 11476 4728
rect 11532 4672 11556 4728
rect 11612 4672 11636 4728
rect 11692 4672 11716 4728
rect 11772 4672 11796 4728
rect 11852 4672 11856 4728
rect 11472 4645 11856 4672
rect 11472 4589 11476 4645
rect 11532 4589 11556 4645
rect 11612 4589 11636 4645
rect 11692 4589 11716 4645
rect 11772 4589 11796 4645
rect 11852 4589 11856 4645
rect 11472 4562 11856 4589
rect 11472 4506 11476 4562
rect 11532 4506 11556 4562
rect 11612 4506 11636 4562
rect 11692 4506 11716 4562
rect 11772 4506 11796 4562
rect 11852 4506 11856 4562
rect 11472 4479 11856 4506
rect 11472 4423 11476 4479
rect 11532 4423 11556 4479
rect 11612 4423 11636 4479
rect 11692 4423 11716 4479
rect 11772 4423 11796 4479
rect 11852 4423 11856 4479
rect 11472 4396 11856 4423
rect 11472 4340 11476 4396
rect 11532 4340 11556 4396
rect 11612 4340 11636 4396
rect 11692 4340 11716 4396
rect 11772 4340 11796 4396
rect 11852 4340 11856 4396
rect 11472 4313 11856 4340
rect 11472 4257 11476 4313
rect 11532 4257 11556 4313
rect 11612 4257 11636 4313
rect 11692 4257 11716 4313
rect 11772 4257 11796 4313
rect 11852 4257 11856 4313
rect 11472 4248 11856 4257
rect 12029 4699 12157 4705
rect 12029 4391 12035 4699
rect 12151 4391 12157 4699
rect 12029 4378 12157 4391
rect 12029 4326 12035 4378
rect 12087 4326 12099 4378
rect 12151 4326 12157 4378
rect 12029 4313 12157 4326
rect 12029 4261 12035 4313
rect 12087 4261 12099 4313
rect 12151 4261 12157 4313
rect 12029 4255 12157 4261
rect 12029 4066 12157 4072
rect 12029 4014 12035 4066
rect 12087 4014 12099 4066
rect 12151 4014 12157 4066
rect 12029 4000 12157 4014
rect 12029 3948 12035 4000
rect 12087 3948 12099 4000
rect 12151 3948 12157 4000
rect 12029 3934 12157 3948
rect 12029 3882 12035 3934
rect 12087 3882 12099 3934
rect 12151 3882 12157 3934
rect 12029 3868 12157 3882
rect 12029 3816 12035 3868
rect 12087 3816 12099 3868
rect 12151 3816 12157 3868
rect 12029 3802 12157 3816
rect 12029 3750 12035 3802
rect 12087 3750 12099 3802
rect 12151 3750 12157 3802
rect 12029 3736 12157 3750
rect 12029 3684 12035 3736
rect 12087 3684 12099 3736
rect 12151 3684 12157 3736
rect 12029 3678 12157 3684
rect 1798 3384 1850 3390
rect 1798 3320 1850 3332
rect 1798 3256 1850 3268
rect 1798 3192 1850 3204
rect 1798 3128 1850 3140
rect 1798 3070 1850 3076
rect 1914 3384 1966 3390
rect 1914 3320 1966 3332
rect 1914 3256 1966 3268
rect 1914 3192 1966 3204
rect 1914 3128 1966 3140
rect 1914 3070 1966 3076
rect 4793 2462 4923 2463
rect 4793 2410 4799 2462
rect 4851 2410 4865 2462
rect 4917 2410 4923 2462
rect 4793 2398 4923 2410
rect 4793 2346 4799 2398
rect 4851 2346 4865 2398
rect 4917 2346 4923 2398
rect 4793 2345 4923 2346
rect 7996 2462 8189 2463
rect 7996 2410 8002 2462
rect 8054 2410 8067 2462
rect 7996 2398 8067 2410
rect 7996 2346 8002 2398
rect 8054 2346 8067 2398
rect 8183 2346 8189 2462
rect 7996 2345 8189 2346
rect 4054 2104 4060 2156
rect 4112 2104 4124 2156
rect 4176 2104 4188 2156
rect 4240 2104 4246 2156
rect 5489 2104 5495 2156
rect 5547 2104 5559 2156
rect 5611 2104 5623 2156
rect 5675 2104 5681 2156
rect 6670 2104 6676 2156
rect 6728 2104 6740 2156
rect 6792 2104 6804 2156
rect 6856 2104 6862 2156
rect 7192 2104 7198 2156
rect 7250 2104 7262 2156
rect 7314 2104 7326 2156
rect 7378 2104 7384 2156
rect 8317 2104 8323 2156
rect 8375 2104 8391 2156
rect 8443 2104 8458 2156
rect 8510 2104 8525 2156
rect 8577 2104 8583 2156
rect 10096 1828 10282 1834
rect 10096 1776 10099 1828
rect 10151 1776 10163 1828
rect 10215 1776 10227 1828
rect 10279 1776 10282 1828
rect 10096 1763 10282 1776
rect 10096 1711 10099 1763
rect 10151 1711 10163 1763
rect 10215 1711 10227 1763
rect 10279 1711 10282 1763
rect 10096 1697 10282 1711
rect 10096 1645 10099 1697
rect 10151 1645 10163 1697
rect 10215 1645 10227 1697
rect 10279 1645 10282 1697
tri 12281 1661 12356 1736 se
rect 12356 1713 12408 2586
tri 12356 1661 12408 1713 nw
rect 10096 1639 10282 1645
tri 12259 1639 12281 1661 se
rect 12281 1639 12309 1661
tri 12234 1614 12259 1639 se
rect 12259 1614 12309 1639
tri 12309 1614 12356 1661 nw
rect 11935 1452 11941 1504
rect 11993 1452 12020 1504
rect 12072 1452 12099 1504
rect 12151 1452 12157 1504
rect 4056 1067 4242 1073
rect 4056 1015 4059 1067
rect 4111 1015 4123 1067
rect 4175 1015 4187 1067
rect 4239 1015 4242 1067
rect 4056 1001 4242 1015
rect 4056 949 4059 1001
rect 4111 949 4123 1001
rect 4175 949 4187 1001
rect 4239 949 4242 1001
rect 4056 935 4242 949
rect 4056 883 4059 935
rect 4111 883 4123 935
rect 4175 883 4187 935
rect 4239 883 4242 935
rect 4056 877 4242 883
rect 5491 1067 5677 1073
rect 5491 1015 5494 1067
rect 5546 1015 5558 1067
rect 5610 1015 5622 1067
rect 5674 1015 5677 1067
rect 5491 1001 5677 1015
rect 5491 949 5494 1001
rect 5546 949 5558 1001
rect 5610 949 5622 1001
rect 5674 949 5677 1001
rect 5491 935 5677 949
rect 5491 883 5494 935
rect 5546 883 5558 935
rect 5610 883 5622 935
rect 5674 883 5677 935
rect 5491 877 5677 883
rect 6672 1067 6858 1073
rect 6672 1015 6675 1067
rect 6727 1015 6739 1067
rect 6791 1015 6803 1067
rect 6855 1015 6858 1067
rect 6672 1001 6858 1015
rect 6672 949 6675 1001
rect 6727 949 6739 1001
rect 6791 949 6803 1001
rect 6855 949 6858 1001
rect 6672 935 6858 949
rect 6672 883 6675 935
rect 6727 883 6739 935
rect 6791 883 6803 935
rect 6855 883 6858 935
rect 6672 877 6858 883
rect 7194 1067 7380 1073
rect 7194 1015 7197 1067
rect 7249 1015 7261 1067
rect 7313 1015 7325 1067
rect 7377 1015 7380 1067
rect 7194 1001 7380 1015
rect 7194 949 7197 1001
rect 7249 949 7261 1001
rect 7313 949 7325 1001
rect 7377 949 7380 1001
rect 7194 935 7380 949
rect 7194 883 7197 935
rect 7249 883 7261 935
rect 7313 883 7325 935
rect 7377 883 7380 935
rect 8321 1067 8579 1071
rect 8321 1015 8327 1067
rect 8379 1015 8392 1067
rect 8444 1015 8457 1067
rect 8321 1003 8457 1015
rect 8321 951 8327 1003
rect 8379 951 8392 1003
rect 8444 951 8457 1003
rect 8321 939 8457 951
rect 8321 887 8327 939
rect 8379 887 8392 939
rect 8444 887 8457 939
rect 8573 887 8579 1067
rect 8321 883 8579 887
rect 7194 877 7380 883
rect 10096 785 10282 791
rect 10096 733 10099 785
rect 10151 733 10163 785
rect 10215 733 10227 785
rect 10279 733 10282 785
rect 10096 720 10282 733
rect 7996 710 8189 711
rect 7996 658 8002 710
rect 8054 658 8067 710
rect 7996 646 8067 658
rect 4795 587 4801 639
rect 4853 587 4865 639
rect 4917 587 4923 639
rect 7996 594 8002 646
rect 8054 594 8067 646
rect 8183 594 8189 710
rect 10096 668 10099 720
rect 10151 668 10163 720
rect 10215 668 10227 720
rect 10279 668 10282 720
rect 10096 654 10282 668
rect 10096 602 10099 654
rect 10151 602 10163 654
rect 10215 602 10227 654
rect 10279 602 10282 654
rect 10096 596 10282 602
rect 7996 593 8189 594
tri 10733 113 10984 364 se
rect 10984 258 11240 870
rect 11935 482 12157 1452
rect 12234 1232 12286 1614
tri 12286 1591 12309 1614 nw
rect 12234 1166 12286 1180
rect 12234 1108 12286 1114
rect 12494 1232 12546 1238
rect 12494 1166 12546 1180
rect 12494 1108 12546 1114
rect 10984 113 11095 258
tri 11095 113 11240 258 nw
rect 1294 61 1300 113
rect 1352 61 1366 113
rect 1418 61 1432 113
rect 1484 61 1498 113
rect 1550 61 1564 113
rect 1616 61 1630 113
rect 1682 61 1696 113
rect 1748 61 1762 113
rect 1814 61 1827 113
rect 1879 61 1892 113
rect 1944 61 1957 113
rect 2009 61 2022 113
rect 2074 61 2087 113
rect 2139 61 2152 113
rect 2204 61 2217 113
rect 2269 61 2282 113
rect 2334 61 2347 113
rect 2399 61 2405 113
rect 4054 61 4060 113
rect 4112 61 4124 113
rect 4176 61 4188 113
rect 4240 61 4246 113
rect 5489 61 5495 113
rect 5547 61 5559 113
rect 5611 61 5623 113
rect 5675 61 5681 113
rect 6670 61 6676 113
rect 6728 61 6740 113
rect 6792 61 6804 113
rect 6856 61 6862 113
rect 7192 61 7198 113
rect 7250 61 7262 113
rect 7314 61 7326 113
rect 7378 61 7384 113
rect 8317 61 8323 113
rect 8375 61 8391 113
rect 8443 61 8458 113
rect 8510 61 8525 113
rect 8577 61 8583 113
tri 10681 61 10733 113 se
rect 10733 61 10751 113
rect 10803 61 10819 113
rect 10871 61 10886 113
rect 10938 61 10953 113
rect 11005 61 11043 113
tri 11043 61 11095 113 nw
tri 10622 2 10681 61 se
rect 10681 2 10984 61
tri 10984 2 11043 61 nw
tri 10578 -42 10622 2 se
rect 10622 -42 10940 2
tri 10940 -42 10984 2 nw
tri 10380 -991 10578 -793 se
rect 10578 -899 10834 -42
tri 10834 -148 10940 -42 nw
rect 10578 -991 10742 -899
tri 10742 -991 10834 -899 nw
rect 10380 -2161 10636 -991
tri 10636 -1097 10742 -991 nw
<< via2 >>
rect 14801 27498 14820 27554
rect 14820 27498 14857 27554
rect 14901 27498 14957 27554
rect 15001 27498 15057 27554
rect 15101 27498 15157 27554
rect 15201 27498 15256 27554
rect 15256 27498 15257 27554
rect 14801 27355 14820 27411
rect 14820 27355 14857 27411
rect 14901 27355 14957 27411
rect 15001 27355 15057 27411
rect 15101 27355 15157 27411
rect 15201 27355 15256 27411
rect 15256 27355 15257 27411
rect 14801 27212 14820 27268
rect 14820 27212 14857 27268
rect 14901 27212 14957 27268
rect 15001 27212 15057 27268
rect 15101 27212 15157 27268
rect 15201 27212 15256 27268
rect 15256 27212 15257 27268
rect 14801 27069 14820 27125
rect 14820 27069 14857 27125
rect 14901 27069 14957 27125
rect 15001 27069 15057 27125
rect 15101 27069 15157 27125
rect 15201 27069 15256 27125
rect 15256 27069 15257 27125
rect 13029 26921 13076 26955
rect 13076 26921 13085 26955
rect 13117 26921 13145 26955
rect 13145 26921 13162 26955
rect 13162 26921 13173 26955
rect 13205 26921 13214 26955
rect 13214 26921 13231 26955
rect 13231 26921 13261 26955
rect 13293 26921 13300 26955
rect 13300 26921 13349 26955
rect 13381 26921 13421 26955
rect 13421 26921 13437 26955
rect 13469 26921 13491 26955
rect 13491 26921 13509 26955
rect 13509 26921 13525 26955
rect 13557 26921 13561 26955
rect 13561 26921 13579 26955
rect 13579 26921 13613 26955
rect 13645 26921 13649 26955
rect 13649 26921 13701 26955
rect 13029 26909 13085 26921
rect 13117 26909 13173 26921
rect 13205 26909 13261 26921
rect 13293 26909 13349 26921
rect 13381 26909 13437 26921
rect 13469 26909 13525 26921
rect 13557 26909 13613 26921
rect 13645 26909 13701 26921
rect 13029 26899 13076 26909
rect 13076 26899 13085 26909
rect 13117 26899 13145 26909
rect 13145 26899 13162 26909
rect 13162 26899 13173 26909
rect 13205 26899 13214 26909
rect 13214 26899 13231 26909
rect 13231 26899 13261 26909
rect 13293 26899 13300 26909
rect 13300 26899 13349 26909
rect 13029 26857 13076 26875
rect 13076 26857 13085 26875
rect 13117 26857 13145 26875
rect 13145 26857 13162 26875
rect 13162 26857 13173 26875
rect 13205 26857 13214 26875
rect 13214 26857 13231 26875
rect 13231 26857 13261 26875
rect 13293 26857 13300 26875
rect 13300 26857 13349 26875
rect 13381 26899 13421 26909
rect 13421 26899 13437 26909
rect 13469 26899 13491 26909
rect 13491 26899 13509 26909
rect 13509 26899 13525 26909
rect 13557 26899 13561 26909
rect 13561 26899 13579 26909
rect 13579 26899 13613 26909
rect 13645 26899 13649 26909
rect 13649 26899 13701 26909
rect 13381 26857 13421 26875
rect 13421 26857 13437 26875
rect 13469 26857 13491 26875
rect 13491 26857 13509 26875
rect 13509 26857 13525 26875
rect 13557 26857 13561 26875
rect 13561 26857 13579 26875
rect 13579 26857 13613 26875
rect 13645 26857 13649 26875
rect 13649 26857 13701 26875
rect 13029 26845 13085 26857
rect 13117 26845 13173 26857
rect 13205 26845 13261 26857
rect 13293 26845 13349 26857
rect 13381 26845 13437 26857
rect 13469 26845 13525 26857
rect 13557 26845 13613 26857
rect 13645 26845 13701 26857
rect 13029 26819 13076 26845
rect 13076 26819 13085 26845
rect 13117 26819 13145 26845
rect 13145 26819 13162 26845
rect 13162 26819 13173 26845
rect 13205 26819 13214 26845
rect 13214 26819 13231 26845
rect 13231 26819 13261 26845
rect 13293 26819 13300 26845
rect 13300 26819 13349 26845
rect 13029 26793 13076 26795
rect 13076 26793 13085 26795
rect 13117 26793 13145 26795
rect 13145 26793 13162 26795
rect 13162 26793 13173 26795
rect 13205 26793 13214 26795
rect 13214 26793 13231 26795
rect 13231 26793 13261 26795
rect 13293 26793 13300 26795
rect 13300 26793 13349 26795
rect 13381 26819 13421 26845
rect 13421 26819 13437 26845
rect 13469 26819 13491 26845
rect 13491 26819 13509 26845
rect 13509 26819 13525 26845
rect 13557 26819 13561 26845
rect 13561 26819 13579 26845
rect 13579 26819 13613 26845
rect 13645 26819 13649 26845
rect 13649 26819 13701 26845
rect 13381 26793 13421 26795
rect 13421 26793 13437 26795
rect 13469 26793 13491 26795
rect 13491 26793 13509 26795
rect 13509 26793 13525 26795
rect 13557 26793 13561 26795
rect 13561 26793 13579 26795
rect 13579 26793 13613 26795
rect 13645 26793 13649 26795
rect 13649 26793 13701 26795
rect 13029 26781 13085 26793
rect 13117 26781 13173 26793
rect 13205 26781 13261 26793
rect 13293 26781 13349 26793
rect 13381 26781 13437 26793
rect 13469 26781 13525 26793
rect 13557 26781 13613 26793
rect 13645 26781 13701 26793
rect 13029 26739 13076 26781
rect 13076 26739 13085 26781
rect 13117 26739 13145 26781
rect 13145 26739 13162 26781
rect 13162 26739 13173 26781
rect 13205 26739 13214 26781
rect 13214 26739 13231 26781
rect 13231 26739 13261 26781
rect 13293 26739 13300 26781
rect 13300 26739 13349 26781
rect 13381 26739 13421 26781
rect 13421 26739 13437 26781
rect 13469 26739 13491 26781
rect 13491 26739 13509 26781
rect 13509 26739 13525 26781
rect 13557 26739 13561 26781
rect 13561 26739 13579 26781
rect 13579 26739 13613 26781
rect 13645 26739 13649 26781
rect 13649 26739 13701 26781
rect 14801 26979 14857 26981
rect 14901 26979 14957 26981
rect 15001 26979 15057 26981
rect 15101 26979 15157 26981
rect 15201 26979 15257 26981
rect 14801 26927 14820 26979
rect 14820 26927 14857 26979
rect 14901 26927 14936 26979
rect 14936 26927 14948 26979
rect 14948 26927 14957 26979
rect 15001 26927 15012 26979
rect 15012 26927 15057 26979
rect 15101 26927 15128 26979
rect 15128 26927 15140 26979
rect 15140 26927 15157 26979
rect 15201 26927 15204 26979
rect 15204 26927 15256 26979
rect 15256 26927 15257 26979
rect 14801 26925 14857 26927
rect 14901 26925 14957 26927
rect 15001 26925 15057 26927
rect 15101 26925 15157 26927
rect 15201 26925 15257 26927
rect 13029 26659 13085 26715
rect 13117 26659 13173 26715
rect 13205 26659 13261 26715
rect 13293 26659 13349 26715
rect 13381 26659 13437 26715
rect 13469 26659 13525 26715
rect 13557 26659 13613 26715
rect 13645 26659 13701 26715
rect 13029 26579 13085 26635
rect 13117 26579 13173 26635
rect 13205 26579 13261 26635
rect 13293 26579 13349 26635
rect 13381 26579 13437 26635
rect 13469 26579 13525 26635
rect 13557 26579 13613 26635
rect 13645 26579 13701 26635
rect 13029 26499 13085 26555
rect 13117 26499 13173 26555
rect 13205 26499 13261 26555
rect 13293 26499 13349 26555
rect 13381 26499 13437 26555
rect 13469 26499 13525 26555
rect 13557 26499 13613 26555
rect 13645 26499 13701 26555
rect 13029 26419 13085 26475
rect 13117 26419 13173 26475
rect 13205 26419 13261 26475
rect 13293 26419 13349 26475
rect 13381 26419 13437 26475
rect 13469 26419 13525 26475
rect 13557 26419 13613 26475
rect 13645 26419 13701 26475
rect 13029 26339 13085 26395
rect 13117 26339 13173 26395
rect 13205 26339 13261 26395
rect 13293 26339 13349 26395
rect 13381 26339 13437 26395
rect 13469 26339 13525 26395
rect 13557 26339 13613 26395
rect 13645 26339 13701 26395
rect 13029 26259 13085 26315
rect 13117 26259 13173 26315
rect 13205 26259 13261 26315
rect 13293 26259 13349 26315
rect 13381 26259 13437 26315
rect 13469 26259 13525 26315
rect 13557 26259 13613 26315
rect 13645 26259 13701 26315
rect 13029 26201 13074 26235
rect 13074 26201 13085 26235
rect 13117 26201 13144 26235
rect 13144 26201 13162 26235
rect 13162 26201 13173 26235
rect 13205 26201 13214 26235
rect 13214 26201 13232 26235
rect 13232 26201 13261 26235
rect 13293 26201 13302 26235
rect 13302 26201 13349 26235
rect 13381 26201 13424 26235
rect 13424 26201 13437 26235
rect 13469 26201 13494 26235
rect 13494 26201 13512 26235
rect 13512 26201 13525 26235
rect 13557 26201 13564 26235
rect 13564 26201 13582 26235
rect 13582 26201 13613 26235
rect 13645 26201 13652 26235
rect 13652 26201 13701 26235
rect 13029 26186 13085 26201
rect 13117 26186 13173 26201
rect 13205 26186 13261 26201
rect 13293 26186 13349 26201
rect 13381 26186 13437 26201
rect 13469 26186 13525 26201
rect 13557 26186 13613 26201
rect 13645 26186 13701 26201
rect 13029 26179 13074 26186
rect 13074 26179 13085 26186
rect 13117 26179 13144 26186
rect 13144 26179 13162 26186
rect 13162 26179 13173 26186
rect 13205 26179 13214 26186
rect 13214 26179 13232 26186
rect 13232 26179 13261 26186
rect 13293 26179 13302 26186
rect 13302 26179 13349 26186
rect 13029 26134 13074 26155
rect 13074 26134 13085 26155
rect 13117 26134 13144 26155
rect 13144 26134 13162 26155
rect 13162 26134 13173 26155
rect 13205 26134 13214 26155
rect 13214 26134 13232 26155
rect 13232 26134 13261 26155
rect 13293 26134 13302 26155
rect 13302 26134 13349 26155
rect 13381 26179 13424 26186
rect 13424 26179 13437 26186
rect 13469 26179 13494 26186
rect 13494 26179 13512 26186
rect 13512 26179 13525 26186
rect 13557 26179 13564 26186
rect 13564 26179 13582 26186
rect 13582 26179 13613 26186
rect 13645 26179 13652 26186
rect 13652 26179 13701 26186
rect 13381 26134 13424 26155
rect 13424 26134 13437 26155
rect 13469 26134 13494 26155
rect 13494 26134 13512 26155
rect 13512 26134 13525 26155
rect 13557 26134 13564 26155
rect 13564 26134 13582 26155
rect 13582 26134 13613 26155
rect 13645 26134 13652 26155
rect 13652 26134 13701 26155
rect 13029 26119 13085 26134
rect 13117 26119 13173 26134
rect 13205 26119 13261 26134
rect 13293 26119 13349 26134
rect 13381 26119 13437 26134
rect 13469 26119 13525 26134
rect 13557 26119 13613 26134
rect 13645 26119 13701 26134
rect 13029 26099 13074 26119
rect 13074 26099 13085 26119
rect 13117 26099 13144 26119
rect 13144 26099 13162 26119
rect 13162 26099 13173 26119
rect 13205 26099 13214 26119
rect 13214 26099 13232 26119
rect 13232 26099 13261 26119
rect 13293 26099 13302 26119
rect 13302 26099 13349 26119
rect 13029 26067 13074 26075
rect 13074 26067 13085 26075
rect 13117 26067 13144 26075
rect 13144 26067 13162 26075
rect 13162 26067 13173 26075
rect 13205 26067 13214 26075
rect 13214 26067 13232 26075
rect 13232 26067 13261 26075
rect 13293 26067 13302 26075
rect 13302 26067 13349 26075
rect 13381 26099 13424 26119
rect 13424 26099 13437 26119
rect 13469 26099 13494 26119
rect 13494 26099 13512 26119
rect 13512 26099 13525 26119
rect 13557 26099 13564 26119
rect 13564 26099 13582 26119
rect 13582 26099 13613 26119
rect 13645 26099 13652 26119
rect 13652 26099 13701 26119
rect 13381 26067 13424 26075
rect 13424 26067 13437 26075
rect 13469 26067 13494 26075
rect 13494 26067 13512 26075
rect 13512 26067 13525 26075
rect 13557 26067 13564 26075
rect 13564 26067 13582 26075
rect 13582 26067 13613 26075
rect 13645 26067 13652 26075
rect 13652 26067 13701 26075
rect 13029 26052 13085 26067
rect 13117 26052 13173 26067
rect 13205 26052 13261 26067
rect 13293 26052 13349 26067
rect 13381 26052 13437 26067
rect 13469 26052 13525 26067
rect 13557 26052 13613 26067
rect 13645 26052 13701 26067
rect 13029 26019 13074 26052
rect 13074 26019 13085 26052
rect 13117 26019 13144 26052
rect 13144 26019 13162 26052
rect 13162 26019 13173 26052
rect 13205 26019 13214 26052
rect 13214 26019 13232 26052
rect 13232 26019 13261 26052
rect 13293 26019 13302 26052
rect 13302 26019 13349 26052
rect 13381 26019 13424 26052
rect 13424 26019 13437 26052
rect 13469 26019 13494 26052
rect 13494 26019 13512 26052
rect 13512 26019 13525 26052
rect 13557 26019 13564 26052
rect 13564 26019 13582 26052
rect 13582 26019 13613 26052
rect 13645 26019 13652 26052
rect 13652 26019 13701 26052
rect 13029 25985 13085 25995
rect 13117 25985 13173 25995
rect 13205 25985 13261 25995
rect 13293 25985 13349 25995
rect 13381 25985 13437 25995
rect 13469 25985 13525 25995
rect 13557 25985 13613 25995
rect 13645 25985 13701 25995
rect 13029 25939 13074 25985
rect 13074 25939 13085 25985
rect 13117 25939 13144 25985
rect 13144 25939 13162 25985
rect 13162 25939 13173 25985
rect 13205 25939 13214 25985
rect 13214 25939 13232 25985
rect 13232 25939 13261 25985
rect 13293 25939 13302 25985
rect 13302 25939 13349 25985
rect 13381 25939 13424 25985
rect 13424 25939 13437 25985
rect 13469 25939 13494 25985
rect 13494 25939 13512 25985
rect 13512 25939 13525 25985
rect 13557 25939 13564 25985
rect 13564 25939 13582 25985
rect 13582 25939 13613 25985
rect 13645 25939 13652 25985
rect 13652 25939 13701 25985
rect 13029 25866 13074 25915
rect 13074 25866 13085 25915
rect 13117 25866 13144 25915
rect 13144 25866 13162 25915
rect 13162 25866 13173 25915
rect 13205 25866 13214 25915
rect 13214 25866 13232 25915
rect 13232 25866 13261 25915
rect 13293 25866 13302 25915
rect 13302 25866 13349 25915
rect 13381 25866 13424 25915
rect 13424 25866 13437 25915
rect 13469 25866 13494 25915
rect 13494 25866 13512 25915
rect 13512 25866 13525 25915
rect 13557 25866 13564 25915
rect 13564 25866 13582 25915
rect 13582 25866 13613 25915
rect 13645 25866 13652 25915
rect 13652 25866 13701 25915
rect 13029 25859 13085 25866
rect 13117 25859 13173 25866
rect 13205 25859 13261 25866
rect 13293 25859 13349 25866
rect 13381 25859 13437 25866
rect 13469 25859 13525 25866
rect 13557 25859 13613 25866
rect 13645 25859 13701 25866
rect 13029 25799 13074 25835
rect 13074 25799 13085 25835
rect 13117 25799 13144 25835
rect 13144 25799 13162 25835
rect 13162 25799 13173 25835
rect 13205 25799 13214 25835
rect 13214 25799 13232 25835
rect 13232 25799 13261 25835
rect 13293 25799 13302 25835
rect 13302 25799 13349 25835
rect 13381 25799 13424 25835
rect 13424 25799 13437 25835
rect 13469 25799 13494 25835
rect 13494 25799 13512 25835
rect 13512 25799 13525 25835
rect 13557 25799 13564 25835
rect 13564 25799 13582 25835
rect 13582 25799 13613 25835
rect 13645 25799 13652 25835
rect 13652 25799 13701 25835
rect 13029 25784 13085 25799
rect 13117 25784 13173 25799
rect 13205 25784 13261 25799
rect 13293 25784 13349 25799
rect 13381 25784 13437 25799
rect 13469 25784 13525 25799
rect 13557 25784 13613 25799
rect 13645 25784 13701 25799
rect 13029 25779 13074 25784
rect 13074 25779 13085 25784
rect 13117 25779 13144 25784
rect 13144 25779 13162 25784
rect 13162 25779 13173 25784
rect 13205 25779 13214 25784
rect 13214 25779 13232 25784
rect 13232 25779 13261 25784
rect 13293 25779 13302 25784
rect 13302 25779 13349 25784
rect 13029 25732 13074 25754
rect 13074 25732 13085 25754
rect 13117 25732 13144 25754
rect 13144 25732 13162 25754
rect 13162 25732 13173 25754
rect 13205 25732 13214 25754
rect 13214 25732 13232 25754
rect 13232 25732 13261 25754
rect 13293 25732 13302 25754
rect 13302 25732 13349 25754
rect 13381 25779 13424 25784
rect 13424 25779 13437 25784
rect 13469 25779 13494 25784
rect 13494 25779 13512 25784
rect 13512 25779 13525 25784
rect 13557 25779 13564 25784
rect 13564 25779 13582 25784
rect 13582 25779 13613 25784
rect 13645 25779 13652 25784
rect 13652 25779 13701 25784
rect 13381 25732 13424 25754
rect 13424 25732 13437 25754
rect 13469 25732 13494 25754
rect 13494 25732 13512 25754
rect 13512 25732 13525 25754
rect 13557 25732 13564 25754
rect 13564 25732 13582 25754
rect 13582 25732 13613 25754
rect 13645 25732 13652 25754
rect 13652 25732 13701 25754
rect 13029 25717 13085 25732
rect 13117 25717 13173 25732
rect 13205 25717 13261 25732
rect 13293 25717 13349 25732
rect 13381 25717 13437 25732
rect 13469 25717 13525 25732
rect 13557 25717 13613 25732
rect 13645 25717 13701 25732
rect 13029 25698 13074 25717
rect 13074 25698 13085 25717
rect 13117 25698 13144 25717
rect 13144 25698 13162 25717
rect 13162 25698 13173 25717
rect 13205 25698 13214 25717
rect 13214 25698 13232 25717
rect 13232 25698 13261 25717
rect 13293 25698 13302 25717
rect 13302 25698 13349 25717
rect 13381 25698 13424 25717
rect 13424 25698 13437 25717
rect 13469 25698 13494 25717
rect 13494 25698 13512 25717
rect 13512 25698 13525 25717
rect 13557 25698 13564 25717
rect 13564 25698 13582 25717
rect 13582 25698 13613 25717
rect 13645 25698 13652 25717
rect 13652 25698 13701 25717
rect 8024 6012 8080 6068
rect 8104 6012 8160 6068
rect 8024 5929 8080 5985
rect 8104 5929 8160 5985
rect 8024 5846 8080 5902
rect 8104 5846 8160 5902
rect 8024 5763 8080 5819
rect 8104 5763 8160 5819
rect 8024 5680 8080 5736
rect 8104 5680 8160 5736
rect 8024 5597 8080 5653
rect 8104 5597 8160 5653
rect 8024 5514 8080 5570
rect 8104 5514 8160 5570
rect 8024 5431 8080 5487
rect 8104 5431 8160 5487
rect 8024 5348 8080 5404
rect 8104 5348 8160 5404
rect 8024 5264 8080 5320
rect 8104 5264 8160 5320
rect 8024 5180 8080 5236
rect 8104 5180 8160 5236
rect 8024 5096 8080 5152
rect 8104 5096 8160 5152
rect 8024 5012 8080 5068
rect 8104 5012 8160 5068
rect 8024 4928 8080 4984
rect 8104 4928 8160 4984
rect 8024 4844 8080 4900
rect 8104 4844 8160 4900
rect 8024 4760 8080 4816
rect 8104 4760 8160 4816
rect 8024 4676 8080 4732
rect 8104 4676 8160 4732
rect 8024 4592 8080 4648
rect 8104 4592 8160 4648
rect 8024 4508 8080 4564
rect 8104 4508 8160 4564
rect 8024 4424 8080 4480
rect 8104 4424 8160 4480
rect 8024 4340 8080 4396
rect 8104 4340 8160 4396
rect 8024 4256 8080 4312
rect 8104 4256 8160 4312
rect 10120 6012 10176 6068
rect 10200 6012 10256 6068
rect 10120 5929 10176 5985
rect 10200 5929 10256 5985
rect 10120 5846 10176 5902
rect 10200 5846 10256 5902
rect 10120 5763 10176 5819
rect 10200 5763 10256 5819
rect 10120 5680 10176 5736
rect 10200 5680 10256 5736
rect 10120 5597 10176 5653
rect 10200 5597 10256 5653
rect 10120 5514 10176 5570
rect 10200 5514 10256 5570
rect 10120 5431 10176 5487
rect 10200 5431 10256 5487
rect 10120 5348 10176 5404
rect 10200 5348 10256 5404
rect 10120 5264 10176 5320
rect 10200 5264 10256 5320
rect 10120 5180 10176 5236
rect 10200 5180 10256 5236
rect 10120 5096 10176 5152
rect 10200 5096 10256 5152
rect 10120 5012 10176 5068
rect 10200 5012 10256 5068
rect 10120 4928 10176 4984
rect 10200 4928 10256 4984
rect 10120 4844 10176 4900
rect 10200 4844 10256 4900
rect 10120 4760 10176 4816
rect 10200 4760 10256 4816
rect 10120 4676 10176 4732
rect 10200 4676 10256 4732
rect 10120 4592 10176 4648
rect 10200 4592 10256 4648
rect 10120 4508 10176 4564
rect 10200 4508 10256 4564
rect 10120 4424 10176 4480
rect 10200 4424 10256 4480
rect 10120 4340 10176 4396
rect 10200 4340 10256 4396
rect 10120 4256 10176 4312
rect 10200 4256 10256 4312
rect 11476 5993 11532 6049
rect 11556 5993 11612 6049
rect 11636 5993 11692 6049
rect 11716 5993 11772 6049
rect 11796 5993 11852 6049
rect 11476 5911 11532 5967
rect 11556 5911 11612 5967
rect 11636 5911 11692 5967
rect 11716 5911 11772 5967
rect 11796 5911 11852 5967
rect 11476 5829 11532 5885
rect 11556 5829 11612 5885
rect 11636 5829 11692 5885
rect 11716 5829 11772 5885
rect 11796 5829 11852 5885
rect 11476 5747 11532 5803
rect 11556 5747 11612 5803
rect 11636 5747 11692 5803
rect 11716 5747 11772 5803
rect 11796 5747 11852 5803
rect 11476 5665 11532 5721
rect 11556 5665 11612 5721
rect 11636 5665 11692 5721
rect 11716 5665 11772 5721
rect 11796 5665 11852 5721
rect 11476 5583 11532 5639
rect 11556 5583 11612 5639
rect 11636 5583 11692 5639
rect 11716 5583 11772 5639
rect 11796 5583 11852 5639
rect 11476 5501 11532 5557
rect 11556 5501 11612 5557
rect 11636 5501 11692 5557
rect 11716 5501 11772 5557
rect 11796 5501 11852 5557
rect 11476 5419 11532 5475
rect 11556 5419 11612 5475
rect 11636 5419 11692 5475
rect 11716 5419 11772 5475
rect 11796 5419 11852 5475
rect 11476 5336 11532 5392
rect 11556 5336 11612 5392
rect 11636 5336 11692 5392
rect 11716 5336 11772 5392
rect 11796 5336 11852 5392
rect 11476 5253 11532 5309
rect 11556 5253 11612 5309
rect 11636 5253 11692 5309
rect 11716 5253 11772 5309
rect 11796 5253 11852 5309
rect 11476 5170 11532 5226
rect 11556 5170 11612 5226
rect 11636 5170 11692 5226
rect 11716 5170 11772 5226
rect 11796 5170 11852 5226
rect 11476 5087 11532 5143
rect 11556 5087 11612 5143
rect 11636 5087 11692 5143
rect 11716 5087 11772 5143
rect 11796 5087 11852 5143
rect 11476 5004 11532 5060
rect 11556 5004 11612 5060
rect 11636 5004 11692 5060
rect 11716 5004 11772 5060
rect 11796 5004 11852 5060
rect 11476 4921 11532 4977
rect 11556 4921 11612 4977
rect 11636 4921 11692 4977
rect 11716 4921 11772 4977
rect 11796 4921 11852 4977
rect 11476 4838 11532 4894
rect 11556 4838 11612 4894
rect 11636 4838 11692 4894
rect 11716 4838 11772 4894
rect 11796 4838 11852 4894
rect 11476 4755 11532 4811
rect 11556 4755 11612 4811
rect 11636 4755 11692 4811
rect 11716 4755 11772 4811
rect 11796 4755 11852 4811
rect 11476 4672 11532 4728
rect 11556 4672 11612 4728
rect 11636 4672 11692 4728
rect 11716 4672 11772 4728
rect 11796 4672 11852 4728
rect 11476 4589 11532 4645
rect 11556 4589 11612 4645
rect 11636 4589 11692 4645
rect 11716 4589 11772 4645
rect 11796 4589 11852 4645
rect 11476 4506 11532 4562
rect 11556 4506 11612 4562
rect 11636 4506 11692 4562
rect 11716 4506 11772 4562
rect 11796 4506 11852 4562
rect 11476 4423 11532 4479
rect 11556 4423 11612 4479
rect 11636 4423 11692 4479
rect 11716 4423 11772 4479
rect 11796 4423 11852 4479
rect 11476 4340 11532 4396
rect 11556 4340 11612 4396
rect 11636 4340 11692 4396
rect 11716 4340 11772 4396
rect 11796 4340 11852 4396
rect 11476 4257 11532 4313
rect 11556 4257 11612 4313
rect 11636 4257 11692 4313
rect 11716 4257 11772 4313
rect 11796 4257 11852 4313
<< metal3 >>
rect 13017 27554 15263 27571
rect 13017 27498 14801 27554
rect 14857 27498 14901 27554
rect 14957 27498 15001 27554
rect 15057 27498 15101 27554
rect 15157 27498 15201 27554
rect 15257 27498 15263 27554
rect 13017 27411 15263 27498
rect 13017 27355 14801 27411
rect 14857 27355 14901 27411
rect 14957 27355 15001 27411
rect 15057 27355 15101 27411
rect 15157 27355 15201 27411
rect 15257 27355 15263 27411
rect 13017 27268 15263 27355
rect 13017 27212 14801 27268
rect 14857 27212 14901 27268
rect 14957 27212 15001 27268
rect 15057 27212 15101 27268
rect 15157 27212 15201 27268
rect 15257 27212 15263 27268
rect 13017 27125 15263 27212
rect 13017 27069 14801 27125
rect 14857 27069 14901 27125
rect 14957 27069 15001 27125
rect 15057 27069 15101 27125
rect 15157 27069 15201 27125
rect 15257 27069 15263 27125
rect 13017 26981 15263 27069
rect 13017 26955 14801 26981
rect 13017 26899 13029 26955
rect 13085 26899 13117 26955
rect 13173 26899 13205 26955
rect 13261 26899 13293 26955
rect 13349 26899 13381 26955
rect 13437 26899 13469 26955
rect 13525 26899 13557 26955
rect 13613 26899 13645 26955
rect 13701 26925 14801 26955
rect 14857 26925 14901 26981
rect 14957 26925 15001 26981
rect 15057 26925 15101 26981
rect 15157 26925 15201 26981
rect 15257 26925 15263 26981
rect 13701 26899 15263 26925
rect 13017 26875 15263 26899
rect 13017 26819 13029 26875
rect 13085 26819 13117 26875
rect 13173 26819 13205 26875
rect 13261 26819 13293 26875
rect 13349 26819 13381 26875
rect 13437 26819 13469 26875
rect 13525 26819 13557 26875
rect 13613 26819 13645 26875
rect 13701 26819 15263 26875
rect 13017 26795 15263 26819
rect 13017 26739 13029 26795
rect 13085 26739 13117 26795
rect 13173 26739 13205 26795
rect 13261 26739 13293 26795
rect 13349 26739 13381 26795
rect 13437 26739 13469 26795
rect 13525 26739 13557 26795
rect 13613 26739 13645 26795
rect 13701 26739 15263 26795
rect 13017 26715 15263 26739
rect 13017 26659 13029 26715
rect 13085 26659 13117 26715
rect 13173 26659 13205 26715
rect 13261 26659 13293 26715
rect 13349 26659 13381 26715
rect 13437 26659 13469 26715
rect 13525 26659 13557 26715
rect 13613 26659 13645 26715
rect 13701 26659 15263 26715
rect 13017 26635 15263 26659
rect 13017 26579 13029 26635
rect 13085 26579 13117 26635
rect 13173 26579 13205 26635
rect 13261 26579 13293 26635
rect 13349 26579 13381 26635
rect 13437 26579 13469 26635
rect 13525 26579 13557 26635
rect 13613 26579 13645 26635
rect 13701 26592 15263 26635
rect 13701 26579 13715 26592
rect 13017 26555 13715 26579
rect 13017 26499 13029 26555
rect 13085 26499 13117 26555
rect 13173 26499 13205 26555
rect 13261 26499 13293 26555
rect 13349 26499 13381 26555
rect 13437 26499 13469 26555
rect 13525 26499 13557 26555
rect 13613 26499 13645 26555
rect 13701 26499 13715 26555
rect 13017 26475 13715 26499
rect 13017 26419 13029 26475
rect 13085 26419 13117 26475
rect 13173 26419 13205 26475
rect 13261 26419 13293 26475
rect 13349 26419 13381 26475
rect 13437 26419 13469 26475
rect 13525 26419 13557 26475
rect 13613 26419 13645 26475
rect 13701 26419 13715 26475
rect 13017 26395 13715 26419
rect 13017 26339 13029 26395
rect 13085 26339 13117 26395
rect 13173 26339 13205 26395
rect 13261 26339 13293 26395
rect 13349 26339 13381 26395
rect 13437 26339 13469 26395
rect 13525 26339 13557 26395
rect 13613 26339 13645 26395
rect 13701 26339 13715 26395
rect 13017 26315 13715 26339
rect 13017 26259 13029 26315
rect 13085 26259 13117 26315
rect 13173 26259 13205 26315
rect 13261 26259 13293 26315
rect 13349 26259 13381 26315
rect 13437 26259 13469 26315
rect 13525 26259 13557 26315
rect 13613 26259 13645 26315
rect 13701 26259 13715 26315
rect 13017 26235 13715 26259
rect 13017 26179 13029 26235
rect 13085 26179 13117 26235
rect 13173 26179 13205 26235
rect 13261 26179 13293 26235
rect 13349 26179 13381 26235
rect 13437 26179 13469 26235
rect 13525 26179 13557 26235
rect 13613 26179 13645 26235
rect 13701 26179 13715 26235
rect 13017 26155 13715 26179
rect 13017 26099 13029 26155
rect 13085 26099 13117 26155
rect 13173 26099 13205 26155
rect 13261 26099 13293 26155
rect 13349 26099 13381 26155
rect 13437 26099 13469 26155
rect 13525 26099 13557 26155
rect 13613 26099 13645 26155
rect 13701 26099 13715 26155
rect 13017 26075 13715 26099
rect 13017 26019 13029 26075
rect 13085 26019 13117 26075
rect 13173 26019 13205 26075
rect 13261 26019 13293 26075
rect 13349 26019 13381 26075
rect 13437 26019 13469 26075
rect 13525 26019 13557 26075
rect 13613 26019 13645 26075
rect 13701 26019 13715 26075
rect 13017 25995 13715 26019
rect 13017 25939 13029 25995
rect 13085 25939 13117 25995
rect 13173 25939 13205 25995
rect 13261 25939 13293 25995
rect 13349 25939 13381 25995
rect 13437 25939 13469 25995
rect 13525 25939 13557 25995
rect 13613 25939 13645 25995
rect 13701 25939 13715 25995
rect 13017 25915 13715 25939
rect 13017 25859 13029 25915
rect 13085 25859 13117 25915
rect 13173 25859 13205 25915
rect 13261 25859 13293 25915
rect 13349 25859 13381 25915
rect 13437 25859 13469 25915
rect 13525 25859 13557 25915
rect 13613 25859 13645 25915
rect 13701 25859 13715 25915
rect 13017 25835 13715 25859
rect 13017 25779 13029 25835
rect 13085 25779 13117 25835
rect 13173 25779 13205 25835
rect 13261 25779 13293 25835
rect 13349 25779 13381 25835
rect 13437 25779 13469 25835
rect 13525 25779 13557 25835
rect 13613 25779 13645 25835
rect 13701 25779 13715 25835
rect 13017 25754 13715 25779
rect 13017 25698 13029 25754
rect 13085 25698 13117 25754
rect 13173 25698 13205 25754
rect 13261 25698 13293 25754
rect 13349 25698 13381 25754
rect 13437 25698 13469 25754
rect 13525 25698 13557 25754
rect 13613 25698 13645 25754
rect 13701 25698 13715 25754
rect 13017 25684 13715 25698
tri 13715 25684 14623 26592 nw
rect 8003 6068 8181 6073
rect 8003 6012 8024 6068
rect 8080 6012 8104 6068
rect 8160 6012 8181 6068
rect 8003 5985 8181 6012
rect 8003 5929 8024 5985
rect 8080 5929 8104 5985
rect 8160 5929 8181 5985
rect 8003 5902 8181 5929
rect 8003 5846 8024 5902
rect 8080 5846 8104 5902
rect 8160 5846 8181 5902
rect 8003 5819 8181 5846
rect 8003 5763 8024 5819
rect 8080 5763 8104 5819
rect 8160 5763 8181 5819
rect 8003 5736 8181 5763
rect 8003 5680 8024 5736
rect 8080 5680 8104 5736
rect 8160 5680 8181 5736
rect 8003 5653 8181 5680
rect 8003 5597 8024 5653
rect 8080 5597 8104 5653
rect 8160 5597 8181 5653
rect 8003 5570 8181 5597
rect 8003 5514 8024 5570
rect 8080 5514 8104 5570
rect 8160 5514 8181 5570
rect 8003 5487 8181 5514
rect 8003 5431 8024 5487
rect 8080 5431 8104 5487
rect 8160 5431 8181 5487
rect 8003 5404 8181 5431
rect 8003 5348 8024 5404
rect 8080 5348 8104 5404
rect 8160 5348 8181 5404
rect 8003 5320 8181 5348
rect 8003 5264 8024 5320
rect 8080 5264 8104 5320
rect 8160 5264 8181 5320
rect 8003 5236 8181 5264
rect 8003 5180 8024 5236
rect 8080 5180 8104 5236
rect 8160 5180 8181 5236
rect 8003 5152 8181 5180
rect 8003 5096 8024 5152
rect 8080 5096 8104 5152
rect 8160 5096 8181 5152
rect 8003 5068 8181 5096
rect 8003 5012 8024 5068
rect 8080 5012 8104 5068
rect 8160 5012 8181 5068
rect 8003 4984 8181 5012
rect 8003 4928 8024 4984
rect 8080 4928 8104 4984
rect 8160 4928 8181 4984
rect 8003 4900 8181 4928
rect 8003 4844 8024 4900
rect 8080 4844 8104 4900
rect 8160 4844 8181 4900
rect 8003 4816 8181 4844
rect 8003 4760 8024 4816
rect 8080 4760 8104 4816
rect 8160 4760 8181 4816
rect 8003 4732 8181 4760
rect 8003 4676 8024 4732
rect 8080 4676 8104 4732
rect 8160 4676 8181 4732
rect 8003 4648 8181 4676
rect 8003 4592 8024 4648
rect 8080 4592 8104 4648
rect 8160 4592 8181 4648
rect 8003 4564 8181 4592
rect 8003 4508 8024 4564
rect 8080 4508 8104 4564
rect 8160 4508 8181 4564
rect 8003 4480 8181 4508
rect 8003 4424 8024 4480
rect 8080 4424 8104 4480
rect 8160 4424 8181 4480
rect 8003 4396 8181 4424
rect 8003 4340 8024 4396
rect 8080 4340 8104 4396
rect 8160 4340 8181 4396
rect 8003 4312 8181 4340
rect 8003 4256 8024 4312
rect 8080 4256 8104 4312
rect 8160 4256 8181 4312
rect 8003 4251 8181 4256
rect 10099 6068 10277 6073
rect 10099 6012 10120 6068
rect 10176 6012 10200 6068
rect 10256 6012 10277 6068
rect 10099 5985 10277 6012
rect 10099 5929 10120 5985
rect 10176 5929 10200 5985
rect 10256 5929 10277 5985
rect 10099 5902 10277 5929
rect 10099 5846 10120 5902
rect 10176 5846 10200 5902
rect 10256 5846 10277 5902
rect 10099 5819 10277 5846
rect 10099 5763 10120 5819
rect 10176 5763 10200 5819
rect 10256 5763 10277 5819
rect 10099 5736 10277 5763
rect 10099 5680 10120 5736
rect 10176 5680 10200 5736
rect 10256 5680 10277 5736
rect 10099 5653 10277 5680
rect 10099 5597 10120 5653
rect 10176 5597 10200 5653
rect 10256 5597 10277 5653
rect 10099 5570 10277 5597
rect 10099 5514 10120 5570
rect 10176 5514 10200 5570
rect 10256 5514 10277 5570
rect 10099 5487 10277 5514
rect 10099 5431 10120 5487
rect 10176 5431 10200 5487
rect 10256 5431 10277 5487
rect 10099 5404 10277 5431
rect 10099 5348 10120 5404
rect 10176 5348 10200 5404
rect 10256 5348 10277 5404
rect 10099 5320 10277 5348
rect 10099 5264 10120 5320
rect 10176 5264 10200 5320
rect 10256 5264 10277 5320
rect 10099 5236 10277 5264
rect 10099 5180 10120 5236
rect 10176 5180 10200 5236
rect 10256 5180 10277 5236
rect 10099 5152 10277 5180
rect 10099 5096 10120 5152
rect 10176 5096 10200 5152
rect 10256 5096 10277 5152
rect 10099 5068 10277 5096
rect 10099 5012 10120 5068
rect 10176 5012 10200 5068
rect 10256 5012 10277 5068
rect 10099 4984 10277 5012
rect 10099 4928 10120 4984
rect 10176 4928 10200 4984
rect 10256 4928 10277 4984
rect 10099 4900 10277 4928
rect 10099 4844 10120 4900
rect 10176 4844 10200 4900
rect 10256 4844 10277 4900
rect 10099 4816 10277 4844
rect 10099 4760 10120 4816
rect 10176 4760 10200 4816
rect 10256 4760 10277 4816
rect 10099 4732 10277 4760
rect 10099 4676 10120 4732
rect 10176 4676 10200 4732
rect 10256 4676 10277 4732
rect 10099 4648 10277 4676
rect 10099 4592 10120 4648
rect 10176 4592 10200 4648
rect 10256 4592 10277 4648
rect 10099 4564 10277 4592
rect 10099 4508 10120 4564
rect 10176 4508 10200 4564
rect 10256 4508 10277 4564
rect 10099 4480 10277 4508
rect 10099 4424 10120 4480
rect 10176 4424 10200 4480
rect 10256 4424 10277 4480
rect 10099 4396 10277 4424
rect 10099 4340 10120 4396
rect 10176 4340 10200 4396
rect 10256 4340 10277 4396
rect 10099 4312 10277 4340
rect 10099 4256 10120 4312
rect 10176 4256 10200 4312
rect 10256 4256 10277 4312
rect 10099 4251 10277 4256
rect 11467 6049 11861 6054
rect 11467 5993 11476 6049
rect 11532 5993 11556 6049
rect 11612 5993 11636 6049
rect 11692 5993 11716 6049
rect 11772 5993 11796 6049
rect 11852 5993 11861 6049
rect 11467 5967 11861 5993
rect 11467 5911 11476 5967
rect 11532 5911 11556 5967
rect 11612 5911 11636 5967
rect 11692 5911 11716 5967
rect 11772 5911 11796 5967
rect 11852 5911 11861 5967
rect 11467 5885 11861 5911
rect 11467 5829 11476 5885
rect 11532 5829 11556 5885
rect 11612 5829 11636 5885
rect 11692 5829 11716 5885
rect 11772 5829 11796 5885
rect 11852 5829 11861 5885
rect 11467 5803 11861 5829
rect 11467 5747 11476 5803
rect 11532 5747 11556 5803
rect 11612 5747 11636 5803
rect 11692 5747 11716 5803
rect 11772 5747 11796 5803
rect 11852 5747 11861 5803
rect 11467 5721 11861 5747
rect 11467 5665 11476 5721
rect 11532 5665 11556 5721
rect 11612 5665 11636 5721
rect 11692 5665 11716 5721
rect 11772 5665 11796 5721
rect 11852 5665 11861 5721
rect 11467 5639 11861 5665
rect 11467 5583 11476 5639
rect 11532 5583 11556 5639
rect 11612 5583 11636 5639
rect 11692 5583 11716 5639
rect 11772 5583 11796 5639
rect 11852 5583 11861 5639
rect 11467 5557 11861 5583
rect 11467 5501 11476 5557
rect 11532 5501 11556 5557
rect 11612 5501 11636 5557
rect 11692 5501 11716 5557
rect 11772 5501 11796 5557
rect 11852 5501 11861 5557
rect 11467 5475 11861 5501
rect 11467 5419 11476 5475
rect 11532 5419 11556 5475
rect 11612 5419 11636 5475
rect 11692 5419 11716 5475
rect 11772 5419 11796 5475
rect 11852 5419 11861 5475
rect 11467 5392 11861 5419
rect 11467 5336 11476 5392
rect 11532 5336 11556 5392
rect 11612 5336 11636 5392
rect 11692 5336 11716 5392
rect 11772 5336 11796 5392
rect 11852 5336 11861 5392
rect 11467 5309 11861 5336
rect 11467 5253 11476 5309
rect 11532 5253 11556 5309
rect 11612 5253 11636 5309
rect 11692 5253 11716 5309
rect 11772 5253 11796 5309
rect 11852 5253 11861 5309
rect 11467 5226 11861 5253
rect 11467 5170 11476 5226
rect 11532 5170 11556 5226
rect 11612 5170 11636 5226
rect 11692 5170 11716 5226
rect 11772 5170 11796 5226
rect 11852 5170 11861 5226
rect 11467 5143 11861 5170
rect 11467 5087 11476 5143
rect 11532 5087 11556 5143
rect 11612 5087 11636 5143
rect 11692 5087 11716 5143
rect 11772 5087 11796 5143
rect 11852 5087 11861 5143
rect 11467 5060 11861 5087
rect 11467 5004 11476 5060
rect 11532 5004 11556 5060
rect 11612 5004 11636 5060
rect 11692 5004 11716 5060
rect 11772 5004 11796 5060
rect 11852 5004 11861 5060
rect 11467 4977 11861 5004
rect 11467 4921 11476 4977
rect 11532 4921 11556 4977
rect 11612 4921 11636 4977
rect 11692 4921 11716 4977
rect 11772 4921 11796 4977
rect 11852 4921 11861 4977
rect 11467 4894 11861 4921
rect 11467 4838 11476 4894
rect 11532 4838 11556 4894
rect 11612 4838 11636 4894
rect 11692 4838 11716 4894
rect 11772 4838 11796 4894
rect 11852 4838 11861 4894
rect 11467 4811 11861 4838
rect 11467 4755 11476 4811
rect 11532 4755 11556 4811
rect 11612 4755 11636 4811
rect 11692 4755 11716 4811
rect 11772 4755 11796 4811
rect 11852 4755 11861 4811
rect 11467 4728 11861 4755
rect 11467 4672 11476 4728
rect 11532 4672 11556 4728
rect 11612 4672 11636 4728
rect 11692 4672 11716 4728
rect 11772 4672 11796 4728
rect 11852 4672 11861 4728
rect 11467 4645 11861 4672
rect 11467 4589 11476 4645
rect 11532 4589 11556 4645
rect 11612 4589 11636 4645
rect 11692 4589 11716 4645
rect 11772 4589 11796 4645
rect 11852 4589 11861 4645
rect 11467 4562 11861 4589
rect 11467 4506 11476 4562
rect 11532 4506 11556 4562
rect 11612 4506 11636 4562
rect 11692 4506 11716 4562
rect 11772 4506 11796 4562
rect 11852 4506 11861 4562
rect 11467 4479 11861 4506
rect 11467 4423 11476 4479
rect 11532 4423 11556 4479
rect 11612 4423 11636 4479
rect 11692 4423 11716 4479
rect 11772 4423 11796 4479
rect 11852 4423 11861 4479
rect 11467 4396 11861 4423
rect 11467 4340 11476 4396
rect 11532 4340 11556 4396
rect 11612 4340 11636 4396
rect 11692 4340 11716 4396
rect 11772 4340 11796 4396
rect 11852 4340 11861 4396
rect 11467 4313 11861 4340
rect 11467 4257 11476 4313
rect 11532 4257 11556 4313
rect 11612 4257 11636 4313
rect 11692 4257 11716 4313
rect 11772 4257 11796 4313
rect 11852 4257 11861 4313
rect 11467 4252 11861 4257
<< metal4 >>
rect -3589 18005 -3164 18876
<< comment >>
tri 13921 17918 13932 17919 se
rect 13932 17918 13952 17919
tri 13952 17918 13963 17919 sw
tri 13911 17917 13921 17918 se
rect 13921 17917 13963 17918
tri 13963 17917 13973 17918 sw
tri 13901 17916 13911 17917 se
rect 13911 17916 13973 17917
tri 13973 17916 13983 17917 sw
tri 13892 17915 13901 17916 se
rect 13901 17915 13983 17916
tri 13983 17915 13992 17916 sw
tri 13883 17913 13892 17915 se
rect 13892 17913 13992 17915
tri 13992 17913 14001 17915 sw
tri 13875 17911 13883 17913 se
rect 13883 17911 14001 17913
tri 14001 17911 14009 17913 sw
tri 13867 17908 13875 17911 se
rect 13875 17908 14009 17911
tri 14009 17908 14017 17911 sw
tri 13860 17906 13867 17908 se
rect 13867 17906 14017 17908
tri 14017 17906 14024 17908 sw
tri 13854 17903 13860 17906 se
rect 13860 17903 14024 17906
tri 14024 17903 14030 17906 sw
tri 13849 17900 13854 17903 se
rect 13854 17900 14030 17903
tri 14030 17900 14035 17903 sw
tri 13844 17897 13849 17900 se
rect 13849 17897 14035 17900
tri 14035 17897 14040 17900 sw
tri 13841 17893 13844 17897 se
rect 13844 17893 14040 17897
tri 14040 17893 14043 17897 sw
tri 13838 17890 13841 17893 se
rect 13841 17890 14043 17893
tri 14043 17890 14046 17893 sw
tri 13837 17887 13838 17890 se
rect 13838 17887 14046 17890
tri 14046 17887 14047 17890 sw
tri 13836 17883 13837 17887 se
tri 13836 17879 13837 17883 ne
rect 13837 17879 14047 17887
tri 14047 17883 14048 17887 sw
tri 14047 17879 14048 17883 nw
tri 13837 17876 13838 17879 ne
rect 13838 17876 14046 17879
tri 14046 17876 14047 17879 nw
tri 13838 17873 13841 17876 ne
rect 13841 17873 14043 17876
tri 14043 17873 14046 17876 nw
tri 13841 17869 13844 17873 ne
rect 13844 17869 14040 17873
tri 14040 17869 14043 17873 nw
tri 13844 17866 13849 17869 ne
rect 13849 17866 14035 17869
tri 14035 17866 14040 17869 nw
tri 13849 17863 13854 17866 ne
rect 13854 17863 14030 17866
tri 14030 17863 14035 17866 nw
tri 13854 17860 13860 17863 ne
rect 13860 17860 14024 17863
tri 14024 17860 14030 17863 nw
tri 13860 17858 13867 17860 ne
rect 13867 17858 14017 17860
tri 14017 17858 14024 17860 nw
tri 13867 17856 13872 17858 ne
rect 13872 17856 14009 17858
tri 13733 17855 13743 17856 se
rect 13743 17855 13765 17856
tri 13765 17855 13773 17856 sw
tri 13873 17855 13875 17856 ne
rect 13875 17855 14009 17856
tri 14009 17855 14017 17858 nw
tri 13722 17854 13733 17855 se
rect 13733 17854 13775 17855
tri 13775 17854 13786 17855 sw
tri 13875 17854 13879 17855 ne
rect 13879 17854 14001 17855
tri 13712 17852 13722 17854 se
rect 13722 17853 13786 17854
tri 13786 17853 13792 17854 sw
tri 13879 17853 13883 17854 ne
rect 13883 17853 14001 17854
tri 14001 17853 14009 17855 nw
rect 13722 17852 13792 17853
tri 13792 17852 13796 17853 sw
tri 13883 17852 13886 17853 ne
rect 13886 17852 13992 17853
tri 13702 17850 13712 17852 se
rect 13712 17851 13796 17852
tri 13796 17851 13802 17852 sw
tri 13886 17851 13892 17852 ne
rect 13892 17851 13992 17852
tri 13992 17851 14001 17853 nw
rect 13712 17850 13802 17851
tri 13802 17850 13806 17851 sw
tri 13892 17850 13897 17851 ne
rect 13897 17850 13983 17851
tri 13983 17850 13992 17851 nw
tri 13693 17848 13702 17850 se
rect 13702 17849 13808 17850
tri 13808 17849 13813 17850 sw
tri 13901 17849 13911 17850 ne
rect 13911 17849 13973 17850
tri 13973 17849 13983 17850 nw
rect 13702 17848 13813 17849
tri 13813 17848 13815 17849 sw
tri 13911 17848 13917 17849 ne
rect 13917 17848 13963 17849
tri 13963 17848 13973 17849 nw
tri 13684 17845 13693 17848 se
rect 13693 17847 13816 17848
tri 13816 17847 13818 17848 sw
tri 13921 17847 13932 17848 ne
rect 13932 17847 13952 17848
tri 13952 17847 13963 17848 nw
rect 13693 17845 13818 17847
tri 13818 17845 13824 17847 sw
tri 13676 17842 13684 17845 se
rect 13684 17842 13824 17845
tri 13824 17842 13832 17845 sw
tri 13669 17838 13676 17842 se
rect 13676 17838 13832 17842
tri 13832 17838 13839 17842 sw
tri 13663 17835 13669 17838 se
rect 13669 17835 13839 17838
tri 13839 17835 13845 17838 sw
tri 13657 17831 13663 17835 se
rect 13663 17831 13845 17835
tri 13845 17831 13851 17835 sw
tri 13652 17826 13657 17831 se
rect 13657 17826 13851 17831
tri 13851 17826 13856 17831 sw
tri 13649 17822 13652 17826 se
rect 13652 17822 13856 17826
tri 13856 17822 13859 17826 sw
tri 13646 17817 13649 17822 se
rect 13649 17817 13859 17822
tri 13859 17817 13862 17822 sw
tri 13645 17813 13646 17817 se
rect 13646 17813 13862 17817
tri 13862 17813 13863 17817 sw
tri 13644 17808 13645 17813 se
tri 13644 17803 13645 17808 ne
rect 13645 17803 13863 17813
tri 13863 17808 13864 17813 sw
tri 13863 17803 13864 17808 nw
tri 13645 17799 13646 17803 ne
rect 13646 17799 13862 17803
tri 13862 17799 13863 17803 nw
tri 13646 17794 13649 17799 ne
rect 13649 17794 13859 17799
tri 13859 17794 13862 17799 nw
tri 13649 17790 13652 17794 ne
rect 13652 17790 13856 17794
tri 13856 17790 13859 17794 nw
tri 13652 17785 13657 17790 ne
rect 13657 17785 13851 17790
tri 13851 17785 13856 17790 nw
tri 13657 17781 13663 17785 ne
rect 13663 17781 13845 17785
tri 13845 17781 13851 17785 nw
tri 13663 17778 13669 17781 ne
rect 13669 17778 13839 17781
tri 13839 17778 13845 17781 nw
tri 13669 17774 13676 17778 ne
rect 13676 17774 13832 17778
tri 13832 17774 13839 17778 nw
tri 13676 17771 13684 17774 ne
rect 13684 17771 13824 17774
tri 13824 17771 13832 17774 nw
tri 13684 17768 13693 17771 ne
rect 13693 17768 13815 17771
tri 13815 17768 13824 17771 nw
tri 13693 17766 13702 17768 ne
rect 13702 17766 13806 17768
tri 13806 17766 13815 17768 nw
tri 13702 17764 13712 17766 ne
rect 13712 17764 13796 17766
tri 13796 17764 13806 17766 nw
tri 13712 17762 13722 17764 ne
rect 13722 17762 13786 17764
tri 13786 17762 13796 17764 nw
tri 13722 17761 13733 17762 ne
rect 13733 17761 13775 17762
tri 13775 17761 13786 17762 nw
tri 13733 17760 13743 17761 ne
rect 13743 17760 13765 17761
tri 13765 17760 13775 17761 nw
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 985 -1 0 3305
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 10945 1 0 17253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1701704242
transform 0 -1 1841 -1 0 11015
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1701704242
transform 0 -1 1957 -1 0 11015
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_2
timestamp 1701704242
transform 0 -1 1957 1 0 3082
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_3
timestamp 1701704242
transform 0 -1 1841 1 0 3082
box 0 0 1 1
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1701704242
transform 0 -1 1957 -1 0 10217
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1701704242
transform 0 -1 1957 1 0 3699
box -12 -6 910 40
use L1M1_CDNS_524688791851017  L1M1_CDNS_524688791851017_0
timestamp 1701704242
transform 0 -1 517 -1 0 10738
box -12 -6 1918 40
use L1M1_CDNS_524688791851017  L1M1_CDNS_524688791851017_1
timestamp 1701704242
transform 0 -1 517 1 0 3178
box -12 -6 1918 40
use L1M1_CDNS_524688791851558  L1M1_CDNS_524688791851558_0
timestamp 1701704242
transform 1 0 9928 0 1 26720
box -12 -6 262 3784
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform -1 0 7686 0 -1 29557
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform -1 0 7686 0 -1 29468
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform -1 0 8126 0 -1 29557
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform -1 0 8126 0 -1 29468
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 1 2098 1 0 29288
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 -1 9060 1 0 29611
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 -1 8980 1 0 29611
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 -1 3413 1 0 5145
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 -1 3413 1 0 8645
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 1 0 5800 0 -1 24989
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 1 0 8491 0 -1 24909
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 1 0 8491 0 -1 25074
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 1 0 5947 0 -1 24909
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 1 0 8427 0 -1 25010
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 1 0 14035 0 1 17859
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform 1 0 6652 0 1 17859
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform 1 0 13335 0 1 17784
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1701704242
transform 1 0 5901 0 1 17784
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1701704242
transform 1 0 4878 0 1 19976
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1701704242
transform 1 0 4878 0 1 19868
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1701704242
transform 1 0 729 0 1 19868
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1701704242
transform 1 0 729 0 1 19976
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1701704242
transform 1 0 4795 0 1 587
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1701704242
transform 0 1 9582 1 0 29478
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1701704242
transform 1 0 10984 0 1 870
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_2
timestamp 1701704242
transform 1 0 6814 0 1 25017
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_3
timestamp 1701704242
transform 1 0 6814 0 1 17939
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_4
timestamp 1701704242
transform 1 0 8317 0 1 6748
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_5
timestamp 1701704242
transform 1 0 9399 0 1 6748
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_6
timestamp 1701704242
transform 1 0 8659 0 1 18091
box 0 0 256 116
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1701704242
transform 1 0 3003 0 1 20732
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1701704242
transform 1 0 3003 0 1 18024
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1701704242
transform 1 0 5489 0 1 6748
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_3
timestamp 1701704242
transform 1 0 6670 0 1 6748
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_4
timestamp 1701704242
transform 1 0 7192 0 1 6748
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform -1 0 7704 0 -1 22110
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1701704242
transform 0 -1 5506 1 0 21982
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1701704242
transform 0 -1 5089 1 0 21794
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1701704242
transform 1 0 4518 0 1 20732
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1701704242
transform 0 1 7760 1 0 21797
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1701704242
transform 1 0 9904 0 1 29946
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1701704242
transform 1 0 12442 0 1 17947
box 0 0 320 116
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1701704242
transform 0 -1 1850 -1 0 11027
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1701704242
transform 0 -1 1966 -1 0 11027
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1701704242
transform 0 -1 1966 1 0 3070
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_3
timestamp 1701704242
transform 0 -1 1850 1 0 3070
box 0 0 1 1
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1701704242
transform 0 -1 8391 1 0 29767
box 0 0 128 244
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 0 1 4679 1 0 29799
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform 0 1 5243 1 0 29799
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1701704242
transform 0 1 5097 1 0 29799
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_0
timestamp 1701704242
transform 1 0 6652 0 1 18308
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1701704242
transform -1 0 2156 0 1 29505
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_1
timestamp 1701704242
transform 0 1 1680 1 0 29477
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_2
timestamp 1701704242
transform 0 1 2034 1 0 29465
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_3
timestamp 1701704242
transform 0 -1 1732 1 0 29334
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_4
timestamp 1701704242
transform 1 0 1727 0 -1 29478
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_5
timestamp 1701704242
transform 1 0 1728 0 1 29285
box 0 0 1 1
use M1M2_CDNS_524688791851557  M1M2_CDNS_524688791851557_0
timestamp 1701704242
transform 0 1 5549 1 0 18037
box 0 0 3008 116
use sky130_fd_io__opamp_biasgen_reg_tsg4  sky130_fd_io__opamp_biasgen_reg_tsg4_0
timestamp 1701704242
transform 1 0 5674 0 1 425
box -5997 -6390 10821 22245
use sky130_fd_io__sio_in_ctl_ls_out_reg  sky130_fd_io__sio_in_ctl_ls_out_reg_0
timestamp 1701704242
transform -1 0 13282 0 -1 1518
box -77 0 1861 1066
use sky130_fd_io__sio_pudrvr_reg_csw  sky130_fd_io__sio_pudrvr_reg_csw_0
timestamp 1701704242
transform 1 0 413 0 1 11283
box -209 -133 14151 7362
use sky130_fd_io__sio_pudrvr_reg_leak  sky130_fd_io__sio_pudrvr_reg_leak_0
timestamp 1701704242
transform 1 0 2800 0 1 636
box -3052 -657 8129 1954
use sky130_fd_io__sio_pudrvr_reg_opamp_c  sky130_fd_io__sio_pudrvr_reg_opamp_c_0
timestamp 1701704242
transform 0 1 -1532 1 0 1384
box 1022 1280 13268 16096
use sky130_fd_io__sio_pudrvr_reg_pu  sky130_fd_io__sio_pudrvr_reg_pu_0
timestamp 1701704242
transform 1 0 -16594 0 1 29585
box -401 -12115 26385 6967
use sky130_fd_io__sio_tk_em1o_b_CDNS_524688791851559  sky130_fd_io__sio_tk_em1o_b_CDNS_524688791851559_0
timestamp 1701704242
transform 1 0 -29 0 -1 548
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_b_CDNS_524688791851560  sky130_fd_io__sio_tk_em1s_b_CDNS_524688791851560_0
timestamp 1701704242
transform 0 1 80 1 0 381
box 0 0 1 1
<< labels >>
flabel comment s 1394 2190 1394 2190 0 FreeSans 1000 0 0 0 condiode
flabel comment s 13943 17888 13943 17888 0 FreeSans 400 0 0 0 ModB1X
flabel comment s 13751 17809 13751 17809 0 FreeSans 400 0 0 0 ModB1Y
flabel comment s 12881 510 12881 510 3 FreeSans 200 90 0 0 drvhi_h
flabel metal1 s 7929 1972 7929 1972 0 FreeSans 200 0 0 0 nbias
flabel metal1 s -16902 29735 -16786 29787 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s -16515 29705 -16414 29772 0 FreeSans 200 0 0 0 vgnd
port 12 nsew
flabel metal1 s -16009 29699 -15957 29734 0 FreeSans 200 90 0 0 nghs_h
port 3 nsew
flabel metal1 s -15929 29699 -15877 29734 0 FreeSans 200 90 0 0 pghs_h
port 4 nsew
flabel metal1 s -102 1819 -16 1871 3 FreeSans 200 0 0 0 pu_h_n<0>
port 5 nsew
flabel metal1 s -102 1705 -16 1757 3 FreeSans 200 0 0 0 pu_h_n<1>
port 6 nsew
flabel metal1 s -102 1580 -15 1632 3 FreeSans 200 0 0 0 en_hicc
port 7 nsew
flabel metal1 s -102 356 -5 408 3 FreeSans 200 0 0 0 puen_reg_h
port 8 nsew
flabel metal1 s -102 588 -35 640 3 FreeSans 200 0 0 0 slow_h_n
port 9 nsew
flabel metal1 s -102 496 -33 548 3 FreeSans 200 0 0 0 vreg_en_h
port 10 nsew
flabel metal1 s -296 29755 450 29809 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -1534 29755 -787 29809 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -4418 29755 -3672 29809 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -5656 29755 -4910 29809 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -8541 29755 -7795 29809 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -9779 29727 -9032 29781 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -10716 29727 -10348 29823 3 FreeSans 200 90 0 0 pad
port 11 nsew
flabel metal1 s -10936 29951 -10744 30003 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 639 29727 1600 29781 0 FreeSans 200 0 0 0 vpb_drvr
port 13 nsew
flabel metal1 s -3493 29727 -1757 29781 0 FreeSans 200 0 0 0 vpb_drvr
port 13 nsew
flabel metal1 s -7622 29727 -5887 29781 0 FreeSans 200 0 0 0 vpb_drvr
port 13 nsew
flabel metal1 s -10112 29907 -9920 29940 0 FreeSans 200 0 0 0 vpb_drvr
port 13 nsew
flabel metal1 s 1699 29465 1751 29510 3 FreeSans 200 90 0 0 pug<0>
port 14 nsew
flabel metal1 s 1698 29326 1750 29371 3 FreeSans 200 90 0 0 pug<1>
port 15 nsew
flabel metal4 s -3589 18005 -3164 18876 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal2 s 7852 17872 7852 17872 3 FreeSans 200 90 0 0 vref_nng
flabel metal2 s 14436 17616 14564 17756 7 FreeSans 200 90 0 0 refleak_bias
port 16 nsew
flabel metal2 s 14250 17616 14378 17756 7 FreeSans 200 90 0 0 voutref
port 17 nsew
flabel metal2 s 5195 7294 5325 7346 0 FreeSans 200 0 0 0 fb_in
port 18 nsew
flabel metal2 s 7677 9068 7807 9198 0 FreeSans 200 0 0 0 fb_out
port 19 nsew
flabel metal2 s -252 7199 68 7353 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal2 s 4727 17756 4987 17809 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 7996 17704 8189 17756 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 10093 17710 10286 17756 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 1783 17709 2109 17756 0 FreeSans 200 0 0 0 vgnd
port 12 nsew
flabel metal2 s 5170 17710 5430 17756 0 FreeSans 200 0 0 0 vgnd
port 12 nsew
flabel metal2 s 8317 17710 8582 17756 0 FreeSans 200 0 0 0 vgnd
port 12 nsew
flabel metal2 s 9399 17710 9657 17756 0 FreeSans 200 0 0 0 vgnd
port 12 nsew
flabel metal2 s 3001 17756 3300 17816 0 FreeSans 200 0 0 0 vgnd_io
port 20 nsew
flabel metal2 s -13399 29062 -12677 29204 0 FreeSans 200 0 0 0 vpb_drvr
port 13 nsew
flabel metal2 s 14026 17621 14170 17756 0 FreeSans 200 0 0 0 vpwr_ka
port 21 nsew
<< properties >>
string GDS_END 98937126
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98210084
string path 202.300 106.275 202.300 151.825 
<< end >>
