magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 319 366
<< mvpmos >>
rect 0 0 200 300
<< mvpdiff >>
rect -53 250 0 300
rect -53 216 -45 250
rect -11 216 0 250
rect -53 182 0 216
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 200 250 253 300
rect 200 216 211 250
rect 245 216 253 250
rect 200 182 253 216
rect 200 148 211 182
rect 245 148 253 182
rect 200 114 253 148
rect 200 80 211 114
rect 245 80 253 114
rect 200 46 253 80
rect 200 12 211 46
rect 245 12 253 46
rect 200 0 253 12
<< mvpdiffc >>
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 211 216 245 250
rect 211 148 245 182
rect 211 80 245 114
rect 211 12 245 46
<< poly >>
rect 0 300 200 332
rect 0 -32 200 0
<< locali >>
rect -45 250 -11 266
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 211 250 245 266
rect 211 182 245 216
rect 211 114 245 148
rect 211 46 245 80
rect 211 -4 245 12
use hvDFL1sd_CDNS_52468879185669  hvDFL1sd_CDNS_52468879185669_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185669  hvDFL1sd_CDNS_52468879185669_1
timestamp 1701704242
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
flabel comment s 228 131 228 131 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87825716
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87824698
<< end >>
