magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< pwell >>
rect -76 -26 199 166
<< mvnmos >>
rect 0 0 120 140
<< mvndiff >>
rect -50 0 0 140
rect 120 114 173 140
rect 120 80 131 114
rect 165 80 173 114
rect 120 46 173 80
rect 120 12 131 46
rect 165 12 173 46
rect 120 0 173 12
<< mvndiffc >>
rect 131 80 165 114
rect 131 12 165 46
<< poly >>
rect 0 140 120 166
rect 0 -26 120 0
<< locali >>
rect 131 114 165 130
rect 131 46 165 80
rect 131 -4 165 12
use DFL1sd_CDNS_559591418088  DFL1sd_CDNS_559591418088_0
timestamp 1701704242
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 148 63 148 63 0 FreeSans 300 0 0 0 D
flabel comment s -25 70 -25 70 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 798696
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 797944
<< end >>
