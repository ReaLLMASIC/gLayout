magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< locali >>
rect 7467 50425 7530 50459
rect 7496 50278 7530 50425
rect 11482 50396 11510 50430
rect 7496 50244 7599 50278
rect 7496 50052 7599 50086
rect 7496 49963 7530 50052
rect 7467 49929 7530 49963
rect 11482 49900 11510 49934
rect 7467 49635 7530 49669
rect 7496 49488 7530 49635
rect 11482 49606 11510 49640
rect 7496 49454 7599 49488
rect 7496 49262 7599 49296
rect 7496 49173 7530 49262
rect 7467 49139 7530 49173
rect 11482 49110 11510 49144
rect 7467 48845 7530 48879
rect 7496 48698 7530 48845
rect 11482 48816 11510 48850
rect 7496 48664 7599 48698
rect 7496 48472 7599 48506
rect 7496 48383 7530 48472
rect 7467 48349 7530 48383
rect 11482 48320 11510 48354
rect 7467 48055 7530 48089
rect 7496 47908 7530 48055
rect 11482 48026 11510 48060
rect 7496 47874 7599 47908
rect 7496 47682 7599 47716
rect 7496 47593 7530 47682
rect 7467 47559 7530 47593
rect 11482 47530 11510 47564
rect 7467 47265 7530 47299
rect 7496 47118 7530 47265
rect 11482 47236 11510 47270
rect 7496 47084 7599 47118
rect 7496 46892 7599 46926
rect 7496 46803 7530 46892
rect 7467 46769 7530 46803
rect 11482 46740 11510 46774
rect 7467 46475 7530 46509
rect 7496 46328 7530 46475
rect 11482 46446 11510 46480
rect 7496 46294 7599 46328
rect 7496 46102 7599 46136
rect 7496 46013 7530 46102
rect 7467 45979 7530 46013
rect 11482 45950 11510 45984
rect 7467 45685 7530 45719
rect 7496 45538 7530 45685
rect 11482 45656 11510 45690
rect 7496 45504 7599 45538
rect 7496 45312 7599 45346
rect 7496 45223 7530 45312
rect 7467 45189 7530 45223
rect 11482 45160 11510 45194
rect 7467 44895 7530 44929
rect 7496 44748 7530 44895
rect 11482 44866 11510 44900
rect 7496 44714 7599 44748
rect 7496 44522 7599 44556
rect 7496 44433 7530 44522
rect 7467 44399 7530 44433
rect 11482 44370 11510 44404
rect 7467 44105 7530 44139
rect 7496 43958 7530 44105
rect 11482 44076 11510 44110
rect 7496 43924 7599 43958
rect 7496 43732 7599 43766
rect 7496 43643 7530 43732
rect 7467 43609 7530 43643
rect 11482 43580 11510 43614
rect 7467 43315 7530 43349
rect 7496 43168 7530 43315
rect 11482 43286 11510 43320
rect 7496 43134 7599 43168
rect 7496 42942 7599 42976
rect 7496 42853 7530 42942
rect 7467 42819 7530 42853
rect 11482 42790 11510 42824
rect 7467 42525 7530 42559
rect 7496 42378 7530 42525
rect 11482 42496 11510 42530
rect 7496 42344 7599 42378
rect 7496 42152 7599 42186
rect 7496 42063 7530 42152
rect 7467 42029 7530 42063
rect 11482 42000 11510 42034
rect 7467 41735 7530 41769
rect 7496 41588 7530 41735
rect 11482 41706 11510 41740
rect 7496 41554 7599 41588
rect 7496 41362 7599 41396
rect 7496 41273 7530 41362
rect 7467 41239 7530 41273
rect 11482 41210 11510 41244
rect 7467 40945 7530 40979
rect 7496 40798 7530 40945
rect 11482 40916 11510 40950
rect 7496 40764 7599 40798
rect 7496 40572 7599 40606
rect 7496 40483 7530 40572
rect 7467 40449 7530 40483
rect 11482 40420 11510 40454
rect 7467 40155 7530 40189
rect 7496 40008 7530 40155
rect 11482 40126 11510 40160
rect 7496 39974 7599 40008
rect 7496 39782 7599 39816
rect 7496 39693 7530 39782
rect 7467 39659 7530 39693
rect 11482 39630 11510 39664
rect 7467 39365 7530 39399
rect 7496 39218 7530 39365
rect 11482 39336 11510 39370
rect 7496 39184 7599 39218
rect 7496 38992 7599 39026
rect 7496 38903 7530 38992
rect 7467 38869 7530 38903
rect 11482 38840 11510 38874
rect 7467 38575 7530 38609
rect 7496 38428 7530 38575
rect 11482 38546 11510 38580
rect 7496 38394 7599 38428
rect 7496 38202 7599 38236
rect 7496 38113 7530 38202
rect 7467 38079 7530 38113
rect 11482 38050 11510 38084
rect 7467 37785 7530 37819
rect 7496 37638 7530 37785
rect 11482 37756 11510 37790
rect 7496 37604 7599 37638
rect 7496 37412 7599 37446
rect 7496 37323 7530 37412
rect 7467 37289 7530 37323
rect 11482 37260 11510 37294
rect 7467 36995 7530 37029
rect 7496 36848 7530 36995
rect 11482 36966 11510 37000
rect 7496 36814 7599 36848
rect 7496 36622 7599 36656
rect 7496 36533 7530 36622
rect 7467 36499 7530 36533
rect 11482 36470 11510 36504
rect 7467 36205 7530 36239
rect 7496 36058 7530 36205
rect 11482 36176 11510 36210
rect 7496 36024 7599 36058
rect 7496 35832 7599 35866
rect 7496 35743 7530 35832
rect 7467 35709 7530 35743
rect 11482 35680 11510 35714
rect 7467 35415 7530 35449
rect 7496 35268 7530 35415
rect 11482 35386 11510 35420
rect 7496 35234 7599 35268
rect 7496 35042 7599 35076
rect 7496 34953 7530 35042
rect 7467 34919 7530 34953
rect 11482 34890 11510 34924
rect 7467 34625 7530 34659
rect 7496 34478 7530 34625
rect 11482 34596 11510 34630
rect 7496 34444 7599 34478
rect 7496 34252 7599 34286
rect 7496 34163 7530 34252
rect 7467 34129 7530 34163
rect 11482 34100 11510 34134
rect 7467 33835 7530 33869
rect 7496 33688 7530 33835
rect 11482 33806 11510 33840
rect 7496 33654 7599 33688
rect 7496 33462 7599 33496
rect 7496 33373 7530 33462
rect 7467 33339 7530 33373
rect 11482 33310 11510 33344
rect 7467 33045 7530 33079
rect 7496 32898 7530 33045
rect 11482 33016 11510 33050
rect 7496 32864 7599 32898
rect 7496 32672 7599 32706
rect 7496 32583 7530 32672
rect 7467 32549 7530 32583
rect 11482 32520 11510 32554
rect 7467 32255 7530 32289
rect 7496 32108 7530 32255
rect 11482 32226 11510 32260
rect 7496 32074 7599 32108
rect 7496 31882 7599 31916
rect 7496 31793 7530 31882
rect 7467 31759 7530 31793
rect 11482 31730 11510 31764
rect 7467 31465 7530 31499
rect 7496 31318 7530 31465
rect 11482 31436 11510 31470
rect 7496 31284 7599 31318
rect 7496 31092 7599 31126
rect 7496 31003 7530 31092
rect 7467 30969 7530 31003
rect 11482 30940 11510 30974
rect 7467 30675 7530 30709
rect 7496 30528 7530 30675
rect 11482 30646 11510 30680
rect 7496 30494 7599 30528
rect 7496 30302 7599 30336
rect 7496 30213 7530 30302
rect 7467 30179 7530 30213
rect 11482 30150 11510 30184
rect 7467 29885 7530 29919
rect 7496 29738 7530 29885
rect 11482 29856 11510 29890
rect 7496 29704 7599 29738
rect 7496 29512 7599 29546
rect 7496 29423 7530 29512
rect 7467 29389 7530 29423
rect 11482 29360 11510 29394
rect 7467 29095 7530 29129
rect 7496 28948 7530 29095
rect 11482 29066 11510 29100
rect 7496 28914 7599 28948
rect 7496 28722 7599 28756
rect 7496 28633 7530 28722
rect 7467 28599 7530 28633
rect 11482 28570 11510 28604
rect 7467 28305 7530 28339
rect 7496 28158 7530 28305
rect 11482 28276 11510 28310
rect 7496 28124 7599 28158
rect 7496 27932 7599 27966
rect 7496 27843 7530 27932
rect 7467 27809 7530 27843
rect 11482 27780 11510 27814
rect 7467 27515 7530 27549
rect 7496 27368 7530 27515
rect 11482 27486 11510 27520
rect 7496 27334 7599 27368
rect 7496 27142 7599 27176
rect 7496 27053 7530 27142
rect 7467 27019 7530 27053
rect 11482 26990 11510 27024
rect 7467 26725 7530 26759
rect 7496 26578 7530 26725
rect 11482 26696 11510 26730
rect 7496 26544 7599 26578
rect 7496 26352 7599 26386
rect 7496 26263 7530 26352
rect 7467 26229 7530 26263
rect 11482 26200 11510 26234
rect 7467 25935 7530 25969
rect 7496 25788 7530 25935
rect 11482 25906 11510 25940
rect 7496 25754 7599 25788
rect 7496 25562 7599 25596
rect 7496 25473 7530 25562
rect 7467 25439 7530 25473
rect 11482 25410 11510 25444
rect 7467 25145 7530 25179
rect 7496 24998 7530 25145
rect 11482 25116 11510 25150
rect 7496 24964 7599 24998
rect 7496 24772 7599 24806
rect 7496 24683 7530 24772
rect 7467 24649 7530 24683
rect 11482 24620 11510 24654
rect 7467 24355 7530 24389
rect 7496 24208 7530 24355
rect 11482 24326 11510 24360
rect 7496 24174 7599 24208
rect 7496 23982 7599 24016
rect 7496 23893 7530 23982
rect 7467 23859 7530 23893
rect 11482 23830 11510 23864
rect 7467 23565 7530 23599
rect 7496 23418 7530 23565
rect 11482 23536 11510 23570
rect 7496 23384 7599 23418
rect 7496 23192 7599 23226
rect 7496 23103 7530 23192
rect 7467 23069 7530 23103
rect 11482 23040 11510 23074
rect 7467 22775 7530 22809
rect 7496 22628 7530 22775
rect 11482 22746 11510 22780
rect 7496 22594 7599 22628
rect 7496 22402 7599 22436
rect 7496 22313 7530 22402
rect 7467 22279 7530 22313
rect 11482 22250 11510 22284
rect 7467 21985 7530 22019
rect 7496 21838 7530 21985
rect 11482 21956 11510 21990
rect 7496 21804 7599 21838
rect 7496 21612 7599 21646
rect 7496 21523 7530 21612
rect 7467 21489 7530 21523
rect 11482 21460 11510 21494
rect 7467 21195 7530 21229
rect 7496 21048 7530 21195
rect 11482 21166 11510 21200
rect 7496 21014 7599 21048
rect 7496 20822 7599 20856
rect 7496 20733 7530 20822
rect 7467 20699 7530 20733
rect 11482 20670 11510 20704
rect 7467 20405 7530 20439
rect 7496 20258 7530 20405
rect 11482 20376 11510 20410
rect 7496 20224 7599 20258
rect 7496 20032 7599 20066
rect 7496 19943 7530 20032
rect 7467 19909 7530 19943
rect 11482 19880 11510 19914
rect 7467 19615 7530 19649
rect 7496 19468 7530 19615
rect 11482 19586 11510 19620
rect 7496 19434 7599 19468
rect 7496 19242 7599 19276
rect 7496 19153 7530 19242
rect 7467 19119 7530 19153
rect 11482 19090 11510 19124
rect 7467 18825 7530 18859
rect 7496 18678 7530 18825
rect 11482 18796 11510 18830
rect 7496 18644 7599 18678
rect 7496 18452 7599 18486
rect 7496 18363 7530 18452
rect 7467 18329 7530 18363
rect 11482 18300 11510 18334
rect 7467 18035 7530 18069
rect 7496 17888 7530 18035
rect 11482 18006 11510 18040
rect 7496 17854 7599 17888
rect 7496 17662 7599 17696
rect 7496 17573 7530 17662
rect 7467 17539 7530 17573
rect 11482 17510 11510 17544
rect 7467 17245 7530 17279
rect 7496 17098 7530 17245
rect 11482 17216 11510 17250
rect 7496 17064 7599 17098
rect 7496 16872 7599 16906
rect 7496 16783 7530 16872
rect 7467 16749 7530 16783
rect 11482 16720 11510 16754
rect 7467 16455 7530 16489
rect 7496 16308 7530 16455
rect 11482 16426 11510 16460
rect 7496 16274 7599 16308
rect 7496 16082 7599 16116
rect 7496 15993 7530 16082
rect 7467 15959 7530 15993
rect 11482 15930 11510 15964
rect 7467 15665 7530 15699
rect 7496 15518 7530 15665
rect 11482 15636 11510 15670
rect 7496 15484 7599 15518
rect 7496 15292 7599 15326
rect 7496 15203 7530 15292
rect 7467 15169 7530 15203
rect 11482 15140 11510 15174
rect 7467 14875 7530 14909
rect 7496 14728 7530 14875
rect 11482 14846 11510 14880
rect 7496 14694 7599 14728
rect 7496 14502 7599 14536
rect 7496 14413 7530 14502
rect 7467 14379 7530 14413
rect 11482 14350 11510 14384
rect 7467 14085 7530 14119
rect 7496 13938 7530 14085
rect 11482 14056 11510 14090
rect 7496 13904 7599 13938
rect 7496 13712 7599 13746
rect 7496 13623 7530 13712
rect 7467 13589 7530 13623
rect 11482 13560 11510 13594
rect 7467 13295 7530 13329
rect 7496 13148 7530 13295
rect 11482 13266 11510 13300
rect 7496 13114 7599 13148
rect 7496 12922 7599 12956
rect 7496 12833 7530 12922
rect 7467 12799 7530 12833
rect 11482 12770 11510 12804
rect 7467 12505 7530 12539
rect 7496 12358 7530 12505
rect 11482 12476 11510 12510
rect 7496 12324 7599 12358
rect 7496 12132 7599 12166
rect 7496 12043 7530 12132
rect 7467 12009 7530 12043
rect 11482 11980 11510 12014
rect 7467 11715 7530 11749
rect 7496 11568 7530 11715
rect 11482 11686 11510 11720
rect 7496 11534 7599 11568
rect 7496 11342 7599 11376
rect 7496 11253 7530 11342
rect 7467 11219 7530 11253
rect 11482 11190 11510 11224
rect 7467 10925 7530 10959
rect 7496 10778 7530 10925
rect 11482 10896 11510 10930
rect 7496 10744 7599 10778
rect 7496 10552 7599 10586
rect 7496 10463 7530 10552
rect 7467 10429 7530 10463
rect 11482 10400 11510 10434
rect 7467 10135 7530 10169
rect 7496 9988 7530 10135
rect 11482 10106 11510 10140
rect 7496 9954 7599 9988
rect 7496 9762 7599 9796
rect 7496 9673 7530 9762
rect 7467 9639 7530 9673
rect 11482 9610 11510 9644
rect 7467 9345 7530 9379
rect 7496 9198 7530 9345
rect 11482 9316 11510 9350
rect 7496 9164 7599 9198
rect 7496 8972 7599 9006
rect 7496 8883 7530 8972
rect 7467 8849 7530 8883
rect 11482 8820 11510 8854
rect 7467 8555 7530 8589
rect 7496 8408 7530 8555
rect 11482 8526 11510 8560
rect 7496 8374 7599 8408
rect 7496 8182 7599 8216
rect 7496 8093 7530 8182
rect 7467 8059 7530 8093
rect 11482 8030 11510 8064
rect 7467 7765 7530 7799
rect 7496 7618 7530 7765
rect 11482 7736 11510 7770
rect 7496 7584 7599 7618
rect 7496 7392 7599 7426
rect 7496 7303 7530 7392
rect 7467 7269 7530 7303
rect 11482 7240 11510 7274
rect 7467 6975 7530 7009
rect 7496 6828 7530 6975
rect 11482 6946 11510 6980
rect 7496 6794 7599 6828
rect 7496 6602 7599 6636
rect 7496 6513 7530 6602
rect 7467 6479 7530 6513
rect 11482 6450 11510 6484
rect 7467 6185 7530 6219
rect 7496 6038 7530 6185
rect 11482 6156 11510 6190
rect 7496 6004 7599 6038
rect 7496 5812 7599 5846
rect 7496 5723 7530 5812
rect 7467 5689 7530 5723
rect 11482 5660 11510 5694
rect 7467 5395 7530 5429
rect 7496 5248 7530 5395
rect 11482 5366 11510 5400
rect 7496 5214 7599 5248
rect 7496 5022 7599 5056
rect 7496 4933 7530 5022
rect 7467 4899 7530 4933
rect 11482 4870 11510 4904
rect 7467 4605 7530 4639
rect 7496 4458 7530 4605
rect 11482 4576 11510 4610
rect 7496 4424 7599 4458
rect 7496 4232 7599 4266
rect 7496 4143 7530 4232
rect 7467 4109 7530 4143
rect 11482 4080 11510 4114
rect 7467 3815 7530 3849
rect 7496 3668 7530 3815
rect 11482 3786 11510 3820
rect 7496 3634 7599 3668
rect 7496 3442 7599 3476
rect 7496 3353 7530 3442
rect 7467 3319 7530 3353
rect 11482 3290 11510 3324
rect 7467 3025 7530 3059
rect 7496 2878 7530 3025
rect 11482 2996 11510 3030
rect 7496 2844 7599 2878
rect 7496 2652 7599 2686
rect 7496 2563 7530 2652
rect 7467 2529 7530 2563
rect 11482 2500 11510 2534
rect 7467 2235 7530 2269
rect 7496 2088 7530 2235
rect 11482 2206 11510 2240
rect 7496 2054 7599 2088
rect 7496 1862 7599 1896
rect 7496 1773 7530 1862
rect 7467 1739 7530 1773
rect 11482 1710 11510 1744
rect 7467 1445 7530 1479
rect 7496 1298 7530 1445
rect 11482 1416 11510 1450
rect 7496 1264 7599 1298
rect 7496 1072 7599 1106
rect 7496 983 7530 1072
rect 7467 949 7530 983
rect 11482 920 11510 954
rect 7467 655 7530 689
rect 7496 508 7530 655
rect 11482 626 11510 660
rect 7496 474 7599 508
rect 7496 282 7599 316
rect 7496 193 7530 282
rect 7467 159 7530 193
rect 11482 130 11510 164
<< metal1 >>
rect 7750 25239 7756 25291
rect 7808 25239 7814 25291
rect 8175 25238 8181 25290
rect 8233 25238 8239 25290
rect 9218 25254 9224 25306
rect 9276 25254 9282 25306
rect 10742 25254 10748 25306
rect 10800 25254 10806 25306
rect 18 29 46 7929
rect 98 29 126 7929
rect 178 29 206 7929
rect 258 29 286 7929
rect 338 29 366 7929
rect 418 29 446 7929
rect 498 29 526 7929
<< via1 >>
rect 7756 25239 7808 25291
rect 8181 25238 8233 25290
rect 9224 25254 9276 25306
rect 10748 25254 10800 25306
<< metal2 >>
rect 7582 0 7610 50560
rect 9222 25308 9278 25317
rect 7754 25293 7810 25302
rect 7754 25228 7810 25237
rect 8179 25292 8235 25301
rect 9222 25243 9278 25252
rect 10746 25308 10802 25317
rect 10746 25243 10802 25252
rect 8179 25227 8235 25236
<< via2 >>
rect 9222 25306 9278 25308
rect 7754 25291 7810 25293
rect 7754 25239 7756 25291
rect 7756 25239 7808 25291
rect 7808 25239 7810 25291
rect 7754 25237 7810 25239
rect 8179 25290 8235 25292
rect 8179 25238 8181 25290
rect 8181 25238 8233 25290
rect 8233 25238 8235 25290
rect 9222 25254 9224 25306
rect 9224 25254 9276 25306
rect 9276 25254 9278 25306
rect 9222 25252 9278 25254
rect 10746 25306 10802 25308
rect 10746 25254 10748 25306
rect 10748 25254 10800 25306
rect 10800 25254 10802 25306
rect 10746 25252 10802 25254
rect 8179 25236 8235 25238
<< metal3 >>
rect 5776 50168 5874 50266
rect 6201 50168 6299 50266
rect 6633 50168 6731 50266
rect 7015 50145 7113 50243
rect 7287 50145 7385 50243
rect 5776 49794 5874 49892
rect 6201 49736 6299 49834
rect 6633 49736 6731 49834
rect 7015 49750 7113 49848
rect 7287 49750 7385 49848
rect 5776 49378 5874 49476
rect 6201 49378 6299 49476
rect 6633 49378 6731 49476
rect 7015 49355 7113 49453
rect 7287 49355 7382 49453
rect 5776 49004 5874 49102
rect 6201 48946 6299 49044
rect 6633 48946 6731 49044
rect 7015 48960 7113 49058
rect 7287 48960 7385 49058
rect 5776 48588 5874 48686
rect 6201 48588 6299 48686
rect 6633 48588 6731 48686
rect 7015 48565 7113 48663
rect 7287 48565 7385 48663
rect 5776 48214 5874 48312
rect 6201 48156 6299 48254
rect 6633 48156 6731 48254
rect 7015 48170 7113 48268
rect 7287 48170 7385 48268
rect 5776 47798 5874 47896
rect 6201 47798 6299 47896
rect 6633 47798 6731 47896
rect 7015 47775 7113 47873
rect 7287 47775 7385 47873
rect 5776 47424 5874 47522
rect 6201 47366 6299 47464
rect 6633 47366 6731 47464
rect 7015 47380 7113 47478
rect 7287 47380 7385 47478
rect 5776 47008 5874 47106
rect 6201 47008 6299 47106
rect 6633 47008 6731 47106
rect 7015 46985 7113 47083
rect 7287 46985 7385 47083
rect 5776 46634 5874 46732
rect 6201 46576 6299 46674
rect 6633 46576 6731 46674
rect 7015 46590 7113 46688
rect 7287 46590 7385 46688
rect 5776 46218 5874 46316
rect 6201 46218 6299 46316
rect 6633 46218 6731 46316
rect 7015 46195 7113 46293
rect 7287 46195 7385 46293
rect 5776 45844 5874 45942
rect 6201 45786 6299 45884
rect 6633 45786 6731 45884
rect 7015 45800 7113 45898
rect 7287 45800 7385 45898
rect 5776 45428 5874 45526
rect 6201 45428 6299 45526
rect 6633 45428 6731 45526
rect 7015 45405 7113 45503
rect 7287 45405 7385 45503
rect 5776 45054 5874 45152
rect 6201 44996 6299 45094
rect 6633 44996 6731 45094
rect 7015 45010 7113 45108
rect 7287 45010 7385 45108
rect 5776 44638 5874 44736
rect 6201 44638 6299 44736
rect 6633 44638 6731 44736
rect 7015 44615 7113 44713
rect 7287 44615 7385 44713
rect 5776 44264 5874 44362
rect 6201 44206 6299 44304
rect 6633 44206 6731 44304
rect 7015 44220 7113 44318
rect 7287 44220 7385 44318
rect 5776 43848 5874 43946
rect 6201 43848 6299 43946
rect 6633 43848 6731 43946
rect 7015 43825 7113 43923
rect 7287 43825 7385 43923
rect 5776 43474 5874 43572
rect 6201 43416 6299 43514
rect 6633 43416 6731 43514
rect 7015 43430 7113 43528
rect 7287 43430 7385 43528
rect 5776 43058 5874 43156
rect 6201 43058 6299 43156
rect 6633 43058 6731 43156
rect 7015 43035 7113 43133
rect 7287 43035 7385 43133
rect 5776 42684 5874 42782
rect 6201 42626 6299 42724
rect 6633 42626 6731 42724
rect 7015 42640 7113 42738
rect 7287 42640 7385 42738
rect 5776 42268 5874 42366
rect 6201 42268 6299 42366
rect 6633 42268 6731 42366
rect 7015 42245 7113 42343
rect 7287 42245 7385 42343
rect 5776 41894 5874 41992
rect 6201 41836 6299 41934
rect 6633 41836 6731 41934
rect 7015 41850 7113 41948
rect 7287 41850 7385 41948
rect 5776 41478 5874 41576
rect 6201 41478 6299 41576
rect 6633 41478 6731 41576
rect 7015 41455 7113 41553
rect 7287 41455 7385 41553
rect 5776 41104 5874 41202
rect 6201 41046 6299 41144
rect 6633 41046 6731 41144
rect 7015 41060 7113 41158
rect 7287 41060 7385 41158
rect 5776 40688 5874 40786
rect 6201 40688 6299 40786
rect 6633 40688 6731 40786
rect 7015 40665 7113 40763
rect 7287 40665 7385 40763
rect 5776 40314 5874 40412
rect 6201 40256 6299 40354
rect 6633 40256 6731 40354
rect 7015 40270 7113 40368
rect 7287 40270 7385 40368
rect 5776 39898 5874 39996
rect 6201 39898 6299 39996
rect 6633 39898 6731 39996
rect 7015 39875 7113 39973
rect 7287 39875 7385 39973
rect 5776 39524 5874 39622
rect 6201 39466 6299 39564
rect 6633 39466 6731 39564
rect 7015 39480 7113 39578
rect 7287 39480 7385 39578
rect 5776 39108 5874 39206
rect 6201 39108 6299 39206
rect 6633 39108 6731 39206
rect 7015 39085 7113 39183
rect 7287 39085 7385 39183
rect 5776 38734 5874 38832
rect 6201 38676 6299 38774
rect 6633 38676 6731 38774
rect 7015 38690 7113 38788
rect 7287 38690 7385 38788
rect 5776 38318 5874 38416
rect 6201 38318 6299 38416
rect 6633 38318 6731 38416
rect 7015 38295 7113 38393
rect 7287 38295 7385 38393
rect 5776 37944 5874 38042
rect 6201 37886 6299 37984
rect 6633 37886 6731 37984
rect 7015 37900 7113 37998
rect 7287 37900 7385 37998
rect 5776 37528 5874 37626
rect 6201 37528 6299 37626
rect 6633 37528 6731 37626
rect 7015 37505 7113 37603
rect 7287 37505 7385 37603
rect 5776 37154 5874 37252
rect 6201 37096 6299 37194
rect 6633 37096 6731 37194
rect 7015 37110 7113 37208
rect 7287 37110 7385 37208
rect 5776 36738 5874 36836
rect 6201 36738 6299 36836
rect 6633 36738 6731 36836
rect 7015 36715 7113 36813
rect 7287 36715 7385 36813
rect 5776 36364 5874 36462
rect 6201 36306 6299 36404
rect 6633 36306 6731 36404
rect 7015 36320 7113 36418
rect 7287 36320 7385 36418
rect 5776 35948 5874 36046
rect 6201 35948 6299 36046
rect 6633 35948 6731 36046
rect 7015 35925 7113 36023
rect 7287 35925 7385 36023
rect 5776 35574 5874 35672
rect 6201 35516 6299 35614
rect 6633 35516 6731 35614
rect 7015 35530 7113 35628
rect 7287 35530 7385 35628
rect 5776 35158 5874 35256
rect 6201 35158 6299 35256
rect 6633 35158 6731 35256
rect 7015 35135 7113 35233
rect 7287 35135 7385 35233
rect 5776 34784 5874 34882
rect 6201 34726 6299 34824
rect 6633 34726 6731 34824
rect 7015 34740 7113 34838
rect 7287 34740 7385 34838
rect 5776 34368 5874 34466
rect 6201 34368 6299 34466
rect 6633 34368 6731 34466
rect 7015 34345 7113 34443
rect 7287 34345 7385 34443
rect 5776 33994 5874 34092
rect 6201 33936 6299 34034
rect 6633 33936 6731 34034
rect 7015 33950 7113 34048
rect 7287 33950 7385 34048
rect 5776 33578 5874 33676
rect 6201 33578 6299 33676
rect 6633 33578 6731 33676
rect 7015 33555 7113 33653
rect 7287 33555 7385 33653
rect 5776 33204 5874 33302
rect 6201 33146 6299 33244
rect 6633 33146 6731 33244
rect 7015 33160 7113 33258
rect 7287 33160 7385 33258
rect 5776 32788 5874 32886
rect 6201 32788 6299 32886
rect 6633 32788 6731 32886
rect 7015 32765 7113 32863
rect 7287 32765 7385 32863
rect 5776 32414 5874 32512
rect 6201 32356 6299 32454
rect 6633 32356 6731 32454
rect 7015 32370 7113 32468
rect 7287 32370 7385 32468
rect 5776 31998 5874 32096
rect 6201 31998 6299 32096
rect 6633 31998 6731 32096
rect 7015 31975 7113 32073
rect 7287 31975 7385 32073
rect 5776 31624 5874 31722
rect 6201 31566 6299 31664
rect 6633 31566 6731 31664
rect 7015 31580 7113 31678
rect 7287 31580 7385 31678
rect 5776 31208 5874 31306
rect 6201 31208 6299 31306
rect 6633 31208 6731 31306
rect 7015 31185 7113 31283
rect 7287 31185 7385 31283
rect 5776 30834 5874 30932
rect 6201 30776 6299 30874
rect 6633 30776 6731 30874
rect 7015 30790 7113 30888
rect 7287 30790 7385 30888
rect 5776 30418 5874 30516
rect 6201 30418 6299 30516
rect 6633 30418 6731 30516
rect 7015 30395 7113 30493
rect 7287 30395 7385 30493
rect 5776 30044 5874 30142
rect 6201 29986 6299 30084
rect 6633 29986 6731 30084
rect 7015 30000 7113 30098
rect 7287 30000 7385 30098
rect 5776 29628 5874 29726
rect 6201 29628 6299 29726
rect 6633 29628 6731 29726
rect 7015 29605 7113 29703
rect 7287 29605 7385 29703
rect 5776 29254 5874 29352
rect 6201 29196 6299 29294
rect 6633 29196 6731 29294
rect 7015 29210 7113 29308
rect 7287 29210 7385 29308
rect 5776 28838 5874 28936
rect 6201 28838 6299 28936
rect 6633 28838 6731 28936
rect 7015 28815 7113 28913
rect 7287 28815 7385 28913
rect 5776 28464 5874 28562
rect 6201 28406 6299 28504
rect 6633 28406 6731 28504
rect 7015 28420 7113 28518
rect 7287 28420 7385 28518
rect 5776 28048 5874 28146
rect 6201 28048 6299 28146
rect 6633 28048 6731 28146
rect 7015 28025 7113 28123
rect 7287 28025 7385 28123
rect 5776 27674 5874 27772
rect 6201 27616 6299 27714
rect 6633 27616 6731 27714
rect 7015 27630 7113 27728
rect 7287 27630 7385 27728
rect 5776 27258 5874 27356
rect 6201 27258 6299 27356
rect 6633 27258 6731 27356
rect 7015 27235 7113 27333
rect 7287 27235 7385 27333
rect 5776 26884 5874 26982
rect 6201 26826 6299 26924
rect 6633 26826 6731 26924
rect 7015 26840 7113 26938
rect 7287 26840 7385 26938
rect 5776 26468 5874 26566
rect 6201 26468 6299 26566
rect 6633 26468 6731 26566
rect 7015 26445 7113 26543
rect 7287 26445 7385 26543
rect 5776 26094 5874 26192
rect 6201 26036 6299 26134
rect 6633 26036 6731 26134
rect 7015 26050 7113 26148
rect 7287 26050 7385 26148
rect 5776 25678 5874 25776
rect 6201 25678 6299 25776
rect 6633 25678 6731 25776
rect 7015 25655 7113 25753
rect 7287 25655 7385 25753
rect 5776 25304 5874 25402
rect 6201 25246 6299 25344
rect 6633 25246 6731 25344
rect 7015 25260 7113 25358
rect 7287 25260 7385 25358
rect 7733 25293 7831 25314
rect 7733 25237 7754 25293
rect 7810 25237 7831 25293
rect 7733 25216 7831 25237
rect 8158 25292 8256 25313
rect 8158 25236 8179 25292
rect 8235 25236 8256 25292
rect 8158 25215 8256 25236
rect 9201 25308 9299 25329
rect 9201 25252 9222 25308
rect 9278 25252 9299 25308
rect 9201 25231 9299 25252
rect 10725 25308 10823 25329
rect 10725 25252 10746 25308
rect 10802 25252 10823 25308
rect 10725 25231 10823 25252
rect 5776 24888 5874 24986
rect 6201 24888 6299 24986
rect 6633 24888 6731 24986
rect 7015 24865 7113 24963
rect 7287 24865 7385 24963
rect 5776 24514 5874 24612
rect 6201 24456 6299 24554
rect 6633 24456 6731 24554
rect 7015 24470 7113 24568
rect 7287 24470 7385 24568
rect 5776 24098 5874 24196
rect 6201 24098 6299 24196
rect 6633 24098 6731 24196
rect 7015 24075 7113 24173
rect 7287 24075 7385 24173
rect 5776 23724 5874 23822
rect 6201 23666 6299 23764
rect 6633 23666 6731 23764
rect 7015 23680 7113 23778
rect 7287 23680 7385 23778
rect 5776 23308 5874 23406
rect 6201 23308 6299 23406
rect 6633 23308 6731 23406
rect 7015 23285 7113 23383
rect 7287 23285 7385 23383
rect 5776 22934 5874 23032
rect 6201 22876 6299 22974
rect 6633 22876 6731 22974
rect 7015 22890 7113 22988
rect 7287 22890 7385 22988
rect 5776 22518 5874 22616
rect 6201 22518 6299 22616
rect 6633 22518 6731 22616
rect 7015 22495 7113 22593
rect 7287 22495 7385 22593
rect 5776 22144 5874 22242
rect 6201 22086 6299 22184
rect 6633 22086 6731 22184
rect 7015 22100 7113 22198
rect 7287 22100 7385 22198
rect 5776 21728 5874 21826
rect 6201 21728 6299 21826
rect 6633 21728 6731 21826
rect 7015 21705 7113 21803
rect 7287 21705 7385 21803
rect 5776 21354 5874 21452
rect 6201 21296 6299 21394
rect 6633 21296 6731 21394
rect 7015 21310 7113 21408
rect 7287 21310 7385 21408
rect 5776 20938 5874 21036
rect 6201 20938 6299 21036
rect 6633 20938 6731 21036
rect 7015 20915 7113 21013
rect 7287 20915 7385 21013
rect 5776 20564 5874 20662
rect 6201 20506 6299 20604
rect 6633 20506 6731 20604
rect 7015 20520 7113 20618
rect 7287 20520 7385 20618
rect 5776 20148 5874 20246
rect 6201 20148 6299 20246
rect 6633 20148 6731 20246
rect 7015 20125 7113 20223
rect 7287 20125 7385 20223
rect 5776 19774 5874 19872
rect 6201 19716 6299 19814
rect 6633 19716 6731 19814
rect 7015 19730 7113 19828
rect 7287 19730 7385 19828
rect 5776 19358 5874 19456
rect 6201 19358 6299 19456
rect 6633 19358 6731 19456
rect 7015 19335 7113 19433
rect 7287 19335 7385 19433
rect 5776 18984 5874 19082
rect 6201 18926 6299 19024
rect 6633 18926 6731 19024
rect 7015 18940 7113 19038
rect 7287 18940 7385 19038
rect 5776 18568 5874 18666
rect 6201 18568 6299 18666
rect 6633 18568 6731 18666
rect 7015 18545 7113 18643
rect 7287 18545 7385 18643
rect 5776 18194 5874 18292
rect 6201 18136 6299 18234
rect 6633 18136 6731 18234
rect 7015 18150 7113 18248
rect 7287 18150 7385 18248
rect 5776 17778 5874 17876
rect 6201 17778 6299 17876
rect 6633 17778 6731 17876
rect 7015 17755 7113 17853
rect 7287 17755 7385 17853
rect 5776 17404 5874 17502
rect 6201 17346 6299 17444
rect 6633 17346 6731 17444
rect 7015 17360 7113 17458
rect 7287 17360 7385 17458
rect 5776 16988 5874 17086
rect 6201 16988 6299 17086
rect 6633 16988 6731 17086
rect 7015 16965 7113 17063
rect 7287 16965 7382 17063
rect 5776 16614 5874 16712
rect 6201 16556 6299 16654
rect 6633 16556 6731 16654
rect 7015 16570 7113 16668
rect 7287 16570 7385 16668
rect 5776 16198 5874 16296
rect 6201 16198 6299 16296
rect 6633 16198 6731 16296
rect 7015 16175 7113 16273
rect 7287 16175 7385 16273
rect 5776 15824 5874 15922
rect 6201 15766 6299 15864
rect 6633 15766 6731 15864
rect 7015 15780 7113 15878
rect 7287 15780 7385 15878
rect 5776 15408 5874 15506
rect 6201 15408 6299 15506
rect 6633 15408 6731 15506
rect 7015 15385 7113 15483
rect 7287 15385 7385 15483
rect 5776 15034 5874 15132
rect 6201 14976 6299 15074
rect 6633 14976 6731 15074
rect 7015 14990 7113 15088
rect 7287 14990 7385 15088
rect 5776 14618 5874 14716
rect 6201 14618 6299 14716
rect 6633 14618 6731 14716
rect 7015 14595 7113 14693
rect 7287 14595 7385 14693
rect 5776 14244 5874 14342
rect 6201 14186 6299 14284
rect 6633 14186 6731 14284
rect 7015 14200 7113 14298
rect 7287 14200 7385 14298
rect 5776 13828 5874 13926
rect 6201 13828 6299 13926
rect 6633 13828 6731 13926
rect 7015 13805 7113 13903
rect 7287 13805 7385 13903
rect 5776 13454 5874 13552
rect 6201 13396 6299 13494
rect 6633 13396 6731 13494
rect 7015 13410 7113 13508
rect 7287 13410 7385 13508
rect 5776 13038 5874 13136
rect 6201 13038 6299 13136
rect 6633 13038 6731 13136
rect 7015 13015 7113 13113
rect 7287 13015 7385 13113
rect 5776 12664 5874 12762
rect 6201 12606 6299 12704
rect 6633 12606 6731 12704
rect 7015 12620 7113 12718
rect 7287 12620 7385 12718
rect 5776 12248 5874 12346
rect 6201 12248 6299 12346
rect 6633 12248 6731 12346
rect 7015 12225 7113 12323
rect 7287 12225 7385 12323
rect 5776 11874 5874 11972
rect 6201 11816 6299 11914
rect 6633 11816 6731 11914
rect 7015 11830 7113 11928
rect 7287 11830 7385 11928
rect 5776 11458 5874 11556
rect 6201 11458 6299 11556
rect 6633 11458 6731 11556
rect 7015 11435 7113 11533
rect 7287 11435 7385 11533
rect 5776 11084 5874 11182
rect 6201 11026 6299 11124
rect 6633 11026 6731 11124
rect 7015 11040 7113 11138
rect 7287 11040 7385 11138
rect 5776 10668 5874 10766
rect 6201 10668 6299 10766
rect 6633 10668 6731 10766
rect 7015 10645 7113 10743
rect 7287 10645 7385 10743
rect 5776 10294 5874 10392
rect 6201 10236 6299 10334
rect 6633 10236 6731 10334
rect 7015 10250 7113 10348
rect 7287 10250 7385 10348
rect 5776 9878 5874 9976
rect 6201 9878 6299 9976
rect 6633 9878 6731 9976
rect 7015 9855 7113 9953
rect 7287 9855 7385 9953
rect 5776 9504 5874 9602
rect 6201 9446 6299 9544
rect 6633 9446 6731 9544
rect 7015 9460 7113 9558
rect 7287 9460 7385 9558
rect 5776 9088 5874 9186
rect 6201 9088 6299 9186
rect 6633 9088 6731 9186
rect 7015 9065 7113 9163
rect 7287 9065 7385 9163
rect 5776 8714 5874 8812
rect 6201 8656 6299 8754
rect 6633 8656 6731 8754
rect 7015 8670 7113 8768
rect 7287 8670 7385 8768
rect 5776 8298 5874 8396
rect 6201 8298 6299 8396
rect 6633 8298 6731 8396
rect 7015 8275 7113 8373
rect 7287 8275 7385 8373
rect 5776 7924 5874 8022
rect 6201 7866 6299 7964
rect 6633 7866 6731 7964
rect 7015 7880 7113 7978
rect 7287 7880 7385 7978
rect 2486 7508 2584 7606
rect 2911 7508 3009 7606
rect 3343 7508 3441 7606
rect 3725 7485 3823 7583
rect 3997 7485 4095 7583
rect 5776 7508 5874 7606
rect 6201 7508 6299 7606
rect 6633 7508 6731 7606
rect 7015 7485 7113 7583
rect 7287 7485 7385 7583
rect 5776 7134 5874 7232
rect 6201 7076 6299 7174
rect 6633 7076 6731 7174
rect 7015 7090 7113 7188
rect 7287 7090 7385 7188
rect 2486 6718 2584 6816
rect 2911 6718 3009 6816
rect 3343 6718 3441 6816
rect 3725 6695 3823 6793
rect 3997 6695 4095 6793
rect 5776 6718 5874 6816
rect 6201 6718 6299 6816
rect 6633 6718 6731 6816
rect 7015 6695 7113 6793
rect 7287 6695 7385 6793
rect 5776 6344 5874 6442
rect 6201 6286 6299 6384
rect 6633 6286 6731 6384
rect 7015 6300 7113 6398
rect 7287 6300 7385 6398
rect 2486 5928 2584 6026
rect 2911 5928 3009 6026
rect 3343 5928 3441 6026
rect 3725 5905 3823 6003
rect 3997 5905 4095 6003
rect 5776 5928 5874 6026
rect 6201 5928 6299 6026
rect 6633 5928 6731 6026
rect 7015 5905 7113 6003
rect 7287 5905 7385 6003
rect 5776 5554 5874 5652
rect 6201 5496 6299 5594
rect 6633 5496 6731 5594
rect 7015 5510 7113 5608
rect 7287 5510 7385 5608
rect 1155 5115 1253 5213
rect 1427 5115 1525 5213
rect 2486 5138 2584 5236
rect 2911 5138 3009 5236
rect 3343 5138 3441 5236
rect 3725 5115 3823 5213
rect 3997 5115 4095 5213
rect 5776 5138 5874 5236
rect 6201 5138 6299 5236
rect 6633 5138 6731 5236
rect 7015 5115 7113 5213
rect 7287 5115 7385 5213
rect 5776 4764 5874 4862
rect 6201 4706 6299 4804
rect 6633 4706 6731 4804
rect 7015 4720 7113 4818
rect 7287 4720 7385 4818
rect 5776 4348 5874 4446
rect 6201 4348 6299 4446
rect 6633 4348 6731 4446
rect 7015 4325 7113 4423
rect 7287 4325 7385 4423
rect 5776 3974 5874 4072
rect 6201 3916 6299 4014
rect 6633 3916 6731 4014
rect 7015 3930 7113 4028
rect 7287 3930 7385 4028
rect 2921 3542 3019 3640
rect 3346 3542 3444 3640
rect 3725 3535 3823 3633
rect 3997 3535 4095 3633
rect 5776 3558 5874 3656
rect 6201 3558 6299 3656
rect 6633 3558 6731 3656
rect 7015 3535 7113 3633
rect 7287 3535 7385 3633
rect 5776 3184 5874 3282
rect 6201 3126 6299 3224
rect 6633 3126 6731 3224
rect 7015 3140 7113 3238
rect 7287 3140 7385 3238
rect 1751 2745 1849 2843
rect 2023 2745 2121 2843
rect 2921 2752 3019 2850
rect 3346 2752 3444 2850
rect 3725 2745 3823 2843
rect 3997 2745 4095 2843
rect 5776 2768 5874 2866
rect 6201 2768 6299 2866
rect 6633 2768 6731 2866
rect 7015 2745 7113 2843
rect 7287 2745 7385 2843
rect 5776 2394 5874 2492
rect 6201 2336 6299 2434
rect 6633 2336 6731 2434
rect 7015 2350 7113 2448
rect 7287 2350 7385 2448
rect 5776 1978 5874 2076
rect 6201 1978 6299 2076
rect 6633 1978 6731 2076
rect 7015 1955 7113 2053
rect 7287 1955 7385 2053
rect 5776 1604 5874 1702
rect 6201 1546 6299 1644
rect 6633 1546 6731 1644
rect 7015 1560 7113 1658
rect 7287 1560 7385 1658
rect 2921 1172 3019 1270
rect 3346 1172 3444 1270
rect 3725 1165 3823 1263
rect 3997 1165 4095 1263
rect 5776 1188 5874 1286
rect 6201 1188 6299 1286
rect 6633 1188 6731 1286
rect 7015 1165 7113 1263
rect 7287 1165 7385 1263
rect 5776 814 5874 912
rect 6201 756 6299 854
rect 6633 756 6731 854
rect 7015 770 7113 868
rect 7287 770 7385 868
rect 1751 375 1849 473
rect 2023 375 2121 473
rect 2921 382 3019 480
rect 3346 382 3444 480
rect 3725 375 3823 473
rect 3997 375 4095 473
rect 5776 398 5874 496
rect 6201 398 6299 496
rect 6633 398 6731 496
rect 7015 375 7113 473
rect 7287 375 7385 473
use contact_8  contact_8_0
timestamp 1701704242
transform 1 0 7750 0 1 25233
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1701704242
transform 1 0 9218 0 1 25248
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1701704242
transform 1 0 8175 0 1 25232
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1701704242
transform 1 0 10742 0 1 25248
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1701704242
transform 1 0 7749 0 1 25228
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1701704242
transform 1 0 9217 0 1 25243
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1701704242
transform 1 0 8174 0 1 25227
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1701704242
transform 1 0 10741 0 1 25243
box 0 0 1 1
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1701704242
transform 1 0 0 0 1 0
box 0 -31 7502 50649
use wordline_driver_array  wordline_driver_array_0
timestamp 1701704242
transform 1 0 7512 0 1 0
box 70 -56 4016 50616
<< labels >>
rlabel locali s 11496 38563 11496 38563 4 wl_97
port 106 nsew
rlabel locali s 11496 34613 11496 34613 4 wl_87
port 96 nsew
rlabel locali s 11496 42017 11496 42017 4 wl_106
port 115 nsew
rlabel locali s 11496 35697 11496 35697 4 wl_90
port 99 nsew
rlabel locali s 11496 42807 11496 42807 4 wl_108
port 117 nsew
rlabel locali s 11496 36983 11496 36983 4 wl_93
port 102 nsew
rlabel locali s 11496 48833 11496 48833 4 wl_123
port 132 nsew
rlabel locali s 11496 28293 11496 28293 4 wl_71
port 80 nsew
rlabel locali s 11496 25923 11496 25923 4 wl_65
port 74 nsew
rlabel locali s 11496 33327 11496 33327 4 wl_84
port 93 nsew
rlabel locali s 11496 39647 11496 39647 4 wl_100
port 109 nsew
rlabel locali s 11496 29083 11496 29083 4 wl_73
port 82 nsew
rlabel locali s 11496 28587 11496 28587 4 wl_72
port 81 nsew
rlabel locali s 11496 41227 11496 41227 4 wl_104
port 113 nsew
rlabel locali s 11496 27007 11496 27007 4 wl_68
port 77 nsew
rlabel locali s 11496 46757 11496 46757 4 wl_118
port 127 nsew
rlabel locali s 11496 45177 11496 45177 4 wl_114
port 123 nsew
rlabel locali s 11496 32243 11496 32243 4 wl_81
port 90 nsew
rlabel locali s 11496 45967 11496 45967 4 wl_116
port 125 nsew
rlabel locali s 11496 43597 11496 43597 4 wl_110
port 119 nsew
rlabel locali s 11496 33823 11496 33823 4 wl_85
port 94 nsew
rlabel locali s 11496 33033 11496 33033 4 wl_83
port 92 nsew
rlabel locali s 11496 39353 11496 39353 4 wl_99
port 108 nsew
rlabel locali s 11496 36193 11496 36193 4 wl_91
port 100 nsew
rlabel locali s 11496 38857 11496 38857 4 wl_98
port 107 nsew
rlabel locali s 11496 42513 11496 42513 4 wl_107
port 116 nsew
rlabel locali s 11496 30663 11496 30663 4 wl_77
port 86 nsew
rlabel locali s 11496 44387 11496 44387 4 wl_112
port 121 nsew
rlabel locali s 11496 38067 11496 38067 4 wl_96
port 105 nsew
rlabel locali s 11496 27503 11496 27503 4 wl_69
port 78 nsew
rlabel locali s 11496 46463 11496 46463 4 wl_117
port 126 nsew
rlabel locali s 11496 37277 11496 37277 4 wl_94
port 103 nsew
rlabel locali s 11496 50413 11496 50413 4 wl_127
port 136 nsew
rlabel locali s 11496 45673 11496 45673 4 wl_115
port 124 nsew
rlabel locali s 11496 26713 11496 26713 4 wl_67
port 76 nsew
rlabel locali s 11496 36487 11496 36487 4 wl_92
port 101 nsew
rlabel locali s 11496 44883 11496 44883 4 wl_113
port 122 nsew
rlabel locali s 11496 48337 11496 48337 4 wl_122
port 131 nsew
rlabel locali s 11496 49917 11496 49917 4 wl_126
port 135 nsew
rlabel locali s 11496 40437 11496 40437 4 wl_102
port 111 nsew
rlabel locali s 11496 30957 11496 30957 4 wl_78
port 87 nsew
rlabel locali s 11496 34117 11496 34117 4 wl_86
port 95 nsew
rlabel locali s 11496 26217 11496 26217 4 wl_66
port 75 nsew
rlabel locali s 11496 31747 11496 31747 4 wl_80
port 89 nsew
rlabel locali s 11496 37773 11496 37773 4 wl_95
port 104 nsew
rlabel locali s 11496 49127 11496 49127 4 wl_124
port 133 nsew
rlabel locali s 11496 25427 11496 25427 4 wl_64
port 73 nsew
rlabel locali s 11496 40933 11496 40933 4 wl_103
port 112 nsew
rlabel locali s 11496 32537 11496 32537 4 wl_82
port 91 nsew
rlabel locali s 11496 47253 11496 47253 4 wl_119
port 128 nsew
rlabel locali s 11496 31453 11496 31453 4 wl_79
port 88 nsew
rlabel locali s 11496 49623 11496 49623 4 wl_125
port 134 nsew
rlabel locali s 11496 29873 11496 29873 4 wl_75
port 84 nsew
rlabel locali s 11496 41723 11496 41723 4 wl_105
port 114 nsew
rlabel locali s 11496 48043 11496 48043 4 wl_121
port 130 nsew
rlabel locali s 11496 30167 11496 30167 4 wl_76
port 85 nsew
rlabel locali s 11496 27797 11496 27797 4 wl_70
port 79 nsew
rlabel locali s 11496 47547 11496 47547 4 wl_120
port 129 nsew
rlabel locali s 11496 44093 11496 44093 4 wl_111
port 120 nsew
rlabel locali s 11496 29377 11496 29377 4 wl_74
port 83 nsew
rlabel locali s 11496 43303 11496 43303 4 wl_109
port 118 nsew
rlabel locali s 11496 35403 11496 35403 4 wl_89
port 98 nsew
rlabel locali s 11496 40143 11496 40143 4 wl_101
port 110 nsew
rlabel locali s 11496 34907 11496 34907 4 wl_88
port 97 nsew
rlabel locali s 11496 11997 11496 11997 4 wl_30
port 39 nsew
rlabel locali s 11496 18023 11496 18023 4 wl_45
port 54 nsew
rlabel locali s 11496 18317 11496 18317 4 wl_46
port 55 nsew
rlabel locali s 11496 21973 11496 21973 4 wl_55
port 64 nsew
rlabel locali s 11496 1433 11496 1433 4 wl_3
port 12 nsew
rlabel locali s 11496 12493 11496 12493 4 wl_31
port 40 nsew
rlabel locali s 11496 11703 11496 11703 4 wl_29
port 38 nsew
rlabel locali s 11496 12787 11496 12787 4 wl_32
port 41 nsew
rlabel locali s 11496 8543 11496 8543 4 wl_21
port 30 nsew
rlabel locali s 11496 15653 11496 15653 4 wl_39
port 48 nsew
rlabel locali s 11496 1727 11496 1727 4 wl_4
port 13 nsew
rlabel locali s 11496 14073 11496 14073 4 wl_35
port 44 nsew
rlabel locali s 11496 937 11496 937 4 wl_2
port 11 nsew
rlabel locali s 11496 8047 11496 8047 4 wl_20
port 29 nsew
rlabel locali s 11496 10913 11496 10913 4 wl_27
port 36 nsew
rlabel locali s 11496 643 11496 643 4 wl_1
port 10 nsew
rlabel locali s 11496 9627 11496 9627 4 wl_24
port 33 nsew
rlabel locali s 11496 20687 11496 20687 4 wl_52
port 61 nsew
rlabel locali s 11496 3307 11496 3307 4 wl_8
port 17 nsew
rlabel locali s 11496 5677 11496 5677 4 wl_14
port 23 nsew
rlabel locali s 11496 147 11496 147 4 wl_0
port 9 nsew
rlabel locali s 11496 23057 11496 23057 4 wl_58
port 67 nsew
rlabel locali s 11496 2223 11496 2223 4 wl_5
port 14 nsew
rlabel locali s 11496 15157 11496 15157 4 wl_38
port 47 nsew
rlabel locali s 11496 20393 11496 20393 4 wl_51
port 60 nsew
rlabel locali s 11496 4887 11496 4887 4 wl_12
port 21 nsew
rlabel locali s 11496 8837 11496 8837 4 wl_22
port 31 nsew
rlabel locali s 11496 21183 11496 21183 4 wl_53
port 62 nsew
rlabel locali s 11496 10417 11496 10417 4 wl_26
port 35 nsew
rlabel locali s 11496 19603 11496 19603 4 wl_49
port 58 nsew
rlabel locali s 11496 4097 11496 4097 4 wl_10
port 19 nsew
rlabel locali s 11496 24343 11496 24343 4 wl_61
port 70 nsew
rlabel locali s 11496 23553 11496 23553 4 wl_59
port 68 nsew
rlabel locali s 11496 22267 11496 22267 4 wl_56
port 65 nsew
rlabel locali s 11496 6963 11496 6963 4 wl_17
port 26 nsew
rlabel locali s 11496 9333 11496 9333 4 wl_23
port 32 nsew
rlabel locali s 11496 3803 11496 3803 4 wl_9
port 18 nsew
rlabel locali s 11496 17233 11496 17233 4 wl_43
port 52 nsew
rlabel locali s 11496 4593 11496 4593 4 wl_11
port 20 nsew
rlabel locali s 11496 15947 11496 15947 4 wl_40
port 49 nsew
rlabel locali s 11496 24637 11496 24637 4 wl_62
port 71 nsew
rlabel locali s 11496 25133 11496 25133 4 wl_63
port 72 nsew
rlabel locali s 11496 6173 11496 6173 4 wl_15
port 24 nsew
rlabel locali s 11496 21477 11496 21477 4 wl_54
port 63 nsew
rlabel locali s 11496 23847 11496 23847 4 wl_60
port 69 nsew
rlabel locali s 11496 18813 11496 18813 4 wl_47
port 56 nsew
rlabel locali s 11496 7753 11496 7753 4 wl_19
port 28 nsew
rlabel locali s 11496 19107 11496 19107 4 wl_48
port 57 nsew
rlabel locali s 11496 2517 11496 2517 4 wl_6
port 15 nsew
rlabel locali s 11496 6467 11496 6467 4 wl_16
port 25 nsew
rlabel locali s 11496 16737 11496 16737 4 wl_42
port 51 nsew
rlabel locali s 11496 22763 11496 22763 4 wl_57
port 66 nsew
rlabel locali s 11496 3013 11496 3013 4 wl_7
port 16 nsew
rlabel locali s 11496 10123 11496 10123 4 wl_25
port 34 nsew
rlabel locali s 11496 11207 11496 11207 4 wl_28
port 37 nsew
rlabel locali s 11496 17527 11496 17527 4 wl_44
port 53 nsew
rlabel locali s 11496 13577 11496 13577 4 wl_34
port 43 nsew
rlabel locali s 11496 16443 11496 16443 4 wl_41
port 50 nsew
rlabel locali s 11496 14863 11496 14863 4 wl_37
port 46 nsew
rlabel locali s 11496 13283 11496 13283 4 wl_33
port 42 nsew
rlabel locali s 11496 19897 11496 19897 4 wl_50
port 59 nsew
rlabel locali s 11496 14367 11496 14367 4 wl_36
port 45 nsew
rlabel locali s 11496 7257 11496 7257 4 wl_18
port 27 nsew
rlabel locali s 11496 5383 11496 5383 4 wl_13
port 22 nsew
rlabel metal1 s 432 3979 432 3979 4 addr_5
port 6 nsew
rlabel metal1 s 272 3979 272 3979 4 addr_3
port 4 nsew
rlabel metal1 s 32 3979 32 3979 4 addr_0
port 1 nsew
rlabel metal1 s 192 3979 192 3979 4 addr_2
port 3 nsew
rlabel metal1 s 112 3979 112 3979 4 addr_1
port 2 nsew
rlabel metal1 s 352 3979 352 3979 4 addr_4
port 5 nsew
rlabel metal1 s 512 3979 512 3979 4 addr_6
port 7 nsew
rlabel metal2 s 7596 25280 7596 25280 4 wl_en
port 8 nsew
rlabel metal3 s 7336 50194 7336 50194 4 vdd
port 137 nsew
rlabel metal3 s 7336 47824 7336 47824 4 vdd
port 137 nsew
rlabel metal3 s 7336 48614 7336 48614 4 vdd
port 137 nsew
rlabel metal3 s 7336 47034 7336 47034 4 vdd
port 137 nsew
rlabel metal3 s 7336 45059 7336 45059 4 vdd
port 137 nsew
rlabel metal3 s 7336 44269 7336 44269 4 vdd
port 137 nsew
rlabel metal3 s 7336 49404 7336 49404 4 vdd
port 137 nsew
rlabel metal3 s 7336 49009 7336 49009 4 vdd
port 137 nsew
rlabel metal3 s 7336 47429 7336 47429 4 vdd
port 137 nsew
rlabel metal3 s 7336 44664 7336 44664 4 vdd
port 137 nsew
rlabel metal3 s 7336 46244 7336 46244 4 vdd
port 137 nsew
rlabel metal3 s 7336 45454 7336 45454 4 vdd
port 137 nsew
rlabel metal3 s 7336 48219 7336 48219 4 vdd
port 137 nsew
rlabel metal3 s 7336 49799 7336 49799 4 vdd
port 137 nsew
rlabel metal3 s 7336 46639 7336 46639 4 vdd
port 137 nsew
rlabel metal3 s 7336 45849 7336 45849 4 vdd
port 137 nsew
rlabel metal3 s 6682 45477 6682 45477 4 vdd
port 137 nsew
rlabel metal3 s 7064 49009 7064 49009 4 gnd
port 138 nsew
rlabel metal3 s 7064 45849 7064 45849 4 gnd
port 138 nsew
rlabel metal3 s 6682 46267 6682 46267 4 vdd
port 137 nsew
rlabel metal3 s 6682 48995 6682 48995 4 vdd
port 137 nsew
rlabel metal3 s 6682 46625 6682 46625 4 vdd
port 137 nsew
rlabel metal3 s 6250 47847 6250 47847 4 vdd
port 137 nsew
rlabel metal3 s 6682 49427 6682 49427 4 vdd
port 137 nsew
rlabel metal3 s 6250 49427 6250 49427 4 vdd
port 137 nsew
rlabel metal3 s 7064 47034 7064 47034 4 gnd
port 138 nsew
rlabel metal3 s 6250 47057 6250 47057 4 vdd
port 137 nsew
rlabel metal3 s 6682 47847 6682 47847 4 vdd
port 137 nsew
rlabel metal3 s 7064 48614 7064 48614 4 gnd
port 138 nsew
rlabel metal3 s 6250 49785 6250 49785 4 vdd
port 137 nsew
rlabel metal3 s 7064 48219 7064 48219 4 gnd
port 138 nsew
rlabel metal3 s 7064 49404 7064 49404 4 gnd
port 138 nsew
rlabel metal3 s 6682 48637 6682 48637 4 vdd
port 137 nsew
rlabel metal3 s 7064 50194 7064 50194 4 gnd
port 138 nsew
rlabel metal3 s 6682 50217 6682 50217 4 vdd
port 137 nsew
rlabel metal3 s 7064 46639 7064 46639 4 gnd
port 138 nsew
rlabel metal3 s 6682 48205 6682 48205 4 vdd
port 137 nsew
rlabel metal3 s 6682 47057 6682 47057 4 vdd
port 137 nsew
rlabel metal3 s 6250 50217 6250 50217 4 vdd
port 137 nsew
rlabel metal3 s 7064 45059 7064 45059 4 gnd
port 138 nsew
rlabel metal3 s 6682 44255 6682 44255 4 vdd
port 137 nsew
rlabel metal3 s 6250 46625 6250 46625 4 vdd
port 137 nsew
rlabel metal3 s 7064 49799 7064 49799 4 gnd
port 138 nsew
rlabel metal3 s 6250 48637 6250 48637 4 vdd
port 137 nsew
rlabel metal3 s 6250 46267 6250 46267 4 vdd
port 137 nsew
rlabel metal3 s 7064 44269 7064 44269 4 gnd
port 138 nsew
rlabel metal3 s 6682 44687 6682 44687 4 vdd
port 137 nsew
rlabel metal3 s 6250 44687 6250 44687 4 vdd
port 137 nsew
rlabel metal3 s 6250 48205 6250 48205 4 vdd
port 137 nsew
rlabel metal3 s 7064 45454 7064 45454 4 gnd
port 138 nsew
rlabel metal3 s 6682 45835 6682 45835 4 vdd
port 137 nsew
rlabel metal3 s 6682 49785 6682 49785 4 vdd
port 137 nsew
rlabel metal3 s 6682 47415 6682 47415 4 vdd
port 137 nsew
rlabel metal3 s 6250 47415 6250 47415 4 vdd
port 137 nsew
rlabel metal3 s 7064 44664 7064 44664 4 gnd
port 138 nsew
rlabel metal3 s 6250 45045 6250 45045 4 vdd
port 137 nsew
rlabel metal3 s 6250 44255 6250 44255 4 vdd
port 137 nsew
rlabel metal3 s 6250 45477 6250 45477 4 vdd
port 137 nsew
rlabel metal3 s 7064 46244 7064 46244 4 gnd
port 138 nsew
rlabel metal3 s 6250 48995 6250 48995 4 vdd
port 137 nsew
rlabel metal3 s 7064 47824 7064 47824 4 gnd
port 138 nsew
rlabel metal3 s 6682 45045 6682 45045 4 vdd
port 137 nsew
rlabel metal3 s 7064 47429 7064 47429 4 gnd
port 138 nsew
rlabel metal3 s 6250 45835 6250 45835 4 vdd
port 137 nsew
rlabel metal3 s 7064 41504 7064 41504 4 gnd
port 138 nsew
rlabel metal3 s 6250 38367 6250 38367 4 vdd
port 137 nsew
rlabel metal3 s 6250 39157 6250 39157 4 vdd
port 137 nsew
rlabel metal3 s 6682 42317 6682 42317 4 vdd
port 137 nsew
rlabel metal3 s 7064 42294 7064 42294 4 gnd
port 138 nsew
rlabel metal3 s 6682 37935 6682 37935 4 vdd
port 137 nsew
rlabel metal3 s 7064 43874 7064 43874 4 gnd
port 138 nsew
rlabel metal3 s 7064 39529 7064 39529 4 gnd
port 138 nsew
rlabel metal3 s 6682 39947 6682 39947 4 vdd
port 137 nsew
rlabel metal3 s 6250 43897 6250 43897 4 vdd
port 137 nsew
rlabel metal3 s 6682 40737 6682 40737 4 vdd
port 137 nsew
rlabel metal3 s 6682 43107 6682 43107 4 vdd
port 137 nsew
rlabel metal3 s 6250 37935 6250 37935 4 vdd
port 137 nsew
rlabel metal3 s 7064 40319 7064 40319 4 gnd
port 138 nsew
rlabel metal3 s 6682 41885 6682 41885 4 vdd
port 137 nsew
rlabel metal3 s 7064 38739 7064 38739 4 gnd
port 138 nsew
rlabel metal3 s 7064 40714 7064 40714 4 gnd
port 138 nsew
rlabel metal3 s 6250 41527 6250 41527 4 vdd
port 137 nsew
rlabel metal3 s 6682 38367 6682 38367 4 vdd
port 137 nsew
rlabel metal3 s 7064 42689 7064 42689 4 gnd
port 138 nsew
rlabel metal3 s 7064 38344 7064 38344 4 gnd
port 138 nsew
rlabel metal3 s 6250 40305 6250 40305 4 vdd
port 137 nsew
rlabel metal3 s 6682 43465 6682 43465 4 vdd
port 137 nsew
rlabel metal3 s 6250 40737 6250 40737 4 vdd
port 137 nsew
rlabel metal3 s 6682 41095 6682 41095 4 vdd
port 137 nsew
rlabel metal3 s 7064 41899 7064 41899 4 gnd
port 138 nsew
rlabel metal3 s 6682 40305 6682 40305 4 vdd
port 137 nsew
rlabel metal3 s 7064 37949 7064 37949 4 gnd
port 138 nsew
rlabel metal3 s 6250 39515 6250 39515 4 vdd
port 137 nsew
rlabel metal3 s 6682 41527 6682 41527 4 vdd
port 137 nsew
rlabel metal3 s 6682 39515 6682 39515 4 vdd
port 137 nsew
rlabel metal3 s 6250 41885 6250 41885 4 vdd
port 137 nsew
rlabel metal3 s 6250 39947 6250 39947 4 vdd
port 137 nsew
rlabel metal3 s 6250 42317 6250 42317 4 vdd
port 137 nsew
rlabel metal3 s 6682 42675 6682 42675 4 vdd
port 137 nsew
rlabel metal3 s 6682 43897 6682 43897 4 vdd
port 137 nsew
rlabel metal3 s 7064 43084 7064 43084 4 gnd
port 138 nsew
rlabel metal3 s 7064 39134 7064 39134 4 gnd
port 138 nsew
rlabel metal3 s 6250 41095 6250 41095 4 vdd
port 137 nsew
rlabel metal3 s 7064 43479 7064 43479 4 gnd
port 138 nsew
rlabel metal3 s 7064 39924 7064 39924 4 gnd
port 138 nsew
rlabel metal3 s 7064 41109 7064 41109 4 gnd
port 138 nsew
rlabel metal3 s 6250 38725 6250 38725 4 vdd
port 137 nsew
rlabel metal3 s 6682 38725 6682 38725 4 vdd
port 137 nsew
rlabel metal3 s 6682 39157 6682 39157 4 vdd
port 137 nsew
rlabel metal3 s 6250 43107 6250 43107 4 vdd
port 137 nsew
rlabel metal3 s 6250 42675 6250 42675 4 vdd
port 137 nsew
rlabel metal3 s 6250 43465 6250 43465 4 vdd
port 137 nsew
rlabel metal3 s 7336 39529 7336 39529 4 vdd
port 137 nsew
rlabel metal3 s 7336 43874 7336 43874 4 vdd
port 137 nsew
rlabel metal3 s 7336 39134 7336 39134 4 vdd
port 137 nsew
rlabel metal3 s 7336 38739 7336 38739 4 vdd
port 137 nsew
rlabel metal3 s 7336 40319 7336 40319 4 vdd
port 137 nsew
rlabel metal3 s 7336 37949 7336 37949 4 vdd
port 137 nsew
rlabel metal3 s 7336 43479 7336 43479 4 vdd
port 137 nsew
rlabel metal3 s 7336 41899 7336 41899 4 vdd
port 137 nsew
rlabel metal3 s 7336 38344 7336 38344 4 vdd
port 137 nsew
rlabel metal3 s 7336 40714 7336 40714 4 vdd
port 137 nsew
rlabel metal3 s 7336 42689 7336 42689 4 vdd
port 137 nsew
rlabel metal3 s 7336 41109 7336 41109 4 vdd
port 137 nsew
rlabel metal3 s 7336 41504 7336 41504 4 vdd
port 137 nsew
rlabel metal3 s 7336 42294 7336 42294 4 vdd
port 137 nsew
rlabel metal3 s 7336 43084 7336 43084 4 vdd
port 137 nsew
rlabel metal3 s 7336 39924 7336 39924 4 vdd
port 137 nsew
rlabel metal3 s 5825 49843 5825 49843 4 gnd
port 138 nsew
rlabel metal3 s 5825 47057 5825 47057 4 gnd
port 138 nsew
rlabel metal3 s 5825 47473 5825 47473 4 gnd
port 138 nsew
rlabel metal3 s 5825 41943 5825 41943 4 gnd
port 138 nsew
rlabel metal3 s 5825 39573 5825 39573 4 gnd
port 138 nsew
rlabel metal3 s 5825 46267 5825 46267 4 gnd
port 138 nsew
rlabel metal3 s 5825 39157 5825 39157 4 gnd
port 138 nsew
rlabel metal3 s 5825 49427 5825 49427 4 gnd
port 138 nsew
rlabel metal3 s 5825 44687 5825 44687 4 gnd
port 138 nsew
rlabel metal3 s 5825 45893 5825 45893 4 gnd
port 138 nsew
rlabel metal3 s 5825 45477 5825 45477 4 gnd
port 138 nsew
rlabel metal3 s 5825 42317 5825 42317 4 gnd
port 138 nsew
rlabel metal3 s 5825 43897 5825 43897 4 gnd
port 138 nsew
rlabel metal3 s 5825 42733 5825 42733 4 gnd
port 138 nsew
rlabel metal3 s 5825 41153 5825 41153 4 gnd
port 138 nsew
rlabel metal3 s 5825 47847 5825 47847 4 gnd
port 138 nsew
rlabel metal3 s 5825 38783 5825 38783 4 gnd
port 138 nsew
rlabel metal3 s 5825 41527 5825 41527 4 gnd
port 138 nsew
rlabel metal3 s 5825 43523 5825 43523 4 gnd
port 138 nsew
rlabel metal3 s 5825 50217 5825 50217 4 gnd
port 138 nsew
rlabel metal3 s 5825 37993 5825 37993 4 gnd
port 138 nsew
rlabel metal3 s 5825 46683 5825 46683 4 gnd
port 138 nsew
rlabel metal3 s 5825 48637 5825 48637 4 gnd
port 138 nsew
rlabel metal3 s 5825 48263 5825 48263 4 gnd
port 138 nsew
rlabel metal3 s 5825 39947 5825 39947 4 gnd
port 138 nsew
rlabel metal3 s 5825 49053 5825 49053 4 gnd
port 138 nsew
rlabel metal3 s 5825 38367 5825 38367 4 gnd
port 138 nsew
rlabel metal3 s 5825 45103 5825 45103 4 gnd
port 138 nsew
rlabel metal3 s 5825 43107 5825 43107 4 gnd
port 138 nsew
rlabel metal3 s 5825 40737 5825 40737 4 gnd
port 138 nsew
rlabel metal3 s 5825 40363 5825 40363 4 gnd
port 138 nsew
rlabel metal3 s 5825 44313 5825 44313 4 gnd
port 138 nsew
rlabel metal3 s 5825 31673 5825 31673 4 gnd
port 138 nsew
rlabel metal3 s 5825 26517 5825 26517 4 gnd
port 138 nsew
rlabel metal3 s 5825 37203 5825 37203 4 gnd
port 138 nsew
rlabel metal3 s 5825 28513 5825 28513 4 gnd
port 138 nsew
rlabel metal3 s 5825 34833 5825 34833 4 gnd
port 138 nsew
rlabel metal3 s 5825 30093 5825 30093 4 gnd
port 138 nsew
rlabel metal3 s 5825 32837 5825 32837 4 gnd
port 138 nsew
rlabel metal3 s 5825 35997 5825 35997 4 gnd
port 138 nsew
rlabel metal3 s 5825 29303 5825 29303 4 gnd
port 138 nsew
rlabel metal3 s 5825 33627 5825 33627 4 gnd
port 138 nsew
rlabel metal3 s 5825 28887 5825 28887 4 gnd
port 138 nsew
rlabel metal3 s 5825 26933 5825 26933 4 gnd
port 138 nsew
rlabel metal3 s 5825 37577 5825 37577 4 gnd
port 138 nsew
rlabel metal3 s 5825 31257 5825 31257 4 gnd
port 138 nsew
rlabel metal3 s 5825 27307 5825 27307 4 gnd
port 138 nsew
rlabel metal3 s 5825 34043 5825 34043 4 gnd
port 138 nsew
rlabel metal3 s 5825 29677 5825 29677 4 gnd
port 138 nsew
rlabel metal3 s 5825 33253 5825 33253 4 gnd
port 138 nsew
rlabel metal3 s 5825 30467 5825 30467 4 gnd
port 138 nsew
rlabel metal3 s 5825 25353 5825 25353 4 gnd
port 138 nsew
rlabel metal3 s 5825 35623 5825 35623 4 gnd
port 138 nsew
rlabel metal3 s 5825 28097 5825 28097 4 gnd
port 138 nsew
rlabel metal3 s 5825 30883 5825 30883 4 gnd
port 138 nsew
rlabel metal3 s 5825 32047 5825 32047 4 gnd
port 138 nsew
rlabel metal3 s 5825 34417 5825 34417 4 gnd
port 138 nsew
rlabel metal3 s 5825 36787 5825 36787 4 gnd
port 138 nsew
rlabel metal3 s 5825 32463 5825 32463 4 gnd
port 138 nsew
rlabel metal3 s 5825 25727 5825 25727 4 gnd
port 138 nsew
rlabel metal3 s 5825 36413 5825 36413 4 gnd
port 138 nsew
rlabel metal3 s 5825 26143 5825 26143 4 gnd
port 138 nsew
rlabel metal3 s 5825 27723 5825 27723 4 gnd
port 138 nsew
rlabel metal3 s 5825 35207 5825 35207 4 gnd
port 138 nsew
rlabel metal3 s 7336 36764 7336 36764 4 vdd
port 137 nsew
rlabel metal3 s 7336 32419 7336 32419 4 vdd
port 137 nsew
rlabel metal3 s 7336 35579 7336 35579 4 vdd
port 137 nsew
rlabel metal3 s 7336 37554 7336 37554 4 vdd
port 137 nsew
rlabel metal3 s 7336 35184 7336 35184 4 vdd
port 137 nsew
rlabel metal3 s 7336 33209 7336 33209 4 vdd
port 137 nsew
rlabel metal3 s 7336 31629 7336 31629 4 vdd
port 137 nsew
rlabel metal3 s 7336 32024 7336 32024 4 vdd
port 137 nsew
rlabel metal3 s 7336 37159 7336 37159 4 vdd
port 137 nsew
rlabel metal3 s 7336 34394 7336 34394 4 vdd
port 137 nsew
rlabel metal3 s 7336 33999 7336 33999 4 vdd
port 137 nsew
rlabel metal3 s 7336 36369 7336 36369 4 vdd
port 137 nsew
rlabel metal3 s 7336 33604 7336 33604 4 vdd
port 137 nsew
rlabel metal3 s 7336 32814 7336 32814 4 vdd
port 137 nsew
rlabel metal3 s 7336 34789 7336 34789 4 vdd
port 137 nsew
rlabel metal3 s 7336 35974 7336 35974 4 vdd
port 137 nsew
rlabel metal3 s 7064 35974 7064 35974 4 gnd
port 138 nsew
rlabel metal3 s 7064 32419 7064 32419 4 gnd
port 138 nsew
rlabel metal3 s 7064 37159 7064 37159 4 gnd
port 138 nsew
rlabel metal3 s 6250 36355 6250 36355 4 vdd
port 137 nsew
rlabel metal3 s 7064 34789 7064 34789 4 gnd
port 138 nsew
rlabel metal3 s 6250 35565 6250 35565 4 vdd
port 137 nsew
rlabel metal3 s 6682 37145 6682 37145 4 vdd
port 137 nsew
rlabel metal3 s 6682 32837 6682 32837 4 vdd
port 137 nsew
rlabel metal3 s 7064 36764 7064 36764 4 gnd
port 138 nsew
rlabel metal3 s 6682 35997 6682 35997 4 vdd
port 137 nsew
rlabel metal3 s 6682 32047 6682 32047 4 vdd
port 137 nsew
rlabel metal3 s 7064 35184 7064 35184 4 gnd
port 138 nsew
rlabel metal3 s 6250 33985 6250 33985 4 vdd
port 137 nsew
rlabel metal3 s 7064 32024 7064 32024 4 gnd
port 138 nsew
rlabel metal3 s 7064 36369 7064 36369 4 gnd
port 138 nsew
rlabel metal3 s 6250 34417 6250 34417 4 vdd
port 137 nsew
rlabel metal3 s 6250 31615 6250 31615 4 vdd
port 137 nsew
rlabel metal3 s 6682 37577 6682 37577 4 vdd
port 137 nsew
rlabel metal3 s 7064 33604 7064 33604 4 gnd
port 138 nsew
rlabel metal3 s 7064 33999 7064 33999 4 gnd
port 138 nsew
rlabel metal3 s 7064 32814 7064 32814 4 gnd
port 138 nsew
rlabel metal3 s 6250 37577 6250 37577 4 vdd
port 137 nsew
rlabel metal3 s 6250 36787 6250 36787 4 vdd
port 137 nsew
rlabel metal3 s 6682 32405 6682 32405 4 vdd
port 137 nsew
rlabel metal3 s 6682 33985 6682 33985 4 vdd
port 137 nsew
rlabel metal3 s 6682 36355 6682 36355 4 vdd
port 137 nsew
rlabel metal3 s 6682 33195 6682 33195 4 vdd
port 137 nsew
rlabel metal3 s 6250 32047 6250 32047 4 vdd
port 137 nsew
rlabel metal3 s 6682 34775 6682 34775 4 vdd
port 137 nsew
rlabel metal3 s 6682 35565 6682 35565 4 vdd
port 137 nsew
rlabel metal3 s 7064 33209 7064 33209 4 gnd
port 138 nsew
rlabel metal3 s 6250 35997 6250 35997 4 vdd
port 137 nsew
rlabel metal3 s 6250 32405 6250 32405 4 vdd
port 137 nsew
rlabel metal3 s 6250 37145 6250 37145 4 vdd
port 137 nsew
rlabel metal3 s 6250 34775 6250 34775 4 vdd
port 137 nsew
rlabel metal3 s 6250 32837 6250 32837 4 vdd
port 137 nsew
rlabel metal3 s 6250 35207 6250 35207 4 vdd
port 137 nsew
rlabel metal3 s 6682 34417 6682 34417 4 vdd
port 137 nsew
rlabel metal3 s 6682 35207 6682 35207 4 vdd
port 137 nsew
rlabel metal3 s 7064 37554 7064 37554 4 gnd
port 138 nsew
rlabel metal3 s 6250 33195 6250 33195 4 vdd
port 137 nsew
rlabel metal3 s 6682 33627 6682 33627 4 vdd
port 137 nsew
rlabel metal3 s 7064 35579 7064 35579 4 gnd
port 138 nsew
rlabel metal3 s 6250 33627 6250 33627 4 vdd
port 137 nsew
rlabel metal3 s 6682 36787 6682 36787 4 vdd
port 137 nsew
rlabel metal3 s 6682 31615 6682 31615 4 vdd
port 137 nsew
rlabel metal3 s 7064 34394 7064 34394 4 gnd
port 138 nsew
rlabel metal3 s 7064 31629 7064 31629 4 gnd
port 138 nsew
rlabel metal3 s 6250 27665 6250 27665 4 vdd
port 137 nsew
rlabel metal3 s 6250 28097 6250 28097 4 vdd
port 137 nsew
rlabel metal3 s 7064 30444 7064 30444 4 gnd
port 138 nsew
rlabel metal3 s 6682 26517 6682 26517 4 vdd
port 137 nsew
rlabel metal3 s 7064 31234 7064 31234 4 gnd
port 138 nsew
rlabel metal3 s 7064 30839 7064 30839 4 gnd
port 138 nsew
rlabel metal3 s 6682 30467 6682 30467 4 vdd
port 137 nsew
rlabel metal3 s 7064 28074 7064 28074 4 gnd
port 138 nsew
rlabel metal3 s 6250 26875 6250 26875 4 vdd
port 137 nsew
rlabel metal3 s 6682 30035 6682 30035 4 vdd
port 137 nsew
rlabel metal3 s 6250 27307 6250 27307 4 vdd
port 137 nsew
rlabel metal3 s 6250 26517 6250 26517 4 vdd
port 137 nsew
rlabel metal3 s 6250 28887 6250 28887 4 vdd
port 137 nsew
rlabel metal3 s 7064 27284 7064 27284 4 gnd
port 138 nsew
rlabel metal3 s 6250 29245 6250 29245 4 vdd
port 137 nsew
rlabel metal3 s 6682 29245 6682 29245 4 vdd
port 137 nsew
rlabel metal3 s 7064 27679 7064 27679 4 gnd
port 138 nsew
rlabel metal3 s 6682 28455 6682 28455 4 vdd
port 137 nsew
rlabel metal3 s 7064 29654 7064 29654 4 gnd
port 138 nsew
rlabel metal3 s 7064 26889 7064 26889 4 gnd
port 138 nsew
rlabel metal3 s 7064 30049 7064 30049 4 gnd
port 138 nsew
rlabel metal3 s 7064 26494 7064 26494 4 gnd
port 138 nsew
rlabel metal3 s 6682 29677 6682 29677 4 vdd
port 137 nsew
rlabel metal3 s 6250 29677 6250 29677 4 vdd
port 137 nsew
rlabel metal3 s 7064 28469 7064 28469 4 gnd
port 138 nsew
rlabel metal3 s 6682 25727 6682 25727 4 vdd
port 137 nsew
rlabel metal3 s 6250 30035 6250 30035 4 vdd
port 137 nsew
rlabel metal3 s 6682 30825 6682 30825 4 vdd
port 137 nsew
rlabel metal3 s 7064 25704 7064 25704 4 gnd
port 138 nsew
rlabel metal3 s 6682 31257 6682 31257 4 vdd
port 137 nsew
rlabel metal3 s 6682 28887 6682 28887 4 vdd
port 137 nsew
rlabel metal3 s 6682 27307 6682 27307 4 vdd
port 137 nsew
rlabel metal3 s 6250 31257 6250 31257 4 vdd
port 137 nsew
rlabel metal3 s 6250 26085 6250 26085 4 vdd
port 137 nsew
rlabel metal3 s 6682 26875 6682 26875 4 vdd
port 137 nsew
rlabel metal3 s 6682 28097 6682 28097 4 vdd
port 137 nsew
rlabel metal3 s 6250 25727 6250 25727 4 vdd
port 137 nsew
rlabel metal3 s 7064 29259 7064 29259 4 gnd
port 138 nsew
rlabel metal3 s 6250 30467 6250 30467 4 vdd
port 137 nsew
rlabel metal3 s 6682 27665 6682 27665 4 vdd
port 137 nsew
rlabel metal3 s 6250 30825 6250 30825 4 vdd
port 137 nsew
rlabel metal3 s 7336 30049 7336 30049 4 vdd
port 137 nsew
rlabel metal3 s 7336 30839 7336 30839 4 vdd
port 137 nsew
rlabel metal3 s 7336 28074 7336 28074 4 vdd
port 137 nsew
rlabel metal3 s 7336 27679 7336 27679 4 vdd
port 137 nsew
rlabel metal3 s 7336 27284 7336 27284 4 vdd
port 137 nsew
rlabel metal3 s 7336 29259 7336 29259 4 vdd
port 137 nsew
rlabel metal3 s 7336 31234 7336 31234 4 vdd
port 137 nsew
rlabel metal3 s 7336 26494 7336 26494 4 vdd
port 137 nsew
rlabel metal3 s 7336 26099 7336 26099 4 vdd
port 137 nsew
rlabel metal3 s 7336 28864 7336 28864 4 vdd
port 137 nsew
rlabel metal3 s 7336 30444 7336 30444 4 vdd
port 137 nsew
rlabel metal3 s 7336 25704 7336 25704 4 vdd
port 137 nsew
rlabel metal3 s 7336 29654 7336 29654 4 vdd
port 137 nsew
rlabel metal3 s 7336 28469 7336 28469 4 vdd
port 137 nsew
rlabel metal3 s 7336 26889 7336 26889 4 vdd
port 137 nsew
rlabel metal3 s 6682 26085 6682 26085 4 vdd
port 137 nsew
rlabel metal3 s 7064 26099 7064 26099 4 gnd
port 138 nsew
rlabel metal3 s 6250 28455 6250 28455 4 vdd
port 137 nsew
rlabel metal3 s 7064 28864 7064 28864 4 gnd
port 138 nsew
rlabel metal3 s 1204 5164 1204 5164 4 gnd
port 138 nsew
rlabel metal3 s 9250 25280 9250 25280 4 gnd
port 138 nsew
rlabel metal3 s 10774 25280 10774 25280 4 vdd
port 137 nsew
rlabel metal3 s 7336 25309 7336 25309 4 vdd
port 137 nsew
rlabel metal3 s 7336 21754 7336 21754 4 vdd
port 137 nsew
rlabel metal3 s 7336 19779 7336 19779 4 vdd
port 137 nsew
rlabel metal3 s 7336 22149 7336 22149 4 vdd
port 137 nsew
rlabel metal3 s 7336 22544 7336 22544 4 vdd
port 137 nsew
rlabel metal3 s 7782 25265 7782 25265 4 gnd
port 138 nsew
rlabel metal3 s 7336 24519 7336 24519 4 vdd
port 137 nsew
rlabel metal3 s 7336 20569 7336 20569 4 vdd
port 137 nsew
rlabel metal3 s 7336 24124 7336 24124 4 vdd
port 137 nsew
rlabel metal3 s 7336 20174 7336 20174 4 vdd
port 137 nsew
rlabel metal3 s 7336 22939 7336 22939 4 vdd
port 137 nsew
rlabel metal3 s 7336 21359 7336 21359 4 vdd
port 137 nsew
rlabel metal3 s 7336 20964 7336 20964 4 vdd
port 137 nsew
rlabel metal3 s 7336 24914 7336 24914 4 vdd
port 137 nsew
rlabel metal3 s 7336 23729 7336 23729 4 vdd
port 137 nsew
rlabel metal3 s 8207 25264 8207 25264 4 vdd
port 137 nsew
rlabel metal3 s 7336 19384 7336 19384 4 vdd
port 137 nsew
rlabel metal3 s 7336 23334 7336 23334 4 vdd
port 137 nsew
rlabel metal3 s 6682 22567 6682 22567 4 vdd
port 137 nsew
rlabel metal3 s 6250 22135 6250 22135 4 vdd
port 137 nsew
rlabel metal3 s 6250 22567 6250 22567 4 vdd
port 137 nsew
rlabel metal3 s 7064 23729 7064 23729 4 gnd
port 138 nsew
rlabel metal3 s 6250 20555 6250 20555 4 vdd
port 137 nsew
rlabel metal3 s 7064 24124 7064 24124 4 gnd
port 138 nsew
rlabel metal3 s 6682 24505 6682 24505 4 vdd
port 137 nsew
rlabel metal3 s 7064 22149 7064 22149 4 gnd
port 138 nsew
rlabel metal3 s 6682 22925 6682 22925 4 vdd
port 137 nsew
rlabel metal3 s 7064 19779 7064 19779 4 gnd
port 138 nsew
rlabel metal3 s 7064 20569 7064 20569 4 gnd
port 138 nsew
rlabel metal3 s 7064 24914 7064 24914 4 gnd
port 138 nsew
rlabel metal3 s 6250 21345 6250 21345 4 vdd
port 137 nsew
rlabel metal3 s 7064 21754 7064 21754 4 gnd
port 138 nsew
rlabel metal3 s 6682 19407 6682 19407 4 vdd
port 137 nsew
rlabel metal3 s 6250 23715 6250 23715 4 vdd
port 137 nsew
rlabel metal3 s 6250 21777 6250 21777 4 vdd
port 137 nsew
rlabel metal3 s 7064 19384 7064 19384 4 gnd
port 138 nsew
rlabel metal3 s 6250 25295 6250 25295 4 vdd
port 137 nsew
rlabel metal3 s 7064 24519 7064 24519 4 gnd
port 138 nsew
rlabel metal3 s 7064 20174 7064 20174 4 gnd
port 138 nsew
rlabel metal3 s 7064 23334 7064 23334 4 gnd
port 138 nsew
rlabel metal3 s 6682 23715 6682 23715 4 vdd
port 137 nsew
rlabel metal3 s 7064 25309 7064 25309 4 gnd
port 138 nsew
rlabel metal3 s 7064 22544 7064 22544 4 gnd
port 138 nsew
rlabel metal3 s 6682 23357 6682 23357 4 vdd
port 137 nsew
rlabel metal3 s 6682 20987 6682 20987 4 vdd
port 137 nsew
rlabel metal3 s 6682 24937 6682 24937 4 vdd
port 137 nsew
rlabel metal3 s 6250 20987 6250 20987 4 vdd
port 137 nsew
rlabel metal3 s 6250 19765 6250 19765 4 vdd
port 137 nsew
rlabel metal3 s 7064 22939 7064 22939 4 gnd
port 138 nsew
rlabel metal3 s 6682 21777 6682 21777 4 vdd
port 137 nsew
rlabel metal3 s 6250 24505 6250 24505 4 vdd
port 137 nsew
rlabel metal3 s 6250 23357 6250 23357 4 vdd
port 137 nsew
rlabel metal3 s 7064 20964 7064 20964 4 gnd
port 138 nsew
rlabel metal3 s 6250 20197 6250 20197 4 vdd
port 137 nsew
rlabel metal3 s 6682 21345 6682 21345 4 vdd
port 137 nsew
rlabel metal3 s 6250 24147 6250 24147 4 vdd
port 137 nsew
rlabel metal3 s 6682 22135 6682 22135 4 vdd
port 137 nsew
rlabel metal3 s 6682 19765 6682 19765 4 vdd
port 137 nsew
rlabel metal3 s 6682 25295 6682 25295 4 vdd
port 137 nsew
rlabel metal3 s 6682 20197 6682 20197 4 vdd
port 137 nsew
rlabel metal3 s 6250 22925 6250 22925 4 vdd
port 137 nsew
rlabel metal3 s 6682 20555 6682 20555 4 vdd
port 137 nsew
rlabel metal3 s 7064 21359 7064 21359 4 gnd
port 138 nsew
rlabel metal3 s 6682 24147 6682 24147 4 vdd
port 137 nsew
rlabel metal3 s 6250 24937 6250 24937 4 vdd
port 137 nsew
rlabel metal3 s 6250 19407 6250 19407 4 vdd
port 137 nsew
rlabel metal3 s 6682 16605 6682 16605 4 vdd
port 137 nsew
rlabel metal3 s 7064 13064 7064 13064 4 gnd
port 138 nsew
rlabel metal3 s 6250 15815 6250 15815 4 vdd
port 137 nsew
rlabel metal3 s 7064 14249 7064 14249 4 gnd
port 138 nsew
rlabel metal3 s 6682 13445 6682 13445 4 vdd
port 137 nsew
rlabel metal3 s 6682 18185 6682 18185 4 vdd
port 137 nsew
rlabel metal3 s 7064 18989 7064 18989 4 gnd
port 138 nsew
rlabel metal3 s 6682 14667 6682 14667 4 vdd
port 137 nsew
rlabel metal3 s 7064 13854 7064 13854 4 gnd
port 138 nsew
rlabel metal3 s 7064 17409 7064 17409 4 gnd
port 138 nsew
rlabel metal3 s 7064 17014 7064 17014 4 gnd
port 138 nsew
rlabel metal3 s 6250 17037 6250 17037 4 vdd
port 137 nsew
rlabel metal3 s 6250 18185 6250 18185 4 vdd
port 137 nsew
rlabel metal3 s 6250 14667 6250 14667 4 vdd
port 137 nsew
rlabel metal3 s 7064 14644 7064 14644 4 gnd
port 138 nsew
rlabel metal3 s 7064 17804 7064 17804 4 gnd
port 138 nsew
rlabel metal3 s 7064 16224 7064 16224 4 gnd
port 138 nsew
rlabel metal3 s 6682 18617 6682 18617 4 vdd
port 137 nsew
rlabel metal3 s 7064 15434 7064 15434 4 gnd
port 138 nsew
rlabel metal3 s 6682 15025 6682 15025 4 vdd
port 137 nsew
rlabel metal3 s 7064 18199 7064 18199 4 gnd
port 138 nsew
rlabel metal3 s 6682 17827 6682 17827 4 vdd
port 137 nsew
rlabel metal3 s 6682 17395 6682 17395 4 vdd
port 137 nsew
rlabel metal3 s 6682 14235 6682 14235 4 vdd
port 137 nsew
rlabel metal3 s 6250 13087 6250 13087 4 vdd
port 137 nsew
rlabel metal3 s 6682 18975 6682 18975 4 vdd
port 137 nsew
rlabel metal3 s 6250 16605 6250 16605 4 vdd
port 137 nsew
rlabel metal3 s 7064 16619 7064 16619 4 gnd
port 138 nsew
rlabel metal3 s 6682 15815 6682 15815 4 vdd
port 137 nsew
rlabel metal3 s 6250 13877 6250 13877 4 vdd
port 137 nsew
rlabel metal3 s 6250 13445 6250 13445 4 vdd
port 137 nsew
rlabel metal3 s 6682 13877 6682 13877 4 vdd
port 137 nsew
rlabel metal3 s 6682 17037 6682 17037 4 vdd
port 137 nsew
rlabel metal3 s 7064 15829 7064 15829 4 gnd
port 138 nsew
rlabel metal3 s 6682 16247 6682 16247 4 vdd
port 137 nsew
rlabel metal3 s 6250 18617 6250 18617 4 vdd
port 137 nsew
rlabel metal3 s 6250 16247 6250 16247 4 vdd
port 137 nsew
rlabel metal3 s 6250 17827 6250 17827 4 vdd
port 137 nsew
rlabel metal3 s 6682 15457 6682 15457 4 vdd
port 137 nsew
rlabel metal3 s 6250 17395 6250 17395 4 vdd
port 137 nsew
rlabel metal3 s 6250 18975 6250 18975 4 vdd
port 137 nsew
rlabel metal3 s 7064 13459 7064 13459 4 gnd
port 138 nsew
rlabel metal3 s 6250 14235 6250 14235 4 vdd
port 137 nsew
rlabel metal3 s 7064 15039 7064 15039 4 gnd
port 138 nsew
rlabel metal3 s 7064 18594 7064 18594 4 gnd
port 138 nsew
rlabel metal3 s 6250 15457 6250 15457 4 vdd
port 137 nsew
rlabel metal3 s 6682 13087 6682 13087 4 vdd
port 137 nsew
rlabel metal3 s 6250 15025 6250 15025 4 vdd
port 137 nsew
rlabel metal3 s 7336 13064 7336 13064 4 vdd
port 137 nsew
rlabel metal3 s 7336 18989 7336 18989 4 vdd
port 137 nsew
rlabel metal3 s 7336 17014 7336 17014 4 vdd
port 137 nsew
rlabel metal3 s 7336 13459 7336 13459 4 vdd
port 137 nsew
rlabel metal3 s 7336 15039 7336 15039 4 vdd
port 137 nsew
rlabel metal3 s 7336 14644 7336 14644 4 vdd
port 137 nsew
rlabel metal3 s 7336 17804 7336 17804 4 vdd
port 137 nsew
rlabel metal3 s 7336 13854 7336 13854 4 vdd
port 137 nsew
rlabel metal3 s 7336 15434 7336 15434 4 vdd
port 137 nsew
rlabel metal3 s 7336 17409 7336 17409 4 vdd
port 137 nsew
rlabel metal3 s 7336 18594 7336 18594 4 vdd
port 137 nsew
rlabel metal3 s 7336 18199 7336 18199 4 vdd
port 137 nsew
rlabel metal3 s 7336 14249 7336 14249 4 vdd
port 137 nsew
rlabel metal3 s 7336 16224 7336 16224 4 vdd
port 137 nsew
rlabel metal3 s 7336 15829 7336 15829 4 vdd
port 137 nsew
rlabel metal3 s 7336 16619 7336 16619 4 vdd
port 137 nsew
rlabel metal3 s 5825 22567 5825 22567 4 gnd
port 138 nsew
rlabel metal3 s 5825 20613 5825 20613 4 gnd
port 138 nsew
rlabel metal3 s 5825 14667 5825 14667 4 gnd
port 138 nsew
rlabel metal3 s 5825 19407 5825 19407 4 gnd
port 138 nsew
rlabel metal3 s 5825 15083 5825 15083 4 gnd
port 138 nsew
rlabel metal3 s 5825 22983 5825 22983 4 gnd
port 138 nsew
rlabel metal3 s 5825 17453 5825 17453 4 gnd
port 138 nsew
rlabel metal3 s 5825 15873 5825 15873 4 gnd
port 138 nsew
rlabel metal3 s 5825 24147 5825 24147 4 gnd
port 138 nsew
rlabel metal3 s 5825 13087 5825 13087 4 gnd
port 138 nsew
rlabel metal3 s 5825 18243 5825 18243 4 gnd
port 138 nsew
rlabel metal3 s 5825 18617 5825 18617 4 gnd
port 138 nsew
rlabel metal3 s 5825 23357 5825 23357 4 gnd
port 138 nsew
rlabel metal3 s 5825 19033 5825 19033 4 gnd
port 138 nsew
rlabel metal3 s 5825 22193 5825 22193 4 gnd
port 138 nsew
rlabel metal3 s 5825 14293 5825 14293 4 gnd
port 138 nsew
rlabel metal3 s 5825 24563 5825 24563 4 gnd
port 138 nsew
rlabel metal3 s 5825 24937 5825 24937 4 gnd
port 138 nsew
rlabel metal3 s 5825 17037 5825 17037 4 gnd
port 138 nsew
rlabel metal3 s 5825 13503 5825 13503 4 gnd
port 138 nsew
rlabel metal3 s 5825 19823 5825 19823 4 gnd
port 138 nsew
rlabel metal3 s 5825 21777 5825 21777 4 gnd
port 138 nsew
rlabel metal3 s 5825 20987 5825 20987 4 gnd
port 138 nsew
rlabel metal3 s 5825 16247 5825 16247 4 gnd
port 138 nsew
rlabel metal3 s 5825 13877 5825 13877 4 gnd
port 138 nsew
rlabel metal3 s 5825 21403 5825 21403 4 gnd
port 138 nsew
rlabel metal3 s 5825 20197 5825 20197 4 gnd
port 138 nsew
rlabel metal3 s 5825 23773 5825 23773 4 gnd
port 138 nsew
rlabel metal3 s 5825 15457 5825 15457 4 gnd
port 138 nsew
rlabel metal3 s 5825 17827 5825 17827 4 gnd
port 138 nsew
rlabel metal3 s 5825 16663 5825 16663 4 gnd
port 138 nsew
rlabel metal3 s 5825 11133 5825 11133 4 gnd
port 138 nsew
rlabel metal3 s 5825 4023 5825 4023 4 gnd
port 138 nsew
rlabel metal3 s 4046 7534 4046 7534 4 vdd
port 137 nsew
rlabel metal3 s 5825 5977 5825 5977 4 gnd
port 138 nsew
rlabel metal3 s 5825 8763 5825 8763 4 gnd
port 138 nsew
rlabel metal3 s 5825 2027 5825 2027 4 gnd
port 138 nsew
rlabel metal3 s 5825 9553 5825 9553 4 gnd
port 138 nsew
rlabel metal3 s 5825 7557 5825 7557 4 gnd
port 138 nsew
rlabel metal3 s 4046 5954 4046 5954 4 vdd
port 137 nsew
rlabel metal3 s 5825 4813 5825 4813 4 gnd
port 138 nsew
rlabel metal3 s 5825 2817 5825 2817 4 gnd
port 138 nsew
rlabel metal3 s 4046 6744 4046 6744 4 vdd
port 137 nsew
rlabel metal3 s 3774 3584 3774 3584 4 gnd
port 138 nsew
rlabel metal3 s 3774 5954 3774 5954 4 gnd
port 138 nsew
rlabel metal3 s 2970 2801 2970 2801 4 gnd
port 138 nsew
rlabel metal3 s 3395 431 3395 431 4 vdd
port 137 nsew
rlabel metal3 s 1800 424 1800 424 4 gnd
port 138 nsew
rlabel metal3 s 2960 7557 2960 7557 4 vdd
port 137 nsew
rlabel metal3 s 3392 5187 3392 5187 4 vdd
port 137 nsew
rlabel metal3 s 1476 5164 1476 5164 4 vdd
port 137 nsew
rlabel metal3 s 2970 1221 2970 1221 4 gnd
port 138 nsew
rlabel metal3 s 3395 1221 3395 1221 4 vdd
port 137 nsew
rlabel metal3 s 2072 424 2072 424 4 vdd
port 137 nsew
rlabel metal3 s 2535 7557 2535 7557 4 gnd
port 138 nsew
rlabel metal3 s 2970 3591 2970 3591 4 gnd
port 138 nsew
rlabel metal3 s 3395 3591 3395 3591 4 vdd
port 137 nsew
rlabel metal3 s 3395 2801 3395 2801 4 vdd
port 137 nsew
rlabel metal3 s 2960 6767 2960 6767 4 vdd
port 137 nsew
rlabel metal3 s 2072 2794 2072 2794 4 vdd
port 137 nsew
rlabel metal3 s 3392 7557 3392 7557 4 vdd
port 137 nsew
rlabel metal3 s 2535 5187 2535 5187 4 gnd
port 138 nsew
rlabel metal3 s 2960 5977 2960 5977 4 vdd
port 137 nsew
rlabel metal3 s 3392 6767 3392 6767 4 vdd
port 137 nsew
rlabel metal3 s 2970 431 2970 431 4 gnd
port 138 nsew
rlabel metal3 s 2535 6767 2535 6767 4 gnd
port 138 nsew
rlabel metal3 s 3392 5977 3392 5977 4 vdd
port 137 nsew
rlabel metal3 s 2960 5187 2960 5187 4 vdd
port 137 nsew
rlabel metal3 s 2535 5977 2535 5977 4 gnd
port 138 nsew
rlabel metal3 s 1800 2794 1800 2794 4 gnd
port 138 nsew
rlabel metal3 s 5825 1653 5825 1653 4 gnd
port 138 nsew
rlabel metal3 s 3774 6744 3774 6744 4 gnd
port 138 nsew
rlabel metal3 s 5825 9927 5825 9927 4 gnd
port 138 nsew
rlabel metal3 s 5825 4397 5825 4397 4 gnd
port 138 nsew
rlabel metal3 s 3774 5164 3774 5164 4 gnd
port 138 nsew
rlabel metal3 s 4046 424 4046 424 4 vdd
port 137 nsew
rlabel metal3 s 5825 11923 5825 11923 4 gnd
port 138 nsew
rlabel metal3 s 5825 8347 5825 8347 4 gnd
port 138 nsew
rlabel metal3 s 5825 1237 5825 1237 4 gnd
port 138 nsew
rlabel metal3 s 5825 10717 5825 10717 4 gnd
port 138 nsew
rlabel metal3 s 4046 2794 4046 2794 4 vdd
port 137 nsew
rlabel metal3 s 4046 5164 4046 5164 4 vdd
port 137 nsew
rlabel metal3 s 5825 3233 5825 3233 4 gnd
port 138 nsew
rlabel metal3 s 5825 5603 5825 5603 4 gnd
port 138 nsew
rlabel metal3 s 5825 2443 5825 2443 4 gnd
port 138 nsew
rlabel metal3 s 5825 6767 5825 6767 4 gnd
port 138 nsew
rlabel metal3 s 5825 9137 5825 9137 4 gnd
port 138 nsew
rlabel metal3 s 5825 6393 5825 6393 4 gnd
port 138 nsew
rlabel metal3 s 5825 12297 5825 12297 4 gnd
port 138 nsew
rlabel metal3 s 5825 7973 5825 7973 4 gnd
port 138 nsew
rlabel metal3 s 5825 447 5825 447 4 gnd
port 138 nsew
rlabel metal3 s 3774 424 3774 424 4 gnd
port 138 nsew
rlabel metal3 s 3774 7534 3774 7534 4 gnd
port 138 nsew
rlabel metal3 s 5825 11507 5825 11507 4 gnd
port 138 nsew
rlabel metal3 s 5825 5187 5825 5187 4 gnd
port 138 nsew
rlabel metal3 s 5825 12713 5825 12713 4 gnd
port 138 nsew
rlabel metal3 s 5825 3607 5825 3607 4 gnd
port 138 nsew
rlabel metal3 s 3774 2794 3774 2794 4 gnd
port 138 nsew
rlabel metal3 s 4046 1214 4046 1214 4 vdd
port 137 nsew
rlabel metal3 s 5825 7183 5825 7183 4 gnd
port 138 nsew
rlabel metal3 s 5825 10343 5825 10343 4 gnd
port 138 nsew
rlabel metal3 s 4046 3584 4046 3584 4 vdd
port 137 nsew
rlabel metal3 s 5825 863 5825 863 4 gnd
port 138 nsew
rlabel metal3 s 3774 1214 3774 1214 4 gnd
port 138 nsew
rlabel metal3 s 7336 12274 7336 12274 4 vdd
port 137 nsew
rlabel metal3 s 7336 10299 7336 10299 4 vdd
port 137 nsew
rlabel metal3 s 7336 11089 7336 11089 4 vdd
port 137 nsew
rlabel metal3 s 7336 8324 7336 8324 4 vdd
port 137 nsew
rlabel metal3 s 7336 10694 7336 10694 4 vdd
port 137 nsew
rlabel metal3 s 7336 7929 7336 7929 4 vdd
port 137 nsew
rlabel metal3 s 7336 11879 7336 11879 4 vdd
port 137 nsew
rlabel metal3 s 7336 7139 7336 7139 4 vdd
port 137 nsew
rlabel metal3 s 7336 8719 7336 8719 4 vdd
port 137 nsew
rlabel metal3 s 7336 6744 7336 6744 4 vdd
port 137 nsew
rlabel metal3 s 7336 9904 7336 9904 4 vdd
port 137 nsew
rlabel metal3 s 7336 11484 7336 11484 4 vdd
port 137 nsew
rlabel metal3 s 7336 12669 7336 12669 4 vdd
port 137 nsew
rlabel metal3 s 7336 7534 7336 7534 4 vdd
port 137 nsew
rlabel metal3 s 7336 9114 7336 9114 4 vdd
port 137 nsew
rlabel metal3 s 7336 9509 7336 9509 4 vdd
port 137 nsew
rlabel metal3 s 7064 12274 7064 12274 4 gnd
port 138 nsew
rlabel metal3 s 6250 7125 6250 7125 4 vdd
port 137 nsew
rlabel metal3 s 6682 11507 6682 11507 4 vdd
port 137 nsew
rlabel metal3 s 6250 12297 6250 12297 4 vdd
port 137 nsew
rlabel metal3 s 7064 11484 7064 11484 4 gnd
port 138 nsew
rlabel metal3 s 6682 10717 6682 10717 4 vdd
port 137 nsew
rlabel metal3 s 6250 7915 6250 7915 4 vdd
port 137 nsew
rlabel metal3 s 7064 7139 7064 7139 4 gnd
port 138 nsew
rlabel metal3 s 6682 9927 6682 9927 4 vdd
port 137 nsew
rlabel metal3 s 6682 8705 6682 8705 4 vdd
port 137 nsew
rlabel metal3 s 7064 7534 7064 7534 4 gnd
port 138 nsew
rlabel metal3 s 6682 10285 6682 10285 4 vdd
port 137 nsew
rlabel metal3 s 7064 11089 7064 11089 4 gnd
port 138 nsew
rlabel metal3 s 6250 9137 6250 9137 4 vdd
port 137 nsew
rlabel metal3 s 6250 8705 6250 8705 4 vdd
port 137 nsew
rlabel metal3 s 7064 9114 7064 9114 4 gnd
port 138 nsew
rlabel metal3 s 6682 9137 6682 9137 4 vdd
port 137 nsew
rlabel metal3 s 6682 12297 6682 12297 4 vdd
port 137 nsew
rlabel metal3 s 6250 7557 6250 7557 4 vdd
port 137 nsew
rlabel metal3 s 6682 8347 6682 8347 4 vdd
port 137 nsew
rlabel metal3 s 6250 11865 6250 11865 4 vdd
port 137 nsew
rlabel metal3 s 7064 9904 7064 9904 4 gnd
port 138 nsew
rlabel metal3 s 6682 7915 6682 7915 4 vdd
port 137 nsew
rlabel metal3 s 7064 6744 7064 6744 4 gnd
port 138 nsew
rlabel metal3 s 7064 12669 7064 12669 4 gnd
port 138 nsew
rlabel metal3 s 6250 9927 6250 9927 4 vdd
port 137 nsew
rlabel metal3 s 6250 11075 6250 11075 4 vdd
port 137 nsew
rlabel metal3 s 7064 8324 7064 8324 4 gnd
port 138 nsew
rlabel metal3 s 6250 12655 6250 12655 4 vdd
port 137 nsew
rlabel metal3 s 6682 7557 6682 7557 4 vdd
port 137 nsew
rlabel metal3 s 6682 6767 6682 6767 4 vdd
port 137 nsew
rlabel metal3 s 6682 11075 6682 11075 4 vdd
port 137 nsew
rlabel metal3 s 6250 6767 6250 6767 4 vdd
port 137 nsew
rlabel metal3 s 7064 11879 7064 11879 4 gnd
port 138 nsew
rlabel metal3 s 6250 8347 6250 8347 4 vdd
port 137 nsew
rlabel metal3 s 7064 8719 7064 8719 4 gnd
port 138 nsew
rlabel metal3 s 6250 11507 6250 11507 4 vdd
port 137 nsew
rlabel metal3 s 6682 7125 6682 7125 4 vdd
port 137 nsew
rlabel metal3 s 7064 9509 7064 9509 4 gnd
port 138 nsew
rlabel metal3 s 6250 10285 6250 10285 4 vdd
port 137 nsew
rlabel metal3 s 6682 9495 6682 9495 4 vdd
port 137 nsew
rlabel metal3 s 7064 7929 7064 7929 4 gnd
port 138 nsew
rlabel metal3 s 6682 11865 6682 11865 4 vdd
port 137 nsew
rlabel metal3 s 6250 9495 6250 9495 4 vdd
port 137 nsew
rlabel metal3 s 6682 12655 6682 12655 4 vdd
port 137 nsew
rlabel metal3 s 7064 10694 7064 10694 4 gnd
port 138 nsew
rlabel metal3 s 6250 10717 6250 10717 4 vdd
port 137 nsew
rlabel metal3 s 7064 10299 7064 10299 4 gnd
port 138 nsew
rlabel metal3 s 6250 1237 6250 1237 4 vdd
port 137 nsew
rlabel metal3 s 7064 819 7064 819 4 gnd
port 138 nsew
rlabel metal3 s 7064 2794 7064 2794 4 gnd
port 138 nsew
rlabel metal3 s 6250 3607 6250 3607 4 vdd
port 137 nsew
rlabel metal3 s 6250 805 6250 805 4 vdd
port 137 nsew
rlabel metal3 s 6250 2027 6250 2027 4 vdd
port 137 nsew
rlabel metal3 s 7064 424 7064 424 4 gnd
port 138 nsew
rlabel metal3 s 6682 5977 6682 5977 4 vdd
port 137 nsew
rlabel metal3 s 6682 6335 6682 6335 4 vdd
port 137 nsew
rlabel metal3 s 6250 4397 6250 4397 4 vdd
port 137 nsew
rlabel metal3 s 7064 1214 7064 1214 4 gnd
port 138 nsew
rlabel metal3 s 6682 3965 6682 3965 4 vdd
port 137 nsew
rlabel metal3 s 6682 447 6682 447 4 vdd
port 137 nsew
rlabel metal3 s 6682 1595 6682 1595 4 vdd
port 137 nsew
rlabel metal3 s 6682 4755 6682 4755 4 vdd
port 137 nsew
rlabel metal3 s 6250 2385 6250 2385 4 vdd
port 137 nsew
rlabel metal3 s 7064 5559 7064 5559 4 gnd
port 138 nsew
rlabel metal3 s 6682 2027 6682 2027 4 vdd
port 137 nsew
rlabel metal3 s 6250 4755 6250 4755 4 vdd
port 137 nsew
rlabel metal3 s 6682 805 6682 805 4 vdd
port 137 nsew
rlabel metal3 s 6250 5977 6250 5977 4 vdd
port 137 nsew
rlabel metal3 s 6682 2385 6682 2385 4 vdd
port 137 nsew
rlabel metal3 s 6682 1237 6682 1237 4 vdd
port 137 nsew
rlabel metal3 s 7064 1609 7064 1609 4 gnd
port 138 nsew
rlabel metal3 s 7064 6349 7064 6349 4 gnd
port 138 nsew
rlabel metal3 s 7064 3584 7064 3584 4 gnd
port 138 nsew
rlabel metal3 s 7064 2399 7064 2399 4 gnd
port 138 nsew
rlabel metal3 s 6250 6335 6250 6335 4 vdd
port 137 nsew
rlabel metal3 s 6250 1595 6250 1595 4 vdd
port 137 nsew
rlabel metal3 s 6250 5187 6250 5187 4 vdd
port 137 nsew
rlabel metal3 s 6682 4397 6682 4397 4 vdd
port 137 nsew
rlabel metal3 s 6682 3175 6682 3175 4 vdd
port 137 nsew
rlabel metal3 s 6250 3175 6250 3175 4 vdd
port 137 nsew
rlabel metal3 s 6250 2817 6250 2817 4 vdd
port 137 nsew
rlabel metal3 s 7064 3189 7064 3189 4 gnd
port 138 nsew
rlabel metal3 s 6682 5545 6682 5545 4 vdd
port 137 nsew
rlabel metal3 s 6682 2817 6682 2817 4 vdd
port 137 nsew
rlabel metal3 s 7064 3979 7064 3979 4 gnd
port 138 nsew
rlabel metal3 s 6250 447 6250 447 4 vdd
port 137 nsew
rlabel metal3 s 6250 5545 6250 5545 4 vdd
port 137 nsew
rlabel metal3 s 7064 4769 7064 4769 4 gnd
port 138 nsew
rlabel metal3 s 6250 3965 6250 3965 4 vdd
port 137 nsew
rlabel metal3 s 7064 5164 7064 5164 4 gnd
port 138 nsew
rlabel metal3 s 6682 3607 6682 3607 4 vdd
port 137 nsew
rlabel metal3 s 7064 2004 7064 2004 4 gnd
port 138 nsew
rlabel metal3 s 7064 5954 7064 5954 4 gnd
port 138 nsew
rlabel metal3 s 6682 5187 6682 5187 4 vdd
port 137 nsew
rlabel metal3 s 7064 4374 7064 4374 4 gnd
port 138 nsew
rlabel metal3 s 7336 3979 7336 3979 4 vdd
port 137 nsew
rlabel metal3 s 7336 2794 7336 2794 4 vdd
port 137 nsew
rlabel metal3 s 7336 5164 7336 5164 4 vdd
port 137 nsew
rlabel metal3 s 7336 1609 7336 1609 4 vdd
port 137 nsew
rlabel metal3 s 7336 424 7336 424 4 vdd
port 137 nsew
rlabel metal3 s 7336 4769 7336 4769 4 vdd
port 137 nsew
rlabel metal3 s 7336 4374 7336 4374 4 vdd
port 137 nsew
rlabel metal3 s 7336 5954 7336 5954 4 vdd
port 137 nsew
rlabel metal3 s 7336 1214 7336 1214 4 vdd
port 137 nsew
rlabel metal3 s 7336 2399 7336 2399 4 vdd
port 137 nsew
rlabel metal3 s 7336 2004 7336 2004 4 vdd
port 137 nsew
rlabel metal3 s 7336 3584 7336 3584 4 vdd
port 137 nsew
rlabel metal3 s 7336 6349 7336 6349 4 vdd
port 137 nsew
rlabel metal3 s 7336 3189 7336 3189 4 vdd
port 137 nsew
rlabel metal3 s 7336 5559 7336 5559 4 vdd
port 137 nsew
rlabel metal3 s 7336 819 7336 819 4 vdd
port 137 nsew
<< properties >>
string FIXED_BBOX 0 0 11546 50588
string GDS_END 5254642
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 5096622
<< end >>
