magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 58
rect 2205 0 2208 58
<< via1 >>
rect 3 0 2205 58
<< metal2 >>
rect 0 0 3 58
rect 2205 0 2208 58
<< properties >>
string GDS_END 78965062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78956098
<< end >>
