magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 287 2982 582
rect -38 261 977 287
rect 1440 261 2982 287
<< pwell >>
rect 1034 157 1427 229
rect 1680 157 1864 201
rect 2449 157 2893 203
rect 1 93 2893 157
rect 1 21 993 93
rect 1287 21 2893 93
rect 29 -17 63 21
<< locali >>
rect 19 195 89 325
rect 339 153 383 344
rect 422 237 465 274
rect 422 153 513 237
rect 1005 221 1050 323
rect 1152 221 1243 333
rect 2551 259 2617 484
rect 2719 259 2785 484
rect 2551 214 2785 259
rect 2551 61 2617 214
rect 2719 61 2785 214
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2944 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 169 393
rect 123 161 169 359
rect 35 127 169 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 493
rect 271 378 357 493
rect 447 378 513 527
rect 271 103 305 378
rect 551 344 617 485
rect 653 365 692 527
rect 825 404 891 493
rect 927 442 993 493
rect 825 364 903 404
rect 499 271 617 344
rect 556 235 617 271
rect 761 264 835 330
rect 556 169 727 235
rect 271 51 357 103
rect 447 17 513 103
rect 556 51 601 169
rect 761 137 795 264
rect 869 230 903 364
rect 829 196 903 230
rect 937 357 993 442
rect 1031 401 1099 493
rect 1133 435 1202 527
rect 1335 430 1401 493
rect 1443 435 1651 475
rect 1031 367 1317 401
rect 637 17 703 122
rect 829 51 883 196
rect 937 165 971 357
rect 1084 187 1118 367
rect 1277 271 1317 367
rect 1351 373 1401 430
rect 1351 237 1385 373
rect 919 129 971 165
rect 919 51 959 129
rect 1052 103 1118 187
rect 993 51 1118 103
rect 1152 17 1202 181
rect 1303 113 1385 237
rect 1419 225 1456 344
rect 1490 331 1583 401
rect 1490 191 1524 331
rect 1617 315 1651 435
rect 1685 367 1732 527
rect 1617 297 1732 315
rect 1423 147 1524 191
rect 1562 263 1732 297
rect 1562 113 1596 263
rect 1698 249 1732 263
rect 1766 275 1832 493
rect 1874 421 1932 527
rect 2045 433 2222 471
rect 1634 213 1674 219
rect 1766 213 1949 275
rect 2018 249 2056 393
rect 1634 209 1949 213
rect 1634 153 1847 209
rect 2090 207 2154 399
rect 1303 51 1427 113
rect 1461 51 1596 113
rect 1649 17 1728 112
rect 1766 51 1847 153
rect 2061 141 2154 207
rect 2188 265 2222 433
rect 2256 427 2308 527
rect 2368 381 2436 493
rect 2256 306 2436 381
rect 2188 199 2362 265
rect 1893 17 1948 123
rect 2188 107 2222 199
rect 2398 165 2436 306
rect 2470 293 2517 527
rect 2651 293 2685 527
rect 2819 293 2871 527
rect 2065 66 2222 107
rect 2270 17 2333 123
rect 2370 60 2436 165
rect 2470 17 2517 180
rect 2651 17 2685 180
rect 2819 17 2871 256
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2944 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
<< metal1 >>
rect 0 561 2944 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2944 561
rect 0 496 2944 527
rect 0 17 2944 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2944 17
rect 0 -48 2944 -17
<< obsm1 >>
rect 115 388 173 397
rect 1490 388 1548 397
rect 2008 388 2066 397
rect 115 360 2066 388
rect 115 351 173 360
rect 1490 351 1548 360
rect 2008 351 2066 360
rect 191 320 249 329
rect 1408 320 1466 329
rect 2092 320 2150 329
rect 191 292 2150 320
rect 191 283 249 292
rect 1408 283 1466 292
rect 2092 283 2150 292
rect 749 184 807 193
rect 2388 184 2446 193
rect 749 156 2446 184
rect 749 147 807 156
rect 2388 147 2446 156
rect 259 116 317 125
rect 825 116 883 125
rect 259 79 883 116
rect 911 116 969 125
rect 1294 116 1352 125
rect 911 79 1352 116
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 339 153 383 344 6 D
port 2 nsew signal input
rlabel locali s 422 153 513 237 6 DE
port 3 nsew signal input
rlabel locali s 422 237 465 274 6 DE
port 3 nsew signal input
rlabel locali s 1152 221 1243 333 6 SCD
port 4 nsew signal input
rlabel locali s 1005 221 1050 323 6 SCE
port 5 nsew signal input
rlabel metal1 s 0 -48 2944 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1287 21 2893 93 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 993 93 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 93 2893 157 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2449 157 2893 203 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1680 157 1864 201 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1034 157 1427 229 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s 1440 261 2982 287 6 VPB
port 8 nsew power bidirectional
rlabel nwell s -38 261 977 287 6 VPB
port 8 nsew power bidirectional
rlabel nwell s -38 287 2982 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2944 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2719 61 2785 214 6 Q
port 10 nsew signal output
rlabel locali s 2551 61 2617 214 6 Q
port 10 nsew signal output
rlabel locali s 2551 214 2785 259 6 Q
port 10 nsew signal output
rlabel locali s 2719 259 2785 484 6 Q
port 10 nsew signal output
rlabel locali s 2551 259 2617 484 6 Q
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2944 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 557420
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 534544
<< end >>
