magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 0 953 7045 1121
rect 0 417 2199 953
rect 2505 417 7045 953
<< pwell >>
rect 82 96 2032 312
rect 2591 96 6970 312
rect 66 10 6979 96
<< mvnmos >>
rect 161 146 281 286
rect 337 146 457 286
rect 623 146 743 286
rect 909 146 1029 286
rect 1085 146 1205 286
rect 1371 146 1491 286
rect 1547 146 1667 286
rect 1833 146 1953 286
rect 2670 146 2790 286
rect 2956 146 3076 286
rect 3132 146 3252 286
rect 3421 146 3541 286
rect 3707 146 3827 286
rect 3883 146 4003 286
rect 4172 146 4292 286
rect 4348 146 4468 286
rect 4634 146 4754 286
rect 4810 146 4930 286
rect 5099 146 5219 286
rect 5275 146 5395 286
rect 5561 146 5681 286
rect 5847 146 5967 286
rect 6023 146 6143 286
rect 6309 146 6429 286
rect 6595 146 6715 286
rect 6771 146 6891 286
<< mvpmos >>
rect 161 752 281 952
rect 337 752 457 952
rect 623 752 743 952
rect 909 752 1029 952
rect 1085 752 1205 952
rect 1371 752 1491 952
rect 1547 752 1667 952
rect 1833 752 1953 952
rect 2670 752 2790 952
rect 2956 752 3076 952
rect 3132 752 3252 952
rect 3421 752 3541 952
rect 3707 752 3827 952
rect 3883 752 4003 952
rect 4172 752 4292 952
rect 4348 752 4468 952
rect 4634 752 4754 952
rect 4810 752 4930 952
rect 5099 752 5219 952
rect 5275 752 5395 952
rect 5561 752 5681 952
rect 5847 752 5967 952
rect 6023 752 6143 952
rect 6309 752 6429 952
rect 6595 752 6715 952
rect 6771 752 6891 952
rect 161 484 281 684
rect 337 484 457 684
rect 623 484 743 684
rect 909 484 1029 684
rect 1085 484 1205 684
rect 1371 484 1491 684
rect 1547 484 1667 684
rect 1833 484 1953 684
rect 2670 484 2790 684
rect 2956 484 3076 684
rect 3132 484 3252 684
rect 3421 484 3541 684
rect 3707 484 3827 684
rect 3883 484 4003 684
rect 4172 484 4292 684
rect 4348 484 4468 684
rect 4634 484 4754 684
rect 4810 484 4930 684
rect 5099 484 5219 684
rect 5275 484 5395 684
rect 5561 484 5681 684
rect 5847 484 5967 684
rect 6023 484 6143 684
rect 6309 484 6429 684
rect 6595 484 6715 684
rect 6771 484 6891 684
<< mvndiff >>
rect 108 274 161 286
rect 108 240 116 274
rect 150 240 161 274
rect 108 206 161 240
rect 108 172 116 206
rect 150 172 161 206
rect 108 146 161 172
rect 281 146 337 286
rect 457 274 510 286
rect 457 240 468 274
rect 502 240 510 274
rect 457 206 510 240
rect 457 172 468 206
rect 502 172 510 206
rect 457 146 510 172
rect 570 274 623 286
rect 570 240 578 274
rect 612 240 623 274
rect 570 206 623 240
rect 570 172 578 206
rect 612 172 623 206
rect 570 146 623 172
rect 743 274 796 286
rect 743 240 754 274
rect 788 240 796 274
rect 743 206 796 240
rect 743 172 754 206
rect 788 172 796 206
rect 743 146 796 172
rect 856 274 909 286
rect 856 240 864 274
rect 898 240 909 274
rect 856 206 909 240
rect 856 172 864 206
rect 898 172 909 206
rect 856 146 909 172
rect 1029 146 1085 286
rect 1205 274 1258 286
rect 1205 240 1216 274
rect 1250 240 1258 274
rect 1205 206 1258 240
rect 1205 172 1216 206
rect 1250 172 1258 206
rect 1205 146 1258 172
rect 1318 274 1371 286
rect 1318 240 1326 274
rect 1360 240 1371 274
rect 1318 206 1371 240
rect 1318 172 1326 206
rect 1360 172 1371 206
rect 1318 146 1371 172
rect 1491 146 1547 286
rect 1667 274 1720 286
rect 1667 240 1678 274
rect 1712 240 1720 274
rect 1667 206 1720 240
rect 1667 172 1678 206
rect 1712 172 1720 206
rect 1667 146 1720 172
rect 1780 274 1833 286
rect 1780 240 1788 274
rect 1822 240 1833 274
rect 1780 206 1833 240
rect 1780 172 1788 206
rect 1822 172 1833 206
rect 1780 146 1833 172
rect 1953 274 2006 286
rect 1953 240 1964 274
rect 1998 240 2006 274
rect 1953 206 2006 240
rect 1953 172 1964 206
rect 1998 172 2006 206
rect 1953 146 2006 172
rect 2617 274 2670 286
rect 2617 240 2625 274
rect 2659 240 2670 274
rect 2617 206 2670 240
rect 2617 172 2625 206
rect 2659 172 2670 206
rect 2617 146 2670 172
rect 2790 274 2843 286
rect 2790 240 2801 274
rect 2835 240 2843 274
rect 2790 206 2843 240
rect 2790 172 2801 206
rect 2835 172 2843 206
rect 2790 146 2843 172
rect 2903 274 2956 286
rect 2903 240 2911 274
rect 2945 240 2956 274
rect 2903 206 2956 240
rect 2903 172 2911 206
rect 2945 172 2956 206
rect 2903 146 2956 172
rect 3076 274 3132 286
rect 3076 240 3087 274
rect 3121 240 3132 274
rect 3076 206 3132 240
rect 3076 172 3087 206
rect 3121 172 3132 206
rect 3076 146 3132 172
rect 3252 274 3308 286
rect 3252 240 3263 274
rect 3297 240 3308 274
rect 3252 206 3308 240
rect 3252 172 3263 206
rect 3297 172 3308 206
rect 3252 146 3308 172
rect 3368 274 3421 286
rect 3368 240 3376 274
rect 3410 240 3421 274
rect 3368 206 3421 240
rect 3368 172 3376 206
rect 3410 172 3421 206
rect 3368 146 3421 172
rect 3541 274 3594 286
rect 3541 240 3552 274
rect 3586 240 3594 274
rect 3541 206 3594 240
rect 3541 172 3552 206
rect 3586 172 3594 206
rect 3541 146 3594 172
rect 3654 274 3707 286
rect 3654 240 3662 274
rect 3696 240 3707 274
rect 3654 206 3707 240
rect 3654 172 3662 206
rect 3696 172 3707 206
rect 3654 146 3707 172
rect 3827 274 3883 286
rect 3827 240 3838 274
rect 3872 240 3883 274
rect 3827 206 3883 240
rect 3827 172 3838 206
rect 3872 172 3883 206
rect 3827 146 3883 172
rect 4003 274 4059 286
rect 4003 240 4014 274
rect 4048 240 4059 274
rect 4003 206 4059 240
rect 4003 172 4014 206
rect 4048 172 4059 206
rect 4003 146 4059 172
rect 4119 274 4172 286
rect 4119 240 4127 274
rect 4161 240 4172 274
rect 4119 206 4172 240
rect 4119 172 4127 206
rect 4161 172 4172 206
rect 4119 146 4172 172
rect 4292 146 4348 286
rect 4468 274 4521 286
rect 4468 240 4479 274
rect 4513 240 4521 274
rect 4468 206 4521 240
rect 4468 172 4479 206
rect 4513 172 4521 206
rect 4468 146 4521 172
rect 4581 274 4634 286
rect 4581 240 4589 274
rect 4623 240 4634 274
rect 4581 206 4634 240
rect 4581 172 4589 206
rect 4623 172 4634 206
rect 4581 146 4634 172
rect 4754 274 4810 286
rect 4754 240 4765 274
rect 4799 240 4810 274
rect 4754 206 4810 240
rect 4754 172 4765 206
rect 4799 172 4810 206
rect 4754 146 4810 172
rect 4930 274 4986 286
rect 4930 240 4941 274
rect 4975 240 4986 274
rect 4930 206 4986 240
rect 4930 172 4941 206
rect 4975 172 4986 206
rect 4930 146 4986 172
rect 5046 274 5099 286
rect 5046 240 5054 274
rect 5088 240 5099 274
rect 5046 206 5099 240
rect 5046 172 5054 206
rect 5088 172 5099 206
rect 5046 146 5099 172
rect 5219 146 5275 286
rect 5395 274 5448 286
rect 5395 240 5406 274
rect 5440 240 5448 274
rect 5395 206 5448 240
rect 5395 172 5406 206
rect 5440 172 5448 206
rect 5395 146 5448 172
rect 5508 274 5561 286
rect 5508 240 5516 274
rect 5550 240 5561 274
rect 5508 206 5561 240
rect 5508 172 5516 206
rect 5550 172 5561 206
rect 5508 146 5561 172
rect 5681 274 5734 286
rect 5681 240 5692 274
rect 5726 240 5734 274
rect 5681 206 5734 240
rect 5681 172 5692 206
rect 5726 172 5734 206
rect 5681 146 5734 172
rect 5794 274 5847 286
rect 5794 240 5802 274
rect 5836 240 5847 274
rect 5794 206 5847 240
rect 5794 172 5802 206
rect 5836 172 5847 206
rect 5794 146 5847 172
rect 5967 146 6023 286
rect 6143 274 6196 286
rect 6143 240 6154 274
rect 6188 240 6196 274
rect 6143 206 6196 240
rect 6143 172 6154 206
rect 6188 172 6196 206
rect 6143 146 6196 172
rect 6256 274 6309 286
rect 6256 240 6264 274
rect 6298 240 6309 274
rect 6256 206 6309 240
rect 6256 172 6264 206
rect 6298 172 6309 206
rect 6256 146 6309 172
rect 6429 274 6482 286
rect 6429 240 6440 274
rect 6474 240 6482 274
rect 6429 206 6482 240
rect 6429 172 6440 206
rect 6474 172 6482 206
rect 6429 146 6482 172
rect 6542 274 6595 286
rect 6542 240 6550 274
rect 6584 240 6595 274
rect 6542 206 6595 240
rect 6542 172 6550 206
rect 6584 172 6595 206
rect 6542 146 6595 172
rect 6715 146 6771 286
rect 6891 274 6944 286
rect 6891 240 6902 274
rect 6936 240 6944 274
rect 6891 206 6944 240
rect 6891 172 6902 206
rect 6936 172 6944 206
rect 6891 146 6944 172
<< mvpdiff >>
rect 108 934 161 952
rect 108 900 116 934
rect 150 900 161 934
rect 108 866 161 900
rect 108 832 116 866
rect 150 832 161 866
rect 108 798 161 832
rect 108 764 116 798
rect 150 764 161 798
rect 108 752 161 764
rect 281 934 337 952
rect 281 900 292 934
rect 326 900 337 934
rect 281 866 337 900
rect 281 832 292 866
rect 326 832 337 866
rect 281 798 337 832
rect 281 764 292 798
rect 326 764 337 798
rect 281 752 337 764
rect 457 934 510 952
rect 457 900 468 934
rect 502 900 510 934
rect 457 866 510 900
rect 457 832 468 866
rect 502 832 510 866
rect 457 798 510 832
rect 457 764 468 798
rect 502 764 510 798
rect 457 752 510 764
rect 570 934 623 952
rect 570 900 578 934
rect 612 900 623 934
rect 570 866 623 900
rect 570 832 578 866
rect 612 832 623 866
rect 570 798 623 832
rect 570 764 578 798
rect 612 764 623 798
rect 570 752 623 764
rect 743 934 796 952
rect 743 900 754 934
rect 788 900 796 934
rect 743 866 796 900
rect 743 832 754 866
rect 788 832 796 866
rect 743 798 796 832
rect 743 764 754 798
rect 788 764 796 798
rect 743 752 796 764
rect 856 934 909 952
rect 856 900 864 934
rect 898 900 909 934
rect 856 866 909 900
rect 856 832 864 866
rect 898 832 909 866
rect 856 798 909 832
rect 856 764 864 798
rect 898 764 909 798
rect 856 752 909 764
rect 1029 934 1085 952
rect 1029 900 1040 934
rect 1074 900 1085 934
rect 1029 866 1085 900
rect 1029 832 1040 866
rect 1074 832 1085 866
rect 1029 798 1085 832
rect 1029 764 1040 798
rect 1074 764 1085 798
rect 1029 752 1085 764
rect 1205 934 1258 952
rect 1205 900 1216 934
rect 1250 900 1258 934
rect 1205 866 1258 900
rect 1205 832 1216 866
rect 1250 832 1258 866
rect 1205 798 1258 832
rect 1205 764 1216 798
rect 1250 764 1258 798
rect 1205 752 1258 764
rect 1318 934 1371 952
rect 1318 900 1326 934
rect 1360 900 1371 934
rect 1318 866 1371 900
rect 1318 832 1326 866
rect 1360 832 1371 866
rect 1318 798 1371 832
rect 1318 764 1326 798
rect 1360 764 1371 798
rect 1318 752 1371 764
rect 1491 934 1547 952
rect 1491 900 1502 934
rect 1536 900 1547 934
rect 1491 866 1547 900
rect 1491 832 1502 866
rect 1536 832 1547 866
rect 1491 798 1547 832
rect 1491 764 1502 798
rect 1536 764 1547 798
rect 1491 752 1547 764
rect 1667 934 1720 952
rect 1667 900 1678 934
rect 1712 900 1720 934
rect 1667 866 1720 900
rect 1667 832 1678 866
rect 1712 832 1720 866
rect 1667 798 1720 832
rect 1667 764 1678 798
rect 1712 764 1720 798
rect 1667 752 1720 764
rect 1780 934 1833 952
rect 1780 900 1788 934
rect 1822 900 1833 934
rect 1780 866 1833 900
rect 1780 832 1788 866
rect 1822 832 1833 866
rect 1780 798 1833 832
rect 1780 764 1788 798
rect 1822 764 1833 798
rect 1780 752 1833 764
rect 1953 934 2006 952
rect 1953 900 1964 934
rect 1998 900 2006 934
rect 1953 866 2006 900
rect 1953 832 1964 866
rect 1998 832 2006 866
rect 1953 798 2006 832
rect 1953 764 1964 798
rect 1998 764 2006 798
rect 1953 752 2006 764
rect 2617 934 2670 952
rect 2617 900 2625 934
rect 2659 900 2670 934
rect 2617 866 2670 900
rect 2617 832 2625 866
rect 2659 832 2670 866
rect 2617 798 2670 832
rect 2617 764 2625 798
rect 2659 764 2670 798
rect 2617 752 2670 764
rect 2790 934 2843 952
rect 2790 900 2801 934
rect 2835 900 2843 934
rect 2790 866 2843 900
rect 2790 832 2801 866
rect 2835 832 2843 866
rect 2790 798 2843 832
rect 2790 764 2801 798
rect 2835 764 2843 798
rect 2790 752 2843 764
rect 2903 934 2956 952
rect 2903 900 2911 934
rect 2945 900 2956 934
rect 2903 866 2956 900
rect 2903 832 2911 866
rect 2945 832 2956 866
rect 2903 798 2956 832
rect 2903 764 2911 798
rect 2945 764 2956 798
rect 2903 752 2956 764
rect 3076 934 3132 952
rect 3076 900 3087 934
rect 3121 900 3132 934
rect 3076 866 3132 900
rect 3076 832 3087 866
rect 3121 832 3132 866
rect 3076 798 3132 832
rect 3076 764 3087 798
rect 3121 764 3132 798
rect 3076 752 3132 764
rect 3252 934 3305 952
rect 3252 900 3263 934
rect 3297 900 3305 934
rect 3252 866 3305 900
rect 3252 832 3263 866
rect 3297 832 3305 866
rect 3252 798 3305 832
rect 3252 764 3263 798
rect 3297 764 3305 798
rect 3252 752 3305 764
rect 3368 934 3421 952
rect 3368 900 3376 934
rect 3410 900 3421 934
rect 3368 866 3421 900
rect 3368 832 3376 866
rect 3410 832 3421 866
rect 3368 798 3421 832
rect 3368 764 3376 798
rect 3410 764 3421 798
rect 3368 752 3421 764
rect 3541 934 3594 952
rect 3541 900 3552 934
rect 3586 900 3594 934
rect 3541 866 3594 900
rect 3541 832 3552 866
rect 3586 832 3594 866
rect 3541 798 3594 832
rect 3541 764 3552 798
rect 3586 764 3594 798
rect 3541 752 3594 764
rect 3654 934 3707 952
rect 3654 900 3662 934
rect 3696 900 3707 934
rect 3654 866 3707 900
rect 3654 832 3662 866
rect 3696 832 3707 866
rect 3654 798 3707 832
rect 3654 764 3662 798
rect 3696 764 3707 798
rect 3654 752 3707 764
rect 3827 934 3883 952
rect 3827 900 3838 934
rect 3872 900 3883 934
rect 3827 866 3883 900
rect 3827 832 3838 866
rect 3872 832 3883 866
rect 3827 798 3883 832
rect 3827 764 3838 798
rect 3872 764 3883 798
rect 3827 752 3883 764
rect 4003 934 4056 952
rect 4003 900 4014 934
rect 4048 900 4056 934
rect 4003 866 4056 900
rect 4003 832 4014 866
rect 4048 832 4056 866
rect 4003 798 4056 832
rect 4003 764 4014 798
rect 4048 764 4056 798
rect 4003 752 4056 764
rect 4119 934 4172 952
rect 4119 900 4127 934
rect 4161 900 4172 934
rect 4119 866 4172 900
rect 4119 832 4127 866
rect 4161 832 4172 866
rect 4119 798 4172 832
rect 4119 764 4127 798
rect 4161 764 4172 798
rect 4119 752 4172 764
rect 4292 934 4348 952
rect 4292 900 4303 934
rect 4337 900 4348 934
rect 4292 866 4348 900
rect 4292 832 4303 866
rect 4337 832 4348 866
rect 4292 798 4348 832
rect 4292 764 4303 798
rect 4337 764 4348 798
rect 4292 752 4348 764
rect 4468 934 4521 952
rect 4468 900 4479 934
rect 4513 900 4521 934
rect 4468 866 4521 900
rect 4468 832 4479 866
rect 4513 832 4521 866
rect 4468 798 4521 832
rect 4468 764 4479 798
rect 4513 764 4521 798
rect 4468 752 4521 764
rect 4581 934 4634 952
rect 4581 900 4589 934
rect 4623 900 4634 934
rect 4581 866 4634 900
rect 4581 832 4589 866
rect 4623 832 4634 866
rect 4581 798 4634 832
rect 4581 764 4589 798
rect 4623 764 4634 798
rect 4581 752 4634 764
rect 4754 934 4810 952
rect 4754 900 4765 934
rect 4799 900 4810 934
rect 4754 866 4810 900
rect 4754 832 4765 866
rect 4799 832 4810 866
rect 4754 798 4810 832
rect 4754 764 4765 798
rect 4799 764 4810 798
rect 4754 752 4810 764
rect 4930 934 4983 952
rect 4930 900 4941 934
rect 4975 900 4983 934
rect 4930 866 4983 900
rect 4930 832 4941 866
rect 4975 832 4983 866
rect 4930 798 4983 832
rect 4930 764 4941 798
rect 4975 764 4983 798
rect 4930 752 4983 764
rect 5046 934 5099 952
rect 5046 900 5054 934
rect 5088 900 5099 934
rect 5046 866 5099 900
rect 5046 832 5054 866
rect 5088 832 5099 866
rect 5046 798 5099 832
rect 5046 764 5054 798
rect 5088 764 5099 798
rect 5046 752 5099 764
rect 5219 934 5275 952
rect 5219 900 5230 934
rect 5264 900 5275 934
rect 5219 866 5275 900
rect 5219 832 5230 866
rect 5264 832 5275 866
rect 5219 798 5275 832
rect 5219 764 5230 798
rect 5264 764 5275 798
rect 5219 752 5275 764
rect 5395 934 5448 952
rect 5395 900 5406 934
rect 5440 900 5448 934
rect 5395 866 5448 900
rect 5395 832 5406 866
rect 5440 832 5448 866
rect 5395 798 5448 832
rect 5395 764 5406 798
rect 5440 764 5448 798
rect 5395 752 5448 764
rect 5508 934 5561 952
rect 5508 900 5516 934
rect 5550 900 5561 934
rect 5508 866 5561 900
rect 5508 832 5516 866
rect 5550 832 5561 866
rect 5508 798 5561 832
rect 5508 764 5516 798
rect 5550 764 5561 798
rect 5508 752 5561 764
rect 5681 934 5734 952
rect 5681 900 5692 934
rect 5726 900 5734 934
rect 5681 866 5734 900
rect 5681 832 5692 866
rect 5726 832 5734 866
rect 5681 798 5734 832
rect 5681 764 5692 798
rect 5726 764 5734 798
rect 5681 752 5734 764
rect 5794 934 5847 952
rect 5794 900 5802 934
rect 5836 900 5847 934
rect 5794 866 5847 900
rect 5794 832 5802 866
rect 5836 832 5847 866
rect 5794 798 5847 832
rect 5794 764 5802 798
rect 5836 764 5847 798
rect 5794 752 5847 764
rect 5967 934 6023 952
rect 5967 900 5978 934
rect 6012 900 6023 934
rect 5967 866 6023 900
rect 5967 832 5978 866
rect 6012 832 6023 866
rect 5967 798 6023 832
rect 5967 764 5978 798
rect 6012 764 6023 798
rect 5967 752 6023 764
rect 6143 934 6196 952
rect 6143 900 6154 934
rect 6188 900 6196 934
rect 6143 866 6196 900
rect 6143 832 6154 866
rect 6188 832 6196 866
rect 6143 798 6196 832
rect 6143 764 6154 798
rect 6188 764 6196 798
rect 6143 752 6196 764
rect 6256 934 6309 952
rect 6256 900 6264 934
rect 6298 900 6309 934
rect 6256 866 6309 900
rect 6256 832 6264 866
rect 6298 832 6309 866
rect 6256 798 6309 832
rect 6256 764 6264 798
rect 6298 764 6309 798
rect 6256 752 6309 764
rect 6429 934 6482 952
rect 6429 900 6440 934
rect 6474 900 6482 934
rect 6429 866 6482 900
rect 6429 832 6440 866
rect 6474 832 6482 866
rect 6429 798 6482 832
rect 6429 764 6440 798
rect 6474 764 6482 798
rect 6429 752 6482 764
rect 6542 934 6595 952
rect 6542 900 6550 934
rect 6584 900 6595 934
rect 6542 866 6595 900
rect 6542 832 6550 866
rect 6584 832 6595 866
rect 6542 798 6595 832
rect 6542 764 6550 798
rect 6584 764 6595 798
rect 6542 752 6595 764
rect 6715 934 6771 952
rect 6715 900 6726 934
rect 6760 900 6771 934
rect 6715 866 6771 900
rect 6715 832 6726 866
rect 6760 832 6771 866
rect 6715 798 6771 832
rect 6715 764 6726 798
rect 6760 764 6771 798
rect 6715 752 6771 764
rect 6891 934 6944 952
rect 6891 900 6902 934
rect 6936 900 6944 934
rect 6891 866 6944 900
rect 6891 832 6902 866
rect 6936 832 6944 866
rect 6891 798 6944 832
rect 6891 764 6902 798
rect 6936 764 6944 798
rect 6891 752 6944 764
rect 108 672 161 684
rect 108 638 116 672
rect 150 638 161 672
rect 108 604 161 638
rect 108 570 116 604
rect 150 570 161 604
rect 108 536 161 570
rect 108 502 116 536
rect 150 502 161 536
rect 108 484 161 502
rect 281 672 337 684
rect 281 638 292 672
rect 326 638 337 672
rect 281 604 337 638
rect 281 570 292 604
rect 326 570 337 604
rect 281 536 337 570
rect 281 502 292 536
rect 326 502 337 536
rect 281 484 337 502
rect 457 672 510 684
rect 457 638 468 672
rect 502 638 510 672
rect 457 604 510 638
rect 457 570 468 604
rect 502 570 510 604
rect 457 536 510 570
rect 457 502 468 536
rect 502 502 510 536
rect 457 484 510 502
rect 570 672 623 684
rect 570 638 578 672
rect 612 638 623 672
rect 570 604 623 638
rect 570 570 578 604
rect 612 570 623 604
rect 570 536 623 570
rect 570 502 578 536
rect 612 502 623 536
rect 570 484 623 502
rect 743 672 796 684
rect 743 638 754 672
rect 788 638 796 672
rect 743 604 796 638
rect 743 570 754 604
rect 788 570 796 604
rect 743 536 796 570
rect 743 502 754 536
rect 788 502 796 536
rect 743 484 796 502
rect 856 672 909 684
rect 856 638 864 672
rect 898 638 909 672
rect 856 604 909 638
rect 856 570 864 604
rect 898 570 909 604
rect 856 536 909 570
rect 856 502 864 536
rect 898 502 909 536
rect 856 484 909 502
rect 1029 672 1085 684
rect 1029 638 1040 672
rect 1074 638 1085 672
rect 1029 604 1085 638
rect 1029 570 1040 604
rect 1074 570 1085 604
rect 1029 536 1085 570
rect 1029 502 1040 536
rect 1074 502 1085 536
rect 1029 484 1085 502
rect 1205 672 1258 684
rect 1205 638 1216 672
rect 1250 638 1258 672
rect 1205 604 1258 638
rect 1205 570 1216 604
rect 1250 570 1258 604
rect 1205 536 1258 570
rect 1205 502 1216 536
rect 1250 502 1258 536
rect 1205 484 1258 502
rect 1318 672 1371 684
rect 1318 638 1326 672
rect 1360 638 1371 672
rect 1318 604 1371 638
rect 1318 570 1326 604
rect 1360 570 1371 604
rect 1318 536 1371 570
rect 1318 502 1326 536
rect 1360 502 1371 536
rect 1318 484 1371 502
rect 1491 672 1547 684
rect 1491 638 1502 672
rect 1536 638 1547 672
rect 1491 604 1547 638
rect 1491 570 1502 604
rect 1536 570 1547 604
rect 1491 536 1547 570
rect 1491 502 1502 536
rect 1536 502 1547 536
rect 1491 484 1547 502
rect 1667 672 1720 684
rect 1667 638 1678 672
rect 1712 638 1720 672
rect 1667 604 1720 638
rect 1667 570 1678 604
rect 1712 570 1720 604
rect 1667 536 1720 570
rect 1667 502 1678 536
rect 1712 502 1720 536
rect 1667 484 1720 502
rect 1780 672 1833 684
rect 1780 638 1788 672
rect 1822 638 1833 672
rect 1780 604 1833 638
rect 1780 570 1788 604
rect 1822 570 1833 604
rect 1780 536 1833 570
rect 1780 502 1788 536
rect 1822 502 1833 536
rect 1780 484 1833 502
rect 1953 672 2006 684
rect 1953 638 1964 672
rect 1998 638 2006 672
rect 1953 604 2006 638
rect 1953 570 1964 604
rect 1998 570 2006 604
rect 1953 536 2006 570
rect 1953 502 1964 536
rect 1998 502 2006 536
rect 1953 484 2006 502
rect 2617 672 2670 684
rect 2617 638 2625 672
rect 2659 638 2670 672
rect 2617 604 2670 638
rect 2617 570 2625 604
rect 2659 570 2670 604
rect 2617 536 2670 570
rect 2617 502 2625 536
rect 2659 502 2670 536
rect 2617 484 2670 502
rect 2790 672 2843 684
rect 2790 638 2801 672
rect 2835 638 2843 672
rect 2790 604 2843 638
rect 2790 570 2801 604
rect 2835 570 2843 604
rect 2790 536 2843 570
rect 2790 502 2801 536
rect 2835 502 2843 536
rect 2790 484 2843 502
rect 2903 672 2956 684
rect 2903 638 2911 672
rect 2945 638 2956 672
rect 2903 604 2956 638
rect 2903 570 2911 604
rect 2945 570 2956 604
rect 2903 536 2956 570
rect 2903 502 2911 536
rect 2945 502 2956 536
rect 2903 484 2956 502
rect 3076 672 3132 684
rect 3076 638 3087 672
rect 3121 638 3132 672
rect 3076 604 3132 638
rect 3076 570 3087 604
rect 3121 570 3132 604
rect 3076 484 3132 570
rect 3252 672 3305 684
rect 3252 638 3263 672
rect 3297 638 3305 672
rect 3252 604 3305 638
rect 3252 570 3263 604
rect 3297 570 3305 604
rect 3252 536 3305 570
rect 3252 502 3263 536
rect 3297 502 3305 536
rect 3252 484 3305 502
rect 3368 672 3421 684
rect 3368 638 3376 672
rect 3410 638 3421 672
rect 3368 604 3421 638
rect 3368 570 3376 604
rect 3410 570 3421 604
rect 3368 536 3421 570
rect 3368 502 3376 536
rect 3410 502 3421 536
rect 3368 484 3421 502
rect 3541 672 3594 684
rect 3541 638 3552 672
rect 3586 638 3594 672
rect 3541 604 3594 638
rect 3541 570 3552 604
rect 3586 570 3594 604
rect 3541 536 3594 570
rect 3541 502 3552 536
rect 3586 502 3594 536
rect 3541 484 3594 502
rect 3654 672 3707 684
rect 3654 638 3662 672
rect 3696 638 3707 672
rect 3654 604 3707 638
rect 3654 570 3662 604
rect 3696 570 3707 604
rect 3654 536 3707 570
rect 3654 502 3662 536
rect 3696 502 3707 536
rect 3654 484 3707 502
rect 3827 672 3883 684
rect 3827 638 3838 672
rect 3872 638 3883 672
rect 3827 604 3883 638
rect 3827 570 3838 604
rect 3872 570 3883 604
rect 3827 484 3883 570
rect 4003 672 4056 684
rect 4003 638 4014 672
rect 4048 638 4056 672
rect 4003 604 4056 638
rect 4003 570 4014 604
rect 4048 570 4056 604
rect 4003 536 4056 570
rect 4003 502 4014 536
rect 4048 502 4056 536
rect 4003 484 4056 502
rect 4119 672 4172 684
rect 4119 638 4127 672
rect 4161 638 4172 672
rect 4119 604 4172 638
rect 4119 570 4127 604
rect 4161 570 4172 604
rect 4119 536 4172 570
rect 4119 502 4127 536
rect 4161 502 4172 536
rect 4119 484 4172 502
rect 4292 672 4348 684
rect 4292 638 4303 672
rect 4337 638 4348 672
rect 4292 604 4348 638
rect 4292 570 4303 604
rect 4337 570 4348 604
rect 4292 536 4348 570
rect 4292 502 4303 536
rect 4337 502 4348 536
rect 4292 484 4348 502
rect 4468 672 4521 684
rect 4468 638 4479 672
rect 4513 638 4521 672
rect 4468 604 4521 638
rect 4468 570 4479 604
rect 4513 570 4521 604
rect 4468 536 4521 570
rect 4468 502 4479 536
rect 4513 502 4521 536
rect 4468 484 4521 502
rect 4581 672 4634 684
rect 4581 638 4589 672
rect 4623 638 4634 672
rect 4581 604 4634 638
rect 4581 570 4589 604
rect 4623 570 4634 604
rect 4581 536 4634 570
rect 4581 502 4589 536
rect 4623 502 4634 536
rect 4581 484 4634 502
rect 4754 672 4810 684
rect 4754 638 4765 672
rect 4799 638 4810 672
rect 4754 604 4810 638
rect 4754 570 4765 604
rect 4799 570 4810 604
rect 4754 484 4810 570
rect 4930 672 4983 684
rect 4930 638 4941 672
rect 4975 638 4983 672
rect 4930 604 4983 638
rect 4930 570 4941 604
rect 4975 570 4983 604
rect 4930 536 4983 570
rect 4930 502 4941 536
rect 4975 502 4983 536
rect 4930 484 4983 502
rect 5046 672 5099 684
rect 5046 638 5054 672
rect 5088 638 5099 672
rect 5046 604 5099 638
rect 5046 570 5054 604
rect 5088 570 5099 604
rect 5046 536 5099 570
rect 5046 502 5054 536
rect 5088 502 5099 536
rect 5046 484 5099 502
rect 5219 672 5275 684
rect 5219 638 5230 672
rect 5264 638 5275 672
rect 5219 604 5275 638
rect 5219 570 5230 604
rect 5264 570 5275 604
rect 5219 536 5275 570
rect 5219 502 5230 536
rect 5264 502 5275 536
rect 5219 484 5275 502
rect 5395 672 5448 684
rect 5395 638 5406 672
rect 5440 638 5448 672
rect 5395 604 5448 638
rect 5395 570 5406 604
rect 5440 570 5448 604
rect 5395 536 5448 570
rect 5395 502 5406 536
rect 5440 502 5448 536
rect 5395 484 5448 502
rect 5508 672 5561 684
rect 5508 638 5516 672
rect 5550 638 5561 672
rect 5508 604 5561 638
rect 5508 570 5516 604
rect 5550 570 5561 604
rect 5508 536 5561 570
rect 5508 502 5516 536
rect 5550 502 5561 536
rect 5508 484 5561 502
rect 5681 672 5734 684
rect 5681 638 5692 672
rect 5726 638 5734 672
rect 5681 604 5734 638
rect 5681 570 5692 604
rect 5726 570 5734 604
rect 5681 536 5734 570
rect 5681 502 5692 536
rect 5726 502 5734 536
rect 5681 484 5734 502
rect 5794 672 5847 684
rect 5794 638 5802 672
rect 5836 638 5847 672
rect 5794 604 5847 638
rect 5794 570 5802 604
rect 5836 570 5847 604
rect 5794 536 5847 570
rect 5794 502 5802 536
rect 5836 502 5847 536
rect 5794 484 5847 502
rect 5967 672 6023 684
rect 5967 638 5978 672
rect 6012 638 6023 672
rect 5967 604 6023 638
rect 5967 570 5978 604
rect 6012 570 6023 604
rect 5967 536 6023 570
rect 5967 502 5978 536
rect 6012 502 6023 536
rect 5967 484 6023 502
rect 6143 672 6196 684
rect 6143 638 6154 672
rect 6188 638 6196 672
rect 6143 604 6196 638
rect 6143 570 6154 604
rect 6188 570 6196 604
rect 6143 536 6196 570
rect 6143 502 6154 536
rect 6188 502 6196 536
rect 6143 484 6196 502
rect 6256 672 6309 684
rect 6256 638 6264 672
rect 6298 638 6309 672
rect 6256 604 6309 638
rect 6256 570 6264 604
rect 6298 570 6309 604
rect 6256 536 6309 570
rect 6256 502 6264 536
rect 6298 502 6309 536
rect 6256 484 6309 502
rect 6429 672 6482 684
rect 6429 638 6440 672
rect 6474 638 6482 672
rect 6429 604 6482 638
rect 6429 570 6440 604
rect 6474 570 6482 604
rect 6429 536 6482 570
rect 6429 502 6440 536
rect 6474 502 6482 536
rect 6429 484 6482 502
rect 6542 672 6595 684
rect 6542 638 6550 672
rect 6584 638 6595 672
rect 6542 604 6595 638
rect 6542 570 6550 604
rect 6584 570 6595 604
rect 6542 536 6595 570
rect 6542 502 6550 536
rect 6584 502 6595 536
rect 6542 484 6595 502
rect 6715 672 6771 684
rect 6715 638 6726 672
rect 6760 638 6771 672
rect 6715 604 6771 638
rect 6715 570 6726 604
rect 6760 570 6771 604
rect 6715 536 6771 570
rect 6715 502 6726 536
rect 6760 502 6771 536
rect 6715 484 6771 502
rect 6891 672 6944 684
rect 6891 638 6902 672
rect 6936 638 6944 672
rect 6891 604 6944 638
rect 6891 570 6902 604
rect 6936 570 6944 604
rect 6891 536 6944 570
rect 6891 502 6902 536
rect 6936 502 6944 536
rect 6891 484 6944 502
<< mvndiffc >>
rect 116 240 150 274
rect 116 172 150 206
rect 468 240 502 274
rect 468 172 502 206
rect 578 240 612 274
rect 578 172 612 206
rect 754 240 788 274
rect 754 172 788 206
rect 864 240 898 274
rect 864 172 898 206
rect 1216 240 1250 274
rect 1216 172 1250 206
rect 1326 240 1360 274
rect 1326 172 1360 206
rect 1678 240 1712 274
rect 1678 172 1712 206
rect 1788 240 1822 274
rect 1788 172 1822 206
rect 1964 240 1998 274
rect 1964 172 1998 206
rect 2625 240 2659 274
rect 2625 172 2659 206
rect 2801 240 2835 274
rect 2801 172 2835 206
rect 2911 240 2945 274
rect 2911 172 2945 206
rect 3087 240 3121 274
rect 3087 172 3121 206
rect 3263 240 3297 274
rect 3263 172 3297 206
rect 3376 240 3410 274
rect 3376 172 3410 206
rect 3552 240 3586 274
rect 3552 172 3586 206
rect 3662 240 3696 274
rect 3662 172 3696 206
rect 3838 240 3872 274
rect 3838 172 3872 206
rect 4014 240 4048 274
rect 4014 172 4048 206
rect 4127 240 4161 274
rect 4127 172 4161 206
rect 4479 240 4513 274
rect 4479 172 4513 206
rect 4589 240 4623 274
rect 4589 172 4623 206
rect 4765 240 4799 274
rect 4765 172 4799 206
rect 4941 240 4975 274
rect 4941 172 4975 206
rect 5054 240 5088 274
rect 5054 172 5088 206
rect 5406 240 5440 274
rect 5406 172 5440 206
rect 5516 240 5550 274
rect 5516 172 5550 206
rect 5692 240 5726 274
rect 5692 172 5726 206
rect 5802 240 5836 274
rect 5802 172 5836 206
rect 6154 240 6188 274
rect 6154 172 6188 206
rect 6264 240 6298 274
rect 6264 172 6298 206
rect 6440 240 6474 274
rect 6440 172 6474 206
rect 6550 240 6584 274
rect 6550 172 6584 206
rect 6902 240 6936 274
rect 6902 172 6936 206
<< mvpdiffc >>
rect 116 900 150 934
rect 116 832 150 866
rect 116 764 150 798
rect 292 900 326 934
rect 292 832 326 866
rect 292 764 326 798
rect 468 900 502 934
rect 468 832 502 866
rect 468 764 502 798
rect 578 900 612 934
rect 578 832 612 866
rect 578 764 612 798
rect 754 900 788 934
rect 754 832 788 866
rect 754 764 788 798
rect 864 900 898 934
rect 864 832 898 866
rect 864 764 898 798
rect 1040 900 1074 934
rect 1040 832 1074 866
rect 1040 764 1074 798
rect 1216 900 1250 934
rect 1216 832 1250 866
rect 1216 764 1250 798
rect 1326 900 1360 934
rect 1326 832 1360 866
rect 1326 764 1360 798
rect 1502 900 1536 934
rect 1502 832 1536 866
rect 1502 764 1536 798
rect 1678 900 1712 934
rect 1678 832 1712 866
rect 1678 764 1712 798
rect 1788 900 1822 934
rect 1788 832 1822 866
rect 1788 764 1822 798
rect 1964 900 1998 934
rect 1964 832 1998 866
rect 1964 764 1998 798
rect 2625 900 2659 934
rect 2625 832 2659 866
rect 2625 764 2659 798
rect 2801 900 2835 934
rect 2801 832 2835 866
rect 2801 764 2835 798
rect 2911 900 2945 934
rect 2911 832 2945 866
rect 2911 764 2945 798
rect 3087 900 3121 934
rect 3087 832 3121 866
rect 3087 764 3121 798
rect 3263 900 3297 934
rect 3263 832 3297 866
rect 3263 764 3297 798
rect 3376 900 3410 934
rect 3376 832 3410 866
rect 3376 764 3410 798
rect 3552 900 3586 934
rect 3552 832 3586 866
rect 3552 764 3586 798
rect 3662 900 3696 934
rect 3662 832 3696 866
rect 3662 764 3696 798
rect 3838 900 3872 934
rect 3838 832 3872 866
rect 3838 764 3872 798
rect 4014 900 4048 934
rect 4014 832 4048 866
rect 4014 764 4048 798
rect 4127 900 4161 934
rect 4127 832 4161 866
rect 4127 764 4161 798
rect 4303 900 4337 934
rect 4303 832 4337 866
rect 4303 764 4337 798
rect 4479 900 4513 934
rect 4479 832 4513 866
rect 4479 764 4513 798
rect 4589 900 4623 934
rect 4589 832 4623 866
rect 4589 764 4623 798
rect 4765 900 4799 934
rect 4765 832 4799 866
rect 4765 764 4799 798
rect 4941 900 4975 934
rect 4941 832 4975 866
rect 4941 764 4975 798
rect 5054 900 5088 934
rect 5054 832 5088 866
rect 5054 764 5088 798
rect 5230 900 5264 934
rect 5230 832 5264 866
rect 5230 764 5264 798
rect 5406 900 5440 934
rect 5406 832 5440 866
rect 5406 764 5440 798
rect 5516 900 5550 934
rect 5516 832 5550 866
rect 5516 764 5550 798
rect 5692 900 5726 934
rect 5692 832 5726 866
rect 5692 764 5726 798
rect 5802 900 5836 934
rect 5802 832 5836 866
rect 5802 764 5836 798
rect 5978 900 6012 934
rect 5978 832 6012 866
rect 5978 764 6012 798
rect 6154 900 6188 934
rect 6154 832 6188 866
rect 6154 764 6188 798
rect 6264 900 6298 934
rect 6264 832 6298 866
rect 6264 764 6298 798
rect 6440 900 6474 934
rect 6440 832 6474 866
rect 6440 764 6474 798
rect 6550 900 6584 934
rect 6550 832 6584 866
rect 6550 764 6584 798
rect 6726 900 6760 934
rect 6726 832 6760 866
rect 6726 764 6760 798
rect 6902 900 6936 934
rect 6902 832 6936 866
rect 6902 764 6936 798
rect 116 638 150 672
rect 116 570 150 604
rect 116 502 150 536
rect 292 638 326 672
rect 292 570 326 604
rect 292 502 326 536
rect 468 638 502 672
rect 468 570 502 604
rect 468 502 502 536
rect 578 638 612 672
rect 578 570 612 604
rect 578 502 612 536
rect 754 638 788 672
rect 754 570 788 604
rect 754 502 788 536
rect 864 638 898 672
rect 864 570 898 604
rect 864 502 898 536
rect 1040 638 1074 672
rect 1040 570 1074 604
rect 1040 502 1074 536
rect 1216 638 1250 672
rect 1216 570 1250 604
rect 1216 502 1250 536
rect 1326 638 1360 672
rect 1326 570 1360 604
rect 1326 502 1360 536
rect 1502 638 1536 672
rect 1502 570 1536 604
rect 1502 502 1536 536
rect 1678 638 1712 672
rect 1678 570 1712 604
rect 1678 502 1712 536
rect 1788 638 1822 672
rect 1788 570 1822 604
rect 1788 502 1822 536
rect 1964 638 1998 672
rect 1964 570 1998 604
rect 1964 502 1998 536
rect 2625 638 2659 672
rect 2625 570 2659 604
rect 2625 502 2659 536
rect 2801 638 2835 672
rect 2801 570 2835 604
rect 2801 502 2835 536
rect 2911 638 2945 672
rect 2911 570 2945 604
rect 2911 502 2945 536
rect 3087 638 3121 672
rect 3087 570 3121 604
rect 3263 638 3297 672
rect 3263 570 3297 604
rect 3263 502 3297 536
rect 3376 638 3410 672
rect 3376 570 3410 604
rect 3376 502 3410 536
rect 3552 638 3586 672
rect 3552 570 3586 604
rect 3552 502 3586 536
rect 3662 638 3696 672
rect 3662 570 3696 604
rect 3662 502 3696 536
rect 3838 638 3872 672
rect 3838 570 3872 604
rect 4014 638 4048 672
rect 4014 570 4048 604
rect 4014 502 4048 536
rect 4127 638 4161 672
rect 4127 570 4161 604
rect 4127 502 4161 536
rect 4303 638 4337 672
rect 4303 570 4337 604
rect 4303 502 4337 536
rect 4479 638 4513 672
rect 4479 570 4513 604
rect 4479 502 4513 536
rect 4589 638 4623 672
rect 4589 570 4623 604
rect 4589 502 4623 536
rect 4765 638 4799 672
rect 4765 570 4799 604
rect 4941 638 4975 672
rect 4941 570 4975 604
rect 4941 502 4975 536
rect 5054 638 5088 672
rect 5054 570 5088 604
rect 5054 502 5088 536
rect 5230 638 5264 672
rect 5230 570 5264 604
rect 5230 502 5264 536
rect 5406 638 5440 672
rect 5406 570 5440 604
rect 5406 502 5440 536
rect 5516 638 5550 672
rect 5516 570 5550 604
rect 5516 502 5550 536
rect 5692 638 5726 672
rect 5692 570 5726 604
rect 5692 502 5726 536
rect 5802 638 5836 672
rect 5802 570 5836 604
rect 5802 502 5836 536
rect 5978 638 6012 672
rect 5978 570 6012 604
rect 5978 502 6012 536
rect 6154 638 6188 672
rect 6154 570 6188 604
rect 6154 502 6188 536
rect 6264 638 6298 672
rect 6264 570 6298 604
rect 6264 502 6298 536
rect 6440 638 6474 672
rect 6440 570 6474 604
rect 6440 502 6474 536
rect 6550 638 6584 672
rect 6550 570 6584 604
rect 6550 502 6584 536
rect 6726 638 6760 672
rect 6726 570 6760 604
rect 6726 502 6760 536
rect 6902 638 6936 672
rect 6902 570 6936 604
rect 6902 502 6936 536
<< mvpsubdiff >>
rect 92 36 116 70
rect 150 36 185 70
rect 219 36 254 70
rect 288 36 323 70
rect 357 36 392 70
rect 426 36 461 70
rect 495 36 530 70
rect 564 36 599 70
rect 633 36 668 70
rect 702 36 737 70
rect 771 36 806 70
rect 840 36 875 70
rect 909 36 944 70
rect 978 36 1013 70
rect 1047 36 1082 70
rect 1116 36 1151 70
rect 1185 36 1220 70
rect 1254 36 1289 70
rect 1323 36 1358 70
rect 1392 36 1427 70
rect 1461 36 1496 70
rect 1530 36 1565 70
rect 1599 36 1634 70
rect 1668 36 1703 70
rect 1737 36 1772 70
rect 1806 36 1841 70
rect 1875 36 1910 70
rect 1944 36 1979 70
rect 2013 36 2048 70
rect 2082 36 2117 70
rect 2151 36 2186 70
rect 2220 36 2255 70
rect 2289 36 2324 70
rect 2358 36 2393 70
rect 2427 36 2462 70
rect 2496 36 2531 70
rect 2565 36 2600 70
rect 2634 36 2669 70
rect 2703 36 2738 70
rect 2772 36 2807 70
rect 2841 36 2876 70
rect 2910 36 2945 70
rect 2979 36 3014 70
rect 3048 36 3083 70
rect 3117 36 3152 70
rect 3186 36 3221 70
rect 3255 36 3290 70
rect 3324 36 3359 70
rect 3393 36 3427 70
rect 3461 36 3495 70
rect 3529 36 3563 70
rect 3597 36 3631 70
rect 3665 36 3699 70
rect 3733 36 3767 70
rect 3801 36 3835 70
rect 3869 36 3903 70
rect 3937 36 3971 70
rect 4005 36 4039 70
rect 4073 36 4107 70
rect 4141 36 4175 70
rect 4209 36 4243 70
rect 4277 36 4311 70
rect 4345 36 4379 70
rect 4413 36 4447 70
rect 4481 36 4515 70
rect 4549 36 4583 70
rect 4617 36 4651 70
rect 4685 36 4719 70
rect 4753 36 4787 70
rect 4821 36 4855 70
rect 4889 36 4923 70
rect 4957 36 4991 70
rect 5025 36 5059 70
rect 5093 36 5127 70
rect 5161 36 5195 70
rect 5229 36 5263 70
rect 5297 36 5331 70
rect 5365 36 5399 70
rect 5433 36 5467 70
rect 5501 36 5535 70
rect 5569 36 5603 70
rect 5637 36 5671 70
rect 5705 36 5739 70
rect 5773 36 5807 70
rect 5841 36 5875 70
rect 5909 36 5943 70
rect 5977 36 6011 70
rect 6045 36 6079 70
rect 6113 36 6147 70
rect 6181 36 6215 70
rect 6249 36 6283 70
rect 6317 36 6351 70
rect 6385 36 6419 70
rect 6453 36 6487 70
rect 6521 36 6555 70
rect 6589 36 6623 70
rect 6657 36 6691 70
rect 6725 36 6759 70
rect 6793 36 6827 70
rect 6861 36 6895 70
rect 6929 36 6953 70
<< mvnsubdiff >>
rect 67 1020 110 1054
rect 144 1020 178 1054
rect 212 1020 246 1054
rect 280 1020 314 1054
rect 348 1020 382 1054
rect 416 1020 450 1054
rect 484 1020 518 1054
rect 552 1020 586 1054
rect 620 1020 654 1054
rect 688 1020 722 1054
rect 756 1020 790 1054
rect 824 1020 858 1054
rect 892 1020 926 1054
rect 960 1020 994 1054
rect 1028 1020 1062 1054
rect 1096 1020 1130 1054
rect 1164 1020 1198 1054
rect 1232 1020 1266 1054
rect 1300 1020 1334 1054
rect 1368 1020 1402 1054
rect 1436 1020 1470 1054
rect 1504 1020 1538 1054
rect 1572 1020 1606 1054
rect 1640 1020 1674 1054
rect 1708 1020 1742 1054
rect 1776 1020 1810 1054
rect 1844 1020 1878 1054
rect 1912 1020 1946 1054
rect 1980 1020 2014 1054
rect 2048 1020 2082 1054
rect 2116 1020 2150 1054
rect 2184 1020 2218 1054
rect 2252 1020 2286 1054
rect 2320 1020 2354 1054
rect 2388 1020 2422 1054
rect 2456 1020 2490 1054
rect 2524 1020 2558 1054
rect 2592 1020 2626 1054
rect 2660 1020 2694 1054
rect 2728 1020 2762 1054
rect 2796 1020 2830 1054
rect 2864 1020 2898 1054
rect 2932 1020 2966 1054
rect 3000 1020 3034 1054
rect 3068 1020 3102 1054
rect 3136 1020 3170 1054
rect 3204 1020 3238 1054
rect 3272 1020 3306 1054
rect 3340 1020 3374 1054
rect 3408 1020 3442 1054
rect 3476 1020 3510 1054
rect 3544 1020 3578 1054
rect 3612 1020 3646 1054
rect 3680 1020 3714 1054
rect 3748 1020 3782 1054
rect 3816 1020 3850 1054
rect 3884 1020 3918 1054
rect 3952 1020 3986 1054
rect 4020 1020 4054 1054
rect 4088 1020 4122 1054
rect 4156 1020 4190 1054
rect 4224 1020 4258 1054
rect 4292 1020 4326 1054
rect 4360 1020 4394 1054
rect 4428 1020 4462 1054
rect 4496 1020 4530 1054
rect 4564 1020 4598 1054
rect 4632 1020 4666 1054
rect 4700 1020 4734 1054
rect 4768 1020 4802 1054
rect 4836 1020 4870 1054
rect 4904 1020 4938 1054
rect 4972 1020 5006 1054
rect 5040 1020 5074 1054
rect 5108 1020 5142 1054
rect 5176 1020 5210 1054
rect 5244 1020 5278 1054
rect 5312 1020 5346 1054
rect 5380 1020 5414 1054
rect 5448 1020 5482 1054
rect 5516 1020 5550 1054
rect 5584 1020 5618 1054
rect 5652 1020 5686 1054
rect 5720 1020 5754 1054
rect 5788 1020 5822 1054
rect 5856 1020 5890 1054
rect 5924 1020 5958 1054
rect 5992 1020 6026 1054
rect 6060 1020 6094 1054
rect 6128 1020 6162 1054
rect 6196 1020 6230 1054
rect 6264 1020 6298 1054
rect 6332 1020 6366 1054
rect 6400 1020 6434 1054
rect 6468 1020 6502 1054
rect 6536 1020 6570 1054
rect 6604 1020 6638 1054
rect 6672 1020 6706 1054
rect 6740 1020 6774 1054
rect 6808 1020 6842 1054
rect 6876 1020 6910 1054
rect 6944 1020 6978 1054
<< mvpsubdiffcont >>
rect 116 36 150 70
rect 185 36 219 70
rect 254 36 288 70
rect 323 36 357 70
rect 392 36 426 70
rect 461 36 495 70
rect 530 36 564 70
rect 599 36 633 70
rect 668 36 702 70
rect 737 36 771 70
rect 806 36 840 70
rect 875 36 909 70
rect 944 36 978 70
rect 1013 36 1047 70
rect 1082 36 1116 70
rect 1151 36 1185 70
rect 1220 36 1254 70
rect 1289 36 1323 70
rect 1358 36 1392 70
rect 1427 36 1461 70
rect 1496 36 1530 70
rect 1565 36 1599 70
rect 1634 36 1668 70
rect 1703 36 1737 70
rect 1772 36 1806 70
rect 1841 36 1875 70
rect 1910 36 1944 70
rect 1979 36 2013 70
rect 2048 36 2082 70
rect 2117 36 2151 70
rect 2186 36 2220 70
rect 2255 36 2289 70
rect 2324 36 2358 70
rect 2393 36 2427 70
rect 2462 36 2496 70
rect 2531 36 2565 70
rect 2600 36 2634 70
rect 2669 36 2703 70
rect 2738 36 2772 70
rect 2807 36 2841 70
rect 2876 36 2910 70
rect 2945 36 2979 70
rect 3014 36 3048 70
rect 3083 36 3117 70
rect 3152 36 3186 70
rect 3221 36 3255 70
rect 3290 36 3324 70
rect 3359 36 3393 70
rect 3427 36 3461 70
rect 3495 36 3529 70
rect 3563 36 3597 70
rect 3631 36 3665 70
rect 3699 36 3733 70
rect 3767 36 3801 70
rect 3835 36 3869 70
rect 3903 36 3937 70
rect 3971 36 4005 70
rect 4039 36 4073 70
rect 4107 36 4141 70
rect 4175 36 4209 70
rect 4243 36 4277 70
rect 4311 36 4345 70
rect 4379 36 4413 70
rect 4447 36 4481 70
rect 4515 36 4549 70
rect 4583 36 4617 70
rect 4651 36 4685 70
rect 4719 36 4753 70
rect 4787 36 4821 70
rect 4855 36 4889 70
rect 4923 36 4957 70
rect 4991 36 5025 70
rect 5059 36 5093 70
rect 5127 36 5161 70
rect 5195 36 5229 70
rect 5263 36 5297 70
rect 5331 36 5365 70
rect 5399 36 5433 70
rect 5467 36 5501 70
rect 5535 36 5569 70
rect 5603 36 5637 70
rect 5671 36 5705 70
rect 5739 36 5773 70
rect 5807 36 5841 70
rect 5875 36 5909 70
rect 5943 36 5977 70
rect 6011 36 6045 70
rect 6079 36 6113 70
rect 6147 36 6181 70
rect 6215 36 6249 70
rect 6283 36 6317 70
rect 6351 36 6385 70
rect 6419 36 6453 70
rect 6487 36 6521 70
rect 6555 36 6589 70
rect 6623 36 6657 70
rect 6691 36 6725 70
rect 6759 36 6793 70
rect 6827 36 6861 70
rect 6895 36 6929 70
<< mvnsubdiffcont >>
rect 110 1020 144 1054
rect 178 1020 212 1054
rect 246 1020 280 1054
rect 314 1020 348 1054
rect 382 1020 416 1054
rect 450 1020 484 1054
rect 518 1020 552 1054
rect 586 1020 620 1054
rect 654 1020 688 1054
rect 722 1020 756 1054
rect 790 1020 824 1054
rect 858 1020 892 1054
rect 926 1020 960 1054
rect 994 1020 1028 1054
rect 1062 1020 1096 1054
rect 1130 1020 1164 1054
rect 1198 1020 1232 1054
rect 1266 1020 1300 1054
rect 1334 1020 1368 1054
rect 1402 1020 1436 1054
rect 1470 1020 1504 1054
rect 1538 1020 1572 1054
rect 1606 1020 1640 1054
rect 1674 1020 1708 1054
rect 1742 1020 1776 1054
rect 1810 1020 1844 1054
rect 1878 1020 1912 1054
rect 1946 1020 1980 1054
rect 2014 1020 2048 1054
rect 2082 1020 2116 1054
rect 2150 1020 2184 1054
rect 2218 1020 2252 1054
rect 2286 1020 2320 1054
rect 2354 1020 2388 1054
rect 2422 1020 2456 1054
rect 2490 1020 2524 1054
rect 2558 1020 2592 1054
rect 2626 1020 2660 1054
rect 2694 1020 2728 1054
rect 2762 1020 2796 1054
rect 2830 1020 2864 1054
rect 2898 1020 2932 1054
rect 2966 1020 3000 1054
rect 3034 1020 3068 1054
rect 3102 1020 3136 1054
rect 3170 1020 3204 1054
rect 3238 1020 3272 1054
rect 3306 1020 3340 1054
rect 3374 1020 3408 1054
rect 3442 1020 3476 1054
rect 3510 1020 3544 1054
rect 3578 1020 3612 1054
rect 3646 1020 3680 1054
rect 3714 1020 3748 1054
rect 3782 1020 3816 1054
rect 3850 1020 3884 1054
rect 3918 1020 3952 1054
rect 3986 1020 4020 1054
rect 4054 1020 4088 1054
rect 4122 1020 4156 1054
rect 4190 1020 4224 1054
rect 4258 1020 4292 1054
rect 4326 1020 4360 1054
rect 4394 1020 4428 1054
rect 4462 1020 4496 1054
rect 4530 1020 4564 1054
rect 4598 1020 4632 1054
rect 4666 1020 4700 1054
rect 4734 1020 4768 1054
rect 4802 1020 4836 1054
rect 4870 1020 4904 1054
rect 4938 1020 4972 1054
rect 5006 1020 5040 1054
rect 5074 1020 5108 1054
rect 5142 1020 5176 1054
rect 5210 1020 5244 1054
rect 5278 1020 5312 1054
rect 5346 1020 5380 1054
rect 5414 1020 5448 1054
rect 5482 1020 5516 1054
rect 5550 1020 5584 1054
rect 5618 1020 5652 1054
rect 5686 1020 5720 1054
rect 5754 1020 5788 1054
rect 5822 1020 5856 1054
rect 5890 1020 5924 1054
rect 5958 1020 5992 1054
rect 6026 1020 6060 1054
rect 6094 1020 6128 1054
rect 6162 1020 6196 1054
rect 6230 1020 6264 1054
rect 6298 1020 6332 1054
rect 6366 1020 6400 1054
rect 6434 1020 6468 1054
rect 6502 1020 6536 1054
rect 6570 1020 6604 1054
rect 6638 1020 6672 1054
rect 6706 1020 6740 1054
rect 6774 1020 6808 1054
rect 6842 1020 6876 1054
rect 6910 1020 6944 1054
<< poly >>
rect 161 952 281 978
rect 337 952 457 978
rect 623 952 743 978
rect 909 952 1029 978
rect 1085 952 1205 978
rect 1371 952 1491 978
rect 1547 952 1667 978
rect 1833 952 1953 978
rect 2670 952 2790 978
rect 2956 952 3076 978
rect 3132 952 3252 978
rect 3421 952 3541 978
rect 3707 952 3827 978
rect 3883 952 4003 978
rect 4172 952 4292 978
rect 4348 952 4468 978
rect 4634 952 4754 978
rect 4810 952 4930 978
rect 5099 952 5219 978
rect 5275 952 5395 978
rect 5561 952 5681 978
rect 5847 952 5967 978
rect 6023 952 6143 978
rect 6309 952 6429 978
rect 6595 952 6715 978
rect 6771 952 6891 978
rect 161 684 281 752
rect 337 684 457 752
rect 623 684 743 752
rect 909 684 1029 752
rect 1085 684 1205 752
rect 1371 684 1491 752
rect 1547 684 1667 752
rect 1833 684 1953 752
rect 2670 684 2790 752
rect 2956 684 3076 752
rect 3132 684 3252 752
rect 3421 684 3541 752
rect 3707 684 3827 752
rect 3883 684 4003 752
rect 4172 684 4292 752
rect 4348 684 4468 752
rect 4634 684 4754 752
rect 4810 684 4930 752
rect 5099 684 5219 752
rect 5275 684 5395 752
rect 5561 684 5681 752
rect 5847 684 5967 752
rect 6023 684 6143 752
rect 6309 684 6429 752
rect 6595 684 6715 752
rect 6771 684 6891 752
rect 161 436 281 484
rect 161 402 207 436
rect 241 402 281 436
rect 161 368 281 402
rect 161 334 207 368
rect 241 334 281 368
rect 161 286 281 334
rect 337 436 457 484
rect 337 402 378 436
rect 412 402 457 436
rect 337 368 457 402
rect 337 334 378 368
rect 412 334 457 368
rect 337 286 457 334
rect 623 436 743 484
rect 623 402 667 436
rect 701 402 743 436
rect 623 368 743 402
rect 623 334 667 368
rect 701 334 743 368
rect 623 286 743 334
rect 909 436 1029 484
rect 909 402 954 436
rect 988 402 1029 436
rect 909 368 1029 402
rect 909 334 954 368
rect 988 334 1029 368
rect 909 286 1029 334
rect 1085 436 1205 484
rect 1085 402 1125 436
rect 1159 402 1205 436
rect 1085 368 1205 402
rect 1085 334 1125 368
rect 1159 334 1205 368
rect 1085 286 1205 334
rect 1371 436 1491 484
rect 1371 402 1417 436
rect 1451 402 1491 436
rect 1371 368 1491 402
rect 1371 334 1417 368
rect 1451 334 1491 368
rect 1371 286 1491 334
rect 1547 436 1667 484
rect 1547 402 1588 436
rect 1622 402 1667 436
rect 1547 368 1667 402
rect 1547 334 1588 368
rect 1622 334 1667 368
rect 1547 286 1667 334
rect 1833 436 1953 484
rect 1833 402 1877 436
rect 1911 402 1953 436
rect 1833 368 1953 402
rect 1833 334 1877 368
rect 1911 334 1953 368
rect 1833 286 1953 334
rect 2670 436 2790 484
rect 2670 402 2714 436
rect 2748 402 2790 436
rect 2670 368 2790 402
rect 2670 334 2714 368
rect 2748 334 2790 368
rect 2670 286 2790 334
rect 2956 436 3076 484
rect 2956 402 2999 436
rect 3033 402 3076 436
rect 2956 368 3076 402
rect 2956 334 2999 368
rect 3033 334 3076 368
rect 2956 286 3076 334
rect 3132 436 3252 484
rect 3132 402 3177 436
rect 3211 402 3252 436
rect 3132 368 3252 402
rect 3132 334 3177 368
rect 3211 334 3252 368
rect 3132 286 3252 334
rect 3421 436 3541 484
rect 3421 402 3465 436
rect 3499 402 3541 436
rect 3421 368 3541 402
rect 3421 334 3465 368
rect 3499 334 3541 368
rect 3421 286 3541 334
rect 3707 436 3827 484
rect 3707 402 3750 436
rect 3784 402 3827 436
rect 3707 368 3827 402
rect 3707 334 3750 368
rect 3784 334 3827 368
rect 3707 286 3827 334
rect 3883 436 4003 484
rect 3883 402 3928 436
rect 3962 402 4003 436
rect 3883 368 4003 402
rect 3883 334 3928 368
rect 3962 334 4003 368
rect 3883 286 4003 334
rect 4172 436 4292 484
rect 4172 402 4217 436
rect 4251 402 4292 436
rect 4172 368 4292 402
rect 4172 334 4217 368
rect 4251 334 4292 368
rect 4172 286 4292 334
rect 4348 436 4468 484
rect 4348 402 4388 436
rect 4422 402 4468 436
rect 4348 368 4468 402
rect 4348 334 4388 368
rect 4422 334 4468 368
rect 4348 286 4468 334
rect 4634 436 4754 484
rect 4634 402 4677 436
rect 4711 402 4754 436
rect 4634 368 4754 402
rect 4634 334 4677 368
rect 4711 334 4754 368
rect 4634 286 4754 334
rect 4810 436 4930 484
rect 4810 402 4855 436
rect 4889 402 4930 436
rect 4810 368 4930 402
rect 4810 334 4855 368
rect 4889 334 4930 368
rect 4810 286 4930 334
rect 5099 436 5219 484
rect 5099 402 5144 436
rect 5178 402 5219 436
rect 5099 368 5219 402
rect 5099 334 5144 368
rect 5178 334 5219 368
rect 5099 286 5219 334
rect 5275 436 5395 484
rect 5275 402 5315 436
rect 5349 402 5395 436
rect 5275 368 5395 402
rect 5275 334 5315 368
rect 5349 334 5395 368
rect 5275 286 5395 334
rect 5561 436 5681 484
rect 5561 402 5603 436
rect 5637 402 5681 436
rect 5561 368 5681 402
rect 5561 334 5603 368
rect 5637 334 5681 368
rect 5561 286 5681 334
rect 5847 436 5967 484
rect 5847 402 5893 436
rect 5927 402 5967 436
rect 5847 368 5967 402
rect 5847 334 5893 368
rect 5927 334 5967 368
rect 5847 286 5967 334
rect 6023 436 6143 484
rect 6023 402 6064 436
rect 6098 402 6143 436
rect 6023 368 6143 402
rect 6023 334 6064 368
rect 6098 334 6143 368
rect 6023 286 6143 334
rect 6309 436 6429 484
rect 6309 402 6353 436
rect 6387 402 6429 436
rect 6309 368 6429 402
rect 6309 334 6353 368
rect 6387 334 6429 368
rect 6309 286 6429 334
rect 6595 436 6715 484
rect 6595 402 6641 436
rect 6675 402 6715 436
rect 6595 368 6715 402
rect 6595 334 6641 368
rect 6675 334 6715 368
rect 6595 286 6715 334
rect 6771 436 6891 484
rect 6771 402 6812 436
rect 6846 402 6891 436
rect 6771 368 6891 402
rect 6771 334 6812 368
rect 6846 334 6891 368
rect 6771 286 6891 334
rect 161 120 281 146
rect 337 120 457 146
rect 623 120 743 146
rect 909 120 1029 146
rect 1085 120 1205 146
rect 1371 120 1491 146
rect 1547 120 1667 146
rect 1833 120 1953 146
rect 2670 120 2790 146
rect 2956 120 3076 146
rect 3132 120 3252 146
rect 3421 120 3541 146
rect 3707 120 3827 146
rect 3883 120 4003 146
rect 4172 120 4292 146
rect 4348 120 4468 146
rect 4634 120 4754 146
rect 4810 120 4930 146
rect 5099 120 5219 146
rect 5275 120 5395 146
rect 5561 120 5681 146
rect 5847 120 5967 146
rect 6023 120 6143 146
rect 6309 120 6429 146
rect 6595 120 6715 146
rect 6771 120 6891 146
<< polycont >>
rect 207 402 241 436
rect 207 334 241 368
rect 378 402 412 436
rect 378 334 412 368
rect 667 402 701 436
rect 667 334 701 368
rect 954 402 988 436
rect 954 334 988 368
rect 1125 402 1159 436
rect 1125 334 1159 368
rect 1417 402 1451 436
rect 1417 334 1451 368
rect 1588 402 1622 436
rect 1588 334 1622 368
rect 1877 402 1911 436
rect 1877 334 1911 368
rect 2714 402 2748 436
rect 2714 334 2748 368
rect 2999 402 3033 436
rect 2999 334 3033 368
rect 3177 402 3211 436
rect 3177 334 3211 368
rect 3465 402 3499 436
rect 3465 334 3499 368
rect 3750 402 3784 436
rect 3750 334 3784 368
rect 3928 402 3962 436
rect 3928 334 3962 368
rect 4217 402 4251 436
rect 4217 334 4251 368
rect 4388 402 4422 436
rect 4388 334 4422 368
rect 4677 402 4711 436
rect 4677 334 4711 368
rect 4855 402 4889 436
rect 4855 334 4889 368
rect 5144 402 5178 436
rect 5144 334 5178 368
rect 5315 402 5349 436
rect 5315 334 5349 368
rect 5603 402 5637 436
rect 5603 334 5637 368
rect 5893 402 5927 436
rect 5893 334 5927 368
rect 6064 402 6098 436
rect 6064 334 6098 368
rect 6353 402 6387 436
rect 6353 334 6387 368
rect 6641 402 6675 436
rect 6641 334 6675 368
rect 6812 402 6846 436
rect 6812 334 6846 368
<< locali >>
rect 67 1020 79 1054
rect 144 1020 152 1054
rect 212 1020 225 1054
rect 280 1020 298 1054
rect 348 1020 371 1054
rect 416 1020 444 1054
rect 484 1020 517 1054
rect 552 1020 586 1054
rect 624 1020 654 1054
rect 697 1020 722 1054
rect 770 1020 790 1054
rect 843 1020 858 1054
rect 916 1020 926 1054
rect 989 1020 994 1054
rect 1096 1020 1101 1054
rect 1164 1020 1173 1054
rect 1232 1020 1245 1054
rect 1300 1020 1317 1054
rect 1368 1020 1389 1054
rect 1436 1020 1461 1054
rect 1504 1020 1533 1054
rect 1572 1020 1605 1054
rect 1640 1020 1674 1054
rect 1711 1020 1742 1054
rect 1783 1020 1810 1054
rect 1855 1020 1878 1054
rect 1927 1020 1946 1054
rect 1999 1020 2014 1054
rect 2071 1020 2082 1054
rect 2143 1020 2150 1054
rect 2215 1020 2218 1054
rect 2252 1020 2253 1054
rect 2320 1020 2325 1054
rect 2388 1020 2397 1054
rect 2456 1020 2469 1054
rect 2524 1020 2541 1054
rect 2592 1020 2613 1054
rect 2660 1020 2685 1054
rect 2728 1020 2757 1054
rect 2796 1020 2829 1054
rect 2864 1020 2898 1054
rect 2935 1020 2966 1054
rect 3007 1020 3034 1054
rect 3079 1020 3102 1054
rect 3151 1020 3170 1054
rect 3223 1020 3238 1054
rect 3295 1020 3306 1054
rect 3367 1020 3374 1054
rect 3439 1020 3442 1054
rect 3476 1020 3477 1054
rect 3544 1020 3549 1054
rect 3612 1020 3621 1054
rect 3680 1020 3693 1054
rect 3748 1020 3765 1054
rect 3816 1020 3837 1054
rect 3884 1020 3909 1054
rect 3952 1020 3981 1054
rect 4020 1020 4053 1054
rect 4088 1020 4122 1054
rect 4159 1020 4190 1054
rect 4231 1020 4258 1054
rect 4303 1020 4326 1054
rect 4375 1020 4394 1054
rect 4447 1020 4462 1054
rect 4519 1020 4530 1054
rect 4591 1020 4598 1054
rect 4663 1020 4666 1054
rect 4700 1020 4701 1054
rect 4768 1020 4773 1054
rect 4836 1020 4845 1054
rect 4904 1020 4917 1054
rect 4972 1020 4989 1054
rect 5040 1020 5061 1054
rect 5108 1020 5133 1054
rect 5176 1020 5205 1054
rect 5244 1020 5277 1054
rect 5312 1020 5346 1054
rect 5383 1020 5414 1054
rect 5455 1020 5482 1054
rect 5527 1020 5550 1054
rect 5599 1020 5618 1054
rect 5671 1020 5686 1054
rect 5743 1020 5754 1054
rect 5815 1020 5822 1054
rect 5887 1020 5890 1054
rect 5924 1020 5925 1054
rect 5992 1020 5997 1054
rect 6060 1020 6069 1054
rect 6128 1020 6141 1054
rect 6196 1020 6213 1054
rect 6264 1020 6285 1054
rect 6332 1020 6357 1054
rect 6400 1020 6429 1054
rect 6468 1020 6501 1054
rect 6536 1020 6570 1054
rect 6607 1020 6638 1054
rect 6679 1020 6706 1054
rect 6751 1020 6774 1054
rect 6823 1020 6842 1054
rect 6895 1020 6910 1054
rect 6967 1020 6978 1054
rect 116 934 150 946
rect 116 866 150 874
rect 116 798 150 832
rect 116 672 150 764
rect 116 604 150 638
rect 116 536 150 570
rect 116 486 150 502
rect 292 934 326 952
rect 292 866 326 900
rect 292 798 326 832
rect 292 672 326 764
rect 292 604 326 638
rect 292 536 326 570
rect 173 402 207 436
rect 245 402 257 436
rect 191 368 257 402
rect 191 334 207 368
rect 241 334 257 368
rect 292 387 326 502
rect 468 934 502 946
rect 468 866 502 874
rect 468 798 502 832
rect 468 672 502 764
rect 468 604 502 638
rect 468 536 502 570
rect 468 486 502 502
rect 578 934 612 946
rect 578 866 612 874
rect 578 798 612 832
rect 578 672 612 764
rect 578 604 612 638
rect 578 536 612 570
rect 578 486 612 502
rect 754 934 788 952
rect 754 866 788 900
rect 754 798 788 832
rect 754 672 788 764
rect 754 604 788 638
rect 754 536 788 570
rect 754 436 788 502
rect 864 934 898 946
rect 864 866 898 874
rect 864 798 898 832
rect 864 672 898 764
rect 864 604 898 638
rect 864 536 898 570
rect 864 486 898 502
rect 1040 934 1074 952
rect 1040 866 1074 900
rect 1040 798 1074 832
rect 1040 672 1074 764
rect 1040 604 1074 638
rect 1040 536 1074 570
rect 292 315 326 353
rect 362 402 374 436
rect 412 402 446 436
rect 651 406 657 436
rect 651 402 667 406
rect 701 402 717 436
rect 362 368 428 402
rect 362 334 378 368
rect 412 334 428 368
rect 651 368 717 402
rect 651 334 657 368
rect 701 334 717 368
rect 754 402 954 436
rect 988 402 1004 436
rect 754 368 1004 402
rect 754 334 954 368
rect 988 334 1004 368
rect 1040 387 1074 502
rect 1216 934 1250 946
rect 1216 866 1250 874
rect 1216 798 1250 832
rect 1216 672 1250 764
rect 1216 604 1250 638
rect 1216 536 1250 570
rect 1216 486 1250 502
rect 1326 934 1360 946
rect 1326 866 1360 874
rect 1326 798 1360 832
rect 1326 672 1360 764
rect 1326 604 1360 638
rect 1326 536 1360 570
rect 1326 486 1360 502
rect 1502 934 1536 952
rect 1502 866 1536 900
rect 1502 798 1536 832
rect 1502 672 1536 764
rect 1502 604 1536 638
rect 1502 536 1536 570
rect 116 274 150 290
rect 116 229 150 240
rect 292 263 326 281
rect 468 274 502 290
rect 292 240 468 263
rect 292 229 502 240
rect 116 157 150 172
rect 463 206 502 229
rect 463 172 468 206
rect 463 156 502 172
rect 578 274 612 290
rect 578 229 612 240
rect 578 157 612 172
rect 754 274 788 334
rect 1040 315 1074 353
rect 1109 430 1125 436
rect 1159 430 1175 436
rect 1109 396 1121 430
rect 1159 402 1193 430
rect 1155 396 1193 402
rect 1401 406 1405 436
rect 1401 402 1417 406
rect 1451 402 1467 436
rect 1109 368 1175 396
rect 1109 334 1125 368
rect 1159 334 1175 368
rect 1401 368 1467 402
rect 1401 334 1405 368
rect 1451 334 1467 368
rect 1502 387 1536 502
rect 1678 934 1712 946
rect 1678 866 1712 874
rect 1678 798 1712 832
rect 1678 672 1712 764
rect 1678 604 1712 638
rect 1678 536 1712 570
rect 1678 486 1712 502
rect 1788 934 1822 946
rect 1788 866 1822 874
rect 1788 798 1822 832
rect 1788 672 1822 764
rect 1788 604 1822 638
rect 1788 536 1822 570
rect 1788 486 1822 502
rect 1964 934 1998 952
rect 1964 866 1998 900
rect 1964 798 1998 832
rect 1964 672 1998 764
rect 1964 604 1998 638
rect 1964 536 1998 570
rect 1964 448 1998 502
rect 2625 934 2659 946
rect 2625 866 2659 874
rect 2625 798 2659 832
rect 2625 672 2659 764
rect 2625 604 2659 638
rect 2625 536 2659 570
rect 2625 486 2659 502
rect 2801 934 2835 952
rect 2801 866 2835 900
rect 2801 798 2835 832
rect 2801 672 2835 764
rect 2801 604 2835 638
rect 2801 536 2835 570
rect 754 206 788 240
rect 754 156 788 172
rect 864 274 898 290
rect 1502 315 1536 353
rect 1572 402 1584 436
rect 1622 402 1656 436
rect 1861 406 1867 436
rect 1861 402 1877 406
rect 1911 402 1927 436
rect 1572 368 1638 402
rect 1572 334 1588 368
rect 1622 334 1638 368
rect 1861 368 1927 402
rect 1861 334 1867 368
rect 1911 334 1927 368
rect 1964 376 1998 414
rect 1040 263 1074 281
rect 898 240 1074 263
rect 864 229 1074 240
rect 1216 274 1250 290
rect 1216 229 1250 240
rect 864 206 903 229
rect 898 172 903 206
rect 864 156 903 172
rect 1216 157 1250 172
rect 1326 274 1360 290
rect 1326 229 1360 240
rect 1502 263 1536 281
rect 1678 274 1712 290
rect 1502 240 1678 263
rect 1502 229 1712 240
rect 1326 157 1360 172
rect 1673 206 1712 229
rect 1673 172 1678 206
rect 1673 156 1712 172
rect 1788 274 1822 290
rect 1788 229 1822 240
rect 1788 157 1822 172
rect 1964 274 1998 342
rect 2698 406 2706 436
rect 2698 402 2714 406
rect 2748 402 2764 436
rect 2698 368 2764 402
rect 2698 334 2706 368
rect 2748 334 2764 368
rect 2801 387 2835 502
rect 2911 934 2945 946
rect 2911 866 2945 874
rect 2911 798 2945 832
rect 2911 672 2945 764
rect 2911 604 2945 638
rect 2911 536 2945 570
rect 3087 934 3121 950
rect 3087 866 3121 900
rect 3087 798 3121 832
rect 3087 672 3121 764
rect 3087 604 3121 638
rect 3087 554 3121 570
rect 3263 934 3297 980
rect 3263 866 3297 900
rect 3263 798 3297 832
rect 3263 672 3297 764
rect 3263 604 3297 638
rect 3263 536 3297 570
rect 2911 486 2945 502
rect 3087 502 3263 520
rect 3087 486 3297 502
rect 3376 934 3410 946
rect 3376 866 3410 874
rect 3376 798 3410 832
rect 3376 672 3410 764
rect 3376 604 3410 638
rect 3376 536 3410 570
rect 3376 486 3410 502
rect 3552 934 3586 952
rect 3552 866 3586 900
rect 3552 798 3586 832
rect 3552 672 3586 764
rect 3552 604 3586 638
rect 3552 536 3586 570
rect 2801 315 2835 353
rect 2983 402 2999 406
rect 3033 402 3049 436
rect 2983 368 3049 402
rect 3033 334 3049 368
rect 3087 387 3121 486
rect 3552 440 3586 502
rect 3662 934 3696 946
rect 3662 866 3696 874
rect 3662 798 3696 832
rect 3662 672 3696 764
rect 3662 604 3696 638
rect 3662 536 3696 570
rect 3838 934 3872 950
rect 3838 866 3872 900
rect 3838 798 3872 832
rect 3838 672 3872 764
rect 3838 604 3872 638
rect 3838 554 3872 570
rect 4014 934 4048 980
rect 4014 866 4048 900
rect 4014 798 4048 832
rect 4014 672 4048 764
rect 4014 604 4048 638
rect 4014 536 4048 570
rect 3662 486 3696 502
rect 3838 502 4014 520
rect 3838 486 4048 502
rect 4127 934 4161 946
rect 4127 866 4161 874
rect 4127 798 4161 832
rect 4127 672 4161 764
rect 4127 604 4161 638
rect 4127 536 4161 570
rect 4127 486 4161 502
rect 4303 934 4337 952
rect 4303 866 4337 900
rect 4303 798 4337 832
rect 4303 672 4337 764
rect 4303 604 4337 638
rect 4303 536 4337 570
rect 1964 206 1998 240
rect 1964 156 1998 172
rect 2625 274 2659 290
rect 2625 229 2659 240
rect 2625 157 2659 172
rect 3087 315 3121 353
rect 3161 430 3177 436
rect 3211 430 3227 436
rect 3161 396 3173 430
rect 3211 402 3245 430
rect 3207 396 3245 402
rect 3448 402 3465 406
rect 3499 402 3515 436
rect 3161 368 3227 396
rect 3161 334 3177 368
rect 3211 334 3227 368
rect 3448 368 3515 402
rect 3499 334 3515 368
rect 3552 368 3586 406
rect 3734 402 3750 418
rect 3784 402 3800 436
rect 3734 380 3800 402
rect 3768 368 3800 380
rect 3734 334 3750 346
rect 3784 334 3800 368
rect 3838 387 3872 486
rect 4303 440 4337 502
rect 4479 934 4513 946
rect 4479 866 4513 874
rect 4479 798 4513 832
rect 4479 672 4513 764
rect 4479 604 4513 638
rect 4479 536 4513 570
rect 4479 486 4513 502
rect 4589 934 4623 946
rect 4589 866 4623 874
rect 4589 798 4623 832
rect 4589 672 4623 764
rect 4589 604 4623 638
rect 4589 536 4623 570
rect 4765 934 4799 950
rect 4765 866 4799 900
rect 4765 798 4799 832
rect 4765 672 4799 764
rect 4765 604 4799 638
rect 4765 554 4799 570
rect 4941 934 4975 980
rect 4941 866 4975 900
rect 4941 798 4975 832
rect 4941 672 4975 764
rect 4941 604 4975 638
rect 4941 536 4975 570
rect 4589 486 4623 502
rect 4765 502 4941 520
rect 4765 486 4975 502
rect 5054 934 5088 946
rect 5054 866 5088 874
rect 5054 798 5088 832
rect 5054 672 5088 764
rect 5054 604 5088 638
rect 5054 536 5088 570
rect 5054 486 5088 502
rect 5230 934 5264 952
rect 5230 866 5264 900
rect 5230 798 5264 832
rect 5230 672 5264 764
rect 5230 604 5264 638
rect 5230 536 5264 570
rect 2801 274 2835 281
rect 2801 206 2835 240
rect 2801 156 2835 172
rect 2911 274 2945 290
rect 2911 229 2945 240
rect 2911 157 2945 172
rect 3087 274 3121 281
rect 3087 206 3121 240
rect 3087 156 3121 172
rect 3263 274 3297 290
rect 3263 229 3297 240
rect 3263 157 3297 172
rect 3376 274 3410 290
rect 3376 229 3410 240
rect 3376 157 3410 172
rect 3552 274 3586 334
rect 3838 315 3872 353
rect 3912 405 3928 436
rect 3962 405 3978 436
rect 3912 371 3924 405
rect 3962 402 3996 405
rect 3958 371 3996 402
rect 4199 402 4217 406
rect 4251 402 4267 436
rect 3912 368 3978 371
rect 3912 334 3928 368
rect 3962 334 3978 368
rect 4199 368 4267 402
rect 4251 334 4267 368
rect 4303 368 4337 406
rect 4372 402 4388 436
rect 4424 406 4438 436
rect 4422 402 4438 406
rect 4372 368 4438 402
rect 4372 334 4388 368
rect 4424 334 4438 368
rect 4661 418 4667 436
rect 4661 402 4677 418
rect 4711 402 4727 436
rect 4661 380 4727 402
rect 4661 346 4667 380
rect 4701 368 4727 380
rect 4661 334 4677 346
rect 4711 334 4727 368
rect 4765 387 4799 486
rect 5230 440 5264 502
rect 5406 934 5440 946
rect 5406 866 5440 874
rect 5406 798 5440 832
rect 5406 672 5440 764
rect 5406 604 5440 638
rect 5406 536 5440 570
rect 5406 486 5440 502
rect 5516 934 5550 952
rect 5516 866 5550 900
rect 5516 798 5550 832
rect 5516 672 5550 764
rect 5516 604 5550 638
rect 5516 536 5550 570
rect 5516 501 5550 502
rect 5692 934 5726 946
rect 5692 866 5726 874
rect 5692 798 5726 832
rect 5692 672 5726 764
rect 5692 604 5726 638
rect 5692 536 5726 570
rect 5692 486 5726 502
rect 5802 934 5836 946
rect 5802 866 5836 874
rect 5802 798 5836 832
rect 5802 672 5836 764
rect 5802 604 5836 638
rect 5802 536 5836 570
rect 5802 486 5836 502
rect 5978 934 6012 952
rect 5978 866 6012 900
rect 5978 798 6012 832
rect 5978 672 6012 764
rect 5978 604 6012 638
rect 5978 536 6012 570
rect 3552 206 3586 240
rect 3552 156 3586 172
rect 3662 274 3696 290
rect 3662 229 3696 240
rect 3662 157 3696 172
rect 3838 274 3872 281
rect 3838 206 3872 240
rect 3838 156 3872 172
rect 4014 274 4048 290
rect 4014 229 4048 240
rect 4014 157 4048 172
rect 4127 274 4161 290
rect 4303 263 4337 334
rect 4765 315 4799 353
rect 4839 430 4855 436
rect 4889 430 4905 436
rect 4839 396 4851 430
rect 4889 402 4923 430
rect 4885 396 4923 402
rect 5128 402 5144 406
rect 5178 402 5194 436
rect 4839 368 4905 396
rect 4839 334 4855 368
rect 4889 334 4905 368
rect 5128 368 5194 402
rect 5178 334 5194 368
rect 5230 368 5264 406
rect 5299 406 5312 436
rect 5299 402 5315 406
rect 5349 402 5365 436
rect 5299 368 5365 402
rect 5299 334 5312 368
rect 5349 334 5365 368
rect 5516 429 5550 467
rect 4161 240 4337 263
rect 4127 229 4337 240
rect 4479 274 4513 290
rect 4479 229 4513 240
rect 4127 206 4166 229
rect 4161 172 4166 206
rect 4127 156 4166 172
rect 4479 157 4513 172
rect 4589 274 4623 290
rect 4589 229 4623 240
rect 4589 157 4623 172
rect 4765 274 4799 281
rect 4765 206 4799 240
rect 4765 156 4799 172
rect 4941 274 4975 290
rect 4941 229 4975 240
rect 4941 157 4975 172
rect 5054 274 5088 290
rect 5230 263 5264 334
rect 5088 240 5264 263
rect 5054 229 5264 240
rect 5406 274 5440 290
rect 5406 229 5440 240
rect 5054 206 5093 229
rect 5088 172 5093 206
rect 5054 156 5093 172
rect 5406 157 5440 172
rect 5516 274 5550 395
rect 5587 402 5603 436
rect 5647 418 5653 436
rect 5637 402 5653 418
rect 5587 380 5653 402
rect 5587 368 5613 380
rect 5587 334 5603 368
rect 5647 346 5653 380
rect 5637 334 5653 346
rect 5877 402 5893 436
rect 5927 402 5943 436
rect 5877 368 5943 402
rect 5877 334 5893 368
rect 5927 334 5943 368
rect 5978 387 6012 502
rect 6154 934 6188 946
rect 6154 866 6188 874
rect 6154 798 6188 832
rect 6154 672 6188 764
rect 6154 604 6188 638
rect 6154 536 6188 570
rect 6154 486 6188 502
rect 6264 934 6298 946
rect 6264 866 6298 874
rect 6264 798 6298 832
rect 6264 672 6298 764
rect 6264 604 6298 638
rect 6264 536 6298 570
rect 6264 486 6298 502
rect 6440 934 6474 952
rect 6440 866 6474 900
rect 6440 798 6474 832
rect 6440 672 6474 764
rect 6440 604 6474 638
rect 6440 536 6474 570
rect 6440 436 6474 502
rect 6550 934 6584 946
rect 6550 866 6584 874
rect 6550 798 6584 832
rect 6550 672 6584 764
rect 6550 604 6584 638
rect 6550 536 6584 570
rect 6550 486 6584 502
rect 6726 934 6760 952
rect 6726 866 6760 900
rect 6726 798 6760 832
rect 6726 672 6760 764
rect 6726 604 6760 638
rect 6726 536 6760 570
rect 6726 440 6760 502
rect 6902 934 6936 946
rect 6902 866 6936 874
rect 6902 798 6936 832
rect 6902 672 6936 764
rect 6902 604 6936 638
rect 6902 536 6936 570
rect 6902 486 6936 502
rect 5978 315 6012 353
rect 6048 402 6060 436
rect 6098 402 6132 436
rect 6336 402 6353 406
rect 6387 402 6403 436
rect 6048 368 6114 402
rect 6048 334 6064 368
rect 6098 334 6114 368
rect 6336 368 6403 402
rect 6387 334 6403 368
rect 6440 402 6641 436
rect 6675 402 6691 436
rect 6440 368 6691 402
rect 6440 334 6641 368
rect 6675 334 6691 368
rect 6726 368 6760 406
rect 6796 402 6812 436
rect 6846 402 6862 406
rect 6796 368 6862 402
rect 6796 334 6812 368
rect 5516 206 5550 240
rect 5516 156 5550 172
rect 5692 274 5726 290
rect 5692 229 5726 240
rect 5692 157 5726 172
rect 5802 274 5836 290
rect 5802 229 5836 240
rect 5978 263 6012 281
rect 6154 274 6188 290
rect 5978 240 6154 263
rect 5978 229 6188 240
rect 5802 157 5836 172
rect 6149 206 6188 229
rect 6149 172 6154 206
rect 6149 156 6188 172
rect 6264 274 6298 290
rect 6264 229 6298 240
rect 6264 157 6298 172
rect 6440 274 6474 334
rect 6440 206 6474 240
rect 6440 156 6474 172
rect 6550 274 6584 290
rect 6550 229 6584 240
rect 6726 263 6760 334
rect 6902 274 6936 290
rect 6726 240 6902 263
rect 6726 229 6936 240
rect 6550 157 6584 172
rect 6897 206 6936 229
rect 6897 172 6902 206
rect 6897 156 6936 172
rect 112 36 116 70
rect 150 36 151 70
rect 219 36 224 70
rect 288 36 297 70
rect 357 36 370 70
rect 426 36 443 70
rect 495 36 516 70
rect 564 36 589 70
rect 633 36 662 70
rect 702 36 735 70
rect 771 36 806 70
rect 842 36 875 70
rect 915 36 944 70
rect 988 36 1013 70
rect 1061 36 1082 70
rect 1134 36 1151 70
rect 1207 36 1220 70
rect 1279 36 1289 70
rect 1351 36 1358 70
rect 1423 36 1427 70
rect 1495 36 1496 70
rect 1530 36 1533 70
rect 1599 36 1605 70
rect 1668 36 1677 70
rect 1737 36 1749 70
rect 1806 36 1821 70
rect 1875 36 1893 70
rect 1944 36 1965 70
rect 2013 36 2037 70
rect 2082 36 2109 70
rect 2151 36 2181 70
rect 2220 36 2253 70
rect 2289 36 2324 70
rect 2359 36 2393 70
rect 2431 36 2462 70
rect 2503 36 2531 70
rect 2575 36 2600 70
rect 2647 36 2669 70
rect 2719 36 2738 70
rect 2791 36 2807 70
rect 2863 36 2876 70
rect 2935 36 2945 70
rect 3007 36 3014 70
rect 3079 36 3083 70
rect 3151 36 3152 70
rect 3186 36 3189 70
rect 3255 36 3261 70
rect 3324 36 3333 70
rect 3393 36 3405 70
rect 3461 36 3477 70
rect 3529 36 3549 70
rect 3597 36 3621 70
rect 3665 36 3693 70
rect 3733 36 3765 70
rect 3801 36 3835 70
rect 3871 36 3903 70
rect 3943 36 3971 70
rect 4015 36 4039 70
rect 4087 36 4107 70
rect 4159 36 4175 70
rect 4231 36 4243 70
rect 4303 36 4311 70
rect 4375 36 4379 70
rect 4481 36 4485 70
rect 4549 36 4557 70
rect 4617 36 4629 70
rect 4685 36 4701 70
rect 4753 36 4773 70
rect 4821 36 4845 70
rect 4889 36 4917 70
rect 4957 36 4989 70
rect 5025 36 5059 70
rect 5095 36 5127 70
rect 5167 36 5195 70
rect 5239 36 5263 70
rect 5311 36 5331 70
rect 5383 36 5399 70
rect 5455 36 5467 70
rect 5527 36 5535 70
rect 5599 36 5603 70
rect 5705 36 5709 70
rect 5773 36 5781 70
rect 5841 36 5853 70
rect 5909 36 5925 70
rect 5977 36 5997 70
rect 6045 36 6069 70
rect 6113 36 6141 70
rect 6181 36 6213 70
rect 6249 36 6283 70
rect 6319 36 6351 70
rect 6391 36 6419 70
rect 6463 36 6487 70
rect 6535 36 6555 70
rect 6607 36 6623 70
rect 6679 36 6691 70
rect 6751 36 6759 70
rect 6823 36 6827 70
rect 6929 36 6933 70
<< viali >>
rect 79 1020 110 1054
rect 110 1020 113 1054
rect 152 1020 178 1054
rect 178 1020 186 1054
rect 225 1020 246 1054
rect 246 1020 259 1054
rect 298 1020 314 1054
rect 314 1020 332 1054
rect 371 1020 382 1054
rect 382 1020 405 1054
rect 444 1020 450 1054
rect 450 1020 478 1054
rect 517 1020 518 1054
rect 518 1020 551 1054
rect 590 1020 620 1054
rect 620 1020 624 1054
rect 663 1020 688 1054
rect 688 1020 697 1054
rect 736 1020 756 1054
rect 756 1020 770 1054
rect 809 1020 824 1054
rect 824 1020 843 1054
rect 882 1020 892 1054
rect 892 1020 916 1054
rect 955 1020 960 1054
rect 960 1020 989 1054
rect 1028 1020 1062 1054
rect 1101 1020 1130 1054
rect 1130 1020 1135 1054
rect 1173 1020 1198 1054
rect 1198 1020 1207 1054
rect 1245 1020 1266 1054
rect 1266 1020 1279 1054
rect 1317 1020 1334 1054
rect 1334 1020 1351 1054
rect 1389 1020 1402 1054
rect 1402 1020 1423 1054
rect 1461 1020 1470 1054
rect 1470 1020 1495 1054
rect 1533 1020 1538 1054
rect 1538 1020 1567 1054
rect 1605 1020 1606 1054
rect 1606 1020 1639 1054
rect 1677 1020 1708 1054
rect 1708 1020 1711 1054
rect 1749 1020 1776 1054
rect 1776 1020 1783 1054
rect 1821 1020 1844 1054
rect 1844 1020 1855 1054
rect 1893 1020 1912 1054
rect 1912 1020 1927 1054
rect 1965 1020 1980 1054
rect 1980 1020 1999 1054
rect 2037 1020 2048 1054
rect 2048 1020 2071 1054
rect 2109 1020 2116 1054
rect 2116 1020 2143 1054
rect 2181 1020 2184 1054
rect 2184 1020 2215 1054
rect 2253 1020 2286 1054
rect 2286 1020 2287 1054
rect 2325 1020 2354 1054
rect 2354 1020 2359 1054
rect 2397 1020 2422 1054
rect 2422 1020 2431 1054
rect 2469 1020 2490 1054
rect 2490 1020 2503 1054
rect 2541 1020 2558 1054
rect 2558 1020 2575 1054
rect 2613 1020 2626 1054
rect 2626 1020 2647 1054
rect 2685 1020 2694 1054
rect 2694 1020 2719 1054
rect 2757 1020 2762 1054
rect 2762 1020 2791 1054
rect 2829 1020 2830 1054
rect 2830 1020 2863 1054
rect 2901 1020 2932 1054
rect 2932 1020 2935 1054
rect 2973 1020 3000 1054
rect 3000 1020 3007 1054
rect 3045 1020 3068 1054
rect 3068 1020 3079 1054
rect 3117 1020 3136 1054
rect 3136 1020 3151 1054
rect 3189 1020 3204 1054
rect 3204 1020 3223 1054
rect 3261 1020 3272 1054
rect 3272 1020 3295 1054
rect 3333 1020 3340 1054
rect 3340 1020 3367 1054
rect 3405 1020 3408 1054
rect 3408 1020 3439 1054
rect 3477 1020 3510 1054
rect 3510 1020 3511 1054
rect 3549 1020 3578 1054
rect 3578 1020 3583 1054
rect 3621 1020 3646 1054
rect 3646 1020 3655 1054
rect 3693 1020 3714 1054
rect 3714 1020 3727 1054
rect 3765 1020 3782 1054
rect 3782 1020 3799 1054
rect 3837 1020 3850 1054
rect 3850 1020 3871 1054
rect 3909 1020 3918 1054
rect 3918 1020 3943 1054
rect 3981 1020 3986 1054
rect 3986 1020 4015 1054
rect 4053 1020 4054 1054
rect 4054 1020 4087 1054
rect 4125 1020 4156 1054
rect 4156 1020 4159 1054
rect 4197 1020 4224 1054
rect 4224 1020 4231 1054
rect 4269 1020 4292 1054
rect 4292 1020 4303 1054
rect 4341 1020 4360 1054
rect 4360 1020 4375 1054
rect 4413 1020 4428 1054
rect 4428 1020 4447 1054
rect 4485 1020 4496 1054
rect 4496 1020 4519 1054
rect 4557 1020 4564 1054
rect 4564 1020 4591 1054
rect 4629 1020 4632 1054
rect 4632 1020 4663 1054
rect 4701 1020 4734 1054
rect 4734 1020 4735 1054
rect 4773 1020 4802 1054
rect 4802 1020 4807 1054
rect 4845 1020 4870 1054
rect 4870 1020 4879 1054
rect 4917 1020 4938 1054
rect 4938 1020 4951 1054
rect 4989 1020 5006 1054
rect 5006 1020 5023 1054
rect 5061 1020 5074 1054
rect 5074 1020 5095 1054
rect 5133 1020 5142 1054
rect 5142 1020 5167 1054
rect 5205 1020 5210 1054
rect 5210 1020 5239 1054
rect 5277 1020 5278 1054
rect 5278 1020 5311 1054
rect 5349 1020 5380 1054
rect 5380 1020 5383 1054
rect 5421 1020 5448 1054
rect 5448 1020 5455 1054
rect 5493 1020 5516 1054
rect 5516 1020 5527 1054
rect 5565 1020 5584 1054
rect 5584 1020 5599 1054
rect 5637 1020 5652 1054
rect 5652 1020 5671 1054
rect 5709 1020 5720 1054
rect 5720 1020 5743 1054
rect 5781 1020 5788 1054
rect 5788 1020 5815 1054
rect 5853 1020 5856 1054
rect 5856 1020 5887 1054
rect 5925 1020 5958 1054
rect 5958 1020 5959 1054
rect 5997 1020 6026 1054
rect 6026 1020 6031 1054
rect 6069 1020 6094 1054
rect 6094 1020 6103 1054
rect 6141 1020 6162 1054
rect 6162 1020 6175 1054
rect 6213 1020 6230 1054
rect 6230 1020 6247 1054
rect 6285 1020 6298 1054
rect 6298 1020 6319 1054
rect 6357 1020 6366 1054
rect 6366 1020 6391 1054
rect 6429 1020 6434 1054
rect 6434 1020 6463 1054
rect 6501 1020 6502 1054
rect 6502 1020 6535 1054
rect 6573 1020 6604 1054
rect 6604 1020 6607 1054
rect 6645 1020 6672 1054
rect 6672 1020 6679 1054
rect 6717 1020 6740 1054
rect 6740 1020 6751 1054
rect 6789 1020 6808 1054
rect 6808 1020 6823 1054
rect 6861 1020 6876 1054
rect 6876 1020 6895 1054
rect 6933 1020 6944 1054
rect 6944 1020 6967 1054
rect 116 946 150 980
rect 116 900 150 908
rect 116 874 150 900
rect 139 402 173 436
rect 211 402 241 436
rect 241 402 245 436
rect 468 946 502 980
rect 468 900 502 908
rect 468 874 502 900
rect 578 946 612 980
rect 578 900 612 908
rect 578 874 612 900
rect 657 436 691 440
rect 864 946 898 980
rect 864 900 898 908
rect 864 874 898 900
rect 292 353 326 387
rect 374 402 378 436
rect 378 402 408 436
rect 446 402 480 436
rect 657 406 667 436
rect 667 406 691 436
rect 657 334 667 368
rect 667 334 691 368
rect 1216 946 1250 980
rect 1216 900 1250 908
rect 1216 874 1250 900
rect 1326 946 1360 980
rect 1326 900 1360 908
rect 1326 874 1360 900
rect 1405 436 1439 440
rect 1040 353 1074 387
rect 292 281 326 315
rect 116 206 150 229
rect 116 195 150 206
rect 116 123 150 157
rect 578 206 612 229
rect 578 195 612 206
rect 578 123 612 157
rect 1121 402 1125 430
rect 1125 402 1155 430
rect 1121 396 1155 402
rect 1193 396 1227 430
rect 1405 406 1417 436
rect 1417 406 1439 436
rect 1405 334 1417 368
rect 1417 334 1439 368
rect 1678 946 1712 980
rect 1678 900 1712 908
rect 1678 874 1712 900
rect 1788 946 1822 980
rect 1788 900 1822 908
rect 1788 874 1822 900
rect 2625 946 2659 980
rect 2625 900 2659 908
rect 2625 874 2659 900
rect 1867 436 1901 440
rect 1502 353 1536 387
rect 1040 281 1074 315
rect 1584 402 1588 436
rect 1588 402 1618 436
rect 1656 402 1690 436
rect 1867 406 1877 436
rect 1877 406 1901 436
rect 1867 334 1877 368
rect 1877 334 1901 368
rect 1964 414 1998 448
rect 2706 436 2740 440
rect 1964 342 1998 376
rect 1216 206 1250 229
rect 1216 195 1250 206
rect 1216 123 1250 157
rect 1502 281 1536 315
rect 1326 206 1360 229
rect 1326 195 1360 206
rect 1326 123 1360 157
rect 1788 206 1822 229
rect 1788 195 1822 206
rect 1788 123 1822 157
rect 2706 406 2714 436
rect 2714 406 2740 436
rect 2706 334 2714 368
rect 2714 334 2740 368
rect 2911 946 2945 980
rect 2911 900 2945 908
rect 2911 874 2945 900
rect 3376 946 3410 980
rect 3376 900 3410 908
rect 3376 874 3410 900
rect 2801 353 2835 387
rect 2983 436 3017 440
rect 2983 406 2999 436
rect 2999 406 3017 436
rect 2983 334 2999 368
rect 2999 334 3017 368
rect 3662 946 3696 980
rect 3662 900 3696 908
rect 3662 874 3696 900
rect 4127 946 4161 980
rect 4127 900 4161 908
rect 4127 874 4161 900
rect 3448 436 3482 440
rect 3087 353 3121 387
rect 2625 206 2659 229
rect 2625 195 2659 206
rect 2625 123 2659 157
rect 2801 281 2835 315
rect 3173 402 3177 430
rect 3177 402 3207 430
rect 3173 396 3207 402
rect 3245 396 3279 430
rect 3448 406 3465 436
rect 3465 406 3482 436
rect 3448 334 3465 368
rect 3465 334 3482 368
rect 3552 406 3586 440
rect 3552 334 3586 368
rect 3734 436 3768 452
rect 3734 418 3750 436
rect 3750 418 3768 436
rect 3734 368 3768 380
rect 3734 346 3750 368
rect 3750 346 3768 368
rect 4479 946 4513 980
rect 4479 900 4513 908
rect 4479 874 4513 900
rect 4589 946 4623 980
rect 4589 900 4623 908
rect 4589 874 4623 900
rect 5054 946 5088 980
rect 5054 900 5088 908
rect 5054 874 5088 900
rect 4199 436 4233 440
rect 3838 353 3872 387
rect 2911 206 2945 229
rect 2911 195 2945 206
rect 2911 123 2945 157
rect 3087 281 3121 315
rect 3263 206 3297 229
rect 3263 195 3297 206
rect 3263 123 3297 157
rect 3376 206 3410 229
rect 3376 195 3410 206
rect 3376 123 3410 157
rect 4199 406 4217 436
rect 4217 406 4233 436
rect 3924 402 3928 405
rect 3928 402 3958 405
rect 3924 371 3958 402
rect 3996 371 4030 405
rect 4199 334 4217 368
rect 4217 334 4233 368
rect 4303 406 4337 440
rect 4390 436 4424 440
rect 4667 436 4701 452
rect 4303 334 4337 368
rect 4390 406 4422 436
rect 4422 406 4424 436
rect 4390 334 4422 368
rect 4422 334 4424 368
rect 4667 418 4677 436
rect 4677 418 4701 436
rect 4667 368 4701 380
rect 4667 346 4677 368
rect 4677 346 4701 368
rect 5406 946 5440 980
rect 5406 900 5440 908
rect 5406 874 5440 900
rect 5516 467 5550 501
rect 5692 946 5726 980
rect 5692 900 5726 908
rect 5692 874 5726 900
rect 5802 946 5836 980
rect 5802 900 5836 908
rect 5802 874 5836 900
rect 5128 436 5162 440
rect 4765 353 4799 387
rect 3662 206 3696 229
rect 3662 195 3696 206
rect 3662 123 3696 157
rect 3838 281 3872 315
rect 4014 206 4048 229
rect 4014 195 4048 206
rect 4014 123 4048 157
rect 4851 402 4855 430
rect 4855 402 4885 430
rect 4851 396 4885 402
rect 4923 396 4957 430
rect 5128 406 5144 436
rect 5144 406 5162 436
rect 5128 334 5144 368
rect 5144 334 5162 368
rect 5230 406 5264 440
rect 5312 436 5346 440
rect 5230 334 5264 368
rect 5312 406 5315 436
rect 5315 406 5346 436
rect 5312 334 5315 368
rect 5315 334 5346 368
rect 5613 436 5647 452
rect 5893 436 5927 440
rect 5516 395 5550 429
rect 4479 206 4513 229
rect 4479 195 4513 206
rect 4479 123 4513 157
rect 4589 206 4623 229
rect 4589 195 4623 206
rect 4589 123 4623 157
rect 4765 281 4799 315
rect 4941 206 4975 229
rect 4941 195 4975 206
rect 4941 123 4975 157
rect 5406 206 5440 229
rect 5406 195 5440 206
rect 5406 123 5440 157
rect 5613 418 5637 436
rect 5637 418 5647 436
rect 5613 368 5647 380
rect 5613 346 5637 368
rect 5637 346 5647 368
rect 5893 406 5927 436
rect 5893 334 5927 368
rect 6154 946 6188 980
rect 6154 900 6188 908
rect 6154 874 6188 900
rect 6264 946 6298 980
rect 6264 900 6298 908
rect 6264 874 6298 900
rect 6336 436 6370 440
rect 6550 946 6584 980
rect 6550 900 6584 908
rect 6550 874 6584 900
rect 6902 946 6936 980
rect 6902 900 6936 908
rect 6902 874 6936 900
rect 5978 353 6012 387
rect 6060 402 6064 436
rect 6064 402 6094 436
rect 6132 402 6166 436
rect 6336 406 6353 436
rect 6353 406 6370 436
rect 6336 334 6353 368
rect 6353 334 6370 368
rect 6726 406 6760 440
rect 6828 436 6862 440
rect 6726 334 6760 368
rect 6828 406 6846 436
rect 6846 406 6862 436
rect 6828 334 6846 368
rect 6846 334 6862 368
rect 5692 206 5726 229
rect 5692 195 5726 206
rect 5692 123 5726 157
rect 5978 281 6012 315
rect 5802 206 5836 229
rect 5802 195 5836 206
rect 5802 123 5836 157
rect 6264 206 6298 229
rect 6264 195 6298 206
rect 6264 123 6298 157
rect 6550 206 6584 229
rect 6550 195 6584 206
rect 6550 123 6584 157
rect 78 36 112 70
rect 151 36 185 70
rect 224 36 254 70
rect 254 36 258 70
rect 297 36 323 70
rect 323 36 331 70
rect 370 36 392 70
rect 392 36 404 70
rect 443 36 461 70
rect 461 36 477 70
rect 516 36 530 70
rect 530 36 550 70
rect 589 36 599 70
rect 599 36 623 70
rect 662 36 668 70
rect 668 36 696 70
rect 735 36 737 70
rect 737 36 769 70
rect 808 36 840 70
rect 840 36 842 70
rect 881 36 909 70
rect 909 36 915 70
rect 954 36 978 70
rect 978 36 988 70
rect 1027 36 1047 70
rect 1047 36 1061 70
rect 1100 36 1116 70
rect 1116 36 1134 70
rect 1173 36 1185 70
rect 1185 36 1207 70
rect 1245 36 1254 70
rect 1254 36 1279 70
rect 1317 36 1323 70
rect 1323 36 1351 70
rect 1389 36 1392 70
rect 1392 36 1423 70
rect 1461 36 1495 70
rect 1533 36 1565 70
rect 1565 36 1567 70
rect 1605 36 1634 70
rect 1634 36 1639 70
rect 1677 36 1703 70
rect 1703 36 1711 70
rect 1749 36 1772 70
rect 1772 36 1783 70
rect 1821 36 1841 70
rect 1841 36 1855 70
rect 1893 36 1910 70
rect 1910 36 1927 70
rect 1965 36 1979 70
rect 1979 36 1999 70
rect 2037 36 2048 70
rect 2048 36 2071 70
rect 2109 36 2117 70
rect 2117 36 2143 70
rect 2181 36 2186 70
rect 2186 36 2215 70
rect 2253 36 2255 70
rect 2255 36 2287 70
rect 2325 36 2358 70
rect 2358 36 2359 70
rect 2397 36 2427 70
rect 2427 36 2431 70
rect 2469 36 2496 70
rect 2496 36 2503 70
rect 2541 36 2565 70
rect 2565 36 2575 70
rect 2613 36 2634 70
rect 2634 36 2647 70
rect 2685 36 2703 70
rect 2703 36 2719 70
rect 2757 36 2772 70
rect 2772 36 2791 70
rect 2829 36 2841 70
rect 2841 36 2863 70
rect 2901 36 2910 70
rect 2910 36 2935 70
rect 2973 36 2979 70
rect 2979 36 3007 70
rect 3045 36 3048 70
rect 3048 36 3079 70
rect 3117 36 3151 70
rect 3189 36 3221 70
rect 3221 36 3223 70
rect 3261 36 3290 70
rect 3290 36 3295 70
rect 3333 36 3359 70
rect 3359 36 3367 70
rect 3405 36 3427 70
rect 3427 36 3439 70
rect 3477 36 3495 70
rect 3495 36 3511 70
rect 3549 36 3563 70
rect 3563 36 3583 70
rect 3621 36 3631 70
rect 3631 36 3655 70
rect 3693 36 3699 70
rect 3699 36 3727 70
rect 3765 36 3767 70
rect 3767 36 3799 70
rect 3837 36 3869 70
rect 3869 36 3871 70
rect 3909 36 3937 70
rect 3937 36 3943 70
rect 3981 36 4005 70
rect 4005 36 4015 70
rect 4053 36 4073 70
rect 4073 36 4087 70
rect 4125 36 4141 70
rect 4141 36 4159 70
rect 4197 36 4209 70
rect 4209 36 4231 70
rect 4269 36 4277 70
rect 4277 36 4303 70
rect 4341 36 4345 70
rect 4345 36 4375 70
rect 4413 36 4447 70
rect 4485 36 4515 70
rect 4515 36 4519 70
rect 4557 36 4583 70
rect 4583 36 4591 70
rect 4629 36 4651 70
rect 4651 36 4663 70
rect 4701 36 4719 70
rect 4719 36 4735 70
rect 4773 36 4787 70
rect 4787 36 4807 70
rect 4845 36 4855 70
rect 4855 36 4879 70
rect 4917 36 4923 70
rect 4923 36 4951 70
rect 4989 36 4991 70
rect 4991 36 5023 70
rect 5061 36 5093 70
rect 5093 36 5095 70
rect 5133 36 5161 70
rect 5161 36 5167 70
rect 5205 36 5229 70
rect 5229 36 5239 70
rect 5277 36 5297 70
rect 5297 36 5311 70
rect 5349 36 5365 70
rect 5365 36 5383 70
rect 5421 36 5433 70
rect 5433 36 5455 70
rect 5493 36 5501 70
rect 5501 36 5527 70
rect 5565 36 5569 70
rect 5569 36 5599 70
rect 5637 36 5671 70
rect 5709 36 5739 70
rect 5739 36 5743 70
rect 5781 36 5807 70
rect 5807 36 5815 70
rect 5853 36 5875 70
rect 5875 36 5887 70
rect 5925 36 5943 70
rect 5943 36 5959 70
rect 5997 36 6011 70
rect 6011 36 6031 70
rect 6069 36 6079 70
rect 6079 36 6103 70
rect 6141 36 6147 70
rect 6147 36 6175 70
rect 6213 36 6215 70
rect 6215 36 6247 70
rect 6285 36 6317 70
rect 6317 36 6319 70
rect 6357 36 6385 70
rect 6385 36 6391 70
rect 6429 36 6453 70
rect 6453 36 6463 70
rect 6501 36 6521 70
rect 6521 36 6535 70
rect 6573 36 6589 70
rect 6589 36 6607 70
rect 6645 36 6657 70
rect 6657 36 6679 70
rect 6717 36 6725 70
rect 6725 36 6751 70
rect 6789 36 6793 70
rect 6793 36 6823 70
rect 6861 36 6895 70
rect 6933 36 6967 70
<< metal1 >>
rect 67 1054 6979 1064
rect 67 1020 79 1054
rect 113 1020 152 1054
rect 186 1020 225 1054
rect 259 1020 298 1054
rect 332 1020 371 1054
rect 405 1020 444 1054
rect 478 1020 517 1054
rect 551 1020 590 1054
rect 624 1020 663 1054
rect 697 1020 736 1054
rect 770 1020 809 1054
rect 843 1020 882 1054
rect 916 1020 955 1054
rect 989 1020 1028 1054
rect 1062 1020 1101 1054
rect 1135 1020 1173 1054
rect 1207 1020 1245 1054
rect 1279 1020 1317 1054
rect 1351 1020 1389 1054
rect 1423 1020 1461 1054
rect 1495 1020 1533 1054
rect 1567 1020 1605 1054
rect 1639 1020 1677 1054
rect 1711 1020 1749 1054
rect 1783 1020 1821 1054
rect 1855 1020 1893 1054
rect 1927 1020 1965 1054
rect 1999 1020 2037 1054
rect 2071 1020 2109 1054
rect 2143 1020 2181 1054
rect 2215 1020 2253 1054
rect 2287 1020 2325 1054
rect 2359 1020 2397 1054
rect 2431 1020 2469 1054
rect 2503 1020 2541 1054
rect 2575 1020 2613 1054
rect 2647 1020 2685 1054
rect 2719 1020 2757 1054
rect 2791 1020 2829 1054
rect 2863 1020 2901 1054
rect 2935 1020 2973 1054
rect 3007 1020 3045 1054
rect 3079 1020 3117 1054
rect 3151 1020 3189 1054
rect 3223 1020 3261 1054
rect 3295 1020 3333 1054
rect 3367 1020 3405 1054
rect 3439 1020 3477 1054
rect 3511 1020 3549 1054
rect 3583 1020 3621 1054
rect 3655 1020 3693 1054
rect 3727 1020 3765 1054
rect 3799 1020 3837 1054
rect 3871 1020 3909 1054
rect 3943 1020 3981 1054
rect 4015 1020 4053 1054
rect 4087 1020 4125 1054
rect 4159 1020 4197 1054
rect 4231 1020 4269 1054
rect 4303 1020 4341 1054
rect 4375 1020 4413 1054
rect 4447 1020 4485 1054
rect 4519 1020 4557 1054
rect 4591 1020 4629 1054
rect 4663 1020 4701 1054
rect 4735 1020 4773 1054
rect 4807 1020 4845 1054
rect 4879 1020 4917 1054
rect 4951 1020 4989 1054
rect 5023 1020 5061 1054
rect 5095 1020 5133 1054
rect 5167 1020 5205 1054
rect 5239 1020 5277 1054
rect 5311 1020 5349 1054
rect 5383 1020 5421 1054
rect 5455 1020 5493 1054
rect 5527 1020 5565 1054
rect 5599 1020 5637 1054
rect 5671 1020 5709 1054
rect 5743 1020 5781 1054
rect 5815 1020 5853 1054
rect 5887 1020 5925 1054
rect 5959 1020 5997 1054
rect 6031 1020 6069 1054
rect 6103 1020 6141 1054
rect 6175 1020 6213 1054
rect 6247 1020 6285 1054
rect 6319 1020 6357 1054
rect 6391 1020 6429 1054
rect 6463 1020 6501 1054
rect 6535 1020 6573 1054
rect 6607 1020 6645 1054
rect 6679 1020 6717 1054
rect 6751 1020 6789 1054
rect 6823 1020 6861 1054
rect 6895 1020 6933 1054
rect 6967 1020 6979 1054
rect 67 980 6979 1020
rect 67 946 116 980
rect 150 946 468 980
rect 502 946 578 980
rect 612 946 864 980
rect 898 946 1216 980
rect 1250 946 1326 980
rect 1360 946 1678 980
rect 1712 946 1788 980
rect 1822 946 2625 980
rect 2659 946 2911 980
rect 2945 946 3376 980
rect 3410 946 3662 980
rect 3696 946 4127 980
rect 4161 946 4479 980
rect 4513 946 4589 980
rect 4623 946 5054 980
rect 5088 946 5406 980
rect 5440 946 5692 980
rect 5726 946 5802 980
rect 5836 946 6154 980
rect 6188 946 6264 980
rect 6298 946 6550 980
rect 6584 946 6902 980
rect 6936 946 6979 980
rect 67 908 6979 946
rect 67 874 116 908
rect 150 874 468 908
rect 502 874 578 908
rect 612 874 864 908
rect 898 874 1216 908
rect 1250 874 1326 908
rect 1360 874 1678 908
rect 1712 874 1788 908
rect 1822 874 2625 908
rect 2659 874 2911 908
rect 2945 874 3376 908
rect 3410 874 3662 908
rect 3696 874 4127 908
rect 4161 874 4479 908
rect 4513 874 4589 908
rect 4623 874 5054 908
rect 5088 874 5406 908
rect 5440 874 5692 908
rect 5726 874 5802 908
rect 5836 874 6154 908
rect 6188 874 6264 908
rect 6298 874 6550 908
rect 6584 874 6902 908
rect 6936 874 6979 908
rect 67 861 6979 874
rect 1958 701 4508 753
tri 4508 701 4514 707 sw
rect 4658 701 4664 753
rect 4716 701 4728 753
rect 4780 701 5583 753
rect 1958 673 2010 701
tri 2010 673 2038 701 nw
tri 4399 673 4427 701 ne
rect 4427 673 4514 701
tri 4514 673 4542 701 sw
rect 127 436 257 442
rect 127 402 139 436
rect 173 402 211 436
rect 245 402 257 436
rect 127 396 257 402
rect 362 436 492 442
rect 362 402 374 436
rect 408 402 446 436
rect 480 402 492 436
rect 286 387 332 399
rect 362 396 492 402
rect 651 440 697 452
rect 651 406 657 440
rect 691 406 697 440
rect 1399 440 1445 452
rect 1861 451 1907 452
rect 286 353 292 387
rect 326 353 332 387
rect 651 368 697 406
rect 1109 430 1239 436
rect 286 334 332 353
tri 332 334 353 355 sw
tri 630 334 651 355 se
rect 651 334 657 368
rect 691 334 697 368
rect 286 321 353 334
tri 353 321 366 334 sw
tri 617 321 630 334 se
rect 630 321 697 334
rect 286 315 697 321
rect 286 281 292 315
rect 326 281 697 315
rect 286 269 697 281
rect 1034 387 1080 399
rect 1109 396 1121 430
rect 1155 396 1193 430
rect 1227 396 1239 430
rect 1109 390 1239 396
rect 1399 406 1405 440
rect 1439 406 1445 440
rect 1034 353 1040 387
rect 1074 353 1080 387
rect 1399 368 1445 406
rect 1572 436 1702 442
rect 1572 402 1584 436
rect 1618 402 1656 436
rect 1690 402 1702 436
rect 1034 334 1080 353
tri 1080 334 1101 355 sw
tri 1378 334 1399 355 se
rect 1399 334 1405 368
rect 1439 334 1445 368
rect 1034 321 1101 334
tri 1101 321 1114 334 sw
tri 1365 321 1378 334 se
rect 1378 321 1445 334
rect 1034 315 1445 321
rect 1034 281 1040 315
rect 1074 281 1445 315
rect 1034 269 1445 281
rect 1496 387 1542 399
rect 1572 396 1702 402
rect 1861 440 1913 451
rect 1861 406 1867 440
rect 1901 406 1913 440
rect 1496 353 1502 387
rect 1536 353 1542 387
rect 1861 368 1913 406
rect 1496 334 1542 353
tri 1542 334 1563 355 sw
tri 1840 334 1861 355 se
rect 1861 334 1867 368
rect 1901 334 1913 368
rect 1496 322 1563 334
tri 1563 322 1575 334 sw
tri 1828 322 1840 334 se
rect 1840 322 1913 334
rect 1958 448 2004 673
tri 2004 667 2010 673 nw
rect 3161 621 4224 673
rect 4276 621 4288 673
rect 4340 621 4346 673
tri 4427 667 4433 673 ne
rect 4433 621 4439 673
rect 4491 621 4503 673
rect 4555 621 5309 673
rect 5361 621 5373 673
rect 5425 621 5856 673
rect 5908 621 5920 673
rect 5972 621 5978 673
rect 3161 593 3233 621
tri 3233 593 3261 621 nw
rect 3161 467 3227 593
tri 3227 587 3233 593 nw
rect 3912 541 3918 593
rect 3970 541 3982 593
rect 4034 569 4040 593
tri 4040 569 4064 593 sw
rect 4034 541 5653 569
tri 5573 513 5601 541 ne
rect 5601 513 5653 541
rect 3728 485 4710 513
tri 5041 501 5053 513 se
rect 5053 501 5556 513
tri 5601 507 5607 513 ne
tri 5025 485 5041 501 se
rect 5041 485 5516 501
tri 3227 467 3230 470 sw
rect 3728 467 3790 485
tri 3790 467 3808 485 nw
tri 4624 467 4642 485 ne
rect 4642 467 4710 485
tri 5007 467 5025 485 se
rect 5025 467 5070 485
tri 5070 467 5088 485 nw
tri 5476 467 5494 485 ne
rect 5494 467 5516 485
rect 5550 467 5556 501
rect 3161 452 3230 467
tri 3230 452 3245 467 sw
rect 3728 452 3775 467
tri 3775 452 3790 467 nw
tri 4642 452 4657 467 ne
rect 4657 456 4710 467
tri 5000 460 5007 467 se
rect 5007 460 5063 467
tri 5063 460 5070 467 nw
tri 5494 460 5501 467 ne
rect 5501 460 5556 467
rect 4657 452 4658 456
tri 4992 452 5000 460 se
rect 5000 452 5055 460
tri 5055 452 5063 460 nw
tri 5501 452 5509 460 ne
rect 5509 452 5556 460
rect 1958 414 1964 448
rect 1998 414 2004 448
rect 1958 376 2004 414
rect 1958 342 1964 376
rect 1998 342 2004 376
rect 1958 330 2004 342
rect 2700 440 2746 452
rect 2700 406 2706 440
rect 2740 406 2746 440
rect 2700 368 2746 406
rect 2977 440 3023 452
rect 2977 406 2983 440
rect 3017 406 3023 440
rect 2700 334 2706 368
rect 2740 334 2746 368
rect 1496 321 1575 322
tri 1575 321 1576 322 sw
tri 1827 321 1828 322 se
rect 1828 321 1913 322
rect 1496 315 1913 321
rect 1496 281 1502 315
rect 1536 281 1913 315
rect 2700 306 2746 334
rect 2795 387 2841 399
rect 2795 353 2801 387
rect 2835 353 2841 387
rect 2977 368 3023 406
rect 3161 440 3245 452
tri 3245 440 3257 452 sw
rect 3442 440 3488 452
rect 3161 436 3257 440
tri 3257 436 3261 440 sw
rect 3161 430 3291 436
rect 2795 334 2841 353
tri 2841 334 2862 355 sw
tri 2956 334 2977 355 se
rect 2977 334 2983 368
rect 3017 334 3023 368
rect 2795 321 2862 334
tri 2862 321 2875 334 sw
tri 2943 321 2956 334 se
rect 2956 321 3023 334
rect 2795 315 3023 321
rect 1496 269 1913 281
rect 2795 281 2801 315
rect 2835 281 3023 315
rect 2795 269 3023 281
rect 3081 387 3127 399
rect 3161 396 3173 430
rect 3207 396 3245 430
rect 3279 396 3291 430
rect 3161 390 3291 396
rect 3442 406 3448 440
rect 3482 406 3488 440
rect 3081 353 3087 387
rect 3121 353 3127 387
rect 3442 368 3488 406
rect 3081 334 3127 353
tri 3127 334 3148 355 sw
tri 3421 334 3442 355 se
rect 3442 334 3448 368
rect 3482 334 3488 368
rect 3081 321 3148 334
tri 3148 321 3161 334 sw
tri 3408 321 3421 334 se
rect 3421 321 3488 334
rect 3546 440 3592 452
rect 3546 406 3552 440
rect 3586 406 3592 440
rect 3546 368 3592 406
rect 3546 334 3552 368
rect 3586 334 3592 368
rect 3728 418 3734 452
rect 3768 418 3774 452
tri 3774 451 3775 452 nw
rect 3728 380 3774 418
rect 4193 440 4239 452
rect 3728 346 3734 380
rect 3768 346 3774 380
rect 3728 334 3774 346
rect 3832 387 3878 399
rect 3832 353 3838 387
rect 3872 353 3878 387
rect 3912 362 3918 414
rect 3970 362 3982 414
rect 4034 362 4042 414
rect 4193 406 4199 440
rect 4233 406 4239 440
rect 4193 368 4239 406
rect 3832 334 3878 353
tri 3878 334 3899 355 sw
tri 4172 334 4193 355 se
rect 4193 334 4199 368
rect 4233 334 4239 368
rect 3546 322 3592 334
rect 3081 315 3488 321
rect 3081 281 3087 315
rect 3121 281 3488 315
rect 3081 269 3488 281
rect 3832 321 3899 334
tri 3899 321 3912 334 sw
tri 4159 321 4172 334 se
rect 4172 321 4239 334
rect 4294 445 4346 452
rect 4294 381 4346 393
rect 4294 322 4346 329
rect 4381 444 4433 452
tri 4657 451 4658 452 ne
rect 4381 380 4433 392
tri 4990 450 4992 452 se
rect 4992 450 5053 452
tri 5053 450 5055 452 nw
tri 4980 440 4990 450 se
rect 4990 440 5043 450
tri 5043 440 5053 450 nw
rect 5122 440 5168 452
tri 4976 436 4980 440 se
rect 4980 436 5039 440
tri 5039 436 5043 440 nw
rect 4658 392 4710 404
rect 4839 430 5009 436
rect 4658 334 4710 340
rect 4759 387 4805 399
rect 4839 396 4851 430
rect 4885 396 4923 430
rect 4957 406 5009 430
tri 5009 406 5039 436 nw
rect 5122 406 5128 440
rect 5162 406 5168 440
rect 4957 396 4998 406
rect 4839 395 4998 396
tri 4998 395 5009 406 nw
rect 4839 390 4993 395
tri 4993 390 4998 395 nw
rect 4759 353 4765 387
rect 4799 353 4805 387
rect 5122 368 5168 406
rect 4759 334 4805 353
tri 4805 334 4826 355 sw
tri 5101 334 5122 355 se
rect 5122 334 5128 368
rect 5162 334 5168 368
rect 4381 322 4433 328
rect 4759 330 4826 334
tri 4826 330 4830 334 sw
tri 5097 330 5101 334 se
rect 5101 330 5168 334
rect 4759 322 4830 330
tri 4830 322 4838 330 sw
tri 5089 322 5097 330 se
rect 5097 322 5168 330
rect 5221 444 5273 452
rect 5221 380 5273 392
rect 5221 322 5273 328
rect 5303 444 5355 452
tri 5509 451 5510 452 ne
rect 5303 380 5355 392
rect 5510 429 5556 452
rect 5510 395 5516 429
rect 5550 395 5556 429
rect 5510 383 5556 395
rect 5607 462 5653 513
tri 5653 462 5659 468 sw
rect 5607 456 5659 462
rect 5607 392 5659 404
rect 5607 334 5659 340
rect 5884 444 5936 452
rect 6050 442 6056 445
rect 5884 380 5936 392
rect 5303 322 5355 328
rect 5884 322 5936 328
rect 5972 387 6018 399
rect 6048 396 6056 442
rect 6050 393 6056 396
rect 6108 393 6120 445
rect 6172 393 6178 445
rect 6330 440 6376 452
rect 6330 406 6336 440
rect 6370 406 6376 440
rect 5972 353 5978 387
rect 6012 353 6018 387
rect 6330 368 6376 406
rect 5972 334 6018 353
tri 6018 334 6039 355 sw
tri 6309 334 6330 355 se
rect 6330 334 6336 368
rect 6370 334 6376 368
rect 3832 315 4239 321
rect 3832 281 3838 315
rect 3872 281 4239 315
rect 3832 269 4239 281
rect 4759 321 4838 322
tri 4838 321 4839 322 sw
tri 5088 321 5089 322 se
rect 5089 321 5168 322
rect 4759 315 5168 321
rect 4759 281 4765 315
rect 4799 281 5168 315
rect 4759 269 5168 281
rect 5972 321 6039 334
tri 6039 321 6052 334 sw
tri 6296 321 6309 334 se
rect 6309 321 6376 334
rect 6720 440 6766 452
rect 6720 406 6726 440
rect 6760 406 6766 440
rect 6720 368 6766 406
rect 6720 334 6726 368
rect 6760 334 6766 368
rect 6720 322 6766 334
rect 6822 440 6868 452
rect 6822 406 6828 440
rect 6862 406 6868 440
rect 6822 368 6868 406
rect 6822 334 6828 368
rect 6862 334 6868 368
rect 6822 322 6868 334
rect 5972 315 6376 321
rect 5972 281 5978 315
rect 6012 281 6376 315
rect 5972 269 6376 281
rect 66 229 6979 241
rect 66 195 116 229
rect 150 195 578 229
rect 612 195 1216 229
rect 1250 195 1326 229
rect 1360 195 1788 229
rect 1822 195 2625 229
rect 2659 195 2911 229
rect 2945 195 3263 229
rect 3297 195 3376 229
rect 3410 195 3662 229
rect 3696 195 4014 229
rect 4048 195 4479 229
rect 4513 195 4589 229
rect 4623 195 4941 229
rect 4975 195 5406 229
rect 5440 195 5692 229
rect 5726 195 5802 229
rect 5836 195 6264 229
rect 6298 195 6550 229
rect 6584 195 6979 229
rect 66 157 6979 195
rect 66 123 116 157
rect 150 123 578 157
rect 612 123 1216 157
rect 1250 123 1326 157
rect 1360 123 1788 157
rect 1822 123 2625 157
rect 2659 123 2911 157
rect 2945 123 3263 157
rect 3297 123 3376 157
rect 3410 123 3662 157
rect 3696 123 4014 157
rect 4048 123 4479 157
rect 4513 123 4589 157
rect 4623 123 4941 157
rect 4975 123 5406 157
rect 5440 123 5692 157
rect 5726 123 5802 157
rect 5836 123 6264 157
rect 6298 123 6550 157
rect 6584 123 6979 157
rect 66 70 6979 123
rect 66 36 78 70
rect 112 36 151 70
rect 185 36 224 70
rect 258 36 297 70
rect 331 36 370 70
rect 404 36 443 70
rect 477 36 516 70
rect 550 36 589 70
rect 623 36 662 70
rect 696 36 735 70
rect 769 36 808 70
rect 842 36 881 70
rect 915 36 954 70
rect 988 36 1027 70
rect 1061 36 1100 70
rect 1134 36 1173 70
rect 1207 36 1245 70
rect 1279 36 1317 70
rect 1351 36 1389 70
rect 1423 36 1461 70
rect 1495 36 1533 70
rect 1567 36 1605 70
rect 1639 36 1677 70
rect 1711 36 1749 70
rect 1783 36 1821 70
rect 1855 36 1893 70
rect 1927 36 1965 70
rect 1999 36 2037 70
rect 2071 36 2109 70
rect 2143 36 2181 70
rect 2215 36 2253 70
rect 2287 36 2325 70
rect 2359 36 2397 70
rect 2431 36 2469 70
rect 2503 36 2541 70
rect 2575 36 2613 70
rect 2647 36 2685 70
rect 2719 36 2757 70
rect 2791 36 2829 70
rect 2863 36 2901 70
rect 2935 36 2973 70
rect 3007 36 3045 70
rect 3079 36 3117 70
rect 3151 36 3189 70
rect 3223 36 3261 70
rect 3295 36 3333 70
rect 3367 36 3405 70
rect 3439 36 3477 70
rect 3511 36 3549 70
rect 3583 36 3621 70
rect 3655 36 3693 70
rect 3727 36 3765 70
rect 3799 36 3837 70
rect 3871 36 3909 70
rect 3943 36 3981 70
rect 4015 36 4053 70
rect 4087 36 4125 70
rect 4159 36 4197 70
rect 4231 36 4269 70
rect 4303 36 4341 70
rect 4375 36 4413 70
rect 4447 36 4485 70
rect 4519 36 4557 70
rect 4591 36 4629 70
rect 4663 36 4701 70
rect 4735 36 4773 70
rect 4807 36 4845 70
rect 4879 36 4917 70
rect 4951 36 4989 70
rect 5023 36 5061 70
rect 5095 36 5133 70
rect 5167 36 5205 70
rect 5239 36 5277 70
rect 5311 36 5349 70
rect 5383 36 5421 70
rect 5455 36 5493 70
rect 5527 36 5565 70
rect 5599 36 5637 70
rect 5671 36 5709 70
rect 5743 36 5781 70
rect 5815 36 5853 70
rect 5887 36 5925 70
rect 5959 36 5997 70
rect 6031 36 6069 70
rect 6103 36 6141 70
rect 6175 36 6213 70
rect 6247 36 6285 70
rect 6319 36 6357 70
rect 6391 36 6429 70
rect 6463 36 6501 70
rect 6535 36 6573 70
rect 6607 36 6645 70
rect 6679 36 6717 70
rect 6751 36 6789 70
rect 6823 36 6861 70
rect 6895 36 6933 70
rect 6967 36 6979 70
rect 66 26 6979 36
rect 6048 -134 6054 -82
rect 6106 -134 6118 -82
rect 6170 -134 6176 -82
<< via1 >>
rect 4664 701 4716 753
rect 4728 701 4780 753
rect 4224 621 4276 673
rect 4288 621 4340 673
rect 4439 621 4491 673
rect 4503 621 4555 673
rect 5309 621 5361 673
rect 5373 621 5425 673
rect 5856 621 5908 673
rect 5920 621 5972 673
rect 3918 541 3970 593
rect 3982 541 4034 593
rect 4658 452 4710 456
rect 3918 405 3970 414
rect 3918 371 3924 405
rect 3924 371 3958 405
rect 3958 371 3970 405
rect 3918 362 3970 371
rect 3982 405 4034 414
rect 3982 371 3996 405
rect 3996 371 4030 405
rect 4030 371 4034 405
rect 3982 362 4034 371
rect 4294 440 4346 445
rect 4294 406 4303 440
rect 4303 406 4337 440
rect 4337 406 4346 440
rect 4294 393 4346 406
rect 4294 368 4346 381
rect 4294 334 4303 368
rect 4303 334 4337 368
rect 4337 334 4346 368
rect 4294 329 4346 334
rect 4381 440 4433 444
rect 4381 406 4390 440
rect 4390 406 4424 440
rect 4424 406 4433 440
rect 4381 392 4433 406
rect 4381 368 4433 380
rect 4381 334 4390 368
rect 4390 334 4424 368
rect 4424 334 4433 368
rect 4658 418 4667 452
rect 4667 418 4701 452
rect 4701 418 4710 452
rect 4658 404 4710 418
rect 4658 380 4710 392
rect 4658 346 4667 380
rect 4667 346 4701 380
rect 4701 346 4710 380
rect 4658 340 4710 346
rect 4381 328 4433 334
rect 5221 440 5273 444
rect 5221 406 5230 440
rect 5230 406 5264 440
rect 5264 406 5273 440
rect 5221 392 5273 406
rect 5221 368 5273 380
rect 5221 334 5230 368
rect 5230 334 5264 368
rect 5264 334 5273 368
rect 5221 328 5273 334
rect 5303 440 5355 444
rect 5303 406 5312 440
rect 5312 406 5346 440
rect 5346 406 5355 440
rect 5303 392 5355 406
rect 5607 452 5659 456
rect 5607 418 5613 452
rect 5613 418 5647 452
rect 5647 418 5659 452
rect 5607 404 5659 418
rect 5303 368 5355 380
rect 5303 334 5312 368
rect 5312 334 5346 368
rect 5346 334 5355 368
rect 5607 380 5659 392
rect 5607 346 5613 380
rect 5613 346 5647 380
rect 5647 346 5659 380
rect 5607 340 5659 346
rect 5884 440 5936 444
rect 5884 406 5893 440
rect 5893 406 5927 440
rect 5927 406 5936 440
rect 5884 392 5936 406
rect 5884 368 5936 380
rect 5884 334 5893 368
rect 5893 334 5927 368
rect 5927 334 5936 368
rect 5303 328 5355 334
rect 5884 328 5936 334
rect 6056 436 6108 445
rect 6056 402 6060 436
rect 6060 402 6094 436
rect 6094 402 6108 436
rect 6056 393 6108 402
rect 6120 436 6172 445
rect 6120 402 6132 436
rect 6132 402 6166 436
rect 6166 402 6172 436
rect 6120 393 6172 402
rect 6054 -134 6106 -82
rect 6118 -134 6170 -82
<< metal2 >>
rect 4658 701 4664 753
rect 4716 701 4728 753
rect 4780 701 4786 753
rect 4658 673 4716 701
tri 4716 673 4744 701 nw
rect 4218 621 4224 673
rect 4276 621 4288 673
rect 4340 621 4346 673
tri 4260 593 4288 621 ne
rect 4288 593 4346 621
rect 3912 541 3918 593
rect 3970 541 3982 593
rect 4034 541 4040 593
tri 4288 587 4294 593 ne
rect 3912 445 3964 541
tri 3964 507 3998 541 nw
tri 3964 445 3967 448 sw
rect 4294 445 4346 593
rect 3912 414 3967 445
tri 3967 414 3998 445 sw
rect 3912 362 3918 414
rect 3970 362 3982 414
rect 4034 362 4040 414
rect 4294 381 4346 393
rect 4294 323 4346 329
rect 4381 621 4439 673
rect 4491 621 4503 673
rect 4555 621 4561 673
rect 4381 444 4433 621
tri 4433 587 4467 621 nw
rect 4381 380 4433 392
rect 4658 456 4710 673
tri 4710 667 4716 673 nw
rect 5303 621 5309 673
rect 5361 621 5373 673
rect 5425 621 5431 673
rect 5850 621 5856 673
rect 5908 621 5920 673
rect 5972 621 5978 673
rect 4658 392 4710 404
rect 4658 334 4710 340
rect 5221 444 5273 450
rect 5221 380 5273 392
rect 4381 322 4433 328
rect 5221 322 5273 328
rect 5303 444 5355 621
tri 5355 587 5389 621 nw
tri 5850 587 5884 621 ne
rect 5303 380 5355 392
rect 5607 456 5659 462
rect 5607 392 5659 404
rect 5607 334 5659 340
rect 5884 444 5936 621
tri 5936 587 5970 621 nw
rect 5884 380 5936 392
rect 5303 322 5355 328
rect 5884 322 5936 328
rect 6048 393 6056 445
rect 6108 393 6120 445
rect 6172 393 6178 445
rect 6048 -82 6100 393
tri 6100 359 6134 393 nw
tri 6100 -82 6143 -39 sw
rect 6048 -134 6054 -82
rect 6106 -134 6118 -82
rect 6170 -134 6176 -82
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1701704242
transform -1 0 5800 0 1 2
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1701704242
transform 1 0 2551 0 1 2
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1701704242
transform 1 0 6190 0 1 2
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_3
timestamp 1701704242
transform 1 0 504 0 1 2
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_4
timestamp 1701704242
transform 1 0 1714 0 1 2
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_5
timestamp 1701704242
transform 1 0 3302 0 1 2
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1701704242
transform 1 0 6476 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1701704242
transform 1 0 1252 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1701704242
transform 1 0 42 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1701704242
transform -1 0 5514 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_4
timestamp 1701704242
transform -1 0 4587 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_5
timestamp 1701704242
transform -1 0 1324 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_6
timestamp 1701704242
transform 1 0 5728 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1701704242
transform 1 0 3588 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1701704242
transform 1 0 4515 0 1 2
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_2
timestamp 1701704242
transform 1 0 2837 0 1 2
box 107 226 460 873
<< labels >>
flabel metal1 s 370 401 484 436 3 FreeSans 200 0 0 0 DM_H_N[0]
port 2 nsew
flabel metal1 s 137 405 237 435 3 FreeSans 100 0 0 0 DM_H_N[1]
port 3 nsew
flabel metal1 s 1592 403 1689 435 3 FreeSans 100 0 0 0 INP_DIS_H_N
port 4 nsew
flabel metal1 s 1871 366 1900 434 3 FreeSans 100 90 0 0 INP_DIS_I_H
port 5 nsew
flabel metal1 s 1968 381 1992 460 3 FreeSans 100 0 0 0 INP_DIS_I_H_N
port 6 nsew
flabel metal1 s 2710 350 2734 419 3 FreeSans 100 90 0 0 VTRIP_SEL_H
port 7 nsew
flabel metal1 s 3449 350 3476 443 3 FreeSans 100 0 0 0 TRIPSEL_I_H
port 8 nsew
flabel metal1 s 3561 350 3588 444 3 FreeSans 100 0 0 0 TRIPSEL_I_H_N
port 9 nsew
flabel metal1 s 3741 364 3768 472 3 FreeSans 100 0 0 0 IBUF_MODE_SEL[1]
port 10 nsew
flabel metal1 s 3941 376 4023 407 3 FreeSans 100 0 0 0 IBUF_MODE_SEL[0]
port 11 nsew
flabel metal1 s 5232 347 5266 432 3 FreeSans 100 0 0 0 MODE_VCCD_N
port 12 nsew
flabel metal1 s 6334 359 6365 436 3 FreeSans 100 0 0 0 MODE_REF_N
port 13 nsew
flabel metal1 s 6831 342 6858 433 3 FreeSans 100 0 0 0 HYS_TRIM
port 14 nsew
flabel metal1 s 6724 344 6759 442 3 FreeSans 100 0 0 0 MODE_REF_3V_N
port 15 nsew
flabel metal1 s 1137 405 1215 431 3 FreeSans 100 0 0 0 DM_H_N[2]
port 16 nsew
flabel metal1 s 4309 345 4337 439 3 FreeSans 100 0 0 0 MODE_NORMAL_N
port 17 nsew
flabel metal1 s 102 885 445 1044 3 FreeSans 100 0 0 0 VDDIO_Q
port 18 nsew
flabel metal1 s 106 46 259 205 3 FreeSans 100 0 0 0 VSSD
port 19 nsew
<< properties >>
string GDS_END 63679252
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 63631630
<< end >>
