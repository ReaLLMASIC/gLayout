magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< locali >>
rect 567 1431 601 1447
rect 567 1381 601 1397
rect 1735 1431 1769 1447
rect 1735 1381 1769 1397
rect 2903 1431 2937 1447
rect 2903 1381 2937 1397
rect 4071 1431 4105 1447
rect 4071 1381 4105 1397
rect 5239 1431 5273 1447
rect 5239 1381 5273 1397
rect 6407 1431 6441 1447
rect 6407 1381 6441 1397
rect 7575 1431 7609 1447
rect 7575 1381 7609 1397
rect 8743 1431 8777 1447
rect 8743 1381 8777 1397
rect 9911 1431 9945 1447
rect 9911 1381 9945 1397
rect 11079 1431 11113 1447
rect 11079 1381 11113 1397
rect 12247 1431 12281 1447
rect 12247 1381 12281 1397
rect 13415 1431 13449 1447
rect 13415 1381 13449 1397
rect 14583 1431 14617 1447
rect 14583 1381 14617 1397
rect 15751 1431 15785 1447
rect 15751 1381 15785 1397
rect 16919 1431 16953 1447
rect 16919 1381 16953 1397
rect 18087 1431 18121 1447
rect 18087 1381 18121 1397
rect 19255 1431 19289 1447
rect 19255 1381 19289 1397
rect 20423 1431 20457 1447
rect 20423 1381 20457 1397
rect 21591 1431 21625 1447
rect 21591 1381 21625 1397
rect 22759 1431 22793 1447
rect 22759 1381 22793 1397
rect 23927 1431 23961 1447
rect 23927 1381 23961 1397
rect 25095 1431 25129 1447
rect 25095 1381 25129 1397
rect 26263 1431 26297 1447
rect 26263 1381 26297 1397
rect 27431 1431 27465 1447
rect 27431 1381 27465 1397
rect 28599 1431 28633 1447
rect 28599 1381 28633 1397
rect 29767 1431 29801 1447
rect 29767 1381 29801 1397
rect 30935 1431 30969 1447
rect 30935 1381 30969 1397
rect 32103 1431 32137 1447
rect 32103 1381 32137 1397
rect 33271 1431 33305 1447
rect 33271 1381 33305 1397
rect 34439 1431 34473 1447
rect 34439 1381 34473 1397
rect 35607 1431 35641 1447
rect 35607 1381 35641 1397
rect 36775 1431 36809 1447
rect 36775 1381 36809 1397
rect 567 17 601 33
rect 567 -33 601 -17
rect 1735 17 1769 33
rect 1735 -33 1769 -17
rect 2903 17 2937 33
rect 2903 -33 2937 -17
rect 4071 17 4105 33
rect 4071 -33 4105 -17
rect 5239 17 5273 33
rect 5239 -33 5273 -17
rect 6407 17 6441 33
rect 6407 -33 6441 -17
rect 7575 17 7609 33
rect 7575 -33 7609 -17
rect 8743 17 8777 33
rect 8743 -33 8777 -17
rect 9911 17 9945 33
rect 9911 -33 9945 -17
rect 11079 17 11113 33
rect 11079 -33 11113 -17
rect 12247 17 12281 33
rect 12247 -33 12281 -17
rect 13415 17 13449 33
rect 13415 -33 13449 -17
rect 14583 17 14617 33
rect 14583 -33 14617 -17
rect 15751 17 15785 33
rect 15751 -33 15785 -17
rect 16919 17 16953 33
rect 16919 -33 16953 -17
rect 18087 17 18121 33
rect 18087 -33 18121 -17
rect 19255 17 19289 33
rect 19255 -33 19289 -17
rect 20423 17 20457 33
rect 20423 -33 20457 -17
rect 21591 17 21625 33
rect 21591 -33 21625 -17
rect 22759 17 22793 33
rect 22759 -33 22793 -17
rect 23927 17 23961 33
rect 23927 -33 23961 -17
rect 25095 17 25129 33
rect 25095 -33 25129 -17
rect 26263 17 26297 33
rect 26263 -33 26297 -17
rect 27431 17 27465 33
rect 27431 -33 27465 -17
rect 28599 17 28633 33
rect 28599 -33 28633 -17
rect 29767 17 29801 33
rect 29767 -33 29801 -17
rect 30935 17 30969 33
rect 30935 -33 30969 -17
rect 32103 17 32137 33
rect 32103 -33 32137 -17
rect 33271 17 33305 33
rect 33271 -33 33305 -17
rect 34439 17 34473 33
rect 34439 -33 34473 -17
rect 35607 17 35641 33
rect 35607 -33 35641 -17
rect 36775 17 36809 33
rect 36775 -33 36809 -17
<< viali >>
rect 567 1397 601 1431
rect 1735 1397 1769 1431
rect 2903 1397 2937 1431
rect 4071 1397 4105 1431
rect 5239 1397 5273 1431
rect 6407 1397 6441 1431
rect 7575 1397 7609 1431
rect 8743 1397 8777 1431
rect 9911 1397 9945 1431
rect 11079 1397 11113 1431
rect 12247 1397 12281 1431
rect 13415 1397 13449 1431
rect 14583 1397 14617 1431
rect 15751 1397 15785 1431
rect 16919 1397 16953 1431
rect 18087 1397 18121 1431
rect 19255 1397 19289 1431
rect 20423 1397 20457 1431
rect 21591 1397 21625 1431
rect 22759 1397 22793 1431
rect 23927 1397 23961 1431
rect 25095 1397 25129 1431
rect 26263 1397 26297 1431
rect 27431 1397 27465 1431
rect 28599 1397 28633 1431
rect 29767 1397 29801 1431
rect 30935 1397 30969 1431
rect 32103 1397 32137 1431
rect 33271 1397 33305 1431
rect 34439 1397 34473 1431
rect 35607 1397 35641 1431
rect 36775 1397 36809 1431
rect 567 -17 601 17
rect 1735 -17 1769 17
rect 2903 -17 2937 17
rect 4071 -17 4105 17
rect 5239 -17 5273 17
rect 6407 -17 6441 17
rect 7575 -17 7609 17
rect 8743 -17 8777 17
rect 9911 -17 9945 17
rect 11079 -17 11113 17
rect 12247 -17 12281 17
rect 13415 -17 13449 17
rect 14583 -17 14617 17
rect 15751 -17 15785 17
rect 16919 -17 16953 17
rect 18087 -17 18121 17
rect 19255 -17 19289 17
rect 20423 -17 20457 17
rect 21591 -17 21625 17
rect 22759 -17 22793 17
rect 23927 -17 23961 17
rect 25095 -17 25129 17
rect 26263 -17 26297 17
rect 27431 -17 27465 17
rect 28599 -17 28633 17
rect 29767 -17 29801 17
rect 30935 -17 30969 17
rect 32103 -17 32137 17
rect 33271 -17 33305 17
rect 34439 -17 34473 17
rect 35607 -17 35641 17
rect 36775 -17 36809 17
<< metal1 >>
rect 552 1388 558 1440
rect 610 1388 616 1440
rect 1720 1388 1726 1440
rect 1778 1388 1784 1440
rect 2888 1388 2894 1440
rect 2946 1388 2952 1440
rect 4056 1388 4062 1440
rect 4114 1388 4120 1440
rect 5224 1388 5230 1440
rect 5282 1388 5288 1440
rect 6392 1388 6398 1440
rect 6450 1388 6456 1440
rect 7560 1388 7566 1440
rect 7618 1388 7624 1440
rect 8728 1388 8734 1440
rect 8786 1388 8792 1440
rect 9896 1388 9902 1440
rect 9954 1388 9960 1440
rect 11064 1388 11070 1440
rect 11122 1388 11128 1440
rect 12232 1388 12238 1440
rect 12290 1388 12296 1440
rect 13400 1388 13406 1440
rect 13458 1388 13464 1440
rect 14568 1388 14574 1440
rect 14626 1388 14632 1440
rect 15736 1388 15742 1440
rect 15794 1388 15800 1440
rect 16904 1388 16910 1440
rect 16962 1388 16968 1440
rect 18072 1388 18078 1440
rect 18130 1388 18136 1440
rect 19240 1388 19246 1440
rect 19298 1388 19304 1440
rect 20408 1388 20414 1440
rect 20466 1388 20472 1440
rect 21576 1388 21582 1440
rect 21634 1388 21640 1440
rect 22744 1388 22750 1440
rect 22802 1388 22808 1440
rect 23912 1388 23918 1440
rect 23970 1388 23976 1440
rect 25080 1388 25086 1440
rect 25138 1388 25144 1440
rect 26248 1388 26254 1440
rect 26306 1388 26312 1440
rect 27416 1388 27422 1440
rect 27474 1388 27480 1440
rect 28584 1388 28590 1440
rect 28642 1388 28648 1440
rect 29752 1388 29758 1440
rect 29810 1388 29816 1440
rect 30920 1388 30926 1440
rect 30978 1388 30984 1440
rect 32088 1388 32094 1440
rect 32146 1388 32152 1440
rect 33256 1388 33262 1440
rect 33314 1388 33320 1440
rect 34424 1388 34430 1440
rect 34482 1388 34488 1440
rect 35592 1388 35598 1440
rect 35650 1388 35656 1440
rect 36760 1388 36766 1440
rect 36818 1388 36824 1440
rect 552 -26 558 26
rect 610 -26 616 26
rect 1720 -26 1726 26
rect 1778 -26 1784 26
rect 2888 -26 2894 26
rect 2946 -26 2952 26
rect 4056 -26 4062 26
rect 4114 -26 4120 26
rect 5224 -26 5230 26
rect 5282 -26 5288 26
rect 6392 -26 6398 26
rect 6450 -26 6456 26
rect 7560 -26 7566 26
rect 7618 -26 7624 26
rect 8728 -26 8734 26
rect 8786 -26 8792 26
rect 9896 -26 9902 26
rect 9954 -26 9960 26
rect 11064 -26 11070 26
rect 11122 -26 11128 26
rect 12232 -26 12238 26
rect 12290 -26 12296 26
rect 13400 -26 13406 26
rect 13458 -26 13464 26
rect 14568 -26 14574 26
rect 14626 -26 14632 26
rect 15736 -26 15742 26
rect 15794 -26 15800 26
rect 16904 -26 16910 26
rect 16962 -26 16968 26
rect 18072 -26 18078 26
rect 18130 -26 18136 26
rect 19240 -26 19246 26
rect 19298 -26 19304 26
rect 20408 -26 20414 26
rect 20466 -26 20472 26
rect 21576 -26 21582 26
rect 21634 -26 21640 26
rect 22744 -26 22750 26
rect 22802 -26 22808 26
rect 23912 -26 23918 26
rect 23970 -26 23976 26
rect 25080 -26 25086 26
rect 25138 -26 25144 26
rect 26248 -26 26254 26
rect 26306 -26 26312 26
rect 27416 -26 27422 26
rect 27474 -26 27480 26
rect 28584 -26 28590 26
rect 28642 -26 28648 26
rect 29752 -26 29758 26
rect 29810 -26 29816 26
rect 30920 -26 30926 26
rect 30978 -26 30984 26
rect 32088 -26 32094 26
rect 32146 -26 32152 26
rect 33256 -26 33262 26
rect 33314 -26 33320 26
rect 34424 -26 34430 26
rect 34482 -26 34488 26
rect 35592 -26 35598 26
rect 35650 -26 35656 26
rect 36760 -26 36766 26
rect 36818 -26 36824 26
<< via1 >>
rect 558 1431 610 1440
rect 558 1397 567 1431
rect 567 1397 601 1431
rect 601 1397 610 1431
rect 558 1388 610 1397
rect 1726 1431 1778 1440
rect 1726 1397 1735 1431
rect 1735 1397 1769 1431
rect 1769 1397 1778 1431
rect 1726 1388 1778 1397
rect 2894 1431 2946 1440
rect 2894 1397 2903 1431
rect 2903 1397 2937 1431
rect 2937 1397 2946 1431
rect 2894 1388 2946 1397
rect 4062 1431 4114 1440
rect 4062 1397 4071 1431
rect 4071 1397 4105 1431
rect 4105 1397 4114 1431
rect 4062 1388 4114 1397
rect 5230 1431 5282 1440
rect 5230 1397 5239 1431
rect 5239 1397 5273 1431
rect 5273 1397 5282 1431
rect 5230 1388 5282 1397
rect 6398 1431 6450 1440
rect 6398 1397 6407 1431
rect 6407 1397 6441 1431
rect 6441 1397 6450 1431
rect 6398 1388 6450 1397
rect 7566 1431 7618 1440
rect 7566 1397 7575 1431
rect 7575 1397 7609 1431
rect 7609 1397 7618 1431
rect 7566 1388 7618 1397
rect 8734 1431 8786 1440
rect 8734 1397 8743 1431
rect 8743 1397 8777 1431
rect 8777 1397 8786 1431
rect 8734 1388 8786 1397
rect 9902 1431 9954 1440
rect 9902 1397 9911 1431
rect 9911 1397 9945 1431
rect 9945 1397 9954 1431
rect 9902 1388 9954 1397
rect 11070 1431 11122 1440
rect 11070 1397 11079 1431
rect 11079 1397 11113 1431
rect 11113 1397 11122 1431
rect 11070 1388 11122 1397
rect 12238 1431 12290 1440
rect 12238 1397 12247 1431
rect 12247 1397 12281 1431
rect 12281 1397 12290 1431
rect 12238 1388 12290 1397
rect 13406 1431 13458 1440
rect 13406 1397 13415 1431
rect 13415 1397 13449 1431
rect 13449 1397 13458 1431
rect 13406 1388 13458 1397
rect 14574 1431 14626 1440
rect 14574 1397 14583 1431
rect 14583 1397 14617 1431
rect 14617 1397 14626 1431
rect 14574 1388 14626 1397
rect 15742 1431 15794 1440
rect 15742 1397 15751 1431
rect 15751 1397 15785 1431
rect 15785 1397 15794 1431
rect 15742 1388 15794 1397
rect 16910 1431 16962 1440
rect 16910 1397 16919 1431
rect 16919 1397 16953 1431
rect 16953 1397 16962 1431
rect 16910 1388 16962 1397
rect 18078 1431 18130 1440
rect 18078 1397 18087 1431
rect 18087 1397 18121 1431
rect 18121 1397 18130 1431
rect 18078 1388 18130 1397
rect 19246 1431 19298 1440
rect 19246 1397 19255 1431
rect 19255 1397 19289 1431
rect 19289 1397 19298 1431
rect 19246 1388 19298 1397
rect 20414 1431 20466 1440
rect 20414 1397 20423 1431
rect 20423 1397 20457 1431
rect 20457 1397 20466 1431
rect 20414 1388 20466 1397
rect 21582 1431 21634 1440
rect 21582 1397 21591 1431
rect 21591 1397 21625 1431
rect 21625 1397 21634 1431
rect 21582 1388 21634 1397
rect 22750 1431 22802 1440
rect 22750 1397 22759 1431
rect 22759 1397 22793 1431
rect 22793 1397 22802 1431
rect 22750 1388 22802 1397
rect 23918 1431 23970 1440
rect 23918 1397 23927 1431
rect 23927 1397 23961 1431
rect 23961 1397 23970 1431
rect 23918 1388 23970 1397
rect 25086 1431 25138 1440
rect 25086 1397 25095 1431
rect 25095 1397 25129 1431
rect 25129 1397 25138 1431
rect 25086 1388 25138 1397
rect 26254 1431 26306 1440
rect 26254 1397 26263 1431
rect 26263 1397 26297 1431
rect 26297 1397 26306 1431
rect 26254 1388 26306 1397
rect 27422 1431 27474 1440
rect 27422 1397 27431 1431
rect 27431 1397 27465 1431
rect 27465 1397 27474 1431
rect 27422 1388 27474 1397
rect 28590 1431 28642 1440
rect 28590 1397 28599 1431
rect 28599 1397 28633 1431
rect 28633 1397 28642 1431
rect 28590 1388 28642 1397
rect 29758 1431 29810 1440
rect 29758 1397 29767 1431
rect 29767 1397 29801 1431
rect 29801 1397 29810 1431
rect 29758 1388 29810 1397
rect 30926 1431 30978 1440
rect 30926 1397 30935 1431
rect 30935 1397 30969 1431
rect 30969 1397 30978 1431
rect 30926 1388 30978 1397
rect 32094 1431 32146 1440
rect 32094 1397 32103 1431
rect 32103 1397 32137 1431
rect 32137 1397 32146 1431
rect 32094 1388 32146 1397
rect 33262 1431 33314 1440
rect 33262 1397 33271 1431
rect 33271 1397 33305 1431
rect 33305 1397 33314 1431
rect 33262 1388 33314 1397
rect 34430 1431 34482 1440
rect 34430 1397 34439 1431
rect 34439 1397 34473 1431
rect 34473 1397 34482 1431
rect 34430 1388 34482 1397
rect 35598 1431 35650 1440
rect 35598 1397 35607 1431
rect 35607 1397 35641 1431
rect 35641 1397 35650 1431
rect 35598 1388 35650 1397
rect 36766 1431 36818 1440
rect 36766 1397 36775 1431
rect 36775 1397 36809 1431
rect 36809 1397 36818 1431
rect 36766 1388 36818 1397
rect 558 17 610 26
rect 558 -17 567 17
rect 567 -17 601 17
rect 601 -17 610 17
rect 558 -26 610 -17
rect 1726 17 1778 26
rect 1726 -17 1735 17
rect 1735 -17 1769 17
rect 1769 -17 1778 17
rect 1726 -26 1778 -17
rect 2894 17 2946 26
rect 2894 -17 2903 17
rect 2903 -17 2937 17
rect 2937 -17 2946 17
rect 2894 -26 2946 -17
rect 4062 17 4114 26
rect 4062 -17 4071 17
rect 4071 -17 4105 17
rect 4105 -17 4114 17
rect 4062 -26 4114 -17
rect 5230 17 5282 26
rect 5230 -17 5239 17
rect 5239 -17 5273 17
rect 5273 -17 5282 17
rect 5230 -26 5282 -17
rect 6398 17 6450 26
rect 6398 -17 6407 17
rect 6407 -17 6441 17
rect 6441 -17 6450 17
rect 6398 -26 6450 -17
rect 7566 17 7618 26
rect 7566 -17 7575 17
rect 7575 -17 7609 17
rect 7609 -17 7618 17
rect 7566 -26 7618 -17
rect 8734 17 8786 26
rect 8734 -17 8743 17
rect 8743 -17 8777 17
rect 8777 -17 8786 17
rect 8734 -26 8786 -17
rect 9902 17 9954 26
rect 9902 -17 9911 17
rect 9911 -17 9945 17
rect 9945 -17 9954 17
rect 9902 -26 9954 -17
rect 11070 17 11122 26
rect 11070 -17 11079 17
rect 11079 -17 11113 17
rect 11113 -17 11122 17
rect 11070 -26 11122 -17
rect 12238 17 12290 26
rect 12238 -17 12247 17
rect 12247 -17 12281 17
rect 12281 -17 12290 17
rect 12238 -26 12290 -17
rect 13406 17 13458 26
rect 13406 -17 13415 17
rect 13415 -17 13449 17
rect 13449 -17 13458 17
rect 13406 -26 13458 -17
rect 14574 17 14626 26
rect 14574 -17 14583 17
rect 14583 -17 14617 17
rect 14617 -17 14626 17
rect 14574 -26 14626 -17
rect 15742 17 15794 26
rect 15742 -17 15751 17
rect 15751 -17 15785 17
rect 15785 -17 15794 17
rect 15742 -26 15794 -17
rect 16910 17 16962 26
rect 16910 -17 16919 17
rect 16919 -17 16953 17
rect 16953 -17 16962 17
rect 16910 -26 16962 -17
rect 18078 17 18130 26
rect 18078 -17 18087 17
rect 18087 -17 18121 17
rect 18121 -17 18130 17
rect 18078 -26 18130 -17
rect 19246 17 19298 26
rect 19246 -17 19255 17
rect 19255 -17 19289 17
rect 19289 -17 19298 17
rect 19246 -26 19298 -17
rect 20414 17 20466 26
rect 20414 -17 20423 17
rect 20423 -17 20457 17
rect 20457 -17 20466 17
rect 20414 -26 20466 -17
rect 21582 17 21634 26
rect 21582 -17 21591 17
rect 21591 -17 21625 17
rect 21625 -17 21634 17
rect 21582 -26 21634 -17
rect 22750 17 22802 26
rect 22750 -17 22759 17
rect 22759 -17 22793 17
rect 22793 -17 22802 17
rect 22750 -26 22802 -17
rect 23918 17 23970 26
rect 23918 -17 23927 17
rect 23927 -17 23961 17
rect 23961 -17 23970 17
rect 23918 -26 23970 -17
rect 25086 17 25138 26
rect 25086 -17 25095 17
rect 25095 -17 25129 17
rect 25129 -17 25138 17
rect 25086 -26 25138 -17
rect 26254 17 26306 26
rect 26254 -17 26263 17
rect 26263 -17 26297 17
rect 26297 -17 26306 17
rect 26254 -26 26306 -17
rect 27422 17 27474 26
rect 27422 -17 27431 17
rect 27431 -17 27465 17
rect 27465 -17 27474 17
rect 27422 -26 27474 -17
rect 28590 17 28642 26
rect 28590 -17 28599 17
rect 28599 -17 28633 17
rect 28633 -17 28642 17
rect 28590 -26 28642 -17
rect 29758 17 29810 26
rect 29758 -17 29767 17
rect 29767 -17 29801 17
rect 29801 -17 29810 17
rect 29758 -26 29810 -17
rect 30926 17 30978 26
rect 30926 -17 30935 17
rect 30935 -17 30969 17
rect 30969 -17 30978 17
rect 30926 -26 30978 -17
rect 32094 17 32146 26
rect 32094 -17 32103 17
rect 32103 -17 32137 17
rect 32137 -17 32146 17
rect 32094 -26 32146 -17
rect 33262 17 33314 26
rect 33262 -17 33271 17
rect 33271 -17 33305 17
rect 33305 -17 33314 17
rect 33262 -26 33314 -17
rect 34430 17 34482 26
rect 34430 -17 34439 17
rect 34439 -17 34473 17
rect 34473 -17 34482 17
rect 34430 -26 34482 -17
rect 35598 17 35650 26
rect 35598 -17 35607 17
rect 35607 -17 35641 17
rect 35641 -17 35650 17
rect 35598 -26 35650 -17
rect 36766 17 36818 26
rect 36766 -17 36775 17
rect 36775 -17 36809 17
rect 36809 -17 36818 17
rect 36766 -26 36818 -17
<< metal2 >>
rect 556 1442 612 1451
rect 137 538 203 590
rect 369 345 397 1414
rect 1724 1442 1780 1451
rect 556 1377 612 1386
rect 1082 609 1148 661
rect 1305 538 1371 590
rect 1537 345 1565 1414
rect 2892 1442 2948 1451
rect 1724 1377 1780 1386
rect 2250 609 2316 661
rect 2473 538 2539 590
rect 2705 345 2733 1414
rect 4060 1442 4116 1451
rect 2892 1377 2948 1386
rect 3418 609 3484 661
rect 3641 538 3707 590
rect 3873 345 3901 1414
rect 5228 1442 5284 1451
rect 4060 1377 4116 1386
rect 4586 609 4652 661
rect 4809 538 4875 590
rect 5041 345 5069 1414
rect 6396 1442 6452 1451
rect 5228 1377 5284 1386
rect 5754 609 5820 661
rect 5977 538 6043 590
rect 6209 345 6237 1414
rect 7564 1442 7620 1451
rect 6396 1377 6452 1386
rect 6922 609 6988 661
rect 7145 538 7211 590
rect 7377 345 7405 1414
rect 8732 1442 8788 1451
rect 7564 1377 7620 1386
rect 8090 609 8156 661
rect 8313 538 8379 590
rect 8545 345 8573 1414
rect 9900 1442 9956 1451
rect 8732 1377 8788 1386
rect 9258 609 9324 661
rect 9481 538 9547 590
rect 9713 345 9741 1414
rect 11068 1442 11124 1451
rect 9900 1377 9956 1386
rect 10426 609 10492 661
rect 10649 538 10715 590
rect 10881 345 10909 1414
rect 12236 1442 12292 1451
rect 11068 1377 11124 1386
rect 11594 609 11660 661
rect 11817 538 11883 590
rect 12049 345 12077 1414
rect 13404 1442 13460 1451
rect 12236 1377 12292 1386
rect 12762 609 12828 661
rect 12985 538 13051 590
rect 13217 345 13245 1414
rect 14572 1442 14628 1451
rect 13404 1377 13460 1386
rect 13930 609 13996 661
rect 14153 538 14219 590
rect 14385 345 14413 1414
rect 15740 1442 15796 1451
rect 14572 1377 14628 1386
rect 15098 609 15164 661
rect 15321 538 15387 590
rect 15553 345 15581 1414
rect 16908 1442 16964 1451
rect 15740 1377 15796 1386
rect 16266 609 16332 661
rect 16489 538 16555 590
rect 16721 345 16749 1414
rect 18076 1442 18132 1451
rect 16908 1377 16964 1386
rect 17434 609 17500 661
rect 17657 538 17723 590
rect 17889 345 17917 1414
rect 19244 1442 19300 1451
rect 18076 1377 18132 1386
rect 18602 609 18668 661
rect 18825 538 18891 590
rect 19057 345 19085 1414
rect 20412 1442 20468 1451
rect 19244 1377 19300 1386
rect 19770 609 19836 661
rect 19993 538 20059 590
rect 20225 345 20253 1414
rect 21580 1442 21636 1451
rect 20412 1377 20468 1386
rect 20938 609 21004 661
rect 21161 538 21227 590
rect 21393 345 21421 1414
rect 22748 1442 22804 1451
rect 21580 1377 21636 1386
rect 22106 609 22172 661
rect 22329 538 22395 590
rect 22561 345 22589 1414
rect 23916 1442 23972 1451
rect 22748 1377 22804 1386
rect 23274 609 23340 661
rect 23497 538 23563 590
rect 23729 345 23757 1414
rect 25084 1442 25140 1451
rect 23916 1377 23972 1386
rect 24442 609 24508 661
rect 24665 538 24731 590
rect 24897 345 24925 1414
rect 26252 1442 26308 1451
rect 25084 1377 25140 1386
rect 25610 609 25676 661
rect 25833 538 25899 590
rect 26065 345 26093 1414
rect 27420 1442 27476 1451
rect 26252 1377 26308 1386
rect 26778 609 26844 661
rect 27001 538 27067 590
rect 27233 345 27261 1414
rect 28588 1442 28644 1451
rect 27420 1377 27476 1386
rect 27946 609 28012 661
rect 28169 538 28235 590
rect 28401 345 28429 1414
rect 29756 1442 29812 1451
rect 28588 1377 28644 1386
rect 29114 609 29180 661
rect 29337 538 29403 590
rect 29569 345 29597 1414
rect 30924 1442 30980 1451
rect 29756 1377 29812 1386
rect 30282 609 30348 661
rect 30505 538 30571 590
rect 30737 345 30765 1414
rect 32092 1442 32148 1451
rect 30924 1377 30980 1386
rect 31450 609 31516 661
rect 31673 538 31739 590
rect 31905 345 31933 1414
rect 33260 1442 33316 1451
rect 32092 1377 32148 1386
rect 32618 609 32684 661
rect 32841 538 32907 590
rect 33073 345 33101 1414
rect 34428 1442 34484 1451
rect 33260 1377 33316 1386
rect 33786 609 33852 661
rect 34009 538 34075 590
rect 34241 345 34269 1414
rect 35596 1442 35652 1451
rect 34428 1377 34484 1386
rect 34954 609 35020 661
rect 35177 538 35243 590
rect 35409 345 35437 1414
rect 36764 1442 36820 1451
rect 35596 1377 35652 1386
rect 36122 609 36188 661
rect 36345 538 36411 590
rect 36577 345 36605 1414
rect 36764 1377 36820 1386
rect 37290 609 37356 661
rect 368 336 424 345
rect 368 271 424 280
rect 1536 336 1592 345
rect 1536 271 1592 280
rect 2704 336 2760 345
rect 2704 271 2760 280
rect 3872 336 3928 345
rect 3872 271 3928 280
rect 5040 336 5096 345
rect 5040 271 5096 280
rect 6208 336 6264 345
rect 6208 271 6264 280
rect 7376 336 7432 345
rect 7376 271 7432 280
rect 8544 336 8600 345
rect 8544 271 8600 280
rect 9712 336 9768 345
rect 9712 271 9768 280
rect 10880 336 10936 345
rect 10880 271 10936 280
rect 12048 336 12104 345
rect 12048 271 12104 280
rect 13216 336 13272 345
rect 13216 271 13272 280
rect 14384 336 14440 345
rect 14384 271 14440 280
rect 15552 336 15608 345
rect 15552 271 15608 280
rect 16720 336 16776 345
rect 16720 271 16776 280
rect 17888 336 17944 345
rect 17888 271 17944 280
rect 19056 336 19112 345
rect 19056 271 19112 280
rect 20224 336 20280 345
rect 20224 271 20280 280
rect 21392 336 21448 345
rect 21392 271 21448 280
rect 22560 336 22616 345
rect 22560 271 22616 280
rect 23728 336 23784 345
rect 23728 271 23784 280
rect 24896 336 24952 345
rect 24896 271 24952 280
rect 26064 336 26120 345
rect 26064 271 26120 280
rect 27232 336 27288 345
rect 27232 271 27288 280
rect 28400 336 28456 345
rect 28400 271 28456 280
rect 29568 336 29624 345
rect 29568 271 29624 280
rect 30736 336 30792 345
rect 30736 271 30792 280
rect 31904 336 31960 345
rect 31904 271 31960 280
rect 33072 336 33128 345
rect 33072 271 33128 280
rect 34240 336 34296 345
rect 34240 271 34296 280
rect 35408 336 35464 345
rect 35408 271 35464 280
rect 36576 336 36632 345
rect 36576 271 36632 280
rect 369 0 397 271
rect 556 28 612 37
rect 1537 0 1565 271
rect 1724 28 1780 37
rect 556 -37 612 -28
rect 2705 0 2733 271
rect 2892 28 2948 37
rect 1724 -37 1780 -28
rect 3873 0 3901 271
rect 4060 28 4116 37
rect 2892 -37 2948 -28
rect 5041 0 5069 271
rect 5228 28 5284 37
rect 4060 -37 4116 -28
rect 6209 0 6237 271
rect 6396 28 6452 37
rect 5228 -37 5284 -28
rect 7377 0 7405 271
rect 7564 28 7620 37
rect 6396 -37 6452 -28
rect 8545 0 8573 271
rect 8732 28 8788 37
rect 7564 -37 7620 -28
rect 9713 0 9741 271
rect 9900 28 9956 37
rect 8732 -37 8788 -28
rect 10881 0 10909 271
rect 11068 28 11124 37
rect 9900 -37 9956 -28
rect 12049 0 12077 271
rect 12236 28 12292 37
rect 11068 -37 11124 -28
rect 13217 0 13245 271
rect 13404 28 13460 37
rect 12236 -37 12292 -28
rect 14385 0 14413 271
rect 14572 28 14628 37
rect 13404 -37 13460 -28
rect 15553 0 15581 271
rect 15740 28 15796 37
rect 14572 -37 14628 -28
rect 16721 0 16749 271
rect 16908 28 16964 37
rect 15740 -37 15796 -28
rect 17889 0 17917 271
rect 18076 28 18132 37
rect 16908 -37 16964 -28
rect 19057 0 19085 271
rect 19244 28 19300 37
rect 18076 -37 18132 -28
rect 20225 0 20253 271
rect 20412 28 20468 37
rect 19244 -37 19300 -28
rect 21393 0 21421 271
rect 21580 28 21636 37
rect 20412 -37 20468 -28
rect 22561 0 22589 271
rect 22748 28 22804 37
rect 21580 -37 21636 -28
rect 23729 0 23757 271
rect 23916 28 23972 37
rect 22748 -37 22804 -28
rect 24897 0 24925 271
rect 25084 28 25140 37
rect 23916 -37 23972 -28
rect 26065 0 26093 271
rect 26252 28 26308 37
rect 25084 -37 25140 -28
rect 27233 0 27261 271
rect 27420 28 27476 37
rect 26252 -37 26308 -28
rect 28401 0 28429 271
rect 28588 28 28644 37
rect 27420 -37 27476 -28
rect 29569 0 29597 271
rect 29756 28 29812 37
rect 28588 -37 28644 -28
rect 30737 0 30765 271
rect 30924 28 30980 37
rect 29756 -37 29812 -28
rect 31905 0 31933 271
rect 32092 28 32148 37
rect 30924 -37 30980 -28
rect 33073 0 33101 271
rect 33260 28 33316 37
rect 32092 -37 32148 -28
rect 34241 0 34269 271
rect 34428 28 34484 37
rect 33260 -37 33316 -28
rect 35409 0 35437 271
rect 35596 28 35652 37
rect 34428 -37 34484 -28
rect 36577 0 36605 271
rect 36764 28 36820 37
rect 35596 -37 35652 -28
rect 36764 -37 36820 -28
<< via2 >>
rect 556 1440 612 1442
rect 556 1388 558 1440
rect 558 1388 610 1440
rect 610 1388 612 1440
rect 1724 1440 1780 1442
rect 556 1386 612 1388
rect 1724 1388 1726 1440
rect 1726 1388 1778 1440
rect 1778 1388 1780 1440
rect 2892 1440 2948 1442
rect 1724 1386 1780 1388
rect 2892 1388 2894 1440
rect 2894 1388 2946 1440
rect 2946 1388 2948 1440
rect 4060 1440 4116 1442
rect 2892 1386 2948 1388
rect 4060 1388 4062 1440
rect 4062 1388 4114 1440
rect 4114 1388 4116 1440
rect 5228 1440 5284 1442
rect 4060 1386 4116 1388
rect 5228 1388 5230 1440
rect 5230 1388 5282 1440
rect 5282 1388 5284 1440
rect 6396 1440 6452 1442
rect 5228 1386 5284 1388
rect 6396 1388 6398 1440
rect 6398 1388 6450 1440
rect 6450 1388 6452 1440
rect 7564 1440 7620 1442
rect 6396 1386 6452 1388
rect 7564 1388 7566 1440
rect 7566 1388 7618 1440
rect 7618 1388 7620 1440
rect 8732 1440 8788 1442
rect 7564 1386 7620 1388
rect 8732 1388 8734 1440
rect 8734 1388 8786 1440
rect 8786 1388 8788 1440
rect 9900 1440 9956 1442
rect 8732 1386 8788 1388
rect 9900 1388 9902 1440
rect 9902 1388 9954 1440
rect 9954 1388 9956 1440
rect 11068 1440 11124 1442
rect 9900 1386 9956 1388
rect 11068 1388 11070 1440
rect 11070 1388 11122 1440
rect 11122 1388 11124 1440
rect 12236 1440 12292 1442
rect 11068 1386 11124 1388
rect 12236 1388 12238 1440
rect 12238 1388 12290 1440
rect 12290 1388 12292 1440
rect 13404 1440 13460 1442
rect 12236 1386 12292 1388
rect 13404 1388 13406 1440
rect 13406 1388 13458 1440
rect 13458 1388 13460 1440
rect 14572 1440 14628 1442
rect 13404 1386 13460 1388
rect 14572 1388 14574 1440
rect 14574 1388 14626 1440
rect 14626 1388 14628 1440
rect 15740 1440 15796 1442
rect 14572 1386 14628 1388
rect 15740 1388 15742 1440
rect 15742 1388 15794 1440
rect 15794 1388 15796 1440
rect 16908 1440 16964 1442
rect 15740 1386 15796 1388
rect 16908 1388 16910 1440
rect 16910 1388 16962 1440
rect 16962 1388 16964 1440
rect 18076 1440 18132 1442
rect 16908 1386 16964 1388
rect 18076 1388 18078 1440
rect 18078 1388 18130 1440
rect 18130 1388 18132 1440
rect 19244 1440 19300 1442
rect 18076 1386 18132 1388
rect 19244 1388 19246 1440
rect 19246 1388 19298 1440
rect 19298 1388 19300 1440
rect 20412 1440 20468 1442
rect 19244 1386 19300 1388
rect 20412 1388 20414 1440
rect 20414 1388 20466 1440
rect 20466 1388 20468 1440
rect 21580 1440 21636 1442
rect 20412 1386 20468 1388
rect 21580 1388 21582 1440
rect 21582 1388 21634 1440
rect 21634 1388 21636 1440
rect 22748 1440 22804 1442
rect 21580 1386 21636 1388
rect 22748 1388 22750 1440
rect 22750 1388 22802 1440
rect 22802 1388 22804 1440
rect 23916 1440 23972 1442
rect 22748 1386 22804 1388
rect 23916 1388 23918 1440
rect 23918 1388 23970 1440
rect 23970 1388 23972 1440
rect 25084 1440 25140 1442
rect 23916 1386 23972 1388
rect 25084 1388 25086 1440
rect 25086 1388 25138 1440
rect 25138 1388 25140 1440
rect 26252 1440 26308 1442
rect 25084 1386 25140 1388
rect 26252 1388 26254 1440
rect 26254 1388 26306 1440
rect 26306 1388 26308 1440
rect 27420 1440 27476 1442
rect 26252 1386 26308 1388
rect 27420 1388 27422 1440
rect 27422 1388 27474 1440
rect 27474 1388 27476 1440
rect 28588 1440 28644 1442
rect 27420 1386 27476 1388
rect 28588 1388 28590 1440
rect 28590 1388 28642 1440
rect 28642 1388 28644 1440
rect 29756 1440 29812 1442
rect 28588 1386 28644 1388
rect 29756 1388 29758 1440
rect 29758 1388 29810 1440
rect 29810 1388 29812 1440
rect 30924 1440 30980 1442
rect 29756 1386 29812 1388
rect 30924 1388 30926 1440
rect 30926 1388 30978 1440
rect 30978 1388 30980 1440
rect 32092 1440 32148 1442
rect 30924 1386 30980 1388
rect 32092 1388 32094 1440
rect 32094 1388 32146 1440
rect 32146 1388 32148 1440
rect 33260 1440 33316 1442
rect 32092 1386 32148 1388
rect 33260 1388 33262 1440
rect 33262 1388 33314 1440
rect 33314 1388 33316 1440
rect 34428 1440 34484 1442
rect 33260 1386 33316 1388
rect 34428 1388 34430 1440
rect 34430 1388 34482 1440
rect 34482 1388 34484 1440
rect 35596 1440 35652 1442
rect 34428 1386 34484 1388
rect 35596 1388 35598 1440
rect 35598 1388 35650 1440
rect 35650 1388 35652 1440
rect 36764 1440 36820 1442
rect 35596 1386 35652 1388
rect 36764 1388 36766 1440
rect 36766 1388 36818 1440
rect 36818 1388 36820 1440
rect 36764 1386 36820 1388
rect 368 280 424 336
rect 1536 280 1592 336
rect 2704 280 2760 336
rect 3872 280 3928 336
rect 5040 280 5096 336
rect 6208 280 6264 336
rect 7376 280 7432 336
rect 8544 280 8600 336
rect 9712 280 9768 336
rect 10880 280 10936 336
rect 12048 280 12104 336
rect 13216 280 13272 336
rect 14384 280 14440 336
rect 15552 280 15608 336
rect 16720 280 16776 336
rect 17888 280 17944 336
rect 19056 280 19112 336
rect 20224 280 20280 336
rect 21392 280 21448 336
rect 22560 280 22616 336
rect 23728 280 23784 336
rect 24896 280 24952 336
rect 26064 280 26120 336
rect 27232 280 27288 336
rect 28400 280 28456 336
rect 29568 280 29624 336
rect 30736 280 30792 336
rect 31904 280 31960 336
rect 33072 280 33128 336
rect 34240 280 34296 336
rect 35408 280 35464 336
rect 36576 280 36632 336
rect 556 26 612 28
rect 556 -26 558 26
rect 558 -26 610 26
rect 610 -26 612 26
rect 1724 26 1780 28
rect 556 -28 612 -26
rect 1724 -26 1726 26
rect 1726 -26 1778 26
rect 1778 -26 1780 26
rect 2892 26 2948 28
rect 1724 -28 1780 -26
rect 2892 -26 2894 26
rect 2894 -26 2946 26
rect 2946 -26 2948 26
rect 4060 26 4116 28
rect 2892 -28 2948 -26
rect 4060 -26 4062 26
rect 4062 -26 4114 26
rect 4114 -26 4116 26
rect 5228 26 5284 28
rect 4060 -28 4116 -26
rect 5228 -26 5230 26
rect 5230 -26 5282 26
rect 5282 -26 5284 26
rect 6396 26 6452 28
rect 5228 -28 5284 -26
rect 6396 -26 6398 26
rect 6398 -26 6450 26
rect 6450 -26 6452 26
rect 7564 26 7620 28
rect 6396 -28 6452 -26
rect 7564 -26 7566 26
rect 7566 -26 7618 26
rect 7618 -26 7620 26
rect 8732 26 8788 28
rect 7564 -28 7620 -26
rect 8732 -26 8734 26
rect 8734 -26 8786 26
rect 8786 -26 8788 26
rect 9900 26 9956 28
rect 8732 -28 8788 -26
rect 9900 -26 9902 26
rect 9902 -26 9954 26
rect 9954 -26 9956 26
rect 11068 26 11124 28
rect 9900 -28 9956 -26
rect 11068 -26 11070 26
rect 11070 -26 11122 26
rect 11122 -26 11124 26
rect 12236 26 12292 28
rect 11068 -28 11124 -26
rect 12236 -26 12238 26
rect 12238 -26 12290 26
rect 12290 -26 12292 26
rect 13404 26 13460 28
rect 12236 -28 12292 -26
rect 13404 -26 13406 26
rect 13406 -26 13458 26
rect 13458 -26 13460 26
rect 14572 26 14628 28
rect 13404 -28 13460 -26
rect 14572 -26 14574 26
rect 14574 -26 14626 26
rect 14626 -26 14628 26
rect 15740 26 15796 28
rect 14572 -28 14628 -26
rect 15740 -26 15742 26
rect 15742 -26 15794 26
rect 15794 -26 15796 26
rect 16908 26 16964 28
rect 15740 -28 15796 -26
rect 16908 -26 16910 26
rect 16910 -26 16962 26
rect 16962 -26 16964 26
rect 18076 26 18132 28
rect 16908 -28 16964 -26
rect 18076 -26 18078 26
rect 18078 -26 18130 26
rect 18130 -26 18132 26
rect 19244 26 19300 28
rect 18076 -28 18132 -26
rect 19244 -26 19246 26
rect 19246 -26 19298 26
rect 19298 -26 19300 26
rect 20412 26 20468 28
rect 19244 -28 19300 -26
rect 20412 -26 20414 26
rect 20414 -26 20466 26
rect 20466 -26 20468 26
rect 21580 26 21636 28
rect 20412 -28 20468 -26
rect 21580 -26 21582 26
rect 21582 -26 21634 26
rect 21634 -26 21636 26
rect 22748 26 22804 28
rect 21580 -28 21636 -26
rect 22748 -26 22750 26
rect 22750 -26 22802 26
rect 22802 -26 22804 26
rect 23916 26 23972 28
rect 22748 -28 22804 -26
rect 23916 -26 23918 26
rect 23918 -26 23970 26
rect 23970 -26 23972 26
rect 25084 26 25140 28
rect 23916 -28 23972 -26
rect 25084 -26 25086 26
rect 25086 -26 25138 26
rect 25138 -26 25140 26
rect 26252 26 26308 28
rect 25084 -28 25140 -26
rect 26252 -26 26254 26
rect 26254 -26 26306 26
rect 26306 -26 26308 26
rect 27420 26 27476 28
rect 26252 -28 26308 -26
rect 27420 -26 27422 26
rect 27422 -26 27474 26
rect 27474 -26 27476 26
rect 28588 26 28644 28
rect 27420 -28 27476 -26
rect 28588 -26 28590 26
rect 28590 -26 28642 26
rect 28642 -26 28644 26
rect 29756 26 29812 28
rect 28588 -28 28644 -26
rect 29756 -26 29758 26
rect 29758 -26 29810 26
rect 29810 -26 29812 26
rect 30924 26 30980 28
rect 29756 -28 29812 -26
rect 30924 -26 30926 26
rect 30926 -26 30978 26
rect 30978 -26 30980 26
rect 32092 26 32148 28
rect 30924 -28 30980 -26
rect 32092 -26 32094 26
rect 32094 -26 32146 26
rect 32146 -26 32148 26
rect 33260 26 33316 28
rect 32092 -28 32148 -26
rect 33260 -26 33262 26
rect 33262 -26 33314 26
rect 33314 -26 33316 26
rect 34428 26 34484 28
rect 33260 -28 33316 -26
rect 34428 -26 34430 26
rect 34430 -26 34482 26
rect 34482 -26 34484 26
rect 35596 26 35652 28
rect 34428 -28 34484 -26
rect 35596 -26 35598 26
rect 35598 -26 35650 26
rect 35650 -26 35652 26
rect 36764 26 36820 28
rect 35596 -28 35652 -26
rect 36764 -26 36766 26
rect 36766 -26 36818 26
rect 36818 -26 36820 26
rect 36764 -28 36820 -26
<< metal3 >>
rect 535 1442 633 1463
rect 535 1386 556 1442
rect 612 1386 633 1442
rect 535 1365 633 1386
rect 1703 1442 1801 1463
rect 1703 1386 1724 1442
rect 1780 1386 1801 1442
rect 1703 1365 1801 1386
rect 2871 1442 2969 1463
rect 2871 1386 2892 1442
rect 2948 1386 2969 1442
rect 2871 1365 2969 1386
rect 4039 1442 4137 1463
rect 4039 1386 4060 1442
rect 4116 1386 4137 1442
rect 4039 1365 4137 1386
rect 5207 1442 5305 1463
rect 5207 1386 5228 1442
rect 5284 1386 5305 1442
rect 5207 1365 5305 1386
rect 6375 1442 6473 1463
rect 6375 1386 6396 1442
rect 6452 1386 6473 1442
rect 6375 1365 6473 1386
rect 7543 1442 7641 1463
rect 7543 1386 7564 1442
rect 7620 1386 7641 1442
rect 7543 1365 7641 1386
rect 8711 1442 8809 1463
rect 8711 1386 8732 1442
rect 8788 1386 8809 1442
rect 8711 1365 8809 1386
rect 9879 1442 9977 1463
rect 9879 1386 9900 1442
rect 9956 1386 9977 1442
rect 9879 1365 9977 1386
rect 11047 1442 11145 1463
rect 11047 1386 11068 1442
rect 11124 1386 11145 1442
rect 11047 1365 11145 1386
rect 12215 1442 12313 1463
rect 12215 1386 12236 1442
rect 12292 1386 12313 1442
rect 12215 1365 12313 1386
rect 13383 1442 13481 1463
rect 13383 1386 13404 1442
rect 13460 1386 13481 1442
rect 13383 1365 13481 1386
rect 14551 1442 14649 1463
rect 14551 1386 14572 1442
rect 14628 1386 14649 1442
rect 14551 1365 14649 1386
rect 15719 1442 15817 1463
rect 15719 1386 15740 1442
rect 15796 1386 15817 1442
rect 15719 1365 15817 1386
rect 16887 1442 16985 1463
rect 16887 1386 16908 1442
rect 16964 1386 16985 1442
rect 16887 1365 16985 1386
rect 18055 1442 18153 1463
rect 18055 1386 18076 1442
rect 18132 1386 18153 1442
rect 18055 1365 18153 1386
rect 19223 1442 19321 1463
rect 19223 1386 19244 1442
rect 19300 1386 19321 1442
rect 19223 1365 19321 1386
rect 20391 1442 20489 1463
rect 20391 1386 20412 1442
rect 20468 1386 20489 1442
rect 20391 1365 20489 1386
rect 21559 1442 21657 1463
rect 21559 1386 21580 1442
rect 21636 1386 21657 1442
rect 21559 1365 21657 1386
rect 22727 1442 22825 1463
rect 22727 1386 22748 1442
rect 22804 1386 22825 1442
rect 22727 1365 22825 1386
rect 23895 1442 23993 1463
rect 23895 1386 23916 1442
rect 23972 1386 23993 1442
rect 23895 1365 23993 1386
rect 25063 1442 25161 1463
rect 25063 1386 25084 1442
rect 25140 1386 25161 1442
rect 25063 1365 25161 1386
rect 26231 1442 26329 1463
rect 26231 1386 26252 1442
rect 26308 1386 26329 1442
rect 26231 1365 26329 1386
rect 27399 1442 27497 1463
rect 27399 1386 27420 1442
rect 27476 1386 27497 1442
rect 27399 1365 27497 1386
rect 28567 1442 28665 1463
rect 28567 1386 28588 1442
rect 28644 1386 28665 1442
rect 28567 1365 28665 1386
rect 29735 1442 29833 1463
rect 29735 1386 29756 1442
rect 29812 1386 29833 1442
rect 29735 1365 29833 1386
rect 30903 1442 31001 1463
rect 30903 1386 30924 1442
rect 30980 1386 31001 1442
rect 30903 1365 31001 1386
rect 32071 1442 32169 1463
rect 32071 1386 32092 1442
rect 32148 1386 32169 1442
rect 32071 1365 32169 1386
rect 33239 1442 33337 1463
rect 33239 1386 33260 1442
rect 33316 1386 33337 1442
rect 33239 1365 33337 1386
rect 34407 1442 34505 1463
rect 34407 1386 34428 1442
rect 34484 1386 34505 1442
rect 34407 1365 34505 1386
rect 35575 1442 35673 1463
rect 35575 1386 35596 1442
rect 35652 1386 35673 1442
rect 35575 1365 35673 1386
rect 36743 1442 36841 1463
rect 36743 1386 36764 1442
rect 36820 1386 36841 1442
rect 36743 1365 36841 1386
rect 363 338 429 341
rect 1531 338 1597 341
rect 2699 338 2765 341
rect 3867 338 3933 341
rect 5035 338 5101 341
rect 6203 338 6269 341
rect 7371 338 7437 341
rect 8539 338 8605 341
rect 9707 338 9773 341
rect 10875 338 10941 341
rect 12043 338 12109 341
rect 13211 338 13277 341
rect 14379 338 14445 341
rect 15547 338 15613 341
rect 16715 338 16781 341
rect 17883 338 17949 341
rect 19051 338 19117 341
rect 20219 338 20285 341
rect 21387 338 21453 341
rect 22555 338 22621 341
rect 23723 338 23789 341
rect 24891 338 24957 341
rect 26059 338 26125 341
rect 27227 338 27293 341
rect 28395 338 28461 341
rect 29563 338 29629 341
rect 30731 338 30797 341
rect 31899 338 31965 341
rect 33067 338 33133 341
rect 34235 338 34301 341
rect 35403 338 35469 341
rect 36571 338 36637 341
rect 0 336 37376 338
rect 0 280 368 336
rect 424 280 1536 336
rect 1592 280 2704 336
rect 2760 280 3872 336
rect 3928 280 5040 336
rect 5096 280 6208 336
rect 6264 280 7376 336
rect 7432 280 8544 336
rect 8600 280 9712 336
rect 9768 280 10880 336
rect 10936 280 12048 336
rect 12104 280 13216 336
rect 13272 280 14384 336
rect 14440 280 15552 336
rect 15608 280 16720 336
rect 16776 280 17888 336
rect 17944 280 19056 336
rect 19112 280 20224 336
rect 20280 280 21392 336
rect 21448 280 22560 336
rect 22616 280 23728 336
rect 23784 280 24896 336
rect 24952 280 26064 336
rect 26120 280 27232 336
rect 27288 280 28400 336
rect 28456 280 29568 336
rect 29624 280 30736 336
rect 30792 280 31904 336
rect 31960 280 33072 336
rect 33128 280 34240 336
rect 34296 280 35408 336
rect 35464 280 36576 336
rect 36632 280 37376 336
rect 0 278 37376 280
rect 363 275 429 278
rect 1531 275 1597 278
rect 2699 275 2765 278
rect 3867 275 3933 278
rect 5035 275 5101 278
rect 6203 275 6269 278
rect 7371 275 7437 278
rect 8539 275 8605 278
rect 9707 275 9773 278
rect 10875 275 10941 278
rect 12043 275 12109 278
rect 13211 275 13277 278
rect 14379 275 14445 278
rect 15547 275 15613 278
rect 16715 275 16781 278
rect 17883 275 17949 278
rect 19051 275 19117 278
rect 20219 275 20285 278
rect 21387 275 21453 278
rect 22555 275 22621 278
rect 23723 275 23789 278
rect 24891 275 24957 278
rect 26059 275 26125 278
rect 27227 275 27293 278
rect 28395 275 28461 278
rect 29563 275 29629 278
rect 30731 275 30797 278
rect 31899 275 31965 278
rect 33067 275 33133 278
rect 34235 275 34301 278
rect 35403 275 35469 278
rect 36571 275 36637 278
rect 535 28 633 49
rect 535 -28 556 28
rect 612 -28 633 28
rect 535 -49 633 -28
rect 1703 28 1801 49
rect 1703 -28 1724 28
rect 1780 -28 1801 28
rect 1703 -49 1801 -28
rect 2871 28 2969 49
rect 2871 -28 2892 28
rect 2948 -28 2969 28
rect 2871 -49 2969 -28
rect 4039 28 4137 49
rect 4039 -28 4060 28
rect 4116 -28 4137 28
rect 4039 -49 4137 -28
rect 5207 28 5305 49
rect 5207 -28 5228 28
rect 5284 -28 5305 28
rect 5207 -49 5305 -28
rect 6375 28 6473 49
rect 6375 -28 6396 28
rect 6452 -28 6473 28
rect 6375 -49 6473 -28
rect 7543 28 7641 49
rect 7543 -28 7564 28
rect 7620 -28 7641 28
rect 7543 -49 7641 -28
rect 8711 28 8809 49
rect 8711 -28 8732 28
rect 8788 -28 8809 28
rect 8711 -49 8809 -28
rect 9879 28 9977 49
rect 9879 -28 9900 28
rect 9956 -28 9977 28
rect 9879 -49 9977 -28
rect 11047 28 11145 49
rect 11047 -28 11068 28
rect 11124 -28 11145 28
rect 11047 -49 11145 -28
rect 12215 28 12313 49
rect 12215 -28 12236 28
rect 12292 -28 12313 28
rect 12215 -49 12313 -28
rect 13383 28 13481 49
rect 13383 -28 13404 28
rect 13460 -28 13481 28
rect 13383 -49 13481 -28
rect 14551 28 14649 49
rect 14551 -28 14572 28
rect 14628 -28 14649 28
rect 14551 -49 14649 -28
rect 15719 28 15817 49
rect 15719 -28 15740 28
rect 15796 -28 15817 28
rect 15719 -49 15817 -28
rect 16887 28 16985 49
rect 16887 -28 16908 28
rect 16964 -28 16985 28
rect 16887 -49 16985 -28
rect 18055 28 18153 49
rect 18055 -28 18076 28
rect 18132 -28 18153 28
rect 18055 -49 18153 -28
rect 19223 28 19321 49
rect 19223 -28 19244 28
rect 19300 -28 19321 28
rect 19223 -49 19321 -28
rect 20391 28 20489 49
rect 20391 -28 20412 28
rect 20468 -28 20489 28
rect 20391 -49 20489 -28
rect 21559 28 21657 49
rect 21559 -28 21580 28
rect 21636 -28 21657 28
rect 21559 -49 21657 -28
rect 22727 28 22825 49
rect 22727 -28 22748 28
rect 22804 -28 22825 28
rect 22727 -49 22825 -28
rect 23895 28 23993 49
rect 23895 -28 23916 28
rect 23972 -28 23993 28
rect 23895 -49 23993 -28
rect 25063 28 25161 49
rect 25063 -28 25084 28
rect 25140 -28 25161 28
rect 25063 -49 25161 -28
rect 26231 28 26329 49
rect 26231 -28 26252 28
rect 26308 -28 26329 28
rect 26231 -49 26329 -28
rect 27399 28 27497 49
rect 27399 -28 27420 28
rect 27476 -28 27497 28
rect 27399 -49 27497 -28
rect 28567 28 28665 49
rect 28567 -28 28588 28
rect 28644 -28 28665 28
rect 28567 -49 28665 -28
rect 29735 28 29833 49
rect 29735 -28 29756 28
rect 29812 -28 29833 28
rect 29735 -49 29833 -28
rect 30903 28 31001 49
rect 30903 -28 30924 28
rect 30980 -28 31001 28
rect 30903 -49 31001 -28
rect 32071 28 32169 49
rect 32071 -28 32092 28
rect 32148 -28 32169 28
rect 32071 -49 32169 -28
rect 33239 28 33337 49
rect 33239 -28 33260 28
rect 33316 -28 33337 28
rect 33239 -49 33337 -28
rect 34407 28 34505 49
rect 34407 -28 34428 28
rect 34484 -28 34505 28
rect 34407 -49 34505 -28
rect 35575 28 35673 49
rect 35575 -28 35596 28
rect 35652 -28 35673 28
rect 35575 -49 35673 -28
rect 36743 28 36841 49
rect 36743 -28 36764 28
rect 36820 -28 36841 28
rect 36743 -49 36841 -28
use contact_7  contact_7_0
timestamp 1701704242
transform 1 0 555 0 1 -33
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1701704242
transform 1 0 7563 0 1 -33
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1701704242
transform 1 0 1723 0 1 -33
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1701704242
transform 1 0 2891 0 1 -33
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1701704242
transform 1 0 5227 0 1 -33
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1701704242
transform 1 0 8731 0 1 -33
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1701704242
transform 1 0 8731 0 1 1381
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1701704242
transform 1 0 7563 0 1 1381
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1701704242
transform 1 0 6395 0 1 1381
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1701704242
transform 1 0 5227 0 1 1381
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1701704242
transform 1 0 4059 0 1 1381
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1701704242
transform 1 0 2891 0 1 1381
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1701704242
transform 1 0 1723 0 1 1381
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1701704242
transform 1 0 555 0 1 1381
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1701704242
transform 1 0 4059 0 1 -33
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1701704242
transform 1 0 6395 0 1 -33
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1701704242
transform 1 0 18075 0 1 1381
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1701704242
transform 1 0 16907 0 1 1381
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1701704242
transform 1 0 15739 0 1 1381
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1701704242
transform 1 0 14571 0 1 1381
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1701704242
transform 1 0 13403 0 1 1381
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1701704242
transform 1 0 12235 0 1 1381
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1701704242
transform 1 0 11067 0 1 1381
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1701704242
transform 1 0 9899 0 1 1381
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1701704242
transform 1 0 9899 0 1 -33
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1701704242
transform 1 0 18075 0 1 -33
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1701704242
transform 1 0 16907 0 1 -33
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1701704242
transform 1 0 15739 0 1 -33
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1701704242
transform 1 0 14571 0 1 -33
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1701704242
transform 1 0 13403 0 1 -33
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1701704242
transform 1 0 12235 0 1 -33
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1701704242
transform 1 0 11067 0 1 -33
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1701704242
transform 1 0 26251 0 1 1381
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1701704242
transform 1 0 25083 0 1 1381
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1701704242
transform 1 0 23915 0 1 1381
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1701704242
transform 1 0 21579 0 1 -33
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1701704242
transform 1 0 22747 0 1 1381
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1701704242
transform 1 0 23915 0 1 -33
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1701704242
transform 1 0 21579 0 1 1381
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1701704242
transform 1 0 19243 0 1 -33
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1701704242
transform 1 0 20411 0 1 1381
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1701704242
transform 1 0 27419 0 1 -33
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1701704242
transform 1 0 19243 0 1 1381
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1701704242
transform 1 0 22747 0 1 -33
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1701704242
transform 1 0 26251 0 1 -33
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1701704242
transform 1 0 20411 0 1 -33
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1701704242
transform 1 0 27419 0 1 1381
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1701704242
transform 1 0 25083 0 1 -33
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1701704242
transform 1 0 30923 0 1 -33
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1701704242
transform 1 0 29755 0 1 -33
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1701704242
transform 1 0 28587 0 1 -33
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1701704242
transform 1 0 36763 0 1 -33
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1701704242
transform 1 0 35595 0 1 -33
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1701704242
transform 1 0 34427 0 1 -33
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1701704242
transform 1 0 33259 0 1 -33
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1701704242
transform 1 0 32091 0 1 -33
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1701704242
transform 1 0 36763 0 1 1381
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1701704242
transform 1 0 35595 0 1 1381
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1701704242
transform 1 0 34427 0 1 1381
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1701704242
transform 1 0 33259 0 1 1381
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1701704242
transform 1 0 32091 0 1 1381
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1701704242
transform 1 0 30923 0 1 1381
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1701704242
transform 1 0 29755 0 1 1381
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1701704242
transform 1 0 28587 0 1 1381
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1701704242
transform 1 0 7560 0 1 -32
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1701704242
transform 1 0 5224 0 1 -32
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1701704242
transform 1 0 2888 0 1 -32
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1701704242
transform 1 0 1720 0 1 -32
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1701704242
transform 1 0 8728 0 1 -32
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1701704242
transform 1 0 552 0 1 -32
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1701704242
transform 1 0 8728 0 1 1382
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1701704242
transform 1 0 7560 0 1 1382
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1701704242
transform 1 0 6392 0 1 1382
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1701704242
transform 1 0 5224 0 1 1382
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1701704242
transform 1 0 4056 0 1 1382
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1701704242
transform 1 0 2888 0 1 1382
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1701704242
transform 1 0 1720 0 1 1382
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1701704242
transform 1 0 552 0 1 1382
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1701704242
transform 1 0 6392 0 1 -32
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1701704242
transform 1 0 4056 0 1 -32
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1701704242
transform 1 0 18072 0 1 1382
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1701704242
transform 1 0 16904 0 1 1382
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1701704242
transform 1 0 15736 0 1 1382
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1701704242
transform 1 0 14568 0 1 1382
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1701704242
transform 1 0 13400 0 1 1382
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1701704242
transform 1 0 12232 0 1 1382
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1701704242
transform 1 0 11064 0 1 1382
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1701704242
transform 1 0 9896 0 1 1382
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1701704242
transform 1 0 9896 0 1 -32
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1701704242
transform 1 0 18072 0 1 -32
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1701704242
transform 1 0 16904 0 1 -32
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1701704242
transform 1 0 15736 0 1 -32
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1701704242
transform 1 0 14568 0 1 -32
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1701704242
transform 1 0 13400 0 1 -32
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1701704242
transform 1 0 12232 0 1 -32
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1701704242
transform 1 0 11064 0 1 -32
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1701704242
transform 1 0 26248 0 1 1382
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1701704242
transform 1 0 25080 0 1 1382
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1701704242
transform 1 0 23912 0 1 1382
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1701704242
transform 1 0 21576 0 1 -32
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1701704242
transform 1 0 22744 0 1 1382
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1701704242
transform 1 0 23912 0 1 -32
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1701704242
transform 1 0 21576 0 1 1382
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1701704242
transform 1 0 19240 0 1 -32
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1701704242
transform 1 0 20408 0 1 1382
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1701704242
transform 1 0 27416 0 1 -32
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1701704242
transform 1 0 19240 0 1 1382
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1701704242
transform 1 0 22744 0 1 -32
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1701704242
transform 1 0 26248 0 1 -32
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1701704242
transform 1 0 20408 0 1 -32
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1701704242
transform 1 0 27416 0 1 1382
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1701704242
transform 1 0 25080 0 1 -32
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1701704242
transform 1 0 29752 0 1 -32
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1701704242
transform 1 0 28584 0 1 -32
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1701704242
transform 1 0 36760 0 1 -32
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1701704242
transform 1 0 35592 0 1 -32
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1701704242
transform 1 0 34424 0 1 -32
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1701704242
transform 1 0 33256 0 1 -32
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1701704242
transform 1 0 32088 0 1 -32
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1701704242
transform 1 0 30920 0 1 -32
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1701704242
transform 1 0 36760 0 1 1382
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1701704242
transform 1 0 35592 0 1 1382
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1701704242
transform 1 0 34424 0 1 1382
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1701704242
transform 1 0 33256 0 1 1382
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1701704242
transform 1 0 32088 0 1 1382
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1701704242
transform 1 0 30920 0 1 1382
box 0 0 1 1
use contact_8  contact_8_62
timestamp 1701704242
transform 1 0 29752 0 1 1382
box 0 0 1 1
use contact_8  contact_8_63
timestamp 1701704242
transform 1 0 28584 0 1 1382
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1701704242
transform 1 0 7559 0 1 -37
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1701704242
transform 1 0 2887 0 1 -37
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1701704242
transform 1 0 1719 0 1 -37
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1701704242
transform 1 0 8539 0 1 271
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1701704242
transform 1 0 7371 0 1 271
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1701704242
transform 1 0 6203 0 1 271
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1701704242
transform 1 0 5035 0 1 271
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1701704242
transform 1 0 3867 0 1 271
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1701704242
transform 1 0 2699 0 1 271
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1701704242
transform 1 0 1531 0 1 271
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1701704242
transform 1 0 363 0 1 271
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1701704242
transform 1 0 8727 0 1 -37
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1701704242
transform 1 0 8727 0 1 1377
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1701704242
transform 1 0 7559 0 1 1377
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1701704242
transform 1 0 6391 0 1 1377
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1701704242
transform 1 0 5223 0 1 1377
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1701704242
transform 1 0 4055 0 1 1377
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1701704242
transform 1 0 2887 0 1 1377
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1701704242
transform 1 0 1719 0 1 1377
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1701704242
transform 1 0 551 0 1 1377
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1701704242
transform 1 0 6391 0 1 -37
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1701704242
transform 1 0 4055 0 1 -37
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1701704242
transform 1 0 551 0 1 -37
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1701704242
transform 1 0 5223 0 1 -37
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1701704242
transform 1 0 18071 0 1 1377
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1701704242
transform 1 0 16903 0 1 1377
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1701704242
transform 1 0 15735 0 1 1377
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1701704242
transform 1 0 14567 0 1 1377
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1701704242
transform 1 0 13399 0 1 1377
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1701704242
transform 1 0 12231 0 1 1377
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1701704242
transform 1 0 11063 0 1 1377
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1701704242
transform 1 0 9895 0 1 1377
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1701704242
transform 1 0 17883 0 1 271
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1701704242
transform 1 0 16715 0 1 271
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1701704242
transform 1 0 15547 0 1 271
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1701704242
transform 1 0 14379 0 1 271
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1701704242
transform 1 0 13211 0 1 271
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1701704242
transform 1 0 12043 0 1 271
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1701704242
transform 1 0 10875 0 1 271
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1701704242
transform 1 0 9707 0 1 271
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1701704242
transform 1 0 18071 0 1 -37
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1701704242
transform 1 0 16903 0 1 -37
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1701704242
transform 1 0 15735 0 1 -37
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1701704242
transform 1 0 14567 0 1 -37
box 0 0 1 1
use contact_9  contact_9_44
timestamp 1701704242
transform 1 0 13399 0 1 -37
box 0 0 1 1
use contact_9  contact_9_45
timestamp 1701704242
transform 1 0 12231 0 1 -37
box 0 0 1 1
use contact_9  contact_9_46
timestamp 1701704242
transform 1 0 11063 0 1 -37
box 0 0 1 1
use contact_9  contact_9_47
timestamp 1701704242
transform 1 0 9895 0 1 -37
box 0 0 1 1
use contact_9  contact_9_48
timestamp 1701704242
transform 1 0 25079 0 1 1377
box 0 0 1 1
use contact_9  contact_9_49
timestamp 1701704242
transform 1 0 23911 0 1 1377
box 0 0 1 1
use contact_9  contact_9_50
timestamp 1701704242
transform 1 0 27227 0 1 271
box 0 0 1 1
use contact_9  contact_9_51
timestamp 1701704242
transform 1 0 26059 0 1 271
box 0 0 1 1
use contact_9  contact_9_52
timestamp 1701704242
transform 1 0 24891 0 1 271
box 0 0 1 1
use contact_9  contact_9_53
timestamp 1701704242
transform 1 0 23723 0 1 271
box 0 0 1 1
use contact_9  contact_9_54
timestamp 1701704242
transform 1 0 22555 0 1 271
box 0 0 1 1
use contact_9  contact_9_55
timestamp 1701704242
transform 1 0 21387 0 1 271
box 0 0 1 1
use contact_9  contact_9_56
timestamp 1701704242
transform 1 0 20219 0 1 271
box 0 0 1 1
use contact_9  contact_9_57
timestamp 1701704242
transform 1 0 19051 0 1 271
box 0 0 1 1
use contact_9  contact_9_58
timestamp 1701704242
transform 1 0 22743 0 1 1377
box 0 0 1 1
use contact_9  contact_9_59
timestamp 1701704242
transform 1 0 21575 0 1 -37
box 0 0 1 1
use contact_9  contact_9_60
timestamp 1701704242
transform 1 0 21575 0 1 1377
box 0 0 1 1
use contact_9  contact_9_61
timestamp 1701704242
transform 1 0 23911 0 1 -37
box 0 0 1 1
use contact_9  contact_9_62
timestamp 1701704242
transform 1 0 20407 0 1 1377
box 0 0 1 1
use contact_9  contact_9_63
timestamp 1701704242
transform 1 0 19239 0 1 -37
box 0 0 1 1
use contact_9  contact_9_64
timestamp 1701704242
transform 1 0 19239 0 1 1377
box 0 0 1 1
use contact_9  contact_9_65
timestamp 1701704242
transform 1 0 27415 0 1 -37
box 0 0 1 1
use contact_9  contact_9_66
timestamp 1701704242
transform 1 0 22743 0 1 -37
box 0 0 1 1
use contact_9  contact_9_67
timestamp 1701704242
transform 1 0 26247 0 1 -37
box 0 0 1 1
use contact_9  contact_9_68
timestamp 1701704242
transform 1 0 27415 0 1 1377
box 0 0 1 1
use contact_9  contact_9_69
timestamp 1701704242
transform 1 0 20407 0 1 -37
box 0 0 1 1
use contact_9  contact_9_70
timestamp 1701704242
transform 1 0 26247 0 1 1377
box 0 0 1 1
use contact_9  contact_9_71
timestamp 1701704242
transform 1 0 25079 0 1 -37
box 0 0 1 1
use contact_9  contact_9_72
timestamp 1701704242
transform 1 0 36571 0 1 271
box 0 0 1 1
use contact_9  contact_9_73
timestamp 1701704242
transform 1 0 35403 0 1 271
box 0 0 1 1
use contact_9  contact_9_74
timestamp 1701704242
transform 1 0 34235 0 1 271
box 0 0 1 1
use contact_9  contact_9_75
timestamp 1701704242
transform 1 0 33067 0 1 271
box 0 0 1 1
use contact_9  contact_9_76
timestamp 1701704242
transform 1 0 31899 0 1 271
box 0 0 1 1
use contact_9  contact_9_77
timestamp 1701704242
transform 1 0 30731 0 1 271
box 0 0 1 1
use contact_9  contact_9_78
timestamp 1701704242
transform 1 0 29563 0 1 271
box 0 0 1 1
use contact_9  contact_9_79
timestamp 1701704242
transform 1 0 28395 0 1 271
box 0 0 1 1
use contact_9  contact_9_80
timestamp 1701704242
transform 1 0 29751 0 1 -37
box 0 0 1 1
use contact_9  contact_9_81
timestamp 1701704242
transform 1 0 28583 0 1 -37
box 0 0 1 1
use contact_9  contact_9_82
timestamp 1701704242
transform 1 0 36759 0 1 -37
box 0 0 1 1
use contact_9  contact_9_83
timestamp 1701704242
transform 1 0 35591 0 1 -37
box 0 0 1 1
use contact_9  contact_9_84
timestamp 1701704242
transform 1 0 34423 0 1 -37
box 0 0 1 1
use contact_9  contact_9_85
timestamp 1701704242
transform 1 0 33255 0 1 -37
box 0 0 1 1
use contact_9  contact_9_86
timestamp 1701704242
transform 1 0 32087 0 1 -37
box 0 0 1 1
use contact_9  contact_9_87
timestamp 1701704242
transform 1 0 30919 0 1 -37
box 0 0 1 1
use contact_9  contact_9_88
timestamp 1701704242
transform 1 0 36759 0 1 1377
box 0 0 1 1
use contact_9  contact_9_89
timestamp 1701704242
transform 1 0 35591 0 1 1377
box 0 0 1 1
use contact_9  contact_9_90
timestamp 1701704242
transform 1 0 34423 0 1 1377
box 0 0 1 1
use contact_9  contact_9_91
timestamp 1701704242
transform 1 0 33255 0 1 1377
box 0 0 1 1
use contact_9  contact_9_92
timestamp 1701704242
transform 1 0 32087 0 1 1377
box 0 0 1 1
use contact_9  contact_9_93
timestamp 1701704242
transform 1 0 30919 0 1 1377
box 0 0 1 1
use contact_9  contact_9_94
timestamp 1701704242
transform 1 0 29751 0 1 1377
box 0 0 1 1
use contact_9  contact_9_95
timestamp 1701704242
transform 1 0 28583 0 1 1377
box 0 0 1 1
use dff  dff_0
timestamp 1701704242
transform 1 0 5840 0 1 0
box -8 -43 1176 1467
use dff  dff_1
timestamp 1701704242
transform 1 0 4672 0 1 0
box -8 -43 1176 1467
use dff  dff_2
timestamp 1701704242
transform 1 0 3504 0 1 0
box -8 -43 1176 1467
use dff  dff_3
timestamp 1701704242
transform 1 0 2336 0 1 0
box -8 -43 1176 1467
use dff  dff_4
timestamp 1701704242
transform 1 0 1168 0 1 0
box -8 -43 1176 1467
use dff  dff_5
timestamp 1701704242
transform 1 0 0 0 1 0
box -8 -43 1176 1467
use dff  dff_6
timestamp 1701704242
transform 1 0 7008 0 1 0
box -8 -43 1176 1467
use dff  dff_7
timestamp 1701704242
transform 1 0 16352 0 1 0
box -8 -43 1176 1467
use dff  dff_8
timestamp 1701704242
transform 1 0 15184 0 1 0
box -8 -43 1176 1467
use dff  dff_9
timestamp 1701704242
transform 1 0 14016 0 1 0
box -8 -43 1176 1467
use dff  dff_10
timestamp 1701704242
transform 1 0 12848 0 1 0
box -8 -43 1176 1467
use dff  dff_11
timestamp 1701704242
transform 1 0 11680 0 1 0
box -8 -43 1176 1467
use dff  dff_12
timestamp 1701704242
transform 1 0 10512 0 1 0
box -8 -43 1176 1467
use dff  dff_13
timestamp 1701704242
transform 1 0 9344 0 1 0
box -8 -43 1176 1467
use dff  dff_14
timestamp 1701704242
transform 1 0 8176 0 1 0
box -8 -43 1176 1467
use dff  dff_15
timestamp 1701704242
transform 1 0 22192 0 1 0
box -8 -43 1176 1467
use dff  dff_16
timestamp 1701704242
transform 1 0 21024 0 1 0
box -8 -43 1176 1467
use dff  dff_17
timestamp 1701704242
transform 1 0 19856 0 1 0
box -8 -43 1176 1467
use dff  dff_18
timestamp 1701704242
transform 1 0 25696 0 1 0
box -8 -43 1176 1467
use dff  dff_19
timestamp 1701704242
transform 1 0 24528 0 1 0
box -8 -43 1176 1467
use dff  dff_20
timestamp 1701704242
transform 1 0 23360 0 1 0
box -8 -43 1176 1467
use dff  dff_21
timestamp 1701704242
transform 1 0 36208 0 1 0
box -8 -43 1176 1467
use dff  dff_22
timestamp 1701704242
transform 1 0 35040 0 1 0
box -8 -43 1176 1467
use dff  dff_23
timestamp 1701704242
transform 1 0 33872 0 1 0
box -8 -43 1176 1467
use dff  dff_24
timestamp 1701704242
transform 1 0 32704 0 1 0
box -8 -43 1176 1467
use dff  dff_25
timestamp 1701704242
transform 1 0 31536 0 1 0
box -8 -43 1176 1467
use dff  dff_26
timestamp 1701704242
transform 1 0 30368 0 1 0
box -8 -43 1176 1467
use dff  dff_27
timestamp 1701704242
transform 1 0 29200 0 1 0
box -8 -43 1176 1467
use dff  dff_28
timestamp 1701704242
transform 1 0 28032 0 1 0
box -8 -43 1176 1467
use dff  dff_29
timestamp 1701704242
transform 1 0 26864 0 1 0
box -8 -43 1176 1467
use dff  dff_30
timestamp 1701704242
transform 1 0 18688 0 1 0
box -8 -43 1176 1467
use dff  dff_31
timestamp 1701704242
transform 1 0 17520 0 1 0
box -8 -43 1176 1467
<< labels >>
rlabel metal2 s 23530 564 23530 564 4 din_20
port 21 nsew
rlabel metal2 s 23307 635 23307 635 4 dout_19
port 52 nsew
rlabel metal2 s 1115 635 1115 635 4 dout_0
port 33 nsew
rlabel metal2 s 34042 564 34042 564 4 din_29
port 30 nsew
rlabel metal2 s 9291 635 9291 635 4 dout_7
port 40 nsew
rlabel metal2 s 24698 564 24698 564 4 din_21
port 22 nsew
rlabel metal2 s 3674 564 3674 564 4 din_3
port 4 nsew
rlabel metal2 s 27034 564 27034 564 4 din_23
port 24 nsew
rlabel metal2 s 18858 564 18858 564 4 din_16
port 17 nsew
rlabel metal2 s 29370 564 29370 564 4 din_25
port 26 nsew
rlabel metal2 s 10682 564 10682 564 4 din_9
port 10 nsew
rlabel metal2 s 24475 635 24475 635 4 dout_20
port 53 nsew
rlabel metal2 s 8346 564 8346 564 4 din_7
port 8 nsew
rlabel metal2 s 2283 635 2283 635 4 dout_1
port 34 nsew
rlabel metal2 s 8123 635 8123 635 4 dout_6
port 39 nsew
rlabel metal2 s 13963 635 13963 635 4 dout_11
port 44 nsew
rlabel metal2 s 10459 635 10459 635 4 dout_8
port 41 nsew
rlabel metal2 s 17690 564 17690 564 4 din_15
port 16 nsew
rlabel metal2 s 37323 635 37323 635 4 dout_31
port 64 nsew
rlabel metal2 s 15131 635 15131 635 4 dout_12
port 45 nsew
rlabel metal2 s 19803 635 19803 635 4 dout_16
port 49 nsew
rlabel metal2 s 36155 635 36155 635 4 dout_30
port 63 nsew
rlabel metal2 s 27979 635 27979 635 4 dout_23
port 56 nsew
rlabel metal2 s 2506 564 2506 564 4 din_2
port 3 nsew
rlabel metal2 s 33819 635 33819 635 4 dout_28
port 61 nsew
rlabel metal2 s 25866 564 25866 564 4 din_22
port 23 nsew
rlabel metal2 s 25643 635 25643 635 4 dout_21
port 54 nsew
rlabel metal2 s 30315 635 30315 635 4 dout_25
port 58 nsew
rlabel metal2 s 32874 564 32874 564 4 din_28
port 29 nsew
rlabel metal2 s 9514 564 9514 564 4 din_8
port 9 nsew
rlabel metal2 s 6955 635 6955 635 4 dout_5
port 38 nsew
rlabel metal2 s 32651 635 32651 635 4 dout_27
port 60 nsew
rlabel metal2 s 4619 635 4619 635 4 dout_3
port 36 nsew
rlabel metal2 s 31483 635 31483 635 4 dout_26
port 59 nsew
rlabel metal2 s 28202 564 28202 564 4 din_24
port 25 nsew
rlabel metal2 s 15354 564 15354 564 4 din_13
port 14 nsew
rlabel metal2 s 20026 564 20026 564 4 din_17
port 18 nsew
rlabel metal2 s 22139 635 22139 635 4 dout_18
port 51 nsew
rlabel metal2 s 14186 564 14186 564 4 din_12
port 13 nsew
rlabel metal2 s 16522 564 16522 564 4 din_14
port 15 nsew
rlabel metal2 s 1338 564 1338 564 4 din_1
port 2 nsew
rlabel metal2 s 12795 635 12795 635 4 dout_10
port 43 nsew
rlabel metal2 s 26811 635 26811 635 4 dout_22
port 55 nsew
rlabel metal2 s 7178 564 7178 564 4 din_6
port 7 nsew
rlabel metal2 s 29147 635 29147 635 4 dout_24
port 57 nsew
rlabel metal2 s 3451 635 3451 635 4 dout_2
port 35 nsew
rlabel metal2 s 5787 635 5787 635 4 dout_4
port 37 nsew
rlabel metal2 s 13018 564 13018 564 4 din_11
port 12 nsew
rlabel metal2 s 31706 564 31706 564 4 din_27
port 28 nsew
rlabel metal2 s 18635 635 18635 635 4 dout_15
port 48 nsew
rlabel metal2 s 21194 564 21194 564 4 din_18
port 19 nsew
rlabel metal2 s 170 564 170 564 4 din_0
port 1 nsew
rlabel metal2 s 11850 564 11850 564 4 din_10
port 11 nsew
rlabel metal2 s 35210 564 35210 564 4 din_30
port 31 nsew
rlabel metal2 s 36378 564 36378 564 4 din_31
port 32 nsew
rlabel metal2 s 17467 635 17467 635 4 dout_14
port 47 nsew
rlabel metal2 s 4842 564 4842 564 4 din_4
port 5 nsew
rlabel metal2 s 6010 564 6010 564 4 din_5
port 6 nsew
rlabel metal2 s 16299 635 16299 635 4 dout_13
port 46 nsew
rlabel metal2 s 11627 635 11627 635 4 dout_9
port 42 nsew
rlabel metal2 s 22362 564 22362 564 4 din_19
port 20 nsew
rlabel metal2 s 34987 635 34987 635 4 dout_29
port 62 nsew
rlabel metal2 s 20971 635 20971 635 4 dout_17
port 50 nsew
rlabel metal2 s 30538 564 30538 564 4 din_26
port 27 nsew
rlabel metal3 s 7592 1414 7592 1414 4 vdd
port 66 nsew
rlabel metal3 s 6424 1414 6424 1414 4 vdd
port 66 nsew
rlabel metal3 s 34456 1414 34456 1414 4 vdd
port 66 nsew
rlabel metal3 s 584 1414 584 1414 4 vdd
port 66 nsew
rlabel metal3 s 1752 1414 1752 1414 4 vdd
port 66 nsew
rlabel metal3 s 21608 1414 21608 1414 4 vdd
port 66 nsew
rlabel metal3 s 2920 1414 2920 1414 4 vdd
port 66 nsew
rlabel metal3 s 14600 1414 14600 1414 4 vdd
port 66 nsew
rlabel metal3 s 27448 1414 27448 1414 4 vdd
port 66 nsew
rlabel metal3 s 18104 1414 18104 1414 4 vdd
port 66 nsew
rlabel metal3 s 13432 1414 13432 1414 4 vdd
port 66 nsew
rlabel metal3 s 4088 1414 4088 1414 4 vdd
port 66 nsew
rlabel metal3 s 11096 1414 11096 1414 4 vdd
port 66 nsew
rlabel metal3 s 19272 1414 19272 1414 4 vdd
port 66 nsew
rlabel metal3 s 9928 1414 9928 1414 4 vdd
port 66 nsew
rlabel metal3 s 5256 1414 5256 1414 4 vdd
port 66 nsew
rlabel metal3 s 15768 1414 15768 1414 4 vdd
port 66 nsew
rlabel metal3 s 26280 1414 26280 1414 4 vdd
port 66 nsew
rlabel metal3 s 16936 1414 16936 1414 4 vdd
port 66 nsew
rlabel metal3 s 12264 1414 12264 1414 4 vdd
port 66 nsew
rlabel metal3 s 30952 1414 30952 1414 4 vdd
port 66 nsew
rlabel metal3 s 28616 1414 28616 1414 4 vdd
port 66 nsew
rlabel metal3 s 35624 1414 35624 1414 4 vdd
port 66 nsew
rlabel metal3 s 23944 1414 23944 1414 4 vdd
port 66 nsew
rlabel metal3 s 8760 1414 8760 1414 4 vdd
port 66 nsew
rlabel metal3 s 32120 1414 32120 1414 4 vdd
port 66 nsew
rlabel metal3 s 25112 1414 25112 1414 4 vdd
port 66 nsew
rlabel metal3 s 20440 1414 20440 1414 4 vdd
port 66 nsew
rlabel metal3 s 22776 1414 22776 1414 4 vdd
port 66 nsew
rlabel metal3 s 29784 1414 29784 1414 4 vdd
port 66 nsew
rlabel metal3 s 33288 1414 33288 1414 4 vdd
port 66 nsew
rlabel metal3 s 36792 1414 36792 1414 4 vdd
port 66 nsew
rlabel metal3 s 23944 0 23944 0 4 gnd
port 67 nsew
rlabel metal3 s 5256 0 5256 0 4 gnd
port 67 nsew
rlabel metal3 s 27448 0 27448 0 4 gnd
port 67 nsew
rlabel metal3 s 30952 0 30952 0 4 gnd
port 67 nsew
rlabel metal3 s 34456 0 34456 0 4 gnd
port 67 nsew
rlabel metal3 s 36792 0 36792 0 4 gnd
port 67 nsew
rlabel metal3 s 26280 0 26280 0 4 gnd
port 67 nsew
rlabel metal3 s 19272 0 19272 0 4 gnd
port 67 nsew
rlabel metal3 s 13432 0 13432 0 4 gnd
port 67 nsew
rlabel metal3 s 1752 0 1752 0 4 gnd
port 67 nsew
rlabel metal3 s 18104 0 18104 0 4 gnd
port 67 nsew
rlabel metal3 s 6424 0 6424 0 4 gnd
port 67 nsew
rlabel metal3 s 25112 0 25112 0 4 gnd
port 67 nsew
rlabel metal3 s 11096 0 11096 0 4 gnd
port 67 nsew
rlabel metal3 s 9928 0 9928 0 4 gnd
port 67 nsew
rlabel metal3 s 584 0 584 0 4 gnd
port 67 nsew
rlabel metal3 s 8760 0 8760 0 4 gnd
port 67 nsew
rlabel metal3 s 21608 0 21608 0 4 gnd
port 67 nsew
rlabel metal3 s 15768 0 15768 0 4 gnd
port 67 nsew
rlabel metal3 s 16936 0 16936 0 4 gnd
port 67 nsew
rlabel metal3 s 14600 0 14600 0 4 gnd
port 67 nsew
rlabel metal3 s 33288 0 33288 0 4 gnd
port 67 nsew
rlabel metal3 s 7592 0 7592 0 4 gnd
port 67 nsew
rlabel metal3 s 29784 0 29784 0 4 gnd
port 67 nsew
rlabel metal3 s 35624 0 35624 0 4 gnd
port 67 nsew
rlabel metal3 s 20440 0 20440 0 4 gnd
port 67 nsew
rlabel metal3 s 12264 0 12264 0 4 gnd
port 67 nsew
rlabel metal3 s 32120 0 32120 0 4 gnd
port 67 nsew
rlabel metal3 s 22776 0 22776 0 4 gnd
port 67 nsew
rlabel metal3 s 28616 0 28616 0 4 gnd
port 67 nsew
rlabel metal3 s 4088 0 4088 0 4 gnd
port 67 nsew
rlabel metal3 s 2920 0 2920 0 4 gnd
port 67 nsew
rlabel metal3 s 18688 308 18688 308 4 clk
port 65 nsew
<< properties >>
string FIXED_BBOX 36759 -37 36825 0
string GDS_END 6489486
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 6454692
<< end >>
