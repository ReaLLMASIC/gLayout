magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect 8566 6529 13654 7090
rect 4468 5098 13654 6529
rect 4468 -484 13004 5098
<< nwell >>
rect 2447 11094 2545 11916
rect 8478 6843 13789 7185
rect 8478 6609 8821 6843
rect 182 4440 880 6322
rect 182 2032 880 3428
rect 4388 6198 8821 6609
rect 1601 267 3181 5231
rect 4388 -251 4748 6198
rect 13396 5372 13789 6843
rect 12797 4970 13789 5372
rect 12797 -251 13170 4970
rect 4388 -593 13170 -251
<< pwell >>
rect 9985 12052 12086 12146
rect 11992 11233 12086 12052
rect 6292 10367 6386 11191
rect 9990 11139 12086 11233
rect 11673 10367 11767 11139
rect 6292 10273 11767 10367
rect 6292 8808 6386 10273
rect 6292 8703 6435 8808
rect 10003 8725 10097 10273
rect 940 6193 1541 6281
rect 940 4338 1028 6193
rect 223 4250 1028 4338
rect 223 3576 311 4250
rect 751 3576 1028 4250
rect 223 3488 1028 3576
rect 940 1972 1028 3488
rect 223 1884 1028 1972
rect 223 396 311 1884
rect 751 396 1028 1884
rect 1453 396 1541 6193
rect 223 308 1541 396
rect 3242 5174 4226 5407
rect 3242 5088 4326 5174
rect 3242 3480 3756 5088
rect 3242 1967 3464 3480
rect 3670 1967 3756 3480
rect 3242 410 3756 1967
rect 4240 410 4326 5088
rect 3242 324 4326 410
rect 4808 5056 12736 5144
rect 4808 3770 4896 5056
rect 6786 4412 7072 4530
rect 6888 4404 7072 4412
rect 6888 4286 7238 4404
rect 9441 3770 9529 5056
rect 4808 3616 9529 3770
rect 4808 1631 4896 3616
rect 9441 1631 9529 3616
rect 4808 1477 9529 1631
rect 4808 271 4896 1477
rect 6888 935 7153 1053
rect 6888 927 7072 935
rect 6803 809 7072 927
rect 9441 516 9529 1477
rect 10270 516 10356 5056
rect 12648 516 12736 5056
rect 9441 428 12736 516
rect 9441 271 9793 428
rect 4808 183 9793 271
rect 9623 170 9793 183
rect 10031 170 10201 428
rect 9623 165 9743 170
rect 10081 165 10201 170
rect 10402 170 10572 428
rect 10402 165 10522 170
rect 10810 165 10980 428
rect 11161 170 11331 428
rect 11569 170 11739 428
rect 11161 165 11281 170
rect 11619 165 11739 170
rect 12128 170 12298 428
rect 12536 170 12706 428
rect 12128 165 12248 170
rect 10810 10 10927 165
rect 6490 -168 6660 10
rect 8273 -168 8443 10
rect 10757 -168 10927 10
rect 12540 10 12706 170
rect 12540 -168 12710 10
<< ndiff >>
rect 6516 -28 6634 -16
rect 6516 -130 6524 -28
rect 6626 -130 6634 -28
rect 6516 -142 6634 -130
rect 8299 -28 8417 -16
rect 8299 -130 8307 -28
rect 8409 -130 8417 -28
rect 8299 -142 8417 -130
rect 10783 -28 10901 -16
rect 10783 -130 10791 -28
rect 10893 -130 10901 -28
rect 10783 -142 10901 -130
rect 12566 -28 12684 -16
rect 12566 -130 12574 -28
rect 12676 -130 12684 -28
rect 12566 -142 12684 -130
<< mvndiff >>
rect 6812 4438 7046 4504
rect 6914 4312 7212 4378
rect 6914 961 7127 1027
rect 6829 835 7046 901
rect 9649 322 9717 327
rect 10107 322 10175 327
rect 9649 310 9767 322
rect 9649 208 9657 310
rect 9759 208 9767 310
rect 9649 196 9767 208
rect 10057 310 10175 322
rect 10057 208 10065 310
rect 10167 208 10175 310
rect 10057 196 10175 208
rect 9649 191 9717 196
rect 10107 191 10175 196
rect 10428 322 10496 327
rect 10886 322 10954 327
rect 10428 310 10546 322
rect 10428 208 10436 310
rect 10538 208 10546 310
rect 10428 196 10546 208
rect 10836 310 10954 322
rect 10836 208 10844 310
rect 10946 208 10954 310
rect 10836 196 10954 208
rect 10428 191 10496 196
rect 10886 191 10954 196
rect 11187 322 11255 327
rect 11645 322 11713 327
rect 11187 310 11305 322
rect 11187 208 11195 310
rect 11297 208 11305 310
rect 11187 196 11305 208
rect 11595 310 11713 322
rect 11595 208 11603 310
rect 11705 208 11713 310
rect 11595 196 11713 208
rect 11187 191 11255 196
rect 11645 191 11713 196
rect 12154 322 12222 327
rect 12612 322 12680 327
rect 12154 310 12272 322
rect 12154 208 12162 310
rect 12264 208 12272 310
rect 12154 196 12272 208
rect 12562 310 12680 322
rect 12562 208 12570 310
rect 12672 208 12680 310
rect 12562 196 12680 208
rect 12154 191 12222 196
rect 12612 191 12680 196
<< ndiffc >>
rect 9725 276 9759 310
rect 9725 208 9759 242
rect 10065 276 10099 310
rect 10065 208 10099 242
rect 10504 276 10538 310
rect 10504 208 10538 242
rect 10844 276 10878 310
rect 10844 208 10878 242
rect 11263 276 11297 310
rect 11263 208 11297 242
rect 11603 276 11637 310
rect 11603 208 11637 242
rect 12230 276 12264 310
rect 12230 208 12264 242
rect 12570 276 12604 310
rect 12570 208 12604 242
rect 6524 -130 6626 -28
rect 8307 -130 8409 -28
rect 10791 -130 10893 -28
rect 12574 -130 12676 -28
<< mvndiffc >>
rect 9657 276 9725 310
rect 9657 242 9759 276
rect 9657 208 9725 242
rect 10099 276 10167 310
rect 10065 242 10167 276
rect 10099 208 10167 242
rect 10436 276 10504 310
rect 10436 242 10538 276
rect 10436 208 10504 242
rect 10878 276 10946 310
rect 10844 242 10946 276
rect 10878 208 10946 242
rect 11195 276 11263 310
rect 11195 242 11297 276
rect 11195 208 11263 242
rect 11637 276 11705 310
rect 11603 242 11705 276
rect 11637 208 11705 242
rect 12162 276 12230 310
rect 12162 242 12264 276
rect 12162 208 12230 242
rect 12604 276 12672 310
rect 12570 242 12672 276
rect 12604 208 12672 242
<< psubdiff >>
rect 966 6254 1515 6255
rect 966 6220 1000 6254
rect 1034 6220 1068 6254
rect 1102 6220 1136 6254
rect 1170 6220 1204 6254
rect 1238 6220 1272 6254
rect 1306 6220 1340 6254
rect 1374 6220 1408 6254
rect 1442 6221 1515 6254
rect 1442 6220 1480 6221
rect 966 6219 1480 6220
rect 966 6136 1002 6219
rect 966 6102 967 6136
rect 1001 6102 1002 6136
rect 966 6068 1002 6102
rect 1479 6187 1480 6219
rect 1514 6187 1515 6221
rect 1479 6153 1515 6187
rect 1479 6119 1480 6153
rect 1514 6119 1515 6153
rect 966 6034 967 6068
rect 1001 6034 1002 6068
rect 966 6000 1002 6034
rect 966 5966 967 6000
rect 1001 5966 1002 6000
rect 966 5932 1002 5966
rect 966 5898 967 5932
rect 1001 5898 1002 5932
rect 966 5864 1002 5898
rect 966 5830 967 5864
rect 1001 5830 1002 5864
rect 966 5796 1002 5830
rect 1479 6085 1515 6119
rect 1479 6051 1480 6085
rect 1514 6051 1515 6085
rect 1479 6017 1515 6051
rect 1479 5983 1480 6017
rect 1514 5983 1515 6017
rect 1479 5949 1515 5983
rect 1479 5915 1480 5949
rect 1514 5915 1515 5949
rect 1479 5881 1515 5915
rect 1479 5847 1480 5881
rect 1514 5847 1515 5881
rect 1479 5813 1515 5847
rect 966 5762 967 5796
rect 1001 5762 1002 5796
rect 966 5728 1002 5762
rect 1479 5779 1480 5813
rect 1514 5779 1515 5813
rect 1479 5745 1515 5779
rect 966 5694 967 5728
rect 1001 5694 1002 5728
rect 966 5660 1002 5694
rect 966 5626 967 5660
rect 1001 5626 1002 5660
rect 966 5592 1002 5626
rect 1479 5711 1480 5745
rect 1514 5711 1515 5745
rect 1479 5677 1515 5711
rect 1479 5643 1480 5677
rect 1514 5643 1515 5677
rect 1479 5609 1515 5643
rect 966 5558 967 5592
rect 1001 5558 1002 5592
rect 966 5524 1002 5558
rect 966 5490 967 5524
rect 1001 5490 1002 5524
rect 966 5456 1002 5490
rect 966 5422 967 5456
rect 1001 5422 1002 5456
rect 1479 5575 1480 5609
rect 1514 5575 1515 5609
rect 1479 5541 1515 5575
rect 1479 5507 1480 5541
rect 1514 5507 1515 5541
rect 1479 5473 1515 5507
rect 966 5388 1002 5422
rect 966 5354 967 5388
rect 1001 5354 1002 5388
rect 966 5320 1002 5354
rect 966 5286 967 5320
rect 1001 5286 1002 5320
rect 966 5252 1002 5286
rect 1479 5439 1480 5473
rect 1514 5439 1515 5473
rect 1479 5405 1515 5439
rect 1479 5371 1480 5405
rect 1514 5371 1515 5405
rect 1479 5337 1515 5371
rect 1479 5303 1480 5337
rect 1514 5303 1515 5337
rect 1479 5269 1515 5303
rect 966 5218 967 5252
rect 1001 5218 1002 5252
rect 966 5184 1002 5218
rect 1479 5235 1480 5269
rect 1514 5235 1515 5269
rect 1479 5201 1515 5235
rect 966 5150 967 5184
rect 1001 5150 1002 5184
rect 966 5116 1002 5150
rect 966 5082 967 5116
rect 1001 5082 1002 5116
rect 966 5048 1002 5082
rect 966 5014 967 5048
rect 1001 5014 1002 5048
rect 966 4980 1002 5014
rect 1479 5167 1480 5201
rect 1514 5167 1515 5201
rect 1479 5133 1515 5167
rect 3268 5357 4200 5381
rect 3268 5355 4137 5357
rect 3268 5352 4069 5355
rect 3268 5318 3292 5352
rect 3326 5318 3362 5352
rect 3396 5318 3433 5352
rect 3467 5318 3504 5352
rect 3538 5318 3575 5352
rect 3609 5318 3646 5352
rect 3680 5318 3717 5352
rect 3751 5318 3788 5352
rect 3822 5318 3859 5352
rect 3893 5318 3930 5352
rect 3964 5318 4001 5352
rect 4035 5321 4069 5352
rect 4103 5323 4137 5355
rect 4171 5323 4200 5357
rect 4103 5321 4200 5323
rect 4035 5318 4200 5321
rect 3268 5289 4200 5318
rect 3268 5284 4137 5289
rect 3268 5250 3292 5284
rect 3326 5250 3362 5284
rect 3396 5250 3432 5284
rect 3466 5250 3502 5284
rect 3536 5250 3572 5284
rect 3606 5250 3643 5284
rect 3677 5250 3714 5284
rect 3748 5250 3785 5284
rect 3819 5250 3856 5284
rect 3890 5250 3927 5284
rect 3961 5250 3998 5284
rect 4032 5250 4069 5284
rect 4103 5255 4137 5284
rect 4171 5255 4200 5289
rect 4103 5250 4200 5255
rect 3268 5216 4200 5250
rect 3268 5182 3292 5216
rect 3326 5182 3362 5216
rect 3396 5182 3432 5216
rect 3466 5182 3502 5216
rect 3536 5182 3572 5216
rect 3606 5182 3642 5216
rect 3676 5182 3712 5216
rect 3746 5182 3782 5216
rect 3816 5182 3852 5216
rect 3886 5182 3922 5216
rect 3956 5182 3992 5216
rect 4026 5182 4062 5216
rect 4096 5182 4132 5216
rect 4166 5182 4200 5216
rect 1479 5099 1480 5133
rect 1514 5099 1515 5133
rect 1479 5065 1515 5099
rect 1479 5031 1480 5065
rect 1514 5031 1515 5065
rect 966 4946 967 4980
rect 1001 4946 1002 4980
rect 966 4912 1002 4946
rect 966 4878 967 4912
rect 1001 4878 1002 4912
rect 966 4844 1002 4878
rect 966 4810 967 4844
rect 1001 4810 1002 4844
rect 1479 4997 1515 5031
rect 1479 4963 1480 4997
rect 1514 4963 1515 4997
rect 1479 4929 1515 4963
rect 1479 4895 1480 4929
rect 1514 4895 1515 4929
rect 1479 4861 1515 4895
rect 966 4776 1002 4810
rect 966 4742 967 4776
rect 1001 4742 1002 4776
rect 966 4708 1002 4742
rect 966 4674 967 4708
rect 1001 4674 1002 4708
rect 966 4640 1002 4674
rect 966 4606 967 4640
rect 1001 4606 1002 4640
rect 966 4572 1002 4606
rect 966 4538 967 4572
rect 1001 4538 1002 4572
rect 966 4504 1002 4538
rect 966 4470 967 4504
rect 1001 4470 1002 4504
rect 966 4436 1002 4470
rect 966 4402 967 4436
rect 1001 4402 1002 4436
rect 966 4368 1002 4402
rect 966 4334 967 4368
rect 1001 4334 1002 4368
rect 249 4311 813 4312
rect 249 4277 283 4311
rect 317 4277 351 4311
rect 385 4277 419 4311
rect 453 4277 487 4311
rect 521 4277 555 4311
rect 589 4277 623 4311
rect 657 4277 691 4311
rect 725 4278 813 4311
rect 725 4277 778 4278
rect 249 4276 778 4277
rect 249 4242 285 4276
rect 249 4208 250 4242
rect 284 4208 285 4242
rect 249 4174 285 4208
rect 249 4140 250 4174
rect 284 4140 285 4174
rect 777 4244 778 4276
rect 812 4244 813 4278
rect 777 4210 813 4244
rect 777 4176 778 4210
rect 812 4176 813 4210
rect 249 4106 285 4140
rect 249 4072 250 4106
rect 284 4072 285 4106
rect 249 4038 285 4072
rect 249 4004 250 4038
rect 284 4004 285 4038
rect 249 3970 285 4004
rect 249 3936 250 3970
rect 284 3936 285 3970
rect 249 3902 285 3936
rect 249 3868 250 3902
rect 284 3868 285 3902
rect 249 3834 285 3868
rect 249 3800 250 3834
rect 284 3800 285 3834
rect 249 3766 285 3800
rect 249 3732 250 3766
rect 284 3732 285 3766
rect 249 3550 285 3732
rect 777 4142 813 4176
rect 777 4108 778 4142
rect 812 4108 813 4142
rect 777 4074 813 4108
rect 777 4040 778 4074
rect 812 4040 813 4074
rect 777 4006 813 4040
rect 777 3972 778 4006
rect 812 3972 813 4006
rect 777 3938 813 3972
rect 777 3904 778 3938
rect 812 3904 813 3938
rect 777 3870 813 3904
rect 777 3836 778 3870
rect 812 3836 813 3870
rect 777 3802 813 3836
rect 777 3768 778 3802
rect 812 3768 813 3802
rect 777 3734 813 3768
rect 777 3700 778 3734
rect 812 3700 813 3734
rect 777 3666 813 3700
rect 777 3632 778 3666
rect 812 3632 813 3666
rect 777 3550 813 3632
rect 249 3549 813 3550
rect 249 3515 337 3549
rect 371 3515 405 3549
rect 439 3515 473 3549
rect 507 3515 541 3549
rect 575 3515 609 3549
rect 643 3515 677 3549
rect 711 3515 745 3549
rect 779 3515 813 3549
rect 249 3514 813 3515
rect 966 4300 1002 4334
rect 966 4266 967 4300
rect 1001 4266 1002 4300
rect 966 4232 1002 4266
rect 966 4198 967 4232
rect 1001 4198 1002 4232
rect 966 4164 1002 4198
rect 966 4130 967 4164
rect 1001 4130 1002 4164
rect 966 4096 1002 4130
rect 966 4062 967 4096
rect 1001 4062 1002 4096
rect 966 4028 1002 4062
rect 966 3994 967 4028
rect 1001 3994 1002 4028
rect 966 3960 1002 3994
rect 966 3926 967 3960
rect 1001 3926 1002 3960
rect 1479 4827 1480 4861
rect 1514 4827 1515 4861
rect 1479 4793 1515 4827
rect 1479 4759 1480 4793
rect 1514 4759 1515 4793
rect 1479 4725 1515 4759
rect 1479 4691 1480 4725
rect 1514 4691 1515 4725
rect 1479 4657 1515 4691
rect 1479 4623 1480 4657
rect 1514 4623 1515 4657
rect 1479 4589 1515 4623
rect 1479 4555 1480 4589
rect 1514 4555 1515 4589
rect 1479 4521 1515 4555
rect 1479 4487 1480 4521
rect 1514 4487 1515 4521
rect 1479 4453 1515 4487
rect 1479 4419 1480 4453
rect 1514 4419 1515 4453
rect 1479 4385 1515 4419
rect 1479 4351 1480 4385
rect 1514 4351 1515 4385
rect 1479 4317 1515 4351
rect 1479 4283 1480 4317
rect 1514 4283 1515 4317
rect 1479 4249 1515 4283
rect 1479 4215 1480 4249
rect 1514 4215 1515 4249
rect 1479 4181 1515 4215
rect 1479 4147 1480 4181
rect 1514 4147 1515 4181
rect 1479 4113 1515 4147
rect 1479 4079 1480 4113
rect 1514 4079 1515 4113
rect 1479 4045 1515 4079
rect 1479 4011 1480 4045
rect 1514 4011 1515 4045
rect 1479 3977 1515 4011
rect 966 3892 1002 3926
rect 966 3858 967 3892
rect 1001 3858 1002 3892
rect 966 3824 1002 3858
rect 966 3790 967 3824
rect 1001 3790 1002 3824
rect 966 3756 1002 3790
rect 966 3722 967 3756
rect 1001 3722 1002 3756
rect 1479 3943 1480 3977
rect 1514 3943 1515 3977
rect 1479 3909 1515 3943
rect 1479 3875 1480 3909
rect 1514 3875 1515 3909
rect 1479 3841 1515 3875
rect 1479 3807 1480 3841
rect 1514 3807 1515 3841
rect 1479 3773 1515 3807
rect 966 3688 1002 3722
rect 966 3654 967 3688
rect 1001 3654 1002 3688
rect 966 3620 1002 3654
rect 966 3586 967 3620
rect 1001 3586 1002 3620
rect 966 3552 1002 3586
rect 966 3518 967 3552
rect 1001 3518 1002 3552
rect 966 3484 1002 3518
rect 966 3450 967 3484
rect 1001 3450 1002 3484
rect 1479 3739 1480 3773
rect 1514 3739 1515 3773
rect 1479 3705 1515 3739
rect 1479 3671 1480 3705
rect 1514 3671 1515 3705
rect 1479 3637 1515 3671
rect 1479 3603 1480 3637
rect 1514 3603 1515 3637
rect 1479 3569 1515 3603
rect 1479 3535 1480 3569
rect 1514 3535 1515 3569
rect 1479 3501 1515 3535
rect 1479 3467 1480 3501
rect 1514 3467 1515 3501
rect 966 3416 1002 3450
rect 966 3382 967 3416
rect 1001 3382 1002 3416
rect 966 3122 1002 3382
rect 1479 3433 1515 3467
rect 1479 3399 1480 3433
rect 1514 3399 1515 3433
rect 1479 3365 1515 3399
rect 1479 3331 1480 3365
rect 1514 3331 1515 3365
rect 1479 3297 1515 3331
rect 1479 3263 1480 3297
rect 1514 3263 1515 3297
rect 1479 3229 1515 3263
rect 1479 3195 1480 3229
rect 1514 3195 1515 3229
rect 966 3088 967 3122
rect 1001 3088 1002 3122
rect 966 3054 1002 3088
rect 966 3020 967 3054
rect 1001 3020 1002 3054
rect 966 2986 1002 3020
rect 966 2952 967 2986
rect 1001 2952 1002 2986
rect 966 2918 1002 2952
rect 1479 3161 1515 3195
rect 1479 3127 1480 3161
rect 1514 3127 1515 3161
rect 1479 3093 1515 3127
rect 1479 3059 1480 3093
rect 1514 3059 1515 3093
rect 1479 3025 1515 3059
rect 1479 2991 1480 3025
rect 1514 2991 1515 3025
rect 1479 2957 1515 2991
rect 966 2884 967 2918
rect 1001 2884 1002 2918
rect 966 2850 1002 2884
rect 966 2816 967 2850
rect 1001 2816 1002 2850
rect 966 2782 1002 2816
rect 966 2748 967 2782
rect 1001 2748 1002 2782
rect 1479 2923 1480 2957
rect 1514 2923 1515 2957
rect 1479 2889 1515 2923
rect 1479 2855 1480 2889
rect 1514 2855 1515 2889
rect 1479 2821 1515 2855
rect 1479 2787 1480 2821
rect 1514 2787 1515 2821
rect 966 2714 1002 2748
rect 966 2680 967 2714
rect 1001 2680 1002 2714
rect 966 2646 1002 2680
rect 966 2612 967 2646
rect 1001 2612 1002 2646
rect 966 2578 1002 2612
rect 966 2544 967 2578
rect 1001 2544 1002 2578
rect 966 2510 1002 2544
rect 1479 2753 1515 2787
rect 1479 2719 1480 2753
rect 1514 2719 1515 2753
rect 1479 2685 1515 2719
rect 1479 2651 1480 2685
rect 1514 2651 1515 2685
rect 1479 2617 1515 2651
rect 1479 2583 1480 2617
rect 1514 2583 1515 2617
rect 1479 2549 1515 2583
rect 966 2476 967 2510
rect 1001 2476 1002 2510
rect 1479 2515 1480 2549
rect 1514 2515 1515 2549
rect 966 2442 1002 2476
rect 966 2408 967 2442
rect 1001 2408 1002 2442
rect 966 2374 1002 2408
rect 966 2340 967 2374
rect 1001 2340 1002 2374
rect 966 2306 1002 2340
rect 966 2272 967 2306
rect 1001 2272 1002 2306
rect 966 2238 1002 2272
rect 1479 2481 1515 2515
rect 1479 2447 1480 2481
rect 1514 2447 1515 2481
rect 1479 2413 1515 2447
rect 1479 2379 1480 2413
rect 1514 2379 1515 2413
rect 1479 2345 1515 2379
rect 1479 2311 1480 2345
rect 1514 2311 1515 2345
rect 1479 2277 1515 2311
rect 966 2204 967 2238
rect 1001 2204 1002 2238
rect 1479 2243 1480 2277
rect 1514 2243 1515 2277
rect 1479 2209 1515 2243
rect 966 2170 1002 2204
rect 966 2136 967 2170
rect 1001 2136 1002 2170
rect 966 2102 1002 2136
rect 966 2068 967 2102
rect 1001 2068 1002 2102
rect 1479 2175 1480 2209
rect 1514 2175 1515 2209
rect 1479 2141 1515 2175
rect 1479 2107 1480 2141
rect 1514 2107 1515 2141
rect 1479 2073 1515 2107
rect 966 2034 1002 2068
rect 966 2000 967 2034
rect 1001 2000 1002 2034
rect 966 1966 1002 2000
rect 249 1945 813 1946
rect 249 1911 283 1945
rect 317 1911 351 1945
rect 385 1911 419 1945
rect 453 1911 487 1945
rect 521 1911 555 1945
rect 589 1911 623 1945
rect 657 1911 691 1945
rect 725 1912 813 1945
rect 725 1911 778 1912
rect 249 1910 778 1911
rect 249 1830 285 1910
rect 249 1796 250 1830
rect 284 1796 285 1830
rect 249 1762 285 1796
rect 777 1878 778 1910
rect 812 1878 813 1912
rect 777 1844 813 1878
rect 777 1810 778 1844
rect 812 1810 813 1844
rect 249 1728 250 1762
rect 284 1728 285 1762
rect 249 1694 285 1728
rect 249 1660 250 1694
rect 284 1660 285 1694
rect 249 1626 285 1660
rect 249 1592 250 1626
rect 284 1592 285 1626
rect 249 1558 285 1592
rect 249 1524 250 1558
rect 284 1524 285 1558
rect 249 1490 285 1524
rect 249 1456 250 1490
rect 284 1456 285 1490
rect 249 1422 285 1456
rect 249 1388 250 1422
rect 284 1388 285 1422
rect 249 1354 285 1388
rect 249 1320 250 1354
rect 284 1320 285 1354
rect 249 1286 285 1320
rect 777 1776 813 1810
rect 777 1742 778 1776
rect 812 1742 813 1776
rect 777 1708 813 1742
rect 777 1674 778 1708
rect 812 1674 813 1708
rect 777 1640 813 1674
rect 777 1606 778 1640
rect 812 1606 813 1640
rect 777 1572 813 1606
rect 777 1538 778 1572
rect 812 1538 813 1572
rect 777 1504 813 1538
rect 777 1470 778 1504
rect 812 1470 813 1504
rect 777 1436 813 1470
rect 777 1402 778 1436
rect 812 1402 813 1436
rect 777 1368 813 1402
rect 777 1334 778 1368
rect 812 1334 813 1368
rect 249 1252 250 1286
rect 284 1252 285 1286
rect 249 1218 285 1252
rect 249 1184 250 1218
rect 284 1184 285 1218
rect 249 1150 285 1184
rect 249 1116 250 1150
rect 284 1116 285 1150
rect 777 1300 813 1334
rect 777 1266 778 1300
rect 812 1266 813 1300
rect 777 1232 813 1266
rect 777 1198 778 1232
rect 812 1198 813 1232
rect 777 1164 813 1198
rect 249 1082 285 1116
rect 249 1048 250 1082
rect 284 1048 285 1082
rect 249 1014 285 1048
rect 249 980 250 1014
rect 284 980 285 1014
rect 249 946 285 980
rect 249 912 250 946
rect 284 912 285 946
rect 249 878 285 912
rect 249 844 250 878
rect 284 844 285 878
rect 249 810 285 844
rect 249 776 250 810
rect 284 776 285 810
rect 249 742 285 776
rect 249 708 250 742
rect 284 708 285 742
rect 249 674 285 708
rect 249 640 250 674
rect 284 640 285 674
rect 249 606 285 640
rect 249 572 250 606
rect 284 572 285 606
rect 249 538 285 572
rect 249 504 250 538
rect 284 504 285 538
rect 249 470 285 504
rect 777 1130 778 1164
rect 812 1130 813 1164
rect 777 1096 813 1130
rect 777 1062 778 1096
rect 812 1062 813 1096
rect 777 1028 813 1062
rect 777 994 778 1028
rect 812 994 813 1028
rect 777 960 813 994
rect 777 926 778 960
rect 812 926 813 960
rect 777 892 813 926
rect 777 858 778 892
rect 812 858 813 892
rect 777 824 813 858
rect 777 790 778 824
rect 812 790 813 824
rect 777 756 813 790
rect 777 722 778 756
rect 812 722 813 756
rect 777 688 813 722
rect 777 654 778 688
rect 812 654 813 688
rect 777 620 813 654
rect 777 586 778 620
rect 812 586 813 620
rect 777 552 813 586
rect 777 518 778 552
rect 812 518 813 552
rect 249 436 250 470
rect 284 436 285 470
rect 249 402 285 436
rect 249 368 250 402
rect 284 370 285 402
rect 777 484 813 518
rect 777 450 778 484
rect 812 450 813 484
rect 777 370 813 450
rect 284 369 813 370
rect 284 368 337 369
rect 249 335 337 368
rect 371 335 405 369
rect 439 335 473 369
rect 507 335 541 369
rect 575 335 609 369
rect 643 335 677 369
rect 711 335 745 369
rect 779 335 813 369
rect 249 334 813 335
rect 966 1932 967 1966
rect 1001 1932 1002 1966
rect 966 1898 1002 1932
rect 966 1864 967 1898
rect 1001 1864 1002 1898
rect 966 1830 1002 1864
rect 1479 2039 1480 2073
rect 1514 2039 1515 2073
rect 1479 2005 1515 2039
rect 1479 1971 1480 2005
rect 1514 1971 1515 2005
rect 1479 1937 1515 1971
rect 1479 1903 1480 1937
rect 1514 1903 1515 1937
rect 1479 1869 1515 1903
rect 966 1796 967 1830
rect 1001 1796 1002 1830
rect 966 1762 1002 1796
rect 966 1728 967 1762
rect 1001 1728 1002 1762
rect 966 1694 1002 1728
rect 966 1660 967 1694
rect 1001 1660 1002 1694
rect 966 1626 1002 1660
rect 966 1592 967 1626
rect 1001 1592 1002 1626
rect 966 1558 1002 1592
rect 1479 1835 1480 1869
rect 1514 1835 1515 1869
rect 1479 1801 1515 1835
rect 1479 1767 1480 1801
rect 1514 1767 1515 1801
rect 1479 1733 1515 1767
rect 1479 1699 1480 1733
rect 1514 1699 1515 1733
rect 1479 1665 1515 1699
rect 1479 1631 1480 1665
rect 1514 1631 1515 1665
rect 1479 1597 1515 1631
rect 966 1524 967 1558
rect 1001 1524 1002 1558
rect 966 1490 1002 1524
rect 966 1456 967 1490
rect 1001 1456 1002 1490
rect 966 1422 1002 1456
rect 966 1388 967 1422
rect 1001 1388 1002 1422
rect 966 1354 1002 1388
rect 1479 1563 1480 1597
rect 1514 1563 1515 1597
rect 1479 1529 1515 1563
rect 1479 1495 1480 1529
rect 1514 1495 1515 1529
rect 1479 1461 1515 1495
rect 1479 1427 1480 1461
rect 1514 1427 1515 1461
rect 1479 1393 1515 1427
rect 966 1320 967 1354
rect 1001 1320 1002 1354
rect 966 1286 1002 1320
rect 966 1252 967 1286
rect 1001 1252 1002 1286
rect 966 1218 1002 1252
rect 966 1184 967 1218
rect 1001 1184 1002 1218
rect 966 1150 1002 1184
rect 966 1116 967 1150
rect 1001 1116 1002 1150
rect 966 1082 1002 1116
rect 966 1048 967 1082
rect 1001 1048 1002 1082
rect 966 1014 1002 1048
rect 966 980 967 1014
rect 1001 980 1002 1014
rect 966 946 1002 980
rect 966 912 967 946
rect 1001 912 1002 946
rect 966 878 1002 912
rect 966 844 967 878
rect 1001 844 1002 878
rect 966 810 1002 844
rect 966 776 967 810
rect 1001 776 1002 810
rect 966 742 1002 776
rect 966 708 967 742
rect 1001 708 1002 742
rect 966 674 1002 708
rect 966 640 967 674
rect 1001 640 1002 674
rect 966 606 1002 640
rect 966 572 967 606
rect 1001 572 1002 606
rect 966 538 1002 572
rect 966 504 967 538
rect 1001 504 1002 538
rect 966 470 1002 504
rect 1479 1359 1480 1393
rect 1514 1359 1515 1393
rect 1479 1325 1515 1359
rect 1479 1291 1480 1325
rect 1514 1291 1515 1325
rect 1479 1257 1515 1291
rect 1479 1223 1480 1257
rect 1514 1223 1515 1257
rect 1479 1189 1515 1223
rect 1479 1155 1480 1189
rect 1514 1155 1515 1189
rect 1479 1121 1515 1155
rect 1479 1087 1480 1121
rect 1514 1087 1515 1121
rect 1479 1053 1515 1087
rect 1479 1019 1480 1053
rect 1514 1019 1515 1053
rect 1479 985 1515 1019
rect 1479 951 1480 985
rect 1514 951 1515 985
rect 1479 917 1515 951
rect 1479 883 1480 917
rect 1514 883 1515 917
rect 1479 849 1515 883
rect 1479 815 1480 849
rect 1514 815 1515 849
rect 1479 781 1515 815
rect 1479 747 1480 781
rect 1514 747 1515 781
rect 1479 713 1515 747
rect 1479 679 1480 713
rect 1514 679 1515 713
rect 1479 645 1515 679
rect 1479 611 1480 645
rect 1514 611 1515 645
rect 1479 577 1515 611
rect 1479 543 1480 577
rect 1514 543 1515 577
rect 1479 509 1515 543
rect 966 436 967 470
rect 1001 436 1002 470
rect 966 402 1002 436
rect 966 368 967 402
rect 1001 370 1002 402
rect 1479 475 1480 509
rect 1514 475 1515 509
rect 1479 370 1515 475
rect 1001 369 1515 370
rect 1001 368 1039 369
rect 966 335 1039 368
rect 1073 335 1107 369
rect 1141 335 1175 369
rect 1209 335 1243 369
rect 1277 335 1311 369
rect 1345 335 1379 369
rect 1413 335 1447 369
rect 1481 335 1515 369
rect 966 334 1515 335
rect 3268 5148 4200 5182
rect 3268 5130 3730 5148
rect 3268 5129 3490 5130
rect 3302 5095 3336 5129
rect 3370 5095 3404 5129
rect 3438 5096 3490 5129
rect 3524 5096 3558 5130
rect 3592 5096 3626 5130
rect 3660 5096 3730 5130
rect 3764 5114 3798 5148
rect 3832 5114 3866 5148
rect 3900 5114 3934 5148
rect 3968 5114 4002 5148
rect 4036 5114 4070 5148
rect 4104 5114 4138 5148
rect 4172 5114 4206 5148
rect 4240 5114 4300 5148
rect 3438 5095 3730 5096
rect 3268 5061 3730 5095
rect 3268 5060 3490 5061
rect 3302 5026 3336 5060
rect 3370 5026 3404 5060
rect 3438 5027 3490 5060
rect 3524 5027 3558 5061
rect 3592 5027 3626 5061
rect 3660 5042 3730 5061
rect 3660 5027 3696 5042
rect 3438 5026 3696 5027
rect 3268 5008 3696 5026
rect 3268 4992 3730 5008
rect 3268 4991 3490 4992
rect 3302 4957 3336 4991
rect 3370 4957 3404 4991
rect 3438 4957 3490 4991
rect 3268 4922 3490 4957
rect 3302 4888 3336 4922
rect 3370 4888 3404 4922
rect 3438 4888 3490 4922
rect 3268 4853 3490 4888
rect 3302 4819 3336 4853
rect 3370 4819 3404 4853
rect 3438 4819 3490 4853
rect 3268 4784 3490 4819
rect 3302 4750 3336 4784
rect 3370 4750 3404 4784
rect 3438 4750 3490 4784
rect 3268 4715 3490 4750
rect 3302 4681 3336 4715
rect 3370 4681 3404 4715
rect 3438 4681 3490 4715
rect 3268 4646 3490 4681
rect 3302 4612 3336 4646
rect 3370 4612 3404 4646
rect 3438 4612 3490 4646
rect 3268 4577 3490 4612
rect 3302 4543 3336 4577
rect 3370 4543 3404 4577
rect 3438 4543 3490 4577
rect 3268 4508 3490 4543
rect 3302 4474 3336 4508
rect 3370 4474 3404 4508
rect 3438 4474 3490 4508
rect 3268 4439 3490 4474
rect 3302 4405 3336 4439
rect 3370 4405 3404 4439
rect 3438 4405 3490 4439
rect 3268 4370 3490 4405
rect 3302 4336 3336 4370
rect 3370 4336 3404 4370
rect 3438 4336 3490 4370
rect 3268 4301 3490 4336
rect 3302 4267 3336 4301
rect 3370 4267 3404 4301
rect 3438 4267 3490 4301
rect 3268 4232 3490 4267
rect 3302 4198 3336 4232
rect 3370 4198 3404 4232
rect 3438 4198 3490 4232
rect 3268 4163 3490 4198
rect 3302 4129 3336 4163
rect 3370 4129 3404 4163
rect 3438 4129 3490 4163
rect 3268 4094 3490 4129
rect 3302 4060 3336 4094
rect 3370 4060 3404 4094
rect 3438 4060 3490 4094
rect 3268 4025 3490 4060
rect 3302 3991 3336 4025
rect 3370 3991 3404 4025
rect 3438 3991 3490 4025
rect 3268 3956 3490 3991
rect 3302 3922 3336 3956
rect 3370 3922 3404 3956
rect 3438 3922 3490 3956
rect 3268 3887 3490 3922
rect 3302 3853 3336 3887
rect 3370 3853 3404 3887
rect 3438 3853 3490 3887
rect 3268 3818 3490 3853
rect 3302 3784 3336 3818
rect 3370 3784 3404 3818
rect 3438 3784 3490 3818
rect 3268 3749 3490 3784
rect 3302 3715 3336 3749
rect 3370 3715 3404 3749
rect 3438 3715 3490 3749
rect 3268 3680 3490 3715
rect 3302 3646 3336 3680
rect 3370 3646 3404 3680
rect 3438 3646 3490 3680
rect 3268 3611 3490 3646
rect 3302 3577 3336 3611
rect 3370 3577 3404 3611
rect 3438 3577 3490 3611
rect 3268 3542 3490 3577
rect 3302 3508 3336 3542
rect 3370 3508 3404 3542
rect 3438 3530 3490 3542
rect 3660 4974 3730 4992
rect 3660 4940 3696 4974
rect 4266 5048 4300 5114
rect 4266 4980 4300 5014
rect 3660 4906 3730 4940
rect 3660 4872 3696 4906
rect 3660 4838 3730 4872
rect 3660 4804 3696 4838
rect 3660 4770 3730 4804
rect 4266 4912 4300 4946
rect 4266 4844 4300 4878
rect 3660 4736 3696 4770
rect 3660 4702 3730 4736
rect 3660 4668 3696 4702
rect 3660 4634 3730 4668
rect 3660 4600 3696 4634
rect 3660 4566 3730 4600
rect 3660 4532 3696 4566
rect 3660 4498 3730 4532
rect 3660 4464 3696 4498
rect 4266 4776 4300 4810
rect 4266 4708 4300 4742
rect 4266 4640 4300 4674
rect 4266 4572 4300 4606
rect 4266 4504 4300 4538
rect 3660 4430 3730 4464
rect 3660 4396 3696 4430
rect 3660 4362 3730 4396
rect 3660 4328 3696 4362
rect 3660 4294 3730 4328
rect 3660 4260 3696 4294
rect 3660 4226 3730 4260
rect 3660 4192 3696 4226
rect 3660 4158 3730 4192
rect 3660 4124 3696 4158
rect 3660 4090 3730 4124
rect 3660 4056 3696 4090
rect 3660 4022 3730 4056
rect 3660 3988 3696 4022
rect 3660 3954 3730 3988
rect 3660 3920 3696 3954
rect 3660 3886 3730 3920
rect 3660 3852 3696 3886
rect 3660 3818 3730 3852
rect 3660 3784 3696 3818
rect 3660 3750 3730 3784
rect 3660 3716 3696 3750
rect 3660 3682 3730 3716
rect 3660 3648 3696 3682
rect 3660 3614 3730 3648
rect 3660 3580 3696 3614
rect 4266 4436 4300 4470
rect 4266 4368 4300 4402
rect 4266 4300 4300 4334
rect 4266 4232 4300 4266
rect 4266 4164 4300 4198
rect 4266 4096 4300 4130
rect 4266 4028 4300 4062
rect 4266 3960 4300 3994
rect 4266 3892 4300 3926
rect 4266 3824 4300 3858
rect 4266 3756 4300 3790
rect 4266 3688 4300 3722
rect 4266 3620 4300 3654
rect 3660 3546 3730 3580
rect 3660 3530 3696 3546
rect 3438 3512 3696 3530
rect 3438 3508 3730 3512
rect 3268 3506 3730 3508
rect 3268 3473 3438 3506
rect 3302 3439 3336 3473
rect 3370 3439 3404 3473
rect 3268 3404 3438 3439
rect 3696 3478 3730 3506
rect 3696 3410 3730 3444
rect 3302 3370 3336 3404
rect 3370 3370 3404 3404
rect 3268 3335 3438 3370
rect 3302 3301 3336 3335
rect 3370 3301 3404 3335
rect 3268 3266 3438 3301
rect 3696 3342 3730 3376
rect 3302 3232 3336 3266
rect 3370 3232 3404 3266
rect 3268 3197 3438 3232
rect 3302 3163 3336 3197
rect 3370 3163 3404 3197
rect 3268 3128 3438 3163
rect 3696 3274 3730 3308
rect 3696 3206 3730 3240
rect 3696 3138 3730 3172
rect 3696 3070 3730 3104
rect 4266 3552 4300 3586
rect 4266 3484 4300 3518
rect 4266 3416 4300 3450
rect 4266 3348 4300 3382
rect 4266 3280 4300 3314
rect 4266 3212 4300 3246
rect 4266 3144 4300 3178
rect 3696 3002 3730 3036
rect 3696 2934 3730 2968
rect 3696 2866 3730 2900
rect 3696 2798 3730 2832
rect 3696 2730 3730 2764
rect 3696 2662 3730 2696
rect 3696 2594 3730 2628
rect 3696 2526 3730 2560
rect 3696 2458 3730 2492
rect 3696 2390 3730 2424
rect 4266 3076 4300 3110
rect 4266 3008 4300 3042
rect 4266 2940 4300 2974
rect 4266 2872 4300 2906
rect 4266 2804 4300 2838
rect 4266 2736 4300 2770
rect 4266 2668 4300 2702
rect 4266 2600 4300 2634
rect 4266 2532 4300 2566
rect 4266 2464 4300 2498
rect 3696 2322 3730 2356
rect 3696 2254 3730 2288
rect 3696 2186 3730 2220
rect 3696 2118 3730 2152
rect 4266 2396 4300 2430
rect 4266 2328 4300 2362
rect 4266 2260 4300 2294
rect 4266 2192 4300 2226
rect 3696 2050 3730 2084
rect 3696 1982 3730 2016
rect 4266 2124 4300 2158
rect 4266 2056 4300 2090
rect 4266 1988 4300 2022
rect 3696 1941 3730 1948
rect 3438 1917 3730 1941
rect 3438 1883 3490 1917
rect 3524 1883 3558 1917
rect 3592 1883 3626 1917
rect 3660 1914 3730 1917
rect 3660 1883 3696 1914
rect 3438 1880 3696 1883
rect 3438 1848 3730 1880
rect 3438 1814 3490 1848
rect 3524 1814 3558 1848
rect 3592 1814 3626 1848
rect 3660 1846 3730 1848
rect 3660 1814 3696 1846
rect 3438 1812 3696 1814
rect 3438 1779 3730 1812
rect 3438 1745 3490 1779
rect 3524 1745 3558 1779
rect 3592 1745 3626 1779
rect 3660 1778 3730 1779
rect 3660 1745 3696 1778
rect 3438 1744 3696 1745
rect 3438 1710 3730 1744
rect 3438 1676 3490 1710
rect 3524 1676 3558 1710
rect 3592 1676 3626 1710
rect 3660 1676 3696 1710
rect 3438 1642 3730 1676
rect 3438 1641 3696 1642
rect 3438 1607 3490 1641
rect 3524 1607 3558 1641
rect 3592 1607 3626 1641
rect 3660 1608 3696 1641
rect 3660 1607 3730 1608
rect 3438 1574 3730 1607
rect 3438 1572 3696 1574
rect 3438 1538 3490 1572
rect 3524 1538 3558 1572
rect 3592 1538 3626 1572
rect 3660 1540 3696 1572
rect 3660 1538 3730 1540
rect 3438 1506 3730 1538
rect 3438 1503 3696 1506
rect 3438 1469 3490 1503
rect 3524 1469 3558 1503
rect 3592 1469 3626 1503
rect 3660 1472 3696 1503
rect 3660 1469 3730 1472
rect 3438 1438 3730 1469
rect 3438 1434 3696 1438
rect 3438 1400 3490 1434
rect 3524 1400 3558 1434
rect 3592 1400 3626 1434
rect 3660 1404 3696 1434
rect 4266 1920 4300 1954
rect 4266 1852 4300 1886
rect 4266 1784 4300 1818
rect 4266 1716 4300 1750
rect 4266 1648 4300 1682
rect 4266 1580 4300 1614
rect 4266 1512 4300 1546
rect 4266 1444 4300 1478
rect 3660 1400 3730 1404
rect 3438 1370 3730 1400
rect 3438 1365 3696 1370
rect 3438 1331 3490 1365
rect 3524 1331 3558 1365
rect 3592 1331 3626 1365
rect 3660 1336 3696 1365
rect 3660 1331 3730 1336
rect 3438 1302 3730 1331
rect 3438 1296 3696 1302
rect 3438 1262 3490 1296
rect 3524 1262 3558 1296
rect 3592 1262 3626 1296
rect 3660 1268 3696 1296
rect 3660 1262 3730 1268
rect 3438 1234 3730 1262
rect 3438 1227 3696 1234
rect 3438 1193 3490 1227
rect 3524 1193 3558 1227
rect 3592 1193 3626 1227
rect 3660 1200 3696 1227
rect 3660 1193 3730 1200
rect 3438 1166 3730 1193
rect 3438 1158 3696 1166
rect 3438 1124 3490 1158
rect 3524 1124 3558 1158
rect 3592 1124 3626 1158
rect 3660 1132 3696 1158
rect 3660 1124 3730 1132
rect 3438 1098 3730 1124
rect 3438 1089 3696 1098
rect 3438 1055 3490 1089
rect 3524 1055 3558 1089
rect 3592 1055 3626 1089
rect 3660 1064 3696 1089
rect 3660 1055 3730 1064
rect 3438 1030 3730 1055
rect 3438 1020 3696 1030
rect 3438 374 3490 1020
rect 3660 996 3696 1020
rect 3660 962 3730 996
rect 3660 928 3696 962
rect 3660 894 3730 928
rect 3660 860 3696 894
rect 3660 826 3730 860
rect 3660 792 3696 826
rect 3660 758 3730 792
rect 3660 724 3696 758
rect 3660 690 3730 724
rect 3660 656 3696 690
rect 3660 622 3730 656
rect 3660 588 3696 622
rect 3660 554 3730 588
rect 3660 520 3696 554
rect 4266 1376 4300 1410
rect 4266 1308 4300 1342
rect 4266 1240 4300 1274
rect 4266 1172 4300 1206
rect 4266 1104 4300 1138
rect 4266 1036 4300 1070
rect 4266 968 4300 1002
rect 4266 900 4300 934
rect 4266 832 4300 866
rect 4266 764 4300 798
rect 4266 696 4300 730
rect 4266 628 4300 662
rect 4266 560 4300 594
rect 3660 486 3730 520
rect 3660 452 3696 486
rect 3660 418 3730 452
rect 3660 384 3696 418
rect 4266 492 4300 526
rect 3660 374 3824 384
rect 3268 350 3824 374
rect 3858 350 3892 384
rect 3926 350 3960 384
rect 3994 350 4028 384
rect 4062 350 4096 384
rect 4130 350 4164 384
rect 4198 350 4232 384
rect 4266 350 4300 458
<< nsubdiff >>
rect 249 3360 813 3361
rect 249 3326 283 3360
rect 317 3326 351 3360
rect 385 3326 419 3360
rect 453 3326 555 3360
rect 589 3326 623 3360
rect 657 3326 691 3360
rect 725 3327 813 3360
rect 725 3326 778 3327
rect 249 3325 778 3326
rect 249 3290 285 3325
rect 249 3256 250 3290
rect 284 3256 285 3290
rect 249 3222 285 3256
rect 249 3188 250 3222
rect 284 3188 285 3222
rect 777 3293 778 3325
rect 812 3293 813 3327
rect 777 3259 813 3293
rect 777 3225 778 3259
rect 812 3225 813 3259
rect 249 3154 285 3188
rect 249 3120 250 3154
rect 284 3120 285 3154
rect 249 3086 285 3120
rect 249 3052 250 3086
rect 284 3052 285 3086
rect 777 3191 813 3225
rect 777 3157 778 3191
rect 812 3157 813 3191
rect 777 3123 813 3157
rect 249 2779 285 3052
rect 777 3089 778 3123
rect 812 3089 813 3123
rect 777 3055 813 3089
rect 777 3021 778 3055
rect 812 3021 813 3055
rect 777 2987 813 3021
rect 777 2953 778 2987
rect 812 2953 813 2987
rect 777 2919 813 2953
rect 249 2745 250 2779
rect 284 2745 285 2779
rect 249 2711 285 2745
rect 249 2677 250 2711
rect 284 2677 285 2711
rect 777 2885 778 2919
rect 812 2885 813 2919
rect 777 2851 813 2885
rect 777 2817 778 2851
rect 812 2817 813 2851
rect 777 2783 813 2817
rect 777 2749 778 2783
rect 812 2749 813 2783
rect 777 2715 813 2749
rect 249 2643 285 2677
rect 249 2609 250 2643
rect 284 2609 285 2643
rect 249 2575 285 2609
rect 249 2541 250 2575
rect 284 2541 285 2575
rect 777 2681 778 2715
rect 812 2681 813 2715
rect 777 2647 813 2681
rect 777 2613 778 2647
rect 812 2613 813 2647
rect 777 2579 813 2613
rect 249 2507 285 2541
rect 249 2473 250 2507
rect 284 2473 285 2507
rect 249 2439 285 2473
rect 249 2405 250 2439
rect 284 2405 285 2439
rect 777 2545 778 2579
rect 812 2545 813 2579
rect 777 2511 813 2545
rect 777 2477 778 2511
rect 812 2477 813 2511
rect 777 2443 813 2477
rect 249 2371 285 2405
rect 249 2337 250 2371
rect 284 2337 285 2371
rect 777 2409 778 2443
rect 812 2409 813 2443
rect 777 2375 813 2409
rect 249 2303 285 2337
rect 249 2269 250 2303
rect 284 2269 285 2303
rect 249 2235 285 2269
rect 249 2201 250 2235
rect 284 2201 285 2235
rect 777 2341 778 2375
rect 812 2341 813 2375
rect 777 2307 813 2341
rect 777 2273 778 2307
rect 812 2273 813 2307
rect 249 2167 285 2201
rect 249 2133 250 2167
rect 284 2135 285 2167
rect 777 2135 813 2273
rect 284 2134 813 2135
rect 284 2133 337 2134
rect 249 2100 337 2133
rect 371 2100 405 2134
rect 439 2100 473 2134
rect 507 2100 541 2134
rect 575 2100 609 2134
rect 643 2100 677 2134
rect 711 2100 745 2134
rect 779 2100 813 2134
rect 249 2099 813 2100
<< mvpsubdiff >>
rect 10011 12116 12060 12120
rect 10011 12082 10070 12116
rect 10104 12082 10155 12116
rect 10189 12082 10240 12116
rect 10274 12082 10325 12116
rect 10359 12082 10410 12116
rect 10444 12082 10495 12116
rect 10529 12082 10580 12116
rect 10614 12082 10665 12116
rect 10699 12082 10750 12116
rect 10784 12082 10835 12116
rect 10869 12082 10920 12116
rect 10954 12082 11005 12116
rect 11039 12082 11090 12116
rect 11124 12082 11175 12116
rect 11209 12082 11260 12116
rect 11294 12082 11345 12116
rect 11379 12082 11430 12116
rect 11464 12082 11515 12116
rect 11549 12082 11600 12116
rect 11634 12082 11685 12116
rect 11719 12082 11770 12116
rect 11804 12082 11856 12116
rect 11890 12082 11942 12116
rect 11976 12082 12060 12116
rect 10011 12078 12060 12082
rect 12018 12027 12060 12078
rect 12018 11993 12022 12027
rect 12056 11993 12060 12027
rect 12018 11934 12060 11993
rect 12018 11900 12022 11934
rect 12056 11900 12060 11934
rect 12018 11841 12060 11900
rect 12018 11807 12022 11841
rect 12056 11807 12060 11841
rect 12018 11748 12060 11807
rect 12018 11714 12022 11748
rect 12056 11714 12060 11748
rect 12018 11655 12060 11714
rect 12018 11621 12022 11655
rect 12056 11621 12060 11655
rect 12018 11562 12060 11621
rect 12018 11528 12022 11562
rect 12056 11528 12060 11562
rect 12018 11469 12060 11528
rect 12018 11435 12022 11469
rect 12056 11435 12060 11469
rect 12018 11376 12060 11435
rect 12018 11342 12022 11376
rect 12056 11342 12060 11376
rect 12018 11283 12060 11342
rect 12018 11249 12022 11283
rect 12056 11249 12060 11283
rect 12018 11207 12060 11249
rect 10016 11203 12060 11207
rect 10016 11169 10066 11203
rect 10100 11169 10152 11203
rect 10186 11169 10238 11203
rect 10272 11169 10324 11203
rect 10358 11169 10410 11203
rect 10444 11169 10496 11203
rect 10530 11169 10582 11203
rect 10616 11169 10668 11203
rect 10702 11169 10754 11203
rect 10788 11169 10840 11203
rect 10874 11169 10927 11203
rect 10961 11169 11014 11203
rect 11048 11169 11101 11203
rect 11135 11169 11188 11203
rect 11222 11169 11275 11203
rect 11309 11169 11362 11203
rect 11396 11169 11449 11203
rect 11483 11169 11536 11203
rect 11570 11169 11623 11203
rect 11657 11169 11765 11203
rect 11799 11169 11852 11203
rect 11886 11169 11939 11203
rect 11973 11169 12060 11203
rect 10016 11165 12060 11169
rect 6318 11108 6360 11165
rect 6318 11074 6322 11108
rect 6356 11074 6360 11108
rect 6318 11023 6360 11074
rect 6318 10989 6322 11023
rect 6356 10989 6360 11023
rect 6318 10937 6360 10989
rect 6318 10903 6322 10937
rect 6356 10903 6360 10937
rect 6318 10851 6360 10903
rect 6318 10817 6322 10851
rect 6356 10817 6360 10851
rect 6318 10765 6360 10817
rect 6318 10731 6322 10765
rect 6356 10731 6360 10765
rect 6318 10679 6360 10731
rect 6318 10645 6322 10679
rect 6356 10645 6360 10679
rect 6318 10593 6360 10645
rect 6318 10559 6322 10593
rect 6356 10559 6360 10593
rect 6318 10507 6360 10559
rect 6318 10473 6322 10507
rect 6356 10473 6360 10507
rect 6318 10421 6360 10473
rect 11699 11120 11741 11165
rect 11699 11086 11703 11120
rect 11737 11086 11741 11120
rect 11699 11033 11741 11086
rect 11699 10999 11703 11033
rect 11737 10999 11741 11033
rect 11699 10945 11741 10999
rect 11699 10911 11703 10945
rect 11737 10911 11741 10945
rect 11699 10857 11741 10911
rect 11699 10823 11703 10857
rect 11737 10823 11741 10857
rect 11699 10769 11741 10823
rect 11699 10735 11703 10769
rect 11737 10735 11741 10769
rect 11699 10681 11741 10735
rect 11699 10647 11703 10681
rect 11737 10647 11741 10681
rect 11699 10593 11741 10647
rect 11699 10559 11703 10593
rect 11737 10559 11741 10593
rect 11699 10505 11741 10559
rect 11699 10471 11703 10505
rect 11737 10471 11741 10505
rect 6318 10387 6322 10421
rect 6356 10387 6360 10421
rect 11699 10417 11741 10471
rect 6318 10341 6360 10387
rect 11699 10383 11703 10417
rect 11737 10383 11741 10417
rect 11699 10341 11741 10383
rect 6318 10337 11741 10341
rect 6318 10335 6417 10337
rect 6318 10301 6322 10335
rect 6356 10303 6417 10335
rect 6451 10303 6503 10337
rect 6537 10303 6589 10337
rect 6623 10303 6675 10337
rect 6709 10303 6761 10337
rect 6795 10303 6847 10337
rect 6881 10303 6933 10337
rect 6967 10303 7019 10337
rect 7053 10303 7105 10337
rect 7139 10303 7191 10337
rect 7225 10303 7277 10337
rect 7311 10303 7363 10337
rect 7397 10303 7449 10337
rect 7483 10303 7535 10337
rect 7569 10303 7621 10337
rect 7655 10303 7707 10337
rect 7741 10303 7793 10337
rect 7827 10303 7879 10337
rect 7913 10303 7965 10337
rect 7999 10303 8051 10337
rect 8085 10303 8137 10337
rect 8171 10303 8222 10337
rect 8256 10303 8307 10337
rect 8341 10303 8392 10337
rect 8426 10303 8477 10337
rect 8511 10303 8562 10337
rect 8596 10303 8647 10337
rect 8681 10303 8732 10337
rect 8766 10303 8817 10337
rect 8851 10303 8902 10337
rect 8936 10303 8987 10337
rect 9021 10303 9072 10337
rect 9106 10303 9157 10337
rect 9191 10303 9242 10337
rect 9276 10303 9327 10337
rect 9361 10303 9412 10337
rect 9446 10303 9497 10337
rect 9531 10303 9582 10337
rect 9616 10303 9667 10337
rect 9701 10303 9752 10337
rect 9786 10303 9837 10337
rect 9871 10303 9922 10337
rect 9956 10303 10007 10337
rect 10041 10303 10092 10337
rect 10126 10303 10177 10337
rect 10211 10303 10262 10337
rect 10296 10303 10347 10337
rect 10381 10303 10432 10337
rect 10466 10303 10517 10337
rect 10551 10303 10602 10337
rect 10636 10303 10687 10337
rect 10721 10303 10772 10337
rect 10806 10303 10857 10337
rect 10891 10303 10942 10337
rect 10976 10303 11027 10337
rect 11061 10303 11112 10337
rect 11146 10303 11197 10337
rect 11231 10303 11282 10337
rect 11316 10303 11367 10337
rect 11401 10303 11452 10337
rect 11486 10303 11537 10337
rect 11571 10303 11622 10337
rect 11656 10303 11741 10337
rect 6356 10301 11741 10303
rect 6318 10299 11741 10301
rect 6318 10249 6360 10299
rect 6318 10215 6322 10249
rect 6356 10215 6360 10249
rect 6318 10163 6360 10215
rect 6318 10129 6322 10163
rect 6356 10129 6360 10163
rect 6318 10077 6360 10129
rect 6318 10043 6322 10077
rect 6356 10043 6360 10077
rect 6318 9991 6360 10043
rect 6318 9957 6322 9991
rect 6356 9957 6360 9991
rect 6318 9905 6360 9957
rect 6318 9871 6322 9905
rect 6356 9871 6360 9905
rect 6318 9819 6360 9871
rect 6318 9785 6322 9819
rect 6356 9785 6360 9819
rect 6318 9733 6360 9785
rect 6318 9699 6322 9733
rect 6356 9699 6360 9733
rect 6318 9647 6360 9699
rect 6318 9613 6322 9647
rect 6356 9613 6360 9647
rect 6318 9561 6360 9613
rect 10029 10238 10071 10299
rect 10029 10204 10033 10238
rect 10067 10204 10071 10238
rect 10029 10153 10071 10204
rect 10029 10119 10033 10153
rect 10067 10119 10071 10153
rect 10029 10068 10071 10119
rect 10029 10034 10033 10068
rect 10067 10034 10071 10068
rect 10029 9983 10071 10034
rect 10029 9949 10033 9983
rect 10067 9949 10071 9983
rect 10029 9898 10071 9949
rect 10029 9864 10033 9898
rect 10067 9864 10071 9898
rect 10029 9812 10071 9864
rect 10029 9778 10033 9812
rect 10067 9778 10071 9812
rect 10029 9726 10071 9778
rect 10029 9692 10033 9726
rect 10067 9692 10071 9726
rect 10029 9640 10071 9692
rect 10029 9606 10033 9640
rect 10067 9606 10071 9640
rect 6318 9527 6322 9561
rect 6356 9527 6360 9561
rect 6318 9475 6360 9527
rect 10029 9554 10071 9606
rect 10029 9520 10033 9554
rect 10067 9520 10071 9554
rect 6318 9441 6322 9475
rect 6356 9441 6360 9475
rect 6318 9389 6360 9441
rect 6318 9355 6322 9389
rect 6356 9355 6360 9389
rect 6318 9303 6360 9355
rect 6318 9269 6322 9303
rect 6356 9269 6360 9303
rect 6318 9217 6360 9269
rect 6318 9183 6322 9217
rect 6356 9183 6360 9217
rect 6318 9131 6360 9183
rect 6318 9097 6322 9131
rect 6356 9097 6360 9131
rect 6318 9045 6360 9097
rect 6318 9011 6322 9045
rect 6356 9011 6360 9045
rect 6318 8959 6360 9011
rect 6318 8925 6322 8959
rect 6356 8925 6360 8959
rect 6318 8873 6360 8925
rect 6318 8839 6322 8873
rect 6356 8839 6360 8873
rect 6318 8787 6360 8839
rect 6318 8753 6322 8787
rect 6356 8782 6360 8787
rect 10029 9468 10071 9520
rect 10029 9434 10033 9468
rect 10067 9434 10071 9468
rect 10029 9382 10071 9434
rect 10029 9348 10033 9382
rect 10067 9348 10071 9382
rect 10029 9296 10071 9348
rect 10029 9262 10033 9296
rect 10067 9262 10071 9296
rect 10029 9210 10071 9262
rect 10029 9176 10033 9210
rect 10067 9176 10071 9210
rect 10029 9124 10071 9176
rect 10029 9090 10033 9124
rect 10067 9090 10071 9124
rect 10029 9038 10071 9090
rect 10029 9004 10033 9038
rect 10067 9004 10071 9038
rect 10029 8952 10071 9004
rect 10029 8918 10033 8952
rect 10067 8918 10071 8952
rect 10029 8866 10071 8918
rect 10029 8832 10033 8866
rect 10067 8832 10071 8866
rect 6356 8753 6409 8782
rect 6318 8729 6409 8753
rect 10029 8751 10071 8832
rect 4834 5117 12710 5118
rect 4834 5083 4868 5117
rect 4902 5083 4936 5117
rect 4970 5083 5004 5117
rect 5038 5083 5072 5117
rect 5106 5083 5140 5117
rect 5174 5083 5208 5117
rect 5242 5083 5276 5117
rect 5310 5083 5344 5117
rect 5378 5083 5412 5117
rect 5446 5083 5480 5117
rect 5514 5083 5548 5117
rect 5582 5083 5616 5117
rect 5650 5083 5684 5117
rect 5718 5083 5752 5117
rect 5786 5083 5820 5117
rect 5854 5083 5888 5117
rect 5922 5083 5956 5117
rect 5990 5083 6024 5117
rect 6058 5083 6092 5117
rect 6126 5083 6160 5117
rect 6194 5083 6228 5117
rect 6262 5083 6296 5117
rect 6330 5083 6364 5117
rect 6398 5083 6432 5117
rect 6466 5083 6500 5117
rect 6534 5083 6568 5117
rect 6602 5083 6636 5117
rect 6670 5083 6704 5117
rect 6738 5083 6772 5117
rect 6806 5083 6840 5117
rect 6874 5083 6908 5117
rect 6942 5083 6976 5117
rect 7010 5083 7044 5117
rect 7078 5083 7112 5117
rect 7146 5083 7180 5117
rect 7214 5083 7248 5117
rect 7282 5083 7316 5117
rect 7350 5083 7384 5117
rect 7418 5083 7452 5117
rect 7486 5083 7520 5117
rect 7554 5083 7588 5117
rect 7622 5083 7656 5117
rect 7690 5083 7724 5117
rect 7758 5083 7792 5117
rect 7826 5083 7860 5117
rect 7894 5083 7928 5117
rect 7962 5083 7996 5117
rect 8030 5083 8064 5117
rect 8098 5083 8132 5117
rect 8166 5083 8200 5117
rect 8234 5083 8268 5117
rect 8302 5083 8336 5117
rect 8370 5083 8404 5117
rect 8438 5083 8472 5117
rect 8506 5083 8540 5117
rect 8574 5083 8608 5117
rect 8642 5083 8676 5117
rect 8710 5083 8744 5117
rect 8778 5083 8812 5117
rect 8846 5083 8880 5117
rect 8914 5083 8948 5117
rect 8982 5083 9016 5117
rect 9050 5083 9084 5117
rect 9118 5083 9152 5117
rect 9186 5083 9220 5117
rect 9254 5083 9288 5117
rect 9322 5083 9356 5117
rect 9390 5083 9424 5117
rect 9458 5083 9492 5117
rect 9526 5083 9560 5117
rect 9594 5083 9628 5117
rect 9662 5083 9696 5117
rect 9730 5083 9764 5117
rect 9798 5083 9832 5117
rect 9866 5083 9900 5117
rect 9934 5083 9968 5117
rect 10002 5083 10036 5117
rect 10070 5083 10104 5117
rect 10138 5083 10172 5117
rect 10206 5083 10240 5117
rect 10274 5083 10308 5117
rect 10342 5083 10376 5117
rect 10410 5083 10444 5117
rect 10478 5083 10512 5117
rect 10546 5083 10580 5117
rect 10614 5083 10648 5117
rect 10682 5083 10716 5117
rect 10750 5083 10784 5117
rect 10818 5083 10852 5117
rect 10886 5083 10920 5117
rect 10954 5083 10988 5117
rect 11022 5083 11056 5117
rect 11090 5083 11124 5117
rect 11158 5083 11192 5117
rect 11226 5083 11260 5117
rect 11294 5083 11328 5117
rect 11362 5083 11396 5117
rect 11430 5083 11464 5117
rect 11498 5083 11532 5117
rect 11566 5083 11600 5117
rect 11634 5083 11668 5117
rect 11702 5083 11736 5117
rect 11770 5083 11804 5117
rect 11838 5083 11872 5117
rect 11906 5083 11940 5117
rect 11974 5083 12008 5117
rect 12042 5083 12076 5117
rect 12110 5083 12144 5117
rect 12178 5083 12212 5117
rect 12246 5083 12280 5117
rect 12314 5083 12348 5117
rect 12382 5083 12416 5117
rect 12450 5083 12484 5117
rect 12518 5083 12552 5117
rect 12586 5084 12710 5117
rect 12586 5083 12675 5084
rect 4834 5082 12675 5083
rect 4834 5037 4870 5082
rect 4834 5003 4835 5037
rect 4869 5003 4870 5037
rect 4834 4969 4870 5003
rect 4834 4935 4835 4969
rect 4869 4935 4870 4969
rect 4834 4901 4870 4935
rect 4834 4867 4835 4901
rect 4869 4867 4870 4901
rect 4834 4833 4870 4867
rect 4834 4799 4835 4833
rect 4869 4799 4870 4833
rect 4834 4765 4870 4799
rect 4834 4731 4835 4765
rect 4869 4731 4870 4765
rect 4834 4697 4870 4731
rect 4834 4663 4835 4697
rect 4869 4663 4870 4697
rect 4834 4629 4870 4663
rect 4834 4595 4835 4629
rect 4869 4595 4870 4629
rect 4834 4561 4870 4595
rect 4834 4527 4835 4561
rect 4869 4527 4870 4561
rect 4834 4493 4870 4527
rect 9467 4987 9503 5082
rect 10296 5046 10330 5082
rect 9467 4953 9468 4987
rect 9502 4953 9503 4987
rect 9467 4919 9503 4953
rect 10296 4978 10330 5012
rect 9467 4885 9468 4919
rect 9502 4885 9503 4919
rect 9467 4851 9503 4885
rect 9467 4817 9468 4851
rect 9502 4817 9503 4851
rect 9467 4783 9503 4817
rect 9467 4749 9468 4783
rect 9502 4749 9503 4783
rect 9467 4715 9503 4749
rect 9467 4681 9468 4715
rect 9502 4681 9503 4715
rect 9467 4647 9503 4681
rect 9467 4613 9468 4647
rect 9502 4613 9503 4647
rect 9467 4579 9503 4613
rect 9467 4545 9468 4579
rect 9502 4545 9503 4579
rect 9467 4511 9503 4545
rect 4834 4459 4835 4493
rect 4869 4459 4870 4493
rect 4834 4425 4870 4459
rect 9467 4477 9468 4511
rect 9502 4477 9503 4511
rect 9467 4443 9503 4477
rect 4834 4391 4835 4425
rect 4869 4391 4870 4425
rect 4834 4357 4870 4391
rect 9467 4409 9468 4443
rect 9502 4409 9503 4443
rect 4834 4323 4835 4357
rect 4869 4323 4870 4357
rect 4834 4289 4870 4323
rect 9467 4375 9503 4409
rect 9467 4341 9468 4375
rect 9502 4341 9503 4375
rect 4834 4255 4835 4289
rect 4869 4255 4870 4289
rect 4834 4221 4870 4255
rect 4834 4187 4835 4221
rect 4869 4187 4870 4221
rect 4834 4153 4870 4187
rect 4834 4119 4835 4153
rect 4869 4119 4870 4153
rect 4834 4085 4870 4119
rect 4834 4051 4835 4085
rect 4869 4051 4870 4085
rect 4834 4017 4870 4051
rect 4834 3983 4835 4017
rect 4869 3983 4870 4017
rect 4834 3949 4870 3983
rect 4834 3915 4835 3949
rect 4869 3915 4870 3949
rect 4834 3881 4870 3915
rect 4834 3847 4835 3881
rect 4869 3847 4870 3881
rect 4834 3813 4870 3847
rect 4834 3779 4835 3813
rect 4869 3779 4870 3813
rect 4834 3745 4870 3779
rect 4834 3711 4835 3745
rect 4869 3744 4870 3745
rect 9467 4307 9503 4341
rect 9467 4273 9468 4307
rect 9502 4273 9503 4307
rect 9467 4239 9503 4273
rect 9467 4205 9468 4239
rect 9502 4205 9503 4239
rect 9467 4171 9503 4205
rect 9467 4137 9468 4171
rect 9502 4137 9503 4171
rect 9467 4103 9503 4137
rect 9467 4069 9468 4103
rect 9502 4069 9503 4103
rect 9467 4035 9503 4069
rect 9467 4001 9468 4035
rect 9502 4001 9503 4035
rect 9467 3967 9503 4001
rect 9467 3933 9468 3967
rect 9502 3933 9503 3967
rect 9467 3899 9503 3933
rect 9467 3865 9468 3899
rect 9502 3865 9503 3899
rect 9467 3831 9503 3865
rect 9467 3797 9468 3831
rect 9502 3797 9503 3831
rect 9467 3763 9503 3797
rect 9467 3744 9468 3763
rect 4869 3711 4963 3744
rect 4834 3710 4963 3711
rect 4997 3710 5032 3744
rect 5066 3710 5101 3744
rect 5135 3710 5170 3744
rect 5204 3710 5239 3744
rect 5273 3710 5308 3744
rect 5342 3710 5377 3744
rect 5411 3710 5446 3744
rect 5480 3710 5515 3744
rect 5549 3710 5584 3744
rect 5618 3710 5653 3744
rect 5687 3710 5722 3744
rect 5756 3710 5791 3744
rect 5825 3710 5860 3744
rect 5894 3710 5929 3744
rect 4834 3677 5929 3710
rect 4834 3643 4835 3677
rect 4869 3676 5929 3677
rect 4869 3643 4963 3676
rect 4834 3642 4963 3643
rect 4997 3642 5032 3676
rect 5066 3642 5101 3676
rect 5135 3642 5170 3676
rect 5204 3642 5239 3676
rect 5273 3642 5308 3676
rect 5342 3642 5377 3676
rect 5411 3642 5446 3676
rect 5480 3642 5515 3676
rect 5549 3642 5584 3676
rect 5618 3642 5653 3676
rect 5687 3642 5722 3676
rect 5756 3642 5791 3676
rect 5825 3642 5860 3676
rect 5894 3642 5929 3676
rect 9363 3729 9468 3744
rect 9502 3729 9503 3763
rect 9363 3695 9503 3729
rect 9363 3661 9468 3695
rect 9502 3661 9503 3695
rect 9363 3642 9503 3661
rect 4834 3609 4870 3642
rect 4834 3575 4835 3609
rect 4869 3575 4870 3609
rect 4834 3541 4870 3575
rect 4834 3507 4835 3541
rect 4869 3507 4870 3541
rect 4834 3473 4870 3507
rect 9467 3627 9503 3642
rect 9467 3593 9468 3627
rect 9502 3593 9503 3627
rect 9467 3559 9503 3593
rect 9467 3525 9468 3559
rect 9502 3525 9503 3559
rect 9467 3491 9503 3525
rect 4834 3439 4835 3473
rect 4869 3439 4870 3473
rect 4834 3405 4870 3439
rect 4834 3371 4835 3405
rect 4869 3371 4870 3405
rect 4834 3337 4870 3371
rect 4834 3303 4835 3337
rect 4869 3303 4870 3337
rect 9467 3457 9468 3491
rect 9502 3457 9503 3491
rect 9467 3423 9503 3457
rect 9467 3389 9468 3423
rect 9502 3389 9503 3423
rect 9467 3355 9503 3389
rect 9467 3321 9468 3355
rect 9502 3321 9503 3355
rect 4834 3269 4870 3303
rect 4834 3235 4835 3269
rect 4869 3235 4870 3269
rect 4834 3201 4870 3235
rect 4834 3167 4835 3201
rect 4869 3167 4870 3201
rect 4834 3133 4870 3167
rect 4834 3099 4835 3133
rect 4869 3099 4870 3133
rect 9467 3287 9503 3321
rect 9467 3253 9468 3287
rect 9502 3253 9503 3287
rect 9467 3219 9503 3253
rect 9467 3185 9468 3219
rect 9502 3185 9503 3219
rect 9467 3151 9503 3185
rect 4834 3065 4870 3099
rect 4834 3031 4835 3065
rect 4869 3031 4870 3065
rect 4834 2997 4870 3031
rect 4834 2963 4835 2997
rect 4869 2963 4870 2997
rect 4834 2929 4870 2963
rect 9467 3117 9468 3151
rect 9502 3117 9503 3151
rect 9467 3083 9503 3117
rect 9467 3049 9468 3083
rect 9502 3049 9503 3083
rect 9467 3015 9503 3049
rect 9467 2981 9468 3015
rect 9502 2981 9503 3015
rect 4834 2895 4835 2929
rect 4869 2895 4870 2929
rect 9467 2947 9503 2981
rect 9467 2913 9468 2947
rect 9502 2913 9503 2947
rect 4834 2861 4870 2895
rect 4834 2827 4835 2861
rect 4869 2827 4870 2861
rect 4834 2793 4870 2827
rect 4834 2759 4835 2793
rect 4869 2759 4870 2793
rect 4834 2725 4870 2759
rect 4834 2691 4835 2725
rect 4869 2691 4870 2725
rect 9467 2879 9503 2913
rect 9467 2845 9468 2879
rect 9502 2845 9503 2879
rect 9467 2811 9503 2845
rect 9467 2777 9468 2811
rect 9502 2777 9503 2811
rect 9467 2743 9503 2777
rect 4834 2657 4870 2691
rect 4834 2623 4835 2657
rect 4869 2623 4870 2657
rect 4834 2589 4870 2623
rect 4834 2555 4835 2589
rect 4869 2555 4870 2589
rect 4834 2521 4870 2555
rect 9467 2709 9468 2743
rect 9502 2709 9503 2743
rect 9467 2675 9503 2709
rect 9467 2641 9468 2675
rect 9502 2641 9503 2675
rect 9467 2607 9503 2641
rect 9467 2573 9468 2607
rect 9502 2573 9503 2607
rect 9467 2539 9503 2573
rect 4834 2487 4835 2521
rect 4869 2487 4870 2521
rect 4834 2453 4870 2487
rect 4834 2419 4835 2453
rect 4869 2419 4870 2453
rect 4834 2385 4870 2419
rect 4834 2351 4835 2385
rect 4869 2351 4870 2385
rect 9467 2505 9468 2539
rect 9502 2505 9503 2539
rect 9467 2471 9503 2505
rect 9467 2437 9468 2471
rect 9502 2437 9503 2471
rect 9467 2402 9503 2437
rect 9467 2368 9468 2402
rect 9502 2368 9503 2402
rect 4834 2317 4870 2351
rect 4834 2283 4835 2317
rect 4869 2283 4870 2317
rect 9467 2333 9503 2368
rect 9467 2299 9468 2333
rect 9502 2299 9503 2333
rect 4834 2249 4870 2283
rect 4834 2215 4835 2249
rect 4869 2215 4870 2249
rect 4834 2181 4870 2215
rect 4834 2147 4835 2181
rect 4869 2147 4870 2181
rect 4834 2113 4870 2147
rect 9467 2264 9503 2299
rect 9467 2230 9468 2264
rect 9502 2230 9503 2264
rect 9467 2195 9503 2230
rect 9467 2161 9468 2195
rect 9502 2161 9503 2195
rect 9467 2126 9503 2161
rect 4834 2079 4835 2113
rect 4869 2079 4870 2113
rect 4834 2045 4870 2079
rect 4834 2011 4835 2045
rect 4869 2011 4870 2045
rect 4834 1977 4870 2011
rect 4834 1943 4835 1977
rect 4869 1943 4870 1977
rect 4834 1909 4870 1943
rect 9467 2092 9468 2126
rect 9502 2092 9503 2126
rect 9467 2057 9503 2092
rect 9467 2023 9468 2057
rect 9502 2023 9503 2057
rect 9467 1988 9503 2023
rect 9467 1954 9468 1988
rect 9502 1954 9503 1988
rect 4834 1875 4835 1909
rect 4869 1875 4870 1909
rect 4834 1841 4870 1875
rect 4834 1807 4835 1841
rect 4869 1807 4870 1841
rect 4834 1773 4870 1807
rect 4834 1739 4835 1773
rect 4869 1739 4870 1773
rect 9467 1919 9503 1954
rect 9467 1885 9468 1919
rect 9502 1885 9503 1919
rect 9467 1850 9503 1885
rect 9467 1816 9468 1850
rect 9502 1816 9503 1850
rect 9467 1781 9503 1816
rect 4834 1705 4870 1739
rect 4834 1671 4835 1705
rect 4869 1671 4870 1705
rect 4834 1637 4870 1671
rect 4834 1603 4835 1637
rect 4869 1605 4870 1637
rect 9467 1747 9468 1781
rect 9502 1747 9503 1781
rect 9467 1712 9503 1747
rect 9467 1678 9468 1712
rect 9502 1678 9503 1712
rect 9467 1643 9503 1678
rect 9467 1609 9468 1643
rect 9502 1609 9503 1643
rect 9467 1605 9503 1609
rect 4869 1603 4963 1605
rect 4834 1571 4963 1603
rect 4997 1571 5032 1605
rect 5066 1571 5101 1605
rect 5135 1571 5170 1605
rect 5204 1571 5239 1605
rect 5273 1571 5308 1605
rect 5342 1571 5377 1605
rect 5411 1571 5446 1605
rect 5480 1571 5515 1605
rect 5549 1571 5584 1605
rect 5618 1571 5653 1605
rect 5687 1571 5722 1605
rect 5756 1571 5791 1605
rect 5825 1571 5860 1605
rect 5894 1571 5929 1605
rect 4834 1569 5929 1571
rect 4834 1535 4835 1569
rect 4869 1537 5929 1569
rect 4869 1535 4963 1537
rect 4834 1503 4963 1535
rect 4997 1503 5032 1537
rect 5066 1503 5101 1537
rect 5135 1503 5170 1537
rect 5204 1503 5239 1537
rect 5273 1503 5308 1537
rect 5342 1503 5377 1537
rect 5411 1503 5446 1537
rect 5480 1503 5515 1537
rect 5549 1503 5584 1537
rect 5618 1503 5653 1537
rect 5687 1503 5722 1537
rect 5756 1503 5791 1537
rect 5825 1503 5860 1537
rect 5894 1503 5929 1537
rect 9363 1574 9503 1605
rect 9363 1540 9468 1574
rect 9502 1540 9503 1574
rect 9363 1505 9503 1540
rect 9363 1503 9468 1505
rect 4834 1501 4870 1503
rect 4834 1467 4835 1501
rect 4869 1467 4870 1501
rect 4834 1433 4870 1467
rect 4834 1399 4835 1433
rect 4869 1399 4870 1433
rect 4834 1365 4870 1399
rect 4834 1331 4835 1365
rect 4869 1331 4870 1365
rect 4834 1297 4870 1331
rect 4834 1263 4835 1297
rect 4869 1263 4870 1297
rect 4834 1229 4870 1263
rect 4834 1195 4835 1229
rect 4869 1195 4870 1229
rect 4834 1161 4870 1195
rect 4834 1127 4835 1161
rect 4869 1127 4870 1161
rect 4834 1093 4870 1127
rect 4834 1059 4835 1093
rect 4869 1059 4870 1093
rect 4834 1025 4870 1059
rect 9467 1471 9468 1503
rect 9502 1471 9503 1505
rect 9467 1436 9503 1471
rect 9467 1402 9468 1436
rect 9502 1402 9503 1436
rect 9467 1367 9503 1402
rect 9467 1333 9468 1367
rect 9502 1333 9503 1367
rect 9467 1298 9503 1333
rect 9467 1264 9468 1298
rect 9502 1264 9503 1298
rect 9467 1229 9503 1264
rect 9467 1195 9468 1229
rect 9502 1195 9503 1229
rect 9467 1160 9503 1195
rect 9467 1126 9468 1160
rect 9502 1126 9503 1160
rect 9467 1091 9503 1126
rect 9467 1057 9468 1091
rect 9502 1057 9503 1091
rect 4834 991 4835 1025
rect 4869 991 4870 1025
rect 4834 957 4870 991
rect 9467 1022 9503 1057
rect 9467 988 9468 1022
rect 9502 988 9503 1022
rect 4834 923 4835 957
rect 4869 923 4870 957
rect 4834 889 4870 923
rect 9467 953 9503 988
rect 9467 919 9468 953
rect 9502 919 9503 953
rect 4834 855 4835 889
rect 4869 855 4870 889
rect 4834 821 4870 855
rect 9467 884 9503 919
rect 9467 850 9468 884
rect 9502 850 9503 884
rect 4834 787 4835 821
rect 4869 787 4870 821
rect 4834 753 4870 787
rect 4834 719 4835 753
rect 4869 719 4870 753
rect 4834 685 4870 719
rect 4834 651 4835 685
rect 4869 651 4870 685
rect 4834 617 4870 651
rect 4834 583 4835 617
rect 4869 583 4870 617
rect 4834 549 4870 583
rect 4834 515 4835 549
rect 4869 515 4870 549
rect 4834 481 4870 515
rect 4834 447 4835 481
rect 4869 447 4870 481
rect 4834 413 4870 447
rect 4834 379 4835 413
rect 4869 379 4870 413
rect 4834 345 4870 379
rect 4834 311 4835 345
rect 4869 311 4870 345
rect 4834 277 4870 311
rect 4834 243 4835 277
rect 4869 245 4870 277
rect 9467 815 9503 850
rect 9467 781 9468 815
rect 9502 781 9503 815
rect 9467 746 9503 781
rect 9467 712 9468 746
rect 9502 712 9503 746
rect 9467 677 9503 712
rect 9467 643 9468 677
rect 9502 643 9503 677
rect 9467 608 9503 643
rect 10296 4910 10330 4944
rect 10296 4842 10330 4876
rect 12674 5050 12675 5082
rect 12709 5050 12710 5084
rect 12674 5016 12710 5050
rect 12674 4982 12675 5016
rect 12709 4982 12710 5016
rect 12674 4948 12710 4982
rect 12674 4914 12675 4948
rect 12709 4914 12710 4948
rect 12674 4880 12710 4914
rect 10296 4774 10330 4808
rect 10296 4706 10330 4740
rect 10296 4638 10330 4672
rect 10296 4570 10330 4604
rect 10296 4502 10330 4536
rect 10296 4434 10330 4468
rect 10296 4366 10330 4400
rect 10296 4298 10330 4332
rect 10296 4230 10330 4264
rect 10296 4162 10330 4196
rect 10296 4094 10330 4128
rect 10296 4026 10330 4060
rect 12674 4846 12675 4880
rect 12709 4846 12710 4880
rect 12674 4812 12710 4846
rect 12674 4778 12675 4812
rect 12709 4778 12710 4812
rect 12674 4744 12710 4778
rect 12674 4710 12675 4744
rect 12709 4710 12710 4744
rect 12674 4676 12710 4710
rect 12674 4642 12675 4676
rect 12709 4642 12710 4676
rect 12674 4608 12710 4642
rect 12674 4574 12675 4608
rect 12709 4574 12710 4608
rect 12674 4540 12710 4574
rect 12674 4506 12675 4540
rect 12709 4506 12710 4540
rect 12674 4472 12710 4506
rect 12674 4438 12675 4472
rect 12709 4438 12710 4472
rect 12674 4404 12710 4438
rect 12674 4370 12675 4404
rect 12709 4370 12710 4404
rect 12674 4336 12710 4370
rect 12674 4302 12675 4336
rect 12709 4302 12710 4336
rect 12674 4268 12710 4302
rect 12674 4234 12675 4268
rect 12709 4234 12710 4268
rect 12674 4200 12710 4234
rect 12674 4166 12675 4200
rect 12709 4166 12710 4200
rect 12674 4132 12710 4166
rect 12674 4098 12675 4132
rect 12709 4098 12710 4132
rect 12674 4064 12710 4098
rect 12674 4030 12675 4064
rect 12709 4030 12710 4064
rect 10296 3958 10330 3992
rect 10296 3890 10330 3924
rect 10296 3822 10330 3856
rect 10296 3754 10330 3788
rect 10296 3686 10330 3720
rect 10296 3618 10330 3652
rect 10296 3550 10330 3584
rect 12674 3996 12710 4030
rect 12674 3962 12675 3996
rect 12709 3962 12710 3996
rect 12674 3928 12710 3962
rect 12674 3894 12675 3928
rect 12709 3894 12710 3928
rect 12674 3860 12710 3894
rect 12674 3826 12675 3860
rect 12709 3826 12710 3860
rect 12674 3792 12710 3826
rect 12674 3758 12675 3792
rect 12709 3758 12710 3792
rect 12674 3724 12710 3758
rect 12674 3690 12675 3724
rect 12709 3690 12710 3724
rect 12674 3656 12710 3690
rect 12674 3622 12675 3656
rect 12709 3622 12710 3656
rect 12674 3588 12710 3622
rect 12674 3554 12675 3588
rect 12709 3554 12710 3588
rect 10296 3482 10330 3516
rect 12674 3520 12710 3554
rect 10296 3414 10330 3448
rect 10296 3346 10330 3380
rect 10296 3278 10330 3312
rect 12674 3486 12675 3520
rect 12709 3486 12710 3520
rect 12674 3452 12710 3486
rect 12674 3418 12675 3452
rect 12709 3418 12710 3452
rect 12674 3384 12710 3418
rect 12674 3350 12675 3384
rect 12709 3350 12710 3384
rect 12674 3316 12710 3350
rect 10296 3210 10330 3244
rect 12674 3282 12675 3316
rect 12709 3282 12710 3316
rect 12674 3248 12710 3282
rect 10296 3142 10330 3176
rect 10296 3074 10330 3108
rect 10296 3006 10330 3040
rect 12674 3214 12675 3248
rect 12709 3214 12710 3248
rect 12674 3180 12710 3214
rect 12674 3146 12675 3180
rect 12709 3146 12710 3180
rect 12674 3112 12710 3146
rect 12674 3078 12675 3112
rect 12709 3078 12710 3112
rect 12674 3044 12710 3078
rect 12674 3010 12675 3044
rect 12709 3010 12710 3044
rect 10296 2938 10330 2972
rect 10296 2870 10330 2904
rect 10296 2802 10330 2836
rect 12674 2976 12710 3010
rect 12674 2942 12675 2976
rect 12709 2942 12710 2976
rect 12674 2908 12710 2942
rect 12674 2874 12675 2908
rect 12709 2874 12710 2908
rect 12674 2840 12710 2874
rect 12674 2806 12675 2840
rect 12709 2806 12710 2840
rect 10296 2734 10330 2768
rect 12674 2772 12710 2806
rect 12674 2738 12675 2772
rect 12709 2738 12710 2772
rect 10296 2666 10330 2700
rect 10296 2598 10330 2632
rect 10296 2530 10330 2564
rect 12674 2704 12710 2738
rect 12674 2670 12675 2704
rect 12709 2670 12710 2704
rect 12674 2636 12710 2670
rect 12674 2602 12675 2636
rect 12709 2602 12710 2636
rect 12674 2568 12710 2602
rect 12674 2534 12675 2568
rect 12709 2534 12710 2568
rect 10296 2462 10330 2496
rect 12674 2500 12710 2534
rect 12674 2466 12675 2500
rect 12709 2466 12710 2500
rect 10296 2394 10330 2428
rect 10296 2326 10330 2360
rect 10296 2258 10330 2292
rect 12674 2432 12710 2466
rect 12674 2398 12675 2432
rect 12709 2398 12710 2432
rect 12674 2364 12710 2398
rect 12674 2330 12675 2364
rect 12709 2330 12710 2364
rect 12674 2296 12710 2330
rect 10296 2190 10330 2224
rect 12674 2262 12675 2296
rect 12709 2262 12710 2296
rect 12674 2228 12710 2262
rect 10296 2122 10330 2156
rect 10296 2054 10330 2088
rect 10296 1986 10330 2020
rect 12674 2194 12675 2228
rect 12709 2194 12710 2228
rect 12674 2160 12710 2194
rect 12674 2126 12675 2160
rect 12709 2126 12710 2160
rect 12674 2092 12710 2126
rect 12674 2058 12675 2092
rect 12709 2058 12710 2092
rect 12674 2024 12710 2058
rect 12674 1990 12675 2024
rect 12709 1990 12710 2024
rect 12674 1956 12710 1990
rect 10296 1918 10330 1952
rect 10296 1850 10330 1884
rect 10296 1782 10330 1816
rect 12674 1922 12675 1956
rect 12709 1922 12710 1956
rect 12674 1888 12710 1922
rect 12674 1854 12675 1888
rect 12709 1854 12710 1888
rect 12674 1820 12710 1854
rect 12674 1786 12675 1820
rect 12709 1786 12710 1820
rect 10296 1714 10330 1748
rect 12674 1752 12710 1786
rect 12674 1718 12675 1752
rect 12709 1718 12710 1752
rect 10296 1646 10330 1680
rect 10296 1578 10330 1612
rect 10296 1510 10330 1544
rect 12674 1684 12710 1718
rect 12674 1650 12675 1684
rect 12709 1650 12710 1684
rect 12674 1616 12710 1650
rect 12674 1582 12675 1616
rect 12709 1582 12710 1616
rect 12674 1548 12710 1582
rect 12674 1514 12675 1548
rect 12709 1514 12710 1548
rect 10296 1442 10330 1476
rect 12674 1480 12710 1514
rect 12674 1446 12675 1480
rect 12709 1446 12710 1480
rect 10296 1374 10330 1408
rect 10296 1306 10330 1340
rect 10296 1238 10330 1272
rect 10296 1170 10330 1204
rect 10296 1102 10330 1136
rect 10296 1034 10330 1068
rect 10296 966 10330 1000
rect 10296 898 10330 932
rect 10296 830 10330 864
rect 10296 762 10330 796
rect 10296 694 10330 728
rect 9467 574 9468 608
rect 9502 574 9503 608
rect 9467 539 9503 574
rect 10296 626 10330 660
rect 12674 1412 12710 1446
rect 12674 1378 12675 1412
rect 12709 1378 12710 1412
rect 12674 1344 12710 1378
rect 12674 1310 12675 1344
rect 12709 1310 12710 1344
rect 12674 1276 12710 1310
rect 12674 1242 12675 1276
rect 12709 1242 12710 1276
rect 12674 1208 12710 1242
rect 12674 1174 12675 1208
rect 12709 1174 12710 1208
rect 12674 1140 12710 1174
rect 12674 1106 12675 1140
rect 12709 1106 12710 1140
rect 12674 1072 12710 1106
rect 12674 1038 12675 1072
rect 12709 1038 12710 1072
rect 12674 1004 12710 1038
rect 12674 970 12675 1004
rect 12709 970 12710 1004
rect 12674 936 12710 970
rect 12674 902 12675 936
rect 12709 902 12710 936
rect 12674 868 12710 902
rect 12674 834 12675 868
rect 12709 834 12710 868
rect 12674 800 12710 834
rect 12674 766 12675 800
rect 12709 766 12710 800
rect 12674 732 12710 766
rect 12674 698 12675 732
rect 12709 698 12710 732
rect 10296 558 10330 592
rect 9467 505 9468 539
rect 9502 505 9503 539
rect 9467 490 9503 505
rect 10296 490 10330 524
rect 12674 608 12710 698
rect 12674 574 12675 608
rect 12709 574 12710 608
rect 12674 490 12710 574
rect 9467 489 12710 490
rect 9467 470 9582 489
rect 9467 436 9468 470
rect 9502 455 9582 470
rect 9616 455 9650 489
rect 9684 455 9718 489
rect 9752 455 9786 489
rect 9820 455 9854 489
rect 9888 455 9922 489
rect 9956 455 9990 489
rect 10024 455 10058 489
rect 10092 455 10126 489
rect 10160 455 10194 489
rect 10228 455 10262 489
rect 10296 455 10330 489
rect 10364 455 10398 489
rect 10432 455 10466 489
rect 10500 455 10534 489
rect 10568 455 10602 489
rect 10636 455 10670 489
rect 10704 455 10738 489
rect 10772 455 10806 489
rect 10840 455 10874 489
rect 10908 455 10942 489
rect 10976 455 11010 489
rect 11044 455 11078 489
rect 11112 455 11146 489
rect 11180 455 11214 489
rect 11248 455 11282 489
rect 11316 455 11350 489
rect 11384 455 11418 489
rect 11452 455 11486 489
rect 11520 455 11554 489
rect 11588 455 11622 489
rect 11656 455 11690 489
rect 11724 455 11758 489
rect 11792 455 11826 489
rect 11860 455 11894 489
rect 11928 455 11962 489
rect 11996 455 12030 489
rect 12064 455 12098 489
rect 12132 455 12166 489
rect 12200 455 12234 489
rect 12268 455 12302 489
rect 12336 455 12370 489
rect 12404 455 12438 489
rect 12472 455 12506 489
rect 12540 455 12574 489
rect 12608 455 12642 489
rect 12676 455 12710 489
rect 9502 454 12710 455
rect 9502 436 9503 454
rect 9467 401 9503 436
rect 9467 367 9468 401
rect 9502 367 9503 401
rect 9467 332 9503 367
rect 9467 298 9468 332
rect 9502 298 9503 332
rect 9467 245 9503 298
rect 4869 244 9503 245
rect 4869 243 4947 244
rect 4834 210 4947 243
rect 4981 210 5015 244
rect 5049 210 5083 244
rect 5117 210 5151 244
rect 5185 210 5219 244
rect 5253 210 5287 244
rect 5321 210 5355 244
rect 5389 210 5423 244
rect 5457 210 5491 244
rect 5525 210 5559 244
rect 5593 210 5627 244
rect 5661 210 5695 244
rect 5729 210 5763 244
rect 5797 210 5831 244
rect 5865 210 5899 244
rect 5933 210 5967 244
rect 6001 210 6035 244
rect 6069 210 6103 244
rect 6137 210 6171 244
rect 6205 210 6239 244
rect 6273 210 6307 244
rect 6341 210 6375 244
rect 6409 210 6443 244
rect 6477 210 6511 244
rect 6545 210 6579 244
rect 6613 210 6647 244
rect 6681 210 6715 244
rect 6749 210 6783 244
rect 6817 210 6851 244
rect 6885 210 6919 244
rect 6953 210 6987 244
rect 7021 210 7055 244
rect 7089 210 7123 244
rect 7157 210 7191 244
rect 7225 210 7259 244
rect 7293 210 7327 244
rect 7361 210 7395 244
rect 7429 210 7463 244
rect 7497 210 7531 244
rect 7565 210 7599 244
rect 7633 210 7667 244
rect 7701 210 7735 244
rect 7769 210 7803 244
rect 7837 210 7871 244
rect 7905 210 7939 244
rect 7973 210 8007 244
rect 8041 210 8075 244
rect 8109 210 8143 244
rect 8177 210 8211 244
rect 8245 210 8279 244
rect 8313 210 8347 244
rect 8381 210 8415 244
rect 8449 210 8483 244
rect 8517 210 8551 244
rect 8585 210 8619 244
rect 8653 210 8687 244
rect 8721 210 8755 244
rect 8789 210 8823 244
rect 8857 210 8891 244
rect 8925 210 8959 244
rect 8993 210 9027 244
rect 9061 210 9095 244
rect 9129 210 9163 244
rect 9197 210 9231 244
rect 9265 210 9299 244
rect 9333 210 9367 244
rect 9401 210 9435 244
rect 9469 210 9503 244
rect 4834 209 9503 210
<< mvnsubdiff >>
rect 8574 6945 13682 6946
rect 8574 6911 8608 6945
rect 8642 6911 8676 6945
rect 8710 6911 8744 6945
rect 8778 6911 8812 6945
rect 8846 6911 8880 6945
rect 8914 6911 8948 6945
rect 8982 6911 9016 6945
rect 9050 6911 9084 6945
rect 9118 6911 9152 6945
rect 9186 6911 9220 6945
rect 9254 6911 9288 6945
rect 9322 6911 9356 6945
rect 9390 6911 9424 6945
rect 9458 6911 9492 6945
rect 9526 6911 9560 6945
rect 9594 6911 9628 6945
rect 9662 6911 9696 6945
rect 9730 6911 9764 6945
rect 9798 6911 9832 6945
rect 9866 6911 9900 6945
rect 9934 6911 9968 6945
rect 10002 6911 10036 6945
rect 10070 6911 10104 6945
rect 10138 6911 10172 6945
rect 10206 6911 10240 6945
rect 10274 6911 10308 6945
rect 10342 6911 10376 6945
rect 10410 6911 10444 6945
rect 10478 6911 10512 6945
rect 10546 6911 10580 6945
rect 10614 6911 10648 6945
rect 10682 6911 10716 6945
rect 10750 6911 10784 6945
rect 10818 6911 10852 6945
rect 10886 6911 10920 6945
rect 10954 6911 10988 6945
rect 11022 6911 11056 6945
rect 11090 6911 11124 6945
rect 11158 6911 11192 6945
rect 11226 6911 11260 6945
rect 11294 6911 11328 6945
rect 11362 6911 11396 6945
rect 11430 6911 11464 6945
rect 11498 6911 11532 6945
rect 11566 6911 11600 6945
rect 11634 6911 11668 6945
rect 11702 6911 11736 6945
rect 11770 6911 11804 6945
rect 11838 6911 11872 6945
rect 11906 6911 11940 6945
rect 11974 6911 12008 6945
rect 12042 6911 12076 6945
rect 12110 6911 12144 6945
rect 12178 6911 12212 6945
rect 12246 6911 12280 6945
rect 12314 6911 12348 6945
rect 12382 6911 12416 6945
rect 12450 6911 12484 6945
rect 12518 6911 12552 6945
rect 12586 6911 12620 6945
rect 12654 6911 12688 6945
rect 12722 6911 12756 6945
rect 12790 6911 12824 6945
rect 12858 6911 12892 6945
rect 12926 6911 12960 6945
rect 12994 6911 13028 6945
rect 13062 6911 13096 6945
rect 13130 6911 13164 6945
rect 13198 6911 13232 6945
rect 13266 6911 13300 6945
rect 13334 6911 13368 6945
rect 13402 6911 13436 6945
rect 13470 6911 13504 6945
rect 13538 6911 13572 6945
rect 13606 6912 13682 6945
rect 13606 6911 13647 6912
rect 8574 6910 13647 6911
rect 8574 6877 8610 6910
rect 8574 6843 8575 6877
rect 8609 6843 8610 6877
rect 8574 6809 8610 6843
rect 8574 6775 8575 6809
rect 8609 6775 8610 6809
rect 8574 6741 8610 6775
rect 8574 6707 8575 6741
rect 8609 6707 8610 6741
rect 8574 6673 8610 6707
rect 8574 6639 8575 6673
rect 8609 6639 8610 6673
rect 8574 6605 8610 6639
rect 8574 6571 8575 6605
rect 8609 6571 8610 6605
rect 8574 6537 8610 6571
rect 8574 6503 8575 6537
rect 8609 6503 8610 6537
rect 8574 6469 8610 6503
rect 8574 6435 8575 6469
rect 8609 6435 8610 6469
rect 8574 6401 8610 6435
rect 8574 6367 8575 6401
rect 8609 6367 8610 6401
rect 8574 6333 8610 6367
rect 8574 6301 8575 6333
rect 4645 6300 8575 6301
rect 4645 6266 4679 6300
rect 4713 6266 4747 6300
rect 4781 6266 4815 6300
rect 4849 6266 4883 6300
rect 4917 6266 4951 6300
rect 4985 6266 5019 6300
rect 5053 6266 5087 6300
rect 5121 6266 5155 6300
rect 5189 6266 5223 6300
rect 5257 6266 5291 6300
rect 5325 6266 5359 6300
rect 5393 6266 5427 6300
rect 5461 6266 5495 6300
rect 5529 6266 5563 6300
rect 5597 6266 5631 6300
rect 5665 6266 5699 6300
rect 5733 6266 5767 6300
rect 5801 6266 5835 6300
rect 5869 6266 5903 6300
rect 5937 6266 5971 6300
rect 6005 6266 6039 6300
rect 6073 6266 6107 6300
rect 6141 6266 6175 6300
rect 6209 6266 6243 6300
rect 6277 6266 6311 6300
rect 6345 6266 6379 6300
rect 6413 6266 6447 6300
rect 6481 6266 6515 6300
rect 6549 6266 6583 6300
rect 6617 6266 6651 6300
rect 6685 6266 6719 6300
rect 6753 6266 6787 6300
rect 6821 6266 6855 6300
rect 6889 6266 6923 6300
rect 6957 6266 6991 6300
rect 7025 6266 7059 6300
rect 7093 6266 7127 6300
rect 7161 6266 7195 6300
rect 7229 6266 7263 6300
rect 7297 6266 7331 6300
rect 7365 6266 7399 6300
rect 7433 6266 7467 6300
rect 7501 6266 7535 6300
rect 7569 6266 7603 6300
rect 7637 6266 7671 6300
rect 7705 6266 7739 6300
rect 7773 6266 7807 6300
rect 7841 6266 7875 6300
rect 7909 6266 7943 6300
rect 7977 6266 8011 6300
rect 8045 6266 8079 6300
rect 8113 6266 8147 6300
rect 8181 6266 8215 6300
rect 8249 6266 8283 6300
rect 8317 6266 8351 6300
rect 8385 6266 8419 6300
rect 8453 6266 8487 6300
rect 8521 6299 8575 6300
rect 8609 6299 8610 6333
rect 8521 6266 8610 6299
rect 4645 6265 8610 6266
rect 13646 6878 13647 6910
rect 13681 6878 13682 6912
rect 13646 6844 13682 6878
rect 13646 6810 13647 6844
rect 13681 6810 13682 6844
rect 13646 6776 13682 6810
rect 13646 6742 13647 6776
rect 13681 6742 13682 6776
rect 13646 6708 13682 6742
rect 13646 6674 13647 6708
rect 13681 6674 13682 6708
rect 13646 6640 13682 6674
rect 13646 6606 13647 6640
rect 13681 6606 13682 6640
rect 13646 6572 13682 6606
rect 13646 6538 13647 6572
rect 13681 6538 13682 6572
rect 13646 6504 13682 6538
rect 13646 6470 13647 6504
rect 13681 6470 13682 6504
rect 13646 6436 13682 6470
rect 13646 6402 13647 6436
rect 13681 6402 13682 6436
rect 13646 6368 13682 6402
rect 13646 6334 13647 6368
rect 13681 6334 13682 6368
rect 13646 6300 13682 6334
rect 13646 6266 13647 6300
rect 13681 6266 13682 6300
rect 249 6254 813 6255
rect 249 6220 283 6254
rect 317 6220 351 6254
rect 385 6220 419 6254
rect 453 6220 487 6254
rect 521 6220 555 6254
rect 589 6220 623 6254
rect 657 6220 691 6254
rect 725 6221 813 6254
rect 725 6220 778 6221
rect 249 6219 778 6220
rect 249 6139 285 6219
rect 249 6105 250 6139
rect 284 6105 285 6139
rect 249 6071 285 6105
rect 777 6187 778 6219
rect 812 6187 813 6221
rect 777 6153 813 6187
rect 777 6119 778 6153
rect 812 6119 813 6153
rect 249 6037 250 6071
rect 284 6037 285 6071
rect 249 6003 285 6037
rect 249 5969 250 6003
rect 284 5969 285 6003
rect 249 5935 285 5969
rect 249 5901 250 5935
rect 284 5901 285 5935
rect 249 5867 285 5901
rect 249 5833 250 5867
rect 284 5833 285 5867
rect 249 5799 285 5833
rect 249 5765 250 5799
rect 284 5765 285 5799
rect 249 5731 285 5765
rect 249 5697 250 5731
rect 284 5697 285 5731
rect 249 5663 285 5697
rect 249 5629 250 5663
rect 284 5629 285 5663
rect 249 5595 285 5629
rect 249 5561 250 5595
rect 284 5561 285 5595
rect 249 5527 285 5561
rect 249 5493 250 5527
rect 284 5493 285 5527
rect 249 5459 285 5493
rect 249 5425 250 5459
rect 284 5425 285 5459
rect 777 6085 813 6119
rect 777 6051 778 6085
rect 812 6051 813 6085
rect 777 6017 813 6051
rect 777 5983 778 6017
rect 812 5983 813 6017
rect 777 5949 813 5983
rect 777 5915 778 5949
rect 812 5915 813 5949
rect 777 5881 813 5915
rect 777 5847 778 5881
rect 812 5847 813 5881
rect 777 5813 813 5847
rect 777 5779 778 5813
rect 812 5779 813 5813
rect 777 5745 813 5779
rect 777 5711 778 5745
rect 812 5711 813 5745
rect 777 5677 813 5711
rect 777 5643 778 5677
rect 812 5643 813 5677
rect 777 5609 813 5643
rect 777 5575 778 5609
rect 812 5575 813 5609
rect 777 5541 813 5575
rect 777 5507 778 5541
rect 812 5507 813 5541
rect 777 5473 813 5507
rect 249 5391 285 5425
rect 249 5357 250 5391
rect 284 5357 285 5391
rect 777 5439 778 5473
rect 812 5439 813 5473
rect 777 5405 813 5439
rect 249 5323 285 5357
rect 249 5289 250 5323
rect 284 5289 285 5323
rect 249 5255 285 5289
rect 249 5221 250 5255
rect 284 5221 285 5255
rect 249 5187 285 5221
rect 249 5153 250 5187
rect 284 5153 285 5187
rect 249 5119 285 5153
rect 249 5085 250 5119
rect 284 5085 285 5119
rect 777 5371 778 5405
rect 812 5371 813 5405
rect 777 5337 813 5371
rect 777 5303 778 5337
rect 812 5303 813 5337
rect 777 5269 813 5303
rect 777 5235 778 5269
rect 812 5235 813 5269
rect 777 5201 813 5235
rect 777 5167 778 5201
rect 812 5167 813 5201
rect 777 5133 813 5167
rect 777 5099 778 5133
rect 812 5099 813 5133
rect 249 5051 285 5085
rect 249 5017 250 5051
rect 284 5017 285 5051
rect 249 4983 285 5017
rect 249 4949 250 4983
rect 284 4949 285 4983
rect 249 4915 285 4949
rect 777 5065 813 5099
rect 777 5031 778 5065
rect 812 5031 813 5065
rect 777 4997 813 5031
rect 777 4963 778 4997
rect 812 4963 813 4997
rect 777 4929 813 4963
rect 249 4881 250 4915
rect 284 4881 285 4915
rect 249 4847 285 4881
rect 249 4813 250 4847
rect 284 4813 285 4847
rect 249 4779 285 4813
rect 777 4895 778 4929
rect 812 4895 813 4929
rect 777 4861 813 4895
rect 777 4827 778 4861
rect 812 4827 813 4861
rect 777 4793 813 4827
rect 249 4745 250 4779
rect 284 4745 285 4779
rect 249 4711 285 4745
rect 249 4677 250 4711
rect 284 4677 285 4711
rect 249 4643 285 4677
rect 249 4609 250 4643
rect 284 4609 285 4643
rect 777 4759 778 4793
rect 812 4759 813 4793
rect 777 4725 813 4759
rect 777 4691 778 4725
rect 812 4691 813 4725
rect 249 4575 285 4609
rect 249 4541 250 4575
rect 284 4543 285 4575
rect 777 4543 813 4691
rect 284 4542 813 4543
rect 284 4541 337 4542
rect 249 4508 337 4541
rect 371 4508 405 4542
rect 439 4508 473 4542
rect 507 4508 541 4542
rect 575 4508 609 4542
rect 643 4508 677 4542
rect 711 4508 745 4542
rect 779 4508 813 4542
rect 249 4507 813 4508
rect 4645 6221 4681 6265
rect 4645 6187 4646 6221
rect 4680 6187 4681 6221
rect 4645 6153 4681 6187
rect 4645 6119 4646 6153
rect 4680 6119 4681 6153
rect 4645 6085 4681 6119
rect 4645 6051 4646 6085
rect 4680 6051 4681 6085
rect 4645 6017 4681 6051
rect 4645 5983 4646 6017
rect 4680 5983 4681 6017
rect 4645 5949 4681 5983
rect 4645 5915 4646 5949
rect 4680 5915 4681 5949
rect 4645 5881 4681 5915
rect 4645 5847 4646 5881
rect 4680 5847 4681 5881
rect 4645 5813 4681 5847
rect 4645 5779 4646 5813
rect 4680 5779 4681 5813
rect 4645 5745 4681 5779
rect 4645 5711 4646 5745
rect 4680 5711 4681 5745
rect 4645 5677 4681 5711
rect 4645 5643 4646 5677
rect 4680 5643 4681 5677
rect 4645 5609 4681 5643
rect 4645 5575 4646 5609
rect 4680 5575 4681 5609
rect 4645 5541 4681 5575
rect 4645 5507 4646 5541
rect 4680 5507 4681 5541
rect 4645 5473 4681 5507
rect 4645 5439 4646 5473
rect 4680 5439 4681 5473
rect 4645 5405 4681 5439
rect 1668 5163 3114 5164
rect 1668 5129 1702 5163
rect 1736 5129 1770 5163
rect 1804 5129 1838 5163
rect 1872 5129 1906 5163
rect 1940 5129 1974 5163
rect 2008 5129 2042 5163
rect 2076 5129 2110 5163
rect 2144 5129 2178 5163
rect 2212 5129 2246 5163
rect 2280 5129 2314 5163
rect 2348 5129 2382 5163
rect 2416 5129 2450 5163
rect 2484 5129 2518 5163
rect 2552 5129 2586 5163
rect 2620 5129 2654 5163
rect 2688 5129 2722 5163
rect 2756 5129 2790 5163
rect 2824 5129 2858 5163
rect 2892 5129 2926 5163
rect 2960 5129 2994 5163
rect 3028 5130 3114 5163
rect 3028 5129 3079 5130
rect 1668 5128 3079 5129
rect 1668 5094 1704 5128
rect 1668 5060 1669 5094
rect 1703 5060 1704 5094
rect 1668 5026 1704 5060
rect 1668 4992 1669 5026
rect 1703 4992 1704 5026
rect 3078 5096 3079 5128
rect 3113 5096 3114 5130
rect 3078 5062 3114 5096
rect 3078 5028 3079 5062
rect 3113 5028 3114 5062
rect 1668 4958 1704 4992
rect 1668 4924 1669 4958
rect 1703 4924 1704 4958
rect 1668 4890 1704 4924
rect 1668 4856 1669 4890
rect 1703 4856 1704 4890
rect 1668 4822 1704 4856
rect 1668 4788 1669 4822
rect 1703 4788 1704 4822
rect 1668 4754 1704 4788
rect 1668 4720 1669 4754
rect 1703 4720 1704 4754
rect 1668 4686 1704 4720
rect 1668 4652 1669 4686
rect 1703 4652 1704 4686
rect 1668 4618 1704 4652
rect 1668 4584 1669 4618
rect 1703 4584 1704 4618
rect 3078 4994 3114 5028
rect 1668 4550 1704 4584
rect 3078 4960 3079 4994
rect 3113 4960 3114 4994
rect 3078 4926 3114 4960
rect 3078 4892 3079 4926
rect 3113 4892 3114 4926
rect 3078 4858 3114 4892
rect 3078 4824 3079 4858
rect 3113 4824 3114 4858
rect 3078 4790 3114 4824
rect 3078 4756 3079 4790
rect 3113 4756 3114 4790
rect 3078 4722 3114 4756
rect 3078 4688 3079 4722
rect 3113 4688 3114 4722
rect 3078 4654 3114 4688
rect 3078 4620 3079 4654
rect 3113 4620 3114 4654
rect 3078 4586 3114 4620
rect 1668 4516 1669 4550
rect 1703 4516 1704 4550
rect 3078 4552 3079 4586
rect 3113 4552 3114 4586
rect 1668 4482 1704 4516
rect 1668 4448 1669 4482
rect 1703 4448 1704 4482
rect 1668 4414 1704 4448
rect 1668 4380 1669 4414
rect 1703 4380 1704 4414
rect 1668 4346 1704 4380
rect 1668 4312 1669 4346
rect 1703 4312 1704 4346
rect 1668 4278 1704 4312
rect 1668 4244 1669 4278
rect 1703 4244 1704 4278
rect 1668 4210 1704 4244
rect 1668 4176 1669 4210
rect 1703 4176 1704 4210
rect 1668 4142 1704 4176
rect 3078 4518 3114 4552
rect 3078 4484 3079 4518
rect 3113 4484 3114 4518
rect 3078 4450 3114 4484
rect 3078 4416 3079 4450
rect 3113 4416 3114 4450
rect 3078 4382 3114 4416
rect 3078 4348 3079 4382
rect 3113 4348 3114 4382
rect 3078 4314 3114 4348
rect 3078 4280 3079 4314
rect 3113 4280 3114 4314
rect 3078 4246 3114 4280
rect 3078 4212 3079 4246
rect 3113 4212 3114 4246
rect 1668 4108 1669 4142
rect 1703 4108 1704 4142
rect 1668 4074 1704 4108
rect 3078 4178 3114 4212
rect 3078 4144 3079 4178
rect 3113 4144 3114 4178
rect 3078 4110 3114 4144
rect 1668 4040 1669 4074
rect 1703 4040 1704 4074
rect 1668 4006 1704 4040
rect 1668 3972 1669 4006
rect 1703 3972 1704 4006
rect 1668 3938 1704 3972
rect 1668 3904 1669 3938
rect 1703 3904 1704 3938
rect 1668 3870 1704 3904
rect 1668 3836 1669 3870
rect 1703 3836 1704 3870
rect 1668 3802 1704 3836
rect 1668 3768 1669 3802
rect 1703 3768 1704 3802
rect 1668 3734 1704 3768
rect 1668 3700 1669 3734
rect 1703 3700 1704 3734
rect 1668 3666 1704 3700
rect 3078 4076 3079 4110
rect 3113 4076 3114 4110
rect 3078 4042 3114 4076
rect 3078 4008 3079 4042
rect 3113 4008 3114 4042
rect 3078 3974 3114 4008
rect 3078 3940 3079 3974
rect 3113 3940 3114 3974
rect 3078 3906 3114 3940
rect 3078 3872 3079 3906
rect 3113 3872 3114 3906
rect 3078 3838 3114 3872
rect 3078 3804 3079 3838
rect 3113 3804 3114 3838
rect 3078 3770 3114 3804
rect 3078 3736 3079 3770
rect 3113 3736 3114 3770
rect 1668 3632 1669 3666
rect 1703 3632 1704 3666
rect 3078 3702 3114 3736
rect 3078 3668 3079 3702
rect 3113 3668 3114 3702
rect 1668 3598 1704 3632
rect 1668 3564 1669 3598
rect 1703 3564 1704 3598
rect 1668 3530 1704 3564
rect 1668 3496 1669 3530
rect 1703 3496 1704 3530
rect 1668 3462 1704 3496
rect 1668 3428 1669 3462
rect 1703 3428 1704 3462
rect 1668 3394 1704 3428
rect 1668 3360 1669 3394
rect 1703 3360 1704 3394
rect 1668 3326 1704 3360
rect 1668 3292 1669 3326
rect 1703 3292 1704 3326
rect 1668 3258 1704 3292
rect 1668 3224 1669 3258
rect 1703 3224 1704 3258
rect 3078 3634 3114 3668
rect 3078 3600 3079 3634
rect 3113 3600 3114 3634
rect 3078 3566 3114 3600
rect 3078 3532 3079 3566
rect 3113 3532 3114 3566
rect 3078 3498 3114 3532
rect 3078 3464 3079 3498
rect 3113 3464 3114 3498
rect 3078 3430 3114 3464
rect 3078 3396 3079 3430
rect 3113 3396 3114 3430
rect 3078 3362 3114 3396
rect 3078 3328 3079 3362
rect 3113 3328 3114 3362
rect 3078 3294 3114 3328
rect 1668 3190 1704 3224
rect 1668 3156 1669 3190
rect 1703 3156 1704 3190
rect 1668 3122 1704 3156
rect 1668 3088 1669 3122
rect 1703 3088 1704 3122
rect 1668 3054 1704 3088
rect 1668 3020 1669 3054
rect 1703 3020 1704 3054
rect 1668 2986 1704 3020
rect 1668 2952 1669 2986
rect 1703 2952 1704 2986
rect 1668 2918 1704 2952
rect 1668 2884 1669 2918
rect 1703 2884 1704 2918
rect 1668 2850 1704 2884
rect 1668 2816 1669 2850
rect 1703 2816 1704 2850
rect 1668 2782 1704 2816
rect 1668 2748 1669 2782
rect 1703 2748 1704 2782
rect 3078 3260 3079 3294
rect 3113 3260 3114 3294
rect 3078 3226 3114 3260
rect 3078 3192 3079 3226
rect 3113 3192 3114 3226
rect 3078 3158 3114 3192
rect 3078 3124 3079 3158
rect 3113 3124 3114 3158
rect 3078 3090 3114 3124
rect 3078 3056 3079 3090
rect 3113 3056 3114 3090
rect 3078 3022 3114 3056
rect 3078 2988 3079 3022
rect 3113 2988 3114 3022
rect 1668 2714 1704 2748
rect 1668 2680 1669 2714
rect 1703 2680 1704 2714
rect 1668 2646 1704 2680
rect 1668 2612 1669 2646
rect 1703 2612 1704 2646
rect 1668 2578 1704 2612
rect 1668 2544 1669 2578
rect 1703 2544 1704 2578
rect 1668 2510 1704 2544
rect 1668 2476 1669 2510
rect 1703 2476 1704 2510
rect 1668 2442 1704 2476
rect 1668 2408 1669 2442
rect 1703 2408 1704 2442
rect 1668 2374 1704 2408
rect 1668 2340 1669 2374
rect 1703 2340 1704 2374
rect 1668 2306 1704 2340
rect 3078 2954 3114 2988
rect 3078 2920 3079 2954
rect 3113 2920 3114 2954
rect 3078 2886 3114 2920
rect 3078 2852 3079 2886
rect 3113 2852 3114 2886
rect 3078 2818 3114 2852
rect 3078 2784 3079 2818
rect 3113 2784 3114 2818
rect 3078 2750 3114 2784
rect 3078 2716 3079 2750
rect 3113 2716 3114 2750
rect 3078 2682 3114 2716
rect 3078 2648 3079 2682
rect 3113 2648 3114 2682
rect 3078 2614 3114 2648
rect 3078 2580 3079 2614
rect 3113 2580 3114 2614
rect 3078 2546 3114 2580
rect 3078 2512 3079 2546
rect 3113 2512 3114 2546
rect 3078 2478 3114 2512
rect 3078 2444 3079 2478
rect 3113 2444 3114 2478
rect 3078 2410 3114 2444
rect 3078 2376 3079 2410
rect 3113 2376 3114 2410
rect 3078 2342 3114 2376
rect 1668 2272 1669 2306
rect 1703 2272 1704 2306
rect 1668 2238 1704 2272
rect 1668 2204 1669 2238
rect 1703 2204 1704 2238
rect 1668 2170 1704 2204
rect 1668 2136 1669 2170
rect 1703 2136 1704 2170
rect 1668 2102 1704 2136
rect 1668 2068 1669 2102
rect 1703 2068 1704 2102
rect 1668 2034 1704 2068
rect 1668 2000 1669 2034
rect 1703 2000 1704 2034
rect 1668 1966 1704 2000
rect 1668 1932 1669 1966
rect 1703 1932 1704 1966
rect 1668 1898 1704 1932
rect 1668 1864 1669 1898
rect 1703 1864 1704 1898
rect 3078 2308 3079 2342
rect 3113 2308 3114 2342
rect 3078 2274 3114 2308
rect 3078 2240 3079 2274
rect 3113 2240 3114 2274
rect 3078 2206 3114 2240
rect 3078 2172 3079 2206
rect 3113 2172 3114 2206
rect 3078 2138 3114 2172
rect 3078 2104 3079 2138
rect 3113 2104 3114 2138
rect 3078 2070 3114 2104
rect 3078 2036 3079 2070
rect 3113 2036 3114 2070
rect 3078 2002 3114 2036
rect 3078 1968 3079 2002
rect 3113 1968 3114 2002
rect 3078 1934 3114 1968
rect 1668 1830 1704 1864
rect 1668 1796 1669 1830
rect 1703 1796 1704 1830
rect 3078 1900 3079 1934
rect 3113 1900 3114 1934
rect 3078 1866 3114 1900
rect 1668 1762 1704 1796
rect 1668 1728 1669 1762
rect 1703 1728 1704 1762
rect 1668 1694 1704 1728
rect 1668 1660 1669 1694
rect 1703 1660 1704 1694
rect 1668 1626 1704 1660
rect 1668 1592 1669 1626
rect 1703 1592 1704 1626
rect 1668 1558 1704 1592
rect 1668 1524 1669 1558
rect 1703 1524 1704 1558
rect 1668 1490 1704 1524
rect 1668 1456 1669 1490
rect 1703 1456 1704 1490
rect 1668 1422 1704 1456
rect 1668 1388 1669 1422
rect 1703 1388 1704 1422
rect 3078 1832 3079 1866
rect 3113 1832 3114 1866
rect 3078 1798 3114 1832
rect 3078 1764 3079 1798
rect 3113 1764 3114 1798
rect 3078 1730 3114 1764
rect 3078 1696 3079 1730
rect 3113 1696 3114 1730
rect 3078 1662 3114 1696
rect 3078 1628 3079 1662
rect 3113 1628 3114 1662
rect 3078 1594 3114 1628
rect 3078 1560 3079 1594
rect 3113 1560 3114 1594
rect 3078 1526 3114 1560
rect 3078 1492 3079 1526
rect 3113 1492 3114 1526
rect 3078 1458 3114 1492
rect 1668 1354 1704 1388
rect 1668 1320 1669 1354
rect 1703 1320 1704 1354
rect 3078 1424 3079 1458
rect 3113 1424 3114 1458
rect 1668 1286 1704 1320
rect 1668 1252 1669 1286
rect 1703 1252 1704 1286
rect 1668 1218 1704 1252
rect 1668 1184 1669 1218
rect 1703 1184 1704 1218
rect 1668 1150 1704 1184
rect 1668 1116 1669 1150
rect 1703 1116 1704 1150
rect 1668 1082 1704 1116
rect 1668 1048 1669 1082
rect 1703 1048 1704 1082
rect 1668 1014 1704 1048
rect 1668 980 1669 1014
rect 1703 980 1704 1014
rect 1668 946 1704 980
rect 3078 1390 3114 1424
rect 3078 1356 3079 1390
rect 3113 1356 3114 1390
rect 3078 1322 3114 1356
rect 3078 1288 3079 1322
rect 3113 1288 3114 1322
rect 3078 1254 3114 1288
rect 3078 1220 3079 1254
rect 3113 1220 3114 1254
rect 3078 1186 3114 1220
rect 3078 1152 3079 1186
rect 3113 1152 3114 1186
rect 3078 1118 3114 1152
rect 3078 1084 3079 1118
rect 3113 1084 3114 1118
rect 3078 1050 3114 1084
rect 3078 1016 3079 1050
rect 3113 1016 3114 1050
rect 3078 982 3114 1016
rect 1668 912 1669 946
rect 1703 912 1704 946
rect 3078 948 3079 982
rect 3113 948 3114 982
rect 1668 878 1704 912
rect 1668 844 1669 878
rect 1703 844 1704 878
rect 1668 810 1704 844
rect 1668 776 1669 810
rect 1703 776 1704 810
rect 1668 742 1704 776
rect 1668 708 1669 742
rect 1703 708 1704 742
rect 1668 674 1704 708
rect 1668 640 1669 674
rect 1703 640 1704 674
rect 1668 606 1704 640
rect 1668 572 1669 606
rect 1703 572 1704 606
rect 1668 538 1704 572
rect 1668 504 1669 538
rect 1703 504 1704 538
rect 1668 470 1704 504
rect 3078 914 3114 948
rect 3078 880 3079 914
rect 3113 880 3114 914
rect 3078 846 3114 880
rect 3078 812 3079 846
rect 3113 812 3114 846
rect 3078 778 3114 812
rect 3078 744 3079 778
rect 3113 744 3114 778
rect 3078 710 3114 744
rect 3078 676 3079 710
rect 3113 676 3114 710
rect 3078 642 3114 676
rect 3078 608 3079 642
rect 3113 608 3114 642
rect 3078 574 3114 608
rect 3078 540 3079 574
rect 3113 540 3114 574
rect 3078 506 3114 540
rect 1668 436 1669 470
rect 1703 436 1704 470
rect 1668 402 1704 436
rect 1668 368 1669 402
rect 1703 370 1704 402
rect 3078 472 3079 506
rect 3113 472 3114 506
rect 3078 370 3114 472
rect 1703 369 3114 370
rect 1703 368 1754 369
rect 1668 335 1754 368
rect 1788 335 1822 369
rect 1856 335 1890 369
rect 1924 335 1958 369
rect 1992 335 2026 369
rect 2060 335 2094 369
rect 2128 335 2162 369
rect 2196 335 2230 369
rect 2264 335 2298 369
rect 2332 335 2366 369
rect 2400 335 2434 369
rect 2468 335 2502 369
rect 2536 335 2570 369
rect 2604 335 2638 369
rect 2672 335 2706 369
rect 2740 335 2774 369
rect 2808 335 2842 369
rect 2876 335 2910 369
rect 2944 335 2978 369
rect 3012 335 3046 369
rect 3080 335 3114 369
rect 4645 5371 4646 5405
rect 4680 5371 4681 5405
rect 4645 5337 4681 5371
rect 4645 5303 4646 5337
rect 4680 5303 4681 5337
rect 4645 5269 4681 5303
rect 4645 5235 4646 5269
rect 4680 5235 4681 5269
rect 4645 5201 4681 5235
rect 4645 5167 4646 5201
rect 4680 5167 4681 5201
rect 4645 5133 4681 5167
rect 4645 5099 4646 5133
rect 4680 5099 4681 5133
rect 13646 6232 13682 6266
rect 13646 6198 13647 6232
rect 13681 6198 13682 6232
rect 13646 6164 13682 6198
rect 13646 6130 13647 6164
rect 13681 6130 13682 6164
rect 13646 6096 13682 6130
rect 13646 6062 13647 6096
rect 13681 6062 13682 6096
rect 13646 6028 13682 6062
rect 13646 5994 13647 6028
rect 13681 5994 13682 6028
rect 13646 5960 13682 5994
rect 13646 5926 13647 5960
rect 13681 5926 13682 5960
rect 13646 5892 13682 5926
rect 13646 5858 13647 5892
rect 13681 5858 13682 5892
rect 13646 5824 13682 5858
rect 13646 5790 13647 5824
rect 13681 5790 13682 5824
rect 13646 5756 13682 5790
rect 13646 5722 13647 5756
rect 13681 5722 13682 5756
rect 13646 5688 13682 5722
rect 13646 5654 13647 5688
rect 13681 5654 13682 5688
rect 13646 5620 13682 5654
rect 13646 5586 13647 5620
rect 13681 5586 13682 5620
rect 13646 5552 13682 5586
rect 13646 5518 13647 5552
rect 13681 5518 13682 5552
rect 13646 5484 13682 5518
rect 13646 5450 13647 5484
rect 13681 5450 13682 5484
rect 13646 5416 13682 5450
rect 13646 5382 13647 5416
rect 13681 5382 13682 5416
rect 13646 5348 13682 5382
rect 13646 5314 13647 5348
rect 13681 5314 13682 5348
rect 13646 5280 13682 5314
rect 13646 5246 13647 5280
rect 13681 5246 13682 5280
rect 13646 5212 13682 5246
rect 13646 5178 13647 5212
rect 13681 5178 13682 5212
rect 4645 5065 4681 5099
rect 4645 5031 4646 5065
rect 4680 5031 4681 5065
rect 4645 4997 4681 5031
rect 4645 4963 4646 4997
rect 4680 4963 4681 4997
rect 4645 4929 4681 4963
rect 4645 4895 4646 4929
rect 4680 4895 4681 4929
rect 4645 4861 4681 4895
rect 4645 4827 4646 4861
rect 4680 4827 4681 4861
rect 4645 4793 4681 4827
rect 4645 4759 4646 4793
rect 4680 4759 4681 4793
rect 4645 4725 4681 4759
rect 4645 4691 4646 4725
rect 4680 4691 4681 4725
rect 4645 4657 4681 4691
rect 4645 4623 4646 4657
rect 4680 4623 4681 4657
rect 4645 4589 4681 4623
rect 4645 4555 4646 4589
rect 4680 4555 4681 4589
rect 4645 4521 4681 4555
rect 4645 4487 4646 4521
rect 4680 4487 4681 4521
rect 4645 4453 4681 4487
rect 4645 4419 4646 4453
rect 4680 4419 4681 4453
rect 4645 4385 4681 4419
rect 4645 4351 4646 4385
rect 4680 4351 4681 4385
rect 4645 4317 4681 4351
rect 4645 4283 4646 4317
rect 4680 4283 4681 4317
rect 4645 4249 4681 4283
rect 4645 4215 4646 4249
rect 4680 4215 4681 4249
rect 4645 4181 4681 4215
rect 4645 4147 4646 4181
rect 4680 4147 4681 4181
rect 4645 4113 4681 4147
rect 4645 4079 4646 4113
rect 4680 4079 4681 4113
rect 4645 4045 4681 4079
rect 4645 4011 4646 4045
rect 4680 4011 4681 4045
rect 4645 3977 4681 4011
rect 4645 3943 4646 3977
rect 4680 3943 4681 3977
rect 4645 3909 4681 3943
rect 4645 3875 4646 3909
rect 4680 3875 4681 3909
rect 4645 3841 4681 3875
rect 4645 3807 4646 3841
rect 4680 3807 4681 3841
rect 4645 3773 4681 3807
rect 4645 3739 4646 3773
rect 4680 3739 4681 3773
rect 4645 3705 4681 3739
rect 4645 3671 4646 3705
rect 4680 3671 4681 3705
rect 4645 3637 4681 3671
rect 4645 3603 4646 3637
rect 4680 3603 4681 3637
rect 4645 3569 4681 3603
rect 4645 3535 4646 3569
rect 4680 3535 4681 3569
rect 4645 3501 4681 3535
rect 4645 3467 4646 3501
rect 4680 3467 4681 3501
rect 4645 3433 4681 3467
rect 4645 3399 4646 3433
rect 4680 3399 4681 3433
rect 4645 3365 4681 3399
rect 4645 3331 4646 3365
rect 4680 3331 4681 3365
rect 4645 3297 4681 3331
rect 4645 3263 4646 3297
rect 4680 3263 4681 3297
rect 4645 3229 4681 3263
rect 4645 3195 4646 3229
rect 4680 3195 4681 3229
rect 4645 3161 4681 3195
rect 4645 3127 4646 3161
rect 4680 3127 4681 3161
rect 4645 3093 4681 3127
rect 4645 3059 4646 3093
rect 4680 3059 4681 3093
rect 4645 3025 4681 3059
rect 4645 2991 4646 3025
rect 4680 2991 4681 3025
rect 4645 2957 4681 2991
rect 4645 2923 4646 2957
rect 4680 2923 4681 2957
rect 4645 2889 4681 2923
rect 4645 2855 4646 2889
rect 4680 2855 4681 2889
rect 4645 2821 4681 2855
rect 4645 2787 4646 2821
rect 4680 2787 4681 2821
rect 4645 2753 4681 2787
rect 4645 2719 4646 2753
rect 4680 2719 4681 2753
rect 4645 2685 4681 2719
rect 4645 2651 4646 2685
rect 4680 2651 4681 2685
rect 4645 2617 4681 2651
rect 4645 2583 4646 2617
rect 4680 2583 4681 2617
rect 4645 2549 4681 2583
rect 4645 2515 4646 2549
rect 4680 2515 4681 2549
rect 4645 2481 4681 2515
rect 4645 2447 4646 2481
rect 4680 2447 4681 2481
rect 4645 2413 4681 2447
rect 4645 2379 4646 2413
rect 4680 2379 4681 2413
rect 4645 2345 4681 2379
rect 4645 2311 4646 2345
rect 4680 2311 4681 2345
rect 4645 2277 4681 2311
rect 4645 2243 4646 2277
rect 4680 2243 4681 2277
rect 4645 2209 4681 2243
rect 4645 2175 4646 2209
rect 4680 2175 4681 2209
rect 4645 2141 4681 2175
rect 4645 2107 4646 2141
rect 4680 2107 4681 2141
rect 4645 2073 4681 2107
rect 4645 2039 4646 2073
rect 4680 2039 4681 2073
rect 4645 2005 4681 2039
rect 4645 1971 4646 2005
rect 4680 1971 4681 2005
rect 4645 1937 4681 1971
rect 4645 1903 4646 1937
rect 4680 1903 4681 1937
rect 4645 1869 4681 1903
rect 4645 1835 4646 1869
rect 4680 1835 4681 1869
rect 4645 1801 4681 1835
rect 4645 1767 4646 1801
rect 4680 1767 4681 1801
rect 4645 1733 4681 1767
rect 4645 1699 4646 1733
rect 4680 1699 4681 1733
rect 4645 1665 4681 1699
rect 4645 1631 4646 1665
rect 4680 1631 4681 1665
rect 4645 1597 4681 1631
rect 4645 1563 4646 1597
rect 4680 1563 4681 1597
rect 4645 1529 4681 1563
rect 4645 1495 4646 1529
rect 4680 1495 4681 1529
rect 4645 1461 4681 1495
rect 4645 1427 4646 1461
rect 4680 1427 4681 1461
rect 4645 1393 4681 1427
rect 4645 1359 4646 1393
rect 4680 1359 4681 1393
rect 4645 1325 4681 1359
rect 4645 1291 4646 1325
rect 4680 1291 4681 1325
rect 4645 1257 4681 1291
rect 4645 1223 4646 1257
rect 4680 1223 4681 1257
rect 4645 1189 4681 1223
rect 4645 1155 4646 1189
rect 4680 1155 4681 1189
rect 4645 1121 4681 1155
rect 4645 1087 4646 1121
rect 4680 1087 4681 1121
rect 4645 1053 4681 1087
rect 4645 1019 4646 1053
rect 4680 1019 4681 1053
rect 4645 985 4681 1019
rect 4645 951 4646 985
rect 4680 951 4681 985
rect 4645 917 4681 951
rect 4645 883 4646 917
rect 4680 883 4681 917
rect 4645 849 4681 883
rect 4645 815 4646 849
rect 4680 815 4681 849
rect 4645 781 4681 815
rect 4645 747 4646 781
rect 4680 747 4681 781
rect 4645 713 4681 747
rect 4645 679 4646 713
rect 4680 679 4681 713
rect 4645 645 4681 679
rect 4645 611 4646 645
rect 4680 611 4681 645
rect 4645 577 4681 611
rect 4645 543 4646 577
rect 4680 543 4681 577
rect 4645 509 4681 543
rect 4645 475 4646 509
rect 4680 475 4681 509
rect 4645 441 4681 475
rect 4645 407 4646 441
rect 4680 407 4681 441
rect 4645 373 4681 407
rect 1668 334 3114 335
rect 4645 339 4646 373
rect 4680 339 4681 373
rect 4645 305 4681 339
rect 4645 271 4646 305
rect 4680 271 4681 305
rect 4645 237 4681 271
rect 4645 203 4646 237
rect 4680 203 4681 237
rect 13646 5080 13682 5178
rect 12945 5079 13682 5080
rect 12945 5046 13070 5079
rect 12945 5012 12946 5046
rect 12980 5045 13070 5046
rect 13104 5045 13138 5079
rect 13172 5045 13206 5079
rect 13240 5045 13274 5079
rect 13308 5045 13342 5079
rect 13376 5045 13410 5079
rect 13444 5045 13478 5079
rect 13512 5045 13546 5079
rect 13580 5045 13614 5079
rect 13648 5045 13682 5079
rect 12980 5044 13682 5045
rect 12980 5012 12981 5044
rect 12945 4978 12981 5012
rect 12945 4944 12946 4978
rect 12980 4944 12981 4978
rect 12945 4910 12981 4944
rect 12945 4876 12946 4910
rect 12980 4876 12981 4910
rect 12945 4842 12981 4876
rect 12945 4808 12946 4842
rect 12980 4808 12981 4842
rect 12945 4774 12981 4808
rect 12945 4740 12946 4774
rect 12980 4740 12981 4774
rect 12945 4706 12981 4740
rect 12945 4672 12946 4706
rect 12980 4672 12981 4706
rect 12945 4638 12981 4672
rect 12945 4604 12946 4638
rect 12980 4604 12981 4638
rect 12945 4570 12981 4604
rect 12945 4536 12946 4570
rect 12980 4536 12981 4570
rect 12945 4502 12981 4536
rect 12945 4468 12946 4502
rect 12980 4468 12981 4502
rect 12945 4434 12981 4468
rect 12945 4400 12946 4434
rect 12980 4400 12981 4434
rect 12945 4366 12981 4400
rect 12945 4332 12946 4366
rect 12980 4332 12981 4366
rect 12945 4298 12981 4332
rect 12945 4264 12946 4298
rect 12980 4264 12981 4298
rect 12945 4230 12981 4264
rect 12945 4196 12946 4230
rect 12980 4196 12981 4230
rect 12945 4162 12981 4196
rect 12945 4128 12946 4162
rect 12980 4128 12981 4162
rect 12945 4094 12981 4128
rect 12945 4060 12946 4094
rect 12980 4060 12981 4094
rect 12945 4026 12981 4060
rect 12945 3992 12946 4026
rect 12980 3992 12981 4026
rect 12945 3958 12981 3992
rect 12945 3924 12946 3958
rect 12980 3924 12981 3958
rect 12945 3890 12981 3924
rect 12945 3856 12946 3890
rect 12980 3856 12981 3890
rect 12945 3822 12981 3856
rect 12945 3788 12946 3822
rect 12980 3788 12981 3822
rect 12945 3754 12981 3788
rect 12945 3720 12946 3754
rect 12980 3720 12981 3754
rect 12945 3686 12981 3720
rect 12945 3652 12946 3686
rect 12980 3652 12981 3686
rect 12945 3618 12981 3652
rect 12945 3584 12946 3618
rect 12980 3584 12981 3618
rect 12945 3550 12981 3584
rect 12945 3516 12946 3550
rect 12980 3516 12981 3550
rect 12945 3482 12981 3516
rect 12945 3448 12946 3482
rect 12980 3448 12981 3482
rect 12945 3414 12981 3448
rect 12945 3380 12946 3414
rect 12980 3380 12981 3414
rect 12945 3346 12981 3380
rect 12945 3312 12946 3346
rect 12980 3312 12981 3346
rect 12945 3278 12981 3312
rect 12945 3244 12946 3278
rect 12980 3244 12981 3278
rect 12945 3210 12981 3244
rect 12945 3176 12946 3210
rect 12980 3176 12981 3210
rect 12945 3142 12981 3176
rect 12945 3108 12946 3142
rect 12980 3108 12981 3142
rect 12945 3074 12981 3108
rect 12945 3040 12946 3074
rect 12980 3040 12981 3074
rect 12945 3006 12981 3040
rect 12945 2972 12946 3006
rect 12980 2972 12981 3006
rect 12945 2938 12981 2972
rect 12945 2904 12946 2938
rect 12980 2904 12981 2938
rect 12945 2870 12981 2904
rect 12945 2836 12946 2870
rect 12980 2836 12981 2870
rect 12945 2802 12981 2836
rect 12945 2768 12946 2802
rect 12980 2768 12981 2802
rect 12945 2734 12981 2768
rect 12945 2700 12946 2734
rect 12980 2700 12981 2734
rect 12945 2666 12981 2700
rect 12945 2632 12946 2666
rect 12980 2632 12981 2666
rect 12945 2598 12981 2632
rect 12945 2564 12946 2598
rect 12980 2564 12981 2598
rect 12945 2530 12981 2564
rect 12945 2496 12946 2530
rect 12980 2496 12981 2530
rect 12945 2462 12981 2496
rect 12945 2428 12946 2462
rect 12980 2428 12981 2462
rect 12945 2394 12981 2428
rect 12945 2360 12946 2394
rect 12980 2360 12981 2394
rect 12945 2326 12981 2360
rect 12945 2292 12946 2326
rect 12980 2292 12981 2326
rect 12945 2258 12981 2292
rect 12945 2224 12946 2258
rect 12980 2224 12981 2258
rect 12945 2190 12981 2224
rect 12945 2156 12946 2190
rect 12980 2156 12981 2190
rect 12945 2122 12981 2156
rect 12945 2088 12946 2122
rect 12980 2088 12981 2122
rect 12945 2054 12981 2088
rect 12945 2020 12946 2054
rect 12980 2020 12981 2054
rect 12945 1986 12981 2020
rect 12945 1952 12946 1986
rect 12980 1952 12981 1986
rect 12945 1918 12981 1952
rect 12945 1884 12946 1918
rect 12980 1884 12981 1918
rect 12945 1850 12981 1884
rect 12945 1816 12946 1850
rect 12980 1816 12981 1850
rect 12945 1782 12981 1816
rect 12945 1748 12946 1782
rect 12980 1748 12981 1782
rect 12945 1714 12981 1748
rect 12945 1680 12946 1714
rect 12980 1680 12981 1714
rect 12945 1646 12981 1680
rect 12945 1612 12946 1646
rect 12980 1612 12981 1646
rect 12945 1578 12981 1612
rect 12945 1544 12946 1578
rect 12980 1544 12981 1578
rect 12945 1510 12981 1544
rect 12945 1476 12946 1510
rect 12980 1476 12981 1510
rect 12945 1442 12981 1476
rect 12945 1408 12946 1442
rect 12980 1408 12981 1442
rect 12945 1374 12981 1408
rect 12945 1340 12946 1374
rect 12980 1340 12981 1374
rect 12945 1306 12981 1340
rect 12945 1272 12946 1306
rect 12980 1272 12981 1306
rect 12945 1238 12981 1272
rect 12945 1204 12946 1238
rect 12980 1204 12981 1238
rect 12945 1170 12981 1204
rect 12945 1136 12946 1170
rect 12980 1136 12981 1170
rect 12945 1102 12981 1136
rect 12945 1068 12946 1102
rect 12980 1068 12981 1102
rect 12945 1034 12981 1068
rect 12945 1000 12946 1034
rect 12980 1000 12981 1034
rect 12945 966 12981 1000
rect 12945 932 12946 966
rect 12980 932 12981 966
rect 12945 898 12981 932
rect 12945 864 12946 898
rect 12980 864 12981 898
rect 12945 830 12981 864
rect 12945 796 12946 830
rect 12980 796 12981 830
rect 12945 762 12981 796
rect 12945 728 12946 762
rect 12980 728 12981 762
rect 12945 694 12981 728
rect 12945 660 12946 694
rect 12980 660 12981 694
rect 12945 626 12981 660
rect 12945 592 12946 626
rect 12980 592 12981 626
rect 12945 558 12981 592
rect 12945 524 12946 558
rect 12980 524 12981 558
rect 12945 490 12981 524
rect 12945 456 12946 490
rect 12980 456 12981 490
rect 12945 422 12981 456
rect 12945 388 12946 422
rect 12980 388 12981 422
rect 12945 354 12981 388
rect 4645 169 4681 203
rect 12945 320 12946 354
rect 12980 320 12981 354
rect 12945 286 12981 320
rect 12945 252 12946 286
rect 12980 252 12981 286
rect 12945 218 12981 252
rect 4645 135 4646 169
rect 4680 135 4681 169
rect 4645 101 4681 135
rect 4645 67 4646 101
rect 4680 67 4681 101
rect 4645 33 4681 67
rect 4645 -1 4646 33
rect 4680 -1 4681 33
rect 4645 -35 4681 -1
rect 12945 184 12946 218
rect 12980 184 12981 218
rect 12945 150 12981 184
rect 12945 116 12946 150
rect 12980 116 12981 150
rect 12945 82 12981 116
rect 12945 48 12946 82
rect 12980 48 12981 82
rect 12945 14 12981 48
rect 4645 -69 4646 -35
rect 4680 -69 4681 -35
rect 4645 -103 4681 -69
rect 4645 -137 4646 -103
rect 4680 -137 4681 -103
rect 4645 -171 4681 -137
rect 12945 -20 12946 14
rect 12980 -20 12981 14
rect 12945 -54 12981 -20
rect 12945 -88 12946 -54
rect 12980 -88 12981 -54
rect 4645 -205 4646 -171
rect 4680 -205 4681 -171
rect 4645 -239 4681 -205
rect 4645 -273 4646 -239
rect 4680 -273 4681 -239
rect 4645 -307 4681 -273
rect 4645 -341 4646 -307
rect 4680 -341 4681 -307
rect 4645 -375 4681 -341
rect 4645 -409 4646 -375
rect 4680 -407 4681 -375
rect 12945 -223 12981 -88
rect 12945 -257 12946 -223
rect 12980 -257 12981 -223
rect 12945 -291 12981 -257
rect 12945 -325 12946 -291
rect 12980 -325 12981 -291
rect 12945 -407 12981 -325
rect 4680 -408 12981 -407
rect 4680 -409 4753 -408
rect 4645 -442 4753 -409
rect 4787 -442 4821 -408
rect 4855 -442 4889 -408
rect 4923 -442 4957 -408
rect 4991 -442 5025 -408
rect 5059 -442 5093 -408
rect 5127 -442 5161 -408
rect 5195 -442 5229 -408
rect 5263 -442 5297 -408
rect 5331 -442 5365 -408
rect 5399 -442 5433 -408
rect 5467 -442 5501 -408
rect 5535 -442 5569 -408
rect 5603 -442 5637 -408
rect 5671 -442 5705 -408
rect 5739 -442 5773 -408
rect 5807 -442 5841 -408
rect 5875 -442 5909 -408
rect 5943 -442 5977 -408
rect 6011 -442 6045 -408
rect 6079 -442 6113 -408
rect 6147 -442 6181 -408
rect 6215 -442 6249 -408
rect 6283 -442 6317 -408
rect 6351 -442 6385 -408
rect 6419 -442 6453 -408
rect 6487 -442 6521 -408
rect 6555 -442 6589 -408
rect 6623 -442 6657 -408
rect 6691 -442 6725 -408
rect 6759 -442 6793 -408
rect 6827 -442 6861 -408
rect 6895 -442 6929 -408
rect 6963 -442 6997 -408
rect 7031 -442 7065 -408
rect 7099 -442 7133 -408
rect 7167 -442 7201 -408
rect 7235 -442 7269 -408
rect 7303 -442 7337 -408
rect 7371 -442 7405 -408
rect 7439 -442 7473 -408
rect 7507 -442 7541 -408
rect 7575 -442 7609 -408
rect 7643 -442 7677 -408
rect 7711 -442 7745 -408
rect 7779 -442 7813 -408
rect 7847 -442 7881 -408
rect 7915 -442 7949 -408
rect 7983 -442 8017 -408
rect 8051 -442 8085 -408
rect 8119 -442 8153 -408
rect 8187 -442 8221 -408
rect 8255 -442 8289 -408
rect 8323 -442 8357 -408
rect 8391 -442 8425 -408
rect 8459 -442 8493 -408
rect 8527 -442 8561 -408
rect 8595 -442 8629 -408
rect 8663 -442 8697 -408
rect 8731 -442 8765 -408
rect 8799 -442 8833 -408
rect 8867 -442 8901 -408
rect 8935 -442 8969 -408
rect 9003 -442 9037 -408
rect 9071 -442 9105 -408
rect 9139 -442 9173 -408
rect 9207 -442 9241 -408
rect 9275 -442 9309 -408
rect 9343 -442 9377 -408
rect 9411 -442 9445 -408
rect 9479 -442 9513 -408
rect 9547 -442 9581 -408
rect 9615 -442 9649 -408
rect 9683 -442 9717 -408
rect 9751 -442 9785 -408
rect 9819 -442 9853 -408
rect 9887 -442 9921 -408
rect 9955 -442 9989 -408
rect 10023 -442 10057 -408
rect 10091 -442 10125 -408
rect 10159 -442 10193 -408
rect 10227 -442 10261 -408
rect 10295 -442 10329 -408
rect 10363 -442 10397 -408
rect 10431 -442 10465 -408
rect 10499 -442 10533 -408
rect 10567 -442 10601 -408
rect 10635 -442 10669 -408
rect 10703 -442 10737 -408
rect 10771 -442 10805 -408
rect 10839 -442 10873 -408
rect 10907 -442 10941 -408
rect 10975 -442 11009 -408
rect 11043 -442 11077 -408
rect 11111 -442 11145 -408
rect 11179 -442 11213 -408
rect 11247 -442 11281 -408
rect 11315 -442 11349 -408
rect 11383 -442 11417 -408
rect 11451 -442 11485 -408
rect 11519 -442 11553 -408
rect 11587 -442 11621 -408
rect 11655 -442 11689 -408
rect 11723 -442 11757 -408
rect 11791 -442 11825 -408
rect 11859 -442 11893 -408
rect 11927 -442 11961 -408
rect 11995 -442 12029 -408
rect 12063 -442 12097 -408
rect 12131 -442 12165 -408
rect 12199 -442 12233 -408
rect 12267 -442 12301 -408
rect 12335 -442 12369 -408
rect 12403 -442 12437 -408
rect 12471 -442 12505 -408
rect 12539 -442 12573 -408
rect 12607 -442 12641 -408
rect 12675 -442 12709 -408
rect 12743 -442 12777 -408
rect 12811 -442 12845 -408
rect 12879 -442 12913 -408
rect 12947 -442 12981 -408
rect 4645 -443 12981 -442
<< psubdiffcont >>
rect 1000 6220 1034 6254
rect 1068 6220 1102 6254
rect 1136 6220 1170 6254
rect 1204 6220 1238 6254
rect 1272 6220 1306 6254
rect 1340 6220 1374 6254
rect 1408 6220 1442 6254
rect 967 6102 1001 6136
rect 1480 6187 1514 6221
rect 1480 6119 1514 6153
rect 967 6034 1001 6068
rect 967 5966 1001 6000
rect 967 5898 1001 5932
rect 967 5830 1001 5864
rect 1480 6051 1514 6085
rect 1480 5983 1514 6017
rect 1480 5915 1514 5949
rect 1480 5847 1514 5881
rect 967 5762 1001 5796
rect 1480 5779 1514 5813
rect 967 5694 1001 5728
rect 967 5626 1001 5660
rect 1480 5711 1514 5745
rect 1480 5643 1514 5677
rect 967 5558 1001 5592
rect 967 5490 1001 5524
rect 967 5422 1001 5456
rect 1480 5575 1514 5609
rect 1480 5507 1514 5541
rect 967 5354 1001 5388
rect 967 5286 1001 5320
rect 1480 5439 1514 5473
rect 1480 5371 1514 5405
rect 1480 5303 1514 5337
rect 967 5218 1001 5252
rect 1480 5235 1514 5269
rect 967 5150 1001 5184
rect 967 5082 1001 5116
rect 967 5014 1001 5048
rect 1480 5167 1514 5201
rect 3292 5318 3326 5352
rect 3362 5318 3396 5352
rect 3433 5318 3467 5352
rect 3504 5318 3538 5352
rect 3575 5318 3609 5352
rect 3646 5318 3680 5352
rect 3717 5318 3751 5352
rect 3788 5318 3822 5352
rect 3859 5318 3893 5352
rect 3930 5318 3964 5352
rect 4001 5318 4035 5352
rect 4069 5321 4103 5355
rect 4137 5323 4171 5357
rect 3292 5250 3326 5284
rect 3362 5250 3396 5284
rect 3432 5250 3466 5284
rect 3502 5250 3536 5284
rect 3572 5250 3606 5284
rect 3643 5250 3677 5284
rect 3714 5250 3748 5284
rect 3785 5250 3819 5284
rect 3856 5250 3890 5284
rect 3927 5250 3961 5284
rect 3998 5250 4032 5284
rect 4069 5250 4103 5284
rect 4137 5255 4171 5289
rect 3292 5182 3326 5216
rect 3362 5182 3396 5216
rect 3432 5182 3466 5216
rect 3502 5182 3536 5216
rect 3572 5182 3606 5216
rect 3642 5182 3676 5216
rect 3712 5182 3746 5216
rect 3782 5182 3816 5216
rect 3852 5182 3886 5216
rect 3922 5182 3956 5216
rect 3992 5182 4026 5216
rect 4062 5182 4096 5216
rect 4132 5182 4166 5216
rect 1480 5099 1514 5133
rect 1480 5031 1514 5065
rect 967 4946 1001 4980
rect 967 4878 1001 4912
rect 967 4810 1001 4844
rect 1480 4963 1514 4997
rect 1480 4895 1514 4929
rect 967 4742 1001 4776
rect 967 4674 1001 4708
rect 967 4606 1001 4640
rect 967 4538 1001 4572
rect 967 4470 1001 4504
rect 967 4402 1001 4436
rect 967 4334 1001 4368
rect 283 4277 317 4311
rect 351 4277 385 4311
rect 419 4277 453 4311
rect 487 4277 521 4311
rect 555 4277 589 4311
rect 623 4277 657 4311
rect 691 4277 725 4311
rect 250 4208 284 4242
rect 250 4140 284 4174
rect 778 4244 812 4278
rect 778 4176 812 4210
rect 250 4072 284 4106
rect 250 4004 284 4038
rect 250 3936 284 3970
rect 250 3868 284 3902
rect 250 3800 284 3834
rect 250 3732 284 3766
rect 778 4108 812 4142
rect 778 4040 812 4074
rect 778 3972 812 4006
rect 778 3904 812 3938
rect 778 3836 812 3870
rect 778 3768 812 3802
rect 778 3700 812 3734
rect 778 3632 812 3666
rect 337 3515 371 3549
rect 405 3515 439 3549
rect 473 3515 507 3549
rect 541 3515 575 3549
rect 609 3515 643 3549
rect 677 3515 711 3549
rect 745 3515 779 3549
rect 967 4266 1001 4300
rect 967 4198 1001 4232
rect 967 4130 1001 4164
rect 967 4062 1001 4096
rect 967 3994 1001 4028
rect 967 3926 1001 3960
rect 1480 4827 1514 4861
rect 1480 4759 1514 4793
rect 1480 4691 1514 4725
rect 1480 4623 1514 4657
rect 1480 4555 1514 4589
rect 1480 4487 1514 4521
rect 1480 4419 1514 4453
rect 1480 4351 1514 4385
rect 1480 4283 1514 4317
rect 1480 4215 1514 4249
rect 1480 4147 1514 4181
rect 1480 4079 1514 4113
rect 1480 4011 1514 4045
rect 967 3858 1001 3892
rect 967 3790 1001 3824
rect 967 3722 1001 3756
rect 1480 3943 1514 3977
rect 1480 3875 1514 3909
rect 1480 3807 1514 3841
rect 967 3654 1001 3688
rect 967 3586 1001 3620
rect 967 3518 1001 3552
rect 967 3450 1001 3484
rect 1480 3739 1514 3773
rect 1480 3671 1514 3705
rect 1480 3603 1514 3637
rect 1480 3535 1514 3569
rect 1480 3467 1514 3501
rect 967 3382 1001 3416
rect 1480 3399 1514 3433
rect 1480 3331 1514 3365
rect 1480 3263 1514 3297
rect 1480 3195 1514 3229
rect 967 3088 1001 3122
rect 967 3020 1001 3054
rect 967 2952 1001 2986
rect 1480 3127 1514 3161
rect 1480 3059 1514 3093
rect 1480 2991 1514 3025
rect 967 2884 1001 2918
rect 967 2816 1001 2850
rect 967 2748 1001 2782
rect 1480 2923 1514 2957
rect 1480 2855 1514 2889
rect 1480 2787 1514 2821
rect 967 2680 1001 2714
rect 967 2612 1001 2646
rect 967 2544 1001 2578
rect 1480 2719 1514 2753
rect 1480 2651 1514 2685
rect 1480 2583 1514 2617
rect 967 2476 1001 2510
rect 1480 2515 1514 2549
rect 967 2408 1001 2442
rect 967 2340 1001 2374
rect 967 2272 1001 2306
rect 1480 2447 1514 2481
rect 1480 2379 1514 2413
rect 1480 2311 1514 2345
rect 967 2204 1001 2238
rect 1480 2243 1514 2277
rect 967 2136 1001 2170
rect 967 2068 1001 2102
rect 1480 2175 1514 2209
rect 1480 2107 1514 2141
rect 967 2000 1001 2034
rect 283 1911 317 1945
rect 351 1911 385 1945
rect 419 1911 453 1945
rect 487 1911 521 1945
rect 555 1911 589 1945
rect 623 1911 657 1945
rect 691 1911 725 1945
rect 250 1796 284 1830
rect 778 1878 812 1912
rect 778 1810 812 1844
rect 250 1728 284 1762
rect 250 1660 284 1694
rect 250 1592 284 1626
rect 250 1524 284 1558
rect 250 1456 284 1490
rect 250 1388 284 1422
rect 250 1320 284 1354
rect 778 1742 812 1776
rect 778 1674 812 1708
rect 778 1606 812 1640
rect 778 1538 812 1572
rect 778 1470 812 1504
rect 778 1402 812 1436
rect 778 1334 812 1368
rect 250 1252 284 1286
rect 250 1184 284 1218
rect 250 1116 284 1150
rect 778 1266 812 1300
rect 778 1198 812 1232
rect 250 1048 284 1082
rect 250 980 284 1014
rect 250 912 284 946
rect 250 844 284 878
rect 250 776 284 810
rect 250 708 284 742
rect 250 640 284 674
rect 250 572 284 606
rect 250 504 284 538
rect 778 1130 812 1164
rect 778 1062 812 1096
rect 778 994 812 1028
rect 778 926 812 960
rect 778 858 812 892
rect 778 790 812 824
rect 778 722 812 756
rect 778 654 812 688
rect 778 586 812 620
rect 778 518 812 552
rect 250 436 284 470
rect 250 368 284 402
rect 778 450 812 484
rect 337 335 371 369
rect 405 335 439 369
rect 473 335 507 369
rect 541 335 575 369
rect 609 335 643 369
rect 677 335 711 369
rect 745 335 779 369
rect 967 1932 1001 1966
rect 967 1864 1001 1898
rect 1480 2039 1514 2073
rect 1480 1971 1514 2005
rect 1480 1903 1514 1937
rect 967 1796 1001 1830
rect 967 1728 1001 1762
rect 967 1660 1001 1694
rect 967 1592 1001 1626
rect 1480 1835 1514 1869
rect 1480 1767 1514 1801
rect 1480 1699 1514 1733
rect 1480 1631 1514 1665
rect 967 1524 1001 1558
rect 967 1456 1001 1490
rect 967 1388 1001 1422
rect 1480 1563 1514 1597
rect 1480 1495 1514 1529
rect 1480 1427 1514 1461
rect 967 1320 1001 1354
rect 967 1252 1001 1286
rect 967 1184 1001 1218
rect 967 1116 1001 1150
rect 967 1048 1001 1082
rect 967 980 1001 1014
rect 967 912 1001 946
rect 967 844 1001 878
rect 967 776 1001 810
rect 967 708 1001 742
rect 967 640 1001 674
rect 967 572 1001 606
rect 967 504 1001 538
rect 1480 1359 1514 1393
rect 1480 1291 1514 1325
rect 1480 1223 1514 1257
rect 1480 1155 1514 1189
rect 1480 1087 1514 1121
rect 1480 1019 1514 1053
rect 1480 951 1514 985
rect 1480 883 1514 917
rect 1480 815 1514 849
rect 1480 747 1514 781
rect 1480 679 1514 713
rect 1480 611 1514 645
rect 1480 543 1514 577
rect 967 436 1001 470
rect 967 368 1001 402
rect 1480 475 1514 509
rect 1039 335 1073 369
rect 1107 335 1141 369
rect 1175 335 1209 369
rect 1243 335 1277 369
rect 1311 335 1345 369
rect 1379 335 1413 369
rect 1447 335 1481 369
rect 3268 5095 3302 5129
rect 3336 5095 3370 5129
rect 3404 5095 3438 5129
rect 3490 5096 3524 5130
rect 3558 5096 3592 5130
rect 3626 5096 3660 5130
rect 3730 5114 3764 5148
rect 3798 5114 3832 5148
rect 3866 5114 3900 5148
rect 3934 5114 3968 5148
rect 4002 5114 4036 5148
rect 4070 5114 4104 5148
rect 4138 5114 4172 5148
rect 4206 5114 4240 5148
rect 3268 5026 3302 5060
rect 3336 5026 3370 5060
rect 3404 5026 3438 5060
rect 3490 5027 3524 5061
rect 3558 5027 3592 5061
rect 3626 5027 3660 5061
rect 3696 5008 3730 5042
rect 3268 4957 3302 4991
rect 3336 4957 3370 4991
rect 3404 4957 3438 4991
rect 3268 4888 3302 4922
rect 3336 4888 3370 4922
rect 3404 4888 3438 4922
rect 3268 4819 3302 4853
rect 3336 4819 3370 4853
rect 3404 4819 3438 4853
rect 3268 4750 3302 4784
rect 3336 4750 3370 4784
rect 3404 4750 3438 4784
rect 3268 4681 3302 4715
rect 3336 4681 3370 4715
rect 3404 4681 3438 4715
rect 3268 4612 3302 4646
rect 3336 4612 3370 4646
rect 3404 4612 3438 4646
rect 3268 4543 3302 4577
rect 3336 4543 3370 4577
rect 3404 4543 3438 4577
rect 3268 4474 3302 4508
rect 3336 4474 3370 4508
rect 3404 4474 3438 4508
rect 3268 4405 3302 4439
rect 3336 4405 3370 4439
rect 3404 4405 3438 4439
rect 3268 4336 3302 4370
rect 3336 4336 3370 4370
rect 3404 4336 3438 4370
rect 3268 4267 3302 4301
rect 3336 4267 3370 4301
rect 3404 4267 3438 4301
rect 3268 4198 3302 4232
rect 3336 4198 3370 4232
rect 3404 4198 3438 4232
rect 3268 4129 3302 4163
rect 3336 4129 3370 4163
rect 3404 4129 3438 4163
rect 3268 4060 3302 4094
rect 3336 4060 3370 4094
rect 3404 4060 3438 4094
rect 3268 3991 3302 4025
rect 3336 3991 3370 4025
rect 3404 3991 3438 4025
rect 3268 3922 3302 3956
rect 3336 3922 3370 3956
rect 3404 3922 3438 3956
rect 3268 3853 3302 3887
rect 3336 3853 3370 3887
rect 3404 3853 3438 3887
rect 3268 3784 3302 3818
rect 3336 3784 3370 3818
rect 3404 3784 3438 3818
rect 3268 3715 3302 3749
rect 3336 3715 3370 3749
rect 3404 3715 3438 3749
rect 3268 3646 3302 3680
rect 3336 3646 3370 3680
rect 3404 3646 3438 3680
rect 3268 3577 3302 3611
rect 3336 3577 3370 3611
rect 3404 3577 3438 3611
rect 3268 3508 3302 3542
rect 3336 3508 3370 3542
rect 3404 3508 3438 3542
rect 3490 3530 3660 4992
rect 3696 4940 3730 4974
rect 4266 5014 4300 5048
rect 3696 4872 3730 4906
rect 3696 4804 3730 4838
rect 4266 4946 4300 4980
rect 4266 4878 4300 4912
rect 4266 4810 4300 4844
rect 3696 4736 3730 4770
rect 3696 4668 3730 4702
rect 3696 4600 3730 4634
rect 3696 4532 3730 4566
rect 3696 4464 3730 4498
rect 4266 4742 4300 4776
rect 4266 4674 4300 4708
rect 4266 4606 4300 4640
rect 4266 4538 4300 4572
rect 3696 4396 3730 4430
rect 3696 4328 3730 4362
rect 3696 4260 3730 4294
rect 3696 4192 3730 4226
rect 3696 4124 3730 4158
rect 3696 4056 3730 4090
rect 3696 3988 3730 4022
rect 3696 3920 3730 3954
rect 3696 3852 3730 3886
rect 3696 3784 3730 3818
rect 3696 3716 3730 3750
rect 3696 3648 3730 3682
rect 3696 3580 3730 3614
rect 4266 4470 4300 4504
rect 4266 4402 4300 4436
rect 4266 4334 4300 4368
rect 4266 4266 4300 4300
rect 4266 4198 4300 4232
rect 4266 4130 4300 4164
rect 4266 4062 4300 4096
rect 4266 3994 4300 4028
rect 4266 3926 4300 3960
rect 4266 3858 4300 3892
rect 4266 3790 4300 3824
rect 4266 3722 4300 3756
rect 4266 3654 4300 3688
rect 3696 3512 3730 3546
rect 3268 3439 3302 3473
rect 3336 3439 3370 3473
rect 3404 3439 3438 3473
rect 3696 3444 3730 3478
rect 3268 3370 3302 3404
rect 3336 3370 3370 3404
rect 3404 3370 3438 3404
rect 3268 3301 3302 3335
rect 3336 3301 3370 3335
rect 3404 3301 3438 3335
rect 3696 3376 3730 3410
rect 3696 3308 3730 3342
rect 3268 3232 3302 3266
rect 3336 3232 3370 3266
rect 3404 3232 3438 3266
rect 3268 3163 3302 3197
rect 3336 3163 3370 3197
rect 3404 3163 3438 3197
rect 3268 374 3438 3128
rect 3696 3240 3730 3274
rect 3696 3172 3730 3206
rect 3696 3104 3730 3138
rect 4266 3586 4300 3620
rect 4266 3518 4300 3552
rect 4266 3450 4300 3484
rect 4266 3382 4300 3416
rect 4266 3314 4300 3348
rect 4266 3246 4300 3280
rect 4266 3178 4300 3212
rect 4266 3110 4300 3144
rect 3696 3036 3730 3070
rect 3696 2968 3730 3002
rect 3696 2900 3730 2934
rect 3696 2832 3730 2866
rect 3696 2764 3730 2798
rect 3696 2696 3730 2730
rect 3696 2628 3730 2662
rect 3696 2560 3730 2594
rect 3696 2492 3730 2526
rect 3696 2424 3730 2458
rect 4266 3042 4300 3076
rect 4266 2974 4300 3008
rect 4266 2906 4300 2940
rect 4266 2838 4300 2872
rect 4266 2770 4300 2804
rect 4266 2702 4300 2736
rect 4266 2634 4300 2668
rect 4266 2566 4300 2600
rect 4266 2498 4300 2532
rect 4266 2430 4300 2464
rect 3696 2356 3730 2390
rect 3696 2288 3730 2322
rect 3696 2220 3730 2254
rect 3696 2152 3730 2186
rect 4266 2362 4300 2396
rect 4266 2294 4300 2328
rect 4266 2226 4300 2260
rect 4266 2158 4300 2192
rect 3696 2084 3730 2118
rect 3696 2016 3730 2050
rect 3696 1948 3730 1982
rect 4266 2090 4300 2124
rect 4266 2022 4300 2056
rect 3490 1883 3524 1917
rect 3558 1883 3592 1917
rect 3626 1883 3660 1917
rect 3696 1880 3730 1914
rect 3490 1814 3524 1848
rect 3558 1814 3592 1848
rect 3626 1814 3660 1848
rect 3696 1812 3730 1846
rect 3490 1745 3524 1779
rect 3558 1745 3592 1779
rect 3626 1745 3660 1779
rect 3696 1744 3730 1778
rect 3490 1676 3524 1710
rect 3558 1676 3592 1710
rect 3626 1676 3660 1710
rect 3696 1676 3730 1710
rect 3490 1607 3524 1641
rect 3558 1607 3592 1641
rect 3626 1607 3660 1641
rect 3696 1608 3730 1642
rect 3490 1538 3524 1572
rect 3558 1538 3592 1572
rect 3626 1538 3660 1572
rect 3696 1540 3730 1574
rect 3490 1469 3524 1503
rect 3558 1469 3592 1503
rect 3626 1469 3660 1503
rect 3696 1472 3730 1506
rect 3490 1400 3524 1434
rect 3558 1400 3592 1434
rect 3626 1400 3660 1434
rect 3696 1404 3730 1438
rect 4266 1954 4300 1988
rect 4266 1886 4300 1920
rect 4266 1818 4300 1852
rect 4266 1750 4300 1784
rect 4266 1682 4300 1716
rect 4266 1614 4300 1648
rect 4266 1546 4300 1580
rect 4266 1478 4300 1512
rect 4266 1410 4300 1444
rect 3490 1331 3524 1365
rect 3558 1331 3592 1365
rect 3626 1331 3660 1365
rect 3696 1336 3730 1370
rect 3490 1262 3524 1296
rect 3558 1262 3592 1296
rect 3626 1262 3660 1296
rect 3696 1268 3730 1302
rect 3490 1193 3524 1227
rect 3558 1193 3592 1227
rect 3626 1193 3660 1227
rect 3696 1200 3730 1234
rect 3490 1124 3524 1158
rect 3558 1124 3592 1158
rect 3626 1124 3660 1158
rect 3696 1132 3730 1166
rect 3490 1055 3524 1089
rect 3558 1055 3592 1089
rect 3626 1055 3660 1089
rect 3696 1064 3730 1098
rect 3490 374 3660 1020
rect 3696 996 3730 1030
rect 3696 928 3730 962
rect 3696 860 3730 894
rect 3696 792 3730 826
rect 3696 724 3730 758
rect 3696 656 3730 690
rect 3696 588 3730 622
rect 3696 520 3730 554
rect 4266 1342 4300 1376
rect 4266 1274 4300 1308
rect 4266 1206 4300 1240
rect 4266 1138 4300 1172
rect 4266 1070 4300 1104
rect 4266 1002 4300 1036
rect 4266 934 4300 968
rect 4266 866 4300 900
rect 4266 798 4300 832
rect 4266 730 4300 764
rect 4266 662 4300 696
rect 4266 594 4300 628
rect 3696 452 3730 486
rect 3696 384 3730 418
rect 4266 526 4300 560
rect 4266 458 4300 492
rect 3824 350 3858 384
rect 3892 350 3926 384
rect 3960 350 3994 384
rect 4028 350 4062 384
rect 4096 350 4130 384
rect 4164 350 4198 384
rect 4232 350 4266 384
rect 12675 4370 12709 4404
rect 12675 4302 12709 4336
rect 12675 4234 12709 4268
rect 12675 4166 12709 4200
rect 12675 4098 12709 4132
rect 12675 4030 12709 4064
rect 12675 3962 12709 3996
rect 12675 3894 12709 3928
rect 12675 3826 12709 3860
rect 12675 3758 12709 3792
rect 12675 3690 12709 3724
rect 12675 3622 12709 3656
rect 12675 3554 12709 3588
rect 12675 3486 12709 3520
rect 12675 3418 12709 3452
rect 12675 3350 12709 3384
rect 12675 3282 12709 3316
rect 12675 3214 12709 3248
rect 12675 3146 12709 3180
rect 12675 3078 12709 3112
rect 12675 3010 12709 3044
rect 12675 2942 12709 2976
rect 12675 2874 12709 2908
rect 12675 2806 12709 2840
rect 12675 2738 12709 2772
rect 12675 2670 12709 2704
rect 12675 2602 12709 2636
rect 12675 2534 12709 2568
rect 12675 2466 12709 2500
rect 12675 2398 12709 2432
rect 12675 2330 12709 2364
rect 12675 2262 12709 2296
rect 12675 2194 12709 2228
rect 12675 2126 12709 2160
rect 12675 2058 12709 2092
rect 12675 1990 12709 2024
rect 12675 1922 12709 1956
rect 12675 1854 12709 1888
rect 12675 1786 12709 1820
rect 12675 1718 12709 1752
rect 12675 1650 12709 1684
rect 12675 1582 12709 1616
rect 12675 1514 12709 1548
rect 12675 1446 12709 1480
rect 12675 1378 12709 1412
rect 12675 1310 12709 1344
rect 12675 1242 12709 1276
rect 12675 1174 12709 1208
rect 12675 1106 12709 1140
rect 12675 1038 12709 1072
rect 12675 970 12709 1004
rect 12675 902 12709 936
rect 12675 834 12709 868
rect 12675 766 12709 800
rect 12675 698 12709 732
<< nsubdiffcont >>
rect 283 3326 317 3360
rect 351 3326 385 3360
rect 419 3326 453 3360
rect 555 3326 589 3360
rect 623 3326 657 3360
rect 691 3326 725 3360
rect 250 3256 284 3290
rect 250 3188 284 3222
rect 778 3293 812 3327
rect 778 3225 812 3259
rect 250 3120 284 3154
rect 250 3052 284 3086
rect 778 3157 812 3191
rect 778 3089 812 3123
rect 778 3021 812 3055
rect 778 2953 812 2987
rect 250 2745 284 2779
rect 250 2677 284 2711
rect 778 2885 812 2919
rect 778 2817 812 2851
rect 778 2749 812 2783
rect 250 2609 284 2643
rect 250 2541 284 2575
rect 778 2681 812 2715
rect 778 2613 812 2647
rect 250 2473 284 2507
rect 250 2405 284 2439
rect 778 2545 812 2579
rect 778 2477 812 2511
rect 250 2337 284 2371
rect 778 2409 812 2443
rect 250 2269 284 2303
rect 250 2201 284 2235
rect 778 2341 812 2375
rect 778 2273 812 2307
rect 250 2133 284 2167
rect 337 2100 371 2134
rect 405 2100 439 2134
rect 473 2100 507 2134
rect 541 2100 575 2134
rect 609 2100 643 2134
rect 677 2100 711 2134
rect 745 2100 779 2134
<< mvpsubdiffcont >>
rect 10070 12082 10104 12116
rect 10155 12082 10189 12116
rect 10240 12082 10274 12116
rect 10325 12082 10359 12116
rect 10410 12082 10444 12116
rect 10495 12082 10529 12116
rect 10580 12082 10614 12116
rect 10665 12082 10699 12116
rect 10750 12082 10784 12116
rect 10835 12082 10869 12116
rect 10920 12082 10954 12116
rect 11005 12082 11039 12116
rect 11090 12082 11124 12116
rect 11175 12082 11209 12116
rect 11260 12082 11294 12116
rect 11345 12082 11379 12116
rect 11430 12082 11464 12116
rect 11515 12082 11549 12116
rect 11600 12082 11634 12116
rect 11685 12082 11719 12116
rect 11770 12082 11804 12116
rect 11856 12082 11890 12116
rect 11942 12082 11976 12116
rect 12022 11993 12056 12027
rect 12022 11900 12056 11934
rect 12022 11807 12056 11841
rect 12022 11714 12056 11748
rect 12022 11621 12056 11655
rect 12022 11528 12056 11562
rect 12022 11435 12056 11469
rect 12022 11342 12056 11376
rect 12022 11249 12056 11283
rect 10066 11169 10100 11203
rect 10152 11169 10186 11203
rect 10238 11169 10272 11203
rect 10324 11169 10358 11203
rect 10410 11169 10444 11203
rect 10496 11169 10530 11203
rect 10582 11169 10616 11203
rect 10668 11169 10702 11203
rect 10754 11169 10788 11203
rect 10840 11169 10874 11203
rect 10927 11169 10961 11203
rect 11014 11169 11048 11203
rect 11101 11169 11135 11203
rect 11188 11169 11222 11203
rect 11275 11169 11309 11203
rect 11362 11169 11396 11203
rect 11449 11169 11483 11203
rect 11536 11169 11570 11203
rect 11623 11169 11657 11203
rect 11765 11169 11799 11203
rect 11852 11169 11886 11203
rect 11939 11169 11973 11203
rect 6322 11074 6356 11108
rect 6322 10989 6356 11023
rect 6322 10903 6356 10937
rect 6322 10817 6356 10851
rect 6322 10731 6356 10765
rect 6322 10645 6356 10679
rect 6322 10559 6356 10593
rect 6322 10473 6356 10507
rect 11703 11086 11737 11120
rect 11703 10999 11737 11033
rect 11703 10911 11737 10945
rect 11703 10823 11737 10857
rect 11703 10735 11737 10769
rect 11703 10647 11737 10681
rect 11703 10559 11737 10593
rect 11703 10471 11737 10505
rect 6322 10387 6356 10421
rect 11703 10383 11737 10417
rect 6322 10301 6356 10335
rect 6417 10303 6451 10337
rect 6503 10303 6537 10337
rect 6589 10303 6623 10337
rect 6675 10303 6709 10337
rect 6761 10303 6795 10337
rect 6847 10303 6881 10337
rect 6933 10303 6967 10337
rect 7019 10303 7053 10337
rect 7105 10303 7139 10337
rect 7191 10303 7225 10337
rect 7277 10303 7311 10337
rect 7363 10303 7397 10337
rect 7449 10303 7483 10337
rect 7535 10303 7569 10337
rect 7621 10303 7655 10337
rect 7707 10303 7741 10337
rect 7793 10303 7827 10337
rect 7879 10303 7913 10337
rect 7965 10303 7999 10337
rect 8051 10303 8085 10337
rect 8137 10303 8171 10337
rect 8222 10303 8256 10337
rect 8307 10303 8341 10337
rect 8392 10303 8426 10337
rect 8477 10303 8511 10337
rect 8562 10303 8596 10337
rect 8647 10303 8681 10337
rect 8732 10303 8766 10337
rect 8817 10303 8851 10337
rect 8902 10303 8936 10337
rect 8987 10303 9021 10337
rect 9072 10303 9106 10337
rect 9157 10303 9191 10337
rect 9242 10303 9276 10337
rect 9327 10303 9361 10337
rect 9412 10303 9446 10337
rect 9497 10303 9531 10337
rect 9582 10303 9616 10337
rect 9667 10303 9701 10337
rect 9752 10303 9786 10337
rect 9837 10303 9871 10337
rect 9922 10303 9956 10337
rect 10007 10303 10041 10337
rect 10092 10303 10126 10337
rect 10177 10303 10211 10337
rect 10262 10303 10296 10337
rect 10347 10303 10381 10337
rect 10432 10303 10466 10337
rect 10517 10303 10551 10337
rect 10602 10303 10636 10337
rect 10687 10303 10721 10337
rect 10772 10303 10806 10337
rect 10857 10303 10891 10337
rect 10942 10303 10976 10337
rect 11027 10303 11061 10337
rect 11112 10303 11146 10337
rect 11197 10303 11231 10337
rect 11282 10303 11316 10337
rect 11367 10303 11401 10337
rect 11452 10303 11486 10337
rect 11537 10303 11571 10337
rect 11622 10303 11656 10337
rect 6322 10215 6356 10249
rect 6322 10129 6356 10163
rect 6322 10043 6356 10077
rect 6322 9957 6356 9991
rect 6322 9871 6356 9905
rect 6322 9785 6356 9819
rect 6322 9699 6356 9733
rect 6322 9613 6356 9647
rect 10033 10204 10067 10238
rect 10033 10119 10067 10153
rect 10033 10034 10067 10068
rect 10033 9949 10067 9983
rect 10033 9864 10067 9898
rect 10033 9778 10067 9812
rect 10033 9692 10067 9726
rect 10033 9606 10067 9640
rect 6322 9527 6356 9561
rect 10033 9520 10067 9554
rect 6322 9441 6356 9475
rect 6322 9355 6356 9389
rect 6322 9269 6356 9303
rect 6322 9183 6356 9217
rect 6322 9097 6356 9131
rect 6322 9011 6356 9045
rect 6322 8925 6356 8959
rect 6322 8839 6356 8873
rect 6322 8753 6356 8787
rect 10033 9434 10067 9468
rect 10033 9348 10067 9382
rect 10033 9262 10067 9296
rect 10033 9176 10067 9210
rect 10033 9090 10067 9124
rect 10033 9004 10067 9038
rect 10033 8918 10067 8952
rect 10033 8832 10067 8866
rect 4868 5083 4902 5117
rect 4936 5083 4970 5117
rect 5004 5083 5038 5117
rect 5072 5083 5106 5117
rect 5140 5083 5174 5117
rect 5208 5083 5242 5117
rect 5276 5083 5310 5117
rect 5344 5083 5378 5117
rect 5412 5083 5446 5117
rect 5480 5083 5514 5117
rect 5548 5083 5582 5117
rect 5616 5083 5650 5117
rect 5684 5083 5718 5117
rect 5752 5083 5786 5117
rect 5820 5083 5854 5117
rect 5888 5083 5922 5117
rect 5956 5083 5990 5117
rect 6024 5083 6058 5117
rect 6092 5083 6126 5117
rect 6160 5083 6194 5117
rect 6228 5083 6262 5117
rect 6296 5083 6330 5117
rect 6364 5083 6398 5117
rect 6432 5083 6466 5117
rect 6500 5083 6534 5117
rect 6568 5083 6602 5117
rect 6636 5083 6670 5117
rect 6704 5083 6738 5117
rect 6772 5083 6806 5117
rect 6840 5083 6874 5117
rect 6908 5083 6942 5117
rect 6976 5083 7010 5117
rect 7044 5083 7078 5117
rect 7112 5083 7146 5117
rect 7180 5083 7214 5117
rect 7248 5083 7282 5117
rect 7316 5083 7350 5117
rect 7384 5083 7418 5117
rect 7452 5083 7486 5117
rect 7520 5083 7554 5117
rect 7588 5083 7622 5117
rect 7656 5083 7690 5117
rect 7724 5083 7758 5117
rect 7792 5083 7826 5117
rect 7860 5083 7894 5117
rect 7928 5083 7962 5117
rect 7996 5083 8030 5117
rect 8064 5083 8098 5117
rect 8132 5083 8166 5117
rect 8200 5083 8234 5117
rect 8268 5083 8302 5117
rect 8336 5083 8370 5117
rect 8404 5083 8438 5117
rect 8472 5083 8506 5117
rect 8540 5083 8574 5117
rect 8608 5083 8642 5117
rect 8676 5083 8710 5117
rect 8744 5083 8778 5117
rect 8812 5083 8846 5117
rect 8880 5083 8914 5117
rect 8948 5083 8982 5117
rect 9016 5083 9050 5117
rect 9084 5083 9118 5117
rect 9152 5083 9186 5117
rect 9220 5083 9254 5117
rect 9288 5083 9322 5117
rect 9356 5083 9390 5117
rect 9424 5083 9458 5117
rect 9492 5083 9526 5117
rect 9560 5083 9594 5117
rect 9628 5083 9662 5117
rect 9696 5083 9730 5117
rect 9764 5083 9798 5117
rect 9832 5083 9866 5117
rect 9900 5083 9934 5117
rect 9968 5083 10002 5117
rect 10036 5083 10070 5117
rect 10104 5083 10138 5117
rect 10172 5083 10206 5117
rect 10240 5083 10274 5117
rect 10308 5083 10342 5117
rect 10376 5083 10410 5117
rect 10444 5083 10478 5117
rect 10512 5083 10546 5117
rect 10580 5083 10614 5117
rect 10648 5083 10682 5117
rect 10716 5083 10750 5117
rect 10784 5083 10818 5117
rect 10852 5083 10886 5117
rect 10920 5083 10954 5117
rect 10988 5083 11022 5117
rect 11056 5083 11090 5117
rect 11124 5083 11158 5117
rect 11192 5083 11226 5117
rect 11260 5083 11294 5117
rect 11328 5083 11362 5117
rect 11396 5083 11430 5117
rect 11464 5083 11498 5117
rect 11532 5083 11566 5117
rect 11600 5083 11634 5117
rect 11668 5083 11702 5117
rect 11736 5083 11770 5117
rect 11804 5083 11838 5117
rect 11872 5083 11906 5117
rect 11940 5083 11974 5117
rect 12008 5083 12042 5117
rect 12076 5083 12110 5117
rect 12144 5083 12178 5117
rect 12212 5083 12246 5117
rect 12280 5083 12314 5117
rect 12348 5083 12382 5117
rect 12416 5083 12450 5117
rect 12484 5083 12518 5117
rect 12552 5083 12586 5117
rect 4835 5003 4869 5037
rect 4835 4935 4869 4969
rect 4835 4867 4869 4901
rect 4835 4799 4869 4833
rect 4835 4731 4869 4765
rect 4835 4663 4869 4697
rect 4835 4595 4869 4629
rect 4835 4527 4869 4561
rect 10296 5012 10330 5046
rect 9468 4953 9502 4987
rect 10296 4944 10330 4978
rect 9468 4885 9502 4919
rect 9468 4817 9502 4851
rect 9468 4749 9502 4783
rect 9468 4681 9502 4715
rect 9468 4613 9502 4647
rect 9468 4545 9502 4579
rect 4835 4459 4869 4493
rect 9468 4477 9502 4511
rect 4835 4391 4869 4425
rect 9468 4409 9502 4443
rect 4835 4323 4869 4357
rect 9468 4341 9502 4375
rect 4835 4255 4869 4289
rect 4835 4187 4869 4221
rect 4835 4119 4869 4153
rect 4835 4051 4869 4085
rect 4835 3983 4869 4017
rect 4835 3915 4869 3949
rect 4835 3847 4869 3881
rect 4835 3779 4869 3813
rect 4835 3711 4869 3745
rect 9468 4273 9502 4307
rect 9468 4205 9502 4239
rect 9468 4137 9502 4171
rect 9468 4069 9502 4103
rect 9468 4001 9502 4035
rect 9468 3933 9502 3967
rect 9468 3865 9502 3899
rect 9468 3797 9502 3831
rect 4963 3710 4997 3744
rect 5032 3710 5066 3744
rect 5101 3710 5135 3744
rect 5170 3710 5204 3744
rect 5239 3710 5273 3744
rect 5308 3710 5342 3744
rect 5377 3710 5411 3744
rect 5446 3710 5480 3744
rect 5515 3710 5549 3744
rect 5584 3710 5618 3744
rect 5653 3710 5687 3744
rect 5722 3710 5756 3744
rect 5791 3710 5825 3744
rect 5860 3710 5894 3744
rect 4835 3643 4869 3677
rect 4963 3642 4997 3676
rect 5032 3642 5066 3676
rect 5101 3642 5135 3676
rect 5170 3642 5204 3676
rect 5239 3642 5273 3676
rect 5308 3642 5342 3676
rect 5377 3642 5411 3676
rect 5446 3642 5480 3676
rect 5515 3642 5549 3676
rect 5584 3642 5618 3676
rect 5653 3642 5687 3676
rect 5722 3642 5756 3676
rect 5791 3642 5825 3676
rect 5860 3642 5894 3676
rect 5929 3642 9363 3744
rect 9468 3729 9502 3763
rect 9468 3661 9502 3695
rect 4835 3575 4869 3609
rect 4835 3507 4869 3541
rect 9468 3593 9502 3627
rect 9468 3525 9502 3559
rect 4835 3439 4869 3473
rect 4835 3371 4869 3405
rect 4835 3303 4869 3337
rect 9468 3457 9502 3491
rect 9468 3389 9502 3423
rect 9468 3321 9502 3355
rect 4835 3235 4869 3269
rect 4835 3167 4869 3201
rect 4835 3099 4869 3133
rect 9468 3253 9502 3287
rect 9468 3185 9502 3219
rect 4835 3031 4869 3065
rect 4835 2963 4869 2997
rect 9468 3117 9502 3151
rect 9468 3049 9502 3083
rect 9468 2981 9502 3015
rect 4835 2895 4869 2929
rect 9468 2913 9502 2947
rect 4835 2827 4869 2861
rect 4835 2759 4869 2793
rect 4835 2691 4869 2725
rect 9468 2845 9502 2879
rect 9468 2777 9502 2811
rect 4835 2623 4869 2657
rect 4835 2555 4869 2589
rect 9468 2709 9502 2743
rect 9468 2641 9502 2675
rect 9468 2573 9502 2607
rect 4835 2487 4869 2521
rect 4835 2419 4869 2453
rect 4835 2351 4869 2385
rect 9468 2505 9502 2539
rect 9468 2437 9502 2471
rect 9468 2368 9502 2402
rect 4835 2283 4869 2317
rect 9468 2299 9502 2333
rect 4835 2215 4869 2249
rect 4835 2147 4869 2181
rect 9468 2230 9502 2264
rect 9468 2161 9502 2195
rect 4835 2079 4869 2113
rect 4835 2011 4869 2045
rect 4835 1943 4869 1977
rect 9468 2092 9502 2126
rect 9468 2023 9502 2057
rect 9468 1954 9502 1988
rect 4835 1875 4869 1909
rect 4835 1807 4869 1841
rect 4835 1739 4869 1773
rect 9468 1885 9502 1919
rect 9468 1816 9502 1850
rect 4835 1671 4869 1705
rect 4835 1603 4869 1637
rect 9468 1747 9502 1781
rect 9468 1678 9502 1712
rect 9468 1609 9502 1643
rect 4963 1571 4997 1605
rect 5032 1571 5066 1605
rect 5101 1571 5135 1605
rect 5170 1571 5204 1605
rect 5239 1571 5273 1605
rect 5308 1571 5342 1605
rect 5377 1571 5411 1605
rect 5446 1571 5480 1605
rect 5515 1571 5549 1605
rect 5584 1571 5618 1605
rect 5653 1571 5687 1605
rect 5722 1571 5756 1605
rect 5791 1571 5825 1605
rect 5860 1571 5894 1605
rect 4835 1535 4869 1569
rect 4963 1503 4997 1537
rect 5032 1503 5066 1537
rect 5101 1503 5135 1537
rect 5170 1503 5204 1537
rect 5239 1503 5273 1537
rect 5308 1503 5342 1537
rect 5377 1503 5411 1537
rect 5446 1503 5480 1537
rect 5515 1503 5549 1537
rect 5584 1503 5618 1537
rect 5653 1503 5687 1537
rect 5722 1503 5756 1537
rect 5791 1503 5825 1537
rect 5860 1503 5894 1537
rect 5929 1503 9363 1605
rect 9468 1540 9502 1574
rect 4835 1467 4869 1501
rect 4835 1399 4869 1433
rect 4835 1331 4869 1365
rect 4835 1263 4869 1297
rect 4835 1195 4869 1229
rect 4835 1127 4869 1161
rect 4835 1059 4869 1093
rect 9468 1471 9502 1505
rect 9468 1402 9502 1436
rect 9468 1333 9502 1367
rect 9468 1264 9502 1298
rect 9468 1195 9502 1229
rect 9468 1126 9502 1160
rect 9468 1057 9502 1091
rect 4835 991 4869 1025
rect 9468 988 9502 1022
rect 4835 923 4869 957
rect 9468 919 9502 953
rect 4835 855 4869 889
rect 9468 850 9502 884
rect 4835 787 4869 821
rect 4835 719 4869 753
rect 4835 651 4869 685
rect 4835 583 4869 617
rect 4835 515 4869 549
rect 4835 447 4869 481
rect 4835 379 4869 413
rect 4835 311 4869 345
rect 4835 243 4869 277
rect 9468 781 9502 815
rect 9468 712 9502 746
rect 9468 643 9502 677
rect 10296 4876 10330 4910
rect 12675 5050 12709 5084
rect 12675 4982 12709 5016
rect 12675 4914 12709 4948
rect 10296 4808 10330 4842
rect 10296 4740 10330 4774
rect 10296 4672 10330 4706
rect 10296 4604 10330 4638
rect 10296 4536 10330 4570
rect 10296 4468 10330 4502
rect 10296 4400 10330 4434
rect 10296 4332 10330 4366
rect 10296 4264 10330 4298
rect 10296 4196 10330 4230
rect 10296 4128 10330 4162
rect 10296 4060 10330 4094
rect 12675 4846 12709 4880
rect 12675 4778 12709 4812
rect 12675 4710 12709 4744
rect 12675 4642 12709 4676
rect 12675 4574 12709 4608
rect 12675 4506 12709 4540
rect 12675 4438 12709 4472
rect 10296 3992 10330 4026
rect 10296 3924 10330 3958
rect 10296 3856 10330 3890
rect 10296 3788 10330 3822
rect 10296 3720 10330 3754
rect 10296 3652 10330 3686
rect 10296 3584 10330 3618
rect 10296 3516 10330 3550
rect 10296 3448 10330 3482
rect 10296 3380 10330 3414
rect 10296 3312 10330 3346
rect 10296 3244 10330 3278
rect 10296 3176 10330 3210
rect 10296 3108 10330 3142
rect 10296 3040 10330 3074
rect 10296 2972 10330 3006
rect 10296 2904 10330 2938
rect 10296 2836 10330 2870
rect 10296 2768 10330 2802
rect 10296 2700 10330 2734
rect 10296 2632 10330 2666
rect 10296 2564 10330 2598
rect 10296 2496 10330 2530
rect 10296 2428 10330 2462
rect 10296 2360 10330 2394
rect 10296 2292 10330 2326
rect 10296 2224 10330 2258
rect 10296 2156 10330 2190
rect 10296 2088 10330 2122
rect 10296 2020 10330 2054
rect 10296 1952 10330 1986
rect 10296 1884 10330 1918
rect 10296 1816 10330 1850
rect 10296 1748 10330 1782
rect 10296 1680 10330 1714
rect 10296 1612 10330 1646
rect 10296 1544 10330 1578
rect 10296 1476 10330 1510
rect 10296 1408 10330 1442
rect 10296 1340 10330 1374
rect 10296 1272 10330 1306
rect 10296 1204 10330 1238
rect 10296 1136 10330 1170
rect 10296 1068 10330 1102
rect 10296 1000 10330 1034
rect 10296 932 10330 966
rect 10296 864 10330 898
rect 10296 796 10330 830
rect 10296 728 10330 762
rect 10296 660 10330 694
rect 9468 574 9502 608
rect 10296 592 10330 626
rect 9468 505 9502 539
rect 10296 524 10330 558
rect 12675 574 12709 608
rect 9468 436 9502 470
rect 9582 455 9616 489
rect 9650 455 9684 489
rect 9718 455 9752 489
rect 9786 455 9820 489
rect 9854 455 9888 489
rect 9922 455 9956 489
rect 9990 455 10024 489
rect 10058 455 10092 489
rect 10126 455 10160 489
rect 10194 455 10228 489
rect 10262 455 10296 489
rect 10330 455 10364 489
rect 10398 455 10432 489
rect 10466 455 10500 489
rect 10534 455 10568 489
rect 10602 455 10636 489
rect 10670 455 10704 489
rect 10738 455 10772 489
rect 10806 455 10840 489
rect 10874 455 10908 489
rect 10942 455 10976 489
rect 11010 455 11044 489
rect 11078 455 11112 489
rect 11146 455 11180 489
rect 11214 455 11248 489
rect 11282 455 11316 489
rect 11350 455 11384 489
rect 11418 455 11452 489
rect 11486 455 11520 489
rect 11554 455 11588 489
rect 11622 455 11656 489
rect 11690 455 11724 489
rect 11758 455 11792 489
rect 11826 455 11860 489
rect 11894 455 11928 489
rect 11962 455 11996 489
rect 12030 455 12064 489
rect 12098 455 12132 489
rect 12166 455 12200 489
rect 12234 455 12268 489
rect 12302 455 12336 489
rect 12370 455 12404 489
rect 12438 455 12472 489
rect 12506 455 12540 489
rect 12574 455 12608 489
rect 12642 455 12676 489
rect 9468 367 9502 401
rect 9468 298 9502 332
rect 4947 210 4981 244
rect 5015 210 5049 244
rect 5083 210 5117 244
rect 5151 210 5185 244
rect 5219 210 5253 244
rect 5287 210 5321 244
rect 5355 210 5389 244
rect 5423 210 5457 244
rect 5491 210 5525 244
rect 5559 210 5593 244
rect 5627 210 5661 244
rect 5695 210 5729 244
rect 5763 210 5797 244
rect 5831 210 5865 244
rect 5899 210 5933 244
rect 5967 210 6001 244
rect 6035 210 6069 244
rect 6103 210 6137 244
rect 6171 210 6205 244
rect 6239 210 6273 244
rect 6307 210 6341 244
rect 6375 210 6409 244
rect 6443 210 6477 244
rect 6511 210 6545 244
rect 6579 210 6613 244
rect 6647 210 6681 244
rect 6715 210 6749 244
rect 6783 210 6817 244
rect 6851 210 6885 244
rect 6919 210 6953 244
rect 6987 210 7021 244
rect 7055 210 7089 244
rect 7123 210 7157 244
rect 7191 210 7225 244
rect 7259 210 7293 244
rect 7327 210 7361 244
rect 7395 210 7429 244
rect 7463 210 7497 244
rect 7531 210 7565 244
rect 7599 210 7633 244
rect 7667 210 7701 244
rect 7735 210 7769 244
rect 7803 210 7837 244
rect 7871 210 7905 244
rect 7939 210 7973 244
rect 8007 210 8041 244
rect 8075 210 8109 244
rect 8143 210 8177 244
rect 8211 210 8245 244
rect 8279 210 8313 244
rect 8347 210 8381 244
rect 8415 210 8449 244
rect 8483 210 8517 244
rect 8551 210 8585 244
rect 8619 210 8653 244
rect 8687 210 8721 244
rect 8755 210 8789 244
rect 8823 210 8857 244
rect 8891 210 8925 244
rect 8959 210 8993 244
rect 9027 210 9061 244
rect 9095 210 9129 244
rect 9163 210 9197 244
rect 9231 210 9265 244
rect 9299 210 9333 244
rect 9367 210 9401 244
rect 9435 210 9469 244
<< mvnsubdiffcont >>
rect 8608 6911 8642 6945
rect 8676 6911 8710 6945
rect 8744 6911 8778 6945
rect 8812 6911 8846 6945
rect 8880 6911 8914 6945
rect 8948 6911 8982 6945
rect 9016 6911 9050 6945
rect 9084 6911 9118 6945
rect 9152 6911 9186 6945
rect 9220 6911 9254 6945
rect 9288 6911 9322 6945
rect 9356 6911 9390 6945
rect 9424 6911 9458 6945
rect 9492 6911 9526 6945
rect 9560 6911 9594 6945
rect 9628 6911 9662 6945
rect 9696 6911 9730 6945
rect 9764 6911 9798 6945
rect 9832 6911 9866 6945
rect 9900 6911 9934 6945
rect 9968 6911 10002 6945
rect 10036 6911 10070 6945
rect 10104 6911 10138 6945
rect 10172 6911 10206 6945
rect 10240 6911 10274 6945
rect 10308 6911 10342 6945
rect 10376 6911 10410 6945
rect 10444 6911 10478 6945
rect 10512 6911 10546 6945
rect 10580 6911 10614 6945
rect 10648 6911 10682 6945
rect 10716 6911 10750 6945
rect 10784 6911 10818 6945
rect 10852 6911 10886 6945
rect 10920 6911 10954 6945
rect 10988 6911 11022 6945
rect 11056 6911 11090 6945
rect 11124 6911 11158 6945
rect 11192 6911 11226 6945
rect 11260 6911 11294 6945
rect 11328 6911 11362 6945
rect 11396 6911 11430 6945
rect 11464 6911 11498 6945
rect 11532 6911 11566 6945
rect 11600 6911 11634 6945
rect 11668 6911 11702 6945
rect 11736 6911 11770 6945
rect 11804 6911 11838 6945
rect 11872 6911 11906 6945
rect 11940 6911 11974 6945
rect 12008 6911 12042 6945
rect 12076 6911 12110 6945
rect 12144 6911 12178 6945
rect 12212 6911 12246 6945
rect 12280 6911 12314 6945
rect 12348 6911 12382 6945
rect 12416 6911 12450 6945
rect 12484 6911 12518 6945
rect 12552 6911 12586 6945
rect 12620 6911 12654 6945
rect 12688 6911 12722 6945
rect 12756 6911 12790 6945
rect 12824 6911 12858 6945
rect 12892 6911 12926 6945
rect 12960 6911 12994 6945
rect 13028 6911 13062 6945
rect 13096 6911 13130 6945
rect 13164 6911 13198 6945
rect 13232 6911 13266 6945
rect 13300 6911 13334 6945
rect 13368 6911 13402 6945
rect 13436 6911 13470 6945
rect 13504 6911 13538 6945
rect 13572 6911 13606 6945
rect 8575 6843 8609 6877
rect 8575 6775 8609 6809
rect 8575 6707 8609 6741
rect 8575 6639 8609 6673
rect 8575 6571 8609 6605
rect 8575 6503 8609 6537
rect 8575 6435 8609 6469
rect 8575 6367 8609 6401
rect 4679 6266 4713 6300
rect 4747 6266 4781 6300
rect 4815 6266 4849 6300
rect 4883 6266 4917 6300
rect 4951 6266 4985 6300
rect 5019 6266 5053 6300
rect 5087 6266 5121 6300
rect 5155 6266 5189 6300
rect 5223 6266 5257 6300
rect 5291 6266 5325 6300
rect 5359 6266 5393 6300
rect 5427 6266 5461 6300
rect 5495 6266 5529 6300
rect 5563 6266 5597 6300
rect 5631 6266 5665 6300
rect 5699 6266 5733 6300
rect 5767 6266 5801 6300
rect 5835 6266 5869 6300
rect 5903 6266 5937 6300
rect 5971 6266 6005 6300
rect 6039 6266 6073 6300
rect 6107 6266 6141 6300
rect 6175 6266 6209 6300
rect 6243 6266 6277 6300
rect 6311 6266 6345 6300
rect 6379 6266 6413 6300
rect 6447 6266 6481 6300
rect 6515 6266 6549 6300
rect 6583 6266 6617 6300
rect 6651 6266 6685 6300
rect 6719 6266 6753 6300
rect 6787 6266 6821 6300
rect 6855 6266 6889 6300
rect 6923 6266 6957 6300
rect 6991 6266 7025 6300
rect 7059 6266 7093 6300
rect 7127 6266 7161 6300
rect 7195 6266 7229 6300
rect 7263 6266 7297 6300
rect 7331 6266 7365 6300
rect 7399 6266 7433 6300
rect 7467 6266 7501 6300
rect 7535 6266 7569 6300
rect 7603 6266 7637 6300
rect 7671 6266 7705 6300
rect 7739 6266 7773 6300
rect 7807 6266 7841 6300
rect 7875 6266 7909 6300
rect 7943 6266 7977 6300
rect 8011 6266 8045 6300
rect 8079 6266 8113 6300
rect 8147 6266 8181 6300
rect 8215 6266 8249 6300
rect 8283 6266 8317 6300
rect 8351 6266 8385 6300
rect 8419 6266 8453 6300
rect 8487 6266 8521 6300
rect 8575 6299 8609 6333
rect 13647 6878 13681 6912
rect 13647 6810 13681 6844
rect 13647 6742 13681 6776
rect 13647 6674 13681 6708
rect 13647 6606 13681 6640
rect 13647 6538 13681 6572
rect 13647 6470 13681 6504
rect 13647 6402 13681 6436
rect 13647 6334 13681 6368
rect 13647 6266 13681 6300
rect 283 6220 317 6254
rect 351 6220 385 6254
rect 419 6220 453 6254
rect 487 6220 521 6254
rect 555 6220 589 6254
rect 623 6220 657 6254
rect 691 6220 725 6254
rect 250 6105 284 6139
rect 778 6187 812 6221
rect 778 6119 812 6153
rect 250 6037 284 6071
rect 250 5969 284 6003
rect 250 5901 284 5935
rect 250 5833 284 5867
rect 250 5765 284 5799
rect 250 5697 284 5731
rect 250 5629 284 5663
rect 250 5561 284 5595
rect 250 5493 284 5527
rect 250 5425 284 5459
rect 778 6051 812 6085
rect 778 5983 812 6017
rect 778 5915 812 5949
rect 778 5847 812 5881
rect 778 5779 812 5813
rect 778 5711 812 5745
rect 778 5643 812 5677
rect 778 5575 812 5609
rect 778 5507 812 5541
rect 250 5357 284 5391
rect 778 5439 812 5473
rect 250 5289 284 5323
rect 250 5221 284 5255
rect 250 5153 284 5187
rect 250 5085 284 5119
rect 778 5371 812 5405
rect 778 5303 812 5337
rect 778 5235 812 5269
rect 778 5167 812 5201
rect 778 5099 812 5133
rect 250 5017 284 5051
rect 250 4949 284 4983
rect 778 5031 812 5065
rect 778 4963 812 4997
rect 250 4881 284 4915
rect 250 4813 284 4847
rect 778 4895 812 4929
rect 778 4827 812 4861
rect 250 4745 284 4779
rect 250 4677 284 4711
rect 250 4609 284 4643
rect 778 4759 812 4793
rect 778 4691 812 4725
rect 250 4541 284 4575
rect 337 4508 371 4542
rect 405 4508 439 4542
rect 473 4508 507 4542
rect 541 4508 575 4542
rect 609 4508 643 4542
rect 677 4508 711 4542
rect 745 4508 779 4542
rect 4646 6187 4680 6221
rect 4646 6119 4680 6153
rect 4646 6051 4680 6085
rect 4646 5983 4680 6017
rect 4646 5915 4680 5949
rect 4646 5847 4680 5881
rect 4646 5779 4680 5813
rect 4646 5711 4680 5745
rect 4646 5643 4680 5677
rect 4646 5575 4680 5609
rect 4646 5507 4680 5541
rect 4646 5439 4680 5473
rect 1702 5129 1736 5163
rect 1770 5129 1804 5163
rect 1838 5129 1872 5163
rect 1906 5129 1940 5163
rect 1974 5129 2008 5163
rect 2042 5129 2076 5163
rect 2110 5129 2144 5163
rect 2178 5129 2212 5163
rect 2246 5129 2280 5163
rect 2314 5129 2348 5163
rect 2382 5129 2416 5163
rect 2450 5129 2484 5163
rect 2518 5129 2552 5163
rect 2586 5129 2620 5163
rect 2654 5129 2688 5163
rect 2722 5129 2756 5163
rect 2790 5129 2824 5163
rect 2858 5129 2892 5163
rect 2926 5129 2960 5163
rect 2994 5129 3028 5163
rect 1669 5060 1703 5094
rect 1669 4992 1703 5026
rect 3079 5096 3113 5130
rect 3079 5028 3113 5062
rect 1669 4924 1703 4958
rect 1669 4856 1703 4890
rect 1669 4788 1703 4822
rect 1669 4720 1703 4754
rect 1669 4652 1703 4686
rect 1669 4584 1703 4618
rect 3079 4960 3113 4994
rect 3079 4892 3113 4926
rect 3079 4824 3113 4858
rect 3079 4756 3113 4790
rect 3079 4688 3113 4722
rect 3079 4620 3113 4654
rect 1669 4516 1703 4550
rect 3079 4552 3113 4586
rect 1669 4448 1703 4482
rect 1669 4380 1703 4414
rect 1669 4312 1703 4346
rect 1669 4244 1703 4278
rect 1669 4176 1703 4210
rect 3079 4484 3113 4518
rect 3079 4416 3113 4450
rect 3079 4348 3113 4382
rect 3079 4280 3113 4314
rect 3079 4212 3113 4246
rect 1669 4108 1703 4142
rect 3079 4144 3113 4178
rect 1669 4040 1703 4074
rect 1669 3972 1703 4006
rect 1669 3904 1703 3938
rect 1669 3836 1703 3870
rect 1669 3768 1703 3802
rect 1669 3700 1703 3734
rect 3079 4076 3113 4110
rect 3079 4008 3113 4042
rect 3079 3940 3113 3974
rect 3079 3872 3113 3906
rect 3079 3804 3113 3838
rect 3079 3736 3113 3770
rect 1669 3632 1703 3666
rect 3079 3668 3113 3702
rect 1669 3564 1703 3598
rect 1669 3496 1703 3530
rect 1669 3428 1703 3462
rect 1669 3360 1703 3394
rect 1669 3292 1703 3326
rect 1669 3224 1703 3258
rect 3079 3600 3113 3634
rect 3079 3532 3113 3566
rect 3079 3464 3113 3498
rect 3079 3396 3113 3430
rect 3079 3328 3113 3362
rect 1669 3156 1703 3190
rect 1669 3088 1703 3122
rect 1669 3020 1703 3054
rect 1669 2952 1703 2986
rect 1669 2884 1703 2918
rect 1669 2816 1703 2850
rect 1669 2748 1703 2782
rect 3079 3260 3113 3294
rect 3079 3192 3113 3226
rect 3079 3124 3113 3158
rect 3079 3056 3113 3090
rect 3079 2988 3113 3022
rect 1669 2680 1703 2714
rect 1669 2612 1703 2646
rect 1669 2544 1703 2578
rect 1669 2476 1703 2510
rect 1669 2408 1703 2442
rect 1669 2340 1703 2374
rect 3079 2920 3113 2954
rect 3079 2852 3113 2886
rect 3079 2784 3113 2818
rect 3079 2716 3113 2750
rect 3079 2648 3113 2682
rect 3079 2580 3113 2614
rect 3079 2512 3113 2546
rect 3079 2444 3113 2478
rect 3079 2376 3113 2410
rect 1669 2272 1703 2306
rect 1669 2204 1703 2238
rect 1669 2136 1703 2170
rect 1669 2068 1703 2102
rect 1669 2000 1703 2034
rect 1669 1932 1703 1966
rect 1669 1864 1703 1898
rect 3079 2308 3113 2342
rect 3079 2240 3113 2274
rect 3079 2172 3113 2206
rect 3079 2104 3113 2138
rect 3079 2036 3113 2070
rect 3079 1968 3113 2002
rect 1669 1796 1703 1830
rect 3079 1900 3113 1934
rect 1669 1728 1703 1762
rect 1669 1660 1703 1694
rect 1669 1592 1703 1626
rect 1669 1524 1703 1558
rect 1669 1456 1703 1490
rect 1669 1388 1703 1422
rect 3079 1832 3113 1866
rect 3079 1764 3113 1798
rect 3079 1696 3113 1730
rect 3079 1628 3113 1662
rect 3079 1560 3113 1594
rect 3079 1492 3113 1526
rect 1669 1320 1703 1354
rect 3079 1424 3113 1458
rect 1669 1252 1703 1286
rect 1669 1184 1703 1218
rect 1669 1116 1703 1150
rect 1669 1048 1703 1082
rect 1669 980 1703 1014
rect 3079 1356 3113 1390
rect 3079 1288 3113 1322
rect 3079 1220 3113 1254
rect 3079 1152 3113 1186
rect 3079 1084 3113 1118
rect 3079 1016 3113 1050
rect 1669 912 1703 946
rect 3079 948 3113 982
rect 1669 844 1703 878
rect 1669 776 1703 810
rect 1669 708 1703 742
rect 1669 640 1703 674
rect 1669 572 1703 606
rect 1669 504 1703 538
rect 3079 880 3113 914
rect 3079 812 3113 846
rect 3079 744 3113 778
rect 3079 676 3113 710
rect 3079 608 3113 642
rect 3079 540 3113 574
rect 1669 436 1703 470
rect 1669 368 1703 402
rect 3079 472 3113 506
rect 1754 335 1788 369
rect 1822 335 1856 369
rect 1890 335 1924 369
rect 1958 335 1992 369
rect 2026 335 2060 369
rect 2094 335 2128 369
rect 2162 335 2196 369
rect 2230 335 2264 369
rect 2298 335 2332 369
rect 2366 335 2400 369
rect 2434 335 2468 369
rect 2502 335 2536 369
rect 2570 335 2604 369
rect 2638 335 2672 369
rect 2706 335 2740 369
rect 2774 335 2808 369
rect 2842 335 2876 369
rect 2910 335 2944 369
rect 2978 335 3012 369
rect 3046 335 3080 369
rect 4646 5371 4680 5405
rect 4646 5303 4680 5337
rect 4646 5235 4680 5269
rect 4646 5167 4680 5201
rect 4646 5099 4680 5133
rect 13647 6198 13681 6232
rect 13647 6130 13681 6164
rect 13647 6062 13681 6096
rect 13647 5994 13681 6028
rect 13647 5926 13681 5960
rect 13647 5858 13681 5892
rect 13647 5790 13681 5824
rect 13647 5722 13681 5756
rect 13647 5654 13681 5688
rect 13647 5586 13681 5620
rect 13647 5518 13681 5552
rect 13647 5450 13681 5484
rect 13647 5382 13681 5416
rect 13647 5314 13681 5348
rect 13647 5246 13681 5280
rect 13647 5178 13681 5212
rect 4646 5031 4680 5065
rect 4646 4963 4680 4997
rect 4646 4895 4680 4929
rect 4646 4827 4680 4861
rect 4646 4759 4680 4793
rect 4646 4691 4680 4725
rect 4646 4623 4680 4657
rect 4646 4555 4680 4589
rect 4646 4487 4680 4521
rect 4646 4419 4680 4453
rect 4646 4351 4680 4385
rect 4646 4283 4680 4317
rect 4646 4215 4680 4249
rect 4646 4147 4680 4181
rect 4646 4079 4680 4113
rect 4646 4011 4680 4045
rect 4646 3943 4680 3977
rect 4646 3875 4680 3909
rect 4646 3807 4680 3841
rect 4646 3739 4680 3773
rect 4646 3671 4680 3705
rect 4646 3603 4680 3637
rect 4646 3535 4680 3569
rect 4646 3467 4680 3501
rect 4646 3399 4680 3433
rect 4646 3331 4680 3365
rect 4646 3263 4680 3297
rect 4646 3195 4680 3229
rect 4646 3127 4680 3161
rect 4646 3059 4680 3093
rect 4646 2991 4680 3025
rect 4646 2923 4680 2957
rect 4646 2855 4680 2889
rect 4646 2787 4680 2821
rect 4646 2719 4680 2753
rect 4646 2651 4680 2685
rect 4646 2583 4680 2617
rect 4646 2515 4680 2549
rect 4646 2447 4680 2481
rect 4646 2379 4680 2413
rect 4646 2311 4680 2345
rect 4646 2243 4680 2277
rect 4646 2175 4680 2209
rect 4646 2107 4680 2141
rect 4646 2039 4680 2073
rect 4646 1971 4680 2005
rect 4646 1903 4680 1937
rect 4646 1835 4680 1869
rect 4646 1767 4680 1801
rect 4646 1699 4680 1733
rect 4646 1631 4680 1665
rect 4646 1563 4680 1597
rect 4646 1495 4680 1529
rect 4646 1427 4680 1461
rect 4646 1359 4680 1393
rect 4646 1291 4680 1325
rect 4646 1223 4680 1257
rect 4646 1155 4680 1189
rect 4646 1087 4680 1121
rect 4646 1019 4680 1053
rect 4646 951 4680 985
rect 4646 883 4680 917
rect 4646 815 4680 849
rect 4646 747 4680 781
rect 4646 679 4680 713
rect 4646 611 4680 645
rect 4646 543 4680 577
rect 4646 475 4680 509
rect 4646 407 4680 441
rect 4646 339 4680 373
rect 4646 271 4680 305
rect 4646 203 4680 237
rect 12946 5012 12980 5046
rect 13070 5045 13104 5079
rect 13138 5045 13172 5079
rect 13206 5045 13240 5079
rect 13274 5045 13308 5079
rect 13342 5045 13376 5079
rect 13410 5045 13444 5079
rect 13478 5045 13512 5079
rect 13546 5045 13580 5079
rect 13614 5045 13648 5079
rect 12946 4944 12980 4978
rect 12946 4876 12980 4910
rect 12946 4808 12980 4842
rect 12946 4740 12980 4774
rect 12946 4672 12980 4706
rect 12946 4604 12980 4638
rect 12946 4536 12980 4570
rect 12946 4468 12980 4502
rect 12946 4400 12980 4434
rect 12946 4332 12980 4366
rect 12946 4264 12980 4298
rect 12946 4196 12980 4230
rect 12946 4128 12980 4162
rect 12946 4060 12980 4094
rect 12946 3992 12980 4026
rect 12946 3924 12980 3958
rect 12946 3856 12980 3890
rect 12946 3788 12980 3822
rect 12946 3720 12980 3754
rect 12946 3652 12980 3686
rect 12946 3584 12980 3618
rect 12946 3516 12980 3550
rect 12946 3448 12980 3482
rect 12946 3380 12980 3414
rect 12946 3312 12980 3346
rect 12946 3244 12980 3278
rect 12946 3176 12980 3210
rect 12946 3108 12980 3142
rect 12946 3040 12980 3074
rect 12946 2972 12980 3006
rect 12946 2904 12980 2938
rect 12946 2836 12980 2870
rect 12946 2768 12980 2802
rect 12946 2700 12980 2734
rect 12946 2632 12980 2666
rect 12946 2564 12980 2598
rect 12946 2496 12980 2530
rect 12946 2428 12980 2462
rect 12946 2360 12980 2394
rect 12946 2292 12980 2326
rect 12946 2224 12980 2258
rect 12946 2156 12980 2190
rect 12946 2088 12980 2122
rect 12946 2020 12980 2054
rect 12946 1952 12980 1986
rect 12946 1884 12980 1918
rect 12946 1816 12980 1850
rect 12946 1748 12980 1782
rect 12946 1680 12980 1714
rect 12946 1612 12980 1646
rect 12946 1544 12980 1578
rect 12946 1476 12980 1510
rect 12946 1408 12980 1442
rect 12946 1340 12980 1374
rect 12946 1272 12980 1306
rect 12946 1204 12980 1238
rect 12946 1136 12980 1170
rect 12946 1068 12980 1102
rect 12946 1000 12980 1034
rect 12946 932 12980 966
rect 12946 864 12980 898
rect 12946 796 12980 830
rect 12946 728 12980 762
rect 12946 660 12980 694
rect 12946 592 12980 626
rect 12946 524 12980 558
rect 12946 456 12980 490
rect 12946 388 12980 422
rect 12946 320 12980 354
rect 12946 252 12980 286
rect 4646 135 4680 169
rect 4646 67 4680 101
rect 4646 -1 4680 33
rect 12946 184 12980 218
rect 12946 116 12980 150
rect 12946 48 12980 82
rect 4646 -69 4680 -35
rect 4646 -137 4680 -103
rect 12946 -20 12980 14
rect 12946 -88 12980 -54
rect 4646 -205 4680 -171
rect 4646 -273 4680 -239
rect 4646 -341 4680 -307
rect 4646 -409 4680 -375
rect 12946 -257 12980 -223
rect 12946 -325 12980 -291
rect 4753 -442 4787 -408
rect 4821 -442 4855 -408
rect 4889 -442 4923 -408
rect 4957 -442 4991 -408
rect 5025 -442 5059 -408
rect 5093 -442 5127 -408
rect 5161 -442 5195 -408
rect 5229 -442 5263 -408
rect 5297 -442 5331 -408
rect 5365 -442 5399 -408
rect 5433 -442 5467 -408
rect 5501 -442 5535 -408
rect 5569 -442 5603 -408
rect 5637 -442 5671 -408
rect 5705 -442 5739 -408
rect 5773 -442 5807 -408
rect 5841 -442 5875 -408
rect 5909 -442 5943 -408
rect 5977 -442 6011 -408
rect 6045 -442 6079 -408
rect 6113 -442 6147 -408
rect 6181 -442 6215 -408
rect 6249 -442 6283 -408
rect 6317 -442 6351 -408
rect 6385 -442 6419 -408
rect 6453 -442 6487 -408
rect 6521 -442 6555 -408
rect 6589 -442 6623 -408
rect 6657 -442 6691 -408
rect 6725 -442 6759 -408
rect 6793 -442 6827 -408
rect 6861 -442 6895 -408
rect 6929 -442 6963 -408
rect 6997 -442 7031 -408
rect 7065 -442 7099 -408
rect 7133 -442 7167 -408
rect 7201 -442 7235 -408
rect 7269 -442 7303 -408
rect 7337 -442 7371 -408
rect 7405 -442 7439 -408
rect 7473 -442 7507 -408
rect 7541 -442 7575 -408
rect 7609 -442 7643 -408
rect 7677 -442 7711 -408
rect 7745 -442 7779 -408
rect 7813 -442 7847 -408
rect 7881 -442 7915 -408
rect 7949 -442 7983 -408
rect 8017 -442 8051 -408
rect 8085 -442 8119 -408
rect 8153 -442 8187 -408
rect 8221 -442 8255 -408
rect 8289 -442 8323 -408
rect 8357 -442 8391 -408
rect 8425 -442 8459 -408
rect 8493 -442 8527 -408
rect 8561 -442 8595 -408
rect 8629 -442 8663 -408
rect 8697 -442 8731 -408
rect 8765 -442 8799 -408
rect 8833 -442 8867 -408
rect 8901 -442 8935 -408
rect 8969 -442 9003 -408
rect 9037 -442 9071 -408
rect 9105 -442 9139 -408
rect 9173 -442 9207 -408
rect 9241 -442 9275 -408
rect 9309 -442 9343 -408
rect 9377 -442 9411 -408
rect 9445 -442 9479 -408
rect 9513 -442 9547 -408
rect 9581 -442 9615 -408
rect 9649 -442 9683 -408
rect 9717 -442 9751 -408
rect 9785 -442 9819 -408
rect 9853 -442 9887 -408
rect 9921 -442 9955 -408
rect 9989 -442 10023 -408
rect 10057 -442 10091 -408
rect 10125 -442 10159 -408
rect 10193 -442 10227 -408
rect 10261 -442 10295 -408
rect 10329 -442 10363 -408
rect 10397 -442 10431 -408
rect 10465 -442 10499 -408
rect 10533 -442 10567 -408
rect 10601 -442 10635 -408
rect 10669 -442 10703 -408
rect 10737 -442 10771 -408
rect 10805 -442 10839 -408
rect 10873 -442 10907 -408
rect 10941 -442 10975 -408
rect 11009 -442 11043 -408
rect 11077 -442 11111 -408
rect 11145 -442 11179 -408
rect 11213 -442 11247 -408
rect 11281 -442 11315 -408
rect 11349 -442 11383 -408
rect 11417 -442 11451 -408
rect 11485 -442 11519 -408
rect 11553 -442 11587 -408
rect 11621 -442 11655 -408
rect 11689 -442 11723 -408
rect 11757 -442 11791 -408
rect 11825 -442 11859 -408
rect 11893 -442 11927 -408
rect 11961 -442 11995 -408
rect 12029 -442 12063 -408
rect 12097 -442 12131 -408
rect 12165 -442 12199 -408
rect 12233 -442 12267 -408
rect 12301 -442 12335 -408
rect 12369 -442 12403 -408
rect 12437 -442 12471 -408
rect 12505 -442 12539 -408
rect 12573 -442 12607 -408
rect 12641 -442 12675 -408
rect 12709 -442 12743 -408
rect 12777 -442 12811 -408
rect 12845 -442 12879 -408
rect 12913 -442 12947 -408
<< poly >>
rect 10205 11328 11861 11344
rect 10205 11294 10221 11328
rect 10255 11294 10291 11328
rect 10325 11294 10361 11328
rect 10395 11294 10431 11328
rect 10465 11294 10500 11328
rect 10534 11294 10569 11328
rect 10603 11294 10638 11328
rect 10672 11294 10707 11328
rect 10741 11294 10776 11328
rect 10810 11294 10845 11328
rect 10879 11294 10914 11328
rect 10948 11294 10983 11328
rect 11017 11294 11052 11328
rect 11086 11294 11121 11328
rect 11155 11294 11190 11328
rect 11224 11294 11259 11328
rect 11293 11294 11328 11328
rect 11362 11294 11397 11328
rect 11431 11294 11466 11328
rect 11500 11294 11535 11328
rect 11569 11294 11604 11328
rect 11638 11294 11673 11328
rect 11707 11294 11742 11328
rect 11776 11294 11811 11328
rect 11845 11294 11861 11328
rect 10205 11278 11861 11294
rect 6488 10437 11568 10453
rect 6488 10403 6504 10437
rect 6538 10403 6573 10437
rect 6607 10403 6642 10437
rect 6676 10403 6711 10437
rect 6745 10403 6780 10437
rect 6814 10403 6849 10437
rect 6883 10403 6918 10437
rect 6952 10403 6987 10437
rect 7021 10403 7056 10437
rect 7090 10403 7125 10437
rect 7159 10403 7194 10437
rect 7228 10403 7263 10437
rect 7297 10403 7332 10437
rect 7366 10403 7401 10437
rect 7435 10403 7470 10437
rect 7504 10403 7539 10437
rect 7573 10403 7608 10437
rect 7642 10403 7677 10437
rect 7711 10403 7746 10437
rect 7780 10403 7815 10437
rect 7849 10403 7884 10437
rect 7918 10403 7953 10437
rect 7987 10403 8022 10437
rect 8056 10403 8091 10437
rect 8125 10403 8160 10437
rect 8194 10403 8229 10437
rect 8263 10403 8298 10437
rect 8332 10403 8367 10437
rect 8401 10403 8436 10437
rect 8470 10403 8505 10437
rect 8539 10403 8574 10437
rect 8608 10403 8643 10437
rect 8677 10403 8712 10437
rect 8746 10403 8781 10437
rect 8815 10403 8850 10437
rect 8884 10403 8919 10437
rect 8953 10403 8988 10437
rect 9022 10403 9057 10437
rect 9091 10403 9126 10437
rect 9160 10403 9195 10437
rect 9229 10403 9264 10437
rect 9298 10403 9333 10437
rect 9367 10403 9402 10437
rect 9436 10403 9471 10437
rect 9505 10403 9540 10437
rect 9574 10403 9609 10437
rect 9643 10403 9678 10437
rect 9712 10403 9747 10437
rect 9781 10403 9816 10437
rect 9850 10403 9885 10437
rect 9919 10403 9954 10437
rect 9988 10403 10022 10437
rect 10056 10403 10090 10437
rect 10124 10403 10158 10437
rect 10192 10403 10226 10437
rect 10260 10403 10294 10437
rect 10328 10403 10362 10437
rect 10396 10403 10430 10437
rect 10464 10403 10498 10437
rect 10532 10403 10566 10437
rect 10600 10403 10634 10437
rect 10668 10403 10702 10437
rect 10736 10403 10770 10437
rect 10804 10403 10838 10437
rect 10872 10403 10906 10437
rect 10940 10403 10974 10437
rect 11008 10403 11042 10437
rect 11076 10403 11110 10437
rect 11144 10403 11178 10437
rect 11212 10403 11246 10437
rect 11280 10403 11314 10437
rect 11348 10403 11382 10437
rect 11416 10403 11450 10437
rect 11484 10403 11518 10437
rect 11552 10403 11568 10437
rect 6488 10387 11568 10403
rect 6487 9553 9856 9576
rect 6487 9519 6504 9553
rect 6538 9519 6573 9553
rect 6607 9519 6642 9553
rect 6676 9519 6711 9553
rect 6745 9519 6780 9553
rect 6814 9519 6849 9553
rect 6883 9519 6918 9553
rect 6952 9519 6987 9553
rect 7021 9519 7056 9553
rect 7090 9519 7125 9553
rect 7159 9519 7194 9553
rect 7228 9519 7263 9553
rect 7297 9519 7332 9553
rect 7366 9519 7401 9553
rect 7435 9519 7470 9553
rect 7504 9519 7539 9553
rect 7573 9519 7608 9553
rect 7642 9519 7677 9553
rect 7711 9519 7746 9553
rect 7780 9519 7815 9553
rect 7849 9519 7884 9553
rect 7918 9519 7953 9553
rect 7987 9519 8022 9553
rect 8056 9519 8091 9553
rect 8125 9519 8160 9553
rect 8194 9519 8229 9553
rect 8263 9519 8298 9553
rect 8332 9519 8367 9553
rect 8401 9519 8436 9553
rect 8470 9519 8505 9553
rect 8539 9519 8574 9553
rect 8608 9519 8643 9553
rect 8677 9519 8712 9553
rect 8746 9519 8781 9553
rect 8815 9519 8850 9553
rect 8884 9519 8918 9553
rect 8952 9519 8986 9553
rect 9020 9519 9054 9553
rect 9088 9519 9122 9553
rect 9156 9519 9190 9553
rect 9224 9519 9258 9553
rect 9292 9519 9326 9553
rect 9360 9519 9394 9553
rect 9428 9519 9462 9553
rect 9496 9519 9530 9553
rect 9564 9519 9598 9553
rect 9632 9519 9666 9553
rect 9700 9519 9734 9553
rect 9768 9519 9802 9553
rect 9836 9519 9856 9553
rect 6487 9498 9856 9519
rect 659 6076 743 6092
rect 659 6042 693 6076
rect 727 6042 743 6076
rect 659 6004 743 6042
rect 659 5972 693 6004
rect 677 5970 693 5972
rect 727 5970 743 6004
rect 677 5932 743 5970
rect 677 5916 693 5932
rect 659 5898 693 5916
rect 727 5898 743 5932
rect 659 5859 743 5898
rect 659 5825 693 5859
rect 727 5825 743 5859
rect 659 5796 743 5825
rect 677 5786 743 5796
rect 677 5752 693 5786
rect 727 5752 743 5786
rect 677 5740 743 5752
rect 659 5713 743 5740
rect 659 5679 693 5713
rect 727 5679 743 5713
rect 659 5640 743 5679
rect 659 5620 693 5640
rect 677 5606 693 5620
rect 727 5606 743 5640
rect 677 5567 743 5606
rect 677 5564 693 5567
rect 659 5533 693 5564
rect 727 5533 743 5567
rect 659 5494 743 5533
rect 659 5460 693 5494
rect 727 5460 743 5494
rect 659 5444 743 5460
rect 319 5372 407 5388
rect 319 5338 335 5372
rect 369 5338 407 5372
rect 319 5295 407 5338
rect 319 5261 335 5295
rect 369 5268 407 5295
rect 369 5261 385 5268
rect 319 5218 385 5261
rect 319 5184 335 5218
rect 369 5212 385 5218
rect 369 5184 407 5212
rect 319 5142 407 5184
rect 319 5108 335 5142
rect 369 5108 407 5142
rect 319 5092 407 5108
rect 609 4910 743 4926
rect 609 4876 693 4910
rect 727 4876 743 4910
rect 609 4842 743 4876
rect 609 4826 693 4842
rect 677 4808 693 4826
rect 727 4808 743 4842
rect 677 4792 743 4808
rect 319 4754 407 4770
rect 319 4720 335 4754
rect 369 4720 407 4754
rect 319 4686 407 4720
rect 319 4652 335 4686
rect 369 4670 407 4686
rect 369 4652 385 4670
rect 319 4636 385 4652
rect 1036 6076 1113 6092
rect 1036 6042 1052 6076
rect 1086 6042 1113 6076
rect 1036 5999 1113 6042
rect 1036 5965 1052 5999
rect 1086 5972 1113 5999
rect 1086 5965 1102 5972
rect 1036 5922 1102 5965
rect 1036 5888 1052 5922
rect 1086 5916 1102 5922
rect 1086 5888 1113 5916
rect 1036 5846 1113 5888
rect 1036 5812 1052 5846
rect 1086 5812 1113 5846
rect 1036 5796 1113 5812
rect 1036 5724 1113 5740
rect 1036 5690 1052 5724
rect 1086 5690 1113 5724
rect 1036 5656 1113 5690
rect 1036 5622 1052 5656
rect 1086 5622 1113 5656
rect 1036 5620 1113 5622
rect 1036 5606 1102 5620
rect 1073 5438 1163 5454
rect 1073 5404 1089 5438
rect 1123 5404 1163 5438
rect 1073 5304 1163 5404
rect 1073 5270 1089 5304
rect 1123 5270 1163 5304
rect 1073 5254 1163 5270
rect 1042 5182 1163 5198
rect 1042 5148 1058 5182
rect 1092 5148 1163 5182
rect 1042 5048 1163 5148
rect 1042 5014 1058 5048
rect 1092 5014 1163 5048
rect 1042 4998 1163 5014
rect 335 4133 407 4149
rect 335 4099 351 4133
rect 385 4099 407 4133
rect 335 4051 407 4099
rect 335 4017 351 4051
rect 385 4029 407 4051
rect 385 4017 401 4029
rect 335 3973 401 4017
rect 335 3970 407 3973
rect 335 3936 351 3970
rect 385 3936 407 3970
rect 335 3889 407 3936
rect 335 3855 351 3889
rect 385 3855 407 3889
rect 335 3853 407 3855
rect 335 3808 401 3853
rect 335 3774 351 3808
rect 385 3797 401 3808
rect 385 3774 407 3797
rect 335 3727 407 3774
rect 335 3693 351 3727
rect 385 3693 407 3727
rect 335 3677 407 3693
rect 1036 4816 1110 4832
rect 1036 4782 1052 4816
rect 1086 4782 1110 4816
rect 1036 4747 1110 4782
rect 1036 4713 1052 4747
rect 1086 4713 1110 4747
rect 1036 4678 1110 4713
rect 1036 4644 1052 4678
rect 1086 4652 1110 4678
rect 1086 4644 1102 4652
rect 1036 4609 1102 4644
rect 1036 4575 1052 4609
rect 1086 4596 1102 4609
rect 1086 4575 1110 4596
rect 1036 4540 1110 4575
rect 1036 4506 1052 4540
rect 1086 4506 1110 4540
rect 1036 4471 1110 4506
rect 1036 4437 1052 4471
rect 1086 4437 1110 4471
rect 1036 4416 1110 4437
rect 1036 4402 1102 4416
rect 1036 4368 1052 4402
rect 1086 4368 1102 4402
rect 1036 4360 1102 4368
rect 1036 4334 1110 4360
rect 1036 4300 1052 4334
rect 1086 4300 1110 4334
rect 1036 4266 1110 4300
rect 1036 4232 1052 4266
rect 1086 4232 1110 4266
rect 1036 4198 1110 4232
rect 1036 4164 1052 4198
rect 1086 4180 1110 4198
rect 1086 4164 1102 4180
rect 1036 4130 1102 4164
rect 1036 4096 1052 4130
rect 1086 4124 1102 4130
rect 1086 4096 1110 4124
rect 1036 4062 1110 4096
rect 1036 4028 1052 4062
rect 1086 4028 1110 4062
rect 1036 3994 1110 4028
rect 1036 3960 1052 3994
rect 1086 3960 1110 3994
rect 1036 3944 1110 3960
rect 1036 3738 1113 3754
rect 1036 3704 1052 3738
rect 1086 3724 1113 3738
rect 1086 3704 1102 3724
rect 1036 3668 1102 3704
rect 1036 3664 1113 3668
rect 1036 3630 1052 3664
rect 1086 3638 1113 3664
rect 1086 3630 1102 3638
rect 1036 3590 1102 3630
rect 1036 3556 1052 3590
rect 1086 3582 1102 3590
rect 1086 3556 1113 3582
rect 1036 3552 1113 3556
rect 1036 3516 1102 3552
rect 1036 3482 1052 3516
rect 1086 3496 1102 3516
rect 1086 3482 1113 3496
rect 1036 3466 1113 3482
rect 333 3182 419 3198
rect 333 3148 349 3182
rect 383 3162 419 3182
rect 383 3148 399 3162
rect 333 3114 399 3148
rect 333 3080 349 3114
rect 383 3080 399 3114
rect 333 3064 399 3080
rect 677 3078 743 3094
rect 677 3044 693 3078
rect 727 3044 743 3078
rect 677 3010 743 3044
rect 677 2996 693 3010
rect 671 2976 693 2996
rect 727 2976 743 3010
rect 671 2960 743 2976
rect 319 2888 419 2904
rect 319 2854 335 2888
rect 369 2868 419 2888
rect 369 2854 385 2868
rect 319 2812 385 2854
rect 319 2811 419 2812
rect 319 2777 335 2811
rect 369 2777 419 2811
rect 319 2776 419 2777
rect 319 2734 385 2776
rect 319 2700 335 2734
rect 369 2720 385 2734
rect 369 2700 419 2720
rect 319 2684 419 2700
rect 677 2536 743 2552
rect 677 2518 693 2536
rect 671 2502 693 2518
rect 727 2502 743 2536
rect 671 2468 743 2502
rect 671 2434 693 2468
rect 727 2434 743 2468
rect 671 2418 743 2434
rect 347 2346 419 2362
rect 347 2312 363 2346
rect 397 2312 419 2346
rect 347 2278 419 2312
rect 347 2244 363 2278
rect 397 2262 419 2278
rect 397 2244 413 2262
rect 347 2228 413 2244
rect 1036 3336 1102 3352
rect 1036 3302 1052 3336
rect 1086 3302 1102 3336
rect 1036 3268 1102 3302
rect 1036 3234 1052 3268
rect 1086 3254 1102 3268
rect 1086 3234 1110 3254
rect 1036 3218 1110 3234
rect 1362 3146 1436 3162
rect 1362 3126 1386 3146
rect 1370 3112 1386 3126
rect 1420 3112 1436 3146
rect 1370 3078 1436 3112
rect 1036 3042 1102 3058
rect 1036 3008 1052 3042
rect 1086 3008 1102 3042
rect 1370 3044 1386 3078
rect 1420 3044 1436 3078
rect 1370 3028 1436 3044
rect 1036 2974 1102 3008
rect 1036 2940 1052 2974
rect 1086 2960 1102 2974
rect 1086 2940 1110 2960
rect 1036 2924 1110 2940
rect 1362 2742 1436 2758
rect 1362 2722 1386 2742
rect 1370 2708 1386 2722
rect 1420 2708 1436 2742
rect 1370 2666 1436 2708
rect 1362 2665 1436 2666
rect 1362 2631 1386 2665
rect 1420 2631 1436 2665
rect 1362 2630 1436 2631
rect 1370 2588 1436 2630
rect 1370 2574 1386 2588
rect 1362 2554 1386 2574
rect 1420 2554 1436 2588
rect 1362 2538 1436 2554
rect 1362 2466 1436 2482
rect 1362 2446 1386 2466
rect 1370 2432 1386 2446
rect 1420 2432 1436 2466
rect 1370 2390 1436 2432
rect 1362 2389 1436 2390
rect 1362 2355 1386 2389
rect 1420 2355 1436 2389
rect 1362 2354 1436 2355
rect 1370 2312 1436 2354
rect 1370 2298 1386 2312
rect 1362 2278 1386 2298
rect 1420 2278 1436 2312
rect 1362 2262 1436 2278
rect 1036 2190 1110 2206
rect 1036 2156 1052 2190
rect 1086 2170 1110 2190
rect 1086 2156 1102 2170
rect 1036 2122 1102 2156
rect 1036 2088 1052 2122
rect 1086 2088 1102 2122
rect 1036 2072 1102 2088
rect 333 1767 407 1783
rect 333 1733 349 1767
rect 383 1733 407 1767
rect 333 1685 407 1733
rect 333 1651 349 1685
rect 383 1651 407 1685
rect 333 1604 407 1651
rect 333 1570 349 1604
rect 383 1570 407 1604
rect 333 1523 407 1570
rect 333 1489 349 1523
rect 383 1489 407 1523
rect 333 1442 407 1489
rect 333 1408 349 1442
rect 383 1408 407 1442
rect 333 1361 407 1408
rect 333 1327 349 1361
rect 383 1327 407 1361
rect 333 1311 407 1327
rect 333 1129 407 1145
rect 333 1095 349 1129
rect 383 1095 407 1129
rect 333 1056 407 1095
rect 333 1022 349 1056
rect 383 1022 407 1056
rect 333 983 407 1022
rect 333 949 349 983
rect 383 949 407 983
rect 333 910 407 949
rect 333 876 349 910
rect 383 876 407 910
rect 333 837 407 876
rect 333 803 349 837
rect 383 803 407 837
rect 333 764 407 803
rect 333 730 349 764
rect 383 730 407 764
rect 333 691 407 730
rect 333 657 349 691
rect 383 657 407 691
rect 333 619 407 657
rect 333 585 349 619
rect 383 585 407 619
rect 333 547 407 585
rect 333 513 349 547
rect 383 513 407 547
rect 333 497 407 513
rect 1036 1847 1113 1863
rect 1036 1813 1052 1847
rect 1086 1833 1113 1847
rect 1086 1813 1102 1833
rect 1036 1777 1102 1813
rect 1036 1773 1113 1777
rect 1036 1739 1052 1773
rect 1086 1747 1113 1773
rect 1086 1739 1102 1747
rect 1036 1699 1102 1739
rect 1036 1665 1052 1699
rect 1086 1691 1102 1699
rect 1086 1665 1113 1691
rect 1036 1661 1113 1665
rect 1036 1625 1102 1661
rect 1036 1591 1052 1625
rect 1086 1605 1102 1625
rect 1086 1591 1113 1605
rect 1036 1575 1113 1591
rect 1036 1369 1110 1385
rect 1036 1335 1052 1369
rect 1086 1335 1110 1369
rect 1036 1300 1110 1335
rect 1036 1266 1052 1300
rect 1086 1266 1110 1300
rect 1036 1231 1110 1266
rect 1036 1197 1052 1231
rect 1086 1205 1110 1231
rect 1086 1197 1102 1205
rect 1036 1162 1102 1197
rect 1036 1128 1052 1162
rect 1086 1149 1102 1162
rect 1086 1128 1110 1149
rect 1036 1093 1110 1128
rect 1036 1059 1052 1093
rect 1086 1059 1110 1093
rect 1036 1024 1110 1059
rect 1036 990 1052 1024
rect 1086 990 1110 1024
rect 1036 969 1110 990
rect 1036 955 1102 969
rect 1036 921 1052 955
rect 1086 921 1102 955
rect 1036 913 1102 921
rect 1036 887 1110 913
rect 1036 853 1052 887
rect 1086 853 1110 887
rect 1036 819 1110 853
rect 1036 785 1052 819
rect 1086 785 1110 819
rect 1036 751 1110 785
rect 1036 717 1052 751
rect 1086 733 1110 751
rect 1086 717 1102 733
rect 1036 683 1102 717
rect 1036 649 1052 683
rect 1086 677 1102 683
rect 1086 649 1110 677
rect 1036 615 1110 649
rect 1036 581 1052 615
rect 1086 581 1110 615
rect 1036 547 1110 581
rect 1036 513 1052 547
rect 1086 513 1110 547
rect 1036 497 1110 513
rect 1738 4985 1810 5001
rect 1738 4951 1754 4985
rect 1788 4951 1810 4985
rect 1738 4902 1810 4951
rect 1738 4868 1754 4902
rect 1788 4868 1810 4902
rect 1738 4819 1810 4868
rect 1738 4785 1754 4819
rect 1788 4785 1810 4819
rect 1738 4735 1810 4785
rect 1738 4701 1754 4735
rect 1788 4701 1810 4735
rect 1738 4651 1810 4701
rect 1738 4617 1754 4651
rect 1788 4617 1810 4651
rect 1738 4601 1810 4617
rect 2462 4985 2534 5001
rect 2462 4951 2484 4985
rect 2518 4971 2534 4985
rect 2518 4951 2540 4971
rect 2462 4902 2540 4951
rect 2462 4868 2484 4902
rect 2518 4868 2540 4902
rect 2462 4819 2540 4868
rect 2462 4785 2484 4819
rect 2518 4785 2540 4819
rect 2462 4735 2540 4785
rect 2462 4701 2484 4735
rect 2518 4701 2540 4735
rect 2462 4651 2540 4701
rect 2462 4617 2484 4651
rect 2518 4617 2540 4651
rect 2462 4601 2540 4617
rect 2534 4571 2540 4601
rect 1738 4529 1810 4545
rect 1738 4495 1754 4529
rect 1788 4495 1810 4529
rect 1738 4446 1810 4495
rect 1738 4412 1754 4446
rect 1788 4412 1810 4446
rect 1738 4363 1810 4412
rect 1738 4329 1754 4363
rect 1788 4329 1810 4363
rect 1738 4279 1810 4329
rect 1738 4245 1754 4279
rect 1788 4245 1810 4279
rect 1738 4195 1810 4245
rect 1738 4161 1754 4195
rect 1788 4161 1810 4195
rect 1738 4145 1810 4161
rect 2462 4359 2468 4545
rect 2892 4482 3032 4515
rect 2892 4448 2914 4482
rect 2948 4448 2982 4482
rect 3016 4448 3032 4482
rect 2892 4415 3032 4448
rect 2462 4343 2540 4359
rect 2462 4309 2484 4343
rect 2518 4309 2540 4343
rect 2462 4272 2540 4309
rect 2462 4238 2484 4272
rect 2518 4259 2540 4272
rect 2518 4238 2534 4259
rect 2462 4203 2534 4238
rect 2462 4201 2540 4203
rect 2462 4167 2484 4201
rect 2518 4167 2540 4201
rect 2462 4145 2540 4167
rect 2468 4130 2540 4145
rect 2468 4096 2484 4130
rect 2518 4103 2540 4130
rect 2518 4096 2534 4103
rect 2468 4089 2534 4096
rect 1738 4073 1810 4089
rect 1738 4039 1754 4073
rect 1788 4039 1810 4073
rect 1738 3990 1810 4039
rect 1738 3956 1754 3990
rect 1788 3956 1810 3990
rect 1738 3907 1810 3956
rect 1738 3873 1754 3907
rect 1788 3873 1810 3907
rect 1738 3823 1810 3873
rect 1738 3789 1754 3823
rect 1788 3789 1810 3823
rect 1738 3739 1810 3789
rect 1738 3705 1754 3739
rect 1788 3705 1810 3739
rect 1738 3689 1810 3705
rect 2462 4059 2534 4089
rect 2462 4025 2484 4059
rect 2518 4047 2534 4059
rect 2518 4025 2540 4047
rect 2462 3988 2540 4025
rect 2462 3954 2484 3988
rect 2518 3954 2540 3988
rect 2462 3947 2540 3954
rect 2462 3917 2534 3947
rect 2462 3883 2484 3917
rect 2518 3891 2534 3917
rect 2518 3883 2540 3891
rect 2462 3845 2540 3883
rect 2462 3811 2484 3845
rect 2518 3811 2540 3845
rect 2462 3791 2540 3811
rect 2462 3773 2534 3791
rect 2462 3739 2484 3773
rect 2518 3739 2534 3773
rect 2462 3735 2534 3739
rect 2462 3701 2540 3735
rect 2462 3689 2484 3701
rect 2468 3667 2484 3689
rect 2518 3667 2540 3701
rect 2468 3635 2540 3667
rect 2468 3633 2534 3635
rect 1738 3617 1810 3633
rect 1738 3583 1754 3617
rect 1788 3583 1810 3617
rect 1738 3534 1810 3583
rect 1738 3500 1754 3534
rect 1788 3500 1810 3534
rect 1738 3451 1810 3500
rect 1738 3417 1754 3451
rect 1788 3417 1810 3451
rect 1738 3367 1810 3417
rect 1738 3333 1754 3367
rect 1788 3333 1810 3367
rect 1738 3283 1810 3333
rect 1738 3249 1754 3283
rect 1788 3249 1810 3283
rect 1738 3233 1810 3249
rect 2462 3629 2534 3633
rect 2462 3595 2484 3629
rect 2518 3595 2534 3629
rect 2462 3579 2534 3595
rect 2462 3557 2540 3579
rect 2462 3523 2484 3557
rect 2518 3523 2540 3557
rect 2462 3485 2540 3523
rect 2462 3451 2484 3485
rect 2518 3479 2540 3485
rect 2518 3451 2534 3479
rect 2462 3423 2534 3451
rect 2462 3413 2540 3423
rect 2462 3379 2484 3413
rect 2518 3379 2540 3413
rect 2462 3341 2540 3379
rect 2462 3307 2484 3341
rect 2518 3323 2540 3341
rect 2518 3307 2534 3323
rect 2462 3269 2534 3307
rect 2462 3235 2484 3269
rect 2518 3267 2534 3269
rect 2518 3235 2540 3267
rect 2462 3233 2540 3235
rect 2468 3219 2540 3233
rect 1738 3161 1810 3177
rect 1738 3127 1754 3161
rect 1788 3127 1810 3161
rect 1738 3078 1810 3127
rect 1738 3044 1754 3078
rect 1788 3044 1810 3078
rect 1738 2995 1810 3044
rect 1738 2961 1754 2995
rect 1788 2961 1810 2995
rect 1738 2911 1810 2961
rect 1738 2877 1754 2911
rect 1788 2877 1810 2911
rect 1738 2827 1810 2877
rect 1738 2793 1754 2827
rect 1788 2793 1810 2827
rect 1738 2777 1810 2793
rect 2462 2955 2468 3177
rect 2534 3167 2540 3219
rect 2892 3078 3032 3111
rect 2892 3044 2914 3078
rect 2948 3044 2982 3078
rect 3016 3044 3032 3078
rect 2892 3011 3032 3044
rect 2462 2939 2540 2955
rect 2462 2905 2484 2939
rect 2518 2905 2540 2939
rect 2462 2855 2540 2905
rect 2892 2855 3032 2955
rect 2462 2813 2534 2855
rect 2462 2779 2484 2813
rect 2518 2799 2534 2813
rect 2898 2799 3032 2855
rect 2518 2779 2540 2799
rect 2462 2777 2540 2779
rect 2468 2763 2540 2777
rect 2510 2737 2540 2763
rect 1738 2705 1810 2721
rect 1738 2671 1754 2705
rect 1788 2671 1810 2705
rect 1738 2622 1810 2671
rect 1738 2588 1754 2622
rect 1788 2588 1810 2622
rect 1738 2539 1810 2588
rect 1738 2505 1754 2539
rect 1788 2505 1810 2539
rect 1738 2455 1810 2505
rect 1738 2421 1754 2455
rect 1788 2421 1810 2455
rect 1738 2371 1810 2421
rect 1738 2337 1754 2371
rect 1788 2337 1810 2371
rect 1738 2321 1810 2337
rect 2462 2321 2468 2721
rect 2534 2699 2540 2737
rect 2892 2699 3032 2799
rect 2892 2616 3032 2643
rect 2892 2582 2914 2616
rect 2948 2582 2982 2616
rect 3016 2582 3032 2616
rect 2892 2543 3032 2582
rect 2892 2470 3032 2487
rect 2892 2436 2914 2470
rect 2948 2436 2982 2470
rect 3016 2436 3032 2470
rect 2892 2387 3032 2436
rect 2534 2291 2540 2331
rect 2498 2265 2540 2291
rect 1738 2249 1810 2265
rect 1738 2215 1754 2249
rect 1788 2215 1810 2249
rect 1738 2166 1810 2215
rect 1738 2132 1754 2166
rect 1788 2132 1810 2166
rect 1738 2083 1810 2132
rect 1738 2049 1754 2083
rect 1788 2049 1810 2083
rect 1738 1999 1810 2049
rect 1738 1965 1754 1999
rect 1788 1965 1810 1999
rect 1738 1915 1810 1965
rect 1738 1881 1754 1915
rect 1788 1881 1810 1915
rect 1738 1865 1810 1881
rect 2462 2249 2540 2265
rect 2462 2215 2484 2249
rect 2518 2231 2540 2249
rect 2518 2215 2534 2231
rect 2462 2179 2534 2215
rect 2462 2145 2484 2179
rect 2518 2175 2534 2179
rect 2518 2145 2540 2175
rect 2462 2109 2540 2145
rect 2462 2075 2484 2109
rect 2518 2075 2540 2109
rect 2462 2039 2534 2075
rect 2462 2005 2484 2039
rect 2518 2019 2534 2039
rect 2518 2005 2540 2019
rect 2462 1969 2540 2005
rect 2462 1935 2484 1969
rect 2518 1935 2540 1969
rect 2462 1919 2540 1935
rect 2462 1899 2534 1919
rect 2462 1865 2484 1899
rect 2518 1865 2534 1899
rect 2468 1863 2534 1865
rect 2468 1828 2540 1863
rect 2468 1809 2484 1828
rect 1738 1793 1810 1809
rect 1738 1759 1754 1793
rect 1788 1759 1810 1793
rect 1738 1710 1810 1759
rect 1738 1676 1754 1710
rect 1788 1676 1810 1710
rect 1738 1627 1810 1676
rect 1738 1593 1754 1627
rect 1788 1593 1810 1627
rect 1738 1543 1810 1593
rect 1738 1509 1754 1543
rect 1788 1509 1810 1543
rect 1738 1459 1810 1509
rect 1738 1425 1754 1459
rect 1788 1425 1810 1459
rect 1738 1409 1810 1425
rect 2462 1794 2484 1809
rect 2518 1794 2540 1828
rect 2462 1763 2540 1794
rect 2462 1757 2534 1763
rect 2462 1723 2484 1757
rect 2518 1723 2534 1757
rect 2462 1707 2534 1723
rect 2462 1686 2540 1707
rect 2462 1652 2484 1686
rect 2518 1652 2540 1686
rect 2462 1615 2540 1652
rect 2462 1581 2484 1615
rect 2518 1607 2540 1615
rect 2518 1581 2534 1607
rect 2462 1551 2534 1581
rect 2462 1544 2540 1551
rect 2462 1510 2484 1544
rect 2518 1510 2540 1544
rect 2462 1473 2540 1510
rect 2462 1439 2484 1473
rect 2518 1451 2540 1473
rect 2518 1439 2534 1451
rect 2462 1409 2534 1439
rect 2468 1402 2534 1409
rect 2468 1368 2484 1402
rect 2518 1395 2534 1402
rect 2518 1368 2540 1395
rect 2468 1353 2540 1368
rect 1738 1337 1810 1353
rect 1738 1303 1754 1337
rect 1788 1303 1810 1337
rect 1738 1254 1810 1303
rect 1738 1220 1754 1254
rect 1788 1220 1810 1254
rect 1738 1171 1810 1220
rect 1738 1137 1754 1171
rect 1788 1137 1810 1171
rect 1738 1087 1810 1137
rect 1738 1053 1754 1087
rect 1788 1053 1810 1087
rect 1738 1003 1810 1053
rect 1738 969 1754 1003
rect 1788 969 1810 1003
rect 1738 953 1810 969
rect 2462 1331 2540 1353
rect 2462 1297 2484 1331
rect 2518 1297 2540 1331
rect 2462 1295 2540 1297
rect 2462 1260 2534 1295
rect 2462 1226 2484 1260
rect 2518 1239 2534 1260
rect 2518 1226 2540 1239
rect 2462 1189 2540 1226
rect 2462 1155 2484 1189
rect 2518 1155 2540 1189
rect 2462 1139 2540 1155
rect 2462 953 2468 1139
rect 2892 1050 3032 1083
rect 2892 1016 2914 1050
rect 2948 1016 2982 1050
rect 3016 1016 3032 1050
rect 2892 983 3032 1016
rect 2534 897 2540 927
rect 1738 881 1810 897
rect 1738 847 1754 881
rect 1788 847 1810 881
rect 1738 798 1810 847
rect 1738 764 1754 798
rect 1788 764 1810 798
rect 1738 715 1810 764
rect 1738 681 1754 715
rect 1788 681 1810 715
rect 1738 631 1810 681
rect 1738 597 1754 631
rect 1788 597 1810 631
rect 1738 547 1810 597
rect 1738 513 1754 547
rect 1788 513 1810 547
rect 1738 497 1810 513
rect 2462 881 2540 897
rect 2462 847 2484 881
rect 2518 847 2540 881
rect 2462 798 2540 847
rect 2462 764 2484 798
rect 2518 764 2540 798
rect 2462 715 2540 764
rect 2462 681 2484 715
rect 2518 681 2540 715
rect 2462 631 2540 681
rect 2462 597 2484 631
rect 2518 597 2540 631
rect 2462 547 2540 597
rect 2462 513 2484 547
rect 2518 527 2540 547
rect 2518 513 2534 527
rect 2462 497 2534 513
rect 3836 4936 3922 4952
rect 3836 4902 3852 4936
rect 3886 4902 3922 4936
rect 3836 4842 3922 4902
rect 3836 4808 3852 4842
rect 3886 4808 3922 4842
rect 3836 4792 3922 4808
rect 4124 4474 4190 4490
rect 4124 4440 4140 4474
rect 4174 4440 4190 4474
rect 4124 4400 4190 4440
rect 4124 4366 4140 4400
rect 4174 4366 4190 4400
rect 4124 4326 4190 4366
rect 4124 4292 4140 4326
rect 4174 4292 4190 4326
rect 4124 4252 4190 4292
rect 4124 4218 4140 4252
rect 4174 4218 4190 4252
rect 4124 4178 4190 4218
rect 4124 4144 4140 4178
rect 4174 4144 4190 4178
rect 4124 4104 4190 4144
rect 4124 4070 4140 4104
rect 4174 4070 4190 4104
rect 4124 4030 4190 4070
rect 4124 3996 4140 4030
rect 4174 3996 4190 4030
rect 4124 3956 4190 3996
rect 4124 3922 4140 3956
rect 4174 3922 4190 3956
rect 4124 3882 4190 3922
rect 4124 3848 4140 3882
rect 4174 3848 4190 3882
rect 4124 3808 4190 3848
rect 4124 3774 4140 3808
rect 4174 3774 4190 3808
rect 4124 3734 4190 3774
rect 4124 3700 4140 3734
rect 4174 3700 4190 3734
rect 4124 3660 4190 3700
rect 4124 3626 4140 3660
rect 4174 3626 4190 3660
rect 4124 3610 4190 3626
rect 3534 3394 3600 3410
rect 3534 3360 3550 3394
rect 3584 3360 3600 3394
rect 3534 3326 3600 3360
rect 3534 3292 3550 3326
rect 3584 3292 3600 3326
rect 3534 3276 3600 3292
rect 3764 3085 3872 3101
rect 3764 3051 3780 3085
rect 3814 3065 3872 3085
rect 3814 3051 3830 3065
rect 3764 3014 3830 3051
rect 3764 2980 3780 3014
rect 3814 2980 3830 3014
rect 3764 2943 3830 2980
rect 3764 2909 3780 2943
rect 3814 2909 3830 2943
rect 3764 2905 3830 2909
rect 3764 2872 3872 2905
rect 3764 2838 3780 2872
rect 3814 2869 3872 2872
rect 3814 2838 3830 2869
rect 3764 2801 3830 2838
rect 3764 2767 3780 2801
rect 3814 2767 3830 2801
rect 3764 2730 3830 2767
rect 3764 2696 3780 2730
rect 3814 2696 3830 2730
rect 3764 2659 3830 2696
rect 3764 2625 3780 2659
rect 3814 2629 3830 2659
rect 3814 2625 3872 2629
rect 3764 2593 3872 2625
rect 3764 2588 3830 2593
rect 3764 2554 3780 2588
rect 3814 2554 3830 2588
rect 3764 2517 3830 2554
rect 3764 2483 3780 2517
rect 3814 2483 3830 2517
rect 3764 2447 3830 2483
rect 3764 2413 3780 2447
rect 3814 2433 3830 2447
rect 3814 2413 3872 2433
rect 3764 2397 3872 2413
rect 3534 2155 3600 2171
rect 3534 2121 3550 2155
rect 3584 2121 3600 2155
rect 3534 2087 3600 2121
rect 3534 2053 3550 2087
rect 3584 2053 3600 2087
rect 3534 2037 3600 2053
rect 3836 2121 3922 2137
rect 3836 2087 3852 2121
rect 3886 2087 3922 2121
rect 3836 2027 3922 2087
rect 3836 1993 3852 2027
rect 3886 1993 3922 2027
rect 3836 1977 3922 1993
rect 4124 1393 4190 1409
rect 4124 1359 4140 1393
rect 4174 1359 4190 1393
rect 4124 1319 4190 1359
rect 4124 1285 4140 1319
rect 4174 1285 4190 1319
rect 4124 1245 4190 1285
rect 4124 1211 4140 1245
rect 4174 1211 4190 1245
rect 4124 1171 4190 1211
rect 4124 1137 4140 1171
rect 4174 1137 4190 1171
rect 4124 1097 4190 1137
rect 4124 1063 4140 1097
rect 4174 1063 4190 1097
rect 4124 1023 4190 1063
rect 4124 989 4140 1023
rect 4174 989 4190 1023
rect 4124 949 4190 989
rect 4124 915 4140 949
rect 4174 915 4190 949
rect 4124 875 4190 915
rect 4124 841 4140 875
rect 4174 841 4190 875
rect 4124 801 4190 841
rect 4124 767 4140 801
rect 4174 767 4190 801
rect 4124 727 4190 767
rect 4124 693 4140 727
rect 4174 693 4190 727
rect 4124 653 4190 693
rect 4124 619 4140 653
rect 4174 619 4190 653
rect 4124 579 4190 619
rect 4124 545 4140 579
rect 4174 545 4190 579
rect 4124 529 4190 545
rect 9668 4987 9848 5009
rect 9668 4953 9708 4987
rect 9742 4953 9776 4987
rect 9810 4953 9848 4987
rect 9668 4931 9848 4953
rect 9904 4987 10084 5009
rect 9904 4953 9944 4987
rect 9978 4953 10012 4987
rect 10046 4953 10084 4987
rect 9904 4931 10084 4953
rect 4930 3452 5002 3491
rect 4930 3418 4946 3452
rect 4980 3418 5002 3452
rect 4930 3384 5002 3418
rect 4930 3350 4946 3384
rect 4980 3350 5002 3384
rect 4930 3311 5002 3350
rect 7054 3311 7126 3491
rect 7168 3311 7240 3491
rect 9292 3452 9433 3491
rect 9292 3418 9314 3452
rect 9348 3418 9433 3452
rect 9292 3384 9433 3418
rect 9292 3350 9314 3384
rect 9348 3350 9433 3384
rect 9292 3311 9433 3350
rect 4930 3097 5002 3131
rect 4930 3063 4946 3097
rect 4980 3063 5002 3097
rect 4930 3029 5002 3063
rect 4930 2995 4946 3029
rect 4980 2995 5002 3029
rect 4930 2951 5002 2995
rect 7054 3092 7126 3131
rect 7054 3058 7076 3092
rect 7110 3058 7126 3092
rect 7054 3024 7126 3058
rect 7054 2990 7076 3024
rect 7110 2990 7126 3024
rect 7054 2951 7126 2990
rect 7168 3092 7240 3131
rect 7168 3058 7184 3092
rect 7218 3058 7240 3092
rect 7168 3024 7240 3058
rect 7168 2990 7184 3024
rect 7218 2990 7240 3024
rect 7168 2951 7240 2990
rect 9292 3092 9433 3131
rect 9292 3058 9314 3092
rect 9348 3058 9433 3092
rect 9292 3024 9433 3058
rect 9292 2990 9314 3024
rect 9348 2990 9433 3024
rect 9292 2951 9433 2990
rect 4930 2861 5002 2895
rect 4930 2827 4946 2861
rect 4980 2827 5002 2861
rect 4930 2793 5002 2827
rect 4930 2759 4946 2793
rect 4980 2759 5002 2793
rect 4930 2715 5002 2759
rect 7054 2856 7126 2895
rect 7054 2822 7076 2856
rect 7110 2822 7126 2856
rect 7054 2788 7126 2822
rect 7054 2754 7076 2788
rect 7110 2754 7126 2788
rect 7054 2715 7126 2754
rect 7168 2856 7240 2895
rect 7168 2822 7184 2856
rect 7218 2822 7240 2856
rect 7168 2788 7240 2822
rect 7168 2754 7184 2788
rect 7218 2754 7240 2788
rect 7168 2715 7240 2754
rect 9292 2856 9433 2895
rect 9292 2822 9314 2856
rect 9348 2822 9433 2856
rect 9292 2788 9433 2822
rect 9292 2754 9314 2788
rect 9348 2754 9433 2788
rect 9292 2715 9433 2754
rect 4930 2494 5002 2533
rect 4930 2460 4946 2494
rect 4980 2460 5002 2494
rect 4930 2426 5002 2460
rect 4930 2392 4946 2426
rect 4980 2392 5002 2426
rect 4930 2353 5002 2392
rect 7054 2494 7126 2533
rect 7054 2460 7076 2494
rect 7110 2460 7126 2494
rect 7054 2426 7126 2460
rect 7054 2392 7076 2426
rect 7110 2392 7126 2426
rect 7054 2353 7126 2392
rect 7168 2494 7240 2533
rect 7168 2460 7184 2494
rect 7218 2460 7240 2494
rect 7168 2426 7240 2460
rect 7168 2392 7184 2426
rect 7218 2392 7240 2426
rect 7168 2353 7240 2392
rect 9292 2494 9433 2533
rect 9292 2460 9314 2494
rect 9348 2460 9433 2494
rect 9292 2426 9433 2460
rect 9292 2392 9314 2426
rect 9348 2392 9433 2426
rect 9292 2353 9433 2392
rect 4930 2258 5002 2297
rect 4930 2224 4946 2258
rect 4980 2224 5002 2258
rect 4930 2190 5002 2224
rect 4930 2156 4946 2190
rect 4980 2156 5002 2190
rect 4930 2117 5002 2156
rect 7054 2258 7126 2297
rect 7054 2224 7076 2258
rect 7110 2224 7126 2258
rect 7054 2190 7126 2224
rect 7054 2156 7076 2190
rect 7110 2156 7126 2190
rect 7054 2117 7126 2156
rect 7168 2258 7240 2297
rect 7168 2224 7184 2258
rect 7218 2224 7240 2258
rect 7168 2190 7240 2224
rect 7168 2156 7184 2190
rect 7218 2156 7240 2190
rect 7168 2117 7240 2156
rect 9292 2258 9433 2297
rect 9292 2224 9314 2258
rect 9348 2224 9433 2258
rect 9292 2190 9433 2224
rect 9292 2156 9314 2190
rect 9348 2156 9433 2190
rect 9292 2117 9433 2156
rect 4930 1898 5002 1937
rect 4930 1864 4946 1898
rect 4980 1864 5002 1898
rect 4930 1830 5002 1864
rect 4930 1796 4946 1830
rect 4980 1796 5002 1830
rect 4930 1757 5002 1796
rect 9292 1898 9433 1937
rect 9292 1864 9314 1898
rect 9348 1864 9433 1898
rect 9292 1830 9433 1864
rect 9292 1796 9314 1830
rect 9348 1796 9433 1830
rect 9292 1757 9433 1796
rect 10384 4057 10456 4857
rect 11108 4057 11186 4857
rect 11838 4057 11916 4857
rect 12568 4057 12640 4857
rect 10384 3952 10456 4001
rect 10384 3918 10400 3952
rect 10434 3918 10456 3952
rect 10384 3884 10456 3918
rect 10384 3850 10400 3884
rect 10434 3850 10456 3884
rect 10384 3801 10456 3850
rect 11108 3952 11186 4001
rect 11108 3918 11130 3952
rect 11164 3918 11186 3952
rect 11108 3884 11186 3918
rect 11108 3850 11130 3884
rect 11164 3850 11186 3884
rect 11108 3801 11186 3850
rect 12568 3892 12640 4001
rect 12568 3858 12590 3892
rect 12624 3858 12640 3892
rect 12568 3824 12640 3858
rect 12568 3790 12590 3824
rect 12624 3790 12640 3824
rect 12568 3756 12640 3790
rect 10384 3696 10456 3745
rect 10384 3662 10400 3696
rect 10434 3662 10456 3696
rect 10384 3628 10456 3662
rect 10384 3594 10400 3628
rect 10434 3594 10456 3628
rect 10384 3545 10456 3594
rect 11108 3696 11186 3745
rect 11108 3662 11130 3696
rect 11164 3662 11186 3696
rect 11108 3628 11186 3662
rect 11108 3594 11130 3628
rect 11164 3594 11186 3628
rect 11108 3545 11186 3594
rect 12568 3722 12590 3756
rect 12624 3722 12640 3756
rect 12568 3688 12640 3722
rect 12568 3654 12590 3688
rect 12624 3654 12640 3688
rect 12568 3545 12640 3654
rect 10384 3440 10456 3489
rect 10384 3406 10400 3440
rect 10434 3406 10456 3440
rect 10384 3372 10456 3406
rect 10384 3338 10400 3372
rect 10434 3338 10456 3372
rect 10384 3289 10456 3338
rect 11108 3440 11186 3489
rect 11108 3406 11130 3440
rect 11164 3406 11186 3440
rect 11108 3372 11186 3406
rect 11108 3338 11130 3372
rect 11164 3338 11186 3372
rect 11108 3289 11186 3338
rect 11838 3440 11916 3489
rect 11838 3406 11860 3440
rect 11894 3406 11916 3440
rect 11838 3372 11916 3406
rect 11838 3338 11860 3372
rect 11894 3338 11916 3372
rect 11838 3289 11916 3338
rect 12568 3440 12640 3489
rect 12568 3406 12590 3440
rect 12624 3406 12640 3440
rect 12568 3372 12640 3406
rect 12568 3338 12590 3372
rect 12624 3338 12640 3372
rect 12568 3289 12640 3338
rect 10384 3184 10456 3233
rect 10384 3150 10400 3184
rect 10434 3150 10456 3184
rect 10384 3116 10456 3150
rect 10384 3082 10400 3116
rect 10434 3082 10456 3116
rect 10384 3033 10456 3082
rect 11108 3184 11186 3233
rect 11108 3150 11130 3184
rect 11164 3150 11186 3184
rect 11108 3116 11186 3150
rect 11108 3082 11130 3116
rect 11164 3082 11186 3116
rect 11108 3033 11186 3082
rect 11838 3184 11916 3233
rect 11838 3150 11860 3184
rect 11894 3150 11916 3184
rect 11838 3116 11916 3150
rect 11838 3082 11860 3116
rect 11894 3082 11916 3116
rect 11838 3033 11916 3082
rect 12568 3184 12640 3233
rect 12568 3150 12590 3184
rect 12624 3150 12640 3184
rect 12568 3116 12640 3150
rect 12568 3082 12590 3116
rect 12624 3082 12640 3116
rect 12568 3033 12640 3082
rect 10384 2928 10456 2977
rect 10384 2894 10400 2928
rect 10434 2894 10456 2928
rect 10384 2860 10456 2894
rect 10384 2826 10400 2860
rect 10434 2826 10456 2860
rect 10384 2777 10456 2826
rect 11108 2928 11186 2977
rect 11108 2894 11130 2928
rect 11164 2894 11186 2928
rect 11108 2860 11186 2894
rect 11108 2826 11130 2860
rect 11164 2826 11186 2860
rect 11108 2777 11186 2826
rect 11838 2928 11916 2977
rect 11838 2894 11860 2928
rect 11894 2894 11916 2928
rect 11838 2860 11916 2894
rect 11838 2826 11860 2860
rect 11894 2826 11916 2860
rect 11838 2777 11916 2826
rect 12568 2928 12640 2977
rect 12568 2894 12590 2928
rect 12624 2894 12640 2928
rect 12568 2860 12640 2894
rect 12568 2826 12590 2860
rect 12624 2826 12640 2860
rect 12568 2777 12640 2826
rect 10384 2672 10456 2721
rect 10384 2638 10400 2672
rect 10434 2638 10456 2672
rect 10384 2604 10456 2638
rect 10384 2570 10400 2604
rect 10434 2570 10456 2604
rect 10384 2521 10456 2570
rect 11108 2672 11186 2721
rect 11108 2638 11130 2672
rect 11164 2638 11186 2672
rect 11108 2604 11186 2638
rect 11108 2570 11130 2604
rect 11164 2570 11186 2604
rect 11108 2521 11186 2570
rect 11838 2672 11916 2721
rect 11838 2638 11860 2672
rect 11894 2638 11916 2672
rect 11838 2604 11916 2638
rect 11838 2570 11860 2604
rect 11894 2570 11916 2604
rect 11838 2521 11916 2570
rect 12568 2672 12640 2721
rect 12568 2638 12590 2672
rect 12624 2638 12640 2672
rect 12568 2604 12640 2638
rect 12568 2570 12590 2604
rect 12624 2570 12640 2604
rect 12568 2521 12640 2570
rect 10384 2416 10456 2465
rect 10384 2382 10400 2416
rect 10434 2382 10456 2416
rect 10384 2348 10456 2382
rect 10384 2314 10400 2348
rect 10434 2314 10456 2348
rect 10384 2265 10456 2314
rect 11108 2416 11186 2465
rect 11108 2382 11130 2416
rect 11164 2382 11186 2416
rect 11108 2348 11186 2382
rect 11108 2314 11130 2348
rect 11164 2314 11186 2348
rect 11108 2265 11186 2314
rect 11838 2416 11916 2465
rect 11838 2382 11860 2416
rect 11894 2382 11916 2416
rect 11838 2348 11916 2382
rect 11838 2314 11860 2348
rect 11894 2314 11916 2348
rect 11838 2265 11916 2314
rect 12568 2265 12640 2465
rect 10384 2160 10456 2209
rect 10384 2126 10400 2160
rect 10434 2126 10456 2160
rect 10384 2092 10456 2126
rect 10384 2058 10400 2092
rect 10434 2058 10456 2092
rect 10384 2009 10456 2058
rect 11108 2160 11186 2209
rect 11108 2126 11130 2160
rect 11164 2126 11186 2160
rect 11108 2092 11186 2126
rect 11108 2058 11130 2092
rect 11164 2058 11186 2092
rect 11108 2009 11186 2058
rect 11838 2160 11916 2209
rect 11838 2126 11860 2160
rect 11894 2126 11916 2160
rect 11838 2092 11916 2126
rect 11838 2058 11860 2092
rect 11894 2058 11916 2092
rect 11838 2009 11916 2058
rect 12568 2160 12640 2209
rect 12568 2126 12590 2160
rect 12624 2126 12640 2160
rect 12568 2092 12640 2126
rect 12568 2058 12590 2092
rect 12624 2058 12640 2092
rect 12568 2009 12640 2058
rect 10384 1904 10456 1953
rect 10384 1870 10400 1904
rect 10434 1870 10456 1904
rect 10384 1836 10456 1870
rect 10384 1802 10400 1836
rect 10434 1802 10456 1836
rect 10384 1753 10456 1802
rect 11108 1904 11186 1953
rect 11108 1870 11130 1904
rect 11164 1870 11186 1904
rect 11108 1836 11186 1870
rect 11108 1802 11130 1836
rect 11164 1802 11186 1836
rect 11108 1753 11186 1802
rect 12568 1904 12640 1953
rect 12568 1870 12590 1904
rect 12624 1870 12640 1904
rect 12568 1836 12640 1870
rect 12568 1802 12590 1836
rect 12624 1802 12640 1836
rect 12568 1753 12640 1802
rect 10384 1648 10456 1697
rect 10384 1614 10400 1648
rect 10434 1614 10456 1648
rect 10384 1580 10456 1614
rect 10384 1546 10400 1580
rect 10434 1546 10456 1580
rect 10384 1497 10456 1546
rect 11108 1648 11186 1697
rect 11108 1614 11130 1648
rect 11164 1614 11186 1648
rect 11108 1580 11186 1614
rect 11108 1546 11130 1580
rect 11164 1546 11186 1580
rect 11108 1497 11186 1546
rect 12568 1648 12640 1697
rect 12568 1614 12590 1648
rect 12624 1614 12640 1648
rect 12568 1580 12640 1614
rect 12568 1546 12590 1580
rect 12624 1546 12640 1580
rect 12568 1497 12640 1546
rect 9668 604 9848 627
rect 9668 570 9708 604
rect 9742 570 9776 604
rect 9810 570 9848 604
rect 9668 549 9848 570
rect 9904 605 10084 627
rect 9904 571 9944 605
rect 9978 571 10012 605
rect 10046 571 10084 605
rect 9904 549 10084 571
rect 10384 641 10456 1441
rect 11108 641 11186 1441
rect 11838 641 11916 1441
rect 12568 641 12640 1441
<< polycont >>
rect 10221 11294 10255 11328
rect 10291 11294 10325 11328
rect 10361 11294 10395 11328
rect 10431 11294 10465 11328
rect 10500 11294 10534 11328
rect 10569 11294 10603 11328
rect 10638 11294 10672 11328
rect 10707 11294 10741 11328
rect 10776 11294 10810 11328
rect 10845 11294 10879 11328
rect 10914 11294 10948 11328
rect 10983 11294 11017 11328
rect 11052 11294 11086 11328
rect 11121 11294 11155 11328
rect 11190 11294 11224 11328
rect 11259 11294 11293 11328
rect 11328 11294 11362 11328
rect 11397 11294 11431 11328
rect 11466 11294 11500 11328
rect 11535 11294 11569 11328
rect 11604 11294 11638 11328
rect 11673 11294 11707 11328
rect 11742 11294 11776 11328
rect 11811 11294 11845 11328
rect 6504 10403 6538 10437
rect 6573 10403 6607 10437
rect 6642 10403 6676 10437
rect 6711 10403 6745 10437
rect 6780 10403 6814 10437
rect 6849 10403 6883 10437
rect 6918 10403 6952 10437
rect 6987 10403 7021 10437
rect 7056 10403 7090 10437
rect 7125 10403 7159 10437
rect 7194 10403 7228 10437
rect 7263 10403 7297 10437
rect 7332 10403 7366 10437
rect 7401 10403 7435 10437
rect 7470 10403 7504 10437
rect 7539 10403 7573 10437
rect 7608 10403 7642 10437
rect 7677 10403 7711 10437
rect 7746 10403 7780 10437
rect 7815 10403 7849 10437
rect 7884 10403 7918 10437
rect 7953 10403 7987 10437
rect 8022 10403 8056 10437
rect 8091 10403 8125 10437
rect 8160 10403 8194 10437
rect 8229 10403 8263 10437
rect 8298 10403 8332 10437
rect 8367 10403 8401 10437
rect 8436 10403 8470 10437
rect 8505 10403 8539 10437
rect 8574 10403 8608 10437
rect 8643 10403 8677 10437
rect 8712 10403 8746 10437
rect 8781 10403 8815 10437
rect 8850 10403 8884 10437
rect 8919 10403 8953 10437
rect 8988 10403 9022 10437
rect 9057 10403 9091 10437
rect 9126 10403 9160 10437
rect 9195 10403 9229 10437
rect 9264 10403 9298 10437
rect 9333 10403 9367 10437
rect 9402 10403 9436 10437
rect 9471 10403 9505 10437
rect 9540 10403 9574 10437
rect 9609 10403 9643 10437
rect 9678 10403 9712 10437
rect 9747 10403 9781 10437
rect 9816 10403 9850 10437
rect 9885 10403 9919 10437
rect 9954 10403 9988 10437
rect 10022 10403 10056 10437
rect 10090 10403 10124 10437
rect 10158 10403 10192 10437
rect 10226 10403 10260 10437
rect 10294 10403 10328 10437
rect 10362 10403 10396 10437
rect 10430 10403 10464 10437
rect 10498 10403 10532 10437
rect 10566 10403 10600 10437
rect 10634 10403 10668 10437
rect 10702 10403 10736 10437
rect 10770 10403 10804 10437
rect 10838 10403 10872 10437
rect 10906 10403 10940 10437
rect 10974 10403 11008 10437
rect 11042 10403 11076 10437
rect 11110 10403 11144 10437
rect 11178 10403 11212 10437
rect 11246 10403 11280 10437
rect 11314 10403 11348 10437
rect 11382 10403 11416 10437
rect 11450 10403 11484 10437
rect 11518 10403 11552 10437
rect 6504 9519 6538 9553
rect 6573 9519 6607 9553
rect 6642 9519 6676 9553
rect 6711 9519 6745 9553
rect 6780 9519 6814 9553
rect 6849 9519 6883 9553
rect 6918 9519 6952 9553
rect 6987 9519 7021 9553
rect 7056 9519 7090 9553
rect 7125 9519 7159 9553
rect 7194 9519 7228 9553
rect 7263 9519 7297 9553
rect 7332 9519 7366 9553
rect 7401 9519 7435 9553
rect 7470 9519 7504 9553
rect 7539 9519 7573 9553
rect 7608 9519 7642 9553
rect 7677 9519 7711 9553
rect 7746 9519 7780 9553
rect 7815 9519 7849 9553
rect 7884 9519 7918 9553
rect 7953 9519 7987 9553
rect 8022 9519 8056 9553
rect 8091 9519 8125 9553
rect 8160 9519 8194 9553
rect 8229 9519 8263 9553
rect 8298 9519 8332 9553
rect 8367 9519 8401 9553
rect 8436 9519 8470 9553
rect 8505 9519 8539 9553
rect 8574 9519 8608 9553
rect 8643 9519 8677 9553
rect 8712 9519 8746 9553
rect 8781 9519 8815 9553
rect 8850 9519 8884 9553
rect 8918 9519 8952 9553
rect 8986 9519 9020 9553
rect 9054 9519 9088 9553
rect 9122 9519 9156 9553
rect 9190 9519 9224 9553
rect 9258 9519 9292 9553
rect 9326 9519 9360 9553
rect 9394 9519 9428 9553
rect 9462 9519 9496 9553
rect 9530 9519 9564 9553
rect 9598 9519 9632 9553
rect 9666 9519 9700 9553
rect 9734 9519 9768 9553
rect 9802 9519 9836 9553
rect 693 6042 727 6076
rect 693 5970 727 6004
rect 693 5898 727 5932
rect 693 5825 727 5859
rect 693 5752 727 5786
rect 693 5679 727 5713
rect 693 5606 727 5640
rect 693 5533 727 5567
rect 693 5460 727 5494
rect 335 5338 369 5372
rect 335 5261 369 5295
rect 335 5184 369 5218
rect 335 5108 369 5142
rect 693 4876 727 4910
rect 693 4808 727 4842
rect 335 4720 369 4754
rect 335 4652 369 4686
rect 1052 6042 1086 6076
rect 1052 5965 1086 5999
rect 1052 5888 1086 5922
rect 1052 5812 1086 5846
rect 1052 5690 1086 5724
rect 1052 5622 1086 5656
rect 1089 5404 1123 5438
rect 1089 5270 1123 5304
rect 1058 5148 1092 5182
rect 1058 5014 1092 5048
rect 351 4099 385 4133
rect 351 4017 385 4051
rect 351 3936 385 3970
rect 351 3855 385 3889
rect 351 3774 385 3808
rect 351 3693 385 3727
rect 1052 4782 1086 4816
rect 1052 4713 1086 4747
rect 1052 4644 1086 4678
rect 1052 4575 1086 4609
rect 1052 4506 1086 4540
rect 1052 4437 1086 4471
rect 1052 4368 1086 4402
rect 1052 4300 1086 4334
rect 1052 4232 1086 4266
rect 1052 4164 1086 4198
rect 1052 4096 1086 4130
rect 1052 4028 1086 4062
rect 1052 3960 1086 3994
rect 1052 3704 1086 3738
rect 1052 3630 1086 3664
rect 1052 3556 1086 3590
rect 1052 3482 1086 3516
rect 349 3148 383 3182
rect 349 3080 383 3114
rect 693 3044 727 3078
rect 693 2976 727 3010
rect 335 2854 369 2888
rect 335 2777 369 2811
rect 335 2700 369 2734
rect 693 2502 727 2536
rect 693 2434 727 2468
rect 363 2312 397 2346
rect 363 2244 397 2278
rect 1052 3302 1086 3336
rect 1052 3234 1086 3268
rect 1386 3112 1420 3146
rect 1052 3008 1086 3042
rect 1386 3044 1420 3078
rect 1052 2940 1086 2974
rect 1386 2708 1420 2742
rect 1386 2631 1420 2665
rect 1386 2554 1420 2588
rect 1386 2432 1420 2466
rect 1386 2355 1420 2389
rect 1386 2278 1420 2312
rect 1052 2156 1086 2190
rect 1052 2088 1086 2122
rect 349 1733 383 1767
rect 349 1651 383 1685
rect 349 1570 383 1604
rect 349 1489 383 1523
rect 349 1408 383 1442
rect 349 1327 383 1361
rect 349 1095 383 1129
rect 349 1022 383 1056
rect 349 949 383 983
rect 349 876 383 910
rect 349 803 383 837
rect 349 730 383 764
rect 349 657 383 691
rect 349 585 383 619
rect 349 513 383 547
rect 1052 1813 1086 1847
rect 1052 1739 1086 1773
rect 1052 1665 1086 1699
rect 1052 1591 1086 1625
rect 1052 1335 1086 1369
rect 1052 1266 1086 1300
rect 1052 1197 1086 1231
rect 1052 1128 1086 1162
rect 1052 1059 1086 1093
rect 1052 990 1086 1024
rect 1052 921 1086 955
rect 1052 853 1086 887
rect 1052 785 1086 819
rect 1052 717 1086 751
rect 1052 649 1086 683
rect 1052 581 1086 615
rect 1052 513 1086 547
rect 1754 4951 1788 4985
rect 1754 4868 1788 4902
rect 1754 4785 1788 4819
rect 1754 4701 1788 4735
rect 1754 4617 1788 4651
rect 2484 4951 2518 4985
rect 2484 4868 2518 4902
rect 2484 4785 2518 4819
rect 2484 4701 2518 4735
rect 2484 4617 2518 4651
rect 1754 4495 1788 4529
rect 1754 4412 1788 4446
rect 1754 4329 1788 4363
rect 1754 4245 1788 4279
rect 1754 4161 1788 4195
rect 2914 4448 2948 4482
rect 2982 4448 3016 4482
rect 2484 4309 2518 4343
rect 2484 4238 2518 4272
rect 2484 4167 2518 4201
rect 2484 4096 2518 4130
rect 1754 4039 1788 4073
rect 1754 3956 1788 3990
rect 1754 3873 1788 3907
rect 1754 3789 1788 3823
rect 1754 3705 1788 3739
rect 2484 4025 2518 4059
rect 2484 3954 2518 3988
rect 2484 3883 2518 3917
rect 2484 3811 2518 3845
rect 2484 3739 2518 3773
rect 2484 3667 2518 3701
rect 1754 3583 1788 3617
rect 1754 3500 1788 3534
rect 1754 3417 1788 3451
rect 1754 3333 1788 3367
rect 1754 3249 1788 3283
rect 2484 3595 2518 3629
rect 2484 3523 2518 3557
rect 2484 3451 2518 3485
rect 2484 3379 2518 3413
rect 2484 3307 2518 3341
rect 2484 3235 2518 3269
rect 1754 3127 1788 3161
rect 1754 3044 1788 3078
rect 1754 2961 1788 2995
rect 1754 2877 1788 2911
rect 1754 2793 1788 2827
rect 2914 3044 2948 3078
rect 2982 3044 3016 3078
rect 2484 2905 2518 2939
rect 2484 2779 2518 2813
rect 1754 2671 1788 2705
rect 1754 2588 1788 2622
rect 1754 2505 1788 2539
rect 1754 2421 1788 2455
rect 1754 2337 1788 2371
rect 2914 2582 2948 2616
rect 2982 2582 3016 2616
rect 2914 2436 2948 2470
rect 2982 2436 3016 2470
rect 1754 2215 1788 2249
rect 1754 2132 1788 2166
rect 1754 2049 1788 2083
rect 1754 1965 1788 1999
rect 1754 1881 1788 1915
rect 2484 2215 2518 2249
rect 2484 2145 2518 2179
rect 2484 2075 2518 2109
rect 2484 2005 2518 2039
rect 2484 1935 2518 1969
rect 2484 1865 2518 1899
rect 1754 1759 1788 1793
rect 1754 1676 1788 1710
rect 1754 1593 1788 1627
rect 1754 1509 1788 1543
rect 1754 1425 1788 1459
rect 2484 1794 2518 1828
rect 2484 1723 2518 1757
rect 2484 1652 2518 1686
rect 2484 1581 2518 1615
rect 2484 1510 2518 1544
rect 2484 1439 2518 1473
rect 2484 1368 2518 1402
rect 1754 1303 1788 1337
rect 1754 1220 1788 1254
rect 1754 1137 1788 1171
rect 1754 1053 1788 1087
rect 1754 969 1788 1003
rect 2484 1297 2518 1331
rect 2484 1226 2518 1260
rect 2484 1155 2518 1189
rect 2914 1016 2948 1050
rect 2982 1016 3016 1050
rect 1754 847 1788 881
rect 1754 764 1788 798
rect 1754 681 1788 715
rect 1754 597 1788 631
rect 1754 513 1788 547
rect 2484 847 2518 881
rect 2484 764 2518 798
rect 2484 681 2518 715
rect 2484 597 2518 631
rect 2484 513 2518 547
rect 3852 4902 3886 4936
rect 3852 4808 3886 4842
rect 4140 4440 4174 4474
rect 4140 4366 4174 4400
rect 4140 4292 4174 4326
rect 4140 4218 4174 4252
rect 4140 4144 4174 4178
rect 4140 4070 4174 4104
rect 4140 3996 4174 4030
rect 4140 3922 4174 3956
rect 4140 3848 4174 3882
rect 4140 3774 4174 3808
rect 4140 3700 4174 3734
rect 4140 3626 4174 3660
rect 3550 3360 3584 3394
rect 3550 3292 3584 3326
rect 3780 3051 3814 3085
rect 3780 2980 3814 3014
rect 3780 2909 3814 2943
rect 3780 2838 3814 2872
rect 3780 2767 3814 2801
rect 3780 2696 3814 2730
rect 3780 2625 3814 2659
rect 3780 2554 3814 2588
rect 3780 2483 3814 2517
rect 3780 2413 3814 2447
rect 3550 2121 3584 2155
rect 3550 2053 3584 2087
rect 3852 2087 3886 2121
rect 3852 1993 3886 2027
rect 4140 1359 4174 1393
rect 4140 1285 4174 1319
rect 4140 1211 4174 1245
rect 4140 1137 4174 1171
rect 4140 1063 4174 1097
rect 4140 989 4174 1023
rect 4140 915 4174 949
rect 4140 841 4174 875
rect 4140 767 4174 801
rect 4140 693 4174 727
rect 4140 619 4174 653
rect 4140 545 4174 579
rect 9708 4953 9742 4987
rect 9776 4953 9810 4987
rect 9944 4953 9978 4987
rect 10012 4953 10046 4987
rect 4946 3418 4980 3452
rect 4946 3350 4980 3384
rect 9314 3418 9348 3452
rect 9314 3350 9348 3384
rect 4946 3063 4980 3097
rect 4946 2995 4980 3029
rect 7076 3058 7110 3092
rect 7076 2990 7110 3024
rect 7184 3058 7218 3092
rect 7184 2990 7218 3024
rect 9314 3058 9348 3092
rect 9314 2990 9348 3024
rect 4946 2827 4980 2861
rect 4946 2759 4980 2793
rect 7076 2822 7110 2856
rect 7076 2754 7110 2788
rect 7184 2822 7218 2856
rect 7184 2754 7218 2788
rect 9314 2822 9348 2856
rect 9314 2754 9348 2788
rect 4946 2460 4980 2494
rect 4946 2392 4980 2426
rect 7076 2460 7110 2494
rect 7076 2392 7110 2426
rect 7184 2460 7218 2494
rect 7184 2392 7218 2426
rect 9314 2460 9348 2494
rect 9314 2392 9348 2426
rect 4946 2224 4980 2258
rect 4946 2156 4980 2190
rect 7076 2224 7110 2258
rect 7076 2156 7110 2190
rect 7184 2224 7218 2258
rect 7184 2156 7218 2190
rect 9314 2224 9348 2258
rect 9314 2156 9348 2190
rect 4946 1864 4980 1898
rect 4946 1796 4980 1830
rect 9314 1864 9348 1898
rect 9314 1796 9348 1830
rect 10400 3918 10434 3952
rect 10400 3850 10434 3884
rect 11130 3918 11164 3952
rect 11130 3850 11164 3884
rect 12590 3858 12624 3892
rect 12590 3790 12624 3824
rect 10400 3662 10434 3696
rect 10400 3594 10434 3628
rect 11130 3662 11164 3696
rect 11130 3594 11164 3628
rect 12590 3722 12624 3756
rect 12590 3654 12624 3688
rect 10400 3406 10434 3440
rect 10400 3338 10434 3372
rect 11130 3406 11164 3440
rect 11130 3338 11164 3372
rect 11860 3406 11894 3440
rect 11860 3338 11894 3372
rect 12590 3406 12624 3440
rect 12590 3338 12624 3372
rect 10400 3150 10434 3184
rect 10400 3082 10434 3116
rect 11130 3150 11164 3184
rect 11130 3082 11164 3116
rect 11860 3150 11894 3184
rect 11860 3082 11894 3116
rect 12590 3150 12624 3184
rect 12590 3082 12624 3116
rect 10400 2894 10434 2928
rect 10400 2826 10434 2860
rect 11130 2894 11164 2928
rect 11130 2826 11164 2860
rect 11860 2894 11894 2928
rect 11860 2826 11894 2860
rect 12590 2894 12624 2928
rect 12590 2826 12624 2860
rect 10400 2638 10434 2672
rect 10400 2570 10434 2604
rect 11130 2638 11164 2672
rect 11130 2570 11164 2604
rect 11860 2638 11894 2672
rect 11860 2570 11894 2604
rect 12590 2638 12624 2672
rect 12590 2570 12624 2604
rect 10400 2382 10434 2416
rect 10400 2314 10434 2348
rect 11130 2382 11164 2416
rect 11130 2314 11164 2348
rect 11860 2382 11894 2416
rect 11860 2314 11894 2348
rect 10400 2126 10434 2160
rect 10400 2058 10434 2092
rect 11130 2126 11164 2160
rect 11130 2058 11164 2092
rect 11860 2126 11894 2160
rect 11860 2058 11894 2092
rect 12590 2126 12624 2160
rect 12590 2058 12624 2092
rect 10400 1870 10434 1904
rect 10400 1802 10434 1836
rect 11130 1870 11164 1904
rect 11130 1802 11164 1836
rect 12590 1870 12624 1904
rect 12590 1802 12624 1836
rect 10400 1614 10434 1648
rect 10400 1546 10434 1580
rect 11130 1614 11164 1648
rect 11130 1546 11164 1580
rect 12590 1614 12624 1648
rect 12590 1546 12624 1580
rect 9708 570 9742 604
rect 9776 570 9810 604
rect 9944 571 9978 605
rect 10012 571 10046 605
<< locali >>
rect 6155 13067 9999 13073
rect 6155 13061 6281 13067
rect 6155 13027 6161 13061
rect 6195 13033 6281 13061
rect 6315 13033 6353 13067
rect 6387 13033 6425 13067
rect 6459 13033 6497 13067
rect 6531 13033 6569 13067
rect 6603 13033 6641 13067
rect 6675 13033 6713 13067
rect 6747 13033 6785 13067
rect 6819 13033 6857 13067
rect 6891 13033 6929 13067
rect 6963 13033 7001 13067
rect 7035 13033 7073 13067
rect 7107 13033 7145 13067
rect 7179 13033 7217 13067
rect 7251 13033 7289 13067
rect 7323 13033 7361 13067
rect 7395 13033 7433 13067
rect 7467 13033 7505 13067
rect 7539 13033 7577 13067
rect 7611 13033 7649 13067
rect 7683 13033 7721 13067
rect 7755 13033 7793 13067
rect 7827 13033 7865 13067
rect 7899 13033 7937 13067
rect 7971 13033 8009 13067
rect 8043 13033 8081 13067
rect 8115 13033 8153 13067
rect 8187 13033 8225 13067
rect 8259 13033 8297 13067
rect 8331 13033 8369 13067
rect 8403 13033 8441 13067
rect 8475 13033 8513 13067
rect 8547 13033 8585 13067
rect 8619 13033 8657 13067
rect 8691 13033 8729 13067
rect 8763 13033 8801 13067
rect 8835 13033 8873 13067
rect 8907 13033 8945 13067
rect 8979 13033 9017 13067
rect 9051 13033 9089 13067
rect 9123 13033 9161 13067
rect 9195 13033 9233 13067
rect 9267 13033 9305 13067
rect 9339 13033 9377 13067
rect 9411 13033 9449 13067
rect 9483 13033 9521 13067
rect 9555 13033 9593 13067
rect 9627 13033 9665 13067
rect 9699 13033 9737 13067
rect 9771 13033 9809 13067
rect 9843 13033 9881 13067
rect 9915 13033 9953 13067
rect 9987 13033 9999 13067
rect 6195 13027 9999 13033
rect 6155 12989 6201 13027
rect 6155 12955 6161 12989
rect 6195 12955 6201 12989
rect 6155 12917 6201 12955
rect 6155 12883 6161 12917
rect 6195 12883 6201 12917
rect 6155 12845 6201 12883
rect 6155 12811 6161 12845
rect 6195 12811 6201 12845
rect 6155 12773 6201 12811
rect 6155 12739 6161 12773
rect 6195 12739 6201 12773
rect 6155 12701 6201 12739
rect 6155 12667 6161 12701
rect 6195 12667 6201 12701
rect 6155 12629 6201 12667
rect 6155 12595 6161 12629
rect 6195 12595 6201 12629
rect 6155 12557 6201 12595
rect 6155 12523 6161 12557
rect 6195 12523 6201 12557
rect 6155 12485 6201 12523
rect 6155 12451 6161 12485
rect 6195 12451 6201 12485
rect 6155 12413 6201 12451
rect 6155 12379 6161 12413
rect 6195 12379 6201 12413
rect 6155 12341 6201 12379
rect 6155 12307 6161 12341
rect 6195 12307 6201 12341
rect 6155 12269 6201 12307
rect 6155 12235 6161 12269
rect 6195 12235 6201 12269
rect 6155 12197 6201 12235
rect 6155 12163 6161 12197
rect 6195 12163 6201 12197
rect 6155 12125 6201 12163
rect 6155 12091 6161 12125
rect 6195 12091 6201 12125
rect 6155 12053 6201 12091
rect 10008 12116 12060 12120
rect 10008 12082 10070 12116
rect 10104 12082 10155 12116
rect 10189 12082 10240 12116
rect 10274 12082 10325 12116
rect 10359 12082 10410 12116
rect 10444 12082 10495 12116
rect 10529 12082 10580 12116
rect 10614 12082 10665 12116
rect 10699 12082 10750 12116
rect 10784 12082 10835 12116
rect 10869 12082 10920 12116
rect 10954 12082 11005 12116
rect 11039 12082 11090 12116
rect 11124 12082 11175 12116
rect 11209 12082 11260 12116
rect 11294 12082 11345 12116
rect 11379 12082 11430 12116
rect 11464 12082 11515 12116
rect 11549 12082 11600 12116
rect 11634 12082 11685 12116
rect 11719 12082 11770 12116
rect 11804 12082 11856 12116
rect 11890 12082 11942 12116
rect 11976 12082 12060 12116
rect 10008 12078 12060 12082
rect 6155 12019 6161 12053
rect 6195 12019 6201 12053
rect 6155 11981 6201 12019
rect 6155 11947 6161 11981
rect 6195 11947 6201 11981
rect 6155 11909 6201 11947
rect 6155 11875 6161 11909
rect 6195 11875 6201 11909
rect 12018 12027 12060 12078
rect 12018 11993 12022 12027
rect 12056 11993 12060 12027
rect 12018 11934 12060 11993
rect 12018 11908 12022 11934
rect 6155 11837 6201 11875
rect 6155 11803 6161 11837
rect 6195 11803 6201 11837
rect 6155 11765 6201 11803
rect 6155 11731 6161 11765
rect 6195 11731 6201 11765
rect 6155 11693 6201 11731
rect 6155 11659 6161 11693
rect 6195 11659 6201 11693
rect 6155 11621 6201 11659
rect 10016 11900 12022 11908
rect 12056 11900 12060 11934
rect 10016 11841 12060 11900
rect 10016 11807 12022 11841
rect 12056 11807 12060 11841
rect 10016 11748 12060 11807
rect 10016 11714 12022 11748
rect 12056 11714 12060 11748
rect 10016 11655 12060 11714
rect 10016 11645 12022 11655
rect 6155 11587 6161 11621
rect 6195 11587 6201 11621
rect 6155 11549 6201 11587
rect 6155 11515 6161 11549
rect 6195 11515 6201 11549
rect 9982 11621 12022 11645
rect 12056 11621 12060 11655
rect 9982 11562 12060 11621
rect 9982 11539 12022 11562
rect 6155 11477 6201 11515
rect 6155 11443 6161 11477
rect 6195 11443 6201 11477
rect 6155 11405 6201 11443
rect 10016 11528 12022 11539
rect 12056 11528 12060 11562
rect 10016 11469 12060 11528
rect 10016 11435 12022 11469
rect 12056 11435 12060 11469
rect 10016 11414 12060 11435
rect 6155 11371 6161 11405
rect 6195 11371 6201 11405
rect 6155 11333 6201 11371
rect 6155 11299 6161 11333
rect 6195 11299 6201 11333
rect 12018 11376 12060 11414
rect 12018 11342 12022 11376
rect 12056 11342 12060 11376
rect 6155 11205 6201 11299
rect 10205 11294 10221 11328
rect 10255 11319 10291 11328
rect 10325 11319 10361 11328
rect 10395 11319 10431 11328
rect 10465 11319 10500 11328
rect 10266 11294 10291 11319
rect 10342 11294 10361 11319
rect 10418 11294 10431 11319
rect 10494 11294 10500 11319
rect 10534 11319 10569 11328
rect 10603 11319 10638 11328
rect 10672 11319 10707 11328
rect 10741 11319 10776 11328
rect 10810 11319 10845 11328
rect 10534 11294 10536 11319
rect 10603 11294 10612 11319
rect 10672 11294 10688 11319
rect 10741 11294 10764 11319
rect 10810 11294 10840 11319
rect 10879 11294 10914 11328
rect 10948 11319 10983 11328
rect 11017 11319 11052 11328
rect 11086 11319 11121 11328
rect 11155 11319 11190 11328
rect 11224 11319 11259 11328
rect 11293 11319 11328 11328
rect 10949 11294 10983 11319
rect 11024 11294 11052 11319
rect 11099 11294 11121 11319
rect 11174 11294 11190 11319
rect 11249 11294 11259 11319
rect 11324 11294 11328 11319
rect 11362 11319 11397 11328
rect 11431 11319 11466 11328
rect 11500 11319 11535 11328
rect 11569 11319 11604 11328
rect 11638 11319 11673 11328
rect 11707 11319 11742 11328
rect 11362 11294 11365 11319
rect 11431 11294 11440 11319
rect 11500 11294 11515 11319
rect 11569 11294 11590 11319
rect 11638 11294 11665 11319
rect 11707 11294 11740 11319
rect 11776 11294 11811 11328
rect 11845 11319 11861 11328
rect 11849 11294 11861 11319
rect 10266 11285 10308 11294
rect 10342 11285 10384 11294
rect 10418 11285 10460 11294
rect 10494 11285 10536 11294
rect 10570 11285 10612 11294
rect 10646 11285 10688 11294
rect 10722 11285 10764 11294
rect 10798 11285 10840 11294
rect 10874 11285 10915 11294
rect 10949 11285 10990 11294
rect 11024 11285 11065 11294
rect 11099 11285 11140 11294
rect 11174 11285 11215 11294
rect 11249 11285 11290 11294
rect 11324 11285 11365 11294
rect 11399 11285 11440 11294
rect 11474 11285 11515 11294
rect 11549 11285 11590 11294
rect 11624 11285 11665 11294
rect 11699 11285 11740 11294
rect 11774 11285 11815 11294
rect 12018 11283 12060 11342
rect 12018 11249 12022 11283
rect 12056 11249 12060 11283
rect 12018 11207 12060 11249
rect 6155 11199 8304 11205
rect 6155 11165 6167 11199
rect 6201 11165 6239 11199
rect 6273 11165 6311 11199
rect 6345 11165 6383 11199
rect 6417 11165 6455 11199
rect 6489 11165 6527 11199
rect 6561 11165 6599 11199
rect 6633 11165 6671 11199
rect 6705 11165 6743 11199
rect 6777 11165 6815 11199
rect 6849 11165 6887 11199
rect 6921 11165 6959 11199
rect 6993 11165 7031 11199
rect 7065 11165 7103 11199
rect 7137 11165 7175 11199
rect 7209 11165 7247 11199
rect 7281 11165 7319 11199
rect 7353 11165 7391 11199
rect 7425 11165 7463 11199
rect 7497 11165 7535 11199
rect 7569 11165 7607 11199
rect 7641 11165 7679 11199
rect 7713 11165 7751 11199
rect 7785 11165 7823 11199
rect 7857 11165 7895 11199
rect 7929 11165 7967 11199
rect 8001 11165 8039 11199
rect 8073 11165 8111 11199
rect 8145 11165 8183 11199
rect 8217 11165 8255 11199
rect 8289 11165 8304 11199
rect 10002 11203 12060 11207
rect 10002 11169 10066 11203
rect 10100 11169 10152 11203
rect 10186 11169 10238 11203
rect 10272 11169 10324 11203
rect 10358 11169 10410 11203
rect 10444 11169 10496 11203
rect 10530 11169 10582 11203
rect 10616 11169 10668 11203
rect 10702 11169 10754 11203
rect 10788 11169 10840 11203
rect 10874 11169 10927 11203
rect 10961 11169 11014 11203
rect 11048 11169 11101 11203
rect 11135 11169 11188 11203
rect 11222 11169 11275 11203
rect 11309 11169 11362 11203
rect 11396 11169 11449 11203
rect 11483 11169 11536 11203
rect 11570 11169 11623 11203
rect 11657 11169 11765 11203
rect 11799 11169 11852 11203
rect 11886 11169 11939 11203
rect 11973 11169 12060 11203
rect 10002 11165 12060 11169
rect 6155 11159 8304 11165
rect 1883 11057 2077 11106
rect 2155 11070 2189 11126
rect 6318 11108 6360 11159
rect 2530 11069 2589 11103
rect 6318 11074 6322 11108
rect 6356 11074 6360 11108
rect 6318 11023 6360 11074
rect 6318 10989 6322 11023
rect 6356 10989 6360 11023
rect 11699 11120 11741 11165
rect 11699 11086 11703 11120
rect 11737 11086 11741 11120
rect 11699 11033 11741 11086
rect 6318 10937 6360 10989
rect 6318 10903 6322 10937
rect 6356 10903 6360 10937
rect 6318 10851 6360 10903
rect 6318 10817 6322 10851
rect 6356 10817 6360 10851
rect 6318 10765 6360 10817
rect 6318 10731 6322 10765
rect 6356 10731 6360 10765
rect 6318 10679 6360 10731
rect 366 10632 1739 10666
rect 332 10600 1739 10632
rect 6318 10645 6322 10679
rect 6356 10645 6360 10679
rect 332 10594 366 10600
rect 6318 10593 6360 10645
rect 6318 10559 6322 10593
rect 6356 10559 6360 10593
rect 6318 10507 6360 10559
rect 6318 10473 6322 10507
rect 6356 10473 6360 10507
rect 6442 11014 11579 11017
rect 6442 10980 7070 11014
rect 7104 10980 7149 11014
rect 7183 10980 7228 11014
rect 7262 10980 7306 11014
rect 7340 10980 7384 11014
rect 7418 10980 7462 11014
rect 7496 10980 11579 11014
rect 6442 10936 11579 10980
rect 6442 10902 7070 10936
rect 7104 10902 7149 10936
rect 7183 10902 7228 10936
rect 7262 10902 7306 10936
rect 7340 10902 7384 10936
rect 7418 10902 7462 10936
rect 7496 10902 11579 10936
rect 6442 10475 11579 10902
rect 11699 10999 11703 11033
rect 11737 10999 11741 11033
rect 11699 10945 11741 10999
rect 11699 10911 11703 10945
rect 11737 10911 11741 10945
rect 11699 10857 11741 10911
rect 11699 10823 11703 10857
rect 11737 10823 11741 10857
rect 11699 10769 11741 10823
rect 11699 10735 11703 10769
rect 11737 10735 11741 10769
rect 11699 10681 11741 10735
rect 11699 10647 11703 10681
rect 11737 10647 11741 10681
rect 11699 10593 11741 10647
rect 11699 10559 11703 10593
rect 11737 10559 11741 10593
rect 11699 10505 11741 10559
rect 6318 10421 6360 10473
rect 11699 10471 11703 10505
rect 11737 10471 11741 10505
rect 6318 10387 6322 10421
rect 6356 10387 6360 10421
rect 6488 10403 6499 10437
rect 6538 10403 6572 10437
rect 6607 10403 6642 10437
rect 6679 10403 6711 10437
rect 6752 10403 6780 10437
rect 6825 10403 6849 10437
rect 6898 10403 6918 10437
rect 6971 10403 6987 10437
rect 7044 10403 7056 10437
rect 7117 10403 7125 10437
rect 7190 10403 7194 10437
rect 7228 10403 7229 10437
rect 7297 10403 7302 10437
rect 7366 10403 7375 10437
rect 7435 10403 7448 10437
rect 7504 10403 7521 10437
rect 7573 10403 7594 10437
rect 7642 10403 7667 10437
rect 7711 10403 7740 10437
rect 7780 10403 7813 10437
rect 7849 10403 7884 10437
rect 7920 10403 7953 10437
rect 7993 10403 8022 10437
rect 8066 10403 8091 10437
rect 8139 10403 8160 10437
rect 8212 10403 8229 10437
rect 8285 10403 8298 10437
rect 8358 10403 8367 10437
rect 8431 10403 8436 10437
rect 8504 10403 8505 10437
rect 8539 10403 8543 10437
rect 8608 10403 8616 10437
rect 8677 10403 8689 10437
rect 8746 10403 8762 10437
rect 8815 10403 8835 10437
rect 8884 10403 8908 10437
rect 8953 10403 8981 10437
rect 9022 10403 9054 10437
rect 9091 10403 9126 10437
rect 9161 10403 9195 10437
rect 9234 10403 9264 10437
rect 9307 10403 9333 10437
rect 9380 10403 9402 10437
rect 9453 10403 9471 10437
rect 9526 10403 9540 10437
rect 9599 10403 9609 10437
rect 9672 10403 9678 10437
rect 9745 10403 9747 10437
rect 9781 10403 9784 10437
rect 9850 10403 9857 10437
rect 9919 10403 9930 10437
rect 9988 10403 10003 10437
rect 10056 10403 10076 10437
rect 10124 10403 10149 10437
rect 10192 10403 10222 10437
rect 10260 10403 10294 10437
rect 10328 10403 10362 10437
rect 10400 10403 10430 10437
rect 10472 10403 10498 10437
rect 10544 10403 10566 10437
rect 10616 10403 10634 10437
rect 10688 10403 10702 10437
rect 10760 10403 10770 10437
rect 10832 10403 10838 10437
rect 10904 10403 10906 10437
rect 10940 10403 10942 10437
rect 11008 10403 11014 10437
rect 11076 10403 11086 10437
rect 11144 10403 11158 10437
rect 11212 10403 11230 10437
rect 11280 10403 11302 10437
rect 11348 10403 11374 10437
rect 11416 10403 11446 10437
rect 11484 10403 11518 10437
rect 11552 10403 11568 10437
rect 11699 10417 11741 10471
rect 6318 10341 6360 10387
rect 11699 10383 11703 10417
rect 11737 10383 11741 10417
rect 11699 10341 11741 10383
rect 6318 10337 11741 10341
rect 6318 10335 6417 10337
rect 6318 10301 6322 10335
rect 6356 10303 6417 10335
rect 6451 10303 6503 10337
rect 6537 10303 6589 10337
rect 6623 10303 6675 10337
rect 6709 10303 6761 10337
rect 6795 10303 6847 10337
rect 6881 10303 6933 10337
rect 6967 10303 7019 10337
rect 7053 10303 7105 10337
rect 7139 10303 7191 10337
rect 7225 10303 7277 10337
rect 7311 10303 7363 10337
rect 7397 10303 7449 10337
rect 7483 10303 7535 10337
rect 7569 10303 7621 10337
rect 7655 10303 7707 10337
rect 7741 10303 7793 10337
rect 7827 10303 7879 10337
rect 7913 10303 7965 10337
rect 7999 10303 8051 10337
rect 8085 10303 8137 10337
rect 8171 10303 8222 10337
rect 8256 10303 8307 10337
rect 8341 10303 8392 10337
rect 8426 10303 8477 10337
rect 8511 10303 8562 10337
rect 8596 10303 8647 10337
rect 8681 10303 8732 10337
rect 8766 10303 8817 10337
rect 8851 10303 8902 10337
rect 8936 10303 8987 10337
rect 9021 10303 9072 10337
rect 9106 10303 9157 10337
rect 9191 10303 9242 10337
rect 9276 10303 9327 10337
rect 9361 10303 9412 10337
rect 9446 10303 9497 10337
rect 9531 10303 9582 10337
rect 9616 10303 9667 10337
rect 9701 10303 9752 10337
rect 9786 10303 9837 10337
rect 9871 10303 9922 10337
rect 9956 10303 10007 10337
rect 10041 10303 10092 10337
rect 10126 10303 10177 10337
rect 10211 10303 10262 10337
rect 10296 10303 10347 10337
rect 10381 10303 10432 10337
rect 10466 10303 10517 10337
rect 10551 10303 10602 10337
rect 10636 10303 10687 10337
rect 10721 10303 10772 10337
rect 10806 10303 10857 10337
rect 10891 10303 10942 10337
rect 10976 10303 11027 10337
rect 11061 10303 11112 10337
rect 11146 10303 11197 10337
rect 11231 10303 11282 10337
rect 11316 10303 11367 10337
rect 11401 10303 11452 10337
rect 11486 10303 11537 10337
rect 11571 10303 11622 10337
rect 11656 10303 11741 10337
rect 6356 10301 11741 10303
rect 6318 10299 11741 10301
rect 6318 10249 6360 10299
rect 6318 10215 6322 10249
rect 6356 10215 6360 10249
rect 6318 10163 6360 10215
rect 6318 10129 6322 10163
rect 6356 10129 6360 10163
rect 10029 10238 10071 10299
rect 10029 10204 10033 10238
rect 10067 10204 10071 10238
rect 10029 10153 10071 10204
rect 6318 10077 6360 10129
rect 6318 10043 6322 10077
rect 6356 10043 6360 10077
rect 6318 9991 6360 10043
rect 6318 9957 6322 9991
rect 6356 9957 6360 9991
rect 6318 9905 6360 9957
rect 6318 9871 6322 9905
rect 6356 9871 6360 9905
rect 6318 9819 6360 9871
rect 6318 9785 6322 9819
rect 6356 9785 6360 9819
rect 6318 9733 6360 9785
rect 6318 9699 6322 9733
rect 6356 9699 6360 9733
rect 6318 9647 6360 9699
rect 6318 9613 6322 9647
rect 6356 9613 6360 9647
rect 6318 9561 6360 9613
rect 6442 10132 9909 10140
rect 6442 10098 7069 10132
rect 7103 10098 7147 10132
rect 7181 10098 7225 10132
rect 7259 10098 7372 10132
rect 7406 10098 7444 10132
rect 7478 10098 9909 10132
rect 6442 10051 9909 10098
rect 6442 10017 7069 10051
rect 7103 10017 7147 10051
rect 7181 10017 7225 10051
rect 7259 10017 7372 10051
rect 7406 10017 7444 10051
rect 7478 10017 9909 10051
rect 6442 9970 9909 10017
rect 6442 9936 7069 9970
rect 7103 9936 7147 9970
rect 7181 9936 7225 9970
rect 7259 9936 7372 9970
rect 7406 9936 7444 9970
rect 7478 9936 9909 9970
rect 6442 9889 9909 9936
rect 6442 9855 7069 9889
rect 7103 9855 7147 9889
rect 7181 9855 7225 9889
rect 7259 9855 7372 9889
rect 7406 9855 7444 9889
rect 7478 9855 9909 9889
rect 6442 9807 9909 9855
rect 6442 9773 7069 9807
rect 7103 9773 7147 9807
rect 7181 9773 7225 9807
rect 7259 9773 7372 9807
rect 7406 9773 7444 9807
rect 7478 9773 9909 9807
rect 6442 9725 9909 9773
rect 6442 9691 7069 9725
rect 7103 9691 7147 9725
rect 7181 9691 7225 9725
rect 7259 9691 7372 9725
rect 7406 9691 7444 9725
rect 7478 9691 9909 9725
rect 6442 9643 9909 9691
rect 6442 9609 7069 9643
rect 7103 9609 7147 9643
rect 7181 9609 7225 9643
rect 7259 9609 7372 9643
rect 7406 9609 7444 9643
rect 7478 9609 9909 9643
rect 6442 9598 9909 9609
rect 10029 10119 10033 10153
rect 10067 10119 10071 10153
rect 10029 10068 10071 10119
rect 10029 10034 10033 10068
rect 10067 10034 10071 10068
rect 10029 9983 10071 10034
rect 10029 9949 10033 9983
rect 10067 9949 10071 9983
rect 10029 9898 10071 9949
rect 10029 9864 10033 9898
rect 10067 9864 10071 9898
rect 10029 9812 10071 9864
rect 10029 9778 10033 9812
rect 10067 9778 10071 9812
rect 10029 9726 10071 9778
rect 10029 9692 10033 9726
rect 10067 9692 10071 9726
rect 10029 9640 10071 9692
rect 10029 9606 10033 9640
rect 10067 9606 10071 9640
rect 6318 9527 6322 9561
rect 6356 9527 6360 9561
rect 10029 9554 10071 9606
rect 6318 9475 6360 9527
rect 6488 9547 6504 9553
rect 6488 9519 6499 9547
rect 6538 9519 6573 9553
rect 6607 9519 6642 9553
rect 6676 9547 6711 9553
rect 6745 9547 6780 9553
rect 6814 9547 6849 9553
rect 6883 9547 6918 9553
rect 6952 9547 6987 9553
rect 7021 9547 7056 9553
rect 6681 9519 6711 9547
rect 6755 9519 6780 9547
rect 6829 9519 6849 9547
rect 6903 9519 6918 9547
rect 6977 9519 6987 9547
rect 7051 9519 7056 9547
rect 7090 9547 7125 9553
rect 7090 9519 7091 9547
rect 6533 9513 6573 9519
rect 6607 9513 6647 9519
rect 6681 9513 6721 9519
rect 6755 9513 6795 9519
rect 6829 9513 6869 9519
rect 6903 9513 6943 9519
rect 6977 9513 7017 9519
rect 7051 9513 7091 9519
rect 7159 9547 7194 9553
rect 7228 9547 7263 9553
rect 7297 9547 7332 9553
rect 7366 9547 7401 9553
rect 7435 9547 7470 9553
rect 7504 9547 7539 9553
rect 7159 9519 7165 9547
rect 7228 9519 7239 9547
rect 7297 9519 7313 9547
rect 7366 9519 7387 9547
rect 7435 9519 7461 9547
rect 7504 9519 7535 9547
rect 7573 9519 7608 9553
rect 7642 9547 7677 9553
rect 7711 9547 7746 9553
rect 7780 9547 7815 9553
rect 7849 9547 7884 9553
rect 7918 9547 7953 9553
rect 7987 9547 8022 9553
rect 8056 9547 8091 9553
rect 7643 9519 7677 9547
rect 7717 9519 7746 9547
rect 7791 9519 7815 9547
rect 7865 9519 7884 9547
rect 7939 9519 7953 9547
rect 8013 9519 8022 9547
rect 8087 9519 8091 9547
rect 8125 9547 8160 9553
rect 8194 9547 8229 9553
rect 8263 9547 8298 9553
rect 8332 9547 8367 9553
rect 8401 9547 8436 9553
rect 8470 9547 8505 9553
rect 8539 9547 8574 9553
rect 8608 9547 8643 9553
rect 8125 9519 8127 9547
rect 8194 9519 8201 9547
rect 8263 9519 8275 9547
rect 8332 9519 8349 9547
rect 8401 9519 8423 9547
rect 8470 9519 8496 9547
rect 8539 9519 8569 9547
rect 8608 9519 8642 9547
rect 8677 9519 8712 9553
rect 8746 9547 8781 9553
rect 8815 9547 8850 9553
rect 8884 9547 8918 9553
rect 8952 9547 8986 9553
rect 9020 9547 9054 9553
rect 9088 9547 9122 9553
rect 9156 9547 9190 9553
rect 8749 9519 8781 9547
rect 8822 9519 8850 9547
rect 8895 9519 8918 9547
rect 8968 9519 8986 9547
rect 9041 9519 9054 9547
rect 9114 9519 9122 9547
rect 9187 9519 9190 9547
rect 9224 9547 9258 9553
rect 9292 9547 9326 9553
rect 9360 9547 9394 9553
rect 9428 9547 9462 9553
rect 9496 9547 9530 9553
rect 9564 9547 9598 9553
rect 9632 9547 9666 9553
rect 9224 9519 9226 9547
rect 9292 9519 9299 9547
rect 9360 9519 9372 9547
rect 9428 9519 9445 9547
rect 9496 9519 9518 9547
rect 9564 9519 9591 9547
rect 9632 9519 9664 9547
rect 9700 9519 9734 9553
rect 9768 9547 9802 9553
rect 9836 9547 9852 9553
rect 9771 9519 9802 9547
rect 9844 9519 9852 9547
rect 10029 9520 10033 9554
rect 10067 9520 10071 9554
rect 7125 9513 7165 9519
rect 7199 9513 7239 9519
rect 7273 9513 7313 9519
rect 7347 9513 7387 9519
rect 7421 9513 7461 9519
rect 7495 9513 7535 9519
rect 7569 9513 7609 9519
rect 7643 9513 7683 9519
rect 7717 9513 7757 9519
rect 7791 9513 7831 9519
rect 7865 9513 7905 9519
rect 7939 9513 7979 9519
rect 8013 9513 8053 9519
rect 8087 9513 8127 9519
rect 8161 9513 8201 9519
rect 8235 9513 8275 9519
rect 8309 9513 8349 9519
rect 8383 9513 8423 9519
rect 8457 9513 8496 9519
rect 8530 9513 8569 9519
rect 8603 9513 8642 9519
rect 8676 9513 8715 9519
rect 8749 9513 8788 9519
rect 8822 9513 8861 9519
rect 8895 9513 8934 9519
rect 8968 9513 9007 9519
rect 9041 9513 9080 9519
rect 9114 9513 9153 9519
rect 9187 9513 9226 9519
rect 9260 9513 9299 9519
rect 9333 9513 9372 9519
rect 9406 9513 9445 9519
rect 9479 9513 9518 9519
rect 9552 9513 9591 9519
rect 9625 9513 9664 9519
rect 9698 9513 9737 9519
rect 9771 9513 9810 9519
rect 6318 9441 6322 9475
rect 6356 9441 6360 9475
rect 6318 9389 6360 9441
rect 10029 9468 10071 9520
rect 10029 9434 10033 9468
rect 10067 9434 10071 9468
rect 6318 9355 6322 9389
rect 6356 9355 6360 9389
rect 6318 9303 6360 9355
rect 6318 9269 6322 9303
rect 6356 9269 6360 9303
rect 6318 9217 6360 9269
rect 6318 9183 6322 9217
rect 6356 9183 6360 9217
rect 6318 9131 6360 9183
rect 6318 9097 6322 9131
rect 6356 9097 6360 9131
rect 6318 9045 6360 9097
rect 6318 9011 6322 9045
rect 6356 9011 6360 9045
rect 6318 8959 6360 9011
rect 6318 8925 6322 8959
rect 6356 8925 6360 8959
rect 6318 8873 6360 8925
rect 6318 8839 6322 8873
rect 6356 8839 6360 8873
rect 6442 9402 9909 9410
rect 6442 9368 7069 9402
rect 7103 9368 7147 9402
rect 7181 9368 7225 9402
rect 7259 9368 7372 9402
rect 7406 9368 7444 9402
rect 7478 9368 9909 9402
rect 6442 9321 9909 9368
rect 6442 9287 7069 9321
rect 7103 9287 7147 9321
rect 7181 9287 7225 9321
rect 7259 9287 7372 9321
rect 7406 9287 7444 9321
rect 7478 9287 9909 9321
rect 6442 9240 9909 9287
rect 6442 9206 7069 9240
rect 7103 9206 7147 9240
rect 7181 9206 7225 9240
rect 7259 9206 7372 9240
rect 7406 9206 7444 9240
rect 7478 9206 9909 9240
rect 6442 9159 9909 9206
rect 6442 9125 7069 9159
rect 7103 9125 7147 9159
rect 7181 9125 7225 9159
rect 7259 9125 7372 9159
rect 7406 9125 7444 9159
rect 7478 9125 9909 9159
rect 6442 9077 9909 9125
rect 6442 9043 7069 9077
rect 7103 9043 7147 9077
rect 7181 9043 7225 9077
rect 7259 9043 7372 9077
rect 7406 9043 7444 9077
rect 7478 9043 9909 9077
rect 6442 8995 9909 9043
rect 6442 8961 7069 8995
rect 7103 8961 7147 8995
rect 7181 8961 7225 8995
rect 7259 8961 7372 8995
rect 7406 8961 7444 8995
rect 7478 8961 9909 8995
rect 6442 8913 9909 8961
rect 6442 8879 7069 8913
rect 7103 8879 7147 8913
rect 7181 8879 7225 8913
rect 7259 8879 7372 8913
rect 7406 8879 7444 8913
rect 7478 8879 9909 8913
rect 6442 8868 9909 8879
rect 10029 9382 10071 9434
rect 10029 9348 10033 9382
rect 10067 9348 10071 9382
rect 10029 9296 10071 9348
rect 10029 9262 10033 9296
rect 10067 9262 10071 9296
rect 10029 9210 10071 9262
rect 10029 9176 10033 9210
rect 10067 9176 10071 9210
rect 10029 9124 10071 9176
rect 10029 9090 10033 9124
rect 10067 9090 10071 9124
rect 10029 9038 10071 9090
rect 10029 9004 10033 9038
rect 10067 9004 10071 9038
rect 10029 8952 10071 9004
rect 10029 8918 10033 8952
rect 10067 8918 10071 8952
rect 6318 8787 6360 8839
rect 6318 8753 6322 8787
rect 6356 8782 6360 8787
rect 10029 8866 10071 8918
rect 10029 8832 10033 8866
rect 10067 8832 10071 8866
rect 6356 8753 6443 8782
rect 10029 8753 10071 8832
rect 6318 8729 6443 8753
rect 6382 8077 6443 8729
rect 11979 8203 12071 8782
rect 8301 6695 8358 7356
rect 13718 7322 13781 8236
rect 8574 6945 13682 6946
rect 8574 6911 8608 6945
rect 8642 6911 8676 6945
rect 8710 6911 8744 6945
rect 8778 6911 8812 6945
rect 8846 6911 8880 6945
rect 8914 6911 8948 6945
rect 8982 6911 9016 6945
rect 9050 6911 9084 6945
rect 9118 6911 9152 6945
rect 9186 6911 9220 6945
rect 9254 6911 9288 6945
rect 9322 6911 9356 6945
rect 9390 6911 9424 6945
rect 9458 6911 9492 6945
rect 9526 6911 9560 6945
rect 9594 6911 9628 6945
rect 9662 6911 9696 6945
rect 9730 6911 9764 6945
rect 9798 6911 9832 6945
rect 9866 6911 9900 6945
rect 9934 6911 9968 6945
rect 10002 6911 10036 6945
rect 10070 6911 10104 6945
rect 10138 6911 10172 6945
rect 10206 6911 10240 6945
rect 10274 6911 10308 6945
rect 10342 6911 10376 6945
rect 10410 6911 10444 6945
rect 10478 6911 10512 6945
rect 10546 6911 10580 6945
rect 10614 6911 10648 6945
rect 10682 6911 10716 6945
rect 10750 6911 10784 6945
rect 10818 6911 10852 6945
rect 10886 6911 10920 6945
rect 10954 6911 10988 6945
rect 11022 6911 11056 6945
rect 11090 6911 11124 6945
rect 11158 6911 11192 6945
rect 11226 6911 11260 6945
rect 11294 6911 11328 6945
rect 11362 6911 11396 6945
rect 11430 6911 11464 6945
rect 11498 6911 11532 6945
rect 11566 6911 11600 6945
rect 11634 6911 11668 6945
rect 11702 6911 11736 6945
rect 11770 6911 11804 6945
rect 11838 6911 11872 6945
rect 11906 6911 11940 6945
rect 11974 6911 12008 6945
rect 12042 6911 12076 6945
rect 12110 6911 12144 6945
rect 12178 6911 12212 6945
rect 12246 6911 12280 6945
rect 12314 6911 12348 6945
rect 12382 6911 12416 6945
rect 12450 6911 12484 6945
rect 12518 6911 12552 6945
rect 12586 6911 12620 6945
rect 12654 6911 12688 6945
rect 12722 6911 12756 6945
rect 12790 6911 12824 6945
rect 12858 6911 12892 6945
rect 12926 6911 12960 6945
rect 12994 6911 13028 6945
rect 13062 6911 13096 6945
rect 13130 6911 13164 6945
rect 13198 6911 13232 6945
rect 13266 6911 13300 6945
rect 13334 6911 13368 6945
rect 13402 6911 13436 6945
rect 13470 6911 13504 6945
rect 13538 6911 13572 6945
rect 13606 6912 13682 6945
rect 13606 6911 13647 6912
rect 8574 6910 13647 6911
rect 8574 6877 8610 6910
rect 8574 6843 8575 6877
rect 8609 6843 8610 6877
rect 8574 6809 8610 6843
rect 8574 6775 8575 6809
rect 8609 6775 8610 6809
rect 8574 6741 8610 6775
rect 8574 6707 8575 6741
rect 8609 6707 8610 6741
rect 8574 6673 8610 6707
rect 8574 6639 8575 6673
rect 8609 6639 8610 6673
rect 8574 6605 8610 6639
rect 8574 6571 8575 6605
rect 8609 6571 8610 6605
rect 8574 6537 8610 6571
rect 8574 6503 8575 6537
rect 8609 6503 8610 6537
rect 8574 6469 8610 6503
rect 8574 6435 8575 6469
rect 8609 6435 8610 6469
rect 8574 6401 8610 6435
rect 8574 6367 8575 6401
rect 8609 6367 8610 6401
rect 8574 6333 8610 6367
rect 8574 6301 8575 6333
rect 4645 6300 8575 6301
rect 4645 6266 4679 6300
rect 4713 6266 4747 6300
rect 4781 6266 4815 6300
rect 4849 6266 4883 6300
rect 4917 6266 4951 6300
rect 4985 6266 5019 6300
rect 5053 6266 5087 6300
rect 5121 6266 5155 6300
rect 5189 6266 5223 6300
rect 5257 6266 5291 6300
rect 5325 6266 5359 6300
rect 5393 6266 5427 6300
rect 5461 6266 5495 6300
rect 5529 6266 5563 6300
rect 5597 6266 5631 6300
rect 5665 6266 5699 6300
rect 5733 6266 5767 6300
rect 5801 6266 5835 6300
rect 5869 6266 5903 6300
rect 5937 6266 5971 6300
rect 6005 6266 6039 6300
rect 6073 6266 6107 6300
rect 6141 6266 6175 6300
rect 6209 6266 6243 6300
rect 6277 6266 6311 6300
rect 6345 6266 6379 6300
rect 6413 6266 6447 6300
rect 6481 6266 6515 6300
rect 6549 6266 6583 6300
rect 6617 6266 6651 6300
rect 6685 6266 6719 6300
rect 6753 6266 6787 6300
rect 6821 6266 6855 6300
rect 6889 6266 6923 6300
rect 6957 6266 6991 6300
rect 7025 6266 7059 6300
rect 7093 6266 7127 6300
rect 7161 6266 7195 6300
rect 7229 6266 7263 6300
rect 7297 6266 7331 6300
rect 7365 6266 7399 6300
rect 7433 6266 7467 6300
rect 7501 6266 7535 6300
rect 7569 6266 7603 6300
rect 7637 6266 7671 6300
rect 7705 6266 7739 6300
rect 7773 6266 7807 6300
rect 7841 6266 7875 6300
rect 7909 6266 7943 6300
rect 7977 6266 8011 6300
rect 8045 6266 8079 6300
rect 8113 6266 8147 6300
rect 8181 6266 8215 6300
rect 8249 6266 8283 6300
rect 8317 6266 8351 6300
rect 8385 6266 8419 6300
rect 8453 6266 8487 6300
rect 8521 6299 8575 6300
rect 8609 6299 8610 6333
rect 8521 6266 8610 6299
rect 4645 6265 8610 6266
rect 13646 6878 13647 6910
rect 13681 6878 13682 6912
rect 13646 6844 13682 6878
rect 13646 6810 13647 6844
rect 13681 6810 13682 6844
rect 13646 6776 13682 6810
rect 13646 6742 13647 6776
rect 13681 6742 13682 6776
rect 13646 6708 13682 6742
rect 13646 6674 13647 6708
rect 13681 6674 13682 6708
rect 13646 6640 13682 6674
rect 13646 6606 13647 6640
rect 13681 6606 13682 6640
rect 13646 6572 13682 6606
rect 13646 6538 13647 6572
rect 13681 6538 13682 6572
rect 13646 6504 13682 6538
rect 13646 6470 13647 6504
rect 13681 6470 13682 6504
rect 13646 6436 13682 6470
rect 13646 6402 13647 6436
rect 13681 6402 13682 6436
rect 13646 6368 13682 6402
rect 13646 6334 13647 6368
rect 13681 6334 13682 6368
rect 13646 6300 13682 6334
rect 13646 6266 13647 6300
rect 13681 6266 13682 6300
rect 249 6254 813 6255
rect 249 6220 283 6254
rect 317 6220 351 6254
rect 385 6220 419 6254
rect 453 6220 487 6254
rect 521 6220 555 6254
rect 589 6220 623 6254
rect 657 6220 691 6254
rect 725 6221 813 6254
rect 725 6220 778 6221
rect 249 6219 778 6220
rect 249 6147 285 6219
rect 249 6105 250 6147
rect 284 6105 285 6147
rect 249 6071 285 6105
rect 777 6187 778 6219
rect 812 6187 813 6221
rect 777 6153 813 6187
rect 777 6113 778 6153
rect 812 6113 813 6153
rect 249 6007 250 6071
rect 284 6007 285 6071
rect 249 6003 285 6007
rect 249 5901 250 6003
rect 284 5901 285 6003
rect 249 5887 285 5901
rect 249 5833 250 5887
rect 284 5833 285 5887
rect 249 5804 285 5833
rect 249 5765 250 5804
rect 284 5765 285 5804
rect 249 5731 285 5765
rect 249 5687 250 5731
rect 284 5687 285 5731
rect 249 5663 285 5687
rect 249 5604 250 5663
rect 284 5604 285 5663
rect 249 5595 285 5604
rect 249 5561 250 5595
rect 284 5561 285 5595
rect 249 5555 285 5561
rect 249 5493 250 5555
rect 284 5493 285 5555
rect 249 5472 285 5493
rect 249 5425 250 5472
rect 284 5425 285 5472
rect 693 6076 727 6092
rect 693 6004 727 6042
rect 693 5932 727 5970
rect 693 5881 727 5898
rect 693 5809 727 5825
rect 693 5737 727 5752
rect 693 5665 727 5679
rect 693 5593 727 5606
rect 693 5521 727 5533
rect 693 5444 727 5460
rect 777 6085 813 6113
rect 777 6027 778 6085
rect 812 6027 813 6085
rect 777 6017 813 6027
rect 777 5983 778 6017
rect 812 5983 813 6017
rect 777 5949 813 5983
rect 777 5915 778 5949
rect 812 5915 813 5949
rect 777 5881 813 5915
rect 777 5847 778 5881
rect 812 5847 813 5881
rect 777 5813 813 5847
rect 777 5752 778 5813
rect 812 5752 813 5813
rect 777 5745 813 5752
rect 777 5711 778 5745
rect 812 5711 813 5745
rect 777 5691 813 5711
rect 777 5643 778 5691
rect 812 5643 813 5691
rect 777 5609 813 5643
rect 777 5575 778 5609
rect 812 5575 813 5609
rect 777 5541 813 5575
rect 777 5492 778 5541
rect 812 5492 813 5541
rect 777 5473 813 5492
rect 249 5391 285 5425
rect 249 5357 250 5391
rect 284 5357 285 5391
rect 777 5439 778 5473
rect 812 5439 813 5473
rect 777 5420 813 5439
rect 249 5323 285 5357
rect 249 5289 250 5323
rect 284 5289 285 5323
rect 249 5255 285 5289
rect 249 5221 250 5255
rect 284 5221 285 5255
rect 249 5187 285 5221
rect 249 5153 250 5187
rect 284 5153 285 5187
rect 249 5119 285 5153
rect 249 5061 250 5119
rect 284 5061 285 5119
rect 249 5051 285 5061
rect 249 4949 250 5051
rect 284 4949 285 5051
rect 335 5372 369 5388
rect 335 5295 369 5338
rect 335 5218 369 5261
rect 335 5142 369 5184
rect 335 5107 369 5108
rect 335 5035 369 5073
rect 777 5371 778 5420
rect 812 5371 813 5420
rect 777 5337 813 5371
rect 777 5281 778 5337
rect 812 5281 813 5337
rect 777 5269 813 5281
rect 777 5235 778 5269
rect 812 5235 813 5269
rect 777 5201 813 5235
rect 777 5167 778 5201
rect 812 5167 813 5201
rect 777 5133 813 5167
rect 777 5099 778 5133
rect 812 5099 813 5133
rect 777 5065 813 5099
rect 777 5031 778 5065
rect 812 5031 813 5065
rect 249 4939 285 4949
rect 249 4881 250 4939
rect 284 4881 285 4939
rect 777 4997 813 5031
rect 777 4963 778 4997
rect 812 4963 813 4997
rect 777 4929 813 4963
rect 249 4861 285 4881
rect 249 4813 250 4861
rect 284 4813 285 4861
rect 249 4782 285 4813
rect 249 4745 250 4782
rect 284 4745 285 4782
rect 693 4910 727 4926
rect 693 4842 727 4853
rect 777 4895 778 4929
rect 812 4895 813 4929
rect 777 4861 813 4895
rect 777 4827 778 4861
rect 812 4827 813 4861
rect 777 4803 813 4827
rect 249 4711 285 4745
rect 249 4669 250 4711
rect 284 4669 285 4711
rect 249 4643 285 4669
rect 249 4590 250 4643
rect 284 4590 285 4643
rect 335 4756 369 4770
rect 335 4686 369 4720
rect 335 4636 369 4650
rect 777 4759 778 4803
rect 812 4759 813 4803
rect 777 4729 813 4759
rect 777 4691 778 4729
rect 812 4691 813 4729
rect 777 4655 813 4691
rect 249 4575 285 4590
rect 249 4511 250 4575
rect 284 4543 285 4575
rect 777 4621 778 4655
rect 812 4621 813 4655
rect 777 4543 813 4621
rect 284 4542 813 4543
rect 284 4511 337 4542
rect 249 4508 337 4511
rect 371 4508 405 4542
rect 449 4508 473 4542
rect 530 4508 541 4542
rect 575 4508 577 4542
rect 643 4508 658 4542
rect 711 4508 740 4542
rect 779 4508 813 4542
rect 249 4507 813 4508
rect 966 6254 1515 6255
rect 966 6220 1000 6254
rect 1034 6220 1068 6254
rect 1102 6220 1136 6254
rect 1170 6220 1204 6254
rect 1238 6220 1272 6254
rect 1306 6220 1340 6254
rect 1374 6220 1408 6254
rect 1442 6221 1515 6254
rect 1442 6220 1480 6221
rect 966 6219 1480 6220
rect 966 6144 1002 6219
rect 966 6102 967 6144
rect 1001 6102 1002 6144
rect 966 6068 1002 6102
rect 1479 6187 1480 6219
rect 1514 6187 1515 6221
rect 1479 6153 1515 6187
rect 1479 6110 1480 6153
rect 1514 6110 1515 6153
rect 966 6022 967 6068
rect 1001 6022 1002 6068
rect 966 6000 1002 6022
rect 966 5966 967 6000
rect 1001 5966 1002 6000
rect 966 5932 1002 5966
rect 966 5898 967 5932
rect 1001 5898 1002 5932
rect 966 5881 1002 5898
rect 966 5830 967 5881
rect 1001 5830 1002 5881
rect 966 5796 1002 5830
rect 966 5752 967 5796
rect 1001 5752 1002 5796
rect 1052 6076 1086 6092
rect 1052 5999 1086 6042
rect 1052 5922 1086 5965
rect 1052 5881 1086 5888
rect 1052 5846 1086 5847
rect 1052 5809 1086 5812
rect 1479 6085 1515 6110
rect 1479 6035 1480 6085
rect 1514 6035 1515 6085
rect 1479 6017 1515 6035
rect 1479 5960 1480 6017
rect 1514 5960 1515 6017
rect 1479 5949 1515 5960
rect 1479 5885 1480 5949
rect 1514 5885 1515 5949
rect 1479 5881 1515 5885
rect 1479 5847 1480 5881
rect 1514 5847 1515 5881
rect 1479 5843 1515 5847
rect 1479 5779 1480 5843
rect 1514 5779 1515 5843
rect 966 5728 1002 5752
rect 1479 5767 1515 5779
rect 966 5694 967 5728
rect 1001 5694 1002 5728
rect 966 5691 1002 5694
rect 966 5626 967 5691
rect 1001 5626 1002 5691
rect 966 5592 1002 5626
rect 966 5558 967 5592
rect 1001 5558 1002 5592
rect 966 5524 1002 5558
rect 966 5490 967 5524
rect 1001 5490 1002 5524
rect 966 5456 1002 5490
rect 1052 5724 1086 5740
rect 1052 5656 1086 5690
rect 1052 5522 1086 5622
rect 1479 5711 1480 5767
rect 1514 5711 1515 5767
rect 1479 5691 1515 5711
rect 1479 5643 1480 5691
rect 1514 5643 1515 5691
rect 1479 5615 1515 5643
rect 1479 5575 1480 5615
rect 1514 5575 1515 5615
rect 1479 5541 1515 5575
rect 1052 5488 1340 5522
rect 966 5413 967 5456
rect 1001 5413 1002 5456
rect 1206 5461 1340 5488
rect 966 5388 1002 5413
rect 966 5323 967 5388
rect 1001 5323 1002 5388
rect 966 5320 1002 5323
rect 966 5286 967 5320
rect 1001 5286 1002 5320
rect 966 5267 1002 5286
rect 966 5218 967 5267
rect 1001 5218 1002 5267
rect 1089 5438 1160 5454
rect 1123 5404 1160 5438
rect 1206 5427 1220 5461
rect 1254 5427 1292 5461
rect 1326 5427 1340 5461
rect 1479 5507 1480 5541
rect 1514 5507 1515 5541
rect 1479 5473 1515 5507
rect 4645 6221 4681 6265
rect 4645 6187 4646 6221
rect 4680 6187 4681 6221
rect 4645 6153 4681 6187
rect 4645 6119 4646 6153
rect 4680 6119 4681 6153
rect 4645 6085 4681 6119
rect 4645 6051 4646 6085
rect 4680 6051 4681 6085
rect 4645 6017 4681 6051
rect 4645 5983 4646 6017
rect 4680 5983 4681 6017
rect 4645 5949 4681 5983
rect 4645 5915 4646 5949
rect 4680 5915 4681 5949
rect 4645 5881 4681 5915
rect 4645 5847 4646 5881
rect 4680 5847 4681 5881
rect 4645 5813 4681 5847
rect 4645 5779 4646 5813
rect 4680 5779 4681 5813
rect 4645 5745 4681 5779
rect 4645 5711 4646 5745
rect 4680 5711 4681 5745
rect 4645 5677 4681 5711
rect 4645 5643 4646 5677
rect 4680 5643 4681 5677
rect 4645 5609 4681 5643
rect 4645 5575 4646 5609
rect 4680 5575 4681 5609
rect 4645 5541 4681 5575
rect 4645 5507 4646 5541
rect 4680 5507 4681 5541
rect 1089 5304 1160 5404
rect 1123 5290 1160 5304
rect 1123 5270 1126 5290
rect 1089 5256 1126 5270
rect 1089 5254 1160 5256
rect 966 5184 1002 5218
rect 1126 5218 1160 5254
rect 966 5144 967 5184
rect 1001 5144 1002 5184
rect 966 5116 1002 5144
rect 966 5055 967 5116
rect 1001 5055 1002 5116
rect 966 5048 1002 5055
rect 966 5014 967 5048
rect 1001 5014 1002 5048
rect 966 4980 1002 5014
rect 1052 5182 1092 5198
rect 1479 5417 1480 5473
rect 1514 5417 1515 5473
rect 1479 5405 1515 5417
rect 1479 5344 1480 5405
rect 1514 5344 1515 5405
rect 3972 5381 4200 5483
rect 1479 5337 1515 5344
rect 1479 5271 1480 5337
rect 1514 5271 1515 5337
rect 1479 5269 1515 5271
rect 1479 5235 1480 5269
rect 1514 5235 1515 5269
rect 1479 5232 1515 5235
rect 1052 5151 1058 5182
rect 1086 5117 1092 5148
rect 1052 5079 1092 5117
rect 1086 5048 1092 5079
rect 1052 5014 1058 5045
rect 1052 4998 1092 5014
rect 1479 5167 1480 5232
rect 1514 5167 1515 5232
rect 1479 5159 1515 5167
rect 3268 5357 4200 5381
rect 3268 5355 4137 5357
rect 3268 5352 4069 5355
rect 3268 5318 3292 5352
rect 3326 5318 3362 5352
rect 3396 5318 3433 5352
rect 3467 5318 3504 5352
rect 3538 5318 3575 5352
rect 3609 5318 3646 5352
rect 3680 5318 3717 5352
rect 3751 5318 3788 5352
rect 3822 5318 3859 5352
rect 3893 5318 3930 5352
rect 3964 5318 4001 5352
rect 4035 5321 4069 5352
rect 4103 5323 4137 5355
rect 4171 5323 4200 5357
rect 4103 5321 4200 5323
rect 4035 5318 4200 5321
rect 3268 5289 4200 5318
rect 3268 5284 4137 5289
rect 3268 5250 3292 5284
rect 3326 5250 3362 5284
rect 3396 5250 3432 5284
rect 3466 5250 3502 5284
rect 3536 5250 3572 5284
rect 3606 5250 3643 5284
rect 3677 5250 3714 5284
rect 3748 5250 3785 5284
rect 3819 5250 3856 5284
rect 3890 5250 3927 5284
rect 3961 5250 3998 5284
rect 4032 5250 4069 5284
rect 4103 5255 4137 5284
rect 4171 5255 4200 5289
rect 4103 5250 4200 5255
rect 3268 5244 4200 5250
rect 3268 5216 3744 5244
rect 3778 5216 3816 5244
rect 3268 5182 3292 5216
rect 3326 5182 3362 5216
rect 3396 5182 3432 5216
rect 3466 5182 3502 5216
rect 3536 5182 3572 5216
rect 3606 5182 3642 5216
rect 3676 5182 3712 5216
rect 3778 5210 3782 5216
rect 3746 5182 3782 5210
rect 3850 5216 3888 5244
rect 3850 5210 3852 5216
rect 3816 5182 3852 5210
rect 3886 5210 3888 5216
rect 3922 5216 3960 5244
rect 3994 5216 4032 5244
rect 4066 5216 4104 5244
rect 4138 5216 4200 5244
rect 3886 5182 3922 5210
rect 3956 5210 3960 5216
rect 4026 5210 4032 5216
rect 4096 5210 4104 5216
rect 3956 5182 3992 5210
rect 4026 5182 4062 5210
rect 4096 5182 4132 5210
rect 4166 5182 4200 5216
rect 1479 5099 1480 5159
rect 1514 5099 1515 5159
rect 1479 5086 1515 5099
rect 1479 5031 1480 5086
rect 1514 5031 1515 5086
rect 1479 5013 1515 5031
rect 966 4946 967 4980
rect 1001 4946 1002 4980
rect 966 4912 1002 4946
rect 966 4878 967 4912
rect 1001 4878 1002 4912
rect 966 4844 1002 4878
rect 966 4810 967 4844
rect 1001 4810 1002 4844
rect 1479 4963 1480 5013
rect 1514 4963 1515 5013
rect 1479 4940 1515 4963
rect 1479 4895 1480 4940
rect 1514 4895 1515 4940
rect 1479 4867 1515 4895
rect 966 4776 1002 4810
rect 966 4742 967 4776
rect 1001 4742 1002 4776
rect 966 4708 1002 4742
rect 966 4674 967 4708
rect 1001 4674 1002 4708
rect 966 4640 1002 4674
rect 966 4601 967 4640
rect 1001 4601 1002 4640
rect 966 4572 1002 4601
rect 966 4524 967 4572
rect 1001 4524 1002 4572
rect 966 4504 1002 4524
rect 966 4447 967 4504
rect 1001 4447 1002 4504
rect 966 4436 1002 4447
rect 966 4371 967 4436
rect 1001 4371 1002 4436
rect 966 4368 1002 4371
rect 966 4334 967 4368
rect 1001 4334 1002 4368
rect 966 4329 1002 4334
rect 249 4311 813 4312
rect 249 4277 250 4311
rect 317 4277 351 4311
rect 385 4277 415 4311
rect 453 4277 487 4311
rect 530 4277 555 4311
rect 611 4277 623 4311
rect 657 4277 658 4311
rect 725 4277 740 4311
rect 774 4278 813 4311
rect 774 4277 778 4278
rect 249 4276 778 4277
rect 249 4242 285 4276
rect 249 4199 250 4242
rect 284 4199 285 4242
rect 249 4174 285 4199
rect 249 4121 250 4174
rect 284 4121 285 4174
rect 777 4244 778 4276
rect 812 4244 813 4278
rect 777 4210 813 4244
rect 777 4176 778 4210
rect 812 4176 813 4210
rect 249 4106 285 4121
rect 249 4044 250 4106
rect 284 4044 285 4106
rect 249 4038 285 4044
rect 249 4004 250 4038
rect 284 4004 285 4038
rect 249 4001 285 4004
rect 249 3936 250 4001
rect 284 3936 285 4001
rect 249 3924 285 3936
rect 249 3868 250 3924
rect 284 3868 285 3924
rect 249 3847 285 3868
rect 249 3800 250 3847
rect 284 3800 285 3847
rect 249 3770 285 3800
rect 249 3732 250 3770
rect 284 3732 285 3770
rect 249 3698 285 3732
rect 351 4133 385 4149
rect 351 4051 385 4099
rect 351 3970 385 4017
rect 351 3889 385 3936
rect 351 3808 385 3855
rect 351 3727 385 3774
rect 14 3664 48 3694
rect 351 3664 385 3693
rect 14 3656 385 3664
rect 48 3622 385 3656
rect 14 3610 385 3622
rect 777 4142 813 4176
rect 777 4108 778 4142
rect 812 4108 813 4142
rect 777 4089 813 4108
rect 777 4040 778 4089
rect 812 4040 813 4089
rect 777 4006 813 4040
rect 777 3969 778 4006
rect 812 3969 813 4006
rect 777 3938 813 3969
rect 777 3883 778 3938
rect 812 3883 813 3938
rect 777 3870 813 3883
rect 777 3836 778 3870
rect 812 3836 813 3870
rect 777 3831 813 3836
rect 777 3768 778 3831
rect 812 3768 813 3831
rect 777 3746 813 3768
rect 777 3700 778 3746
rect 812 3700 813 3746
rect 777 3666 813 3700
rect 777 3632 778 3666
rect 812 3632 813 3666
rect 249 3550 285 3576
rect 777 3550 813 3632
rect 249 3549 813 3550
rect 249 3515 337 3549
rect 371 3515 399 3549
rect 439 3515 473 3549
rect 507 3515 541 3549
rect 581 3515 609 3549
rect 655 3515 677 3549
rect 729 3515 745 3549
rect 779 3515 813 3549
rect 249 3514 813 3515
rect 966 4266 967 4329
rect 1001 4266 1002 4329
rect 966 4253 1002 4266
rect 966 4198 967 4253
rect 1001 4198 1002 4253
rect 966 4164 1002 4198
rect 966 4130 967 4164
rect 1001 4130 1002 4164
rect 966 4096 1002 4130
rect 966 4062 967 4096
rect 1001 4062 1002 4096
rect 966 4028 1002 4062
rect 966 3994 967 4028
rect 1001 3994 1002 4028
rect 966 3960 1002 3994
rect 966 3926 967 3960
rect 1001 3926 1002 3960
rect 966 3892 1002 3926
rect 1052 4816 1086 4832
rect 1052 4747 1086 4759
rect 1052 4678 1086 4687
rect 1052 4609 1086 4644
rect 1052 4540 1086 4575
rect 1052 4471 1086 4506
rect 1052 4402 1086 4437
rect 1052 4334 1086 4368
rect 1052 4266 1086 4300
rect 1052 4198 1086 4232
rect 1052 4130 1086 4164
rect 1052 4089 1086 4096
rect 1052 4017 1086 4028
rect 1052 3921 1086 3960
rect 1479 4827 1480 4867
rect 1514 4827 1515 4867
rect 1479 4794 1515 4827
rect 1479 4759 1480 4794
rect 1514 4759 1515 4794
rect 1479 4725 1515 4759
rect 1479 4687 1480 4725
rect 1514 4687 1515 4725
rect 1479 4657 1515 4687
rect 1479 4614 1480 4657
rect 1514 4614 1515 4657
rect 1479 4589 1515 4614
rect 1479 4541 1480 4589
rect 1514 4541 1515 4589
rect 1479 4521 1515 4541
rect 1479 4468 1480 4521
rect 1514 4468 1515 4521
rect 1479 4453 1515 4468
rect 1479 4395 1480 4453
rect 1514 4395 1515 4453
rect 1479 4385 1515 4395
rect 1479 4322 1480 4385
rect 1514 4322 1515 4385
rect 1479 4317 1515 4322
rect 1479 4215 1480 4317
rect 1514 4215 1515 4317
rect 1479 4210 1515 4215
rect 1479 4147 1480 4210
rect 1514 4147 1515 4210
rect 1479 4137 1515 4147
rect 1479 4079 1480 4137
rect 1514 4079 1515 4137
rect 1479 4064 1515 4079
rect 1479 4011 1480 4064
rect 1514 4011 1515 4064
rect 1479 3991 1515 4011
rect 1479 3943 1480 3991
rect 1514 3943 1515 3991
rect 966 3825 967 3892
rect 1001 3825 1002 3892
rect 966 3824 1002 3825
rect 966 3790 967 3824
rect 1001 3790 1002 3824
rect 966 3785 1002 3790
rect 966 3722 967 3785
rect 1001 3722 1002 3785
rect 1479 3918 1515 3943
rect 1479 3875 1480 3918
rect 1514 3875 1515 3918
rect 1479 3845 1515 3875
rect 1479 3807 1480 3845
rect 1514 3807 1515 3845
rect 1479 3773 1515 3807
rect 966 3711 1002 3722
rect 966 3654 967 3711
rect 1001 3654 1002 3711
rect 966 3638 1002 3654
rect 966 3586 967 3638
rect 1001 3586 1002 3638
rect 966 3565 1002 3586
rect 966 3518 967 3565
rect 1001 3518 1002 3565
rect 966 3492 1002 3518
rect 966 3450 967 3492
rect 1001 3450 1002 3492
rect 1052 3738 1086 3754
rect 1479 3738 1480 3773
rect 1514 3738 1515 3773
rect 1052 3664 1086 3694
rect 1196 3679 1234 3713
rect 1268 3679 1306 3713
rect 1479 3705 1515 3738
rect 1052 3590 1086 3622
rect 1052 3516 1086 3550
rect 1479 3665 1480 3705
rect 1514 3665 1515 3705
rect 1479 3637 1515 3665
rect 1479 3592 1480 3637
rect 1514 3592 1515 3637
rect 1479 3569 1515 3592
rect 1196 3501 1234 3535
rect 1268 3501 1306 3535
rect 1479 3519 1480 3569
rect 1514 3519 1515 3569
rect 1479 3501 1515 3519
rect 1052 3466 1086 3478
rect 966 3416 1002 3450
rect 966 3382 967 3416
rect 1001 3382 1002 3416
rect 249 3360 813 3361
rect 249 3326 283 3360
rect 317 3326 351 3360
rect 385 3338 419 3360
rect 453 3338 555 3360
rect 589 3338 623 3360
rect 657 3338 691 3360
rect 725 3338 813 3360
rect 966 3348 1002 3382
rect 1479 3446 1480 3501
rect 1514 3446 1515 3501
rect 1479 3433 1515 3446
rect 1479 3373 1480 3433
rect 1514 3373 1515 3433
rect 1479 3365 1515 3373
rect 406 3326 419 3338
rect 249 3304 372 3326
rect 406 3304 450 3326
rect 484 3304 528 3338
rect 589 3326 606 3338
rect 657 3326 684 3338
rect 725 3326 762 3338
rect 796 3327 813 3338
rect 562 3304 606 3326
rect 640 3304 684 3326
rect 718 3304 762 3326
rect 249 3300 285 3304
rect 249 3256 250 3300
rect 284 3256 285 3300
rect 249 3222 285 3256
rect 249 3187 250 3222
rect 284 3187 285 3222
rect 777 3293 778 3304
rect 812 3293 813 3327
rect 1052 3336 1086 3352
rect 777 3259 813 3293
rect 777 3225 778 3259
rect 812 3225 813 3259
rect 249 3154 285 3187
rect 249 3108 250 3154
rect 284 3108 285 3154
rect 249 3086 285 3108
rect 249 3030 250 3086
rect 284 3030 285 3086
rect 249 3018 285 3030
rect 349 3182 383 3198
rect 349 3114 383 3148
rect 777 3191 813 3225
rect 1012 3302 1052 3314
rect 1012 3280 1086 3302
rect 978 3268 1086 3280
rect 978 3242 1052 3268
rect 1012 3234 1052 3242
rect 1012 3208 1086 3234
rect 1479 3299 1480 3365
rect 1514 3299 1515 3365
rect 1479 3297 1515 3299
rect 1479 3263 1480 3297
rect 1514 3263 1515 3297
rect 1479 3259 1515 3263
rect 777 3157 778 3191
rect 812 3157 813 3191
rect 1479 3195 1480 3259
rect 1514 3195 1515 3259
rect 1479 3185 1515 3195
rect 777 3123 813 3157
rect 349 3041 383 3080
rect 693 3078 727 3094
rect 349 3007 441 3041
rect 693 3010 727 3044
rect 249 2904 283 2939
rect 249 2901 369 2904
rect 283 2888 369 2901
rect 283 2867 335 2888
rect 249 2787 285 2824
rect 267 2779 285 2787
rect 233 2745 250 2753
rect 284 2745 285 2779
rect 233 2714 285 2745
rect 267 2711 285 2714
rect 233 2677 250 2680
rect 284 2677 285 2711
rect 335 2811 369 2854
rect 475 2823 513 2857
rect 335 2734 369 2777
rect 693 2797 727 2976
rect 547 2731 585 2765
rect 335 2684 369 2700
rect 693 2725 727 2763
rect 777 3089 778 3123
rect 812 3089 813 3123
rect 777 3055 813 3089
rect 777 3021 778 3055
rect 812 3021 813 3055
rect 777 2987 813 3021
rect 777 2953 778 2987
rect 812 2953 813 2987
rect 777 2919 813 2953
rect 777 2885 778 2919
rect 812 2885 813 2919
rect 777 2851 813 2885
rect 777 2817 778 2851
rect 812 2817 813 2851
rect 777 2783 813 2817
rect 777 2749 778 2783
rect 812 2749 813 2783
rect 777 2715 813 2749
rect 233 2643 285 2677
rect 233 2641 250 2643
rect 284 2609 285 2643
rect 267 2607 285 2609
rect 249 2575 285 2607
rect 249 2541 250 2575
rect 284 2541 285 2575
rect 777 2680 778 2715
rect 812 2680 813 2715
rect 777 2647 813 2680
rect 777 2603 778 2647
rect 812 2603 813 2647
rect 777 2579 813 2603
rect 249 2507 285 2541
rect 249 2473 250 2507
rect 284 2473 285 2507
rect 249 2439 285 2473
rect 249 2405 250 2439
rect 284 2405 285 2439
rect 249 2371 285 2405
rect 249 2337 250 2371
rect 284 2337 285 2371
rect 249 2324 285 2337
rect 267 2303 285 2324
rect 233 2269 250 2290
rect 284 2269 285 2303
rect 233 2235 285 2269
rect 233 2234 250 2235
rect 284 2201 285 2235
rect 363 2529 513 2545
rect 547 2529 585 2563
rect 619 2529 643 2545
rect 363 2511 643 2529
rect 693 2536 727 2552
rect 363 2346 397 2511
rect 363 2278 397 2312
rect 693 2468 727 2502
rect 693 2269 727 2434
rect 363 2228 397 2244
rect 441 2235 727 2269
rect 777 2526 778 2579
rect 812 2526 813 2579
rect 777 2511 813 2526
rect 777 2449 778 2511
rect 812 2449 813 2511
rect 777 2443 813 2449
rect 777 2409 778 2443
rect 812 2409 813 2443
rect 777 2407 813 2409
rect 777 2341 778 2407
rect 812 2341 813 2407
rect 777 2331 813 2341
rect 777 2273 778 2331
rect 812 2273 813 2331
rect 267 2200 285 2201
rect 233 2167 285 2200
rect 233 2145 250 2167
rect 284 2135 285 2167
rect 777 2135 813 2273
rect 284 2134 813 2135
rect 284 2133 333 2134
rect 267 2111 333 2133
rect 249 2100 333 2111
rect 371 2100 405 2134
rect 448 2100 473 2134
rect 529 2100 541 2134
rect 575 2100 576 2134
rect 643 2100 658 2134
rect 711 2100 740 2134
rect 779 2100 813 2134
rect 249 2099 813 2100
rect 966 3122 1002 3174
rect 966 3088 967 3122
rect 1001 3088 1002 3122
rect 966 3054 1002 3088
rect 1386 3146 1420 3162
rect 1386 3078 1420 3112
rect 966 3020 967 3054
rect 1001 3020 1002 3054
rect 966 2986 1002 3020
rect 966 2952 967 2986
rect 1001 2952 1002 2986
rect 966 2919 1002 2952
rect 966 2884 967 2919
rect 1001 2884 1002 2919
rect 966 2850 1002 2884
rect 966 2816 967 2850
rect 1001 2816 1002 2850
rect 966 2782 1002 2816
rect 966 2748 967 2782
rect 1001 2748 1002 2782
rect 966 2714 1002 2748
rect 966 2680 967 2714
rect 1001 2680 1002 2714
rect 1052 3042 1086 3058
rect 1052 2974 1086 3008
rect 1386 3005 1420 3044
rect 1340 2971 1420 3005
rect 1479 3127 1480 3185
rect 1514 3127 1515 3185
rect 1479 3111 1515 3127
rect 1479 3059 1480 3111
rect 1514 3059 1515 3111
rect 1479 3037 1515 3059
rect 1479 2991 1480 3037
rect 1514 2991 1515 3037
rect 1052 2797 1086 2940
rect 1052 2725 1086 2763
rect 1479 2963 1515 2991
rect 1479 2923 1480 2963
rect 1514 2923 1515 2963
rect 1479 2889 1515 2923
rect 1479 2855 1480 2889
rect 1514 2855 1515 2889
rect 1479 2821 1515 2855
rect 1479 2787 1480 2821
rect 1514 2787 1515 2821
rect 1386 2742 1420 2758
rect 966 2646 1002 2680
rect 966 2605 967 2646
rect 1001 2605 1002 2646
rect 966 2578 1002 2605
rect 966 2530 967 2578
rect 1001 2530 1002 2578
rect 1386 2665 1420 2703
rect 1386 2593 1420 2631
rect 966 2510 1002 2530
rect 966 2455 967 2510
rect 1001 2455 1002 2510
rect 966 2442 1002 2455
rect 966 2380 967 2442
rect 1001 2380 1002 2442
rect 966 2374 1002 2380
rect 966 2340 967 2374
rect 1001 2340 1002 2374
rect 966 2339 1002 2340
rect 966 2272 967 2339
rect 1001 2272 1002 2339
rect 966 2238 1002 2272
rect 966 2204 967 2238
rect 1001 2204 1002 2238
rect 966 2170 1002 2204
rect 966 2136 967 2170
rect 1001 2136 1002 2170
rect 966 2102 1002 2136
rect 966 2068 967 2102
rect 1001 2068 1002 2102
rect 1386 2538 1420 2554
rect 1479 2753 1515 2787
rect 1479 2719 1480 2753
rect 1514 2719 1515 2753
rect 1479 2685 1515 2719
rect 1479 2647 1480 2685
rect 1514 2647 1515 2685
rect 1479 2617 1515 2647
rect 1479 2583 1480 2617
rect 1514 2583 1515 2617
rect 1479 2568 1515 2583
rect 1052 2492 1086 2530
rect 1479 2515 1480 2568
rect 1514 2515 1515 2568
rect 1052 2190 1086 2458
rect 1386 2466 1420 2482
rect 1386 2389 1420 2427
rect 1386 2312 1420 2355
rect 1386 2262 1420 2278
rect 1479 2481 1515 2515
rect 1479 2447 1480 2481
rect 1514 2447 1515 2481
rect 1479 2413 1515 2447
rect 1479 2359 1480 2413
rect 1514 2359 1515 2413
rect 1479 2345 1515 2359
rect 1479 2285 1480 2345
rect 1514 2285 1515 2345
rect 1479 2277 1515 2285
rect 1052 2122 1086 2156
rect 1052 2072 1086 2088
rect 1479 2211 1480 2277
rect 1514 2211 1515 2277
rect 1479 2209 1515 2211
rect 1479 2175 1480 2209
rect 1514 2175 1515 2209
rect 1479 2171 1515 2175
rect 1479 2107 1480 2171
rect 1514 2107 1515 2171
rect 1479 2097 1515 2107
rect 966 2034 1002 2068
rect 966 2000 967 2034
rect 1001 2000 1002 2034
rect 966 1966 1002 2000
rect 249 1945 345 1946
rect 379 1945 423 1946
rect 457 1945 501 1946
rect 535 1945 579 1946
rect 613 1945 657 1946
rect 249 1911 283 1945
rect 317 1912 345 1945
rect 317 1911 351 1912
rect 385 1911 419 1945
rect 457 1912 487 1945
rect 535 1912 555 1945
rect 613 1912 623 1945
rect 453 1911 487 1912
rect 521 1911 555 1912
rect 589 1911 623 1912
rect 691 1945 813 1946
rect 657 1911 691 1912
rect 725 1912 813 1945
rect 725 1911 778 1912
rect 249 1910 778 1911
rect 249 1830 285 1910
rect 249 1796 250 1830
rect 284 1796 285 1830
rect 777 1874 778 1910
rect 812 1874 813 1912
rect 777 1844 813 1874
rect 249 1762 285 1796
rect 249 1696 250 1762
rect 284 1696 285 1762
rect 249 1694 285 1696
rect 249 1660 250 1694
rect 284 1660 285 1694
rect 249 1657 285 1660
rect 249 1592 250 1657
rect 284 1592 285 1657
rect 249 1584 285 1592
rect 249 1524 250 1584
rect 284 1524 285 1584
rect 249 1511 285 1524
rect 249 1456 250 1511
rect 284 1456 285 1511
rect 249 1438 285 1456
rect 249 1388 250 1438
rect 284 1388 285 1438
rect 249 1365 285 1388
rect 249 1320 250 1365
rect 284 1320 285 1365
rect 249 1292 285 1320
rect 349 1767 383 1770
rect 349 1732 383 1733
rect 349 1685 383 1698
rect 349 1604 383 1651
rect 349 1523 383 1570
rect 349 1442 383 1489
rect 349 1361 383 1408
rect 349 1311 383 1327
rect 777 1791 778 1844
rect 812 1791 813 1844
rect 777 1776 813 1791
rect 777 1709 778 1776
rect 812 1709 813 1776
rect 777 1708 813 1709
rect 777 1674 778 1708
rect 812 1674 813 1708
rect 777 1661 813 1674
rect 777 1606 778 1661
rect 812 1606 813 1661
rect 777 1579 813 1606
rect 777 1538 778 1579
rect 812 1538 813 1579
rect 777 1504 813 1538
rect 777 1470 778 1504
rect 812 1470 813 1504
rect 777 1436 813 1470
rect 777 1402 778 1436
rect 812 1402 813 1436
rect 777 1368 813 1402
rect 777 1334 778 1368
rect 812 1334 813 1368
rect 777 1315 813 1334
rect 249 1252 250 1292
rect 284 1252 285 1292
rect 249 1219 285 1252
rect 249 1184 250 1219
rect 284 1184 285 1219
rect 249 1150 285 1184
rect 249 1116 250 1150
rect 284 1116 285 1150
rect 777 1266 778 1315
rect 812 1266 813 1315
rect 777 1232 813 1266
rect 777 1198 778 1232
rect 812 1198 813 1232
rect 777 1176 813 1198
rect 249 1082 285 1116
rect 249 1048 250 1082
rect 284 1048 285 1082
rect 249 1014 285 1048
rect 249 980 250 1014
rect 284 980 285 1014
rect 249 946 285 980
rect 249 912 250 946
rect 284 912 285 946
rect 249 878 285 912
rect 249 844 250 878
rect 284 844 285 878
rect 249 810 285 844
rect 249 766 250 810
rect 284 766 285 810
rect 249 742 285 766
rect 249 688 250 742
rect 284 688 285 742
rect 249 674 285 688
rect 249 610 250 674
rect 284 610 285 674
rect 249 606 285 610
rect 249 572 250 606
rect 284 572 285 606
rect 249 565 285 572
rect 249 504 250 565
rect 284 504 285 565
rect 249 486 285 504
rect 349 1133 383 1145
rect 349 1061 383 1095
rect 349 983 383 1022
rect 349 910 383 949
rect 349 871 383 876
rect 349 799 383 803
rect 349 764 383 765
rect 349 727 383 730
rect 349 691 383 693
rect 349 655 383 657
rect 349 619 383 621
rect 349 583 383 585
rect 349 547 383 549
rect 349 497 383 513
rect 777 1130 778 1176
rect 812 1130 813 1176
rect 777 1096 813 1130
rect 777 1062 778 1096
rect 812 1062 813 1096
rect 777 1028 813 1062
rect 777 994 778 1028
rect 812 994 813 1028
rect 777 960 813 994
rect 777 926 778 960
rect 812 926 813 960
rect 777 892 813 926
rect 777 858 778 892
rect 812 876 813 892
rect 966 1904 967 1966
rect 1001 1904 1002 1966
rect 966 1898 1002 1904
rect 966 1864 967 1898
rect 1001 1864 1002 1898
rect 966 1859 1002 1864
rect 1479 2039 1480 2097
rect 1514 2039 1515 2097
rect 1479 2023 1515 2039
rect 1479 1971 1480 2023
rect 1514 1971 1515 2023
rect 1479 1949 1515 1971
rect 1479 1903 1480 1949
rect 1514 1903 1515 1949
rect 1479 1875 1515 1903
rect 966 1796 967 1859
rect 1001 1796 1002 1859
rect 966 1780 1002 1796
rect 966 1728 967 1780
rect 1001 1728 1002 1780
rect 966 1701 1002 1728
rect 966 1660 967 1701
rect 1001 1660 1002 1701
rect 966 1626 1002 1660
rect 966 1588 967 1626
rect 1001 1588 1002 1626
rect 966 1558 1002 1588
rect 1052 1851 1086 1863
rect 1479 1835 1480 1875
rect 1514 1835 1515 1875
rect 1138 1822 1162 1828
rect 1052 1779 1086 1813
rect 1196 1794 1234 1828
rect 1268 1794 1306 1828
rect 1479 1801 1515 1835
rect 1052 1707 1086 1739
rect 1052 1635 1086 1665
rect 1479 1767 1480 1801
rect 1514 1767 1515 1801
rect 1479 1733 1515 1767
rect 1479 1693 1480 1733
rect 1514 1693 1515 1733
rect 1479 1665 1515 1693
rect 1196 1616 1234 1650
rect 1268 1616 1306 1650
rect 1479 1619 1480 1665
rect 1514 1619 1515 1665
rect 1052 1575 1086 1591
rect 1479 1597 1515 1619
rect 966 1510 967 1558
rect 1001 1510 1002 1558
rect 966 1490 1002 1510
rect 966 1456 967 1490
rect 1001 1456 1002 1490
rect 966 1422 1002 1456
rect 966 1366 967 1422
rect 1001 1366 1002 1422
rect 1479 1545 1480 1597
rect 1514 1545 1515 1597
rect 1479 1529 1515 1545
rect 1479 1471 1480 1529
rect 1514 1471 1515 1529
rect 1479 1461 1515 1471
rect 1479 1397 1480 1461
rect 1514 1397 1515 1461
rect 1479 1393 1515 1397
rect 966 1354 1002 1366
rect 966 1287 967 1354
rect 1001 1287 1002 1354
rect 966 1286 1002 1287
rect 966 1252 967 1286
rect 1001 1252 1002 1286
rect 966 1218 1002 1252
rect 966 1184 967 1218
rect 1001 1184 1002 1218
rect 966 1150 1002 1184
rect 966 1116 967 1150
rect 1001 1116 1002 1150
rect 966 1106 1002 1116
rect 966 1048 967 1106
rect 1001 1048 1002 1106
rect 966 1030 1002 1048
rect 966 980 967 1030
rect 1001 980 1002 1030
rect 966 946 1002 980
rect 966 912 967 946
rect 1001 912 1002 946
rect 966 878 1002 912
rect 777 842 789 858
rect 823 842 861 876
rect 777 824 813 842
rect 777 790 778 824
rect 812 790 813 824
rect 777 756 813 790
rect 777 722 778 756
rect 812 722 813 756
rect 777 688 813 722
rect 777 654 778 688
rect 812 654 813 688
rect 777 620 813 654
rect 777 586 778 620
rect 812 586 813 620
rect 777 582 813 586
rect 777 518 778 582
rect 812 518 813 582
rect 777 499 813 518
rect 249 436 250 486
rect 284 436 285 486
rect 249 407 285 436
rect 249 368 250 407
rect 284 370 285 407
rect 777 450 778 499
rect 812 450 813 499
rect 777 370 813 450
rect 284 369 813 370
rect 284 368 337 369
rect 249 335 337 368
rect 399 335 405 369
rect 439 335 440 369
rect 507 335 515 369
rect 575 335 590 369
rect 643 335 665 369
rect 711 335 740 369
rect 779 335 813 369
rect 249 334 813 335
rect 966 836 967 878
rect 1001 836 1002 878
rect 966 810 1002 836
rect 966 776 967 810
rect 1001 776 1002 810
rect 966 742 1002 776
rect 966 694 967 742
rect 1001 694 1002 742
rect 966 674 1002 694
rect 966 640 967 674
rect 1001 640 1002 674
rect 966 606 1002 640
rect 966 572 967 606
rect 1001 572 1002 606
rect 966 538 1002 572
rect 966 504 967 538
rect 1001 504 1002 538
rect 966 484 1002 504
rect 1052 1373 1086 1385
rect 1052 1301 1086 1335
rect 1052 1231 1086 1266
rect 1052 1162 1086 1197
rect 1052 1093 1086 1128
rect 1052 1024 1086 1059
rect 1052 955 1086 990
rect 1479 1359 1480 1393
rect 1514 1359 1515 1393
rect 1479 1357 1515 1359
rect 1479 1291 1480 1357
rect 1514 1291 1515 1357
rect 1479 1284 1515 1291
rect 1479 1223 1480 1284
rect 1514 1223 1515 1284
rect 1479 1211 1515 1223
rect 1479 1155 1480 1211
rect 1514 1155 1515 1211
rect 1479 1138 1515 1155
rect 1479 1087 1480 1138
rect 1514 1087 1515 1138
rect 1479 1065 1515 1087
rect 1479 1019 1480 1065
rect 1514 1019 1515 1065
rect 1479 992 1515 1019
rect 1243 924 1319 958
rect 1479 951 1480 992
rect 1514 951 1515 992
rect 1052 887 1086 921
rect 1052 819 1086 853
rect 1052 751 1086 785
rect 1052 683 1086 717
rect 1052 642 1086 649
rect 1052 570 1086 581
rect 1052 497 1086 513
rect 1479 919 1515 951
rect 1479 883 1480 919
rect 1514 883 1515 919
rect 1479 849 1515 883
rect 1479 812 1480 849
rect 1514 812 1515 849
rect 1479 781 1515 812
rect 1479 739 1480 781
rect 1514 739 1515 781
rect 1479 713 1515 739
rect 1479 666 1480 713
rect 1514 666 1515 713
rect 1479 645 1515 666
rect 1479 593 1480 645
rect 1514 593 1515 645
rect 1479 577 1515 593
rect 1479 520 1480 577
rect 1514 520 1515 577
rect 1479 509 1515 520
rect 966 436 967 484
rect 1001 436 1002 484
rect 966 407 1002 436
rect 966 368 967 407
rect 1001 370 1002 407
rect 1479 447 1480 509
rect 1514 447 1515 509
rect 1479 370 1515 447
rect 1001 369 1515 370
rect 1001 368 1039 369
rect 966 335 1039 368
rect 1073 335 1077 369
rect 1141 335 1150 369
rect 1209 335 1223 369
rect 1277 335 1296 369
rect 1345 335 1369 369
rect 1413 335 1442 369
rect 1481 335 1515 369
rect 966 334 1515 335
rect 1668 5163 3114 5164
rect 1668 5129 1702 5163
rect 1736 5129 1770 5163
rect 1819 5129 1838 5163
rect 1894 5129 1906 5163
rect 1969 5129 1974 5163
rect 2008 5129 2010 5163
rect 2076 5129 2085 5163
rect 2144 5129 2160 5163
rect 2212 5129 2235 5163
rect 2280 5129 2310 5163
rect 2348 5129 2382 5163
rect 2419 5129 2450 5163
rect 2494 5129 2518 5163
rect 2570 5129 2586 5163
rect 2646 5129 2654 5163
rect 2756 5129 2764 5163
rect 2824 5129 2840 5163
rect 2892 5129 2916 5163
rect 2960 5129 2992 5163
rect 3028 5129 3068 5163
rect 3102 5130 3114 5163
rect 1668 5128 3079 5129
rect 1668 5125 1704 5128
rect 1668 5060 1669 5125
rect 1703 5060 1704 5125
rect 1668 5051 1704 5060
rect 1668 4992 1669 5051
rect 1703 4992 1704 5051
rect 3078 5096 3079 5128
rect 3113 5096 3114 5130
rect 3078 5091 3114 5096
rect 3078 5028 3079 5091
rect 3113 5028 3114 5091
rect 1668 4977 1704 4992
rect 1668 4924 1669 4977
rect 1703 4924 1704 4977
rect 1668 4903 1704 4924
rect 1668 4856 1669 4903
rect 1703 4856 1704 4903
rect 1668 4829 1704 4856
rect 1668 4788 1669 4829
rect 1703 4788 1704 4829
rect 1668 4755 1704 4788
rect 1668 4720 1669 4755
rect 1703 4720 1704 4755
rect 1668 4686 1704 4720
rect 1668 4647 1669 4686
rect 1703 4647 1704 4686
rect 1668 4618 1704 4647
rect 1668 4573 1669 4618
rect 1703 4573 1704 4618
rect 1668 4550 1704 4573
rect 1668 4499 1669 4550
rect 1703 4499 1704 4550
rect 1668 4482 1704 4499
rect 1668 4425 1669 4482
rect 1703 4425 1704 4482
rect 1668 4414 1704 4425
rect 1668 4351 1669 4414
rect 1703 4351 1704 4414
rect 1668 4346 1704 4351
rect 1668 4312 1669 4346
rect 1703 4312 1704 4346
rect 1668 4311 1704 4312
rect 1668 4244 1669 4311
rect 1703 4244 1704 4311
rect 1668 4237 1704 4244
rect 1668 4176 1669 4237
rect 1703 4176 1704 4237
rect 1668 4163 1704 4176
rect 1668 4108 1669 4163
rect 1703 4108 1704 4163
rect 1668 4089 1704 4108
rect 1668 4040 1669 4089
rect 1703 4040 1704 4089
rect 1668 4015 1704 4040
rect 1668 3972 1669 4015
rect 1703 3972 1704 4015
rect 1668 3941 1704 3972
rect 1668 3904 1669 3941
rect 1703 3904 1704 3941
rect 1668 3870 1704 3904
rect 1668 3833 1669 3870
rect 1703 3833 1704 3870
rect 1668 3802 1704 3833
rect 1668 3759 1669 3802
rect 1703 3759 1704 3802
rect 1668 3734 1704 3759
rect 1668 3685 1669 3734
rect 1703 3685 1704 3734
rect 1668 3666 1704 3685
rect 1668 3612 1669 3666
rect 1703 3612 1704 3666
rect 1668 3598 1704 3612
rect 1668 3539 1669 3598
rect 1703 3539 1704 3598
rect 1668 3530 1704 3539
rect 1668 3466 1669 3530
rect 1703 3466 1704 3530
rect 1668 3462 1704 3466
rect 1668 3428 1669 3462
rect 1703 3428 1704 3462
rect 1668 3427 1704 3428
rect 1668 3360 1669 3427
rect 1703 3360 1704 3427
rect 1668 3354 1704 3360
rect 1668 3292 1669 3354
rect 1703 3292 1704 3354
rect 1668 3281 1704 3292
rect 1668 3224 1669 3281
rect 1703 3224 1704 3281
rect 1668 3208 1704 3224
rect 1668 3156 1669 3208
rect 1703 3156 1704 3208
rect 1668 3135 1704 3156
rect 1668 3088 1669 3135
rect 1703 3088 1704 3135
rect 1668 3062 1704 3088
rect 1668 3020 1669 3062
rect 1703 3020 1704 3062
rect 1668 2989 1704 3020
rect 1668 2952 1669 2989
rect 1703 2952 1704 2989
rect 1668 2918 1704 2952
rect 1668 2884 1669 2918
rect 1703 2884 1704 2918
rect 1668 2850 1704 2884
rect 1668 2816 1669 2850
rect 1703 2816 1704 2850
rect 1668 2782 1704 2816
rect 1668 2748 1669 2782
rect 1703 2748 1704 2782
rect 1668 2714 1704 2748
rect 1668 2680 1669 2714
rect 1703 2680 1704 2714
rect 1668 2646 1704 2680
rect 1668 2612 1669 2646
rect 1703 2612 1704 2646
rect 1668 2578 1704 2612
rect 1668 2544 1669 2578
rect 1703 2544 1704 2578
rect 1668 2524 1704 2544
rect 1668 2476 1669 2524
rect 1703 2476 1704 2524
rect 1668 2451 1704 2476
rect 1668 2408 1669 2451
rect 1703 2408 1704 2451
rect 1668 2378 1704 2408
rect 1668 2340 1669 2378
rect 1703 2340 1704 2378
rect 1668 2306 1704 2340
rect 1668 2271 1669 2306
rect 1703 2271 1704 2306
rect 1668 2238 1704 2271
rect 1668 2198 1669 2238
rect 1703 2198 1704 2238
rect 1668 2170 1704 2198
rect 1668 2125 1669 2170
rect 1703 2125 1704 2170
rect 1668 2102 1704 2125
rect 1668 2052 1669 2102
rect 1703 2052 1704 2102
rect 1668 2034 1704 2052
rect 1668 1979 1669 2034
rect 1703 1979 1704 2034
rect 1668 1966 1704 1979
rect 1668 1906 1669 1966
rect 1703 1906 1704 1966
rect 1668 1898 1704 1906
rect 1668 1833 1669 1898
rect 1703 1833 1704 1898
rect 1668 1830 1704 1833
rect 1668 1796 1669 1830
rect 1703 1796 1704 1830
rect 1668 1794 1704 1796
rect 1668 1728 1669 1794
rect 1703 1728 1704 1794
rect 1668 1721 1704 1728
rect 1668 1660 1669 1721
rect 1703 1660 1704 1721
rect 1668 1648 1704 1660
rect 1668 1592 1669 1648
rect 1703 1592 1704 1648
rect 1668 1575 1704 1592
rect 1668 1524 1669 1575
rect 1703 1524 1704 1575
rect 1668 1502 1704 1524
rect 1668 1456 1669 1502
rect 1703 1456 1704 1502
rect 1668 1429 1704 1456
rect 1668 1388 1669 1429
rect 1703 1388 1704 1429
rect 1668 1356 1704 1388
rect 1668 1320 1669 1356
rect 1703 1320 1704 1356
rect 1668 1286 1704 1320
rect 1668 1249 1669 1286
rect 1703 1249 1704 1286
rect 1668 1218 1704 1249
rect 1668 1176 1669 1218
rect 1703 1176 1704 1218
rect 1668 1150 1704 1176
rect 1668 1103 1669 1150
rect 1703 1103 1704 1150
rect 1668 1082 1704 1103
rect 1668 1030 1669 1082
rect 1703 1030 1704 1082
rect 1668 1014 1704 1030
rect 1668 957 1669 1014
rect 1703 957 1704 1014
rect 1668 946 1704 957
rect 1668 884 1669 946
rect 1703 884 1704 946
rect 1668 878 1704 884
rect 1668 811 1669 878
rect 1703 811 1704 878
rect 1668 810 1704 811
rect 1668 776 1669 810
rect 1703 776 1704 810
rect 1668 772 1704 776
rect 1668 708 1669 772
rect 1703 708 1704 772
rect 1668 699 1704 708
rect 1668 640 1669 699
rect 1703 640 1704 699
rect 1668 626 1704 640
rect 1668 572 1669 626
rect 1703 572 1704 626
rect 1668 553 1704 572
rect 1668 504 1669 553
rect 1703 504 1704 553
rect 1668 480 1704 504
rect 1752 4985 1788 5017
rect 3078 5015 3114 5028
rect 1752 4951 1754 4985
rect 1752 4902 1788 4951
rect 1752 4868 1754 4902
rect 1752 4819 1788 4868
rect 1752 4785 1754 4819
rect 1752 4735 1788 4785
rect 1752 4701 1754 4735
rect 1752 4651 1788 4701
rect 1752 4617 1754 4651
rect 1752 4529 1788 4617
rect 2484 4985 2518 5001
rect 2484 4902 2518 4951
rect 2484 4819 2518 4868
rect 2484 4735 2518 4785
rect 2484 4651 2518 4701
rect 2484 4601 2518 4617
rect 3078 4960 3079 5015
rect 3113 4960 3114 5015
rect 3078 4939 3114 4960
rect 3078 4892 3079 4939
rect 3113 4892 3114 4939
rect 3078 4863 3114 4892
rect 3078 4824 3079 4863
rect 3113 4824 3114 4863
rect 3078 4790 3114 4824
rect 3078 4753 3079 4790
rect 3113 4753 3114 4790
rect 3078 4722 3114 4753
rect 3078 4677 3079 4722
rect 3113 4677 3114 4722
rect 3078 4654 3114 4677
rect 3078 4601 3079 4654
rect 3113 4601 3114 4654
rect 3078 4586 3114 4601
rect 3078 4560 3079 4586
rect 1752 4495 1754 4529
rect 2870 4526 3079 4560
rect 1752 4446 1788 4495
rect 1752 4412 1754 4446
rect 2914 4525 3079 4526
rect 3113 4525 3114 4586
rect 2914 4518 3114 4525
rect 2914 4484 3079 4518
rect 3113 4484 3114 4518
rect 2914 4482 3114 4484
rect 2948 4448 2982 4482
rect 3016 4448 3079 4482
rect 2914 4432 3079 4448
rect 1752 4363 1788 4412
rect 1752 4329 1754 4363
rect 3078 4416 3079 4432
rect 3113 4416 3114 4482
rect 3078 4405 3114 4416
rect 1752 4279 1788 4329
rect 1752 4245 1754 4279
rect 1752 4195 1788 4245
rect 1752 4161 1754 4195
rect 1752 4073 1788 4161
rect 1752 4039 1754 4073
rect 1752 3990 1788 4039
rect 1752 3956 1754 3990
rect 1752 3907 1788 3956
rect 1752 3873 1754 3907
rect 1752 3823 1788 3873
rect 1752 3789 1754 3823
rect 1752 3739 1788 3789
rect 1752 3705 1754 3739
rect 1752 3617 1788 3705
rect 1752 3583 1754 3617
rect 1752 3534 1788 3583
rect 1752 3500 1754 3534
rect 1752 3451 1788 3500
rect 1752 3417 1754 3451
rect 1752 3367 1788 3417
rect 1752 3333 1754 3367
rect 1752 3283 1788 3333
rect 1752 3249 1754 3283
rect 1752 3161 1788 3249
rect 2484 4343 2518 4359
rect 2484 4272 2518 4309
rect 2484 4201 2518 4238
rect 2484 4130 2518 4167
rect 2484 4059 2518 4096
rect 2484 3988 2518 4025
rect 2484 3917 2518 3954
rect 3078 4348 3079 4405
rect 3113 4348 3114 4405
rect 3078 4328 3114 4348
rect 3078 4280 3079 4328
rect 3113 4280 3114 4328
rect 3078 4246 3114 4280
rect 3078 4212 3079 4246
rect 3113 4212 3114 4246
rect 3078 4178 3114 4212
rect 3078 4134 3079 4178
rect 3113 4134 3114 4178
rect 3078 4110 3114 4134
rect 3078 4058 3079 4110
rect 3113 4058 3114 4110
rect 3078 4042 3114 4058
rect 3078 3983 3079 4042
rect 3113 3983 3114 4042
rect 3078 3974 3114 3983
rect 2654 3902 2692 3936
rect 2726 3902 2764 3936
rect 3078 3908 3079 3974
rect 3113 3908 3114 3974
rect 3078 3906 3114 3908
rect 2484 3845 2518 3883
rect 2484 3773 2518 3811
rect 2484 3701 2518 3739
rect 2484 3629 2518 3667
rect 3078 3872 3079 3906
rect 3113 3872 3114 3906
rect 3078 3838 3114 3872
rect 3078 3804 3079 3838
rect 3113 3804 3114 3838
rect 3078 3770 3114 3804
rect 3078 3709 3079 3770
rect 3113 3709 3114 3770
rect 3078 3702 3114 3709
rect 3078 3668 3079 3702
rect 3113 3668 3114 3702
rect 3078 3645 3114 3668
rect 2484 3557 2518 3595
rect 2600 3578 2620 3590
rect 2654 3578 2692 3612
rect 2726 3578 2764 3612
rect 2798 3578 2836 3612
rect 3078 3600 3079 3645
rect 3113 3600 3114 3645
rect 2484 3485 2518 3523
rect 2484 3413 2518 3451
rect 2484 3341 2518 3379
rect 3078 3566 3114 3600
rect 3078 3514 3079 3566
rect 3113 3514 3114 3566
rect 3078 3498 3114 3514
rect 3078 3464 3079 3498
rect 3113 3464 3114 3498
rect 3078 3430 3114 3464
rect 3078 3396 3079 3430
rect 3113 3396 3114 3430
rect 3078 3388 3114 3396
rect 3078 3328 3079 3388
rect 3113 3328 3114 3388
rect 2484 3269 2518 3307
rect 2654 3278 2692 3312
rect 2726 3278 2764 3312
rect 3078 3302 3114 3328
rect 2484 3219 2518 3235
rect 3078 3260 3079 3302
rect 3113 3260 3114 3302
rect 3078 3226 3114 3260
rect 1752 3127 1754 3161
rect 1752 3078 1788 3127
rect 3078 3182 3079 3226
rect 3113 3182 3114 3226
rect 3078 3158 3114 3182
rect 3078 3097 3079 3158
rect 3113 3097 3114 3158
rect 3078 3094 3114 3097
rect 1752 3044 1754 3078
rect 1752 2995 1788 3044
rect 2914 3090 3114 3094
rect 2914 3078 3079 3090
rect 2948 3044 2982 3078
rect 3016 3056 3079 3078
rect 3113 3056 3114 3090
rect 3016 3046 3114 3056
rect 3016 3044 3079 3046
rect 2914 3028 3079 3044
rect 1752 2961 1754 2995
rect 1752 2911 1788 2961
rect 3078 2988 3079 3028
rect 3113 2988 3114 3046
rect 3078 2961 3114 2988
rect 1752 2877 1754 2911
rect 1752 2838 1788 2877
rect 1786 2827 1788 2838
rect 1752 2793 1754 2804
rect 1752 2766 1788 2793
rect 1786 2732 1788 2766
rect 1752 2705 1788 2732
rect 1752 2694 1754 2705
rect 1786 2660 1788 2671
rect 2484 2939 2518 2955
rect 2484 2838 2518 2905
rect 2484 2766 2518 2779
rect 2484 2694 2518 2732
rect 3078 2920 3079 2961
rect 3113 2920 3114 2961
rect 3078 2886 3114 2920
rect 3078 2852 3079 2886
rect 3113 2852 3114 2886
rect 3078 2818 3114 2852
rect 3078 2784 3079 2818
rect 3113 2784 3114 2818
rect 3078 2750 3114 2784
rect 3078 2716 3079 2750
rect 3113 2716 3114 2750
rect 3078 2682 3114 2716
rect 1752 2622 1788 2660
rect 3078 2648 3079 2682
rect 3113 2648 3114 2682
rect 1752 2588 1754 2622
rect 1752 2539 1788 2588
rect 1752 2505 1754 2539
rect 2914 2616 3044 2632
rect 2948 2582 2982 2616
rect 3016 2582 3044 2616
rect 2914 2545 3044 2582
rect 2914 2511 2922 2545
rect 2956 2511 2994 2545
rect 3028 2511 3044 2545
rect 3078 2614 3114 2648
rect 3078 2560 3079 2614
rect 3113 2560 3114 2614
rect 3078 2546 3114 2560
rect 1752 2455 1788 2505
rect 1752 2421 1754 2455
rect 2600 2470 2870 2498
rect 3078 2485 3079 2546
rect 3113 2485 3114 2546
rect 3078 2478 3114 2485
rect 3078 2470 3079 2478
rect 2600 2436 2914 2470
rect 2948 2436 2982 2470
rect 3016 2436 3079 2470
rect 1752 2371 1788 2421
rect 2914 2404 3079 2436
rect 1752 2337 1754 2371
rect 1752 2249 1788 2337
rect 3078 2376 3079 2404
rect 3113 2376 3114 2478
rect 3078 2369 3114 2376
rect 3078 2308 3079 2369
rect 3113 2308 3114 2369
rect 3078 2294 3114 2308
rect 1752 2215 1754 2249
rect 1752 2166 1788 2215
rect 1752 2132 1754 2166
rect 1752 2083 1788 2132
rect 1752 2049 1754 2083
rect 1752 1999 1788 2049
rect 1752 1965 1754 1999
rect 1752 1915 1788 1965
rect 1752 1881 1754 1915
rect 1752 1793 1788 1881
rect 1752 1759 1754 1793
rect 1752 1710 1788 1759
rect 1752 1676 1754 1710
rect 1752 1627 1788 1676
rect 1752 1593 1754 1627
rect 1752 1543 1788 1593
rect 1752 1509 1754 1543
rect 1752 1459 1788 1509
rect 1752 1425 1754 1459
rect 1752 1337 1788 1425
rect 1752 1303 1754 1337
rect 1752 1254 1788 1303
rect 1752 1220 1754 1254
rect 1752 1171 1788 1220
rect 1752 1137 1754 1171
rect 2484 2249 2518 2265
rect 2484 2179 2518 2215
rect 2484 2109 2518 2145
rect 2484 2039 2518 2075
rect 2484 1969 2518 2005
rect 2484 1899 2518 1935
rect 2484 1828 2518 1865
rect 2484 1757 2518 1794
rect 2484 1686 2518 1723
rect 2484 1615 2518 1652
rect 2484 1544 2518 1581
rect 2484 1473 2518 1510
rect 2484 1402 2518 1439
rect 2484 1331 2518 1368
rect 2484 1260 2518 1297
rect 3078 2240 3079 2294
rect 3113 2240 3114 2294
rect 3078 2219 3114 2240
rect 3078 2172 3079 2219
rect 3113 2172 3114 2219
rect 3078 2144 3114 2172
rect 3078 2104 3079 2144
rect 3113 2104 3114 2144
rect 3078 2070 3114 2104
rect 3078 2036 3079 2070
rect 3113 2036 3114 2070
rect 3078 2002 3114 2036
rect 3078 1950 3079 2002
rect 3113 1950 3114 2002
rect 3078 1934 3114 1950
rect 3078 1900 3079 1934
rect 3113 1900 3114 1934
rect 3078 1886 3114 1900
rect 3078 1832 3079 1886
rect 3113 1832 3114 1886
rect 3078 1798 3114 1832
rect 3078 1755 3079 1798
rect 3113 1755 3114 1798
rect 3078 1730 3114 1755
rect 3078 1696 3079 1730
rect 3113 1696 3114 1730
rect 3078 1662 3114 1696
rect 3078 1628 3079 1662
rect 3113 1628 3114 1662
rect 3078 1594 3114 1628
rect 3078 1556 3079 1594
rect 3113 1556 3114 1594
rect 3078 1526 3114 1556
rect 3078 1480 3079 1526
rect 3113 1480 3114 1526
rect 3078 1458 3114 1480
rect 3078 1405 3079 1458
rect 3113 1405 3114 1458
rect 3078 1390 3114 1405
rect 3078 1330 3079 1390
rect 3113 1330 3114 1390
rect 3078 1322 3114 1330
rect 3078 1288 3079 1322
rect 3113 1288 3114 1322
rect 2654 1250 2692 1284
rect 2726 1250 2764 1284
rect 3078 1254 3114 1288
rect 2484 1189 2518 1226
rect 2484 1139 2518 1155
rect 3078 1220 3079 1254
rect 3113 1220 3114 1254
rect 3078 1204 3114 1220
rect 3078 1152 3079 1204
rect 3113 1152 3114 1204
rect 1752 1087 1788 1137
rect 1752 1053 1754 1087
rect 3078 1130 3114 1152
rect 3078 1084 3079 1130
rect 3113 1084 3114 1130
rect 3078 1066 3114 1084
rect 1752 1003 1788 1053
rect 1752 969 1754 1003
rect 2914 1057 3114 1066
rect 2914 1050 3079 1057
rect 2948 1016 2982 1050
rect 3016 1016 3079 1050
rect 3113 1016 3114 1057
rect 2914 984 3114 1016
rect 2914 972 3079 984
rect 1752 881 1788 969
rect 2870 948 3079 972
rect 3113 948 3114 984
rect 2870 938 3114 948
rect 3078 914 3114 938
rect 1752 847 1754 881
rect 1752 798 1788 847
rect 1752 764 1754 798
rect 1752 715 1788 764
rect 1752 681 1754 715
rect 1752 631 1788 681
rect 1752 597 1754 631
rect 1752 547 1788 597
rect 1752 513 1754 547
rect 1752 481 1788 513
rect 2484 881 2518 897
rect 2484 798 2518 847
rect 2484 715 2518 764
rect 2484 631 2518 681
rect 2484 547 2518 597
rect 2484 497 2518 513
rect 3078 880 3079 914
rect 3113 880 3114 914
rect 3078 846 3114 880
rect 3078 812 3079 846
rect 3113 812 3114 846
rect 3078 778 3114 812
rect 3078 744 3079 778
rect 3113 744 3114 778
rect 3078 710 3114 744
rect 3078 661 3079 710
rect 3113 661 3114 710
rect 3078 642 3114 661
rect 3078 589 3079 642
rect 3113 589 3114 642
rect 3078 574 3114 589
rect 3078 517 3079 574
rect 3113 517 3114 574
rect 3078 506 3114 517
rect 1668 436 1669 480
rect 1703 436 1704 480
rect 1668 407 1704 436
rect 1668 368 1669 407
rect 1703 370 1704 407
rect 3078 445 3079 506
rect 3113 445 3114 506
rect 3078 370 3114 445
rect 1703 369 3114 370
rect 1703 368 1754 369
rect 1668 335 1754 368
rect 1817 335 1822 369
rect 1856 335 1857 369
rect 1924 335 1931 369
rect 1992 335 2005 369
rect 2060 335 2079 369
rect 2128 335 2153 369
rect 2196 335 2227 369
rect 2264 335 2298 369
rect 2335 335 2366 369
rect 2409 335 2434 369
rect 2483 335 2502 369
rect 2557 335 2570 369
rect 2631 335 2638 369
rect 2705 335 2706 369
rect 2740 335 2745 369
rect 2808 335 2819 369
rect 2876 335 2893 369
rect 2944 335 2967 369
rect 3012 335 3041 369
rect 3080 335 3114 369
rect 3268 5153 4200 5182
rect 3268 5130 3713 5153
rect 3747 5148 3792 5153
rect 3826 5148 3870 5153
rect 3904 5148 3948 5153
rect 3982 5148 4026 5153
rect 4060 5148 4104 5153
rect 3268 5129 3490 5130
rect 3302 5095 3336 5129
rect 3370 5095 3404 5129
rect 3438 5096 3490 5129
rect 3524 5096 3558 5130
rect 3592 5096 3626 5130
rect 3660 5119 3713 5130
rect 3764 5119 3792 5148
rect 3660 5096 3730 5119
rect 3764 5114 3798 5119
rect 3832 5114 3866 5148
rect 3904 5119 3934 5148
rect 3982 5119 4002 5148
rect 4060 5119 4070 5148
rect 3900 5114 3934 5119
rect 3968 5114 4002 5119
rect 4036 5114 4070 5119
rect 4138 5148 4200 5153
rect 4645 5473 4681 5507
rect 4645 5439 4646 5473
rect 4680 5439 4681 5473
rect 4645 5405 4681 5439
rect 4645 5371 4646 5405
rect 4680 5371 4681 5405
rect 4645 5337 4681 5371
rect 4645 5303 4646 5337
rect 4680 5303 4681 5337
rect 4645 5269 4681 5303
rect 4645 5235 4646 5269
rect 4680 5235 4681 5269
rect 4645 5201 4681 5235
rect 4645 5167 4646 5201
rect 4680 5167 4681 5201
rect 4104 5114 4138 5119
rect 4172 5114 4206 5148
rect 4240 5114 4300 5148
rect 3438 5095 3730 5096
rect 3268 5061 3730 5095
rect 3268 5060 3490 5061
rect 3302 5026 3336 5060
rect 3370 5026 3404 5060
rect 3438 5027 3490 5060
rect 3524 5027 3558 5061
rect 3592 5027 3626 5061
rect 3660 5042 3730 5061
rect 3660 5027 3696 5042
rect 3438 5026 3696 5027
rect 3268 5008 3696 5026
rect 3268 4992 3730 5008
rect 4266 5058 4300 5114
rect 3268 4991 3490 4992
rect 3302 4957 3336 4991
rect 3370 4957 3404 4991
rect 3438 4957 3490 4991
rect 3268 4922 3490 4957
rect 3302 4888 3336 4922
rect 3370 4888 3404 4922
rect 3438 4888 3490 4922
rect 3268 4853 3490 4888
rect 3302 4819 3336 4853
rect 3370 4819 3404 4853
rect 3438 4819 3490 4853
rect 3268 4784 3490 4819
rect 3302 4750 3336 4784
rect 3370 4750 3404 4784
rect 3438 4750 3490 4784
rect 3268 4715 3490 4750
rect 3302 4681 3336 4715
rect 3370 4681 3404 4715
rect 3438 4681 3490 4715
rect 3268 4646 3490 4681
rect 3302 4612 3336 4646
rect 3370 4612 3404 4646
rect 3438 4612 3490 4646
rect 3268 4577 3490 4612
rect 3302 4543 3336 4577
rect 3370 4543 3404 4577
rect 3438 4543 3490 4577
rect 3268 4508 3490 4543
rect 3302 4474 3336 4508
rect 3370 4474 3404 4508
rect 3438 4474 3490 4508
rect 3268 4439 3490 4474
rect 3302 4405 3336 4439
rect 3370 4405 3404 4439
rect 3438 4405 3490 4439
rect 3268 4370 3490 4405
rect 3302 4336 3336 4370
rect 3370 4336 3404 4370
rect 3438 4336 3490 4370
rect 3268 4301 3490 4336
rect 3302 4267 3336 4301
rect 3370 4267 3404 4301
rect 3438 4267 3490 4301
rect 3268 4232 3490 4267
rect 3302 4198 3336 4232
rect 3370 4198 3404 4232
rect 3438 4198 3490 4232
rect 3268 4163 3490 4198
rect 3302 4129 3336 4163
rect 3370 4129 3404 4163
rect 3438 4129 3490 4163
rect 3268 4094 3490 4129
rect 3302 4060 3336 4094
rect 3370 4060 3404 4094
rect 3438 4060 3490 4094
rect 3268 4025 3490 4060
rect 3302 3991 3336 4025
rect 3370 3991 3404 4025
rect 3438 3991 3490 4025
rect 3268 3956 3490 3991
rect 3302 3922 3336 3956
rect 3370 3922 3404 3956
rect 3438 3922 3490 3956
rect 3268 3887 3490 3922
rect 3302 3853 3336 3887
rect 3370 3853 3404 3887
rect 3438 3853 3490 3887
rect 3268 3818 3490 3853
rect 3302 3784 3336 3818
rect 3370 3784 3404 3818
rect 3438 3784 3490 3818
rect 3268 3749 3490 3784
rect 3302 3715 3336 3749
rect 3370 3715 3404 3749
rect 3438 3715 3490 3749
rect 3268 3680 3490 3715
rect 3302 3646 3336 3680
rect 3370 3646 3404 3680
rect 3438 3646 3490 3680
rect 3268 3611 3490 3646
rect 3302 3577 3336 3611
rect 3370 3577 3404 3611
rect 3438 3577 3490 3611
rect 3268 3542 3490 3577
rect 3302 3508 3336 3542
rect 3370 3508 3404 3542
rect 3438 3530 3490 3542
rect 3660 4974 3730 4992
rect 3660 4940 3696 4974
rect 3660 4906 3730 4940
rect 3660 4872 3696 4906
rect 3660 4838 3730 4872
rect 3660 4804 3696 4838
rect 3660 4770 3730 4804
rect 3852 4963 3944 4997
rect 4266 4980 4300 5014
rect 3852 4936 3886 4963
rect 3852 4842 3886 4902
rect 3852 4792 3886 4808
rect 4266 4912 4300 4920
rect 4266 4850 4300 4878
rect 3660 4736 3696 4770
rect 3660 4702 3730 4736
rect 3660 4668 3696 4702
rect 3660 4634 3730 4668
rect 3660 4600 3696 4634
rect 3660 4566 3730 4600
rect 3660 4532 3696 4566
rect 4266 4776 4300 4810
rect 4266 4708 4300 4742
rect 4266 4640 4300 4674
rect 4645 5133 4681 5167
rect 4645 5099 4646 5133
rect 4680 5099 4681 5133
rect 13646 6232 13682 6266
rect 13646 6198 13647 6232
rect 13681 6198 13682 6232
rect 13646 6164 13682 6198
rect 13646 6130 13647 6164
rect 13681 6130 13682 6164
rect 13646 6096 13682 6130
rect 13646 6062 13647 6096
rect 13681 6062 13682 6096
rect 13646 6028 13682 6062
rect 13646 5994 13647 6028
rect 13681 5994 13682 6028
rect 13646 5960 13682 5994
rect 13646 5926 13647 5960
rect 13681 5926 13682 5960
rect 13646 5892 13682 5926
rect 13646 5858 13647 5892
rect 13681 5858 13682 5892
rect 13646 5824 13682 5858
rect 13646 5790 13647 5824
rect 13681 5790 13682 5824
rect 13646 5756 13682 5790
rect 13646 5722 13647 5756
rect 13681 5722 13682 5756
rect 13646 5688 13682 5722
rect 13646 5654 13647 5688
rect 13681 5654 13682 5688
rect 13646 5620 13682 5654
rect 13646 5586 13647 5620
rect 13681 5586 13682 5620
rect 13646 5552 13682 5586
rect 13646 5518 13647 5552
rect 13681 5518 13682 5552
rect 13774 5540 13812 5574
rect 13846 5540 14063 5574
rect 13646 5484 13682 5518
rect 13646 5450 13647 5484
rect 13681 5450 13682 5484
rect 13774 5466 13812 5500
rect 13846 5466 13991 5500
rect 13646 5416 13682 5450
rect 13646 5382 13647 5416
rect 13681 5382 13682 5416
rect 13646 5348 13682 5382
rect 13646 5314 13647 5348
rect 13681 5314 13682 5348
rect 13646 5280 13682 5314
rect 13646 5246 13647 5280
rect 13681 5246 13682 5280
rect 13646 5212 13682 5246
rect 13646 5178 13647 5212
rect 13681 5178 13682 5212
rect 13957 5237 13991 5466
rect 14029 5305 14063 5540
rect 14029 5271 14355 5305
rect 14389 5271 14427 5305
rect 14547 5271 14585 5305
rect 14513 5237 14619 5271
rect 13957 5203 14619 5237
rect 4645 5065 4681 5099
rect 4645 5031 4646 5065
rect 4680 5031 4681 5065
rect 4645 4997 4681 5031
rect 4645 4963 4646 4997
rect 4680 4963 4681 4997
rect 4645 4929 4681 4963
rect 4645 4895 4646 4929
rect 4680 4895 4681 4929
rect 4645 4861 4681 4895
rect 4645 4827 4646 4861
rect 4680 4827 4681 4861
rect 4645 4793 4681 4827
rect 4645 4759 4646 4793
rect 4680 4759 4681 4793
rect 4645 4725 4681 4759
rect 4645 4691 4646 4725
rect 4680 4691 4681 4725
rect 4645 4657 4681 4691
rect 4645 4623 4646 4657
rect 4680 4623 4681 4657
rect 4645 4607 4681 4623
rect 4266 4572 4300 4606
rect 3660 4498 3730 4532
rect 4096 4501 4174 4535
rect 3660 4464 3696 4498
rect 3660 4430 3730 4464
rect 3660 4396 3696 4430
rect 3660 4362 3730 4396
rect 3660 4328 3696 4362
rect 3660 4294 3730 4328
rect 3660 4260 3696 4294
rect 3660 4226 3730 4260
rect 3660 4192 3696 4226
rect 3660 4158 3730 4192
rect 3660 4124 3696 4158
rect 3660 4090 3730 4124
rect 3660 4056 3696 4090
rect 3660 4022 3730 4056
rect 3660 3988 3696 4022
rect 3660 3954 3730 3988
rect 3660 3920 3696 3954
rect 3660 3886 3730 3920
rect 3660 3852 3696 3886
rect 3660 3818 3730 3852
rect 3660 3784 3696 3818
rect 3660 3750 3730 3784
rect 3660 3716 3696 3750
rect 3660 3682 3730 3716
rect 3660 3648 3696 3682
rect 3660 3614 3730 3648
rect 3660 3580 3696 3614
rect 4140 4474 4174 4501
rect 4140 4400 4174 4440
rect 4140 4332 4174 4366
rect 4140 4259 4174 4292
rect 4140 4186 4174 4218
rect 4140 4113 4174 4144
rect 4140 4040 4174 4070
rect 4140 3956 4174 3996
rect 4140 3882 4174 3922
rect 4140 3808 4174 3848
rect 4140 3734 4174 3774
rect 4140 3660 4174 3700
rect 4140 3610 4174 3626
rect 4266 4504 4300 4538
rect 4565 4595 4681 4607
rect 4565 4561 4574 4595
rect 4608 4561 4646 4595
rect 4565 4555 4646 4561
rect 4680 4555 4681 4595
rect 4565 4528 4681 4555
rect 4266 4436 4300 4470
rect 4266 4368 4300 4402
rect 4266 4330 4300 4334
rect 4266 4232 4300 4266
rect 4266 4164 4300 4188
rect 4266 4096 4300 4130
rect 4266 4028 4300 4062
rect 4266 3960 4300 3994
rect 4266 3892 4300 3926
rect 4266 3824 4300 3858
rect 4266 3756 4300 3790
rect 4266 3688 4300 3709
rect 4266 3645 4300 3654
rect 3660 3546 3730 3580
rect 3660 3530 3696 3546
rect 3438 3512 3696 3530
rect 3438 3508 3730 3512
rect 3268 3506 3730 3508
rect 3268 3473 3438 3506
rect 3302 3439 3336 3473
rect 3370 3439 3404 3473
rect 3268 3404 3438 3439
rect 3302 3370 3336 3404
rect 3370 3370 3404 3404
rect 3696 3478 3730 3506
rect 3696 3410 3730 3444
rect 3268 3335 3438 3370
rect 3302 3301 3336 3335
rect 3370 3301 3404 3335
rect 3268 3266 3438 3301
rect 3302 3232 3336 3266
rect 3370 3232 3404 3266
rect 3534 3360 3550 3394
rect 3584 3360 3600 3394
rect 3534 3347 3600 3360
rect 3534 3292 3550 3347
rect 3584 3292 3600 3347
rect 3534 3275 3600 3292
rect 3534 3241 3550 3275
rect 3584 3241 3600 3275
rect 3696 3342 3730 3376
rect 3696 3274 3730 3308
rect 3268 3197 3438 3232
rect 3302 3163 3336 3197
rect 3370 3163 3404 3197
rect 3268 3128 3438 3163
rect 3696 3206 3730 3240
rect 3696 3138 3730 3172
rect 3696 3070 3730 3104
rect 4266 3552 4300 3586
rect 4266 3484 4300 3514
rect 4266 3416 4300 3450
rect 4266 3348 4300 3382
rect 4266 3280 4300 3314
rect 4266 3212 4300 3239
rect 4266 3144 4300 3166
rect 3696 3002 3730 3036
rect 3696 2934 3730 2968
rect 3696 2866 3730 2900
rect 3696 2798 3730 2832
rect 3696 2730 3730 2764
rect 3696 2662 3730 2696
rect 3696 2594 3730 2628
rect 3696 2526 3730 2560
rect 3696 2458 3730 2492
rect 3696 2390 3730 2424
rect 3780 3085 3814 3101
rect 3780 3036 3814 3051
rect 3780 2943 3814 2980
rect 4266 3076 4300 3093
rect 4266 3008 4300 3020
rect 3928 2916 3966 2950
rect 4266 2940 4300 2947
rect 3780 2872 3814 2904
rect 4266 2872 4300 2874
rect 3780 2801 3814 2838
rect 3928 2824 3966 2858
rect 4000 2824 4059 2858
rect 4266 2835 4300 2838
rect 3780 2730 3814 2767
rect 3780 2659 3814 2696
rect 3780 2588 3814 2625
rect 4266 2763 4300 2770
rect 4266 2691 4300 2702
rect 4266 2619 4300 2634
rect 3780 2517 3814 2554
rect 3928 2548 3966 2582
rect 3780 2447 3814 2483
rect 3780 2397 3814 2413
rect 4266 2547 4300 2566
rect 4266 2475 4300 2498
rect 4266 2403 4300 2430
rect 3696 2322 3730 2356
rect 3534 2223 3550 2257
rect 3584 2223 3600 2257
rect 3534 2185 3600 2223
rect 3534 2121 3550 2185
rect 3584 2121 3600 2185
rect 3534 2087 3600 2121
rect 3534 2053 3550 2087
rect 3584 2053 3600 2087
rect 3696 2254 3730 2288
rect 3696 2186 3730 2220
rect 3696 2118 3730 2152
rect 4266 2331 4300 2362
rect 4266 2260 4300 2294
rect 4266 2192 4300 2225
rect 3696 2050 3730 2084
rect 3696 1982 3730 2016
rect 3696 1941 3730 1948
rect 3438 1917 3730 1941
rect 3852 2121 3886 2137
rect 3852 2027 3886 2087
rect 3852 1966 3886 1993
rect 4266 2124 4300 2158
rect 4266 2056 4300 2090
rect 4266 1988 4300 2022
rect 3852 1932 3944 1966
rect 3438 1883 3490 1917
rect 3524 1883 3558 1917
rect 3592 1883 3626 1917
rect 3660 1914 3730 1917
rect 3660 1883 3696 1914
rect 3438 1880 3696 1883
rect 3438 1848 3730 1880
rect 3438 1814 3490 1848
rect 3524 1814 3558 1848
rect 3592 1814 3626 1848
rect 3660 1846 3730 1848
rect 3660 1814 3696 1846
rect 3438 1812 3696 1814
rect 3438 1779 3730 1812
rect 3438 1745 3490 1779
rect 3524 1745 3558 1779
rect 3592 1745 3626 1779
rect 3660 1778 3730 1779
rect 3660 1745 3696 1778
rect 3438 1744 3696 1745
rect 3438 1710 3730 1744
rect 3438 1676 3490 1710
rect 3524 1676 3558 1710
rect 3592 1676 3626 1710
rect 3660 1676 3696 1710
rect 3438 1642 3730 1676
rect 3438 1641 3696 1642
rect 3438 1607 3490 1641
rect 3524 1607 3558 1641
rect 3592 1607 3626 1641
rect 3660 1608 3696 1641
rect 3660 1607 3730 1608
rect 3438 1574 3730 1607
rect 3438 1572 3696 1574
rect 3438 1538 3490 1572
rect 3524 1538 3558 1572
rect 3592 1538 3626 1572
rect 3660 1540 3696 1572
rect 3660 1538 3730 1540
rect 3438 1506 3730 1538
rect 3438 1503 3696 1506
rect 3438 1469 3490 1503
rect 3524 1469 3558 1503
rect 3592 1469 3626 1503
rect 3660 1472 3696 1503
rect 3660 1469 3730 1472
rect 3438 1438 3730 1469
rect 3438 1434 3696 1438
rect 3438 1400 3490 1434
rect 3524 1400 3558 1434
rect 3592 1400 3626 1434
rect 3660 1404 3696 1434
rect 4266 1920 4300 1950
rect 4266 1863 4300 1886
rect 4266 1784 4300 1818
rect 4266 1716 4300 1750
rect 4266 1648 4300 1682
rect 4266 1580 4300 1614
rect 4266 1512 4300 1546
rect 4266 1444 4300 1478
rect 3660 1400 3730 1404
rect 3438 1370 3730 1400
rect 3438 1365 3696 1370
rect 3438 1331 3490 1365
rect 3524 1331 3558 1365
rect 3592 1331 3626 1365
rect 3660 1336 3696 1365
rect 3660 1331 3730 1336
rect 3438 1302 3730 1331
rect 3438 1296 3696 1302
rect 3438 1262 3490 1296
rect 3524 1262 3558 1296
rect 3592 1262 3626 1296
rect 3660 1268 3696 1296
rect 3660 1262 3730 1268
rect 3438 1234 3730 1262
rect 3438 1227 3696 1234
rect 3438 1193 3490 1227
rect 3524 1193 3558 1227
rect 3592 1193 3626 1227
rect 3660 1200 3696 1227
rect 3660 1193 3730 1200
rect 3438 1166 3730 1193
rect 3438 1158 3696 1166
rect 3438 1124 3490 1158
rect 3524 1124 3558 1158
rect 3592 1124 3626 1158
rect 3660 1132 3696 1158
rect 3660 1124 3730 1132
rect 3438 1098 3730 1124
rect 3438 1089 3696 1098
rect 3438 1055 3490 1089
rect 3524 1055 3558 1089
rect 3592 1055 3626 1089
rect 3660 1064 3696 1089
rect 3660 1055 3730 1064
rect 3438 1030 3730 1055
rect 3438 1020 3696 1030
rect 3438 374 3490 1020
rect 3660 996 3696 1020
rect 3660 962 3730 996
rect 3660 928 3696 962
rect 3660 894 3730 928
rect 3660 860 3696 894
rect 3660 826 3730 860
rect 3660 792 3696 826
rect 3660 758 3730 792
rect 3660 724 3696 758
rect 3660 690 3730 724
rect 3660 656 3696 690
rect 3660 622 3730 656
rect 3660 588 3696 622
rect 3660 554 3730 588
rect 3660 520 3696 554
rect 4140 1400 4174 1409
rect 4140 1319 4174 1359
rect 4140 1245 4174 1279
rect 4140 1171 4174 1191
rect 4140 1097 4174 1103
rect 4140 1023 4174 1063
rect 4140 949 4174 989
rect 4140 875 4174 915
rect 4140 801 4174 841
rect 4140 727 4174 767
rect 4140 653 4174 693
rect 4140 579 4174 619
rect 4140 529 4174 545
rect 4266 1376 4300 1410
rect 4266 1308 4300 1330
rect 4266 1250 4300 1274
rect 4266 1172 4300 1206
rect 4266 1104 4300 1138
rect 4266 1036 4300 1070
rect 4266 968 4300 1002
rect 4266 900 4300 934
rect 4266 832 4300 866
rect 4266 764 4300 798
rect 4266 696 4300 730
rect 4266 628 4300 658
rect 4266 560 4300 582
rect 3660 486 3730 520
rect 3660 452 3696 486
rect 3660 418 3730 452
rect 3660 384 3696 418
rect 4266 492 4300 506
rect 3660 377 3824 384
rect 3858 377 3892 384
rect 3926 377 3960 384
rect 3994 377 4028 384
rect 3660 374 3738 377
rect 3268 343 3738 374
rect 3772 343 3810 377
rect 3858 350 3882 377
rect 3926 350 3954 377
rect 3994 350 4026 377
rect 4062 350 4096 384
rect 4130 377 4164 384
rect 4132 350 4164 377
rect 4198 350 4232 384
rect 4266 350 4300 431
rect 3844 343 3882 350
rect 3916 343 3954 350
rect 3988 343 4026 350
rect 4060 343 4098 350
rect 4132 343 4300 350
rect 3268 341 4300 343
rect 4645 4521 4681 4528
rect 4645 4487 4646 4521
rect 4680 4487 4681 4521
rect 4645 4453 4681 4487
rect 4645 4419 4646 4453
rect 4680 4419 4681 4453
rect 4645 4402 4681 4419
rect 4645 4351 4646 4402
rect 4680 4351 4681 4402
rect 4645 4317 4681 4351
rect 4645 4265 4646 4317
rect 4680 4265 4681 4317
rect 4645 4249 4681 4265
rect 4645 4215 4646 4249
rect 4680 4215 4681 4249
rect 4645 4196 4681 4215
rect 4645 4147 4646 4196
rect 4680 4147 4681 4196
rect 4645 4113 4681 4147
rect 4645 4079 4646 4113
rect 4680 4079 4681 4113
rect 4645 4045 4681 4079
rect 4645 3990 4646 4045
rect 4680 3990 4681 4045
rect 4645 3977 4681 3990
rect 4645 3910 4646 3977
rect 4680 3910 4681 3977
rect 4645 3909 4681 3910
rect 4645 3875 4646 3909
rect 4680 3875 4681 3909
rect 4645 3864 4681 3875
rect 4645 3807 4646 3864
rect 4680 3807 4681 3864
rect 4645 3785 4681 3807
rect 4645 3739 4646 3785
rect 4680 3739 4681 3785
rect 4645 3706 4681 3739
rect 4645 3671 4646 3706
rect 4680 3671 4681 3706
rect 4645 3637 4681 3671
rect 4645 3593 4646 3637
rect 4680 3593 4681 3637
rect 4645 3569 4681 3593
rect 4645 3514 4646 3569
rect 4680 3514 4681 3569
rect 4645 3501 4681 3514
rect 4645 3467 4646 3501
rect 4680 3467 4681 3501
rect 4645 3433 4681 3467
rect 4645 3399 4646 3433
rect 4680 3399 4681 3433
rect 4645 3388 4681 3399
rect 4645 3331 4646 3388
rect 4680 3331 4681 3388
rect 4645 3309 4681 3331
rect 4645 3263 4646 3309
rect 4680 3263 4681 3309
rect 4645 3230 4681 3263
rect 4645 3195 4646 3230
rect 4680 3195 4681 3230
rect 4645 3161 4681 3195
rect 4645 3127 4646 3161
rect 4680 3127 4681 3161
rect 4645 3093 4681 3127
rect 4645 3036 4646 3093
rect 4680 3036 4681 3093
rect 4645 3025 4681 3036
rect 4645 2960 4646 3025
rect 4680 2960 4681 3025
rect 4645 2957 4681 2960
rect 4645 2923 4646 2957
rect 4680 2923 4681 2957
rect 4645 2918 4681 2923
rect 4645 2855 4646 2918
rect 4680 2855 4681 2918
rect 4645 2842 4681 2855
rect 4645 2787 4646 2842
rect 4680 2787 4681 2842
rect 4645 2766 4681 2787
rect 4645 2719 4646 2766
rect 4680 2719 4681 2766
rect 4645 2690 4681 2719
rect 4645 2651 4646 2690
rect 4680 2651 4681 2690
rect 4645 2617 4681 2651
rect 4645 2580 4646 2617
rect 4680 2580 4681 2617
rect 4645 2549 4681 2580
rect 4645 2504 4646 2549
rect 4680 2504 4681 2549
rect 4645 2481 4681 2504
rect 4645 2428 4646 2481
rect 4680 2428 4681 2481
rect 4645 2413 4681 2428
rect 4645 2379 4646 2413
rect 4680 2379 4681 2413
rect 4645 2345 4681 2379
rect 4645 2311 4646 2345
rect 4680 2311 4681 2345
rect 4645 2277 4681 2311
rect 4645 2243 4646 2277
rect 4680 2243 4681 2277
rect 4645 2209 4681 2243
rect 4645 2175 4646 2209
rect 4680 2175 4681 2209
rect 4645 2141 4681 2175
rect 4645 2107 4646 2141
rect 4680 2107 4681 2141
rect 4645 2073 4681 2107
rect 4645 2039 4646 2073
rect 4680 2039 4681 2073
rect 4645 2005 4681 2039
rect 4645 1971 4646 2005
rect 4680 1971 4681 2005
rect 4645 1937 4681 1971
rect 4645 1903 4646 1937
rect 4680 1903 4681 1937
rect 4645 1869 4681 1903
rect 4645 1835 4646 1869
rect 4680 1835 4681 1869
rect 4645 1801 4681 1835
rect 4645 1767 4646 1801
rect 4680 1767 4681 1801
rect 4645 1733 4681 1767
rect 4645 1699 4646 1733
rect 4680 1699 4681 1733
rect 4645 1681 4681 1699
rect 4645 1631 4646 1681
rect 4680 1631 4681 1681
rect 4645 1600 4681 1631
rect 4645 1563 4646 1600
rect 4680 1563 4681 1600
rect 4645 1529 4681 1563
rect 4645 1486 4646 1529
rect 4680 1486 4681 1529
rect 4645 1461 4681 1486
rect 4645 1406 4646 1461
rect 4680 1406 4681 1461
rect 4645 1393 4681 1406
rect 4645 1326 4646 1393
rect 4680 1326 4681 1393
rect 4645 1325 4681 1326
rect 4645 1291 4646 1325
rect 4680 1291 4681 1325
rect 4645 1257 4681 1291
rect 4645 1223 4646 1257
rect 4680 1223 4681 1257
rect 4645 1189 4681 1223
rect 4645 1155 4646 1189
rect 4680 1155 4681 1189
rect 4645 1121 4681 1155
rect 4645 1087 4646 1121
rect 4680 1087 4681 1121
rect 4645 1053 4681 1087
rect 4645 1019 4646 1053
rect 4680 1019 4681 1053
rect 4645 985 4681 1019
rect 4645 951 4646 985
rect 4680 951 4681 985
rect 4645 917 4681 951
rect 4645 883 4646 917
rect 4680 883 4681 917
rect 4645 849 4681 883
rect 4645 815 4646 849
rect 4680 815 4681 849
rect 4645 781 4681 815
rect 4645 747 4646 781
rect 4680 747 4681 781
rect 4645 713 4681 747
rect 4645 679 4646 713
rect 4680 679 4681 713
rect 4645 645 4681 679
rect 4645 611 4646 645
rect 4680 611 4681 645
rect 4645 577 4681 611
rect 4645 543 4646 577
rect 4680 543 4681 577
rect 4645 509 4681 543
rect 4645 475 4646 509
rect 4680 475 4681 509
rect 4645 448 4681 475
rect 4645 407 4646 448
rect 4680 407 4681 448
rect 4645 373 4681 407
rect 1668 334 3114 335
rect 4645 339 4646 373
rect 4680 339 4681 373
rect 4645 330 4681 339
rect 4645 271 4646 330
rect 4680 271 4681 330
rect 4645 237 4681 271
rect 4645 203 4646 237
rect 4680 203 4681 237
rect 4834 5086 4841 5118
rect 4875 5117 4913 5120
rect 4947 5117 4985 5120
rect 5019 5117 5057 5120
rect 5091 5117 5129 5120
rect 5163 5117 5201 5120
rect 5235 5117 5273 5120
rect 5307 5117 5345 5120
rect 5379 5117 5417 5120
rect 5451 5117 5489 5120
rect 5523 5117 5561 5120
rect 5595 5117 5633 5120
rect 5667 5117 5705 5120
rect 5739 5117 5777 5120
rect 5811 5117 5849 5120
rect 5883 5117 5921 5120
rect 5955 5117 5993 5120
rect 6027 5117 6065 5120
rect 6099 5117 6137 5120
rect 6171 5117 6209 5120
rect 6243 5117 6281 5120
rect 6315 5117 6353 5120
rect 6387 5117 6425 5120
rect 6459 5117 6497 5120
rect 6531 5117 6569 5120
rect 6603 5117 6641 5120
rect 6675 5117 6713 5120
rect 6747 5117 6785 5120
rect 6819 5117 6858 5120
rect 6892 5117 6931 5120
rect 6965 5117 7004 5120
rect 7038 5117 7077 5120
rect 7111 5117 7150 5120
rect 7184 5117 7223 5120
rect 7257 5117 7296 5120
rect 7330 5117 7369 5120
rect 7403 5117 7442 5120
rect 7476 5117 7515 5120
rect 7549 5117 7588 5120
rect 7622 5117 7661 5120
rect 7695 5117 7734 5120
rect 7768 5117 7807 5120
rect 7841 5117 7880 5120
rect 7914 5117 7953 5120
rect 7987 5117 8026 5120
rect 8060 5117 8099 5120
rect 8133 5117 8172 5120
rect 8206 5117 8245 5120
rect 8279 5117 8318 5120
rect 8352 5117 8391 5120
rect 8425 5117 8464 5120
rect 8498 5117 8537 5120
rect 8571 5117 8610 5120
rect 8644 5117 8683 5120
rect 8717 5117 8756 5120
rect 8790 5117 8829 5120
rect 8863 5117 8902 5120
rect 8936 5117 8975 5120
rect 9009 5117 9048 5120
rect 9082 5117 9121 5120
rect 9155 5117 9194 5120
rect 9228 5117 9267 5120
rect 9301 5117 9340 5120
rect 9374 5117 9413 5120
rect 9447 5117 12710 5118
rect 4902 5086 4913 5117
rect 4970 5086 4985 5117
rect 5038 5086 5057 5117
rect 5106 5086 5129 5117
rect 5174 5086 5201 5117
rect 5242 5086 5273 5117
rect 4834 5083 4868 5086
rect 4902 5083 4936 5086
rect 4970 5083 5004 5086
rect 5038 5083 5072 5086
rect 5106 5083 5140 5086
rect 5174 5083 5208 5086
rect 5242 5083 5276 5086
rect 5310 5083 5344 5117
rect 5379 5086 5412 5117
rect 5451 5086 5480 5117
rect 5523 5086 5548 5117
rect 5595 5086 5616 5117
rect 5667 5086 5684 5117
rect 5739 5086 5752 5117
rect 5811 5086 5820 5117
rect 5883 5086 5888 5117
rect 5955 5086 5956 5117
rect 5378 5083 5412 5086
rect 5446 5083 5480 5086
rect 5514 5083 5548 5086
rect 5582 5083 5616 5086
rect 5650 5083 5684 5086
rect 5718 5083 5752 5086
rect 5786 5083 5820 5086
rect 5854 5083 5888 5086
rect 5922 5083 5956 5086
rect 5990 5086 5993 5117
rect 6058 5086 6065 5117
rect 6126 5086 6137 5117
rect 6194 5086 6209 5117
rect 6262 5086 6281 5117
rect 6330 5086 6353 5117
rect 6398 5086 6425 5117
rect 6466 5086 6497 5117
rect 5990 5083 6024 5086
rect 6058 5083 6092 5086
rect 6126 5083 6160 5086
rect 6194 5083 6228 5086
rect 6262 5083 6296 5086
rect 6330 5083 6364 5086
rect 6398 5083 6432 5086
rect 6466 5083 6500 5086
rect 6534 5083 6568 5117
rect 6603 5086 6636 5117
rect 6675 5086 6704 5117
rect 6747 5086 6772 5117
rect 6819 5086 6840 5117
rect 6892 5086 6908 5117
rect 6965 5086 6976 5117
rect 7038 5086 7044 5117
rect 7111 5086 7112 5117
rect 6602 5083 6636 5086
rect 6670 5083 6704 5086
rect 6738 5083 6772 5086
rect 6806 5083 6840 5086
rect 6874 5083 6908 5086
rect 6942 5083 6976 5086
rect 7010 5083 7044 5086
rect 7078 5083 7112 5086
rect 7146 5086 7150 5117
rect 7214 5086 7223 5117
rect 7282 5086 7296 5117
rect 7350 5086 7369 5117
rect 7418 5086 7442 5117
rect 7486 5086 7515 5117
rect 7146 5083 7180 5086
rect 7214 5083 7248 5086
rect 7282 5083 7316 5086
rect 7350 5083 7384 5086
rect 7418 5083 7452 5086
rect 7486 5083 7520 5086
rect 7554 5083 7588 5117
rect 7622 5083 7656 5117
rect 7695 5086 7724 5117
rect 7768 5086 7792 5117
rect 7841 5086 7860 5117
rect 7914 5086 7928 5117
rect 7987 5086 7996 5117
rect 8060 5086 8064 5117
rect 7690 5083 7724 5086
rect 7758 5083 7792 5086
rect 7826 5083 7860 5086
rect 7894 5083 7928 5086
rect 7962 5083 7996 5086
rect 8030 5083 8064 5086
rect 8098 5086 8099 5117
rect 8166 5086 8172 5117
rect 8234 5086 8245 5117
rect 8302 5086 8318 5117
rect 8370 5086 8391 5117
rect 8438 5086 8464 5117
rect 8506 5086 8537 5117
rect 8098 5083 8132 5086
rect 8166 5083 8200 5086
rect 8234 5083 8268 5086
rect 8302 5083 8336 5086
rect 8370 5083 8404 5086
rect 8438 5083 8472 5086
rect 8506 5083 8540 5086
rect 8574 5083 8608 5117
rect 8644 5086 8676 5117
rect 8717 5086 8744 5117
rect 8790 5086 8812 5117
rect 8863 5086 8880 5117
rect 8936 5086 8948 5117
rect 9009 5086 9016 5117
rect 9082 5086 9084 5117
rect 8642 5083 8676 5086
rect 8710 5083 8744 5086
rect 8778 5083 8812 5086
rect 8846 5083 8880 5086
rect 8914 5083 8948 5086
rect 8982 5083 9016 5086
rect 9050 5083 9084 5086
rect 9118 5086 9121 5117
rect 9186 5086 9194 5117
rect 9254 5086 9267 5117
rect 9322 5086 9340 5117
rect 9390 5086 9413 5117
rect 9118 5083 9152 5086
rect 9186 5083 9220 5086
rect 9254 5083 9288 5086
rect 9322 5083 9356 5086
rect 9390 5083 9424 5086
rect 9458 5083 9492 5117
rect 9540 5083 9560 5117
rect 9614 5083 9628 5117
rect 9688 5083 9696 5117
rect 9762 5083 9764 5117
rect 9798 5083 9802 5117
rect 9866 5083 9876 5117
rect 9934 5083 9950 5117
rect 10002 5083 10024 5117
rect 10070 5083 10098 5117
rect 10138 5083 10172 5117
rect 10206 5083 10240 5117
rect 10280 5083 10308 5117
rect 10354 5083 10376 5117
rect 10428 5083 10444 5117
rect 10502 5083 10512 5117
rect 10576 5083 10580 5117
rect 10614 5083 10616 5117
rect 10682 5083 10690 5117
rect 10750 5083 10764 5117
rect 10818 5083 10838 5117
rect 10886 5083 10912 5117
rect 10954 5083 10986 5117
rect 11022 5083 11056 5117
rect 11094 5083 11124 5117
rect 11168 5083 11192 5117
rect 11241 5083 11260 5117
rect 11314 5083 11328 5117
rect 11387 5083 11396 5117
rect 11430 5083 11464 5117
rect 11498 5083 11532 5117
rect 11566 5083 11600 5117
rect 11643 5083 11668 5117
rect 11717 5083 11736 5117
rect 11791 5083 11804 5117
rect 11866 5083 11872 5117
rect 11906 5083 11907 5117
rect 11974 5083 11982 5117
rect 12042 5083 12057 5117
rect 12110 5083 12132 5117
rect 12178 5083 12207 5117
rect 12246 5083 12280 5117
rect 12316 5083 12348 5117
rect 12391 5083 12416 5117
rect 12466 5083 12484 5117
rect 12541 5083 12552 5117
rect 12586 5106 12710 5117
rect 12586 5083 12675 5106
rect 4834 5082 12675 5083
rect 4834 5037 4870 5082
rect 4834 4990 4835 5037
rect 4869 4990 4870 5037
rect 4834 4969 4870 4990
rect 4834 4918 4835 4969
rect 4869 4918 4870 4969
rect 4834 4901 4870 4918
rect 4834 4867 4835 4901
rect 4869 4867 4870 4901
rect 4834 4833 4870 4867
rect 4834 4799 4835 4833
rect 4869 4799 4870 4833
rect 4834 4771 4870 4799
rect 4834 4731 4835 4771
rect 4869 4731 4870 4771
rect 4834 4697 4870 4731
rect 4834 4656 4835 4697
rect 4869 4656 4870 4697
rect 4834 4629 4870 4656
rect 4834 4576 4835 4629
rect 4869 4576 4870 4629
rect 4834 4561 4870 4576
rect 4834 4496 4835 4561
rect 4869 4496 4870 4561
rect 4834 4493 4870 4496
rect 4834 4459 4835 4493
rect 4869 4459 4870 4493
rect 4834 4450 4870 4459
rect 4834 4391 4835 4450
rect 4869 4391 4870 4450
rect 4834 4370 4870 4391
rect 4834 4323 4835 4370
rect 4869 4323 4870 4370
rect 4834 4290 4870 4323
rect 4834 4255 4835 4290
rect 4869 4255 4870 4290
rect 4834 4221 4870 4255
rect 4834 4176 4835 4221
rect 4869 4176 4870 4221
rect 4834 4153 4870 4176
rect 4834 4119 4835 4153
rect 4869 4119 4870 4153
rect 4834 4085 4870 4119
rect 4834 4051 4835 4085
rect 4869 4051 4870 4085
rect 4834 4017 4870 4051
rect 4834 3983 4835 4017
rect 4869 3983 4870 4017
rect 4834 3949 4870 3983
rect 4834 3915 4835 3949
rect 4869 3915 4870 3949
rect 4834 3881 4870 3915
rect 4834 3847 4835 3881
rect 4869 3847 4870 3881
rect 4834 3813 4870 3847
rect 4834 3779 4835 3813
rect 4869 3779 4870 3813
rect 4834 3745 4870 3779
rect 9467 5005 9503 5082
rect 9467 4953 9468 5005
rect 9502 4953 9503 5005
rect 10296 5046 10330 5082
rect 9467 4932 9503 4953
rect 9467 4885 9468 4932
rect 9502 4885 9503 4932
rect 9692 4953 9708 4987
rect 9742 4953 9776 4987
rect 9810 4953 9826 4987
rect 9692 4921 9826 4953
rect 9692 4887 9706 4921
rect 9740 4887 9778 4921
rect 9812 4887 9826 4921
rect 9928 4953 9944 4987
rect 9978 4953 10012 4987
rect 10046 4953 10062 4987
rect 9928 4921 10062 4953
rect 9928 4887 9942 4921
rect 9976 4887 10014 4921
rect 10048 4887 10062 4921
rect 10296 4978 10330 5012
rect 10296 4910 10330 4944
rect 9467 4859 9503 4885
rect 9467 4817 9468 4859
rect 9502 4817 9503 4859
rect 10296 4842 10330 4876
rect 12674 5050 12675 5082
rect 12709 5050 12710 5106
rect 13646 5080 13682 5178
rect 12674 5032 12710 5050
rect 12674 4982 12675 5032
rect 12709 4982 12710 5032
rect 12674 4958 12710 4982
rect 12674 4914 12675 4958
rect 12709 4914 12710 4958
rect 12674 4884 12710 4914
rect 9467 4786 9503 4817
rect 9467 4749 9468 4786
rect 9502 4749 9503 4786
rect 9467 4715 9503 4749
rect 9467 4679 9468 4715
rect 9502 4679 9503 4715
rect 9467 4647 9503 4679
rect 9467 4606 9468 4647
rect 9502 4606 9503 4647
rect 9467 4579 9503 4606
rect 9467 4533 9468 4579
rect 9502 4533 9503 4579
rect 9467 4511 9503 4533
rect 9467 4460 9468 4511
rect 9502 4460 9503 4511
rect 9467 4443 9503 4460
rect 9467 4387 9468 4443
rect 9502 4387 9503 4443
rect 9467 4375 9503 4387
rect 9467 4314 9468 4375
rect 9502 4314 9503 4375
rect 9467 4307 9503 4314
rect 9467 4241 9468 4307
rect 9502 4241 9503 4307
rect 9467 4239 9503 4241
rect 9467 4205 9468 4239
rect 9502 4205 9503 4239
rect 9467 4202 9503 4205
rect 9467 4137 9468 4202
rect 9502 4137 9503 4202
rect 9467 4128 9503 4137
rect 9467 4069 9468 4128
rect 9502 4069 9503 4128
rect 9467 4054 9503 4069
rect 9467 4001 9468 4054
rect 9502 4001 9503 4054
rect 9467 3980 9503 4001
rect 9467 3933 9468 3980
rect 9502 3933 9503 3980
rect 9467 3906 9503 3933
rect 9467 3865 9468 3906
rect 9502 3865 9503 3906
rect 9467 3832 9503 3865
rect 9467 3797 9468 3832
rect 9502 3797 9503 3832
rect 9467 3763 9503 3797
rect 4834 3711 4835 3745
rect 4869 3744 4870 3745
rect 8971 3744 9010 3746
rect 9044 3744 9083 3746
rect 9117 3744 9156 3746
rect 9190 3744 9229 3746
rect 9263 3744 9302 3746
rect 9336 3744 9375 3746
rect 4869 3711 4963 3744
rect 4834 3710 4963 3711
rect 4997 3710 5032 3744
rect 4834 3677 5049 3710
rect 4834 3643 4835 3677
rect 4869 3676 5049 3677
rect 4869 3643 4963 3676
rect 4834 3642 4963 3643
rect 4997 3642 5032 3676
rect 9363 3712 9375 3744
rect 9467 3744 9468 3763
rect 9409 3724 9468 3744
rect 9502 3724 9503 3763
rect 9409 3712 9503 3724
rect 9363 3695 9503 3712
rect 9363 3674 9468 3695
rect 9363 3642 9375 3674
rect 4834 3609 4870 3642
rect 8971 3640 9010 3642
rect 9044 3640 9083 3642
rect 9117 3640 9156 3642
rect 9190 3640 9229 3642
rect 9263 3640 9302 3642
rect 9336 3640 9375 3642
rect 9409 3650 9468 3674
rect 9502 3650 9503 3695
rect 9409 3642 9503 3650
rect 4834 3575 4835 3609
rect 4869 3575 4870 3609
rect 4834 3541 4870 3575
rect 4834 3507 4835 3541
rect 4869 3507 4870 3541
rect 4834 3473 4870 3507
rect 4834 3439 4835 3473
rect 4869 3468 4870 3473
rect 9467 3627 9503 3642
rect 9467 3576 9468 3627
rect 9502 3576 9503 3627
rect 9467 3559 9503 3576
rect 9467 3502 9468 3559
rect 9502 3502 9503 3559
rect 9467 3491 9503 3502
rect 9467 3468 9468 3491
rect 4869 3452 4980 3468
rect 4869 3439 4946 3452
rect 4834 3418 4946 3439
rect 4834 3405 4980 3418
rect 4834 3371 4835 3405
rect 4869 3384 4980 3405
rect 4869 3371 4946 3384
rect 4834 3350 4946 3371
rect 4834 3337 4980 3350
rect 4834 3299 4835 3337
rect 4869 3334 4980 3337
rect 9314 3457 9468 3468
rect 9502 3457 9503 3491
rect 9314 3452 9503 3457
rect 9348 3423 9503 3452
rect 9348 3418 9468 3423
rect 9314 3389 9468 3418
rect 9502 3389 9503 3423
rect 9314 3384 9503 3389
rect 9348 3355 9503 3384
rect 9348 3350 9468 3355
rect 9314 3334 9468 3350
rect 4869 3299 4870 3334
rect 4834 3269 4870 3299
rect 4834 3221 4835 3269
rect 4869 3221 4870 3269
rect 4834 3201 4870 3221
rect 4834 3143 4835 3201
rect 4869 3143 4870 3201
rect 4834 3133 4870 3143
rect 4834 3031 4835 3133
rect 4869 3031 4870 3133
rect 9467 3316 9468 3334
rect 9502 3316 9503 3355
rect 9467 3287 9503 3316
rect 9467 3227 9468 3287
rect 9502 3227 9503 3287
rect 9467 3219 9503 3227
rect 9467 3185 9468 3219
rect 9502 3185 9503 3219
rect 9467 3151 9503 3185
rect 9467 3117 9468 3151
rect 9502 3117 9503 3151
rect 4834 3021 4870 3031
rect 4834 2963 4835 3021
rect 4869 2963 4870 3021
rect 4946 3097 4980 3113
rect 4946 3058 4980 3063
rect 7004 3062 7042 3096
rect 7076 3092 7110 3108
rect 4946 3029 4958 3058
rect 4992 3024 5030 3058
rect 7076 3024 7110 3058
rect 4946 2979 4980 2995
rect 4834 2943 4870 2963
rect 4834 2895 4835 2943
rect 4869 2895 4870 2943
rect 4834 2865 4870 2895
rect 4834 2827 4835 2865
rect 4869 2827 4870 2865
rect 4834 2793 4870 2827
rect 4834 2753 4835 2793
rect 4869 2753 4870 2793
rect 4834 2725 4870 2753
rect 4946 2861 4980 2877
rect 4946 2793 4980 2827
rect 7076 2856 7110 2990
rect 7076 2788 7110 2822
rect 4946 2749 4958 2759
rect 4992 2749 5030 2783
rect 7004 2749 7042 2783
rect 4946 2743 4980 2749
rect 7076 2738 7110 2754
rect 7184 3092 7218 3108
rect 9314 3092 9348 3108
rect 7184 3024 7218 3058
rect 7252 3031 7290 3065
rect 9242 3031 9280 3065
rect 7184 2856 7218 2990
rect 9314 3024 9348 3058
rect 9314 2974 9348 2990
rect 9467 3083 9503 3117
rect 9467 3049 9468 3083
rect 9502 3049 9503 3083
rect 9467 3015 9503 3049
rect 9623 4767 9657 4806
rect 9623 4694 9657 4733
rect 9623 4621 9657 4660
rect 9623 4548 9657 4587
rect 9623 4475 9657 4514
rect 9623 4402 9657 4441
rect 9623 4329 9657 4368
rect 9623 4256 9657 4295
rect 9623 4182 9657 4222
rect 9623 4108 9657 4148
rect 9623 4034 9657 4074
rect 9623 3960 9657 4000
rect 9623 3886 9657 3926
rect 9623 3812 9657 3852
rect 9623 3738 9657 3778
rect 9623 3664 9657 3704
rect 9623 3590 9657 3630
rect 9623 3516 9657 3556
rect 9623 3442 9657 3482
rect 9623 3368 9657 3408
rect 9623 3294 9657 3334
rect 9623 3220 9657 3260
rect 9623 3146 9657 3186
rect 9623 3072 9657 3112
rect 9859 4767 9893 4806
rect 9859 4694 9893 4733
rect 9859 4621 9893 4660
rect 9859 4548 9893 4587
rect 9859 4475 9893 4514
rect 9859 4402 9893 4441
rect 9859 4329 9893 4368
rect 9859 4256 9893 4295
rect 9859 4183 9893 4222
rect 9859 4110 9893 4149
rect 9859 4037 9893 4076
rect 9859 3964 9893 4003
rect 9859 3891 9893 3930
rect 9859 3817 9893 3857
rect 9859 3743 9893 3783
rect 9859 3669 9893 3709
rect 9859 3595 9893 3635
rect 9859 3521 9893 3561
rect 9859 3447 9893 3487
rect 9859 3373 9893 3413
rect 9859 3299 9893 3339
rect 9859 3225 9893 3265
rect 9859 3151 9893 3191
rect 9859 3077 9893 3117
rect 10095 4729 10129 4767
rect 10095 4657 10129 4695
rect 10095 4585 10129 4623
rect 10095 4513 10129 4551
rect 10095 4441 10129 4479
rect 10095 4369 10129 4407
rect 10095 4297 10129 4335
rect 10095 4225 10129 4263
rect 10095 4153 10129 4191
rect 10095 4081 10129 4119
rect 10095 4009 10129 4047
rect 10095 3937 10129 3975
rect 10095 3865 10129 3903
rect 10095 3793 10129 3831
rect 10095 3721 10129 3759
rect 10095 3649 10129 3687
rect 10095 3577 10129 3615
rect 10095 3505 10129 3543
rect 10095 3433 10129 3471
rect 10095 3361 10129 3399
rect 10095 3289 10129 3327
rect 10095 3217 10129 3255
rect 10095 3145 10129 3183
rect 10095 3072 10129 3111
rect 9467 2981 9468 3015
rect 9502 2981 9503 3015
rect 9467 2947 9503 2981
rect 10095 2999 10129 3038
rect 10296 4774 10330 4808
rect 10296 4706 10330 4740
rect 10296 4638 10330 4672
rect 10296 4570 10330 4604
rect 10296 4502 10330 4536
rect 10296 4434 10330 4468
rect 10296 4366 10330 4400
rect 10296 4298 10330 4332
rect 10296 4230 10330 4264
rect 10296 4162 10330 4196
rect 10296 4094 10330 4128
rect 10423 4711 10457 4757
rect 10423 4631 10457 4677
rect 10423 4552 10457 4597
rect 10423 4473 10457 4518
rect 10423 4394 10457 4439
rect 10423 4315 10457 4360
rect 10423 4236 10457 4281
rect 10423 4157 10457 4202
rect 11130 4711 11164 4757
rect 11130 4631 11164 4677
rect 11130 4552 11164 4597
rect 11130 4473 11164 4518
rect 11130 4394 11164 4439
rect 11130 4315 11164 4360
rect 11130 4236 11164 4281
rect 11130 4157 11164 4202
rect 11274 4784 11751 4868
rect 12674 4846 12675 4884
rect 12709 4846 12710 4884
rect 12674 4812 12710 4846
rect 11274 4750 11290 4784
rect 11324 4750 11372 4784
rect 11406 4750 11454 4784
rect 11488 4750 11536 4784
rect 11570 4750 11618 4784
rect 11652 4750 11700 4784
rect 11734 4750 11751 4784
rect 11274 4708 11751 4750
rect 11274 4674 11290 4708
rect 11324 4674 11372 4708
rect 11406 4674 11454 4708
rect 11488 4674 11536 4708
rect 11570 4674 11618 4708
rect 11652 4674 11700 4708
rect 11734 4674 11751 4708
rect 11274 4632 11751 4674
rect 11274 4598 11290 4632
rect 11324 4598 11372 4632
rect 11406 4598 11454 4632
rect 11488 4598 11536 4632
rect 11570 4598 11618 4632
rect 11652 4598 11700 4632
rect 11734 4598 11751 4632
rect 11274 4555 11751 4598
rect 11274 4521 11290 4555
rect 11324 4521 11372 4555
rect 11406 4521 11454 4555
rect 11488 4521 11536 4555
rect 11570 4521 11618 4555
rect 11652 4521 11700 4555
rect 11734 4521 11751 4555
rect 11274 4478 11751 4521
rect 11274 4444 11290 4478
rect 11324 4444 11372 4478
rect 11406 4444 11454 4478
rect 11488 4444 11536 4478
rect 11570 4444 11618 4478
rect 11652 4444 11700 4478
rect 11734 4444 11751 4478
rect 11274 4401 11751 4444
rect 11274 4367 11290 4401
rect 11324 4367 11372 4401
rect 11406 4367 11454 4401
rect 11488 4367 11536 4401
rect 11570 4367 11618 4401
rect 11652 4367 11700 4401
rect 11734 4367 11751 4401
rect 11274 4324 11751 4367
rect 11274 4290 11290 4324
rect 11324 4290 11372 4324
rect 11406 4290 11454 4324
rect 11488 4290 11536 4324
rect 11570 4290 11618 4324
rect 11652 4290 11700 4324
rect 11734 4290 11751 4324
rect 11274 4247 11751 4290
rect 11274 4213 11290 4247
rect 11324 4213 11372 4247
rect 11406 4213 11454 4247
rect 11488 4213 11536 4247
rect 11570 4213 11618 4247
rect 11652 4213 11700 4247
rect 11734 4213 11751 4247
rect 11274 4170 11751 4213
rect 11274 4136 11290 4170
rect 11324 4136 11372 4170
rect 11406 4136 11454 4170
rect 11488 4136 11536 4170
rect 11570 4136 11618 4170
rect 11652 4136 11700 4170
rect 11734 4136 11751 4170
rect 10296 4026 10330 4060
rect 10296 3958 10330 3992
rect 10296 3890 10330 3924
rect 10296 3822 10330 3856
rect 10296 3754 10330 3788
rect 10296 3686 10330 3720
rect 10296 3618 10330 3652
rect 10296 3550 10330 3584
rect 10296 3482 10330 3516
rect 10296 3414 10330 3448
rect 10296 3346 10330 3380
rect 10296 3278 10330 3312
rect 10296 3210 10330 3244
rect 10296 3142 10330 3176
rect 10296 3074 10330 3108
rect 10296 3006 10330 3040
rect 9467 2913 9468 2947
rect 9502 2913 9503 2947
rect 9467 2879 9503 2913
rect 7184 2788 7218 2822
rect 9253 2856 9348 2872
rect 9253 2822 9314 2856
rect 9253 2788 9348 2822
rect 7184 2738 7218 2754
rect 7252 2751 7290 2785
rect 9181 2751 9219 2785
rect 9253 2754 9314 2788
rect 9253 2738 9348 2754
rect 9467 2845 9468 2879
rect 9502 2845 9503 2879
rect 9467 2811 9503 2845
rect 9467 2777 9468 2811
rect 9502 2777 9503 2811
rect 9467 2743 9503 2777
rect 4834 2675 4835 2725
rect 4869 2675 4870 2725
rect 4834 2657 4870 2675
rect 4834 2597 4835 2657
rect 4869 2597 4870 2657
rect 4834 2589 4870 2597
rect 4834 2555 4835 2589
rect 4869 2555 4870 2589
rect 4834 2553 4870 2555
rect 4834 2487 4835 2553
rect 4869 2487 4870 2553
rect 9467 2709 9468 2743
rect 9502 2709 9503 2743
rect 9467 2675 9503 2709
rect 9467 2641 9468 2675
rect 9502 2641 9503 2675
rect 9467 2607 9503 2641
rect 9467 2573 9468 2607
rect 9502 2573 9503 2607
rect 9467 2539 9503 2573
rect 4834 2476 4870 2487
rect 4834 2419 4835 2476
rect 4869 2419 4870 2476
rect 4834 2385 4870 2419
rect 4834 2351 4835 2385
rect 4869 2351 4870 2385
rect 4946 2494 4980 2510
rect 4946 2445 4980 2460
rect 7076 2494 7110 2510
rect 4946 2426 4958 2445
rect 4992 2411 5030 2445
rect 7076 2426 7110 2460
rect 4946 2376 4980 2392
rect 7004 2390 7042 2424
rect 4834 2317 4870 2351
rect 4834 2283 4835 2317
rect 4869 2283 4870 2317
rect 4834 2249 4870 2283
rect 4834 2215 4835 2249
rect 4869 2215 4870 2249
rect 4834 2181 4870 2215
rect 4834 2147 4835 2181
rect 4869 2147 4870 2181
rect 4834 2113 4870 2147
rect 4946 2258 5173 2274
rect 4980 2224 5173 2258
rect 4946 2207 5173 2224
rect 4946 2190 5067 2207
rect 4980 2173 5067 2190
rect 5101 2173 5139 2207
rect 7076 2258 7110 2392
rect 7076 2190 7110 2224
rect 4980 2156 5173 2173
rect 4946 2140 5173 2156
rect 7004 2152 7042 2186
rect 7076 2140 7110 2156
rect 7184 2494 7218 2510
rect 7252 2464 7290 2498
rect 9314 2494 9348 2510
rect 7184 2426 7218 2460
rect 9242 2426 9280 2460
rect 9314 2426 9348 2460
rect 7184 2258 7218 2392
rect 9314 2376 9348 2392
rect 9467 2505 9468 2539
rect 9502 2505 9503 2539
rect 9467 2471 9503 2505
rect 9467 2437 9468 2471
rect 9502 2437 9503 2471
rect 9467 2402 9503 2437
rect 9467 2368 9468 2402
rect 9502 2368 9503 2402
rect 9467 2333 9503 2368
rect 9467 2299 9468 2333
rect 9502 2299 9503 2333
rect 7184 2190 7218 2224
rect 9314 2258 9348 2274
rect 9314 2190 9348 2224
rect 7184 2140 7218 2156
rect 7252 2148 7290 2182
rect 9264 2148 9302 2182
rect 9336 2148 9348 2156
rect 9314 2140 9348 2148
rect 9467 2264 9503 2299
rect 9467 2230 9468 2264
rect 9502 2230 9503 2264
rect 9467 2195 9503 2230
rect 10296 2938 10330 2972
rect 10296 2870 10330 2904
rect 10296 2802 10330 2836
rect 10296 2734 10330 2768
rect 10296 2666 10330 2700
rect 10296 2598 10330 2632
rect 10296 2530 10330 2564
rect 10296 2462 10330 2496
rect 10296 2394 10330 2428
rect 10296 2326 10330 2360
rect 10296 2258 10330 2292
rect 9467 2161 9468 2195
rect 9502 2161 9503 2195
rect 4834 2079 4835 2113
rect 4869 2079 4870 2113
rect 4834 2045 4870 2079
rect 4834 2011 4835 2045
rect 4869 2011 4870 2045
rect 4834 1977 4870 2011
rect 4834 1943 4835 1977
rect 4869 1943 4870 1977
rect 4834 1914 4870 1943
rect 9467 2126 9503 2161
rect 9859 2152 9893 2193
rect 9467 2092 9468 2126
rect 9502 2092 9503 2126
rect 9467 2057 9503 2092
rect 9467 2023 9468 2057
rect 9502 2023 9503 2057
rect 9467 1988 9503 2023
rect 9467 1954 9468 1988
rect 9502 1954 9503 1988
rect 9467 1919 9503 1954
rect 9467 1914 9468 1919
rect 4834 1909 4980 1914
rect 4834 1875 4835 1909
rect 4869 1898 4980 1909
rect 4869 1875 4946 1898
rect 4834 1864 4946 1875
rect 4834 1841 4980 1864
rect 4834 1807 4835 1841
rect 4869 1830 4980 1841
rect 4869 1807 4946 1830
rect 4834 1796 4946 1807
rect 4834 1780 4980 1796
rect 9314 1898 9468 1914
rect 9348 1885 9468 1898
rect 9502 1885 9503 1919
rect 9348 1864 9503 1885
rect 9314 1850 9503 1864
rect 9314 1830 9468 1850
rect 9348 1816 9468 1830
rect 9502 1816 9503 1850
rect 9348 1796 9503 1816
rect 9314 1781 9503 1796
rect 9314 1780 9468 1781
rect 4834 1773 4870 1780
rect 4834 1739 4835 1773
rect 4869 1739 4870 1773
rect 4834 1705 4870 1739
rect 4834 1671 4835 1705
rect 4869 1671 4870 1705
rect 4834 1637 4870 1671
rect 4834 1603 4835 1637
rect 4869 1605 4870 1637
rect 9467 1747 9468 1780
rect 9502 1747 9503 1781
rect 9467 1712 9503 1747
rect 9467 1678 9468 1712
rect 9502 1678 9503 1712
rect 9467 1643 9503 1678
rect 9467 1609 9468 1643
rect 9502 1609 9503 1643
rect 9467 1605 9503 1609
rect 4869 1603 4963 1605
rect 4834 1571 4963 1603
rect 4997 1571 5032 1605
rect 5066 1572 5101 1605
rect 5135 1572 5170 1605
rect 5204 1572 5239 1605
rect 5273 1572 5308 1605
rect 5342 1572 5377 1605
rect 5411 1572 5446 1605
rect 5083 1571 5101 1572
rect 5155 1571 5170 1572
rect 5227 1571 5239 1572
rect 5299 1571 5308 1572
rect 5371 1571 5377 1572
rect 5443 1571 5446 1572
rect 5480 1572 5515 1605
rect 5480 1571 5481 1572
rect 4834 1569 5049 1571
rect 4834 1535 4835 1569
rect 4869 1538 5049 1569
rect 5083 1538 5121 1571
rect 5155 1538 5193 1571
rect 5227 1538 5265 1571
rect 5299 1538 5337 1571
rect 5371 1538 5409 1571
rect 5443 1538 5481 1571
rect 5549 1572 5584 1605
rect 5618 1572 5653 1605
rect 5687 1572 5722 1605
rect 5756 1572 5791 1605
rect 5825 1572 5860 1605
rect 5894 1572 5929 1605
rect 9363 1574 9503 1605
rect 9363 1572 9468 1574
rect 5549 1571 5553 1572
rect 5618 1571 5625 1572
rect 5687 1571 5697 1572
rect 5756 1571 5769 1572
rect 5825 1571 5841 1572
rect 5894 1571 5913 1572
rect 5515 1538 5553 1571
rect 5587 1538 5625 1571
rect 5659 1538 5697 1571
rect 5731 1538 5769 1571
rect 5803 1538 5841 1571
rect 5875 1538 5913 1571
rect 9363 1538 9375 1572
rect 9409 1540 9468 1572
rect 9502 1540 9503 1574
rect 9409 1538 9503 1540
rect 4869 1537 5929 1538
rect 4869 1535 4963 1537
rect 4834 1503 4963 1535
rect 4997 1503 5032 1537
rect 5066 1503 5101 1537
rect 5135 1503 5170 1537
rect 5204 1503 5239 1537
rect 5273 1503 5308 1537
rect 5342 1503 5377 1537
rect 5411 1503 5446 1537
rect 5480 1503 5515 1537
rect 5549 1503 5584 1537
rect 5618 1503 5653 1537
rect 5687 1503 5722 1537
rect 5756 1503 5791 1537
rect 5825 1503 5860 1537
rect 5894 1503 5929 1537
rect 9363 1505 9503 1538
rect 9363 1503 9468 1505
rect 4834 1501 4870 1503
rect 4834 1467 4835 1501
rect 4869 1467 4870 1501
rect 4834 1433 4870 1467
rect 4834 1399 4835 1433
rect 4869 1399 4870 1433
rect 4834 1365 4870 1399
rect 4834 1331 4835 1365
rect 4869 1331 4870 1365
rect 4834 1297 4870 1331
rect 4834 1263 4835 1297
rect 4869 1263 4870 1297
rect 4834 1229 4870 1263
rect 4834 1195 4835 1229
rect 4869 1195 4870 1229
rect 4834 1161 4870 1195
rect 4834 1127 4835 1161
rect 4869 1127 4870 1161
rect 4834 1093 4870 1127
rect 4834 1059 4835 1093
rect 4869 1059 4870 1093
rect 4834 1025 4870 1059
rect 4834 991 4835 1025
rect 4869 991 4870 1025
rect 4834 957 4870 991
rect 4834 923 4835 957
rect 4869 923 4870 957
rect 4834 889 4870 923
rect 4834 855 4835 889
rect 4869 855 4870 889
rect 4834 821 4870 855
rect 4834 787 4835 821
rect 4869 787 4870 821
rect 4834 753 4870 787
rect 4834 719 4835 753
rect 4869 719 4870 753
rect 4834 685 4870 719
rect 4834 651 4835 685
rect 4869 651 4870 685
rect 4834 617 4870 651
rect 4834 583 4835 617
rect 4869 583 4870 617
rect 4834 549 4870 583
rect 4834 515 4835 549
rect 4869 515 4870 549
rect 4834 481 4870 515
rect 4834 447 4835 481
rect 4869 447 4870 481
rect 4834 436 4870 447
rect 4834 379 4835 436
rect 4869 379 4870 436
rect 4834 345 4870 379
rect 4834 294 4835 345
rect 4869 294 4870 345
rect 4834 277 4870 294
rect 4834 243 4835 277
rect 4869 245 4870 277
rect 9467 1468 9468 1503
rect 9502 1468 9503 1505
rect 9467 1436 9503 1468
rect 9467 1394 9468 1436
rect 9502 1394 9503 1436
rect 9467 1367 9503 1394
rect 9467 1320 9468 1367
rect 9502 1320 9503 1367
rect 9467 1298 9503 1320
rect 9467 1246 9468 1298
rect 9502 1246 9503 1298
rect 9467 1229 9503 1246
rect 9467 1172 9468 1229
rect 9502 1172 9503 1229
rect 9467 1160 9503 1172
rect 9467 1098 9468 1160
rect 9502 1098 9503 1160
rect 9467 1091 9503 1098
rect 9467 1024 9468 1091
rect 9502 1024 9503 1091
rect 9467 1022 9503 1024
rect 9467 988 9468 1022
rect 9502 988 9503 1022
rect 9467 984 9503 988
rect 9467 919 9468 984
rect 9502 919 9503 984
rect 9467 910 9503 919
rect 9467 850 9468 910
rect 9502 850 9503 910
rect 9467 836 9503 850
rect 9467 781 9468 836
rect 9502 781 9503 836
rect 9467 763 9503 781
rect 9467 712 9468 763
rect 9502 712 9503 763
rect 9467 690 9503 712
rect 9467 643 9468 690
rect 9502 643 9503 690
rect 9623 2062 9657 2102
rect 9623 1988 9657 2028
rect 9623 1914 9657 1954
rect 9623 1840 9657 1880
rect 9623 1766 9657 1806
rect 9623 1692 9657 1732
rect 9623 1618 9657 1658
rect 9623 1544 9657 1584
rect 9623 1470 9657 1510
rect 9623 1395 9657 1436
rect 9623 1320 9657 1361
rect 9623 1245 9657 1286
rect 9623 1170 9657 1211
rect 9623 1095 9657 1136
rect 9623 1020 9657 1061
rect 9623 945 9657 986
rect 9623 870 9657 911
rect 9623 795 9657 836
rect 9623 720 9657 761
rect 9859 2077 9893 2118
rect 10296 2190 10330 2224
rect 10296 2122 10330 2156
rect 9859 2002 9893 2043
rect 9859 1927 9893 1968
rect 9859 1852 9893 1893
rect 9859 1777 9893 1818
rect 9859 1702 9893 1743
rect 9859 1627 9893 1668
rect 9859 1552 9893 1593
rect 9859 1477 9893 1518
rect 9859 1402 9893 1443
rect 9859 1327 9893 1368
rect 9859 1252 9893 1293
rect 9859 1176 9893 1218
rect 9859 1100 9893 1142
rect 9859 1024 9893 1066
rect 9859 948 9893 990
rect 9859 872 9893 914
rect 9859 796 9893 838
rect 9859 720 9893 762
rect 10095 1989 10129 2029
rect 10095 1915 10129 1955
rect 10095 1841 10129 1881
rect 10095 1767 10129 1807
rect 10095 1693 10129 1733
rect 10095 1619 10129 1659
rect 10095 1545 10129 1585
rect 10095 1470 10129 1511
rect 10095 1395 10129 1436
rect 10095 1320 10129 1361
rect 10095 1245 10129 1286
rect 10095 1170 10129 1211
rect 10095 1095 10129 1136
rect 10095 1020 10129 1061
rect 10095 945 10129 986
rect 10095 870 10129 911
rect 10095 795 10129 836
rect 10095 720 10129 761
rect 10296 2054 10330 2088
rect 10296 1986 10330 2020
rect 10296 1918 10330 1952
rect 10296 1850 10330 1884
rect 10296 1782 10330 1816
rect 10296 1714 10330 1748
rect 10296 1646 10330 1680
rect 10296 1578 10330 1612
rect 10296 1510 10330 1544
rect 10296 1442 10330 1476
rect 10400 3954 10434 4084
rect 10400 3884 10434 3918
rect 10400 3698 10434 3848
rect 11130 3954 11164 4084
rect 11130 3884 11164 3918
rect 10654 3756 10692 3790
rect 10726 3756 10764 3790
rect 10798 3756 10836 3790
rect 10870 3756 10908 3790
rect 10942 3756 10980 3790
rect 11014 3756 11052 3790
rect 10400 3628 10434 3662
rect 10400 3442 10434 3592
rect 10400 3372 10434 3406
rect 10400 3184 10434 3336
rect 11130 3698 11164 3848
rect 11274 3790 11751 4136
rect 11860 4711 11894 4757
rect 11860 4631 11894 4677
rect 11860 4552 11894 4597
rect 11860 4473 11894 4518
rect 11860 4394 11894 4439
rect 11860 4315 11894 4360
rect 11860 4236 11894 4281
rect 11860 4157 11894 4202
rect 12565 4711 12599 4757
rect 12565 4631 12599 4677
rect 12565 4552 12599 4597
rect 12565 4473 12599 4518
rect 12565 4394 12599 4439
rect 12565 4315 12599 4360
rect 12565 4236 12599 4281
rect 12565 4157 12599 4202
rect 12674 4776 12675 4812
rect 12709 4776 12710 4812
rect 12674 4744 12710 4776
rect 12674 4702 12675 4744
rect 12709 4702 12710 4744
rect 12674 4676 12710 4702
rect 12674 4628 12675 4676
rect 12709 4628 12710 4676
rect 12674 4608 12710 4628
rect 12674 4554 12675 4608
rect 12709 4554 12710 4608
rect 12674 4540 12710 4554
rect 12674 4480 12675 4540
rect 12709 4480 12710 4540
rect 12674 4472 12710 4480
rect 12674 4406 12675 4472
rect 12709 4406 12710 4472
rect 12674 4365 12710 4406
rect 12674 4331 12675 4365
rect 12709 4331 12710 4365
rect 12674 4290 12710 4331
rect 12674 4256 12675 4290
rect 12709 4256 12710 4290
rect 12674 4215 12710 4256
rect 12674 4181 12675 4215
rect 12709 4181 12710 4215
rect 12674 4140 12710 4181
rect 12674 4106 12675 4140
rect 12709 4106 12710 4140
rect 11130 3628 11164 3662
rect 11130 3442 11164 3592
rect 11130 3372 11164 3406
rect 10654 3244 10692 3278
rect 10726 3244 10764 3278
rect 10798 3244 10836 3278
rect 10870 3244 10908 3278
rect 10942 3244 10980 3278
rect 11014 3244 11052 3278
rect 10400 3116 10434 3150
rect 11130 3184 11164 3336
rect 11130 3116 11164 3150
rect 11860 3442 11894 4084
rect 12674 4065 12710 4106
rect 12674 4031 12675 4065
rect 12709 4031 12710 4065
rect 12674 3990 12710 4031
rect 12674 3956 12675 3990
rect 12709 3956 12710 3990
rect 12674 3915 12710 3956
rect 12590 3892 12624 3908
rect 12590 3829 12624 3858
rect 12674 3881 12675 3915
rect 12709 3881 12710 3915
rect 12590 3824 12592 3829
rect 12624 3790 12626 3795
rect 12590 3756 12626 3790
rect 12590 3688 12624 3722
rect 12590 3638 12624 3654
rect 12674 3670 12710 3881
rect 12674 3636 12675 3670
rect 12709 3636 12710 3670
rect 12674 3590 12710 3636
rect 12674 3556 12675 3590
rect 12709 3556 12710 3590
rect 11860 3372 11894 3406
rect 11860 3184 11894 3336
rect 12590 3442 12624 3512
rect 12590 3372 12624 3406
rect 12042 3244 12080 3278
rect 12114 3244 12152 3278
rect 12186 3244 12224 3278
rect 12258 3244 12296 3278
rect 12330 3244 12368 3278
rect 11860 3116 11894 3150
rect 10400 3058 10434 3082
rect 11080 3066 11118 3100
rect 11152 3066 11164 3082
rect 11810 3066 11848 3100
rect 11882 3066 11894 3082
rect 10400 2986 10434 3024
rect 10400 2928 10434 2952
rect 11130 2944 11164 3066
rect 11860 2944 11894 3066
rect 11080 2910 11118 2944
rect 11152 2928 11164 2944
rect 11810 2910 11848 2944
rect 11882 2928 11894 2944
rect 10400 2860 10434 2894
rect 10400 2672 10434 2826
rect 11130 2860 11164 2894
rect 10654 2732 10692 2766
rect 10726 2732 10764 2766
rect 10798 2732 10836 2766
rect 10870 2732 10908 2766
rect 10942 2732 10980 2766
rect 11014 2732 11052 2766
rect 10400 2604 10434 2638
rect 11130 2672 11164 2826
rect 11130 2604 11164 2638
rect 11860 2860 11894 2894
rect 11860 2672 11894 2826
rect 12590 3186 12624 3336
rect 12590 3116 12624 3150
rect 12590 2928 12624 3080
rect 12590 2860 12624 2894
rect 12590 2802 12624 2826
rect 12674 3510 12710 3556
rect 12674 3476 12675 3510
rect 12709 3476 12710 3510
rect 12674 3430 12710 3476
rect 12674 3396 12675 3430
rect 12709 3396 12710 3430
rect 12674 3350 12710 3396
rect 12674 3316 12675 3350
rect 12709 3316 12710 3350
rect 12674 3270 12710 3316
rect 12674 3236 12675 3270
rect 12709 3236 12710 3270
rect 12674 3190 12710 3236
rect 12674 3156 12675 3190
rect 12709 3156 12710 3190
rect 12674 3109 12710 3156
rect 12674 3075 12675 3109
rect 12709 3075 12710 3109
rect 12674 3028 12710 3075
rect 12674 2994 12675 3028
rect 12709 2994 12710 3028
rect 12674 2789 12710 2994
rect 12042 2732 12080 2766
rect 12114 2732 12152 2766
rect 12186 2732 12224 2766
rect 12258 2732 12296 2766
rect 12330 2732 12368 2766
rect 12402 2732 12440 2766
rect 11860 2604 11894 2638
rect 10400 2546 10434 2570
rect 11080 2554 11118 2588
rect 11152 2554 11164 2570
rect 11810 2554 11848 2588
rect 11882 2554 11894 2570
rect 10400 2474 10434 2512
rect 10400 2416 10434 2440
rect 11130 2432 11164 2554
rect 11860 2432 11894 2554
rect 11080 2398 11118 2432
rect 11152 2416 11164 2432
rect 11810 2398 11848 2432
rect 11882 2416 11894 2432
rect 10400 2348 10434 2382
rect 10400 2277 10434 2314
rect 11130 2348 11164 2382
rect 10400 2205 10434 2243
rect 10654 2220 10692 2254
rect 10726 2220 10764 2254
rect 10798 2220 10836 2254
rect 10870 2220 10908 2254
rect 10942 2220 10980 2254
rect 11014 2220 11052 2254
rect 10400 2160 10434 2171
rect 10400 2092 10434 2126
rect 10400 1906 10434 2058
rect 10400 1836 10434 1870
rect 10400 1650 10434 1800
rect 11130 2160 11164 2314
rect 11130 2092 11164 2126
rect 11130 1906 11164 2058
rect 11860 2348 11894 2382
rect 11860 2160 11894 2314
rect 12590 2730 12624 2768
rect 12590 2672 12624 2696
rect 12590 2604 12624 2638
rect 12042 2220 12080 2254
rect 12114 2220 12152 2254
rect 12186 2220 12224 2254
rect 12258 2220 12296 2254
rect 12330 2220 12368 2254
rect 11860 2092 11894 2126
rect 11860 2042 11894 2058
rect 12590 2160 12624 2570
rect 12704 2755 12710 2789
rect 12670 2706 12710 2755
rect 12704 2672 12710 2706
rect 12670 2622 12710 2672
rect 12704 2588 12710 2622
rect 12670 2538 12710 2588
rect 12704 2504 12710 2538
rect 12590 2092 12624 2126
rect 12590 2040 12624 2058
rect 12674 2249 12710 2504
rect 12674 2215 12675 2249
rect 12709 2215 12710 2249
rect 12674 2174 12710 2215
rect 12674 2140 12675 2174
rect 12709 2140 12710 2174
rect 12674 2099 12710 2140
rect 12674 2065 12675 2099
rect 12709 2065 12710 2099
rect 12674 2024 12710 2065
rect 11130 1836 11164 1870
rect 10654 1708 10692 1742
rect 10726 1708 10764 1742
rect 10798 1708 10836 1742
rect 10870 1708 10908 1742
rect 10942 1708 10980 1742
rect 11014 1708 11052 1742
rect 10400 1580 10434 1614
rect 10400 1414 10434 1544
rect 11130 1650 11164 1800
rect 11130 1580 11164 1614
rect 11130 1414 11164 1544
rect 10296 1374 10330 1408
rect 10296 1306 10330 1340
rect 10296 1238 10330 1272
rect 10296 1170 10330 1204
rect 10296 1102 10330 1136
rect 10296 1034 10330 1068
rect 10296 966 10330 1000
rect 10296 898 10330 932
rect 10296 830 10330 864
rect 10296 762 10330 796
rect 10296 694 10330 728
rect 10423 1295 10457 1341
rect 10423 1215 10457 1261
rect 10423 1136 10457 1181
rect 10423 1057 10457 1102
rect 10423 978 10457 1023
rect 10423 899 10457 944
rect 10423 820 10457 865
rect 10423 741 10457 786
rect 11130 1295 11164 1341
rect 11130 1215 11164 1261
rect 11130 1136 11164 1181
rect 11130 1057 11164 1102
rect 11130 978 11164 1023
rect 11130 899 11164 944
rect 11130 820 11164 865
rect 11130 741 11164 786
rect 9467 617 9503 643
rect 9467 574 9468 617
rect 9502 574 9503 617
rect 10296 626 10330 660
rect 9467 544 9503 574
rect 9692 570 9706 604
rect 9742 570 9776 604
rect 9812 570 9826 604
rect 9928 571 9942 605
rect 9978 571 10012 605
rect 10048 571 10062 605
rect 11274 593 11763 1998
rect 12674 1990 12675 2024
rect 12709 1990 12710 2024
rect 12674 1949 12710 1990
rect 12590 1906 12624 1920
rect 12590 1836 12624 1870
rect 12590 1650 12624 1800
rect 12590 1580 12624 1614
rect 12590 1528 12624 1544
rect 12674 1915 12675 1949
rect 12709 1915 12710 1949
rect 12674 1874 12710 1915
rect 12674 1840 12675 1874
rect 12709 1840 12710 1874
rect 12674 1799 12710 1840
rect 12674 1765 12675 1799
rect 12709 1765 12710 1799
rect 12674 1724 12710 1765
rect 12674 1690 12675 1724
rect 12709 1690 12710 1724
rect 12674 1649 12710 1690
rect 12674 1615 12675 1649
rect 12709 1615 12710 1649
rect 12674 1574 12710 1615
rect 12674 1540 12675 1574
rect 12709 1540 12710 1574
rect 12674 1499 12710 1540
rect 12674 1465 12675 1499
rect 12709 1465 12710 1499
rect 12674 1424 12710 1465
rect 12674 1390 12675 1424
rect 12709 1390 12710 1424
rect 12570 1375 12590 1390
rect 11860 1295 11894 1341
rect 11860 1215 11894 1261
rect 11860 1136 11894 1181
rect 11860 1057 11894 1102
rect 11860 978 11894 1023
rect 11860 899 11894 944
rect 11860 820 11894 865
rect 11860 741 11894 786
rect 12565 1295 12599 1341
rect 12565 1215 12599 1261
rect 12565 1136 12599 1181
rect 12565 1057 12599 1102
rect 12565 978 12599 1023
rect 12565 899 12599 944
rect 12565 820 12599 865
rect 12565 741 12599 786
rect 12674 1349 12710 1390
rect 12674 1315 12675 1349
rect 12709 1315 12710 1349
rect 12674 1274 12710 1315
rect 12674 1240 12675 1274
rect 12709 1240 12710 1274
rect 12674 1199 12710 1240
rect 12674 1165 12675 1199
rect 12709 1165 12710 1199
rect 12674 1124 12710 1165
rect 12674 1090 12675 1124
rect 12709 1090 12710 1124
rect 12674 1049 12710 1090
rect 12674 1015 12675 1049
rect 12709 1015 12710 1049
rect 12674 974 12710 1015
rect 12674 940 12675 974
rect 12709 940 12710 974
rect 12674 899 12710 940
rect 12674 865 12675 899
rect 12709 865 12710 899
rect 12674 825 12710 865
rect 12674 791 12675 825
rect 12709 791 12710 825
rect 12674 751 12710 791
rect 12674 717 12675 751
rect 12709 717 12710 751
rect 12570 668 12590 707
rect 12674 677 12710 717
rect 12674 643 12675 677
rect 12709 643 12710 677
rect 12674 608 12710 643
rect 9467 505 9468 544
rect 9502 505 9503 544
rect 9467 490 9503 505
rect 10296 558 10330 592
rect 10296 490 10330 524
rect 12674 569 12675 608
rect 12709 569 12710 608
rect 12674 490 12710 569
rect 9467 489 12710 490
rect 9467 471 9582 489
rect 9467 436 9468 471
rect 9502 455 9582 471
rect 9616 455 9650 489
rect 9684 455 9718 489
rect 9752 455 9786 489
rect 9820 455 9854 489
rect 9888 455 9922 489
rect 9956 455 9990 489
rect 10024 455 10058 489
rect 10092 455 10126 489
rect 10160 455 10194 489
rect 10228 455 10262 489
rect 10296 455 10330 489
rect 10364 455 10398 489
rect 10432 455 10466 489
rect 10500 455 10534 489
rect 10568 455 10602 489
rect 10636 455 10670 489
rect 10704 455 10738 489
rect 10772 455 10806 489
rect 10840 455 10874 489
rect 10908 455 10942 489
rect 10976 455 11010 489
rect 11044 455 11078 489
rect 11112 455 11146 489
rect 11180 455 11212 489
rect 11248 455 11282 489
rect 11321 455 11350 489
rect 11396 455 11418 489
rect 11471 455 11486 489
rect 11546 455 11554 489
rect 11621 455 11622 489
rect 11656 455 11662 489
rect 11724 455 11737 489
rect 11792 455 11812 489
rect 11860 455 11887 489
rect 11928 455 11962 489
rect 11996 455 12030 489
rect 12071 455 12098 489
rect 12146 455 12166 489
rect 12221 455 12234 489
rect 12296 455 12302 489
rect 12336 455 12337 489
rect 12404 455 12412 489
rect 12472 455 12487 489
rect 12540 455 12562 489
rect 12608 455 12637 489
rect 12676 455 12710 489
rect 9502 454 12710 455
rect 12945 5079 13682 5080
rect 12945 5046 13070 5079
rect 12945 5012 12946 5046
rect 12980 5045 13070 5046
rect 13104 5045 13138 5079
rect 13172 5045 13206 5079
rect 13240 5045 13274 5079
rect 13308 5045 13342 5079
rect 13376 5045 13410 5079
rect 13444 5045 13478 5079
rect 13512 5045 13546 5079
rect 13580 5045 13614 5079
rect 13648 5045 13682 5079
rect 12980 5044 13682 5045
rect 12980 5012 12981 5044
rect 12945 4978 12981 5012
rect 12945 4944 12946 4978
rect 12980 4944 12981 4978
rect 12945 4910 12981 4944
rect 12945 4876 12946 4910
rect 12980 4876 12981 4910
rect 12945 4842 12981 4876
rect 12945 4808 12946 4842
rect 12980 4808 12981 4842
rect 12945 4774 12981 4808
rect 12945 4740 12946 4774
rect 12980 4740 12981 4774
rect 12945 4706 12981 4740
rect 12945 4672 12946 4706
rect 12980 4672 12981 4706
rect 12945 4638 12981 4672
rect 12945 4604 12946 4638
rect 12980 4604 12981 4638
rect 12945 4570 12981 4604
rect 12945 4536 12946 4570
rect 12980 4536 12981 4570
rect 12945 4502 12981 4536
rect 12945 4468 12946 4502
rect 12980 4468 12981 4502
rect 12945 4434 12981 4468
rect 12945 4400 12946 4434
rect 12980 4400 12981 4434
rect 12945 4366 12981 4400
rect 12945 4332 12946 4366
rect 12980 4332 12981 4366
rect 12945 4298 12981 4332
rect 12945 4264 12946 4298
rect 12980 4264 12981 4298
rect 12945 4230 12981 4264
rect 12945 4196 12946 4230
rect 12980 4196 12981 4230
rect 12945 4162 12981 4196
rect 12945 4128 12946 4162
rect 12980 4128 12981 4162
rect 12945 4094 12981 4128
rect 12945 4060 12946 4094
rect 12980 4060 12981 4094
rect 12945 4026 12981 4060
rect 12945 3992 12946 4026
rect 12980 3992 12981 4026
rect 12945 3958 12981 3992
rect 12945 3924 12946 3958
rect 12980 3924 12981 3958
rect 12945 3890 12981 3924
rect 12945 3856 12946 3890
rect 12980 3856 12981 3890
rect 12945 3822 12981 3856
rect 12945 3788 12946 3822
rect 12980 3788 12981 3822
rect 12945 3754 12981 3788
rect 12945 3720 12946 3754
rect 12980 3720 12981 3754
rect 12945 3686 12981 3720
rect 12945 3652 12946 3686
rect 12980 3652 12981 3686
rect 12945 3618 12981 3652
rect 12945 3584 12946 3618
rect 12980 3584 12981 3618
rect 12945 3550 12981 3584
rect 12945 3516 12946 3550
rect 12980 3516 12981 3550
rect 12945 3482 12981 3516
rect 12945 3448 12946 3482
rect 12980 3448 12981 3482
rect 12945 3414 12981 3448
rect 12945 3380 12946 3414
rect 12980 3380 12981 3414
rect 12945 3346 12981 3380
rect 12945 3312 12946 3346
rect 12980 3312 12981 3346
rect 12945 3278 12981 3312
rect 12945 3244 12946 3278
rect 12980 3244 12981 3278
rect 12945 3210 12981 3244
rect 12945 3176 12946 3210
rect 12980 3176 12981 3210
rect 12945 3142 12981 3176
rect 12945 3108 12946 3142
rect 12980 3108 12981 3142
rect 12945 3074 12981 3108
rect 12945 3040 12946 3074
rect 12980 3040 12981 3074
rect 12945 3006 12981 3040
rect 12945 2972 12946 3006
rect 12980 2972 12981 3006
rect 12945 2938 12981 2972
rect 12945 2904 12946 2938
rect 12980 2904 12981 2938
rect 12945 2870 12981 2904
rect 12945 2836 12946 2870
rect 12980 2836 12981 2870
rect 12945 2802 12981 2836
rect 12945 2768 12946 2802
rect 12980 2768 12981 2802
rect 12945 2734 12981 2768
rect 12945 2700 12946 2734
rect 12980 2700 12981 2734
rect 12945 2666 12981 2700
rect 12945 2632 12946 2666
rect 12980 2632 12981 2666
rect 12945 2598 12981 2632
rect 12945 2564 12946 2598
rect 12980 2564 12981 2598
rect 12945 2530 12981 2564
rect 12945 2496 12946 2530
rect 12980 2496 12981 2530
rect 12945 2462 12981 2496
rect 12945 2428 12946 2462
rect 12980 2428 12981 2462
rect 12945 2394 12981 2428
rect 12945 2360 12946 2394
rect 12980 2360 12981 2394
rect 12945 2326 12981 2360
rect 12945 2292 12946 2326
rect 12980 2292 12981 2326
rect 12945 2258 12981 2292
rect 12945 2224 12946 2258
rect 12980 2224 12981 2258
rect 12945 2190 12981 2224
rect 12945 2156 12946 2190
rect 12980 2156 12981 2190
rect 12945 2122 12981 2156
rect 12945 2088 12946 2122
rect 12980 2088 12981 2122
rect 12945 2054 12981 2088
rect 12945 2020 12946 2054
rect 12980 2020 12981 2054
rect 12945 1986 12981 2020
rect 12945 1952 12946 1986
rect 12980 1952 12981 1986
rect 12945 1918 12981 1952
rect 12945 1884 12946 1918
rect 12980 1884 12981 1918
rect 12945 1850 12981 1884
rect 12945 1816 12946 1850
rect 12980 1816 12981 1850
rect 12945 1782 12981 1816
rect 12945 1748 12946 1782
rect 12980 1748 12981 1782
rect 12945 1714 12981 1748
rect 12945 1680 12946 1714
rect 12980 1680 12981 1714
rect 12945 1646 12981 1680
rect 12945 1612 12946 1646
rect 12980 1612 12981 1646
rect 12945 1578 12981 1612
rect 12945 1544 12946 1578
rect 12980 1544 12981 1578
rect 12945 1510 12981 1544
rect 12945 1476 12946 1510
rect 12980 1476 12981 1510
rect 12945 1442 12981 1476
rect 12945 1408 12946 1442
rect 12980 1408 12981 1442
rect 12945 1374 12981 1408
rect 12945 1340 12946 1374
rect 12980 1340 12981 1374
rect 12945 1306 12981 1340
rect 12945 1272 12946 1306
rect 12980 1272 12981 1306
rect 12945 1238 12981 1272
rect 12945 1204 12946 1238
rect 12980 1204 12981 1238
rect 12945 1170 12981 1204
rect 12945 1136 12946 1170
rect 12980 1136 12981 1170
rect 12945 1102 12981 1136
rect 12945 1068 12946 1102
rect 12980 1068 12981 1102
rect 12945 1034 12981 1068
rect 12945 1000 12946 1034
rect 12980 1000 12981 1034
rect 12945 966 12981 1000
rect 12945 932 12946 966
rect 12980 932 12981 966
rect 12945 898 12981 932
rect 12945 864 12946 898
rect 12980 864 12981 898
rect 12945 830 12981 864
rect 12945 796 12946 830
rect 12980 796 12981 830
rect 12945 762 12981 796
rect 12945 728 12946 762
rect 12980 728 12981 762
rect 12945 694 12981 728
rect 12945 660 12946 694
rect 12980 660 12981 694
rect 12945 626 12981 660
rect 12945 592 12946 626
rect 12980 592 12981 626
rect 12945 558 12981 592
rect 12945 524 12946 558
rect 12980 524 12981 558
rect 12945 490 12981 524
rect 12945 456 12946 490
rect 12980 456 12981 490
rect 9502 436 9503 454
rect 9467 401 9503 436
rect 9467 364 9468 401
rect 9502 364 9503 401
rect 9467 332 9503 364
rect 9467 291 9468 332
rect 9502 291 9503 332
rect 12945 422 12981 456
rect 12945 388 12946 422
rect 12980 388 12981 422
rect 12945 354 12981 388
rect 9467 245 9503 291
rect 4834 211 4844 243
rect 4878 211 4917 245
rect 4951 244 4990 245
rect 5024 244 5063 245
rect 5097 244 5136 245
rect 5170 244 5209 245
rect 5243 244 5282 245
rect 5316 244 5355 245
rect 5389 244 5428 245
rect 5462 244 5501 245
rect 5535 244 5574 245
rect 5608 244 5646 245
rect 5680 244 5718 245
rect 5752 244 5790 245
rect 5824 244 5862 245
rect 5896 244 5934 245
rect 5968 244 6006 245
rect 6040 244 6078 245
rect 6112 244 6150 245
rect 6184 244 6222 245
rect 6256 244 6294 245
rect 6328 244 6366 245
rect 6400 244 6438 245
rect 6472 244 6510 245
rect 6544 244 6582 245
rect 6616 244 6654 245
rect 6688 244 6726 245
rect 6760 244 6798 245
rect 6832 244 6870 245
rect 6904 244 6942 245
rect 6976 244 7014 245
rect 7048 244 7086 245
rect 7120 244 7158 245
rect 7192 244 7230 245
rect 7264 244 7302 245
rect 7336 244 7374 245
rect 7408 244 7446 245
rect 7480 244 7518 245
rect 7552 244 7590 245
rect 7624 244 7662 245
rect 7696 244 7734 245
rect 7768 244 7806 245
rect 7840 244 7878 245
rect 7912 244 7950 245
rect 7984 244 8022 245
rect 8056 244 8094 245
rect 8128 244 8166 245
rect 8200 244 8238 245
rect 8272 244 8310 245
rect 8344 244 8382 245
rect 8416 244 8454 245
rect 8488 244 8526 245
rect 8560 244 8598 245
rect 8632 244 8670 245
rect 8704 244 8742 245
rect 8776 244 8814 245
rect 8848 244 8886 245
rect 8920 244 8958 245
rect 8992 244 9030 245
rect 9064 244 9102 245
rect 9136 244 9174 245
rect 9208 244 9246 245
rect 9280 244 9318 245
rect 9352 244 9390 245
rect 9424 244 9462 245
rect 4981 211 4990 244
rect 5049 211 5063 244
rect 5117 211 5136 244
rect 5185 211 5209 244
rect 5253 211 5282 244
rect 4834 210 4947 211
rect 4981 210 5015 211
rect 5049 210 5083 211
rect 5117 210 5151 211
rect 5185 210 5219 211
rect 5253 210 5287 211
rect 5321 210 5355 244
rect 5389 210 5423 244
rect 5462 211 5491 244
rect 5535 211 5559 244
rect 5608 211 5627 244
rect 5680 211 5695 244
rect 5752 211 5763 244
rect 5824 211 5831 244
rect 5896 211 5899 244
rect 5457 210 5491 211
rect 5525 210 5559 211
rect 5593 210 5627 211
rect 5661 210 5695 211
rect 5729 210 5763 211
rect 5797 210 5831 211
rect 5865 210 5899 211
rect 5933 211 5934 244
rect 6001 211 6006 244
rect 6069 211 6078 244
rect 6137 211 6150 244
rect 6205 211 6222 244
rect 6273 211 6294 244
rect 6341 211 6366 244
rect 6409 211 6438 244
rect 6477 211 6510 244
rect 5933 210 5967 211
rect 6001 210 6035 211
rect 6069 210 6103 211
rect 6137 210 6171 211
rect 6205 210 6239 211
rect 6273 210 6307 211
rect 6341 210 6375 211
rect 6409 210 6443 211
rect 6477 210 6511 211
rect 6545 210 6579 244
rect 6616 211 6647 244
rect 6688 211 6715 244
rect 6760 211 6783 244
rect 6832 211 6851 244
rect 6904 211 6919 244
rect 6976 211 6987 244
rect 7048 211 7055 244
rect 7120 211 7123 244
rect 6613 210 6647 211
rect 6681 210 6715 211
rect 6749 210 6783 211
rect 6817 210 6851 211
rect 6885 210 6919 211
rect 6953 210 6987 211
rect 7021 210 7055 211
rect 7089 210 7123 211
rect 7157 211 7158 244
rect 7225 211 7230 244
rect 7293 211 7302 244
rect 7361 211 7374 244
rect 7429 211 7446 244
rect 7497 211 7518 244
rect 7565 211 7590 244
rect 7633 211 7662 244
rect 7701 211 7734 244
rect 7157 210 7191 211
rect 7225 210 7259 211
rect 7293 210 7327 211
rect 7361 210 7395 211
rect 7429 210 7463 211
rect 7497 210 7531 211
rect 7565 210 7599 211
rect 7633 210 7667 211
rect 7701 210 7735 211
rect 7769 210 7803 244
rect 7840 211 7871 244
rect 7912 211 7939 244
rect 7984 211 8007 244
rect 8056 211 8075 244
rect 8128 211 8143 244
rect 8200 211 8211 244
rect 8272 211 8279 244
rect 8344 211 8347 244
rect 7837 210 7871 211
rect 7905 210 7939 211
rect 7973 210 8007 211
rect 8041 210 8075 211
rect 8109 210 8143 211
rect 8177 210 8211 211
rect 8245 210 8279 211
rect 8313 210 8347 211
rect 8381 211 8382 244
rect 8449 211 8454 244
rect 8517 211 8526 244
rect 8585 211 8598 244
rect 8653 211 8670 244
rect 8721 211 8742 244
rect 8789 211 8814 244
rect 8857 211 8886 244
rect 8925 211 8958 244
rect 8381 210 8415 211
rect 8449 210 8483 211
rect 8517 210 8551 211
rect 8585 210 8619 211
rect 8653 210 8687 211
rect 8721 210 8755 211
rect 8789 210 8823 211
rect 8857 210 8891 211
rect 8925 210 8959 211
rect 8993 210 9027 244
rect 9064 211 9095 244
rect 9136 211 9163 244
rect 9208 211 9231 244
rect 9280 211 9299 244
rect 9352 211 9367 244
rect 9424 211 9435 244
rect 9496 211 9503 245
rect 9061 210 9095 211
rect 9129 210 9163 211
rect 9197 210 9231 211
rect 9265 210 9299 211
rect 9333 210 9367 211
rect 9401 210 9435 211
rect 9469 210 9503 211
rect 4834 209 9503 210
rect 9650 310 9759 326
rect 9650 281 9657 310
rect 9725 281 9759 310
rect 9756 276 9759 281
rect 4645 169 4681 203
rect 9650 208 9657 247
rect 9725 208 9759 242
rect 9650 192 9759 208
rect 10065 310 10196 326
rect 10065 281 10099 310
rect 10167 281 10196 310
rect 10065 276 10090 281
rect 10065 208 10099 242
rect 10167 208 10196 247
rect 10065 192 10196 208
rect 10436 310 10573 326
rect 10504 281 10573 310
rect 10504 276 10539 281
rect 10538 247 10539 276
rect 10538 242 10573 247
rect 10504 208 10573 242
rect 10436 192 10573 208
rect 10844 310 10999 326
rect 10844 276 10878 310
rect 10946 281 10999 310
rect 10946 247 10965 281
rect 10844 208 10878 242
rect 10946 208 10999 247
rect 10844 192 10999 208
rect 11195 314 11334 326
rect 11195 310 11300 314
rect 11263 280 11300 310
rect 11263 276 11334 280
rect 11297 242 11334 276
rect 11263 208 11300 242
rect 11195 192 11334 208
rect 11603 310 12264 326
rect 11603 276 11637 310
rect 11705 267 12162 310
rect 12230 276 12264 310
rect 11603 208 11637 242
rect 11705 233 11846 267
rect 11880 233 11925 267
rect 11959 233 12004 267
rect 12038 233 12082 267
rect 12116 233 12162 267
rect 11705 208 12162 233
rect 12230 208 12264 242
rect 11603 192 12264 208
rect 12570 314 12672 326
rect 12570 280 12574 314
rect 12608 310 12672 314
rect 12570 276 12604 280
rect 12570 208 12574 242
rect 12570 192 12672 208
rect 12945 320 12946 354
rect 12980 320 12981 354
rect 12945 286 12981 320
rect 12945 252 12946 286
rect 12980 252 12981 286
rect 12945 218 12981 252
rect 4645 135 4646 169
rect 4680 135 4681 169
rect 4645 101 4681 135
rect 4645 67 4646 101
rect 4680 67 4681 101
rect 4645 33 4681 67
rect 4645 -1 4646 33
rect 4680 -1 4681 33
rect 12945 184 12946 218
rect 12980 184 12981 218
rect 12945 150 12981 184
rect 12945 116 12946 150
rect 12980 116 12981 150
rect 12945 82 12981 116
rect 12945 48 12946 82
rect 12980 48 12981 82
rect 12945 14 12981 48
rect 4645 -35 4681 -1
rect 4645 -69 4646 -35
rect 4680 -69 4681 -35
rect 4645 -103 4681 -69
rect 4645 -137 4646 -103
rect 4680 -137 4681 -103
rect 4645 -171 4681 -137
rect 4645 -205 4646 -171
rect 4680 -205 4681 -171
rect 4645 -239 4681 -205
rect 6465 -28 6627 4
rect 6465 -130 6524 -28
rect 6626 -130 6627 -28
rect 6465 -172 6627 -130
rect 8341 -28 8379 -8
rect 10791 -28 10893 -12
rect 12574 -28 12676 -12
rect 8307 -146 8409 -130
rect 10791 -146 10893 -130
rect 12608 -134 12676 -130
rect 12574 -146 12676 -134
rect 12945 -20 12946 14
rect 12980 -20 12981 14
rect 12945 -54 12981 -20
rect 12945 -88 12946 -54
rect 12980 -88 12981 -54
rect 6465 -206 6508 -172
rect 6542 -206 6580 -172
rect 6614 -206 6627 -172
rect 6465 -216 6627 -206
rect 4645 -273 4646 -239
rect 4680 -273 4681 -239
rect 4645 -307 4681 -273
rect 4645 -341 4646 -307
rect 4680 -341 4681 -307
rect 4645 -375 4681 -341
rect 4645 -409 4646 -375
rect 4680 -407 4681 -375
rect 12945 -223 12981 -88
rect 12945 -257 12946 -223
rect 12980 -257 12981 -223
rect 12945 -291 12981 -257
rect 12945 -325 12946 -291
rect 12980 -325 12981 -291
rect 12945 -407 12981 -325
rect 4680 -408 12981 -407
rect 4680 -409 4753 -408
rect 4645 -442 4753 -409
rect 4787 -442 4821 -408
rect 4855 -442 4889 -408
rect 4923 -442 4957 -408
rect 4991 -442 5025 -408
rect 5059 -442 5093 -408
rect 5127 -442 5161 -408
rect 5195 -442 5229 -408
rect 5263 -442 5297 -408
rect 5331 -442 5365 -408
rect 5399 -442 5433 -408
rect 5467 -442 5501 -408
rect 5535 -442 5569 -408
rect 5603 -442 5637 -408
rect 5671 -442 5705 -408
rect 5739 -442 5773 -408
rect 5807 -442 5841 -408
rect 5875 -442 5909 -408
rect 5943 -442 5977 -408
rect 6011 -442 6045 -408
rect 6079 -442 6113 -408
rect 6147 -442 6181 -408
rect 6215 -442 6249 -408
rect 6283 -442 6317 -408
rect 6351 -442 6385 -408
rect 6419 -442 6453 -408
rect 6487 -442 6521 -408
rect 6555 -442 6589 -408
rect 6623 -442 6657 -408
rect 6691 -442 6725 -408
rect 6759 -442 6793 -408
rect 6827 -442 6861 -408
rect 6895 -442 6929 -408
rect 6963 -442 6997 -408
rect 7031 -442 7065 -408
rect 7099 -442 7133 -408
rect 7167 -442 7201 -408
rect 7235 -442 7269 -408
rect 7303 -442 7337 -408
rect 7371 -442 7405 -408
rect 7439 -442 7473 -408
rect 7507 -442 7541 -408
rect 7575 -442 7609 -408
rect 7643 -442 7677 -408
rect 7711 -442 7745 -408
rect 7779 -442 7813 -408
rect 7847 -442 7881 -408
rect 7915 -442 7949 -408
rect 7983 -442 8017 -408
rect 8051 -442 8085 -408
rect 8119 -442 8153 -408
rect 8187 -442 8221 -408
rect 8255 -442 8289 -408
rect 8323 -442 8357 -408
rect 8391 -442 8425 -408
rect 8459 -442 8493 -408
rect 8527 -442 8561 -408
rect 8595 -442 8629 -408
rect 8663 -442 8697 -408
rect 8731 -442 8765 -408
rect 8799 -442 8833 -408
rect 8867 -442 8901 -408
rect 8935 -442 8969 -408
rect 9003 -442 9037 -408
rect 9071 -442 9105 -408
rect 9139 -442 9173 -408
rect 9207 -442 9241 -408
rect 9275 -442 9309 -408
rect 9343 -442 9377 -408
rect 9411 -442 9445 -408
rect 9479 -442 9513 -408
rect 9547 -442 9581 -408
rect 9615 -442 9649 -408
rect 9683 -442 9717 -408
rect 9751 -442 9785 -408
rect 9819 -442 9853 -408
rect 9887 -442 9921 -408
rect 9955 -442 9989 -408
rect 10023 -442 10057 -408
rect 10091 -442 10125 -408
rect 10159 -442 10193 -408
rect 10227 -442 10261 -408
rect 10295 -442 10329 -408
rect 10363 -442 10397 -408
rect 10431 -442 10465 -408
rect 10499 -442 10533 -408
rect 10567 -442 10601 -408
rect 10635 -442 10669 -408
rect 10703 -442 10737 -408
rect 10771 -442 10805 -408
rect 10839 -442 10873 -408
rect 10907 -442 10941 -408
rect 10975 -442 11009 -408
rect 11043 -442 11077 -408
rect 11111 -442 11145 -408
rect 11179 -442 11213 -408
rect 11247 -442 11281 -408
rect 11315 -442 11349 -408
rect 11383 -442 11417 -408
rect 11451 -442 11485 -408
rect 11519 -442 11553 -408
rect 11587 -442 11621 -408
rect 11655 -442 11689 -408
rect 11723 -442 11757 -408
rect 11791 -442 11825 -408
rect 11859 -442 11893 -408
rect 11927 -442 11961 -408
rect 11995 -442 12029 -408
rect 12063 -442 12097 -408
rect 12131 -442 12165 -408
rect 12199 -442 12233 -408
rect 12267 -442 12301 -408
rect 12335 -442 12369 -408
rect 12403 -442 12437 -408
rect 12471 -442 12505 -408
rect 12539 -442 12573 -408
rect 12607 -442 12641 -408
rect 12675 -442 12709 -408
rect 12743 -442 12777 -408
rect 12811 -442 12845 -408
rect 12879 -442 12913 -408
rect 12947 -442 12981 -408
rect 4645 -443 12981 -442
<< viali >>
rect 6161 13027 6195 13061
rect 6281 13033 6315 13067
rect 6353 13033 6387 13067
rect 6425 13033 6459 13067
rect 6497 13033 6531 13067
rect 6569 13033 6603 13067
rect 6641 13033 6675 13067
rect 6713 13033 6747 13067
rect 6785 13033 6819 13067
rect 6857 13033 6891 13067
rect 6929 13033 6963 13067
rect 7001 13033 7035 13067
rect 7073 13033 7107 13067
rect 7145 13033 7179 13067
rect 7217 13033 7251 13067
rect 7289 13033 7323 13067
rect 7361 13033 7395 13067
rect 7433 13033 7467 13067
rect 7505 13033 7539 13067
rect 7577 13033 7611 13067
rect 7649 13033 7683 13067
rect 7721 13033 7755 13067
rect 7793 13033 7827 13067
rect 7865 13033 7899 13067
rect 7937 13033 7971 13067
rect 8009 13033 8043 13067
rect 8081 13033 8115 13067
rect 8153 13033 8187 13067
rect 8225 13033 8259 13067
rect 8297 13033 8331 13067
rect 8369 13033 8403 13067
rect 8441 13033 8475 13067
rect 8513 13033 8547 13067
rect 8585 13033 8619 13067
rect 8657 13033 8691 13067
rect 8729 13033 8763 13067
rect 8801 13033 8835 13067
rect 8873 13033 8907 13067
rect 8945 13033 8979 13067
rect 9017 13033 9051 13067
rect 9089 13033 9123 13067
rect 9161 13033 9195 13067
rect 9233 13033 9267 13067
rect 9305 13033 9339 13067
rect 9377 13033 9411 13067
rect 9449 13033 9483 13067
rect 9521 13033 9555 13067
rect 9593 13033 9627 13067
rect 9665 13033 9699 13067
rect 9737 13033 9771 13067
rect 9809 13033 9843 13067
rect 9881 13033 9915 13067
rect 9953 13033 9987 13067
rect 6161 12955 6195 12989
rect 6161 12883 6195 12917
rect 6161 12811 6195 12845
rect 6161 12739 6195 12773
rect 6161 12667 6195 12701
rect 6161 12595 6195 12629
rect 6161 12523 6195 12557
rect 6161 12451 6195 12485
rect 6161 12379 6195 12413
rect 6161 12307 6195 12341
rect 6161 12235 6195 12269
rect 6161 12163 6195 12197
rect 6161 12091 6195 12125
rect 6161 12019 6195 12053
rect 6161 11947 6195 11981
rect 6161 11875 6195 11909
rect 6161 11803 6195 11837
rect 6161 11731 6195 11765
rect 6161 11659 6195 11693
rect 6161 11587 6195 11621
rect 6161 11515 6195 11549
rect 6161 11443 6195 11477
rect 6161 11371 6195 11405
rect 6161 11299 6195 11333
rect 10232 11294 10255 11319
rect 10255 11294 10266 11319
rect 10308 11294 10325 11319
rect 10325 11294 10342 11319
rect 10384 11294 10395 11319
rect 10395 11294 10418 11319
rect 10460 11294 10465 11319
rect 10465 11294 10494 11319
rect 10536 11294 10569 11319
rect 10569 11294 10570 11319
rect 10612 11294 10638 11319
rect 10638 11294 10646 11319
rect 10688 11294 10707 11319
rect 10707 11294 10722 11319
rect 10764 11294 10776 11319
rect 10776 11294 10798 11319
rect 10840 11294 10845 11319
rect 10845 11294 10874 11319
rect 10915 11294 10948 11319
rect 10948 11294 10949 11319
rect 10990 11294 11017 11319
rect 11017 11294 11024 11319
rect 11065 11294 11086 11319
rect 11086 11294 11099 11319
rect 11140 11294 11155 11319
rect 11155 11294 11174 11319
rect 11215 11294 11224 11319
rect 11224 11294 11249 11319
rect 11290 11294 11293 11319
rect 11293 11294 11324 11319
rect 11365 11294 11397 11319
rect 11397 11294 11399 11319
rect 11440 11294 11466 11319
rect 11466 11294 11474 11319
rect 11515 11294 11535 11319
rect 11535 11294 11549 11319
rect 11590 11294 11604 11319
rect 11604 11294 11624 11319
rect 11665 11294 11673 11319
rect 11673 11294 11699 11319
rect 11740 11294 11742 11319
rect 11742 11294 11774 11319
rect 11815 11294 11845 11319
rect 11845 11294 11849 11319
rect 10232 11285 10266 11294
rect 10308 11285 10342 11294
rect 10384 11285 10418 11294
rect 10460 11285 10494 11294
rect 10536 11285 10570 11294
rect 10612 11285 10646 11294
rect 10688 11285 10722 11294
rect 10764 11285 10798 11294
rect 10840 11285 10874 11294
rect 10915 11285 10949 11294
rect 10990 11285 11024 11294
rect 11065 11285 11099 11294
rect 11140 11285 11174 11294
rect 11215 11285 11249 11294
rect 11290 11285 11324 11294
rect 11365 11285 11399 11294
rect 11440 11285 11474 11294
rect 11515 11285 11549 11294
rect 11590 11285 11624 11294
rect 11665 11285 11699 11294
rect 11740 11285 11774 11294
rect 11815 11285 11849 11294
rect 6167 11165 6201 11199
rect 6239 11165 6273 11199
rect 6311 11165 6345 11199
rect 6383 11165 6417 11199
rect 6455 11165 6489 11199
rect 6527 11165 6561 11199
rect 6599 11165 6633 11199
rect 6671 11165 6705 11199
rect 6743 11165 6777 11199
rect 6815 11165 6849 11199
rect 6887 11165 6921 11199
rect 6959 11165 6993 11199
rect 7031 11165 7065 11199
rect 7103 11165 7137 11199
rect 7175 11165 7209 11199
rect 7247 11165 7281 11199
rect 7319 11165 7353 11199
rect 7391 11165 7425 11199
rect 7463 11165 7497 11199
rect 7535 11165 7569 11199
rect 7607 11165 7641 11199
rect 7679 11165 7713 11199
rect 7751 11165 7785 11199
rect 7823 11165 7857 11199
rect 7895 11165 7929 11199
rect 7967 11165 8001 11199
rect 8039 11165 8073 11199
rect 8111 11165 8145 11199
rect 8183 11165 8217 11199
rect 8255 11165 8289 11199
rect 2155 11036 2189 11070
rect 2496 11069 2530 11103
rect 2589 11069 2623 11103
rect 332 10632 366 10666
rect 332 10560 366 10594
rect 7070 10980 7104 11014
rect 7149 10980 7183 11014
rect 7228 10980 7262 11014
rect 7306 10980 7340 11014
rect 7384 10980 7418 11014
rect 7462 10980 7496 11014
rect 7070 10902 7104 10936
rect 7149 10902 7183 10936
rect 7228 10902 7262 10936
rect 7306 10902 7340 10936
rect 7384 10902 7418 10936
rect 7462 10902 7496 10936
rect 6499 10403 6504 10437
rect 6504 10403 6533 10437
rect 6572 10403 6573 10437
rect 6573 10403 6606 10437
rect 6645 10403 6676 10437
rect 6676 10403 6679 10437
rect 6718 10403 6745 10437
rect 6745 10403 6752 10437
rect 6791 10403 6814 10437
rect 6814 10403 6825 10437
rect 6864 10403 6883 10437
rect 6883 10403 6898 10437
rect 6937 10403 6952 10437
rect 6952 10403 6971 10437
rect 7010 10403 7021 10437
rect 7021 10403 7044 10437
rect 7083 10403 7090 10437
rect 7090 10403 7117 10437
rect 7156 10403 7159 10437
rect 7159 10403 7190 10437
rect 7229 10403 7263 10437
rect 7302 10403 7332 10437
rect 7332 10403 7336 10437
rect 7375 10403 7401 10437
rect 7401 10403 7409 10437
rect 7448 10403 7470 10437
rect 7470 10403 7482 10437
rect 7521 10403 7539 10437
rect 7539 10403 7555 10437
rect 7594 10403 7608 10437
rect 7608 10403 7628 10437
rect 7667 10403 7677 10437
rect 7677 10403 7701 10437
rect 7740 10403 7746 10437
rect 7746 10403 7774 10437
rect 7813 10403 7815 10437
rect 7815 10403 7847 10437
rect 7886 10403 7918 10437
rect 7918 10403 7920 10437
rect 7959 10403 7987 10437
rect 7987 10403 7993 10437
rect 8032 10403 8056 10437
rect 8056 10403 8066 10437
rect 8105 10403 8125 10437
rect 8125 10403 8139 10437
rect 8178 10403 8194 10437
rect 8194 10403 8212 10437
rect 8251 10403 8263 10437
rect 8263 10403 8285 10437
rect 8324 10403 8332 10437
rect 8332 10403 8358 10437
rect 8397 10403 8401 10437
rect 8401 10403 8431 10437
rect 8470 10403 8504 10437
rect 8543 10403 8574 10437
rect 8574 10403 8577 10437
rect 8616 10403 8643 10437
rect 8643 10403 8650 10437
rect 8689 10403 8712 10437
rect 8712 10403 8723 10437
rect 8762 10403 8781 10437
rect 8781 10403 8796 10437
rect 8835 10403 8850 10437
rect 8850 10403 8869 10437
rect 8908 10403 8919 10437
rect 8919 10403 8942 10437
rect 8981 10403 8988 10437
rect 8988 10403 9015 10437
rect 9054 10403 9057 10437
rect 9057 10403 9088 10437
rect 9127 10403 9160 10437
rect 9160 10403 9161 10437
rect 9200 10403 9229 10437
rect 9229 10403 9234 10437
rect 9273 10403 9298 10437
rect 9298 10403 9307 10437
rect 9346 10403 9367 10437
rect 9367 10403 9380 10437
rect 9419 10403 9436 10437
rect 9436 10403 9453 10437
rect 9492 10403 9505 10437
rect 9505 10403 9526 10437
rect 9565 10403 9574 10437
rect 9574 10403 9599 10437
rect 9638 10403 9643 10437
rect 9643 10403 9672 10437
rect 9711 10403 9712 10437
rect 9712 10403 9745 10437
rect 9784 10403 9816 10437
rect 9816 10403 9818 10437
rect 9857 10403 9885 10437
rect 9885 10403 9891 10437
rect 9930 10403 9954 10437
rect 9954 10403 9964 10437
rect 10003 10403 10022 10437
rect 10022 10403 10037 10437
rect 10076 10403 10090 10437
rect 10090 10403 10110 10437
rect 10149 10403 10158 10437
rect 10158 10403 10183 10437
rect 10222 10403 10226 10437
rect 10226 10403 10256 10437
rect 10294 10403 10328 10437
rect 10366 10403 10396 10437
rect 10396 10403 10400 10437
rect 10438 10403 10464 10437
rect 10464 10403 10472 10437
rect 10510 10403 10532 10437
rect 10532 10403 10544 10437
rect 10582 10403 10600 10437
rect 10600 10403 10616 10437
rect 10654 10403 10668 10437
rect 10668 10403 10688 10437
rect 10726 10403 10736 10437
rect 10736 10403 10760 10437
rect 10798 10403 10804 10437
rect 10804 10403 10832 10437
rect 10870 10403 10872 10437
rect 10872 10403 10904 10437
rect 10942 10403 10974 10437
rect 10974 10403 10976 10437
rect 11014 10403 11042 10437
rect 11042 10403 11048 10437
rect 11086 10403 11110 10437
rect 11110 10403 11120 10437
rect 11158 10403 11178 10437
rect 11178 10403 11192 10437
rect 11230 10403 11246 10437
rect 11246 10403 11264 10437
rect 11302 10403 11314 10437
rect 11314 10403 11336 10437
rect 11374 10403 11382 10437
rect 11382 10403 11408 10437
rect 11446 10403 11450 10437
rect 11450 10403 11480 10437
rect 11518 10403 11552 10437
rect 7069 10098 7103 10132
rect 7147 10098 7181 10132
rect 7225 10098 7259 10132
rect 7372 10098 7406 10132
rect 7444 10098 7478 10132
rect 7069 10017 7103 10051
rect 7147 10017 7181 10051
rect 7225 10017 7259 10051
rect 7372 10017 7406 10051
rect 7444 10017 7478 10051
rect 7069 9936 7103 9970
rect 7147 9936 7181 9970
rect 7225 9936 7259 9970
rect 7372 9936 7406 9970
rect 7444 9936 7478 9970
rect 7069 9855 7103 9889
rect 7147 9855 7181 9889
rect 7225 9855 7259 9889
rect 7372 9855 7406 9889
rect 7444 9855 7478 9889
rect 7069 9773 7103 9807
rect 7147 9773 7181 9807
rect 7225 9773 7259 9807
rect 7372 9773 7406 9807
rect 7444 9773 7478 9807
rect 7069 9691 7103 9725
rect 7147 9691 7181 9725
rect 7225 9691 7259 9725
rect 7372 9691 7406 9725
rect 7444 9691 7478 9725
rect 7069 9609 7103 9643
rect 7147 9609 7181 9643
rect 7225 9609 7259 9643
rect 7372 9609 7406 9643
rect 7444 9609 7478 9643
rect 6499 9519 6504 9547
rect 6504 9519 6533 9547
rect 6573 9519 6607 9547
rect 6647 9519 6676 9547
rect 6676 9519 6681 9547
rect 6721 9519 6745 9547
rect 6745 9519 6755 9547
rect 6795 9519 6814 9547
rect 6814 9519 6829 9547
rect 6869 9519 6883 9547
rect 6883 9519 6903 9547
rect 6943 9519 6952 9547
rect 6952 9519 6977 9547
rect 7017 9519 7021 9547
rect 7021 9519 7051 9547
rect 6499 9513 6533 9519
rect 6573 9513 6607 9519
rect 6647 9513 6681 9519
rect 6721 9513 6755 9519
rect 6795 9513 6829 9519
rect 6869 9513 6903 9519
rect 6943 9513 6977 9519
rect 7017 9513 7051 9519
rect 7091 9513 7125 9547
rect 7165 9519 7194 9547
rect 7194 9519 7199 9547
rect 7239 9519 7263 9547
rect 7263 9519 7273 9547
rect 7313 9519 7332 9547
rect 7332 9519 7347 9547
rect 7387 9519 7401 9547
rect 7401 9519 7421 9547
rect 7461 9519 7470 9547
rect 7470 9519 7495 9547
rect 7535 9519 7539 9547
rect 7539 9519 7569 9547
rect 7609 9519 7642 9547
rect 7642 9519 7643 9547
rect 7683 9519 7711 9547
rect 7711 9519 7717 9547
rect 7757 9519 7780 9547
rect 7780 9519 7791 9547
rect 7831 9519 7849 9547
rect 7849 9519 7865 9547
rect 7905 9519 7918 9547
rect 7918 9519 7939 9547
rect 7979 9519 7987 9547
rect 7987 9519 8013 9547
rect 8053 9519 8056 9547
rect 8056 9519 8087 9547
rect 8127 9519 8160 9547
rect 8160 9519 8161 9547
rect 8201 9519 8229 9547
rect 8229 9519 8235 9547
rect 8275 9519 8298 9547
rect 8298 9519 8309 9547
rect 8349 9519 8367 9547
rect 8367 9519 8383 9547
rect 8423 9519 8436 9547
rect 8436 9519 8457 9547
rect 8496 9519 8505 9547
rect 8505 9519 8530 9547
rect 8569 9519 8574 9547
rect 8574 9519 8603 9547
rect 8642 9519 8643 9547
rect 8643 9519 8676 9547
rect 8715 9519 8746 9547
rect 8746 9519 8749 9547
rect 8788 9519 8815 9547
rect 8815 9519 8822 9547
rect 8861 9519 8884 9547
rect 8884 9519 8895 9547
rect 8934 9519 8952 9547
rect 8952 9519 8968 9547
rect 9007 9519 9020 9547
rect 9020 9519 9041 9547
rect 9080 9519 9088 9547
rect 9088 9519 9114 9547
rect 9153 9519 9156 9547
rect 9156 9519 9187 9547
rect 9226 9519 9258 9547
rect 9258 9519 9260 9547
rect 9299 9519 9326 9547
rect 9326 9519 9333 9547
rect 9372 9519 9394 9547
rect 9394 9519 9406 9547
rect 9445 9519 9462 9547
rect 9462 9519 9479 9547
rect 9518 9519 9530 9547
rect 9530 9519 9552 9547
rect 9591 9519 9598 9547
rect 9598 9519 9625 9547
rect 9664 9519 9666 9547
rect 9666 9519 9698 9547
rect 9737 9519 9768 9547
rect 9768 9519 9771 9547
rect 9810 9519 9836 9547
rect 9836 9519 9844 9547
rect 7165 9513 7199 9519
rect 7239 9513 7273 9519
rect 7313 9513 7347 9519
rect 7387 9513 7421 9519
rect 7461 9513 7495 9519
rect 7535 9513 7569 9519
rect 7609 9513 7643 9519
rect 7683 9513 7717 9519
rect 7757 9513 7791 9519
rect 7831 9513 7865 9519
rect 7905 9513 7939 9519
rect 7979 9513 8013 9519
rect 8053 9513 8087 9519
rect 8127 9513 8161 9519
rect 8201 9513 8235 9519
rect 8275 9513 8309 9519
rect 8349 9513 8383 9519
rect 8423 9513 8457 9519
rect 8496 9513 8530 9519
rect 8569 9513 8603 9519
rect 8642 9513 8676 9519
rect 8715 9513 8749 9519
rect 8788 9513 8822 9519
rect 8861 9513 8895 9519
rect 8934 9513 8968 9519
rect 9007 9513 9041 9519
rect 9080 9513 9114 9519
rect 9153 9513 9187 9519
rect 9226 9513 9260 9519
rect 9299 9513 9333 9519
rect 9372 9513 9406 9519
rect 9445 9513 9479 9519
rect 9518 9513 9552 9519
rect 9591 9513 9625 9519
rect 9664 9513 9698 9519
rect 9737 9513 9771 9519
rect 9810 9513 9844 9519
rect 7069 9368 7103 9402
rect 7147 9368 7181 9402
rect 7225 9368 7259 9402
rect 7372 9368 7406 9402
rect 7444 9368 7478 9402
rect 7069 9287 7103 9321
rect 7147 9287 7181 9321
rect 7225 9287 7259 9321
rect 7372 9287 7406 9321
rect 7444 9287 7478 9321
rect 7069 9206 7103 9240
rect 7147 9206 7181 9240
rect 7225 9206 7259 9240
rect 7372 9206 7406 9240
rect 7444 9206 7478 9240
rect 7069 9125 7103 9159
rect 7147 9125 7181 9159
rect 7225 9125 7259 9159
rect 7372 9125 7406 9159
rect 7444 9125 7478 9159
rect 7069 9043 7103 9077
rect 7147 9043 7181 9077
rect 7225 9043 7259 9077
rect 7372 9043 7406 9077
rect 7444 9043 7478 9077
rect 7069 8961 7103 8995
rect 7147 8961 7181 8995
rect 7225 8961 7259 8995
rect 7372 8961 7406 8995
rect 7444 8961 7478 8995
rect 7069 8879 7103 8913
rect 7147 8879 7181 8913
rect 7225 8879 7259 8913
rect 7372 8879 7406 8913
rect 7444 8879 7478 8913
rect 250 6139 284 6147
rect 250 6113 284 6139
rect 778 6119 812 6147
rect 778 6113 812 6119
rect 250 6037 284 6041
rect 250 6007 284 6037
rect 250 5935 284 5969
rect 250 5867 284 5887
rect 250 5853 284 5867
rect 250 5799 284 5804
rect 250 5770 284 5799
rect 250 5697 284 5721
rect 250 5687 284 5697
rect 250 5629 284 5638
rect 250 5604 284 5629
rect 250 5527 284 5555
rect 250 5521 284 5527
rect 250 5459 284 5472
rect 250 5438 284 5459
rect 693 5859 727 5881
rect 693 5847 727 5859
rect 693 5786 727 5809
rect 693 5775 727 5786
rect 693 5713 727 5737
rect 693 5703 727 5713
rect 693 5640 727 5665
rect 693 5631 727 5640
rect 693 5567 727 5593
rect 693 5559 727 5567
rect 693 5494 727 5521
rect 693 5487 727 5494
rect 778 6051 812 6061
rect 778 6027 812 6051
rect 778 5847 812 5881
rect 778 5779 812 5786
rect 778 5752 812 5779
rect 778 5677 812 5691
rect 778 5657 812 5677
rect 778 5507 812 5526
rect 778 5492 812 5507
rect 250 5085 284 5095
rect 250 5061 284 5085
rect 250 4983 284 5017
rect 335 5073 369 5107
rect 335 5001 369 5035
rect 778 5405 812 5420
rect 778 5386 812 5405
rect 778 5303 812 5315
rect 778 5281 812 5303
rect 250 4915 284 4939
rect 250 4905 284 4915
rect 250 4847 284 4861
rect 250 4827 284 4847
rect 250 4779 284 4782
rect 250 4748 284 4779
rect 693 4876 727 4887
rect 693 4853 727 4876
rect 693 4808 727 4815
rect 693 4781 727 4808
rect 250 4677 284 4703
rect 250 4669 284 4677
rect 250 4609 284 4624
rect 250 4590 284 4609
rect 335 4754 369 4756
rect 335 4722 369 4754
rect 335 4652 369 4684
rect 335 4650 369 4652
rect 778 4793 812 4803
rect 778 4769 812 4793
rect 778 4725 812 4729
rect 778 4695 812 4725
rect 250 4541 284 4545
rect 778 4621 812 4655
rect 250 4511 284 4541
rect 415 4508 439 4542
rect 439 4508 449 4542
rect 496 4508 507 4542
rect 507 4508 530 4542
rect 577 4508 609 4542
rect 609 4508 611 4542
rect 658 4508 677 4542
rect 677 4508 692 4542
rect 740 4508 745 4542
rect 745 4508 774 4542
rect 967 6136 1001 6144
rect 967 6110 1001 6136
rect 1480 6119 1514 6144
rect 1480 6110 1514 6119
rect 967 6034 1001 6056
rect 967 6022 1001 6034
rect 967 5864 1001 5881
rect 967 5847 1001 5864
rect 967 5762 1001 5786
rect 967 5752 1001 5762
rect 1052 5847 1086 5881
rect 1052 5775 1086 5809
rect 1480 6051 1514 6069
rect 1480 6035 1514 6051
rect 1480 5983 1514 5994
rect 1480 5960 1514 5983
rect 1480 5915 1514 5919
rect 1480 5885 1514 5915
rect 1480 5813 1514 5843
rect 1480 5809 1514 5813
rect 967 5660 1001 5691
rect 967 5657 1001 5660
rect 1480 5745 1514 5767
rect 1480 5733 1514 5745
rect 1480 5677 1514 5691
rect 1480 5657 1514 5677
rect 1480 5609 1514 5615
rect 1480 5581 1514 5609
rect 967 5422 1001 5447
rect 967 5413 1001 5422
rect 967 5354 1001 5357
rect 967 5323 1001 5354
rect 967 5252 1001 5267
rect 967 5233 1001 5252
rect 1220 5427 1254 5461
rect 1292 5427 1326 5461
rect 1126 5256 1160 5290
rect 967 5150 1001 5178
rect 967 5144 1001 5150
rect 967 5082 1001 5089
rect 967 5055 1001 5082
rect 1126 5184 1160 5218
rect 1480 5439 1514 5451
rect 1480 5417 1514 5439
rect 1480 5371 1514 5378
rect 1480 5344 1514 5371
rect 1480 5303 1514 5305
rect 1480 5271 1514 5303
rect 1052 5148 1058 5151
rect 1058 5148 1086 5151
rect 1052 5117 1086 5148
rect 1052 5048 1086 5079
rect 1052 5045 1058 5048
rect 1058 5045 1086 5048
rect 1480 5201 1514 5232
rect 1480 5198 1514 5201
rect 3744 5216 3778 5244
rect 3744 5210 3746 5216
rect 3746 5210 3778 5216
rect 3816 5210 3850 5244
rect 3888 5210 3922 5244
rect 3960 5216 3994 5244
rect 4032 5216 4066 5244
rect 4104 5216 4138 5244
rect 3960 5210 3992 5216
rect 3992 5210 3994 5216
rect 4032 5210 4062 5216
rect 4062 5210 4066 5216
rect 4104 5210 4132 5216
rect 4132 5210 4138 5216
rect 1480 5133 1514 5159
rect 1480 5125 1514 5133
rect 1480 5065 1514 5086
rect 1480 5052 1514 5065
rect 1480 4997 1514 5013
rect 1480 4979 1514 4997
rect 1480 4929 1514 4940
rect 1480 4906 1514 4929
rect 967 4606 1001 4635
rect 967 4601 1001 4606
rect 967 4538 1001 4558
rect 967 4524 1001 4538
rect 967 4470 1001 4481
rect 967 4447 1001 4470
rect 967 4402 1001 4405
rect 967 4371 1001 4402
rect 250 4277 283 4311
rect 283 4277 284 4311
rect 415 4277 419 4311
rect 419 4277 449 4311
rect 496 4277 521 4311
rect 521 4277 530 4311
rect 577 4277 589 4311
rect 589 4277 611 4311
rect 658 4277 691 4311
rect 691 4277 692 4311
rect 740 4277 774 4311
rect 250 4208 284 4233
rect 250 4199 284 4208
rect 250 4140 284 4155
rect 250 4121 284 4140
rect 250 4072 284 4078
rect 250 4044 284 4072
rect 250 3970 284 4001
rect 250 3967 284 3970
rect 250 3902 284 3924
rect 250 3890 284 3902
rect 250 3834 284 3847
rect 250 3813 284 3834
rect 250 3766 284 3770
rect 250 3736 284 3766
rect 14 3694 48 3728
rect 14 3622 48 3656
rect 778 4074 812 4089
rect 778 4055 812 4074
rect 778 3972 812 4003
rect 778 3969 812 3972
rect 778 3904 812 3917
rect 778 3883 812 3904
rect 778 3802 812 3831
rect 778 3797 812 3802
rect 778 3734 812 3746
rect 778 3712 812 3734
rect 399 3515 405 3549
rect 405 3515 433 3549
rect 473 3515 507 3549
rect 547 3515 575 3549
rect 575 3515 581 3549
rect 621 3515 643 3549
rect 643 3515 655 3549
rect 695 3515 711 3549
rect 711 3515 729 3549
rect 967 4300 1001 4329
rect 967 4295 1001 4300
rect 967 4232 1001 4253
rect 967 4219 1001 4232
rect 1052 4782 1086 4793
rect 1052 4759 1086 4782
rect 1052 4713 1086 4721
rect 1052 4687 1086 4713
rect 1052 4062 1086 4089
rect 1052 4055 1086 4062
rect 1052 3994 1086 4017
rect 1052 3983 1086 3994
rect 1480 4861 1514 4867
rect 1480 4833 1514 4861
rect 1480 4793 1514 4794
rect 1480 4760 1514 4793
rect 1480 4691 1514 4721
rect 1480 4687 1514 4691
rect 1480 4623 1514 4648
rect 1480 4614 1514 4623
rect 1480 4555 1514 4575
rect 1480 4541 1514 4555
rect 1480 4487 1514 4502
rect 1480 4468 1514 4487
rect 1480 4419 1514 4429
rect 1480 4395 1514 4419
rect 1480 4351 1514 4356
rect 1480 4322 1514 4351
rect 1480 4249 1514 4283
rect 1480 4181 1514 4210
rect 1480 4176 1514 4181
rect 1480 4113 1514 4137
rect 1480 4103 1514 4113
rect 1480 4045 1514 4064
rect 1480 4030 1514 4045
rect 1480 3977 1514 3991
rect 1480 3957 1514 3977
rect 967 3858 1001 3859
rect 967 3825 1001 3858
rect 967 3756 1001 3785
rect 967 3751 1001 3756
rect 1480 3909 1514 3918
rect 1480 3884 1514 3909
rect 1480 3841 1514 3845
rect 1480 3811 1514 3841
rect 967 3688 1001 3711
rect 967 3677 1001 3688
rect 967 3620 1001 3638
rect 967 3604 1001 3620
rect 967 3552 1001 3565
rect 967 3531 1001 3552
rect 967 3484 1001 3492
rect 967 3458 1001 3484
rect 1052 3704 1086 3728
rect 1480 3739 1514 3772
rect 1480 3738 1514 3739
rect 1052 3694 1086 3704
rect 1162 3679 1196 3713
rect 1234 3679 1268 3713
rect 1306 3679 1340 3713
rect 1052 3630 1086 3656
rect 1052 3622 1086 3630
rect 1052 3556 1086 3584
rect 1052 3550 1086 3556
rect 1480 3671 1514 3699
rect 1480 3665 1514 3671
rect 1480 3603 1514 3626
rect 1480 3592 1514 3603
rect 1052 3482 1086 3512
rect 1162 3501 1196 3535
rect 1234 3501 1268 3535
rect 1306 3501 1340 3535
rect 1480 3535 1514 3553
rect 1480 3519 1514 3535
rect 1052 3478 1086 3482
rect 1480 3467 1514 3480
rect 1480 3446 1514 3467
rect 1480 3399 1514 3407
rect 1480 3373 1514 3399
rect 372 3326 385 3338
rect 385 3326 406 3338
rect 450 3326 453 3338
rect 453 3326 484 3338
rect 372 3304 406 3326
rect 450 3304 484 3326
rect 528 3326 555 3338
rect 555 3326 562 3338
rect 606 3326 623 3338
rect 623 3326 640 3338
rect 684 3326 691 3338
rect 691 3326 718 3338
rect 762 3327 796 3338
rect 528 3304 562 3326
rect 606 3304 640 3326
rect 684 3304 718 3326
rect 762 3304 778 3327
rect 778 3304 796 3327
rect 250 3290 284 3300
rect 250 3266 284 3290
rect 250 3188 284 3221
rect 250 3187 284 3188
rect 250 3120 284 3142
rect 250 3108 284 3120
rect 250 3052 284 3064
rect 250 3030 284 3052
rect 978 3280 1012 3314
rect 978 3208 1012 3242
rect 1480 3331 1514 3333
rect 1480 3299 1514 3331
rect 1480 3229 1514 3259
rect 1480 3225 1514 3229
rect 249 2939 283 2973
rect 249 2867 283 2901
rect 233 2779 267 2787
rect 233 2753 250 2779
rect 250 2753 267 2779
rect 233 2711 267 2714
rect 233 2680 250 2711
rect 250 2680 267 2711
rect 441 2823 475 2857
rect 513 2823 547 2857
rect 513 2731 547 2765
rect 585 2731 619 2765
rect 693 2763 727 2797
rect 693 2691 727 2725
rect 233 2609 250 2641
rect 250 2609 267 2641
rect 233 2607 267 2609
rect 778 2681 812 2714
rect 778 2680 812 2681
rect 778 2613 812 2637
rect 778 2603 812 2613
rect 233 2303 267 2324
rect 233 2290 250 2303
rect 250 2290 267 2303
rect 233 2201 250 2234
rect 250 2201 267 2234
rect 513 2529 547 2563
rect 585 2529 619 2563
rect 778 2545 812 2560
rect 778 2526 812 2545
rect 778 2477 812 2483
rect 778 2449 812 2477
rect 778 2375 812 2407
rect 778 2373 812 2375
rect 778 2307 812 2331
rect 778 2297 812 2307
rect 233 2200 267 2201
rect 233 2133 250 2145
rect 250 2133 267 2145
rect 233 2111 267 2133
rect 333 2100 337 2134
rect 337 2100 367 2134
rect 414 2100 439 2134
rect 439 2100 448 2134
rect 495 2100 507 2134
rect 507 2100 529 2134
rect 576 2100 609 2134
rect 609 2100 610 2134
rect 658 2100 677 2134
rect 677 2100 692 2134
rect 740 2100 745 2134
rect 745 2100 774 2134
rect 967 2918 1001 2919
rect 967 2885 1001 2918
rect 967 2680 1001 2714
rect 1480 3161 1514 3185
rect 1480 3151 1514 3161
rect 1480 3093 1514 3111
rect 1480 3077 1514 3093
rect 1480 3025 1514 3037
rect 1480 3003 1514 3025
rect 1052 2763 1086 2797
rect 1480 2957 1514 2963
rect 1480 2929 1514 2957
rect 1480 2855 1514 2889
rect 1052 2691 1086 2725
rect 1386 2708 1420 2737
rect 1386 2703 1420 2708
rect 967 2612 1001 2639
rect 967 2605 1001 2612
rect 967 2544 1001 2564
rect 967 2530 1001 2544
rect 1386 2631 1420 2665
rect 1386 2588 1420 2593
rect 967 2476 1001 2489
rect 967 2455 1001 2476
rect 967 2408 1001 2414
rect 967 2380 1001 2408
rect 967 2306 1001 2339
rect 967 2305 1001 2306
rect 1052 2530 1086 2564
rect 1386 2559 1420 2588
rect 1480 2651 1514 2681
rect 1480 2647 1514 2651
rect 1052 2458 1086 2492
rect 1480 2549 1514 2568
rect 1480 2534 1514 2549
rect 1386 2432 1420 2461
rect 1386 2427 1420 2432
rect 1386 2355 1420 2389
rect 1480 2379 1514 2393
rect 1480 2359 1514 2379
rect 1480 2311 1514 2319
rect 1480 2285 1514 2311
rect 1480 2243 1514 2245
rect 1480 2211 1514 2243
rect 1480 2141 1514 2171
rect 1480 2137 1514 2141
rect 345 1945 379 1946
rect 423 1945 457 1946
rect 501 1945 535 1946
rect 579 1945 613 1946
rect 345 1912 351 1945
rect 351 1912 379 1945
rect 423 1912 453 1945
rect 453 1912 457 1945
rect 501 1912 521 1945
rect 521 1912 535 1945
rect 579 1912 589 1945
rect 589 1912 613 1945
rect 657 1912 691 1946
rect 778 1878 812 1908
rect 778 1874 812 1878
rect 250 1728 284 1730
rect 250 1696 284 1728
rect 250 1626 284 1657
rect 250 1623 284 1626
rect 250 1558 284 1584
rect 250 1550 284 1558
rect 250 1490 284 1511
rect 250 1477 284 1490
rect 250 1422 284 1438
rect 250 1404 284 1422
rect 250 1354 284 1365
rect 250 1331 284 1354
rect 349 1770 383 1804
rect 349 1698 383 1732
rect 778 1810 812 1825
rect 778 1791 812 1810
rect 778 1742 812 1743
rect 778 1709 812 1742
rect 778 1640 812 1661
rect 778 1627 812 1640
rect 778 1572 812 1579
rect 778 1545 812 1572
rect 250 1286 284 1292
rect 250 1258 284 1286
rect 250 1218 284 1219
rect 250 1185 284 1218
rect 778 1300 812 1315
rect 778 1281 812 1300
rect 250 844 284 878
rect 250 776 284 800
rect 250 766 284 776
rect 250 708 284 722
rect 250 688 284 708
rect 250 640 284 644
rect 250 610 284 640
rect 250 538 284 565
rect 250 531 284 538
rect 349 1129 383 1133
rect 349 1099 383 1129
rect 349 1056 383 1061
rect 349 1027 383 1056
rect 349 837 383 871
rect 349 765 383 799
rect 349 693 383 727
rect 349 621 383 655
rect 349 549 383 583
rect 778 1164 812 1176
rect 778 1142 812 1164
rect 967 1932 1001 1938
rect 967 1904 1001 1932
rect 1480 2073 1514 2097
rect 1480 2063 1514 2073
rect 1480 2005 1514 2023
rect 1480 1989 1514 2005
rect 1480 1937 1514 1949
rect 1480 1915 1514 1937
rect 967 1830 1001 1859
rect 967 1825 1001 1830
rect 967 1762 1001 1780
rect 967 1746 1001 1762
rect 967 1694 1001 1701
rect 967 1667 1001 1694
rect 967 1592 1001 1622
rect 967 1588 1001 1592
rect 1052 1847 1086 1851
rect 1052 1817 1086 1847
rect 1480 1869 1514 1875
rect 1480 1841 1514 1869
rect 1162 1794 1196 1828
rect 1234 1794 1268 1828
rect 1306 1794 1340 1828
rect 1052 1773 1086 1779
rect 1052 1745 1086 1773
rect 1052 1699 1086 1707
rect 1052 1673 1086 1699
rect 1480 1767 1514 1801
rect 1480 1699 1514 1727
rect 1480 1693 1514 1699
rect 1052 1625 1086 1635
rect 1052 1601 1086 1625
rect 1162 1616 1196 1650
rect 1234 1616 1268 1650
rect 1306 1616 1340 1650
rect 1480 1631 1514 1653
rect 1480 1619 1514 1631
rect 967 1524 1001 1544
rect 967 1510 1001 1524
rect 967 1388 1001 1400
rect 967 1366 1001 1388
rect 1480 1563 1514 1579
rect 1480 1545 1514 1563
rect 1480 1495 1514 1505
rect 1480 1471 1514 1495
rect 1480 1427 1514 1431
rect 1480 1397 1514 1427
rect 967 1320 1001 1321
rect 967 1287 1001 1320
rect 967 1082 1001 1106
rect 967 1072 1001 1082
rect 967 1014 1001 1030
rect 967 996 1001 1014
rect 789 858 812 876
rect 812 858 823 876
rect 789 842 823 858
rect 861 842 895 876
rect 778 552 812 582
rect 778 548 812 552
rect 250 470 284 486
rect 250 452 284 470
rect 250 402 284 407
rect 250 373 284 402
rect 778 484 812 499
rect 778 465 812 484
rect 365 335 371 369
rect 371 335 399 369
rect 440 335 473 369
rect 473 335 474 369
rect 515 335 541 369
rect 541 335 549 369
rect 590 335 609 369
rect 609 335 624 369
rect 665 335 677 369
rect 677 335 699 369
rect 740 335 745 369
rect 745 335 774 369
rect 967 844 1001 870
rect 967 836 1001 844
rect 967 708 1001 728
rect 967 694 1001 708
rect 1052 1369 1086 1373
rect 1052 1339 1086 1369
rect 1052 1300 1086 1301
rect 1052 1267 1086 1300
rect 1480 1325 1514 1357
rect 1480 1323 1514 1325
rect 1480 1257 1514 1284
rect 1480 1250 1514 1257
rect 1480 1189 1514 1211
rect 1480 1177 1514 1189
rect 1480 1121 1514 1138
rect 1480 1104 1514 1121
rect 1480 1053 1514 1065
rect 1480 1031 1514 1053
rect 1209 924 1243 958
rect 1319 924 1353 958
rect 1480 985 1514 992
rect 1480 958 1514 985
rect 1052 615 1086 642
rect 1052 608 1086 615
rect 1052 547 1086 570
rect 1052 536 1086 547
rect 1480 917 1514 919
rect 1480 885 1514 917
rect 1480 815 1514 846
rect 1480 812 1514 815
rect 1480 747 1514 773
rect 1480 739 1514 747
rect 1480 679 1514 700
rect 1480 666 1514 679
rect 1480 611 1514 627
rect 1480 593 1514 611
rect 1480 543 1514 554
rect 1480 520 1514 543
rect 967 470 1001 484
rect 967 450 1001 470
rect 967 402 1001 407
rect 967 373 1001 402
rect 1480 475 1514 481
rect 1480 447 1514 475
rect 1077 335 1107 369
rect 1107 335 1111 369
rect 1150 335 1175 369
rect 1175 335 1184 369
rect 1223 335 1243 369
rect 1243 335 1257 369
rect 1296 335 1311 369
rect 1311 335 1330 369
rect 1369 335 1379 369
rect 1379 335 1403 369
rect 1442 335 1447 369
rect 1447 335 1476 369
rect 1785 5129 1804 5163
rect 1804 5129 1819 5163
rect 1860 5129 1872 5163
rect 1872 5129 1894 5163
rect 1935 5129 1940 5163
rect 1940 5129 1969 5163
rect 2010 5129 2042 5163
rect 2042 5129 2044 5163
rect 2085 5129 2110 5163
rect 2110 5129 2119 5163
rect 2160 5129 2178 5163
rect 2178 5129 2194 5163
rect 2235 5129 2246 5163
rect 2246 5129 2269 5163
rect 2310 5129 2314 5163
rect 2314 5129 2344 5163
rect 2385 5129 2416 5163
rect 2416 5129 2419 5163
rect 2460 5129 2484 5163
rect 2484 5129 2494 5163
rect 2536 5129 2552 5163
rect 2552 5129 2570 5163
rect 2612 5129 2620 5163
rect 2620 5129 2646 5163
rect 2688 5129 2722 5163
rect 2764 5129 2790 5163
rect 2790 5129 2798 5163
rect 2840 5129 2858 5163
rect 2858 5129 2874 5163
rect 2916 5129 2926 5163
rect 2926 5129 2950 5163
rect 2992 5129 2994 5163
rect 2994 5129 3026 5163
rect 3068 5130 3102 5163
rect 3068 5129 3079 5130
rect 3079 5129 3102 5130
rect 1669 5094 1703 5125
rect 1669 5091 1703 5094
rect 1669 5026 1703 5051
rect 1669 5017 1703 5026
rect 3079 5062 3113 5091
rect 3079 5057 3113 5062
rect 1669 4958 1703 4977
rect 1669 4943 1703 4958
rect 1669 4890 1703 4903
rect 1669 4869 1703 4890
rect 1669 4822 1703 4829
rect 1669 4795 1703 4822
rect 1669 4754 1703 4755
rect 1669 4721 1703 4754
rect 1669 4652 1703 4681
rect 1669 4647 1703 4652
rect 1669 4584 1703 4607
rect 1669 4573 1703 4584
rect 1669 4516 1703 4533
rect 1669 4499 1703 4516
rect 1669 4448 1703 4459
rect 1669 4425 1703 4448
rect 1669 4380 1703 4385
rect 1669 4351 1703 4380
rect 1669 4278 1703 4311
rect 1669 4277 1703 4278
rect 1669 4210 1703 4237
rect 1669 4203 1703 4210
rect 1669 4142 1703 4163
rect 1669 4129 1703 4142
rect 1669 4074 1703 4089
rect 1669 4055 1703 4074
rect 1669 4006 1703 4015
rect 1669 3981 1703 4006
rect 1669 3938 1703 3941
rect 1669 3907 1703 3938
rect 1669 3836 1703 3867
rect 1669 3833 1703 3836
rect 1669 3768 1703 3793
rect 1669 3759 1703 3768
rect 1669 3700 1703 3719
rect 1669 3685 1703 3700
rect 1669 3632 1703 3646
rect 1669 3612 1703 3632
rect 1669 3564 1703 3573
rect 1669 3539 1703 3564
rect 1669 3496 1703 3500
rect 1669 3466 1703 3496
rect 1669 3394 1703 3427
rect 1669 3393 1703 3394
rect 1669 3326 1703 3354
rect 1669 3320 1703 3326
rect 1669 3258 1703 3281
rect 1669 3247 1703 3258
rect 1669 3190 1703 3208
rect 1669 3174 1703 3190
rect 1669 3122 1703 3135
rect 1669 3101 1703 3122
rect 1669 3054 1703 3062
rect 1669 3028 1703 3054
rect 1669 2986 1703 2989
rect 1669 2955 1703 2986
rect 1669 2510 1703 2524
rect 1669 2490 1703 2510
rect 1669 2442 1703 2451
rect 1669 2417 1703 2442
rect 1669 2374 1703 2378
rect 1669 2344 1703 2374
rect 1669 2272 1703 2305
rect 1669 2271 1703 2272
rect 1669 2204 1703 2232
rect 1669 2198 1703 2204
rect 1669 2136 1703 2159
rect 1669 2125 1703 2136
rect 1669 2068 1703 2086
rect 1669 2052 1703 2068
rect 1669 2000 1703 2013
rect 1669 1979 1703 2000
rect 1669 1932 1703 1940
rect 1669 1906 1703 1932
rect 1669 1864 1703 1867
rect 1669 1833 1703 1864
rect 1669 1762 1703 1794
rect 1669 1760 1703 1762
rect 1669 1694 1703 1721
rect 1669 1687 1703 1694
rect 1669 1626 1703 1648
rect 1669 1614 1703 1626
rect 1669 1558 1703 1575
rect 1669 1541 1703 1558
rect 1669 1490 1703 1502
rect 1669 1468 1703 1490
rect 1669 1422 1703 1429
rect 1669 1395 1703 1422
rect 1669 1354 1703 1356
rect 1669 1322 1703 1354
rect 1669 1252 1703 1283
rect 1669 1249 1703 1252
rect 1669 1184 1703 1210
rect 1669 1176 1703 1184
rect 1669 1116 1703 1137
rect 1669 1103 1703 1116
rect 1669 1048 1703 1064
rect 1669 1030 1703 1048
rect 1669 980 1703 991
rect 1669 957 1703 980
rect 1669 912 1703 918
rect 1669 884 1703 912
rect 1669 844 1703 845
rect 1669 811 1703 844
rect 1669 742 1703 772
rect 1669 738 1703 742
rect 1669 674 1703 699
rect 1669 665 1703 674
rect 1669 606 1703 626
rect 1669 592 1703 606
rect 1669 538 1703 553
rect 1669 519 1703 538
rect 3079 4994 3113 5015
rect 3079 4981 3113 4994
rect 3079 4926 3113 4939
rect 3079 4905 3113 4926
rect 3079 4858 3113 4863
rect 3079 4829 3113 4858
rect 3079 4756 3113 4787
rect 3079 4753 3113 4756
rect 3079 4688 3113 4711
rect 3079 4677 3113 4688
rect 3079 4620 3113 4635
rect 3079 4601 3113 4620
rect 3079 4552 3113 4559
rect 3079 4525 3113 4552
rect 3079 4450 3113 4482
rect 3079 4448 3113 4450
rect 3079 4382 3113 4405
rect 3079 4371 3113 4382
rect 3079 4314 3113 4328
rect 3079 4294 3113 4314
rect 3079 4144 3113 4168
rect 3079 4134 3113 4144
rect 3079 4076 3113 4092
rect 3079 4058 3113 4076
rect 3079 4008 3113 4017
rect 3079 3983 3113 4008
rect 2620 3902 2654 3936
rect 2692 3902 2726 3936
rect 2764 3902 2798 3936
rect 3079 3940 3113 3942
rect 3079 3908 3113 3940
rect 3079 3736 3113 3743
rect 3079 3709 3113 3736
rect 2620 3578 2654 3612
rect 2692 3578 2726 3612
rect 2764 3578 2798 3612
rect 2836 3578 2870 3612
rect 3079 3634 3113 3645
rect 3079 3611 3113 3634
rect 3079 3532 3113 3548
rect 3079 3514 3113 3532
rect 3079 3362 3113 3388
rect 3079 3354 3113 3362
rect 2620 3278 2654 3312
rect 2692 3278 2726 3312
rect 2764 3278 2798 3312
rect 3079 3294 3113 3302
rect 3079 3268 3113 3294
rect 3079 3192 3113 3216
rect 3079 3182 3113 3192
rect 3079 3124 3113 3131
rect 3079 3097 3113 3124
rect 3079 3022 3113 3046
rect 3079 3012 3113 3022
rect 1752 2827 1786 2838
rect 1752 2804 1754 2827
rect 1754 2804 1786 2827
rect 1752 2732 1786 2766
rect 1752 2671 1754 2694
rect 1754 2671 1786 2694
rect 1752 2660 1786 2671
rect 2484 2813 2518 2838
rect 2484 2804 2518 2813
rect 2484 2732 2518 2766
rect 2484 2660 2518 2694
rect 3079 2954 3113 2961
rect 3079 2927 3113 2954
rect 2922 2511 2956 2545
rect 2994 2511 3028 2545
rect 3079 2580 3113 2594
rect 3079 2560 3113 2580
rect 3079 2512 3113 2519
rect 3079 2485 3113 2512
rect 3079 2410 3113 2444
rect 3079 2342 3113 2369
rect 3079 2335 3113 2342
rect 3079 2274 3113 2294
rect 3079 2260 3113 2274
rect 3079 2206 3113 2219
rect 3079 2185 3113 2206
rect 3079 2138 3113 2144
rect 3079 2110 3113 2138
rect 3079 1968 3113 1984
rect 3079 1950 3113 1968
rect 3079 1866 3113 1886
rect 3079 1852 3113 1866
rect 3079 1764 3113 1789
rect 3079 1755 3113 1764
rect 3079 1560 3113 1590
rect 3079 1556 3113 1560
rect 3079 1492 3113 1514
rect 3079 1480 3113 1492
rect 3079 1424 3113 1439
rect 3079 1405 3113 1424
rect 3079 1356 3113 1364
rect 3079 1330 3113 1356
rect 2620 1250 2654 1284
rect 2692 1250 2726 1284
rect 2764 1250 2798 1284
rect 3079 1186 3113 1204
rect 3079 1170 3113 1186
rect 3079 1118 3113 1130
rect 3079 1096 3113 1118
rect 3079 1050 3113 1057
rect 3079 1023 3113 1050
rect 3079 982 3113 984
rect 3079 950 3113 982
rect 3079 676 3113 695
rect 3079 661 3113 676
rect 3079 608 3113 623
rect 3079 589 3113 608
rect 3079 540 3113 551
rect 3079 517 3113 540
rect 1669 470 1703 480
rect 1669 446 1703 470
rect 1669 402 1703 407
rect 1669 373 1703 402
rect 3079 472 3113 479
rect 3079 445 3113 472
rect 1783 335 1788 369
rect 1788 335 1817 369
rect 1857 335 1890 369
rect 1890 335 1891 369
rect 1931 335 1958 369
rect 1958 335 1965 369
rect 2005 335 2026 369
rect 2026 335 2039 369
rect 2079 335 2094 369
rect 2094 335 2113 369
rect 2153 335 2162 369
rect 2162 335 2187 369
rect 2227 335 2230 369
rect 2230 335 2261 369
rect 2301 335 2332 369
rect 2332 335 2335 369
rect 2375 335 2400 369
rect 2400 335 2409 369
rect 2449 335 2468 369
rect 2468 335 2483 369
rect 2523 335 2536 369
rect 2536 335 2557 369
rect 2597 335 2604 369
rect 2604 335 2631 369
rect 2671 335 2672 369
rect 2672 335 2705 369
rect 2745 335 2774 369
rect 2774 335 2779 369
rect 2819 335 2842 369
rect 2842 335 2853 369
rect 2893 335 2910 369
rect 2910 335 2927 369
rect 2967 335 2978 369
rect 2978 335 3001 369
rect 3041 335 3046 369
rect 3046 335 3075 369
rect 3713 5148 3747 5153
rect 3792 5148 3826 5153
rect 3870 5148 3904 5153
rect 3948 5148 3982 5153
rect 4026 5148 4060 5153
rect 3713 5119 3730 5148
rect 3730 5119 3747 5148
rect 3792 5119 3798 5148
rect 3798 5119 3826 5148
rect 3870 5119 3900 5148
rect 3900 5119 3904 5148
rect 3948 5119 3968 5148
rect 3968 5119 3982 5148
rect 4026 5119 4036 5148
rect 4036 5119 4060 5148
rect 4104 5119 4138 5153
rect 4266 5048 4300 5058
rect 4266 5024 4300 5048
rect 4266 4946 4300 4954
rect 4266 4920 4300 4946
rect 4266 4844 4300 4850
rect 4266 4816 4300 4844
rect 13740 5540 13774 5574
rect 13812 5540 13846 5574
rect 13740 5466 13774 5500
rect 13812 5466 13846 5500
rect 14355 5271 14389 5305
rect 14427 5271 14461 5305
rect 14513 5271 14547 5305
rect 14585 5271 14619 5305
rect 4140 4326 4174 4332
rect 4140 4298 4174 4326
rect 4140 4252 4174 4259
rect 4140 4225 4174 4252
rect 4140 4178 4174 4186
rect 4140 4152 4174 4178
rect 4140 4104 4174 4113
rect 4140 4079 4174 4104
rect 4140 4030 4174 4040
rect 4140 4006 4174 4030
rect 4574 4561 4608 4595
rect 4646 4589 4680 4595
rect 4646 4561 4680 4589
rect 4266 4300 4300 4330
rect 4266 4296 4300 4300
rect 4266 4198 4300 4222
rect 4266 4188 4300 4198
rect 4266 3722 4300 3743
rect 4266 3709 4300 3722
rect 4266 3620 4300 3645
rect 4266 3611 4300 3620
rect 3550 3326 3584 3347
rect 3550 3313 3584 3326
rect 3550 3241 3584 3275
rect 4266 3518 4300 3548
rect 4266 3514 4300 3518
rect 4266 3246 4300 3273
rect 4266 3239 4300 3246
rect 4266 3178 4300 3200
rect 4266 3166 4300 3178
rect 4266 3110 4300 3127
rect 3780 3014 3814 3036
rect 3780 3002 3814 3014
rect 4266 3093 4300 3110
rect 4266 3042 4300 3054
rect 4266 3020 4300 3042
rect 4266 2974 4300 2981
rect 3780 2909 3814 2938
rect 3894 2916 3928 2950
rect 3966 2916 4000 2950
rect 4266 2947 4300 2974
rect 3780 2904 3814 2909
rect 4266 2906 4300 2908
rect 4266 2874 4300 2906
rect 3894 2824 3928 2858
rect 3966 2824 4000 2858
rect 4266 2804 4300 2835
rect 4266 2801 4300 2804
rect 4266 2736 4300 2763
rect 4266 2729 4300 2736
rect 4266 2668 4300 2691
rect 4266 2657 4300 2668
rect 4266 2600 4300 2619
rect 4266 2585 4300 2600
rect 3894 2548 3928 2582
rect 3966 2548 4000 2582
rect 4266 2532 4300 2547
rect 4266 2513 4300 2532
rect 4266 2464 4300 2475
rect 4266 2441 4300 2464
rect 3550 2223 3584 2257
rect 3550 2155 3584 2185
rect 3550 2151 3584 2155
rect 4266 2396 4300 2403
rect 4266 2369 4300 2396
rect 4266 2328 4300 2331
rect 4266 2297 4300 2328
rect 4266 2226 4300 2259
rect 4266 2225 4300 2226
rect 4266 1954 4300 1984
rect 4266 1950 4300 1954
rect 4266 1852 4300 1863
rect 4266 1829 4300 1852
rect 4140 1393 4174 1400
rect 4140 1366 4174 1393
rect 4140 1285 4174 1313
rect 4140 1279 4174 1285
rect 4140 1211 4174 1225
rect 4140 1191 4174 1211
rect 4140 1103 4174 1137
rect 4266 1342 4300 1364
rect 4266 1330 4300 1342
rect 4266 1240 4300 1250
rect 4266 1216 4300 1240
rect 4266 662 4300 692
rect 4266 658 4300 662
rect 4266 594 4300 616
rect 4266 582 4300 594
rect 4266 526 4300 540
rect 4266 506 4300 526
rect 4266 458 4300 465
rect 4266 431 4300 458
rect 3738 343 3772 377
rect 3810 350 3824 377
rect 3824 350 3844 377
rect 3882 350 3892 377
rect 3892 350 3916 377
rect 3954 350 3960 377
rect 3960 350 3988 377
rect 4026 350 4028 377
rect 4028 350 4060 377
rect 4098 350 4130 377
rect 4130 350 4132 377
rect 3810 343 3844 350
rect 3882 343 3916 350
rect 3954 343 3988 350
rect 4026 343 4060 350
rect 4098 343 4132 350
rect 4646 4385 4680 4402
rect 4646 4368 4680 4385
rect 4646 4283 4680 4299
rect 4646 4265 4680 4283
rect 4646 4181 4680 4196
rect 4646 4162 4680 4181
rect 4646 4011 4680 4024
rect 4646 3990 4680 4011
rect 4646 3943 4680 3944
rect 4646 3910 4680 3943
rect 4646 3841 4680 3864
rect 4646 3830 4680 3841
rect 4646 3773 4680 3785
rect 4646 3751 4680 3773
rect 4646 3705 4680 3706
rect 4646 3672 4680 3705
rect 4646 3603 4680 3627
rect 4646 3593 4680 3603
rect 4646 3535 4680 3548
rect 4646 3514 4680 3535
rect 4646 3365 4680 3388
rect 4646 3354 4680 3365
rect 4646 3297 4680 3309
rect 4646 3275 4680 3297
rect 4646 3229 4680 3230
rect 4646 3196 4680 3229
rect 4646 3059 4680 3070
rect 4646 3036 4680 3059
rect 4646 2991 4680 2994
rect 4646 2960 4680 2991
rect 4646 2889 4680 2918
rect 4646 2884 4680 2889
rect 4646 2821 4680 2842
rect 4646 2808 4680 2821
rect 4646 2753 4680 2766
rect 4646 2732 4680 2753
rect 4646 2685 4680 2690
rect 4646 2656 4680 2685
rect 4646 2583 4680 2614
rect 4646 2580 4680 2583
rect 4646 2515 4680 2538
rect 4646 2504 4680 2515
rect 4646 2447 4680 2462
rect 4646 2428 4680 2447
rect 4646 1665 4680 1681
rect 4646 1647 4680 1665
rect 4646 1597 4680 1600
rect 4646 1566 4680 1597
rect 4646 1495 4680 1520
rect 4646 1486 4680 1495
rect 4646 1427 4680 1440
rect 4646 1406 4680 1427
rect 4646 1359 4680 1360
rect 4646 1326 4680 1359
rect 4646 441 4680 448
rect 4646 414 4680 441
rect 4646 305 4680 330
rect 4646 296 4680 305
rect 4841 5117 4875 5120
rect 4913 5117 4947 5120
rect 4985 5117 5019 5120
rect 5057 5117 5091 5120
rect 5129 5117 5163 5120
rect 5201 5117 5235 5120
rect 5273 5117 5307 5120
rect 5345 5117 5379 5120
rect 5417 5117 5451 5120
rect 5489 5117 5523 5120
rect 5561 5117 5595 5120
rect 5633 5117 5667 5120
rect 5705 5117 5739 5120
rect 5777 5117 5811 5120
rect 5849 5117 5883 5120
rect 5921 5117 5955 5120
rect 5993 5117 6027 5120
rect 6065 5117 6099 5120
rect 6137 5117 6171 5120
rect 6209 5117 6243 5120
rect 6281 5117 6315 5120
rect 6353 5117 6387 5120
rect 6425 5117 6459 5120
rect 6497 5117 6531 5120
rect 6569 5117 6603 5120
rect 6641 5117 6675 5120
rect 6713 5117 6747 5120
rect 6785 5117 6819 5120
rect 6858 5117 6892 5120
rect 6931 5117 6965 5120
rect 7004 5117 7038 5120
rect 7077 5117 7111 5120
rect 7150 5117 7184 5120
rect 7223 5117 7257 5120
rect 7296 5117 7330 5120
rect 7369 5117 7403 5120
rect 7442 5117 7476 5120
rect 7515 5117 7549 5120
rect 7588 5117 7622 5120
rect 7661 5117 7695 5120
rect 7734 5117 7768 5120
rect 7807 5117 7841 5120
rect 7880 5117 7914 5120
rect 7953 5117 7987 5120
rect 8026 5117 8060 5120
rect 8099 5117 8133 5120
rect 8172 5117 8206 5120
rect 8245 5117 8279 5120
rect 8318 5117 8352 5120
rect 8391 5117 8425 5120
rect 8464 5117 8498 5120
rect 8537 5117 8571 5120
rect 8610 5117 8644 5120
rect 8683 5117 8717 5120
rect 8756 5117 8790 5120
rect 8829 5117 8863 5120
rect 8902 5117 8936 5120
rect 8975 5117 9009 5120
rect 9048 5117 9082 5120
rect 9121 5117 9155 5120
rect 9194 5117 9228 5120
rect 9267 5117 9301 5120
rect 9340 5117 9374 5120
rect 9413 5117 9447 5120
rect 4841 5086 4868 5117
rect 4868 5086 4875 5117
rect 4913 5086 4936 5117
rect 4936 5086 4947 5117
rect 4985 5086 5004 5117
rect 5004 5086 5019 5117
rect 5057 5086 5072 5117
rect 5072 5086 5091 5117
rect 5129 5086 5140 5117
rect 5140 5086 5163 5117
rect 5201 5086 5208 5117
rect 5208 5086 5235 5117
rect 5273 5086 5276 5117
rect 5276 5086 5307 5117
rect 5345 5086 5378 5117
rect 5378 5086 5379 5117
rect 5417 5086 5446 5117
rect 5446 5086 5451 5117
rect 5489 5086 5514 5117
rect 5514 5086 5523 5117
rect 5561 5086 5582 5117
rect 5582 5086 5595 5117
rect 5633 5086 5650 5117
rect 5650 5086 5667 5117
rect 5705 5086 5718 5117
rect 5718 5086 5739 5117
rect 5777 5086 5786 5117
rect 5786 5086 5811 5117
rect 5849 5086 5854 5117
rect 5854 5086 5883 5117
rect 5921 5086 5922 5117
rect 5922 5086 5955 5117
rect 5993 5086 6024 5117
rect 6024 5086 6027 5117
rect 6065 5086 6092 5117
rect 6092 5086 6099 5117
rect 6137 5086 6160 5117
rect 6160 5086 6171 5117
rect 6209 5086 6228 5117
rect 6228 5086 6243 5117
rect 6281 5086 6296 5117
rect 6296 5086 6315 5117
rect 6353 5086 6364 5117
rect 6364 5086 6387 5117
rect 6425 5086 6432 5117
rect 6432 5086 6459 5117
rect 6497 5086 6500 5117
rect 6500 5086 6531 5117
rect 6569 5086 6602 5117
rect 6602 5086 6603 5117
rect 6641 5086 6670 5117
rect 6670 5086 6675 5117
rect 6713 5086 6738 5117
rect 6738 5086 6747 5117
rect 6785 5086 6806 5117
rect 6806 5086 6819 5117
rect 6858 5086 6874 5117
rect 6874 5086 6892 5117
rect 6931 5086 6942 5117
rect 6942 5086 6965 5117
rect 7004 5086 7010 5117
rect 7010 5086 7038 5117
rect 7077 5086 7078 5117
rect 7078 5086 7111 5117
rect 7150 5086 7180 5117
rect 7180 5086 7184 5117
rect 7223 5086 7248 5117
rect 7248 5086 7257 5117
rect 7296 5086 7316 5117
rect 7316 5086 7330 5117
rect 7369 5086 7384 5117
rect 7384 5086 7403 5117
rect 7442 5086 7452 5117
rect 7452 5086 7476 5117
rect 7515 5086 7520 5117
rect 7520 5086 7549 5117
rect 7588 5086 7622 5117
rect 7661 5086 7690 5117
rect 7690 5086 7695 5117
rect 7734 5086 7758 5117
rect 7758 5086 7768 5117
rect 7807 5086 7826 5117
rect 7826 5086 7841 5117
rect 7880 5086 7894 5117
rect 7894 5086 7914 5117
rect 7953 5086 7962 5117
rect 7962 5086 7987 5117
rect 8026 5086 8030 5117
rect 8030 5086 8060 5117
rect 8099 5086 8132 5117
rect 8132 5086 8133 5117
rect 8172 5086 8200 5117
rect 8200 5086 8206 5117
rect 8245 5086 8268 5117
rect 8268 5086 8279 5117
rect 8318 5086 8336 5117
rect 8336 5086 8352 5117
rect 8391 5086 8404 5117
rect 8404 5086 8425 5117
rect 8464 5086 8472 5117
rect 8472 5086 8498 5117
rect 8537 5086 8540 5117
rect 8540 5086 8571 5117
rect 8610 5086 8642 5117
rect 8642 5086 8644 5117
rect 8683 5086 8710 5117
rect 8710 5086 8717 5117
rect 8756 5086 8778 5117
rect 8778 5086 8790 5117
rect 8829 5086 8846 5117
rect 8846 5086 8863 5117
rect 8902 5086 8914 5117
rect 8914 5086 8936 5117
rect 8975 5086 8982 5117
rect 8982 5086 9009 5117
rect 9048 5086 9050 5117
rect 9050 5086 9082 5117
rect 9121 5086 9152 5117
rect 9152 5086 9155 5117
rect 9194 5086 9220 5117
rect 9220 5086 9228 5117
rect 9267 5086 9288 5117
rect 9288 5086 9301 5117
rect 9340 5086 9356 5117
rect 9356 5086 9374 5117
rect 9413 5086 9424 5117
rect 9424 5086 9447 5117
rect 9506 5083 9526 5117
rect 9526 5083 9540 5117
rect 9580 5083 9594 5117
rect 9594 5083 9614 5117
rect 9654 5083 9662 5117
rect 9662 5083 9688 5117
rect 9728 5083 9730 5117
rect 9730 5083 9762 5117
rect 9802 5083 9832 5117
rect 9832 5083 9836 5117
rect 9876 5083 9900 5117
rect 9900 5083 9910 5117
rect 9950 5083 9968 5117
rect 9968 5083 9984 5117
rect 10024 5083 10036 5117
rect 10036 5083 10058 5117
rect 10098 5083 10104 5117
rect 10104 5083 10132 5117
rect 10172 5083 10206 5117
rect 10246 5083 10274 5117
rect 10274 5083 10280 5117
rect 10320 5083 10342 5117
rect 10342 5083 10354 5117
rect 10394 5083 10410 5117
rect 10410 5083 10428 5117
rect 10468 5083 10478 5117
rect 10478 5083 10502 5117
rect 10542 5083 10546 5117
rect 10546 5083 10576 5117
rect 10616 5083 10648 5117
rect 10648 5083 10650 5117
rect 10690 5083 10716 5117
rect 10716 5083 10724 5117
rect 10764 5083 10784 5117
rect 10784 5083 10798 5117
rect 10838 5083 10852 5117
rect 10852 5083 10872 5117
rect 10912 5083 10920 5117
rect 10920 5083 10946 5117
rect 10986 5083 10988 5117
rect 10988 5083 11020 5117
rect 11060 5083 11090 5117
rect 11090 5083 11094 5117
rect 11134 5083 11158 5117
rect 11158 5083 11168 5117
rect 11207 5083 11226 5117
rect 11226 5083 11241 5117
rect 11280 5083 11294 5117
rect 11294 5083 11314 5117
rect 11353 5083 11362 5117
rect 11362 5083 11387 5117
rect 11609 5083 11634 5117
rect 11634 5083 11643 5117
rect 11683 5083 11702 5117
rect 11702 5083 11717 5117
rect 11757 5083 11770 5117
rect 11770 5083 11791 5117
rect 11832 5083 11838 5117
rect 11838 5083 11866 5117
rect 11907 5083 11940 5117
rect 11940 5083 11941 5117
rect 11982 5083 12008 5117
rect 12008 5083 12016 5117
rect 12057 5083 12076 5117
rect 12076 5083 12091 5117
rect 12132 5083 12144 5117
rect 12144 5083 12166 5117
rect 12207 5083 12212 5117
rect 12212 5083 12241 5117
rect 12282 5083 12314 5117
rect 12314 5083 12316 5117
rect 12357 5083 12382 5117
rect 12382 5083 12391 5117
rect 12432 5083 12450 5117
rect 12450 5083 12466 5117
rect 12507 5083 12518 5117
rect 12518 5083 12541 5117
rect 12675 5084 12709 5106
rect 4835 5003 4869 5024
rect 4835 4990 4869 5003
rect 4835 4935 4869 4952
rect 4835 4918 4869 4935
rect 4835 4765 4869 4771
rect 4835 4737 4869 4765
rect 4835 4663 4869 4690
rect 4835 4656 4869 4663
rect 4835 4595 4869 4610
rect 4835 4576 4869 4595
rect 4835 4527 4869 4530
rect 4835 4496 4869 4527
rect 4835 4425 4869 4450
rect 4835 4416 4869 4425
rect 4835 4357 4869 4370
rect 4835 4336 4869 4357
rect 4835 4289 4869 4290
rect 4835 4256 4869 4289
rect 4835 4187 4869 4210
rect 4835 4176 4869 4187
rect 9468 4987 9502 5005
rect 9468 4971 9502 4987
rect 9468 4919 9502 4932
rect 9468 4898 9502 4919
rect 9706 4887 9740 4921
rect 9778 4887 9812 4921
rect 9942 4887 9976 4921
rect 10014 4887 10048 4921
rect 9468 4851 9502 4859
rect 9468 4825 9502 4851
rect 12675 5072 12709 5084
rect 12675 5016 12709 5032
rect 12675 4998 12709 5016
rect 12675 4948 12709 4958
rect 12675 4924 12709 4948
rect 9468 4783 9502 4786
rect 9468 4752 9502 4783
rect 9468 4681 9502 4713
rect 9468 4679 9502 4681
rect 9468 4613 9502 4640
rect 9468 4606 9502 4613
rect 9468 4545 9502 4567
rect 9468 4533 9502 4545
rect 9468 4477 9502 4494
rect 9468 4460 9502 4477
rect 9468 4409 9502 4421
rect 9468 4387 9502 4409
rect 9468 4341 9502 4348
rect 9468 4314 9502 4341
rect 9468 4273 9502 4275
rect 9468 4241 9502 4273
rect 9468 4171 9502 4202
rect 9468 4168 9502 4171
rect 9468 4103 9502 4128
rect 9468 4094 9502 4103
rect 9468 4035 9502 4054
rect 9468 4020 9502 4035
rect 9468 3967 9502 3980
rect 9468 3946 9502 3967
rect 9468 3899 9502 3906
rect 9468 3872 9502 3899
rect 9468 3831 9502 3832
rect 9468 3798 9502 3831
rect 5049 3744 8971 3746
rect 9010 3744 9044 3746
rect 9083 3744 9117 3746
rect 9156 3744 9190 3746
rect 9229 3744 9263 3746
rect 9302 3744 9336 3746
rect 5049 3710 5066 3744
rect 5066 3710 5101 3744
rect 5101 3710 5135 3744
rect 5135 3710 5170 3744
rect 5170 3710 5204 3744
rect 5204 3710 5239 3744
rect 5239 3710 5273 3744
rect 5273 3710 5308 3744
rect 5308 3710 5342 3744
rect 5342 3710 5377 3744
rect 5377 3710 5411 3744
rect 5411 3710 5446 3744
rect 5446 3710 5480 3744
rect 5480 3710 5515 3744
rect 5515 3710 5549 3744
rect 5549 3710 5584 3744
rect 5584 3710 5618 3744
rect 5618 3710 5653 3744
rect 5653 3710 5687 3744
rect 5687 3710 5722 3744
rect 5722 3710 5756 3744
rect 5756 3710 5791 3744
rect 5791 3710 5825 3744
rect 5825 3710 5860 3744
rect 5860 3710 5894 3744
rect 5894 3710 5929 3744
rect 5049 3676 5929 3710
rect 5049 3642 5066 3676
rect 5066 3642 5101 3676
rect 5101 3642 5135 3676
rect 5135 3642 5170 3676
rect 5170 3642 5204 3676
rect 5204 3642 5239 3676
rect 5239 3642 5273 3676
rect 5273 3642 5308 3676
rect 5308 3642 5342 3676
rect 5342 3642 5377 3676
rect 5377 3642 5411 3676
rect 5411 3642 5446 3676
rect 5446 3642 5480 3676
rect 5480 3642 5515 3676
rect 5515 3642 5549 3676
rect 5549 3642 5584 3676
rect 5584 3642 5618 3676
rect 5618 3642 5653 3676
rect 5653 3642 5687 3676
rect 5687 3642 5722 3676
rect 5722 3642 5756 3676
rect 5756 3642 5791 3676
rect 5791 3642 5825 3676
rect 5825 3642 5860 3676
rect 5860 3642 5894 3676
rect 5894 3642 5929 3676
rect 5929 3642 8971 3744
rect 9010 3712 9044 3744
rect 9083 3712 9117 3744
rect 9156 3712 9190 3744
rect 9229 3712 9263 3744
rect 9302 3712 9336 3744
rect 9375 3712 9409 3746
rect 9468 3729 9502 3758
rect 9468 3724 9502 3729
rect 9010 3642 9044 3674
rect 9083 3642 9117 3674
rect 9156 3642 9190 3674
rect 9229 3642 9263 3674
rect 9302 3642 9336 3674
rect 5049 3640 8971 3642
rect 9010 3640 9044 3642
rect 9083 3640 9117 3642
rect 9156 3640 9190 3642
rect 9229 3640 9263 3642
rect 9302 3640 9336 3642
rect 9375 3640 9409 3674
rect 9468 3661 9502 3684
rect 9468 3650 9502 3661
rect 9468 3593 9502 3610
rect 9468 3576 9502 3593
rect 9468 3525 9502 3536
rect 9468 3502 9502 3525
rect 4835 3303 4869 3333
rect 4835 3299 4869 3303
rect 4835 3235 4869 3255
rect 4835 3221 4869 3235
rect 4835 3167 4869 3177
rect 4835 3143 4869 3167
rect 4835 3065 4869 3099
rect 9468 3321 9502 3350
rect 9468 3316 9502 3321
rect 9468 3253 9502 3261
rect 9468 3227 9502 3253
rect 4835 2997 4869 3021
rect 4835 2987 4869 2997
rect 6970 3062 7004 3096
rect 7042 3062 7076 3096
rect 4958 3029 4992 3058
rect 4958 3024 4980 3029
rect 4980 3024 4992 3029
rect 5030 3024 5064 3058
rect 4835 2929 4869 2943
rect 4835 2909 4869 2929
rect 4835 2861 4869 2865
rect 4835 2831 4869 2861
rect 4835 2759 4869 2787
rect 4835 2753 4869 2759
rect 4958 2759 4980 2783
rect 4980 2759 4992 2783
rect 4958 2749 4992 2759
rect 5030 2749 5064 2783
rect 6970 2749 7004 2783
rect 7042 2749 7076 2783
rect 7218 3031 7252 3065
rect 7290 3031 7324 3065
rect 9208 3031 9242 3065
rect 9280 3031 9314 3065
rect 9623 4806 9657 4840
rect 9623 4733 9657 4767
rect 9623 4660 9657 4694
rect 9623 4587 9657 4621
rect 9623 4514 9657 4548
rect 9623 4441 9657 4475
rect 9623 4368 9657 4402
rect 9623 4295 9657 4329
rect 9623 4222 9657 4256
rect 9623 4148 9657 4182
rect 9623 4074 9657 4108
rect 9623 4000 9657 4034
rect 9623 3926 9657 3960
rect 9623 3852 9657 3886
rect 9623 3778 9657 3812
rect 9623 3704 9657 3738
rect 9623 3630 9657 3664
rect 9623 3556 9657 3590
rect 9623 3482 9657 3516
rect 9623 3408 9657 3442
rect 9623 3334 9657 3368
rect 9623 3260 9657 3294
rect 9623 3186 9657 3220
rect 9623 3112 9657 3146
rect 9623 3038 9657 3072
rect 9859 4806 9893 4840
rect 9859 4733 9893 4767
rect 9859 4660 9893 4694
rect 9859 4587 9893 4621
rect 9859 4514 9893 4548
rect 9859 4441 9893 4475
rect 9859 4368 9893 4402
rect 9859 4295 9893 4329
rect 9859 4222 9893 4256
rect 9859 4149 9893 4183
rect 9859 4076 9893 4110
rect 9859 4003 9893 4037
rect 9859 3930 9893 3964
rect 9859 3857 9893 3891
rect 9859 3783 9893 3817
rect 9859 3709 9893 3743
rect 9859 3635 9893 3669
rect 9859 3561 9893 3595
rect 9859 3487 9893 3521
rect 9859 3413 9893 3447
rect 9859 3339 9893 3373
rect 9859 3265 9893 3299
rect 9859 3191 9893 3225
rect 9859 3117 9893 3151
rect 9859 3043 9893 3077
rect 10095 4767 10129 4801
rect 10095 4695 10129 4729
rect 10095 4623 10129 4657
rect 10095 4551 10129 4585
rect 10095 4479 10129 4513
rect 10095 4407 10129 4441
rect 10095 4335 10129 4369
rect 10095 4263 10129 4297
rect 10095 4191 10129 4225
rect 10095 4119 10129 4153
rect 10095 4047 10129 4081
rect 10095 3975 10129 4009
rect 10095 3903 10129 3937
rect 10095 3831 10129 3865
rect 10095 3759 10129 3793
rect 10095 3687 10129 3721
rect 10095 3615 10129 3649
rect 10095 3543 10129 3577
rect 10095 3471 10129 3505
rect 10095 3399 10129 3433
rect 10095 3327 10129 3361
rect 10095 3255 10129 3289
rect 10095 3183 10129 3217
rect 10095 3111 10129 3145
rect 10095 3038 10129 3072
rect 10095 2965 10129 2999
rect 10423 4757 10457 4791
rect 10423 4677 10457 4711
rect 10423 4597 10457 4631
rect 10423 4518 10457 4552
rect 10423 4439 10457 4473
rect 10423 4360 10457 4394
rect 10423 4281 10457 4315
rect 10423 4202 10457 4236
rect 10423 4123 10457 4157
rect 11130 4757 11164 4791
rect 11130 4677 11164 4711
rect 11130 4597 11164 4631
rect 11130 4518 11164 4552
rect 11130 4439 11164 4473
rect 11130 4360 11164 4394
rect 11130 4281 11164 4315
rect 11130 4202 11164 4236
rect 11130 4123 11164 4157
rect 12675 4880 12709 4884
rect 12675 4850 12709 4880
rect 11290 4750 11324 4784
rect 11372 4750 11406 4784
rect 11454 4750 11488 4784
rect 11536 4750 11570 4784
rect 11618 4750 11652 4784
rect 11700 4750 11734 4784
rect 11290 4674 11324 4708
rect 11372 4674 11406 4708
rect 11454 4674 11488 4708
rect 11536 4674 11570 4708
rect 11618 4674 11652 4708
rect 11700 4674 11734 4708
rect 11290 4598 11324 4632
rect 11372 4598 11406 4632
rect 11454 4598 11488 4632
rect 11536 4598 11570 4632
rect 11618 4598 11652 4632
rect 11700 4598 11734 4632
rect 11290 4521 11324 4555
rect 11372 4521 11406 4555
rect 11454 4521 11488 4555
rect 11536 4521 11570 4555
rect 11618 4521 11652 4555
rect 11700 4521 11734 4555
rect 11290 4444 11324 4478
rect 11372 4444 11406 4478
rect 11454 4444 11488 4478
rect 11536 4444 11570 4478
rect 11618 4444 11652 4478
rect 11700 4444 11734 4478
rect 11290 4367 11324 4401
rect 11372 4367 11406 4401
rect 11454 4367 11488 4401
rect 11536 4367 11570 4401
rect 11618 4367 11652 4401
rect 11700 4367 11734 4401
rect 11290 4290 11324 4324
rect 11372 4290 11406 4324
rect 11454 4290 11488 4324
rect 11536 4290 11570 4324
rect 11618 4290 11652 4324
rect 11700 4290 11734 4324
rect 11290 4213 11324 4247
rect 11372 4213 11406 4247
rect 11454 4213 11488 4247
rect 11536 4213 11570 4247
rect 11618 4213 11652 4247
rect 11700 4213 11734 4247
rect 11290 4136 11324 4170
rect 11372 4136 11406 4170
rect 11454 4136 11488 4170
rect 11536 4136 11570 4170
rect 11618 4136 11652 4170
rect 11700 4136 11734 4170
rect 7218 2751 7252 2785
rect 7290 2751 7324 2785
rect 9147 2751 9181 2785
rect 9219 2751 9253 2785
rect 4835 2691 4869 2709
rect 4835 2675 4869 2691
rect 4835 2623 4869 2631
rect 4835 2597 4869 2623
rect 4835 2521 4869 2553
rect 4835 2519 4869 2521
rect 4835 2453 4869 2476
rect 4835 2442 4869 2453
rect 4958 2426 4992 2445
rect 4958 2411 4980 2426
rect 4980 2411 4992 2426
rect 5030 2411 5064 2445
rect 6970 2390 7004 2424
rect 7042 2390 7076 2424
rect 5067 2173 5101 2207
rect 5139 2173 5173 2207
rect 6970 2152 7004 2186
rect 7042 2152 7076 2186
rect 7218 2464 7252 2498
rect 7290 2464 7324 2498
rect 9208 2426 9242 2460
rect 9280 2426 9314 2460
rect 7218 2148 7252 2182
rect 7290 2148 7324 2182
rect 9230 2148 9264 2182
rect 9302 2156 9314 2182
rect 9314 2156 9336 2182
rect 9302 2148 9336 2156
rect 9859 2193 9893 2227
rect 5049 1571 5066 1572
rect 5066 1571 5083 1572
rect 5121 1571 5135 1572
rect 5135 1571 5155 1572
rect 5193 1571 5204 1572
rect 5204 1571 5227 1572
rect 5265 1571 5273 1572
rect 5273 1571 5299 1572
rect 5337 1571 5342 1572
rect 5342 1571 5371 1572
rect 5409 1571 5411 1572
rect 5411 1571 5443 1572
rect 5049 1538 5083 1571
rect 5121 1538 5155 1571
rect 5193 1538 5227 1571
rect 5265 1538 5299 1571
rect 5337 1538 5371 1571
rect 5409 1538 5443 1571
rect 5481 1538 5515 1572
rect 5553 1571 5584 1572
rect 5584 1571 5587 1572
rect 5625 1571 5653 1572
rect 5653 1571 5659 1572
rect 5697 1571 5722 1572
rect 5722 1571 5731 1572
rect 5769 1571 5791 1572
rect 5791 1571 5803 1572
rect 5841 1571 5860 1572
rect 5860 1571 5875 1572
rect 5553 1538 5587 1571
rect 5625 1538 5659 1571
rect 5697 1538 5731 1571
rect 5769 1538 5803 1571
rect 5841 1538 5875 1571
rect 5913 1538 5929 1572
rect 5929 1538 5947 1572
rect 5985 1538 6019 1572
rect 6057 1538 6091 1572
rect 6129 1538 6163 1572
rect 6201 1538 6235 1572
rect 6273 1538 6307 1572
rect 6345 1538 6379 1572
rect 6417 1538 6451 1572
rect 6489 1538 6523 1572
rect 6561 1538 6595 1572
rect 6633 1538 6667 1572
rect 6705 1538 6739 1572
rect 6777 1538 6811 1572
rect 6849 1538 6883 1572
rect 6921 1538 6955 1572
rect 6993 1538 7027 1572
rect 7065 1538 7099 1572
rect 7137 1538 7171 1572
rect 7209 1538 7243 1572
rect 7281 1538 7315 1572
rect 7353 1538 7387 1572
rect 7425 1538 7459 1572
rect 7497 1538 7531 1572
rect 7569 1538 7603 1572
rect 7641 1538 7675 1572
rect 7713 1538 7747 1572
rect 7785 1538 7819 1572
rect 7857 1538 7891 1572
rect 7929 1538 7963 1572
rect 8001 1538 8035 1572
rect 8073 1538 8107 1572
rect 8145 1538 8179 1572
rect 8217 1538 8251 1572
rect 8289 1538 8323 1572
rect 8361 1538 8395 1572
rect 8433 1538 8467 1572
rect 8505 1538 8539 1572
rect 8577 1538 8611 1572
rect 8649 1538 8683 1572
rect 8721 1538 8755 1572
rect 8793 1538 8827 1572
rect 8865 1538 8899 1572
rect 8937 1538 8971 1572
rect 9010 1538 9044 1572
rect 9083 1538 9117 1572
rect 9156 1538 9190 1572
rect 9229 1538 9263 1572
rect 9302 1538 9336 1572
rect 9375 1538 9409 1572
rect 4835 413 4869 436
rect 4835 402 4869 413
rect 4835 311 4869 328
rect 4835 294 4869 311
rect 9468 1471 9502 1502
rect 9468 1468 9502 1471
rect 9468 1402 9502 1428
rect 9468 1394 9502 1402
rect 9468 1333 9502 1354
rect 9468 1320 9502 1333
rect 9468 1264 9502 1280
rect 9468 1246 9502 1264
rect 9468 1195 9502 1206
rect 9468 1172 9502 1195
rect 9468 1126 9502 1132
rect 9468 1098 9502 1126
rect 9468 1057 9502 1058
rect 9468 1024 9502 1057
rect 9468 953 9502 984
rect 9468 950 9502 953
rect 9468 884 9502 910
rect 9468 876 9502 884
rect 9468 815 9502 836
rect 9468 802 9502 815
rect 9468 746 9502 763
rect 9468 729 9502 746
rect 9468 677 9502 690
rect 9468 656 9502 677
rect 9623 2102 9657 2136
rect 9623 2028 9657 2062
rect 9623 1954 9657 1988
rect 9623 1880 9657 1914
rect 9623 1806 9657 1840
rect 9623 1732 9657 1766
rect 9623 1658 9657 1692
rect 9623 1584 9657 1618
rect 9623 1510 9657 1544
rect 9623 1436 9657 1470
rect 9623 1361 9657 1395
rect 9623 1286 9657 1320
rect 9623 1211 9657 1245
rect 9623 1136 9657 1170
rect 9623 1061 9657 1095
rect 9623 986 9657 1020
rect 9623 911 9657 945
rect 9623 836 9657 870
rect 9623 761 9657 795
rect 9623 686 9657 720
rect 9859 2118 9893 2152
rect 9859 2043 9893 2077
rect 9859 1968 9893 2002
rect 9859 1893 9893 1927
rect 9859 1818 9893 1852
rect 9859 1743 9893 1777
rect 9859 1668 9893 1702
rect 9859 1593 9893 1627
rect 9859 1518 9893 1552
rect 9859 1443 9893 1477
rect 9859 1368 9893 1402
rect 9859 1293 9893 1327
rect 9859 1218 9893 1252
rect 9859 1142 9893 1176
rect 9859 1066 9893 1100
rect 9859 990 9893 1024
rect 9859 914 9893 948
rect 9859 838 9893 872
rect 9859 762 9893 796
rect 9859 686 9893 720
rect 10095 2029 10129 2063
rect 10095 1955 10129 1989
rect 10095 1881 10129 1915
rect 10095 1807 10129 1841
rect 10095 1733 10129 1767
rect 10095 1659 10129 1693
rect 10095 1585 10129 1619
rect 10095 1511 10129 1545
rect 10095 1436 10129 1470
rect 10095 1361 10129 1395
rect 10095 1286 10129 1320
rect 10095 1211 10129 1245
rect 10095 1136 10129 1170
rect 10095 1061 10129 1095
rect 10095 986 10129 1020
rect 10095 911 10129 945
rect 10095 836 10129 870
rect 10095 761 10129 795
rect 10095 686 10129 720
rect 10400 3952 10434 3954
rect 10400 3920 10434 3952
rect 10400 3850 10434 3882
rect 10400 3848 10434 3850
rect 11130 3952 11164 3954
rect 11130 3920 11164 3952
rect 11130 3850 11164 3882
rect 11130 3848 11164 3850
rect 10620 3756 10654 3790
rect 10692 3756 10726 3790
rect 10764 3756 10798 3790
rect 10836 3756 10870 3790
rect 10908 3756 10942 3790
rect 10980 3756 11014 3790
rect 11052 3756 11086 3790
rect 10400 3696 10434 3698
rect 10400 3664 10434 3696
rect 10400 3594 10434 3626
rect 10400 3592 10434 3594
rect 10400 3440 10434 3442
rect 10400 3408 10434 3440
rect 10400 3338 10434 3370
rect 10400 3336 10434 3338
rect 11860 4757 11894 4791
rect 11860 4677 11894 4711
rect 11860 4597 11894 4631
rect 11860 4518 11894 4552
rect 11860 4439 11894 4473
rect 11860 4360 11894 4394
rect 11860 4281 11894 4315
rect 11860 4202 11894 4236
rect 11860 4123 11894 4157
rect 12565 4757 12599 4791
rect 12565 4677 12599 4711
rect 12565 4597 12599 4631
rect 12565 4518 12599 4552
rect 12565 4439 12599 4473
rect 12565 4360 12599 4394
rect 12565 4281 12599 4315
rect 12565 4202 12599 4236
rect 12565 4123 12599 4157
rect 12675 4778 12709 4810
rect 12675 4776 12709 4778
rect 12675 4710 12709 4736
rect 12675 4702 12709 4710
rect 12675 4642 12709 4662
rect 12675 4628 12709 4642
rect 12675 4574 12709 4588
rect 12675 4554 12709 4574
rect 12675 4506 12709 4514
rect 12675 4480 12709 4506
rect 12675 4438 12709 4440
rect 12675 4406 12709 4438
rect 12675 4331 12709 4365
rect 12675 4256 12709 4290
rect 12675 4181 12709 4215
rect 12675 4106 12709 4140
rect 11130 3696 11164 3698
rect 11130 3664 11164 3696
rect 11130 3594 11164 3626
rect 11130 3592 11164 3594
rect 11130 3440 11164 3442
rect 11130 3408 11164 3440
rect 11130 3338 11164 3370
rect 11130 3336 11164 3338
rect 10620 3244 10654 3278
rect 10692 3244 10726 3278
rect 10764 3244 10798 3278
rect 10836 3244 10870 3278
rect 10908 3244 10942 3278
rect 10980 3244 11014 3278
rect 11052 3244 11086 3278
rect 12675 4031 12709 4065
rect 12675 3956 12709 3990
rect 12675 3881 12709 3915
rect 12592 3824 12626 3829
rect 12592 3795 12624 3824
rect 12624 3795 12626 3824
rect 12592 3722 12624 3756
rect 12624 3722 12626 3756
rect 12675 3636 12709 3670
rect 12675 3556 12709 3590
rect 11860 3440 11894 3442
rect 11860 3408 11894 3440
rect 11860 3338 11894 3370
rect 11860 3336 11894 3338
rect 12590 3440 12624 3442
rect 12590 3408 12624 3440
rect 12590 3338 12624 3370
rect 12590 3336 12624 3338
rect 12008 3244 12042 3278
rect 12080 3244 12114 3278
rect 12152 3244 12186 3278
rect 12224 3244 12258 3278
rect 12296 3244 12330 3278
rect 12368 3244 12402 3278
rect 11046 3066 11080 3100
rect 11118 3082 11130 3100
rect 11130 3082 11152 3100
rect 11118 3066 11152 3082
rect 11776 3066 11810 3100
rect 11848 3082 11860 3100
rect 11860 3082 11882 3100
rect 11848 3066 11882 3082
rect 10400 3024 10434 3058
rect 10400 2952 10434 2986
rect 11046 2910 11080 2944
rect 11118 2928 11152 2944
rect 11118 2910 11130 2928
rect 11130 2910 11152 2928
rect 11776 2910 11810 2944
rect 11848 2928 11882 2944
rect 11848 2910 11860 2928
rect 11860 2910 11882 2928
rect 10620 2732 10654 2766
rect 10692 2732 10726 2766
rect 10764 2732 10798 2766
rect 10836 2732 10870 2766
rect 10908 2732 10942 2766
rect 10980 2732 11014 2766
rect 11052 2732 11086 2766
rect 12590 3184 12624 3186
rect 12590 3152 12624 3184
rect 12590 3082 12624 3114
rect 12590 3080 12624 3082
rect 12590 2768 12624 2802
rect 12675 3476 12709 3510
rect 12675 3396 12709 3430
rect 12675 3316 12709 3350
rect 12675 3236 12709 3270
rect 12675 3156 12709 3190
rect 12675 3075 12709 3109
rect 12675 2994 12709 3028
rect 12008 2732 12042 2766
rect 12080 2732 12114 2766
rect 12152 2732 12186 2766
rect 12224 2732 12258 2766
rect 12296 2732 12330 2766
rect 12368 2732 12402 2766
rect 12440 2732 12474 2766
rect 11046 2554 11080 2588
rect 11118 2570 11130 2588
rect 11130 2570 11152 2588
rect 11118 2554 11152 2570
rect 11776 2554 11810 2588
rect 11848 2570 11860 2588
rect 11860 2570 11882 2588
rect 11848 2554 11882 2570
rect 10400 2512 10434 2546
rect 10400 2440 10434 2474
rect 11046 2398 11080 2432
rect 11118 2416 11152 2432
rect 11118 2398 11130 2416
rect 11130 2398 11152 2416
rect 11776 2398 11810 2432
rect 11848 2416 11882 2432
rect 11848 2398 11860 2416
rect 11860 2398 11882 2416
rect 10400 2243 10434 2277
rect 10620 2220 10654 2254
rect 10692 2220 10726 2254
rect 10764 2220 10798 2254
rect 10836 2220 10870 2254
rect 10908 2220 10942 2254
rect 10980 2220 11014 2254
rect 11052 2220 11086 2254
rect 10400 2171 10434 2205
rect 10400 1904 10434 1906
rect 10400 1872 10434 1904
rect 10400 1802 10434 1834
rect 10400 1800 10434 1802
rect 12590 2696 12624 2730
rect 12008 2220 12042 2254
rect 12080 2220 12114 2254
rect 12152 2220 12186 2254
rect 12224 2220 12258 2254
rect 12296 2220 12330 2254
rect 12368 2220 12402 2254
rect 12670 2755 12704 2789
rect 12670 2672 12704 2706
rect 12670 2588 12704 2622
rect 12670 2504 12704 2538
rect 12675 2215 12709 2249
rect 12675 2140 12709 2174
rect 12675 2065 12709 2099
rect 11130 1904 11164 1906
rect 11130 1872 11164 1904
rect 11130 1802 11164 1834
rect 11130 1800 11164 1802
rect 10620 1708 10654 1742
rect 10692 1708 10726 1742
rect 10764 1708 10798 1742
rect 10836 1708 10870 1742
rect 10908 1708 10942 1742
rect 10980 1708 11014 1742
rect 11052 1708 11086 1742
rect 10400 1648 10434 1650
rect 10400 1616 10434 1648
rect 10400 1546 10434 1578
rect 10400 1544 10434 1546
rect 11130 1648 11164 1650
rect 11130 1616 11164 1648
rect 11130 1546 11164 1578
rect 11130 1544 11164 1546
rect 10423 1341 10457 1375
rect 10423 1261 10457 1295
rect 10423 1181 10457 1215
rect 10423 1102 10457 1136
rect 10423 1023 10457 1057
rect 10423 944 10457 978
rect 10423 865 10457 899
rect 10423 786 10457 820
rect 10423 707 10457 741
rect 11130 1341 11164 1375
rect 11130 1261 11164 1295
rect 11130 1181 11164 1215
rect 11130 1102 11164 1136
rect 11130 1023 11164 1057
rect 11130 944 11164 978
rect 11130 865 11164 899
rect 11130 786 11164 820
rect 11130 707 11164 741
rect 9468 608 9502 617
rect 9468 583 9502 608
rect 9706 570 9708 604
rect 9708 570 9740 604
rect 9778 570 9810 604
rect 9810 570 9812 604
rect 9942 571 9944 605
rect 9944 571 9976 605
rect 10014 571 10046 605
rect 10046 571 10048 605
rect 12675 1990 12709 2024
rect 12590 1904 12624 1906
rect 12590 1872 12624 1904
rect 12590 1802 12624 1834
rect 12590 1800 12624 1802
rect 12590 1648 12624 1650
rect 12590 1616 12624 1648
rect 12590 1546 12624 1578
rect 12590 1544 12624 1546
rect 12675 1915 12709 1949
rect 12675 1840 12709 1874
rect 12675 1765 12709 1799
rect 12675 1690 12709 1724
rect 12675 1615 12709 1649
rect 12675 1540 12709 1574
rect 12675 1465 12709 1499
rect 12675 1390 12709 1424
rect 11860 1341 11894 1375
rect 11860 1261 11894 1295
rect 11860 1181 11894 1215
rect 11860 1102 11894 1136
rect 11860 1023 11894 1057
rect 11860 944 11894 978
rect 11860 865 11894 899
rect 11860 786 11894 820
rect 11860 707 11894 741
rect 12565 1341 12599 1375
rect 12565 1261 12599 1295
rect 12565 1181 12599 1215
rect 12565 1102 12599 1136
rect 12565 1023 12599 1057
rect 12565 944 12599 978
rect 12565 865 12599 899
rect 12565 786 12599 820
rect 12565 707 12599 741
rect 12675 1315 12709 1349
rect 12675 1240 12709 1274
rect 12675 1165 12709 1199
rect 12675 1090 12709 1124
rect 12675 1015 12709 1049
rect 12675 940 12709 974
rect 12675 865 12709 899
rect 12675 791 12709 825
rect 12675 717 12709 751
rect 12675 643 12709 677
rect 9468 539 9502 544
rect 9468 510 9502 539
rect 12675 574 12709 603
rect 12675 569 12709 574
rect 9468 470 9502 471
rect 9468 437 9502 470
rect 11212 455 11214 489
rect 11214 455 11246 489
rect 11287 455 11316 489
rect 11316 455 11321 489
rect 11362 455 11384 489
rect 11384 455 11396 489
rect 11437 455 11452 489
rect 11452 455 11471 489
rect 11512 455 11520 489
rect 11520 455 11546 489
rect 11587 455 11588 489
rect 11588 455 11621 489
rect 11662 455 11690 489
rect 11690 455 11696 489
rect 11737 455 11758 489
rect 11758 455 11771 489
rect 11812 455 11826 489
rect 11826 455 11846 489
rect 11887 455 11894 489
rect 11894 455 11921 489
rect 11962 455 11996 489
rect 12037 455 12064 489
rect 12064 455 12071 489
rect 12112 455 12132 489
rect 12132 455 12146 489
rect 12187 455 12200 489
rect 12200 455 12221 489
rect 12262 455 12268 489
rect 12268 455 12296 489
rect 12337 455 12370 489
rect 12370 455 12371 489
rect 12412 455 12438 489
rect 12438 455 12446 489
rect 12487 455 12506 489
rect 12506 455 12521 489
rect 12562 455 12574 489
rect 12574 455 12596 489
rect 12637 455 12642 489
rect 12642 455 12671 489
rect 9468 367 9502 398
rect 9468 364 9502 367
rect 9468 298 9502 325
rect 9468 291 9502 298
rect 4844 243 4869 245
rect 4869 243 4878 245
rect 4844 211 4878 243
rect 4917 244 4951 245
rect 4990 244 5024 245
rect 5063 244 5097 245
rect 5136 244 5170 245
rect 5209 244 5243 245
rect 5282 244 5316 245
rect 5355 244 5389 245
rect 5428 244 5462 245
rect 5501 244 5535 245
rect 5574 244 5608 245
rect 5646 244 5680 245
rect 5718 244 5752 245
rect 5790 244 5824 245
rect 5862 244 5896 245
rect 5934 244 5968 245
rect 6006 244 6040 245
rect 6078 244 6112 245
rect 6150 244 6184 245
rect 6222 244 6256 245
rect 6294 244 6328 245
rect 6366 244 6400 245
rect 6438 244 6472 245
rect 6510 244 6544 245
rect 6582 244 6616 245
rect 6654 244 6688 245
rect 6726 244 6760 245
rect 6798 244 6832 245
rect 6870 244 6904 245
rect 6942 244 6976 245
rect 7014 244 7048 245
rect 7086 244 7120 245
rect 7158 244 7192 245
rect 7230 244 7264 245
rect 7302 244 7336 245
rect 7374 244 7408 245
rect 7446 244 7480 245
rect 7518 244 7552 245
rect 7590 244 7624 245
rect 7662 244 7696 245
rect 7734 244 7768 245
rect 7806 244 7840 245
rect 7878 244 7912 245
rect 7950 244 7984 245
rect 8022 244 8056 245
rect 8094 244 8128 245
rect 8166 244 8200 245
rect 8238 244 8272 245
rect 8310 244 8344 245
rect 8382 244 8416 245
rect 8454 244 8488 245
rect 8526 244 8560 245
rect 8598 244 8632 245
rect 8670 244 8704 245
rect 8742 244 8776 245
rect 8814 244 8848 245
rect 8886 244 8920 245
rect 8958 244 8992 245
rect 9030 244 9064 245
rect 9102 244 9136 245
rect 9174 244 9208 245
rect 9246 244 9280 245
rect 9318 244 9352 245
rect 9390 244 9424 245
rect 9462 244 9496 245
rect 4917 211 4947 244
rect 4947 211 4951 244
rect 4990 211 5015 244
rect 5015 211 5024 244
rect 5063 211 5083 244
rect 5083 211 5097 244
rect 5136 211 5151 244
rect 5151 211 5170 244
rect 5209 211 5219 244
rect 5219 211 5243 244
rect 5282 211 5287 244
rect 5287 211 5316 244
rect 5355 211 5389 244
rect 5428 211 5457 244
rect 5457 211 5462 244
rect 5501 211 5525 244
rect 5525 211 5535 244
rect 5574 211 5593 244
rect 5593 211 5608 244
rect 5646 211 5661 244
rect 5661 211 5680 244
rect 5718 211 5729 244
rect 5729 211 5752 244
rect 5790 211 5797 244
rect 5797 211 5824 244
rect 5862 211 5865 244
rect 5865 211 5896 244
rect 5934 211 5967 244
rect 5967 211 5968 244
rect 6006 211 6035 244
rect 6035 211 6040 244
rect 6078 211 6103 244
rect 6103 211 6112 244
rect 6150 211 6171 244
rect 6171 211 6184 244
rect 6222 211 6239 244
rect 6239 211 6256 244
rect 6294 211 6307 244
rect 6307 211 6328 244
rect 6366 211 6375 244
rect 6375 211 6400 244
rect 6438 211 6443 244
rect 6443 211 6472 244
rect 6510 211 6511 244
rect 6511 211 6544 244
rect 6582 211 6613 244
rect 6613 211 6616 244
rect 6654 211 6681 244
rect 6681 211 6688 244
rect 6726 211 6749 244
rect 6749 211 6760 244
rect 6798 211 6817 244
rect 6817 211 6832 244
rect 6870 211 6885 244
rect 6885 211 6904 244
rect 6942 211 6953 244
rect 6953 211 6976 244
rect 7014 211 7021 244
rect 7021 211 7048 244
rect 7086 211 7089 244
rect 7089 211 7120 244
rect 7158 211 7191 244
rect 7191 211 7192 244
rect 7230 211 7259 244
rect 7259 211 7264 244
rect 7302 211 7327 244
rect 7327 211 7336 244
rect 7374 211 7395 244
rect 7395 211 7408 244
rect 7446 211 7463 244
rect 7463 211 7480 244
rect 7518 211 7531 244
rect 7531 211 7552 244
rect 7590 211 7599 244
rect 7599 211 7624 244
rect 7662 211 7667 244
rect 7667 211 7696 244
rect 7734 211 7735 244
rect 7735 211 7768 244
rect 7806 211 7837 244
rect 7837 211 7840 244
rect 7878 211 7905 244
rect 7905 211 7912 244
rect 7950 211 7973 244
rect 7973 211 7984 244
rect 8022 211 8041 244
rect 8041 211 8056 244
rect 8094 211 8109 244
rect 8109 211 8128 244
rect 8166 211 8177 244
rect 8177 211 8200 244
rect 8238 211 8245 244
rect 8245 211 8272 244
rect 8310 211 8313 244
rect 8313 211 8344 244
rect 8382 211 8415 244
rect 8415 211 8416 244
rect 8454 211 8483 244
rect 8483 211 8488 244
rect 8526 211 8551 244
rect 8551 211 8560 244
rect 8598 211 8619 244
rect 8619 211 8632 244
rect 8670 211 8687 244
rect 8687 211 8704 244
rect 8742 211 8755 244
rect 8755 211 8776 244
rect 8814 211 8823 244
rect 8823 211 8848 244
rect 8886 211 8891 244
rect 8891 211 8920 244
rect 8958 211 8959 244
rect 8959 211 8992 244
rect 9030 211 9061 244
rect 9061 211 9064 244
rect 9102 211 9129 244
rect 9129 211 9136 244
rect 9174 211 9197 244
rect 9197 211 9208 244
rect 9246 211 9265 244
rect 9265 211 9280 244
rect 9318 211 9333 244
rect 9333 211 9352 244
rect 9390 211 9401 244
rect 9401 211 9424 244
rect 9462 211 9469 244
rect 9469 211 9496 244
rect 9650 247 9657 281
rect 9657 247 9684 281
rect 9722 276 9725 281
rect 9725 276 9756 281
rect 9722 247 9756 276
rect 10090 276 10099 281
rect 10099 276 10124 281
rect 10090 247 10124 276
rect 10162 247 10167 281
rect 10167 247 10196 281
rect 10467 247 10501 281
rect 10539 247 10573 281
rect 10893 247 10927 281
rect 10965 247 10999 281
rect 11300 280 11334 314
rect 11300 208 11334 242
rect 11846 233 11880 267
rect 11925 233 11959 267
rect 12004 233 12038 267
rect 12082 233 12116 267
rect 12574 310 12608 314
rect 12574 280 12604 310
rect 12604 280 12608 310
rect 12574 208 12604 242
rect 12604 208 12608 242
rect 8307 -28 8341 -8
rect 8379 -28 8413 -8
rect 8307 -42 8341 -28
rect 8379 -42 8409 -28
rect 8409 -42 8413 -28
rect 12574 -62 12608 -28
rect 10789 -126 10791 -92
rect 10791 -126 10823 -92
rect 10861 -126 10893 -92
rect 10893 -126 10895 -92
rect 12574 -130 12608 -100
rect 12574 -134 12608 -130
rect 6508 -206 6542 -172
rect 6580 -206 6614 -172
<< metal1 >>
rect 15265 13446 15325 13492
rect 10102 13224 10154 13230
tri 2379 13194 2391 13206 se
tri 2511 13194 2523 13206 sw
rect 2379 13188 2431 13194
rect 2379 13124 2431 13136
rect 2379 13066 2431 13072
rect 2471 13188 2523 13194
tri 10068 13150 10102 13184 ne
rect 10102 13160 10154 13172
rect 2471 13124 2523 13136
tri 10154 13150 10188 13184 nw
rect 10102 13102 10154 13108
rect 2471 13066 2523 13072
rect 6152 13067 9999 13073
rect 6204 13033 6281 13067
rect 6315 13033 6353 13067
rect 6387 13033 6425 13067
rect 6459 13033 6497 13067
rect 6531 13033 6569 13067
rect 6603 13033 6641 13067
rect 6675 13033 6713 13067
rect 6747 13033 6785 13067
rect 6819 13033 6857 13067
rect 6891 13033 6929 13067
rect 6963 13033 7001 13067
rect 7035 13033 7073 13067
rect 7107 13033 7145 13067
rect 7179 13033 7217 13067
rect 7251 13033 7289 13067
rect 7323 13033 7361 13067
rect 7395 13033 7433 13067
rect 7467 13033 7505 13067
rect 7539 13033 7577 13067
rect 7611 13033 7649 13067
rect 7683 13033 7721 13067
rect 7755 13033 7793 13067
rect 7827 13033 7865 13067
rect 7899 13033 7937 13067
rect 7971 13033 8009 13067
rect 8043 13033 8081 13067
rect 8115 13033 8153 13067
rect 8187 13033 8225 13067
rect 8259 13033 8297 13067
rect 8331 13033 8369 13067
rect 8403 13033 8441 13067
rect 8475 13033 8513 13067
rect 8547 13033 8585 13067
rect 8619 13033 8657 13067
rect 8691 13033 8729 13067
rect 8763 13033 8801 13067
rect 8835 13033 8873 13067
rect 8907 13033 8945 13067
rect 8979 13033 9017 13067
rect 9051 13033 9089 13067
rect 9123 13033 9161 13067
rect 9195 13033 9233 13067
rect 9267 13033 9305 13067
rect 9339 13033 9377 13067
rect 9411 13033 9449 13067
rect 9483 13033 9521 13067
rect 9555 13033 9593 13067
rect 9627 13033 9665 13067
rect 9699 13033 9737 13067
rect 9771 13033 9809 13067
rect 9843 13033 9881 13067
rect 9915 13033 9953 13067
rect 9987 13033 9999 13067
rect 6204 13027 9999 13033
rect 212 12980 272 13026
rect 6152 13001 6204 13015
rect 6152 12935 6204 12949
tri 6204 12940 6291 13027 nw
rect 6152 12869 6204 12883
rect 6152 12811 6161 12817
rect 6195 12811 6204 12817
rect 6152 12803 6204 12811
rect 6152 12739 6161 12751
rect 6195 12739 6204 12751
rect 6152 12737 6204 12739
rect 6152 12671 6161 12685
rect 6195 12671 6204 12685
rect 6152 12605 6161 12619
rect 6195 12605 6204 12619
rect 6152 12539 6161 12553
rect 6195 12539 6204 12553
rect 6152 12485 6204 12487
rect 6152 12473 6161 12485
rect 6195 12473 6204 12485
rect 6152 12413 6204 12421
rect 6152 12407 6161 12413
rect 6195 12407 6204 12413
rect 6152 12341 6204 12355
rect 6152 12275 6204 12289
rect 6152 12209 6204 12223
rect 6152 12143 6204 12157
rect 6152 12077 6204 12091
rect 6152 12019 6161 12025
rect 6195 12019 6204 12025
rect 6152 12011 6204 12019
rect 6152 11947 6161 11959
rect 6195 11947 6204 11959
rect 6152 11945 6204 11947
rect 6152 11879 6161 11893
rect 6195 11879 6204 11893
rect 6152 11813 6161 11827
rect 6195 11813 6204 11827
rect 6152 11747 6161 11761
rect 6195 11747 6204 11761
rect 6152 11693 6204 11695
rect 2471 11679 2523 11685
rect 6152 11681 6161 11693
rect 6195 11681 6204 11693
rect 2471 11621 2523 11627
tri 2523 11621 2541 11639 sw
rect 6152 11621 6204 11629
rect 2471 11615 2541 11621
rect 2523 11603 2541 11615
tri 2541 11603 2559 11621 sw
rect 6152 11615 6161 11621
rect 6195 11615 6204 11621
rect 2523 11595 3385 11603
tri 3385 11595 3393 11603 sw
rect 2523 11587 3393 11595
tri 3393 11587 3401 11595 sw
rect 2523 11563 3401 11587
rect 2471 11557 3401 11563
tri 3365 11549 3373 11557 ne
rect 3373 11549 3401 11557
tri 3401 11549 3439 11587 sw
tri 3373 11529 3393 11549 ne
rect 3393 11529 3439 11549
tri 3439 11529 3459 11549 sw
tri 3393 11515 3407 11529 ne
rect 3407 11515 3459 11529
tri 3459 11515 3473 11529 sw
tri 3407 11477 3445 11515 ne
rect 3445 11477 3473 11515
tri 3473 11477 3511 11515 sw
tri 3445 11463 3459 11477 ne
rect 3459 11463 3511 11477
tri 3511 11463 3525 11477 sw
tri 3459 11448 3474 11463 ne
rect 3474 11448 3525 11463
rect 5786 11457 5878 11563
rect 6152 11549 6204 11563
rect 6152 11483 6204 11497
rect 1673 11172 3305 11448
tri 3474 11443 3479 11448 ne
tri 3471 11138 3479 11146 se
rect 3479 11138 3525 11448
rect 6152 11417 6204 11431
rect 6152 11351 6204 11365
rect 6152 11285 6204 11299
rect 10220 11319 11266 11325
rect 11318 11319 11330 11325
rect 11382 11319 11861 11325
tri 6204 11285 6211 11292 sw
rect 10220 11285 10232 11319
rect 10266 11285 10308 11319
rect 10342 11285 10384 11319
rect 10418 11285 10460 11319
rect 10494 11285 10536 11319
rect 10570 11285 10612 11319
rect 10646 11285 10688 11319
rect 10722 11285 10764 11319
rect 10798 11285 10840 11319
rect 10874 11285 10915 11319
rect 10949 11285 10990 11319
rect 11024 11285 11065 11319
rect 11099 11285 11140 11319
rect 11174 11285 11215 11319
rect 11249 11285 11266 11319
rect 11324 11285 11330 11319
rect 11399 11285 11440 11319
rect 11474 11285 11515 11319
rect 11549 11285 11590 11319
rect 11624 11285 11665 11319
rect 11699 11285 11740 11319
rect 11774 11285 11815 11319
rect 11849 11285 11861 11319
rect 6152 11284 6211 11285
rect 6204 11232 6211 11284
rect 6152 11217 6211 11232
rect 6204 11205 6211 11217
tri 6211 11205 6291 11285 sw
rect 10220 11279 11266 11285
tri 11254 11273 11260 11279 ne
rect 11260 11273 11266 11279
rect 11318 11273 11330 11285
rect 11382 11279 11861 11285
rect 11382 11273 11388 11279
tri 11388 11273 11394 11279 nw
rect 6204 11199 8304 11205
rect 6204 11165 6239 11199
rect 6273 11165 6311 11199
rect 6345 11165 6383 11199
rect 6417 11165 6455 11199
rect 6489 11165 6527 11199
rect 6561 11165 6599 11199
rect 6633 11165 6671 11199
rect 6705 11165 6743 11199
rect 6777 11165 6815 11199
rect 6849 11165 6887 11199
rect 6921 11165 6959 11199
rect 6993 11165 7031 11199
rect 7065 11165 7103 11199
rect 7137 11165 7175 11199
rect 7209 11165 7247 11199
rect 7281 11165 7319 11199
rect 7353 11165 7391 11199
rect 7425 11165 7463 11199
rect 7497 11165 7535 11199
rect 7569 11165 7607 11199
rect 7641 11165 7679 11199
rect 7713 11165 7751 11199
rect 7785 11165 7823 11199
rect 7857 11165 7895 11199
rect 7929 11165 7967 11199
rect 8001 11165 8039 11199
rect 8073 11165 8111 11199
rect 8145 11165 8183 11199
rect 8217 11165 8255 11199
rect 8289 11165 8304 11199
rect 6152 11159 8304 11165
rect 2149 11126 2195 11138
tri 2195 11126 2207 11138 sw
tri 3459 11126 3471 11138 se
rect 3471 11126 3525 11138
rect 2149 11113 2207 11126
tri 2207 11113 2220 11126 sw
tri 3446 11113 3459 11126 se
rect 3459 11113 3512 11126
tri 3512 11113 3525 11126 nw
rect 2149 11110 2220 11113
tri 2220 11110 2223 11113 sw
tri 2274 11110 2277 11113 se
rect 2277 11110 2350 11113
rect 2149 11070 2350 11110
rect 2149 11036 2155 11070
rect 2189 11061 2350 11070
rect 2402 11061 2414 11113
rect 2466 11103 2635 11113
tri 3443 11110 3446 11113 se
rect 3446 11110 3509 11113
tri 3509 11110 3512 11113 nw
rect 2466 11069 2496 11103
rect 2530 11069 2589 11103
rect 2623 11069 2635 11103
tri 3423 11090 3443 11110 se
rect 3443 11090 3489 11110
tri 3489 11090 3509 11110 nw
tri 3403 11070 3423 11090 se
rect 2466 11061 2635 11069
rect 2189 11036 2195 11061
rect 2149 11024 2195 11036
tri 2195 11027 2229 11061 nw
rect 3129 11024 3423 11070
tri 3423 11024 3489 11090 nw
rect 7058 11017 7508 11020
rect 1673 10720 3305 10996
rect 7058 10965 7068 11017
rect 7120 10965 7144 11017
rect 7196 10965 7220 11017
rect 7272 10965 7296 11017
rect 7348 10965 7372 11017
rect 7424 10965 7447 11017
rect 7499 10965 7508 11017
tri 10109 10996 10128 11015 ne
rect 10128 10996 10143 11015
tri 10128 10981 10143 10996 ne
rect 7058 10953 7508 10965
rect 7058 10901 7068 10953
rect 7120 10901 7144 10953
rect 7196 10901 7220 10953
rect 7272 10901 7296 10953
rect 7348 10901 7372 10953
rect 7424 10901 7447 10953
rect 7499 10901 7508 10953
rect 7058 10896 7508 10901
tri 15237 10774 15240 10777 ne
rect 5587 10701 11489 10753
rect 326 10672 378 10678
rect 326 10608 378 10620
rect 326 10548 378 10556
tri 15206 10494 15240 10528 se
rect 6487 10437 11266 10443
rect 11318 10437 11330 10443
rect 11382 10437 11564 10443
rect 6487 10403 6499 10437
rect 6533 10403 6572 10437
rect 6606 10403 6645 10437
rect 6679 10403 6718 10437
rect 6752 10403 6791 10437
rect 6825 10403 6864 10437
rect 6898 10403 6937 10437
rect 6971 10403 7010 10437
rect 7044 10403 7083 10437
rect 7117 10403 7156 10437
rect 7190 10403 7229 10437
rect 7263 10403 7302 10437
rect 7336 10403 7375 10437
rect 7409 10403 7448 10437
rect 7482 10403 7521 10437
rect 7555 10403 7594 10437
rect 7628 10403 7667 10437
rect 7701 10403 7740 10437
rect 7774 10403 7813 10437
rect 7847 10403 7886 10437
rect 7920 10403 7959 10437
rect 7993 10403 8032 10437
rect 8066 10403 8105 10437
rect 8139 10403 8178 10437
rect 8212 10403 8251 10437
rect 8285 10403 8324 10437
rect 8358 10403 8397 10437
rect 8431 10403 8470 10437
rect 8504 10403 8543 10437
rect 8577 10403 8616 10437
rect 8650 10403 8689 10437
rect 8723 10403 8762 10437
rect 8796 10403 8835 10437
rect 8869 10403 8908 10437
rect 8942 10403 8981 10437
rect 9015 10403 9054 10437
rect 9088 10403 9127 10437
rect 9161 10403 9200 10437
rect 9234 10403 9273 10437
rect 9307 10403 9346 10437
rect 9380 10403 9419 10437
rect 9453 10403 9492 10437
rect 9526 10403 9565 10437
rect 9599 10403 9638 10437
rect 9672 10403 9711 10437
rect 9745 10403 9784 10437
rect 9818 10403 9857 10437
rect 9891 10403 9930 10437
rect 9964 10403 10003 10437
rect 10037 10403 10076 10437
rect 10110 10403 10149 10437
rect 10183 10403 10222 10437
rect 10256 10403 10294 10437
rect 10328 10403 10366 10437
rect 10400 10403 10438 10437
rect 10472 10403 10510 10437
rect 10544 10403 10582 10437
rect 10616 10403 10654 10437
rect 10688 10403 10726 10437
rect 10760 10403 10798 10437
rect 10832 10403 10870 10437
rect 10904 10403 10942 10437
rect 10976 10403 11014 10437
rect 11048 10403 11086 10437
rect 11120 10403 11158 10437
rect 11192 10403 11230 10437
rect 11264 10403 11266 10437
rect 11408 10403 11446 10437
rect 11480 10403 11518 10437
rect 11552 10403 11564 10437
rect 6487 10397 11266 10403
tri 11254 10391 11260 10397 ne
rect 11260 10391 11266 10397
rect 11318 10391 11330 10403
rect 11382 10397 11564 10403
rect 11382 10391 11388 10397
tri 11388 10391 11394 10397 nw
rect 15240 10378 15446 10777
tri 15446 10494 15480 10528 sw
rect 7063 10132 7506 10148
rect 7063 10080 7067 10132
rect 7119 10080 7131 10132
rect 7183 10080 7195 10132
rect 7247 10080 7259 10098
rect 7311 10080 7323 10132
rect 7439 10098 7444 10132
rect 7375 10080 7387 10098
rect 7439 10080 7451 10098
rect 7503 10080 7506 10132
rect 7063 10065 7506 10080
rect 7063 10013 7067 10065
rect 7119 10013 7131 10065
rect 7183 10013 7195 10065
rect 7247 10051 7259 10065
rect 7247 10013 7259 10017
rect 7311 10013 7323 10065
rect 7375 10051 7387 10065
rect 7439 10051 7451 10065
rect 7439 10017 7444 10051
rect 7375 10013 7387 10017
rect 7439 10013 7451 10017
rect 7503 10013 7506 10065
rect 7063 9998 7506 10013
rect 7063 9946 7067 9998
rect 7119 9946 7131 9998
rect 7183 9946 7195 9998
rect 7247 9970 7259 9998
rect 7311 9946 7323 9998
rect 7375 9970 7387 9998
rect 7439 9970 7451 9998
rect 7439 9946 7444 9970
rect 7503 9946 7506 9998
rect 7063 9936 7069 9946
rect 7103 9936 7147 9946
rect 7181 9936 7225 9946
rect 7259 9936 7372 9946
rect 7406 9936 7444 9946
rect 7478 9936 7506 9946
rect 7063 9930 7506 9936
rect 7063 9878 7067 9930
rect 7119 9878 7131 9930
rect 7183 9878 7195 9930
rect 7247 9889 7259 9930
rect 7311 9878 7323 9930
rect 7375 9889 7387 9930
rect 7439 9889 7451 9930
rect 7439 9878 7444 9889
rect 7503 9878 7506 9930
rect 7063 9862 7069 9878
rect 7103 9862 7147 9878
rect 7181 9862 7225 9878
rect 7259 9862 7372 9878
rect 7406 9862 7444 9878
rect 7478 9862 7506 9878
rect 7063 9810 7067 9862
rect 7119 9810 7131 9862
rect 7183 9810 7195 9862
rect 7247 9810 7259 9855
rect 7311 9810 7323 9862
rect 7439 9855 7444 9862
rect 7375 9810 7387 9855
rect 7439 9810 7451 9855
rect 7503 9810 7506 9862
rect 7063 9807 7506 9810
rect 7063 9794 7069 9807
rect 7103 9794 7147 9807
rect 7181 9794 7225 9807
rect 7259 9794 7372 9807
rect 7406 9794 7444 9807
rect 7478 9794 7506 9807
rect 7063 9742 7067 9794
rect 7119 9742 7131 9794
rect 7183 9742 7195 9794
rect 7247 9742 7259 9773
rect 7311 9742 7323 9794
rect 7439 9773 7444 9794
rect 7375 9742 7387 9773
rect 7439 9742 7451 9773
rect 7503 9742 7506 9794
rect 7063 9726 7506 9742
rect 7063 9674 7067 9726
rect 7119 9674 7131 9726
rect 7183 9674 7195 9726
rect 7247 9725 7259 9726
rect 7247 9674 7259 9691
rect 7311 9674 7323 9726
rect 7375 9725 7387 9726
rect 7439 9725 7451 9726
rect 7439 9691 7444 9725
rect 7375 9674 7387 9691
rect 7439 9674 7451 9691
rect 7503 9674 7506 9726
rect 7063 9658 7506 9674
rect 7063 9606 7067 9658
rect 7119 9606 7131 9658
rect 7183 9606 7195 9658
rect 7247 9643 7259 9658
rect 7247 9606 7259 9609
rect 7311 9606 7323 9658
rect 7375 9643 7387 9658
rect 7439 9643 7451 9658
rect 7439 9609 7444 9643
rect 7375 9606 7387 9609
rect 7439 9606 7451 9609
rect 7503 9606 7506 9658
rect 7063 9586 7506 9606
tri 10292 9559 10299 9566 se
rect 10299 9559 10453 9566
tri 10453 9559 10460 9566 sw
tri 10286 9553 10292 9559 se
rect 10292 9553 10331 9559
rect 6487 9547 10331 9553
rect 6487 9513 6499 9547
rect 6533 9513 6573 9547
rect 6607 9513 6647 9547
rect 6681 9513 6721 9547
rect 6755 9513 6795 9547
rect 6829 9513 6869 9547
rect 6903 9513 6943 9547
rect 6977 9513 7017 9547
rect 7051 9513 7091 9547
rect 7125 9513 7165 9547
rect 7199 9513 7239 9547
rect 7273 9513 7313 9547
rect 7347 9513 7387 9547
rect 7421 9513 7461 9547
rect 7495 9513 7535 9547
rect 7569 9513 7609 9547
rect 7643 9513 7683 9547
rect 7717 9513 7757 9547
rect 7791 9513 7831 9547
rect 7865 9513 7905 9547
rect 7939 9513 7979 9547
rect 8013 9513 8053 9547
rect 8087 9513 8127 9547
rect 8161 9513 8201 9547
rect 8235 9513 8275 9547
rect 8309 9513 8349 9547
rect 8383 9513 8423 9547
rect 8457 9513 8496 9547
rect 8530 9513 8569 9547
rect 8603 9513 8642 9547
rect 8676 9513 8715 9547
rect 8749 9513 8788 9547
rect 8822 9513 8861 9547
rect 8895 9513 8934 9547
rect 8968 9513 9007 9547
rect 9041 9513 9080 9547
rect 9114 9513 9153 9547
rect 9187 9513 9226 9547
rect 9260 9513 9299 9547
rect 9333 9513 9372 9547
rect 9406 9513 9445 9547
rect 9479 9513 9518 9547
rect 9552 9513 9591 9547
rect 9625 9513 9664 9547
rect 9698 9513 9737 9547
rect 9771 9513 9810 9547
rect 9844 9513 10331 9547
rect 6487 9507 10331 9513
rect 10383 9507 10395 9559
rect 10447 9553 10460 9559
tri 10460 9553 10466 9559 sw
tri 11254 9553 11260 9559 se
rect 11260 9553 11266 9559
rect 10447 9507 11266 9553
rect 11318 9507 11330 9559
rect 11382 9553 11388 9559
tri 11388 9553 11394 9559 sw
rect 11382 9514 12197 9553
tri 12197 9514 12236 9553 sw
rect 11382 9507 12236 9514
tri 12134 9462 12179 9507 ne
rect 7063 9402 7506 9418
rect 7063 9350 7067 9402
rect 7119 9350 7131 9402
rect 7183 9350 7195 9402
rect 7247 9350 7259 9368
rect 7311 9350 7323 9402
rect 7439 9368 7444 9402
rect 7375 9350 7387 9368
rect 7439 9350 7451 9368
rect 7503 9350 7506 9402
rect 7063 9335 7506 9350
rect 7063 9283 7067 9335
rect 7119 9283 7131 9335
rect 7183 9283 7195 9335
rect 7247 9321 7259 9335
rect 7247 9283 7259 9287
rect 7311 9283 7323 9335
rect 7375 9321 7387 9335
rect 7439 9321 7451 9335
rect 7439 9287 7444 9321
rect 7375 9283 7387 9287
rect 7439 9283 7451 9287
rect 7503 9283 7506 9335
rect 7063 9268 7506 9283
rect 7063 9216 7067 9268
rect 7119 9216 7131 9268
rect 7183 9216 7195 9268
rect 7247 9240 7259 9268
rect 7311 9216 7323 9268
rect 7375 9240 7387 9268
rect 7439 9240 7451 9268
rect 7439 9216 7444 9240
rect 7503 9216 7506 9268
rect 7063 9206 7069 9216
rect 7103 9206 7147 9216
rect 7181 9206 7225 9216
rect 7259 9206 7372 9216
rect 7406 9206 7444 9216
rect 7478 9206 7506 9216
rect 7063 9200 7506 9206
rect 7063 9148 7067 9200
rect 7119 9148 7131 9200
rect 7183 9148 7195 9200
rect 7247 9159 7259 9200
rect 7311 9148 7323 9200
rect 7375 9159 7387 9200
rect 7439 9159 7451 9200
rect 7439 9148 7444 9159
rect 7503 9148 7506 9200
rect 7063 9132 7069 9148
rect 7103 9132 7147 9148
rect 7181 9132 7225 9148
rect 7259 9132 7372 9148
rect 7406 9132 7444 9148
rect 7478 9132 7506 9148
rect 7063 9080 7067 9132
rect 7119 9080 7131 9132
rect 7183 9080 7195 9132
rect 7247 9080 7259 9125
rect 7311 9080 7323 9132
rect 7439 9125 7444 9132
rect 7375 9080 7387 9125
rect 7439 9080 7451 9125
rect 7503 9080 7506 9132
rect 7063 9077 7506 9080
rect 7063 9064 7069 9077
rect 7103 9064 7147 9077
rect 7181 9064 7225 9077
rect 7259 9064 7372 9077
rect 7406 9064 7444 9077
rect 7478 9064 7506 9077
rect 7063 9012 7067 9064
rect 7119 9012 7131 9064
rect 7183 9012 7195 9064
rect 7247 9012 7259 9043
rect 7311 9012 7323 9064
rect 7439 9043 7444 9064
rect 7375 9012 7387 9043
rect 7439 9012 7451 9043
rect 7503 9012 7506 9064
rect 7063 8996 7506 9012
rect 7063 8944 7067 8996
rect 7119 8944 7131 8996
rect 7183 8944 7195 8996
rect 7247 8995 7259 8996
rect 7247 8944 7259 8961
rect 7311 8944 7323 8996
rect 7375 8995 7387 8996
rect 7439 8995 7451 8996
rect 7439 8961 7444 8995
rect 7375 8944 7387 8961
rect 7439 8944 7451 8961
rect 7503 8944 7506 8996
rect 10715 8983 10775 9029
rect 7063 8928 7506 8944
rect 7063 8876 7067 8928
rect 7119 8876 7131 8928
rect 7183 8876 7195 8928
rect 7247 8913 7259 8928
rect 7247 8876 7259 8879
rect 7311 8876 7323 8928
rect 7375 8913 7387 8928
rect 7439 8913 7451 8928
rect 7439 8879 7444 8913
rect 7375 8876 7387 8879
rect 7439 8876 7451 8879
rect 7503 8876 7506 8928
rect 7063 8856 7506 8876
rect 9586 8742 9678 8788
tri 4813 8557 4825 8569 se
rect 4825 8517 4831 8569
rect 4883 8517 4895 8569
rect 4947 8517 4953 8569
tri 4953 8557 4965 8569 sw
rect 12179 8329 12236 9507
tri 12179 8325 12183 8329 ne
rect 12183 8325 12236 8329
tri 12236 8325 12270 8359 sw
tri 12183 8320 12188 8325 ne
rect 12188 8320 12462 8325
tri 12462 8320 12467 8325 sw
tri 12646 8320 12651 8325 se
rect 12651 8320 13697 8325
tri 12188 8279 12229 8320 ne
rect 12229 8279 13697 8320
tri 13685 8273 13691 8279 ne
rect 13691 8273 13697 8279
rect 13749 8273 13761 8325
rect 13813 8273 13819 8325
rect 147 7797 153 7849
rect 205 7797 217 7849
rect 269 7797 884 7849
rect 936 7797 948 7849
rect 1000 7797 1006 7849
tri 12988 7486 12991 7489 se
tri 12988 7437 12991 7440 ne
rect 13343 7437 13641 7489
rect 12643 7194 12649 7246
rect 12701 7194 12733 7246
rect 12785 7194 12818 7246
rect 12870 7194 12903 7246
rect 12955 7194 12961 7246
rect 12991 7194 12997 7246
rect 13049 7194 13069 7246
rect 13121 7194 13141 7246
rect 13193 7194 13213 7246
rect 13265 7194 13286 7246
rect 13338 7194 13344 7246
rect 2705 7051 2824 7122
tri 2824 7051 2895 7122 sw
rect 2705 6968 2895 7051
tri 2813 6886 2895 6968 ne
tri 2895 6907 3039 7051 sw
rect 2895 6886 3039 6907
tri 3039 6886 3060 6907 sw
tri 8726 6886 8747 6907 se
rect 8747 6886 13879 6907
tri 2895 6721 3060 6886 ne
tri 3060 6796 3150 6886 sw
tri 8636 6796 8726 6886 se
rect 8726 6796 13879 6886
rect 3060 6721 3150 6796
tri 3150 6721 3225 6796 sw
tri 3060 6690 3091 6721 ne
rect 3091 6690 3225 6721
tri 8530 6690 8636 6796 se
rect 8636 6791 8795 6796
tri 8795 6791 8800 6796 nw
tri 13868 6791 13873 6796 ne
rect 13873 6791 13879 6796
rect 13995 6791 14001 6907
rect 8636 6690 8694 6791
tri 8694 6690 8795 6791 nw
tri 14008 6753 14033 6778 se
rect 13767 6747 14033 6753
rect 13819 6695 14033 6747
tri 3091 6672 3109 6690 ne
rect 3109 6526 3225 6690
tri 8375 6535 8530 6690 se
tri 3225 6526 3234 6535 sw
tri 8366 6526 8375 6535 se
rect 8375 6526 8530 6535
tri 8530 6526 8694 6690 nw
rect 13767 6683 13819 6695
tri 13819 6645 13869 6695 nw
tri 14008 6670 14033 6695 ne
rect 13767 6625 13819 6631
rect 8847 6526 8899 6544
tri 8899 6526 8911 6538 sw
tri 10977 6526 10989 6538 se
rect 10989 6526 11217 6544
tri 11217 6526 11229 6538 sw
tri 13295 6526 13307 6538 se
rect 13307 6526 13359 6544
rect 3109 6487 3234 6526
tri 3234 6487 3273 6526 sw
tri 8327 6487 8366 6526 se
rect 8366 6487 8491 6526
tri 8491 6487 8530 6526 nw
rect 8847 6504 8911 6526
tri 8911 6504 8933 6526 sw
tri 10955 6504 10977 6526 se
rect 10977 6504 11229 6526
tri 11229 6504 11251 6526 sw
tri 13273 6504 13295 6526 se
rect 13295 6504 13359 6526
tri 3109 6362 3234 6487 ne
rect 3234 6478 3273 6487
tri 3273 6478 3282 6487 sw
tri 8318 6478 8327 6487 se
rect 8327 6478 8366 6487
rect 3234 6362 8366 6478
tri 8366 6362 8491 6487 nw
rect 8847 6458 13359 6504
rect 8847 6414 8899 6458
tri 8899 6424 8933 6458 nw
tri 10955 6424 10989 6458 ne
rect 10989 6414 11217 6458
tri 11217 6424 11251 6458 nw
tri 13273 6424 13307 6458 ne
rect 13307 6414 13359 6458
rect 2918 6340 2958 6341
tri 2958 6340 2959 6341 sw
rect 10960 6340 11276 6386
rect 2918 6316 2959 6340
tri 2959 6316 2983 6340 sw
rect 2918 6313 2983 6316
tri 2918 6308 2923 6313 ne
rect 2923 6308 2983 6313
tri 2923 6300 2931 6308 ne
rect 2931 6289 2983 6308
rect -87 6233 2712 6239
rect -35 6221 2712 6233
tri 2712 6221 2730 6239 sw
rect 2931 6221 2983 6237
rect 8847 6268 8899 6308
tri 8899 6268 8933 6302 sw
tri 10955 6268 10989 6302 se
rect 10989 6268 11217 6308
tri 11217 6268 11251 6302 sw
tri 13273 6268 13307 6302 se
rect 13307 6268 13359 6308
rect 8847 6222 13359 6268
rect 8847 6221 8932 6222
tri 8932 6221 8933 6222 nw
tri 10955 6221 10956 6222 ne
rect 10956 6221 11217 6222
rect -35 6189 2730 6221
tri 2730 6189 2762 6221 sw
rect -35 6187 2762 6189
rect -35 6181 1 6187
rect -87 6169 1 6181
rect -35 6147 1 6169
tri 1 6147 41 6187 nw
tri 2698 6159 2726 6187 ne
rect 2726 6159 2762 6187
rect 244 6153 296 6159
rect -35 6146 0 6147
tri 0 6146 1 6147 nw
rect -35 6117 -33 6146
rect -87 6113 -33 6117
tri -33 6113 0 6146 nw
rect 766 6153 818 6159
tri 2726 6156 2729 6159 ne
rect 2729 6156 2762 6159
rect -87 6111 -35 6113
tri -35 6111 -33 6113 nw
rect 244 6086 296 6101
rect 417 6094 445 6146
rect 497 6094 509 6146
rect 561 6094 573 6146
rect 625 6094 631 6146
rect 244 6019 250 6034
rect 284 6019 296 6034
rect 766 6073 818 6101
rect 958 6150 1010 6156
rect 1471 6150 1523 6156
rect 958 6068 1010 6098
rect 1150 6094 1156 6146
rect 1208 6094 1225 6146
rect 1277 6094 1294 6146
rect 1346 6094 1352 6146
tri 2729 6146 2739 6156 ne
rect 2739 6146 2762 6156
tri 2762 6146 2805 6189 sw
rect 2931 6163 2983 6169
rect 4637 6215 4689 6221
rect 8847 6178 8899 6221
tri 8899 6188 8932 6221 nw
tri 10956 6188 10989 6221 ne
rect 10989 6178 11217 6221
tri 11217 6188 11251 6222 nw
tri 13273 6188 13307 6222 ne
rect 13307 6178 13359 6222
rect 4637 6146 4689 6163
tri 2739 6123 2762 6146 ne
rect 2762 6123 2805 6146
tri 2805 6123 2828 6146 sw
rect 766 6015 818 6021
rect 878 6044 930 6050
rect 958 6010 1010 6016
rect 1471 6085 1523 6098
tri 2274 6094 2303 6123 se
rect 2303 6094 2705 6123
tri 2234 6054 2274 6094 se
rect 2274 6054 2705 6094
tri 2762 6077 2808 6123 ne
rect 2808 6117 3075 6123
rect 2808 6077 3023 6117
rect 1471 6020 1523 6033
tri 853 5967 878 5992 se
rect 878 5979 930 5992
rect 244 5952 250 5967
rect 284 5952 296 5967
rect 244 5887 296 5900
rect 244 5885 250 5887
rect 284 5885 296 5887
rect 244 5818 296 5833
rect 244 5751 296 5766
rect 244 5687 250 5699
rect 284 5687 296 5699
rect 244 5684 296 5687
rect 244 5617 250 5632
rect 284 5617 296 5632
rect 244 5555 296 5565
rect 244 5550 250 5555
rect 284 5550 296 5555
rect 244 5484 296 5498
rect 244 5426 296 5432
rect 329 5921 463 5967
rect 619 5927 878 5967
tri 930 5967 955 5992 sw
rect 930 5927 1150 5967
rect 619 5921 1150 5927
rect 1471 5960 1480 5968
rect 1514 5960 1523 5968
rect 1471 5955 1523 5960
rect 329 5919 398 5921
tri 398 5919 400 5921 nw
rect 329 5631 375 5919
tri 375 5896 398 5919 nw
rect 687 5881 733 5893
rect 687 5847 693 5881
rect 727 5847 733 5881
rect 687 5809 733 5847
rect 417 5742 445 5794
rect 497 5742 509 5794
rect 561 5742 573 5794
rect 625 5742 631 5794
rect 687 5775 693 5809
rect 727 5775 733 5809
rect 687 5737 733 5775
rect 687 5703 693 5737
rect 727 5703 733 5737
rect 687 5665 733 5703
tri 375 5631 384 5640 sw
rect 687 5631 693 5665
rect 727 5631 733 5665
rect 769 5887 821 5893
rect 769 5795 821 5835
rect 769 5703 821 5743
rect 769 5645 821 5651
rect 958 5887 1010 5893
rect 958 5795 1010 5835
rect 958 5703 1010 5743
rect 958 5645 1010 5651
rect 1046 5881 1092 5893
rect 1046 5847 1052 5881
rect 1086 5847 1092 5881
rect 1046 5809 1092 5847
rect 1046 5775 1052 5809
rect 1086 5775 1092 5809
rect 1471 5890 1480 5903
rect 1514 5890 1523 5903
rect 1570 5887 2096 6054
rect 2132 5982 2705 6054
tri 2998 6052 3023 6077 ne
rect 3023 6049 3075 6065
rect 3023 5991 3075 5997
rect 10960 6104 11276 6150
rect 4637 6077 4689 6094
rect 4637 6008 4689 6025
rect 2132 5887 2610 5982
tri 2610 5887 2705 5982 nw
rect 4637 5939 4689 5956
rect 8847 6028 8899 6076
tri 8899 6028 8933 6062 sw
tri 10955 6028 10989 6062 se
rect 10989 6059 11217 6072
tri 11217 6059 11220 6062 sw
rect 10989 6028 11220 6059
tri 11220 6028 11251 6059 sw
tri 13273 6028 13304 6059 se
rect 13304 6028 13356 6072
rect 8847 5982 13356 6028
rect 8847 5946 8899 5982
tri 8899 5948 8933 5982 nw
tri 10955 5948 10989 5982 ne
rect 10989 5942 11217 5982
tri 11217 5948 11251 5982 nw
tri 13273 5951 13304 5982 ne
rect 13304 5942 13356 5982
rect 1471 5825 1480 5838
rect 1514 5825 1523 5838
rect 329 5615 384 5631
tri 384 5615 400 5631 sw
rect 687 5615 733 5631
tri 733 5615 758 5640 sw
tri 1021 5615 1046 5640 se
rect 1046 5615 1092 5775
rect 1150 5742 1156 5794
rect 1208 5742 1225 5794
rect 1277 5742 1294 5794
rect 1346 5742 1352 5794
rect 1471 5767 1523 5773
rect 1471 5759 1480 5767
rect 1514 5759 1523 5767
rect 1686 5763 1704 5887
tri 1704 5763 1828 5887 nw
rect 4637 5870 4689 5887
rect 10960 5868 11276 5914
rect 4637 5801 4689 5818
tri 1686 5745 1704 5763 nw
rect 1471 5693 1523 5707
rect 4637 5731 4689 5749
rect 8847 5791 8899 5836
tri 8899 5791 8933 5825 sw
tri 10955 5791 10989 5825 se
rect 10989 5791 11217 5836
tri 11217 5791 11251 5825 sw
tri 13273 5791 13307 5825 se
rect 13307 5791 13359 5836
rect 8847 5745 13359 5791
rect 8847 5706 8899 5745
tri 8899 5711 8933 5745 nw
tri 10955 5711 10989 5745 ne
rect 10989 5706 11217 5745
tri 11217 5711 11251 5745 nw
tri 13273 5711 13307 5745 ne
rect 13307 5706 13359 5745
rect 4637 5673 4689 5679
tri 1092 5615 1117 5640 sw
rect 1471 5627 1523 5641
rect 329 5569 463 5615
rect 687 5593 1150 5615
rect 329 5559 399 5569
tri 399 5559 409 5569 nw
rect 687 5559 693 5593
rect 727 5569 1150 5593
rect 3023 5656 3075 5662
rect 3023 5592 3075 5604
tri 2298 5580 2303 5585 se
rect 2303 5580 2705 5585
rect 1471 5569 1523 5575
tri 2292 5574 2298 5580 se
rect 2298 5574 2705 5580
tri 2287 5569 2292 5574 se
rect 2292 5569 2705 5574
rect 727 5559 733 5569
rect 329 5540 380 5559
tri 380 5540 399 5559 nw
rect 160 5402 212 5408
tri 318 5360 329 5371 se
rect 329 5360 375 5540
tri 375 5535 380 5540 nw
rect 687 5521 733 5559
tri 733 5544 758 5569 nw
tri 2262 5544 2287 5569 se
rect 2287 5544 2705 5569
tri 2259 5541 2262 5544 se
rect 2262 5541 2705 5544
rect 687 5487 693 5521
rect 727 5487 733 5521
rect 417 5390 445 5442
rect 497 5390 509 5442
rect 561 5390 573 5442
rect 625 5390 631 5442
tri 212 5357 215 5360 sw
tri 315 5357 318 5360 se
rect 318 5357 375 5360
tri 673 5357 687 5371 se
rect 687 5357 733 5487
rect 212 5355 215 5357
tri 215 5355 217 5357 sw
tri 313 5355 315 5357 se
rect 315 5355 375 5357
tri 671 5355 673 5357 se
rect 673 5355 733 5357
rect 212 5350 217 5355
rect 160 5338 217 5350
rect 212 5326 217 5338
tri 217 5326 246 5355 sw
tri 284 5326 313 5355 se
rect 313 5351 375 5355
rect 313 5326 350 5351
tri 350 5326 375 5351 nw
tri 642 5326 671 5355 se
rect 671 5351 733 5355
rect 671 5326 705 5351
rect 212 5323 347 5326
tri 347 5323 350 5326 nw
tri 639 5323 642 5326 se
rect 642 5323 705 5326
tri 705 5323 733 5351 nw
rect 769 5532 821 5538
rect 769 5467 821 5480
rect 769 5403 778 5415
rect 812 5403 821 5415
rect 769 5339 821 5351
rect 212 5315 339 5323
tri 339 5315 347 5323 nw
tri 631 5315 639 5323 se
rect 639 5315 697 5323
tri 697 5315 705 5323 nw
rect 212 5286 305 5315
rect 160 5281 305 5286
tri 305 5281 339 5315 nw
tri 621 5305 631 5315 se
rect 631 5305 687 5315
tri 687 5305 697 5315 nw
tri 597 5281 621 5305 se
rect 621 5281 663 5305
tri 663 5281 687 5305 nw
rect 769 5281 778 5287
rect 812 5281 821 5287
rect 160 5280 304 5281
tri 304 5280 305 5281 nw
tri 596 5280 597 5281 se
rect 597 5280 649 5281
tri 583 5267 596 5280 se
rect 596 5267 649 5280
tri 649 5267 663 5281 nw
rect 769 5275 821 5281
tri 579 5263 583 5267 se
rect 583 5263 645 5267
tri 645 5263 649 5267 nw
rect 619 5217 645 5263
rect 769 5217 821 5223
rect 870 5535 1603 5541
tri 2258 5540 2259 5541 se
rect 2259 5540 2705 5541
rect 870 5495 1043 5535
tri 845 5189 870 5214 se
rect 870 5189 912 5495
tri 912 5470 937 5495 nw
tri 1018 5470 1043 5495 ne
rect 1095 5495 1603 5535
tri 2252 5534 2258 5540 se
rect 2258 5534 2705 5540
tri 3075 5585 3152 5662 sw
rect 7927 5624 8019 5670
tri 11852 5585 11853 5586 se
rect 11853 5585 11859 5586
rect 3075 5580 3152 5585
tri 3152 5580 3157 5585 sw
tri 11847 5580 11852 5585 se
rect 11852 5580 11859 5585
rect 3075 5574 3157 5580
tri 3157 5574 3163 5580 sw
tri 11841 5574 11847 5580 se
rect 11847 5574 11859 5580
rect 3075 5570 3163 5574
tri 3163 5570 3167 5574 sw
tri 11837 5570 11841 5574 se
rect 11841 5570 11859 5574
rect 3075 5540 4611 5570
tri 4611 5540 4641 5570 sw
tri 8575 5540 8605 5570 se
rect 8605 5540 11859 5570
rect 3023 5539 4641 5540
tri 4641 5539 4642 5540 sw
tri 8574 5539 8575 5540 se
rect 8575 5539 11859 5540
rect 3023 5534 11859 5539
rect 11911 5534 11923 5586
rect 11975 5580 11981 5586
tri 11981 5580 11987 5586 sw
rect 11975 5574 11987 5580
tri 11987 5574 11993 5580 sw
tri 13722 5574 13728 5580 se
rect 13728 5574 13858 5580
rect 11975 5570 11993 5574
tri 11993 5570 11997 5574 sw
tri 13718 5570 13722 5574 se
rect 13722 5570 13740 5574
rect 11975 5540 13740 5570
rect 13774 5540 13812 5574
rect 13846 5540 13858 5574
rect 11975 5534 13858 5540
tri 2240 5522 2252 5534 se
rect 2252 5522 2705 5534
tri 4597 5522 4609 5534 ne
rect 4609 5522 8591 5534
tri 2234 5516 2240 5522 se
rect 2240 5516 2705 5522
rect 1043 5471 1095 5483
rect 0 5147 912 5189
rect 958 5453 1010 5459
tri 1095 5470 1120 5495 nw
tri 1532 5470 1557 5495 ne
tri 1188 5466 1189 5467 se
rect 1189 5466 1338 5467
tri 1183 5461 1188 5466 se
rect 1188 5461 1338 5466
tri 1149 5427 1183 5461 se
rect 1183 5427 1220 5461
rect 1254 5427 1292 5461
rect 1326 5427 1338 5461
tri 1143 5421 1149 5427 se
rect 1149 5421 1338 5427
rect 1471 5458 1523 5464
rect 1043 5413 1095 5419
tri 1139 5417 1143 5421 se
rect 1143 5417 1195 5421
tri 1195 5417 1199 5421 nw
tri 1135 5413 1139 5417 se
rect 1139 5413 1189 5417
tri 1133 5411 1135 5413 se
rect 1135 5411 1189 5413
tri 1189 5411 1195 5417 nw
rect 958 5382 1010 5401
tri 1112 5390 1133 5411 se
rect 1133 5390 1156 5411
tri 1100 5378 1112 5390 se
rect 1112 5378 1156 5390
tri 1156 5378 1189 5411 nw
rect 1471 5393 1523 5406
tri 1077 5355 1100 5378 se
rect 1100 5355 1133 5378
tri 1133 5355 1156 5378 nw
tri 1066 5344 1077 5355 se
rect 1077 5344 1122 5355
tri 1122 5344 1133 5355 nw
rect 958 5323 967 5330
rect 1001 5323 1010 5330
rect 958 5311 1010 5323
rect 958 5241 967 5259
rect 1001 5241 1010 5259
rect 958 5178 1010 5189
rect 958 5171 967 5178
rect 1001 5171 1010 5178
rect 329 5107 375 5119
rect 244 5101 296 5107
rect 244 5033 296 5049
rect 244 4965 296 4981
rect 244 4905 250 4913
rect 284 4905 296 4913
rect 244 4897 296 4905
rect 244 4829 250 4845
rect 284 4829 296 4845
rect 244 4761 250 4777
rect 284 4761 296 4777
rect 244 4703 296 4709
rect 244 4693 250 4703
rect 284 4693 296 4703
rect 244 4625 296 4641
rect 244 4557 296 4573
rect 244 4499 296 4505
rect 329 5073 335 5107
rect 369 5073 375 5107
rect 958 5101 1010 5119
rect 329 5035 375 5073
rect 417 5038 445 5090
rect 497 5038 509 5090
rect 561 5038 573 5090
rect 625 5038 631 5090
rect 958 5043 1010 5049
tri 1046 5324 1066 5344 se
rect 1066 5324 1102 5344
tri 1102 5324 1122 5344 nw
rect 1471 5328 1523 5341
rect 1046 5151 1092 5324
tri 1092 5314 1102 5324 nw
rect 1046 5117 1052 5151
rect 1086 5117 1092 5151
rect 1046 5079 1092 5117
rect 1046 5045 1052 5079
rect 1086 5045 1092 5079
rect 329 5001 335 5035
rect 369 5013 375 5035
tri 1045 5017 1046 5018 se
rect 1046 5017 1092 5045
tri 1043 5015 1045 5017 se
rect 1045 5015 1092 5017
tri 375 5013 377 5015 sw
tri 1041 5013 1043 5015 se
rect 1043 5013 1092 5015
rect 369 5001 377 5013
rect 329 4989 377 5001
tri 377 4989 401 5013 sw
tri 1017 4989 1041 5013 se
rect 1041 4998 1092 5013
rect 1041 4989 1077 4998
rect 329 4983 401 4989
tri 401 4983 407 4989 sw
tri 1011 4983 1017 4989 se
rect 1017 4983 1077 4989
tri 1077 4983 1092 4998 nw
rect 1120 5290 1166 5302
rect 1120 5256 1126 5290
rect 1160 5256 1166 5290
rect 1120 5218 1166 5256
rect 1471 5271 1480 5276
rect 1514 5271 1523 5276
rect 1471 5263 1523 5271
rect 1120 5184 1126 5218
rect 1160 5184 1166 5218
rect 1215 5200 1221 5252
rect 1273 5200 1285 5252
rect 1337 5200 1352 5252
rect 1557 5283 1603 5495
rect 1769 5510 2705 5516
rect 1885 5444 2705 5510
rect 1885 5394 2655 5444
tri 2655 5394 2705 5444 nw
rect 2750 5516 2802 5522
tri 2802 5506 2818 5522 sw
tri 4609 5506 4625 5522 ne
rect 4625 5506 8591 5522
tri 8591 5506 8619 5534 nw
rect 2802 5503 4584 5506
tri 4584 5503 4587 5506 sw
tri 4625 5503 4628 5506 ne
rect 4628 5503 8588 5506
tri 8588 5503 8591 5506 nw
tri 8629 5503 8632 5506 se
rect 8632 5503 13858 5506
rect 2802 5500 4587 5503
tri 4587 5500 4590 5503 sw
tri 8626 5500 8629 5503 se
rect 8629 5500 13858 5503
rect 2802 5475 4590 5500
tri 4590 5475 4615 5500 sw
tri 8601 5475 8626 5500 se
rect 8626 5475 13740 5500
rect 2802 5470 13740 5475
rect 2802 5466 2823 5470
tri 2823 5466 2827 5470 nw
tri 4570 5466 4574 5470 ne
rect 4574 5466 8642 5470
tri 8642 5466 8646 5470 nw
tri 13718 5466 13722 5470 ne
rect 13722 5466 13740 5470
rect 13774 5466 13812 5500
rect 13846 5466 13858 5500
rect 2802 5464 2817 5466
rect 2750 5460 2817 5464
tri 2817 5460 2823 5466 nw
tri 4574 5460 4580 5466 ne
rect 4580 5460 8636 5466
tri 8636 5460 8642 5466 nw
tri 13722 5460 13728 5466 ne
rect 13728 5460 13858 5466
rect 2750 5452 2802 5460
tri 2802 5445 2817 5460 nw
tri 4580 5445 4595 5460 ne
rect 4595 5445 8615 5460
tri 4595 5439 4601 5445 ne
rect 4601 5439 8615 5445
tri 8615 5439 8636 5460 nw
tri 13947 5430 13953 5436 se
rect 13953 5430 14005 5945
rect 1885 5347 2608 5394
tri 2608 5347 2655 5394 nw
rect 2750 5392 2802 5400
rect 2931 5378 2937 5430
rect 2989 5378 3005 5430
rect 3057 5411 4463 5430
tri 4463 5411 4482 5430 sw
tri 13928 5411 13947 5430 se
rect 13947 5411 14005 5430
rect 3057 5378 4831 5411
tri 4449 5359 4468 5378 ne
rect 4468 5359 4831 5378
rect 4883 5359 4895 5411
rect 4947 5401 14005 5411
rect 4947 5359 13963 5401
tri 13963 5359 14005 5401 nw
tri 14818 5359 14823 5364 se
rect 14823 5359 16424 5364
tri 16424 5359 16429 5364 sw
tri 14806 5347 14818 5359 se
rect 14818 5347 16429 5359
tri 16429 5347 16441 5359 sw
rect 1885 5330 2585 5347
rect 1769 5324 2585 5330
tri 2585 5324 2608 5347 nw
rect 2830 5295 2836 5347
rect 2888 5295 2900 5347
rect 2952 5324 4386 5347
tri 4386 5324 4409 5347 sw
tri 14803 5344 14806 5347 se
rect 14806 5344 16441 5347
tri 16441 5344 16444 5347 sw
tri 14019 5330 14033 5344 se
rect 2952 5311 4409 5324
tri 4409 5311 4422 5324 sw
rect 2952 5305 4422 5311
tri 4422 5305 4428 5311 sw
rect 2952 5302 4428 5305
tri 4428 5302 4431 5305 sw
tri 10264 5302 10267 5305 se
rect 10267 5302 10319 5305
rect 2952 5295 4431 5302
tri 4360 5291 4364 5295 ne
rect 4364 5291 4431 5295
tri 1603 5283 1611 5291 sw
tri 4364 5283 4372 5291 ne
rect 4372 5283 4431 5291
tri 4431 5283 4450 5302 sw
tri 10245 5283 10264 5302 se
rect 10264 5299 10319 5302
rect 10264 5283 10267 5299
rect 1557 5271 1611 5283
tri 1611 5271 1623 5283 sw
tri 4372 5271 4384 5283 ne
rect 4384 5271 6780 5283
rect 1557 5269 1623 5271
tri 1623 5269 1625 5271 sw
tri 4384 5269 4386 5271 ne
rect 4386 5269 6780 5271
rect 1557 5266 1625 5269
tri 1625 5266 1628 5269 sw
tri 4386 5266 4389 5269 ne
rect 4389 5266 6780 5269
rect 1557 5260 3642 5266
tri 4389 5265 4390 5266 ne
rect 4390 5265 6780 5266
rect 1557 5220 3590 5260
rect 1120 5017 1166 5184
rect 1471 5198 1480 5211
rect 1514 5198 1523 5211
tri 3565 5210 3575 5220 ne
rect 3575 5210 3590 5220
tri 3575 5200 3585 5210 ne
rect 3585 5208 3590 5210
tri 4390 5252 4403 5265 ne
rect 4403 5252 6780 5265
rect 3585 5200 3642 5208
tri 3585 5195 3590 5200 ne
rect 3590 5192 3642 5200
rect 1471 5133 1480 5146
rect 1514 5133 1523 5146
rect 1471 5068 1480 5081
rect 1514 5068 1523 5081
tri 1166 5017 1167 5018 sw
rect 1120 5015 1167 5017
tri 1167 5015 1169 5017 sw
rect 1120 5013 1169 5015
tri 1169 5013 1171 5015 sw
rect 1471 5013 1523 5016
rect 1120 4993 1171 5013
tri 1171 4993 1191 5013 sw
rect 1471 5003 1480 5013
rect 1514 5003 1523 5013
rect 329 4931 699 4983
rect 751 4931 763 4983
rect 815 4979 1073 4983
tri 1073 4979 1077 4983 nw
rect 815 4977 1071 4979
tri 1071 4977 1073 4979 nw
rect 815 4963 1057 4977
tri 1057 4963 1071 4977 nw
rect 815 4962 1056 4963
tri 1056 4962 1057 4963 nw
tri 1119 4962 1120 4963 se
rect 1120 4962 1225 4993
rect 815 4943 1037 4962
tri 1037 4943 1056 4962 nw
tri 1100 4943 1119 4962 se
rect 1119 4947 1225 4962
rect 1119 4943 1166 4947
tri 1166 4943 1170 4947 nw
rect 815 4940 1034 4943
tri 1034 4940 1037 4943 nw
tri 1097 4940 1100 4943 se
rect 1100 4940 1163 4943
tri 1163 4940 1166 4943 nw
rect 1471 4940 1523 4951
rect 815 4931 1025 4940
tri 1025 4931 1034 4940 nw
tri 1088 4931 1097 4940 se
rect 1097 4931 1129 4940
rect 329 4906 388 4931
tri 388 4906 413 4931 nw
tri 1063 4906 1088 4931 se
rect 1088 4906 1129 4931
tri 1129 4906 1163 4940 nw
rect 1471 4938 1480 4940
rect 1514 4938 1523 4940
rect 329 4905 387 4906
tri 387 4905 388 4906 nw
tri 1062 4905 1063 4906 se
rect 1063 4905 1128 4906
tri 1128 4905 1129 4906 nw
rect 329 4903 385 4905
tri 385 4903 387 4905 nw
tri 1060 4903 1062 4905 se
rect 1062 4903 1126 4905
tri 1126 4903 1128 4905 nw
rect 329 4899 381 4903
tri 381 4899 385 4903 nw
tri 1056 4899 1060 4903 se
rect 1060 4899 1122 4903
tri 1122 4899 1126 4903 nw
rect 329 4756 375 4899
tri 375 4893 381 4899 nw
rect 687 4887 1092 4899
rect 687 4853 693 4887
rect 727 4869 1092 4887
tri 1092 4869 1122 4899 nw
rect 727 4867 1090 4869
tri 1090 4867 1092 4869 nw
rect 727 4853 1076 4867
tri 1076 4853 1090 4867 nw
rect 687 4833 744 4853
tri 744 4833 764 4853 nw
rect 1352 4837 1426 4883
tri 1352 4833 1356 4837 ne
rect 1356 4833 1426 4837
rect 687 4829 740 4833
tri 740 4829 744 4833 nw
tri 1356 4829 1360 4833 ne
rect 1360 4829 1426 4833
rect 439 4772 445 4824
rect 497 4772 509 4824
rect 561 4772 573 4824
rect 625 4772 631 4824
rect 687 4815 739 4829
tri 739 4828 740 4829 nw
tri 1360 4828 1361 4829 ne
rect 1361 4828 1426 4829
tri 1361 4815 1374 4828 ne
rect 1374 4815 1426 4828
rect 687 4781 693 4815
rect 727 4781 739 4815
rect 329 4722 335 4756
rect 369 4722 375 4756
rect 329 4684 375 4722
rect 687 4741 739 4781
tri 684 4687 687 4690 se
rect 687 4687 739 4689
rect 329 4650 335 4684
rect 369 4650 375 4684
tri 678 4681 684 4687 se
rect 684 4681 739 4687
tri 662 4665 678 4681 se
rect 678 4677 739 4681
rect 678 4665 687 4677
rect 244 4311 290 4323
rect 244 4277 250 4311
rect 284 4277 290 4311
rect 244 4233 290 4277
rect 244 4199 250 4233
rect 284 4199 290 4233
rect 244 4155 290 4199
rect 244 4121 250 4155
rect 284 4121 290 4155
rect 244 4078 290 4121
rect 244 4044 250 4078
rect 284 4044 290 4078
rect 244 4001 290 4044
rect 244 3967 250 4001
rect 284 3967 290 4001
rect 244 3924 290 3967
rect 244 3890 250 3924
rect 284 3890 290 3924
rect 244 3847 290 3890
rect 244 3813 250 3847
rect 284 3813 290 3847
rect 244 3770 290 3813
rect 8 3728 54 3740
rect 8 3694 14 3728
rect 48 3694 54 3728
rect 8 3656 54 3694
rect 8 3622 14 3656
rect 48 3622 54 3656
rect 8 3610 54 3622
rect 244 3736 250 3770
rect 284 3736 290 3770
rect 329 4055 375 4650
rect 599 4625 687 4665
rect 599 4619 739 4625
rect 772 4803 818 4815
tri 1374 4809 1380 4815 ne
rect 772 4769 778 4803
rect 812 4769 818 4803
rect 772 4729 818 4769
rect 772 4695 778 4729
rect 812 4695 818 4729
rect 772 4655 818 4695
rect 849 4799 1092 4805
rect 901 4793 1092 4799
rect 901 4759 1052 4793
rect 1086 4759 1092 4793
rect 901 4747 1092 4759
rect 849 4735 1092 4747
rect 901 4721 1092 4735
rect 901 4687 1052 4721
rect 1086 4687 1092 4721
rect 901 4683 1092 4687
rect 849 4675 1092 4683
rect 772 4621 778 4655
rect 812 4621 818 4655
tri 771 4575 772 4576 se
rect 772 4575 818 4621
tri 754 4558 771 4575 se
rect 771 4558 818 4575
tri 747 4551 754 4558 se
rect 754 4551 818 4558
rect 403 4499 409 4551
rect 461 4499 495 4551
rect 547 4542 582 4551
rect 634 4542 818 4551
rect 547 4508 577 4542
rect 634 4508 658 4542
rect 692 4508 740 4542
rect 774 4508 818 4542
rect 547 4499 582 4508
rect 634 4499 818 4508
rect 958 4641 1010 4647
rect 958 4565 1010 4589
rect 958 4490 1010 4513
rect 958 4415 1010 4438
tri 945 4329 958 4342 se
rect 958 4340 1010 4363
tri 933 4317 945 4329 se
rect 945 4317 958 4329
rect 403 4311 958 4317
rect 403 4277 415 4311
rect 449 4277 496 4311
rect 530 4277 577 4311
rect 611 4277 658 4311
rect 692 4277 740 4311
rect 774 4288 958 4311
rect 774 4277 1010 4288
rect 403 4271 1010 4277
tri 747 4253 765 4271 ne
rect 765 4265 1010 4271
rect 765 4253 958 4265
tri 765 4246 772 4253 ne
rect 772 4213 958 4253
rect 772 4207 1010 4213
rect 1046 4601 1150 4647
rect 1046 4575 1094 4601
tri 1094 4575 1120 4601 nw
rect 619 4176 669 4200
tri 669 4176 693 4200 sw
tri 1022 4176 1046 4200 se
rect 1046 4176 1092 4575
tri 1092 4573 1094 4575 nw
tri 1370 4429 1380 4439 se
rect 1380 4429 1426 4815
tri 1352 4411 1370 4429 se
rect 1370 4411 1426 4429
rect 1352 4365 1426 4411
tri 1352 4356 1361 4365 ne
rect 1361 4356 1426 4365
tri 1361 4337 1380 4356 ne
tri 1092 4176 1119 4203 sw
rect 619 4175 693 4176
tri 693 4175 694 4176 sw
tri 1021 4175 1022 4176 se
rect 1022 4175 1119 4176
tri 1119 4175 1120 4176 sw
rect 619 4154 1150 4175
tri 649 4137 666 4154 ne
rect 666 4137 1150 4154
tri 666 4116 687 4137 ne
rect 687 4129 1150 4137
rect 687 4116 745 4129
tri 745 4116 758 4129 nw
tri 375 4055 382 4062 sw
rect 329 4030 382 4055
tri 382 4030 407 4055 sw
rect 329 4024 407 4030
tri 407 4024 413 4030 sw
rect 329 3978 443 4024
rect 329 3969 404 3978
tri 404 3969 413 3978 nw
rect 329 3957 392 3969
tri 392 3957 404 3969 nw
rect 329 3946 381 3957
tri 381 3946 392 3957 nw
rect 329 3944 379 3946
tri 379 3944 381 3946 nw
rect 329 3942 377 3944
tri 377 3942 379 3944 nw
rect 329 3941 376 3942
tri 376 3941 377 3942 nw
rect 329 3793 375 3941
tri 375 3940 376 3941 nw
tri 684 3883 687 3886 se
rect 687 3883 733 4116
tri 733 4104 745 4116 nw
tri 673 3872 684 3883 se
rect 684 3872 733 3883
tri 668 3867 673 3872 se
rect 673 3867 733 3872
tri 660 3859 668 3867 se
rect 668 3859 733 3867
tri 649 3848 660 3859 se
rect 660 3848 733 3859
rect 619 3802 733 3848
rect 772 4089 818 4101
rect 772 4055 778 4089
rect 812 4055 818 4089
rect 772 4003 818 4055
rect 772 3969 778 4003
rect 812 3969 818 4003
rect 772 3917 818 3969
rect 772 3883 778 3917
rect 812 3884 818 3917
rect 849 4095 1096 4101
rect 901 4089 1096 4095
rect 901 4055 1052 4089
rect 1086 4055 1096 4089
rect 901 4043 1096 4055
rect 849 4031 1096 4043
rect 901 4017 1096 4031
rect 901 3983 1052 4017
rect 1086 3983 1096 4017
rect 901 3979 1096 3983
rect 849 3967 1096 3979
rect 901 3915 1096 3967
tri 1370 3957 1380 3967 se
rect 1380 3957 1426 4356
tri 1359 3946 1370 3957 se
rect 1370 3946 1426 3957
tri 1357 3944 1359 3946 se
rect 1359 3944 1426 3946
tri 1355 3942 1357 3944 se
rect 1357 3942 1426 3944
tri 1354 3941 1355 3942 se
rect 1355 3941 1426 3942
rect 849 3909 1096 3915
tri 1352 3939 1354 3941 se
rect 1354 3939 1426 3941
tri 818 3884 830 3896 sw
rect 1352 3893 1426 3939
tri 1352 3884 1361 3893 ne
rect 1361 3884 1426 3893
rect 812 3883 830 3884
rect 772 3872 830 3883
tri 830 3872 842 3884 sw
tri 1361 3872 1373 3884 ne
rect 1373 3872 1426 3884
rect 772 3871 842 3872
tri 842 3871 843 3872 sw
tri 1373 3871 1374 3872 ne
rect 1374 3871 1426 3872
rect 772 3865 1010 3871
tri 1374 3867 1378 3871 ne
rect 1378 3867 1426 3871
tri 1378 3865 1380 3867 ne
rect 772 3831 958 3865
rect 772 3797 778 3831
rect 812 3813 958 3831
rect 812 3797 1010 3813
tri 375 3793 379 3797 sw
rect 329 3785 379 3793
tri 379 3785 387 3793 sw
rect 772 3792 1010 3797
rect 329 3777 387 3785
tri 387 3777 395 3785 sw
tri 329 3759 347 3777 ne
rect 347 3759 395 3777
tri 395 3759 413 3777 sw
tri 347 3751 355 3759 ne
rect 355 3755 413 3759
tri 413 3755 417 3759 sw
rect 355 3751 417 3755
tri 417 3751 421 3755 sw
tri 355 3746 360 3751 ne
rect 360 3746 421 3751
tri 421 3746 426 3751 sw
rect 772 3746 958 3792
rect 1150 3759 1156 3811
rect 1208 3759 1220 3811
rect 1272 3759 1284 3811
rect 1336 3759 1352 3811
tri 360 3740 366 3746 ne
rect 366 3740 426 3746
tri 426 3740 432 3746 sw
rect 244 3689 290 3736
tri 366 3712 394 3740 ne
rect 394 3712 432 3740
tri 432 3712 460 3740 sw
rect 772 3712 778 3746
rect 812 3740 958 3746
tri 1373 3740 1380 3747 se
rect 1380 3740 1426 3867
rect 812 3720 1010 3740
rect 812 3712 958 3720
tri 394 3711 395 3712 ne
rect 395 3711 460 3712
tri 460 3711 461 3712 sw
tri 395 3704 402 3711 ne
rect 402 3704 461 3711
tri 290 3689 305 3704 sw
tri 402 3689 417 3704 ne
rect 417 3689 461 3704
tri 461 3689 483 3711 sw
rect 772 3700 958 3712
tri 933 3689 944 3700 ne
rect 944 3689 958 3700
rect 244 3677 305 3689
tri 305 3677 317 3689 sw
rect 417 3677 483 3689
tri 483 3677 495 3689 sw
tri 944 3677 956 3689 ne
rect 956 3677 958 3689
rect 244 3672 317 3677
tri 317 3672 322 3677 sw
rect 417 3672 495 3677
tri 495 3672 500 3677 sw
tri 956 3675 958 3677 ne
rect 244 3665 322 3672
tri 322 3665 329 3672 sw
rect 619 3666 821 3672
rect 244 3664 329 3665
tri 329 3664 330 3665 sw
rect 244 3656 330 3664
tri 330 3656 338 3664 sw
rect 244 3638 338 3656
tri 338 3638 356 3656 sw
rect 244 3626 356 3638
tri 356 3626 368 3638 sw
rect 619 3626 769 3666
rect 244 3610 368 3626
tri 368 3610 384 3626 sw
tri 744 3610 760 3626 ne
rect 760 3614 769 3626
rect 760 3610 821 3614
rect 244 3604 384 3610
tri 384 3604 390 3610 sw
tri 760 3604 766 3610 ne
rect 766 3604 821 3610
rect 244 3601 390 3604
tri 390 3601 393 3604 sw
tri 766 3601 769 3604 ne
rect 769 3602 821 3604
rect 244 3595 393 3601
tri 244 3592 247 3595 ne
rect 247 3592 393 3595
tri 393 3592 402 3601 sw
tri 247 3584 255 3592 ne
rect 255 3584 402 3592
tri 402 3584 410 3592 sw
tri 255 3565 274 3584 ne
rect 274 3565 410 3584
tri 410 3565 429 3584 sw
tri 274 3549 290 3565 ne
rect 290 3555 429 3565
tri 429 3555 439 3565 sw
rect 290 3549 741 3555
tri 290 3515 324 3549 ne
rect 324 3515 399 3549
rect 433 3515 473 3549
rect 507 3515 547 3549
rect 581 3515 621 3549
rect 655 3515 695 3549
rect 729 3531 741 3549
rect 769 3544 821 3550
rect 958 3648 1010 3668
rect 958 3576 1010 3596
tri 956 3532 958 3534 se
tri 741 3531 742 3532 sw
tri 955 3531 956 3532 se
rect 956 3531 958 3532
rect 729 3515 742 3531
tri 324 3512 327 3515 ne
rect 327 3512 742 3515
tri 742 3512 761 3531 sw
tri 936 3512 955 3531 se
rect 955 3524 958 3531
rect 955 3512 1010 3524
tri 327 3509 330 3512 ne
rect 330 3509 761 3512
tri 761 3509 764 3512 sw
tri 933 3509 936 3512 se
rect 936 3509 1010 3512
tri 330 3507 332 3509 ne
rect 332 3507 764 3509
tri 764 3507 766 3509 sw
tri 931 3507 933 3509 se
rect 933 3507 1010 3509
tri 332 3500 339 3507 ne
rect 339 3504 1010 3507
rect 339 3500 958 3504
rect 240 3494 292 3500
tri 339 3492 347 3500 ne
rect 347 3492 958 3500
tri 347 3458 381 3492 ne
rect 381 3458 958 3492
tri 381 3446 393 3458 ne
rect 393 3452 958 3458
rect 393 3446 1010 3452
rect 1046 3728 1092 3740
tri 1371 3738 1373 3740 se
rect 1373 3738 1426 3740
rect 1046 3694 1052 3728
rect 1086 3694 1092 3728
tri 1352 3719 1371 3738 se
rect 1371 3719 1426 3738
rect 1046 3656 1092 3694
rect 1150 3713 1426 3719
rect 1150 3679 1162 3713
rect 1196 3679 1234 3713
rect 1268 3679 1306 3713
rect 1340 3679 1426 3713
rect 1150 3673 1426 3679
tri 1352 3665 1360 3673 ne
rect 1360 3665 1426 3673
rect 1046 3622 1052 3656
rect 1086 3622 1092 3656
tri 1360 3646 1379 3665 ne
rect 1379 3646 1426 3665
tri 1379 3645 1380 3646 ne
rect 1046 3584 1092 3622
rect 1046 3550 1052 3584
rect 1086 3550 1092 3584
rect 1150 3581 1156 3633
rect 1208 3581 1220 3633
rect 1272 3581 1284 3633
rect 1336 3581 1352 3633
tri 1364 3553 1380 3569 se
rect 1380 3553 1426 3646
rect 1046 3512 1092 3550
tri 1352 3541 1364 3553 se
rect 1364 3541 1426 3553
rect 1046 3478 1052 3512
rect 1086 3478 1092 3512
rect 1150 3535 1426 3541
rect 1150 3501 1162 3535
rect 1196 3501 1234 3535
rect 1268 3501 1306 3535
rect 1340 3501 1426 3535
rect 1150 3495 1426 3501
rect 1471 4873 1523 4886
rect 1471 4808 1523 4821
rect 1471 4743 1523 4756
rect 1471 4687 1480 4691
rect 1514 4687 1523 4691
rect 1471 4678 1523 4687
rect 1471 4614 1480 4626
rect 1514 4614 1523 4626
rect 1471 4613 1523 4614
rect 1471 4548 1480 4561
rect 1514 4548 1523 4561
rect 1471 4483 1480 4496
rect 1514 4483 1523 4496
rect 1471 4429 1523 4431
rect 1471 4418 1480 4429
rect 1514 4418 1523 4429
rect 1471 4356 1523 4366
rect 1471 4353 1480 4356
rect 1514 4353 1523 4356
rect 1471 4287 1523 4301
rect 1471 4221 1523 4235
rect 1471 4155 1523 4169
rect 1471 4089 1523 4103
rect 1471 4030 1480 4037
rect 1514 4030 1523 4037
rect 1471 4023 1523 4030
rect 1471 3957 1480 3971
rect 1514 3957 1523 3971
rect 1471 3891 1480 3905
rect 1514 3891 1523 3905
rect 1471 3825 1480 3839
rect 1514 3825 1523 3839
rect 1471 3772 1523 3773
rect 1471 3759 1480 3772
rect 1514 3759 1523 3772
rect 1471 3699 1523 3707
rect 1471 3693 1480 3699
rect 1514 3693 1523 3699
rect 1471 3627 1523 3641
rect 1471 3561 1523 3575
rect 1471 3495 1523 3509
tri 292 3442 293 3443 sw
rect 240 3430 293 3442
rect 292 3427 293 3430
tri 293 3427 308 3442 sw
rect 292 3418 308 3427
tri 308 3418 317 3427 sw
rect 292 3378 1018 3418
rect 240 3372 1018 3378
tri 947 3354 965 3372 ne
rect 965 3354 1018 3372
tri 965 3347 972 3354 ne
rect 0 3338 808 3344
rect 0 3304 372 3338
rect 406 3304 450 3338
rect 484 3304 528 3338
rect 562 3304 606 3338
rect 640 3304 684 3338
rect 718 3304 762 3338
rect 796 3304 808 3338
rect 0 3300 808 3304
rect 0 3266 250 3300
rect 284 3298 808 3300
rect 849 3325 901 3331
rect 284 3280 297 3298
tri 297 3280 315 3298 nw
tri 834 3280 849 3295 se
rect 284 3266 290 3280
tri 290 3273 297 3280 nw
tri 827 3273 834 3280 se
rect 834 3273 849 3280
tri 824 3270 827 3273 se
rect 827 3270 901 3273
rect 0 3221 290 3266
rect 0 3187 250 3221
rect 284 3187 290 3221
rect 0 3142 290 3187
rect 0 3108 250 3142
rect 284 3108 290 3142
rect 0 3064 290 3108
rect 0 3030 250 3064
rect 284 3030 290 3064
rect 0 3018 290 3030
rect 329 3261 901 3270
rect 329 3252 849 3261
rect 329 3200 445 3252
rect 497 3200 509 3252
rect 561 3200 573 3252
rect 625 3209 849 3252
rect 625 3200 901 3209
rect 972 3314 1018 3354
rect 972 3280 978 3314
rect 1012 3280 1018 3314
rect 972 3242 1018 3280
rect 972 3208 978 3242
rect 1012 3208 1018 3242
rect 329 3196 428 3200
tri 428 3196 432 3200 nw
rect 972 3196 1018 3208
rect 329 3185 417 3196
tri 417 3185 428 3196 nw
rect 240 2977 292 2985
rect 240 2913 292 2925
rect 240 2855 292 2861
rect 329 2885 401 3185
tri 401 3169 417 3185 nw
tri 1033 3169 1046 3182 se
rect 1046 3169 1092 3478
rect 1150 3412 1156 3464
rect 1208 3412 1220 3464
rect 1272 3412 1284 3464
rect 1336 3412 1352 3464
rect 1471 3429 1523 3443
rect 1471 3373 1480 3377
rect 1514 3373 1523 3377
rect 1471 3363 1523 3373
rect 1352 3259 1426 3305
tri 1352 3231 1380 3259 ne
tri 1028 3164 1033 3169 se
rect 1033 3164 1092 3169
rect 1150 3164 1156 3216
rect 1208 3164 1220 3216
rect 1272 3164 1284 3216
rect 1336 3164 1352 3216
tri 1021 3157 1028 3164 se
rect 1028 3157 1092 3164
rect 631 3151 1092 3157
tri 1092 3151 1098 3157 sw
rect 631 3143 1098 3151
tri 1098 3143 1106 3151 sw
rect 631 3135 1106 3143
tri 1106 3135 1114 3143 sw
rect 631 3121 1114 3135
tri 1114 3121 1128 3135 sw
rect 631 3111 1150 3121
tri 1072 3077 1106 3111 ne
rect 1106 3077 1150 3111
tri 1106 3075 1108 3077 ne
rect 1108 3075 1150 3077
rect 631 3041 901 3047
rect 631 3001 849 3041
tri 819 2994 826 3001 ne
rect 826 2994 849 3001
tri 826 2989 831 2994 ne
rect 831 2989 849 2994
tri 901 3039 909 3047 sw
rect 901 3037 909 3039
tri 909 3037 911 3039 sw
tri 1378 3037 1380 3039 se
rect 1380 3037 1426 3259
rect 901 3011 911 3037
tri 911 3011 937 3037 sw
tri 1352 3011 1378 3037 se
rect 1378 3011 1426 3037
rect 901 2989 1150 3011
tri 831 2971 849 2989 ne
rect 849 2977 1150 2989
rect 557 2909 631 2950
rect 901 2965 1150 2977
rect 1352 2965 1426 3011
rect 1471 3299 1480 3311
rect 1514 3299 1523 3311
rect 1471 3297 1523 3299
rect 1471 3231 1480 3245
rect 1514 3231 1523 3245
rect 1471 3165 1480 3179
rect 1514 3165 1523 3179
rect 1471 3111 1523 3113
rect 1471 3099 1480 3111
rect 1514 3099 1523 3111
rect 1471 3037 1523 3047
rect 1471 3033 1480 3037
rect 1514 3033 1523 3037
rect 1471 2967 1523 2981
rect 901 2963 945 2965
tri 945 2963 947 2965 nw
rect 901 2931 913 2963
tri 913 2931 945 2963 nw
rect 901 2929 911 2931
tri 911 2929 913 2931 nw
rect 901 2927 909 2929
tri 909 2927 911 2929 nw
rect 849 2919 901 2925
tri 901 2919 909 2927 nw
rect 958 2925 1010 2931
rect 1663 5163 3020 5172
rect 3072 5163 3122 5172
rect 1663 5129 1785 5163
rect 1819 5129 1860 5163
rect 1894 5129 1935 5163
rect 1969 5129 2010 5163
rect 2044 5129 2085 5163
rect 2119 5129 2160 5163
rect 2194 5129 2235 5163
rect 2269 5129 2310 5163
rect 2344 5129 2385 5163
rect 2419 5129 2460 5163
rect 2494 5129 2536 5163
rect 2570 5129 2612 5163
rect 2646 5129 2688 5163
rect 2722 5129 2764 5163
rect 2798 5129 2840 5163
rect 2874 5129 2916 5163
rect 2950 5129 2992 5163
rect 3102 5129 3122 5163
rect 3590 5134 3642 5140
rect 3670 5244 4124 5252
rect 3670 5210 3744 5244
rect 3778 5210 3816 5244
rect 3850 5210 3888 5244
rect 3922 5210 3960 5244
rect 3994 5210 4032 5244
rect 4066 5210 4104 5244
rect 3670 5200 4124 5210
rect 4176 5200 4188 5252
rect 4240 5200 4246 5252
tri 4403 5227 4428 5252 ne
rect 4428 5231 6780 5252
rect 6832 5231 6844 5283
rect 6896 5247 10267 5283
rect 11853 5278 11859 5330
rect 11911 5278 11926 5330
rect 11978 5278 12407 5330
rect 12459 5278 12474 5330
rect 12526 5278 12532 5330
tri 14008 5319 14019 5330 se
rect 14019 5319 14033 5330
tri 14778 5319 14803 5344 se
rect 14803 5319 16444 5344
tri 16444 5319 16469 5344 sw
rect 12587 5270 14085 5319
tri 14777 5318 14778 5319 se
rect 14778 5318 16469 5319
tri 16469 5318 16470 5319 sw
tri 14770 5311 14777 5318 se
rect 14777 5311 14823 5318
rect 14343 5305 14473 5311
rect 14343 5271 14355 5305
rect 14389 5271 14427 5305
rect 14461 5271 14473 5305
rect 12587 5265 12661 5270
tri 12661 5265 12666 5270 nw
rect 14343 5265 14473 5271
rect 14501 5305 14631 5311
rect 14501 5271 14513 5305
rect 14547 5271 14585 5305
rect 14619 5271 14631 5305
tri 14757 5298 14770 5311 se
rect 14770 5298 14823 5311
tri 14823 5298 14843 5318 nw
tri 16404 5298 16424 5318 ne
rect 16424 5298 16491 5318
rect 14501 5265 14631 5271
tri 14724 5265 14757 5298 se
rect 14757 5265 14762 5298
rect 12587 5251 12647 5265
tri 12647 5251 12661 5265 nw
tri 14710 5251 14724 5265 se
rect 14724 5251 14762 5265
rect 6896 5235 10319 5247
rect 6896 5231 10267 5235
rect 4428 5227 10267 5231
tri 10221 5200 10248 5227 ne
rect 10248 5200 10267 5227
rect 3670 5172 4168 5200
tri 4168 5172 4196 5200 nw
tri 10248 5181 10267 5200 ne
rect 10267 5177 10319 5183
rect 11455 5245 11507 5251
rect 11507 5193 12234 5227
rect 11455 5178 12234 5193
rect 3670 5162 4158 5172
tri 4158 5162 4168 5172 nw
rect 3670 5153 4150 5162
tri 4150 5154 4158 5162 nw
rect 1663 5125 3020 5129
rect 1663 5091 1669 5125
rect 1703 5120 3020 5125
rect 3072 5120 3122 5129
rect 1703 5119 1733 5120
tri 1733 5119 1734 5120 nw
tri 3045 5119 3046 5120 ne
rect 3046 5119 3122 5120
rect 1703 5091 1709 5119
tri 1709 5095 1733 5119 nw
tri 3046 5095 3070 5119 ne
rect 1663 5051 1709 5091
rect 3070 5091 3122 5119
rect 3670 5119 3713 5153
rect 3747 5119 3792 5153
rect 3826 5119 3870 5153
rect 3904 5119 3948 5153
rect 3982 5119 4026 5153
rect 4060 5119 4104 5153
rect 4138 5119 4150 5153
rect 11507 5175 12234 5178
rect 12286 5175 12301 5227
rect 12353 5175 12359 5227
rect 4829 5124 9554 5126
rect 3070 5079 3079 5091
rect 3113 5079 3122 5091
tri 3643 5089 3670 5116 se
rect 3670 5113 4150 5119
rect 4637 5118 4689 5124
rect 3670 5089 3737 5113
tri 3737 5089 3761 5113 nw
rect 4258 5108 4310 5114
tri 3234 5086 3237 5089 se
rect 3237 5086 3300 5089
tri 3231 5083 3234 5086 se
rect 3234 5083 3300 5086
tri 3220 5072 3231 5083 se
rect 3231 5072 3300 5083
rect 3706 5086 3734 5089
tri 3734 5086 3737 5089 nw
rect 3706 5085 3733 5086
tri 3733 5085 3734 5086 nw
rect 3706 5083 3731 5085
tri 3731 5083 3733 5085 nw
rect 3706 5072 3720 5083
tri 3720 5072 3731 5083 nw
rect 3932 5079 4150 5085
tri 3706 5058 3720 5072 nw
rect 1663 5017 1669 5051
rect 1703 5017 1709 5051
rect 1663 4977 1709 5017
rect 1820 5003 2032 5055
rect 2084 5003 2096 5055
rect 2148 5003 2160 5055
rect 2212 5003 2224 5055
rect 2276 5003 2288 5055
rect 2340 5003 2403 5055
rect 1663 4943 1669 4977
rect 1703 4943 1709 4977
rect 1663 4903 1709 4943
rect 1663 4869 1669 4903
rect 1703 4869 1709 4903
rect 1663 4829 1709 4869
rect 1663 4795 1669 4829
rect 1703 4795 1709 4829
rect 1663 4755 1709 4795
rect 1663 4721 1669 4755
rect 1703 4721 1709 4755
rect 1663 4681 1709 4721
rect 1663 4647 1669 4681
rect 1703 4647 1709 4681
rect 1663 4607 1709 4647
tri 1792 4981 1794 4983 sw
tri 2476 4981 2478 4983 se
rect 2478 4981 2527 5017
rect 1792 4973 1794 4981
tri 1794 4973 1802 4981 sw
tri 2468 4973 2476 4981 se
rect 2476 4973 2527 4981
rect 2566 4973 2572 5025
rect 2624 4973 2636 5025
rect 2688 4973 2882 5025
rect 3070 5015 3122 5027
rect 3070 5012 3079 5015
rect 3113 5012 3122 5015
rect 1792 4971 1802 4973
tri 1802 4971 1804 4973 sw
tri 2466 4971 2468 4973 se
rect 2468 4971 2527 4973
rect 1792 4958 1804 4971
tri 1804 4958 1817 4971 sw
tri 2453 4958 2466 4971 se
rect 2466 4958 2527 4971
rect 1792 4952 2527 4958
rect 1792 4900 1946 4952
rect 1998 4900 2527 4952
rect 1792 4868 2527 4900
rect 1792 4816 1946 4868
rect 1998 4816 2527 4868
rect 1792 4785 2527 4816
rect 1792 4733 1946 4785
rect 1998 4733 2527 4785
rect 1792 4702 2527 4733
rect 1792 4650 1946 4702
rect 1998 4650 2527 4702
rect 1792 4644 2527 4650
rect 1792 4640 1813 4644
tri 1813 4640 1817 4644 nw
tri 2453 4640 2457 4644 ne
rect 2457 4640 2527 4644
rect 1792 4635 1808 4640
tri 1808 4635 1813 4640 nw
tri 2457 4635 2462 4640 ne
rect 2462 4635 2527 4640
tri 1792 4619 1808 4635 nw
tri 2462 4619 2478 4635 ne
rect 1663 4573 1669 4607
rect 1703 4573 1709 4607
rect 1663 4533 1709 4573
rect 1820 4547 2032 4599
rect 2084 4547 2096 4599
rect 2148 4547 2160 4599
rect 2212 4547 2224 4599
rect 2276 4547 2288 4599
rect 2340 4547 2403 4599
rect 1663 4499 1669 4533
rect 1703 4499 1709 4533
rect 1663 4459 1709 4499
rect 1663 4425 1669 4459
rect 1703 4425 1709 4459
rect 1663 4385 1709 4425
rect 1663 4351 1669 4385
rect 1703 4351 1709 4385
rect 1663 4311 1709 4351
rect 1663 4277 1669 4311
rect 1703 4277 1709 4311
rect 1663 4237 1709 4277
rect 1663 4203 1669 4237
rect 1703 4203 1709 4237
rect 1663 4163 1709 4203
tri 1792 4525 1794 4527 sw
tri 2476 4525 2478 4527 se
rect 2478 4525 2527 4635
rect 3070 4945 3122 4960
rect 3932 5027 4098 5079
rect 3932 5015 4150 5027
rect 3932 4963 4098 5015
rect 3932 4957 4150 4963
rect 4258 5026 4266 5056
rect 4300 5026 4310 5056
rect 3070 4878 3122 4893
rect 3070 4811 3122 4826
rect 4258 4954 4310 4974
rect 4258 4944 4266 4954
rect 4300 4944 4310 4954
rect 4258 4862 4310 4892
rect 4258 4804 4310 4810
rect 4637 5049 4689 5066
rect 4637 4980 4689 4997
rect 4637 4911 4689 4928
rect 4829 5120 5034 5124
rect 5086 5120 5100 5124
rect 5152 5120 5166 5124
rect 5218 5120 5232 5124
rect 5284 5120 5298 5124
rect 5350 5120 5364 5124
rect 5416 5120 5430 5124
rect 5482 5120 5496 5124
rect 5548 5120 5562 5124
rect 4829 5086 4841 5120
rect 4875 5086 4913 5120
rect 4947 5086 4985 5120
rect 5019 5086 5034 5120
rect 5091 5086 5100 5120
rect 5163 5086 5166 5120
rect 5416 5086 5417 5120
rect 5482 5086 5489 5120
rect 5548 5086 5561 5120
rect 4829 5072 5034 5086
rect 5086 5072 5100 5086
rect 5152 5072 5166 5086
rect 5218 5072 5232 5086
rect 5284 5072 5298 5086
rect 5350 5072 5364 5086
rect 5416 5072 5430 5086
rect 5482 5072 5496 5086
rect 5548 5072 5562 5086
rect 5614 5072 5628 5124
rect 5680 5072 5694 5124
rect 5746 5072 5760 5124
rect 5812 5072 5826 5124
rect 5878 5120 5892 5124
rect 5944 5120 5959 5124
rect 6011 5120 6142 5124
rect 5883 5086 5892 5120
rect 5955 5086 5959 5120
rect 6027 5086 6065 5120
rect 6099 5086 6137 5120
rect 5878 5072 5892 5086
rect 5944 5072 5959 5086
rect 6011 5072 6142 5086
rect 6194 5072 6206 5124
rect 6258 5072 6270 5124
rect 6322 5072 6334 5124
rect 6386 5120 6399 5124
rect 6451 5120 6464 5124
rect 6516 5120 6529 5124
rect 6581 5120 6594 5124
rect 6646 5120 6969 5124
rect 7021 5120 7045 5124
rect 7097 5120 7121 5124
rect 7173 5120 7197 5124
rect 7249 5120 7273 5124
rect 7325 5120 7393 5124
rect 7445 5120 7461 5124
rect 7513 5120 7529 5124
rect 7581 5120 7598 5124
rect 7650 5120 7667 5124
rect 7719 5120 7736 5124
rect 6387 5086 6399 5120
rect 6459 5086 6464 5120
rect 6675 5086 6713 5120
rect 6747 5086 6785 5120
rect 6819 5086 6858 5120
rect 6892 5086 6931 5120
rect 6965 5086 6969 5120
rect 7038 5086 7045 5120
rect 7111 5086 7121 5120
rect 7184 5086 7197 5120
rect 7257 5086 7273 5120
rect 7330 5086 7369 5120
rect 7513 5086 7515 5120
rect 7581 5086 7588 5120
rect 7650 5086 7661 5120
rect 7719 5086 7734 5120
rect 6386 5072 6399 5086
rect 6451 5072 6464 5086
rect 6516 5072 6529 5086
rect 6581 5072 6594 5086
rect 6646 5072 6969 5086
rect 7021 5072 7045 5086
rect 7097 5072 7121 5086
rect 7173 5072 7197 5086
rect 7249 5072 7273 5086
rect 7325 5072 7393 5086
rect 7445 5072 7461 5086
rect 7513 5072 7529 5086
rect 7581 5072 7598 5086
rect 7650 5072 7667 5086
rect 7719 5072 7736 5086
rect 7788 5072 7805 5124
rect 7857 5072 7874 5124
rect 7926 5072 7943 5124
rect 7995 5072 8012 5124
rect 8064 5120 8187 5124
rect 8239 5120 8255 5124
rect 8307 5120 8323 5124
rect 8064 5086 8099 5120
rect 8133 5086 8172 5120
rect 8239 5086 8245 5120
rect 8307 5086 8318 5120
rect 8064 5072 8187 5086
rect 8239 5072 8255 5086
rect 8307 5072 8323 5086
rect 8375 5072 8391 5124
rect 8443 5072 8459 5124
rect 8511 5072 8528 5124
rect 8580 5072 8597 5124
rect 8649 5072 8666 5124
rect 8718 5072 8735 5124
rect 8787 5120 8804 5124
rect 8856 5120 8873 5124
rect 8925 5120 8942 5124
rect 8994 5120 9011 5124
rect 9063 5120 9080 5124
rect 9132 5120 9554 5124
rect 8790 5086 8804 5120
rect 8863 5086 8873 5120
rect 8936 5086 8942 5120
rect 9009 5086 9011 5120
rect 9155 5086 9194 5120
rect 9228 5086 9267 5120
rect 9301 5086 9340 5120
rect 9374 5086 9413 5120
rect 9447 5117 9554 5120
rect 9606 5117 9622 5126
rect 9674 5117 9690 5126
rect 9742 5117 9759 5126
rect 9811 5117 9828 5126
rect 9880 5117 9897 5126
rect 9949 5117 9966 5126
rect 10018 5117 10490 5126
rect 10542 5117 10554 5126
rect 10606 5117 10618 5126
rect 9447 5103 9506 5117
rect 9447 5086 9459 5103
rect 8787 5072 8804 5086
rect 8856 5072 8873 5086
rect 8925 5072 8942 5086
rect 8994 5072 9011 5086
rect 9063 5072 9080 5086
rect 9132 5072 9459 5086
rect 9540 5083 9554 5117
rect 9614 5083 9622 5117
rect 9688 5083 9690 5117
rect 9949 5083 9950 5117
rect 10018 5083 10024 5117
rect 10058 5083 10098 5117
rect 10132 5083 10172 5117
rect 10206 5083 10246 5117
rect 10280 5083 10320 5117
rect 10354 5083 10394 5117
rect 10428 5083 10468 5117
rect 10606 5083 10616 5117
rect 4829 5066 4892 5072
rect 4829 5024 4840 5066
tri 4892 5047 4917 5072 nw
tri 9434 5047 9459 5072 ne
rect 9511 5074 9554 5083
rect 9606 5074 9622 5083
rect 9674 5074 9690 5083
rect 9742 5074 9759 5083
rect 9811 5074 9828 5083
rect 9880 5074 9897 5083
rect 9949 5074 9966 5083
rect 10018 5074 10490 5083
rect 10542 5074 10554 5083
rect 10606 5074 10618 5083
rect 10670 5074 10682 5126
rect 10734 5074 10747 5126
rect 10799 5074 10812 5126
rect 10864 5117 10877 5126
rect 10929 5117 10942 5126
rect 10994 5117 11007 5126
rect 11059 5117 11207 5126
rect 10872 5083 10877 5117
rect 11059 5083 11060 5117
rect 11094 5083 11134 5117
rect 11168 5083 11207 5117
rect 10864 5074 10877 5083
rect 10929 5074 10942 5083
rect 10994 5074 11007 5083
rect 11059 5074 11207 5083
rect 11259 5074 11274 5126
rect 11326 5074 11341 5126
rect 11393 5074 11399 5126
rect 11455 5120 11507 5126
rect 11597 5074 11603 5126
rect 11655 5074 11670 5126
rect 11722 5074 11737 5126
rect 11789 5117 11965 5126
rect 11791 5083 11832 5117
rect 11866 5083 11907 5117
rect 11941 5083 11965 5117
rect 11789 5074 11965 5083
rect 12017 5074 12029 5126
rect 12081 5117 12093 5126
rect 12145 5117 12157 5126
rect 12209 5117 12221 5126
rect 12273 5117 12399 5126
rect 12451 5117 12495 5126
rect 12091 5083 12093 5117
rect 12273 5083 12282 5117
rect 12316 5083 12357 5117
rect 12391 5083 12399 5117
rect 12466 5083 12495 5117
rect 12081 5074 12093 5083
rect 12145 5074 12157 5083
rect 12209 5074 12221 5083
rect 12273 5074 12399 5083
rect 12451 5074 12495 5083
rect 12547 5074 12553 5126
rect 9511 5072 9536 5074
tri 9536 5072 9538 5074 nw
rect 4829 4990 4835 5024
rect 4869 4990 4892 5014
rect 4829 4964 4892 4990
rect 4829 4952 4840 4964
rect 4829 4918 4835 4952
rect 4829 4912 4840 4918
rect 4829 4906 4892 4912
rect 9459 5038 9511 5051
tri 9511 5047 9536 5072 nw
tri 9600 5032 9614 5046 se
rect 9614 5032 10323 5046
tri 9568 5000 9600 5032 se
rect 9600 5000 10323 5032
tri 9566 4998 9568 5000 se
rect 9568 4998 9632 5000
tri 9632 4998 9634 5000 nw
tri 10243 4998 10245 5000 ne
rect 10245 4998 10323 5000
rect 9459 4973 9468 4986
rect 9502 4973 9511 4986
tri 9548 4980 9566 4998 se
rect 9566 4980 9614 4998
tri 9614 4980 9632 4998 nw
tri 10245 4980 10263 4998 ne
rect 10263 4980 10323 4998
rect 9459 4908 9468 4921
rect 9502 4908 9511 4921
tri 4972 4887 4980 4895 se
tri 4969 4884 4972 4887 se
rect 4972 4884 4980 4887
tri 4955 4870 4969 4884 se
rect 4969 4870 4980 4884
rect 4637 4842 4689 4859
rect 3070 4753 3079 4759
rect 3113 4753 3122 4759
rect 3070 4744 3122 4753
tri 3220 4743 3229 4752 ne
rect 3229 4743 3300 4752
rect 3878 4738 3884 4790
rect 3936 4738 3948 4790
rect 4000 4738 4012 4790
rect 4064 4738 4070 4790
rect 4637 4773 4689 4790
rect 4637 4715 4689 4721
rect 4749 4864 4980 4870
rect 4801 4820 4980 4864
rect 9459 4843 9468 4856
rect 9502 4843 9511 4856
rect 4801 4812 4812 4820
rect 4749 4806 4812 4812
tri 4812 4806 4826 4820 nw
rect 4749 4801 4807 4806
tri 4807 4801 4812 4806 nw
rect 4749 4779 4801 4801
tri 4801 4795 4807 4801 nw
rect 9459 4786 9511 4791
rect 3070 4677 3079 4692
rect 3113 4690 3122 4692
tri 3122 4690 3144 4712 sw
tri 4727 4690 4749 4712 se
rect 4749 4693 4801 4727
rect 3113 4687 3144 4690
tri 3144 4687 3147 4690 sw
tri 4724 4687 4727 4690 se
rect 4727 4687 4749 4690
rect 3113 4677 4749 4687
rect 3122 4641 4749 4677
rect 3122 4635 4801 4641
rect 4829 4777 4892 4783
rect 4829 4771 4840 4777
rect 4829 4737 4835 4771
rect 4829 4725 4840 4737
rect 4829 4708 4892 4725
rect 4829 4690 4840 4708
rect 4829 4656 4835 4690
rect 4829 4639 4892 4656
rect 3070 4610 3079 4625
rect 3113 4610 3122 4625
tri 3122 4610 3147 4635 nw
rect 4829 4610 4840 4639
rect 1792 4517 1794 4525
tri 1794 4517 1802 4525 sw
tri 2468 4517 2476 4525 se
rect 2476 4517 2527 4525
rect 2566 4517 2572 4569
rect 2624 4517 2636 4569
rect 2688 4517 2882 4569
rect 4565 4595 4689 4607
rect 4565 4586 4574 4595
rect 4608 4586 4646 4595
rect 4680 4586 4689 4595
tri 3220 4575 3229 4584 se
rect 3229 4575 3300 4584
rect 3070 4543 3079 4558
rect 3113 4543 3122 4558
rect 4617 4534 4637 4586
rect 4565 4528 4689 4534
rect 4829 4576 4835 4610
rect 4869 4576 4892 4587
rect 4829 4570 4892 4576
rect 4829 4530 4840 4570
rect 1792 4502 1802 4517
tri 1802 4502 1817 4517 sw
tri 2453 4502 2468 4517 se
rect 2468 4502 2527 4517
rect 1792 4188 2527 4502
rect 3070 4482 3122 4491
rect 3070 4476 3079 4482
rect 3113 4476 3122 4482
rect 4829 4496 4835 4530
rect 4869 4501 4892 4518
rect 2830 4404 2882 4410
tri 2789 4336 2817 4364 ne
rect 2817 4352 2830 4364
rect 2817 4340 2882 4352
rect 2817 4336 2830 4340
tri 2817 4332 2821 4336 ne
rect 2821 4332 2830 4336
tri 2821 4328 2825 4332 ne
rect 2825 4328 2830 4332
tri 2825 4323 2830 4328 ne
rect 2830 4282 2882 4288
rect 3070 4408 3122 4424
rect 3070 4340 3122 4356
rect 3784 4417 4180 4461
rect 3784 4416 3865 4417
tri 3865 4416 3866 4417 nw
tri 4100 4416 4101 4417 ne
rect 4101 4416 4180 4417
rect 3784 4402 3851 4416
tri 3851 4402 3865 4416 nw
tri 4101 4402 4115 4416 ne
rect 4115 4402 4180 4416
rect 4829 4450 4840 4496
rect 4829 4416 4835 4450
rect 4869 4432 4892 4449
rect 3784 4389 3838 4402
tri 3838 4389 3851 4402 nw
tri 4115 4389 4128 4402 ne
rect 4128 4389 4180 4402
tri 3220 4310 3229 4319 ne
rect 3229 4310 3300 4319
rect 3070 4282 3122 4288
tri 3770 4265 3784 4279 se
rect 3784 4265 3826 4389
tri 3826 4377 3838 4389 nw
rect 3878 4337 3884 4389
rect 3936 4337 3948 4389
rect 4000 4337 4012 4389
rect 4064 4337 4084 4389
tri 4128 4383 4134 4389 ne
tri 3764 4259 3770 4265 se
rect 3770 4259 3826 4265
rect 4134 4332 4180 4389
rect 4637 4408 4689 4414
rect 4637 4342 4689 4356
rect 4134 4298 4140 4332
rect 4174 4298 4180 4332
tri 4130 4259 4134 4263 se
rect 4134 4259 4180 4298
tri 3759 4254 3764 4259 se
rect 3764 4254 3826 4259
rect 2882 4208 3826 4254
tri 4100 4229 4130 4259 se
rect 4130 4229 4140 4259
tri 2894 4188 2914 4208 ne
rect 2914 4188 2970 4208
tri 2970 4188 2990 4208 nw
tri 3759 4188 3779 4208 ne
rect 3779 4188 3826 4208
rect 1792 4186 1815 4188
tri 1815 4186 1817 4188 nw
tri 2453 4186 2455 4188 ne
rect 2455 4186 2527 4188
tri 2914 4186 2916 4188 ne
rect 2916 4186 2968 4188
tri 2968 4186 2970 4188 nw
tri 3779 4186 3781 4188 ne
rect 3781 4186 3826 4188
rect 1792 4183 1812 4186
tri 1812 4183 1815 4186 nw
tri 2455 4183 2458 4186 ne
rect 2458 4183 2527 4186
tri 2916 4183 2919 4186 ne
rect 1792 4168 1797 4183
tri 1797 4168 1812 4183 nw
tri 2458 4168 2473 4183 ne
rect 2473 4168 2527 4183
tri 1792 4163 1797 4168 nw
tri 2473 4163 2478 4168 ne
rect 1663 4129 1669 4163
rect 1703 4129 1709 4163
rect 1663 4089 1709 4129
rect 1820 4091 2032 4143
rect 2084 4091 2096 4143
rect 2148 4091 2160 4143
rect 2212 4091 2224 4143
rect 2276 4091 2288 4143
rect 2340 4091 2403 4143
rect 1663 4055 1669 4089
rect 1703 4055 1709 4089
rect 1663 4015 1709 4055
rect 1663 3981 1669 4015
rect 1703 3981 1709 4015
rect 1663 3941 1709 3981
rect 1663 3907 1669 3941
rect 1703 3907 1709 3941
rect 1663 3867 1709 3907
rect 1663 3833 1669 3867
rect 1703 3833 1709 3867
rect 1663 3793 1709 3833
rect 1663 3759 1669 3793
rect 1703 3759 1709 3793
rect 1663 3719 1709 3759
rect 1663 3685 1669 3719
rect 1703 3685 1709 3719
tri 1792 4058 1805 4071 sw
tri 2465 4058 2478 4071 se
rect 2478 4058 2527 4168
tri 2825 4134 2830 4139 se
rect 2830 4134 2882 4139
tri 2819 4128 2825 4134 se
rect 2825 4133 2882 4134
rect 2825 4128 2830 4133
tri 2804 4113 2819 4128 se
rect 2819 4113 2830 4128
rect 1792 4054 1805 4058
tri 1805 4054 1809 4058 sw
tri 2461 4054 2465 4058 se
rect 2465 4054 2527 4058
rect 1792 4046 1809 4054
tri 1809 4046 1817 4054 sw
tri 2453 4046 2461 4054 se
rect 2461 4046 2527 4054
rect 1792 3885 2527 4046
tri 2789 4098 2804 4113 se
rect 2804 4098 2830 4113
rect 2789 4081 2830 4098
rect 2789 4069 2882 4081
rect 2789 4052 2830 4069
tri 2789 4040 2801 4052 ne
rect 2801 4040 2830 4052
tri 2801 4017 2824 4040 ne
rect 2824 4017 2830 4040
tri 2824 4011 2830 4017 ne
rect 2830 4011 2882 4017
tri 2898 3946 2919 3967 se
rect 2919 3946 2965 4186
tri 2965 4183 2968 4186 nw
tri 3781 4183 3784 4186 ne
rect 3784 4183 3826 4186
rect 4084 4225 4140 4229
rect 4174 4225 4180 4259
rect 4084 4186 4180 4225
rect 4084 4183 4140 4186
tri 4100 4180 4103 4183 ne
rect 4103 4180 4140 4183
tri 2896 3944 2898 3946 se
rect 2898 3944 2965 3946
tri 2894 3942 2896 3944 se
rect 2896 3942 2965 3944
rect 2608 3936 2842 3942
rect 2608 3902 2620 3936
rect 2654 3902 2692 3936
rect 2726 3902 2764 3936
rect 2798 3902 2842 3936
rect 2608 3896 2842 3902
rect 2843 3897 2844 3941
rect 2880 3897 2881 3941
rect 2882 3896 2965 3942
rect 3070 4174 3122 4180
tri 4103 4159 4124 4180 ne
rect 4124 4159 4140 4180
tri 3226 4156 3229 4159 se
rect 3229 4156 3300 4159
tri 3222 4152 3226 4156 se
rect 3226 4152 3300 4156
tri 4124 4152 4131 4159 ne
rect 4131 4152 4140 4159
rect 4174 4152 4180 4186
rect 4258 4336 4310 4342
rect 4258 4234 4310 4284
rect 4258 4176 4310 4182
rect 4637 4275 4646 4290
rect 4680 4275 4689 4290
rect 4637 4208 4689 4223
rect 4829 4380 4840 4416
rect 4829 4370 4892 4380
rect 9459 4778 9468 4786
rect 9502 4778 9511 4786
rect 9459 4713 9511 4726
rect 9459 4648 9511 4661
rect 9459 4583 9511 4596
rect 9459 4518 9511 4531
rect 9459 4460 9468 4466
rect 9502 4460 9511 4466
rect 9459 4453 9511 4460
rect 9459 4388 9468 4401
rect 9502 4388 9511 4401
rect 6892 4373 6902 4374
rect 4829 4336 4835 4370
rect 4869 4362 4892 4370
rect 4829 4310 4840 4336
rect 6774 4321 6780 4373
rect 6832 4321 6844 4373
rect 6896 4321 6902 4373
rect 6892 4316 6902 4321
rect 9459 4323 9468 4336
rect 9502 4323 9511 4336
rect 4829 4292 4892 4310
rect 4829 4290 4840 4292
rect 4829 4256 4835 4290
rect 4829 4240 4840 4256
rect 4829 4222 4892 4240
rect 4829 4210 4840 4222
rect 4829 4176 4835 4210
rect 4829 4170 4840 4176
rect 4829 4164 4892 4170
rect 9459 4258 9468 4271
rect 9502 4258 9511 4271
rect 9459 4202 9511 4206
rect 9459 4193 9468 4202
rect 9502 4193 9511 4202
tri 3220 4150 3222 4152 se
rect 3222 4150 3300 4152
tri 4131 4150 4133 4152 ne
rect 4133 4150 4180 4152
tri 4133 4149 4134 4150 ne
rect 3070 4100 3122 4122
rect 4134 4148 4180 4150
tri 4180 4148 4188 4156 sw
rect 4637 4150 4689 4156
tri 9265 4150 9268 4153 se
tri 9263 4148 9265 4150 se
rect 9265 4148 9268 4150
rect 4134 4139 4188 4148
tri 4188 4139 4197 4148 sw
tri 9254 4139 9263 4148 se
rect 9263 4139 9268 4148
rect 4134 4128 4197 4139
tri 4197 4128 4208 4139 sw
tri 9243 4128 9254 4139 se
rect 9254 4128 9268 4139
rect 4134 4122 4208 4128
tri 4208 4122 4214 4128 sw
tri 9237 4122 9243 4128 se
rect 9243 4122 9268 4128
rect 9459 4128 9511 4141
rect 4134 4116 4230 4122
rect 4134 4113 4178 4116
rect 4134 4079 4140 4113
rect 4174 4079 4178 4113
rect 3070 4027 3122 4048
rect 3878 4021 3884 4073
rect 3936 4021 3948 4073
rect 4000 4021 4012 4073
rect 4064 4021 4084 4073
rect 4134 4064 4178 4079
rect 4134 4052 4230 4064
tri 9241 4054 9251 4064 ne
rect 9251 4054 9268 4064
rect 4134 4040 4178 4052
rect 4134 4006 4140 4040
rect 4174 4006 4178 4040
rect 4134 4000 4178 4006
tri 9251 4037 9268 4054 ne
rect 9459 4063 9511 4076
rect 4134 3994 4230 4000
rect 4637 4030 4689 4036
rect 3070 3954 3122 3975
rect 9459 3998 9511 4011
rect 4637 3963 4689 3978
tri 4086 3917 4098 3929 se
rect 4098 3923 4150 3929
rect 3070 3896 3122 3902
tri 3220 3893 3221 3894 ne
rect 3221 3893 3300 3894
tri 2527 3885 2535 3893 sw
tri 3221 3885 3229 3893 ne
rect 3229 3885 3300 3893
rect 1792 3874 2535 3885
tri 2535 3874 2546 3885 sw
rect 1792 3872 2546 3874
tri 2546 3872 2548 3874 sw
rect 1792 3868 2548 3872
tri 2548 3868 2552 3872 sw
rect 4084 3871 4098 3917
tri 4092 3868 4095 3871 ne
rect 4095 3868 4150 3871
rect 1792 3864 3096 3868
tri 3096 3864 3100 3868 sw
tri 4095 3865 4098 3868 ne
rect 4098 3865 4150 3868
rect 4637 3910 4646 3911
rect 4680 3910 4689 3911
rect 4637 3896 4689 3910
rect 1792 3840 3100 3864
tri 3100 3840 3124 3864 sw
rect 1792 3837 3124 3840
tri 3124 3837 3127 3840 sw
rect 1792 3831 4470 3837
rect 1792 3814 4418 3831
rect 1792 3798 2536 3814
tri 2536 3798 2552 3814 nw
tri 3071 3798 3087 3814 ne
rect 3087 3798 4418 3814
rect 1792 3732 2527 3798
tri 2527 3789 2536 3798 nw
tri 3087 3791 3094 3798 ne
rect 3094 3791 4418 3798
tri 4385 3789 4387 3791 ne
rect 4387 3789 4418 3791
tri 4387 3786 4390 3789 ne
rect 4390 3786 4418 3789
rect 2830 3780 2882 3786
tri 4390 3785 4391 3786 ne
rect 4391 3785 4418 3786
rect 1792 3709 1794 3732
tri 1794 3709 1817 3732 nw
tri 2453 3709 2476 3732 ne
rect 2476 3709 2527 3732
tri 2789 3709 2820 3740 ne
rect 2820 3728 2830 3740
tri 4391 3763 4413 3785 ne
rect 4413 3779 4418 3785
rect 4413 3767 4470 3779
rect 4413 3763 4418 3767
rect 2820 3716 2882 3728
rect 2820 3709 2830 3716
tri 1792 3707 1794 3709 nw
tri 2476 3707 2478 3709 ne
rect 1663 3646 1709 3685
rect 1663 3612 1669 3646
rect 1703 3612 1709 3646
rect 1820 3635 2032 3687
rect 2084 3635 2096 3687
rect 2148 3635 2160 3687
rect 2212 3635 2224 3687
rect 2276 3635 2288 3687
rect 2340 3635 2403 3687
rect 1663 3573 1709 3612
rect 1663 3539 1669 3573
rect 1703 3539 1709 3573
rect 1663 3500 1709 3539
rect 1663 3466 1669 3500
rect 1703 3466 1709 3500
rect 1663 3427 1709 3466
rect 1663 3393 1669 3427
rect 1703 3393 1709 3427
rect 1663 3354 1709 3393
rect 1663 3320 1669 3354
rect 1703 3320 1709 3354
rect 1663 3281 1709 3320
rect 1663 3247 1669 3281
rect 1703 3247 1709 3281
tri 1792 3612 1795 3615 sw
tri 2475 3612 2478 3615 se
rect 2478 3612 2527 3709
tri 2820 3706 2823 3709 ne
rect 2823 3706 2830 3709
tri 2823 3699 2830 3706 ne
rect 2830 3658 2882 3664
rect 3070 3749 3122 3755
rect 3878 3711 3884 3763
rect 3936 3711 3948 3763
rect 4000 3711 4012 3763
rect 4064 3711 4084 3763
tri 4413 3758 4418 3763 ne
rect 4258 3749 4310 3755
rect 2910 3653 2962 3659
tri 2909 3645 2910 3646 se
tri 2899 3635 2909 3645 se
rect 2909 3635 2910 3645
tri 2882 3618 2899 3635 se
rect 2899 3618 2910 3635
rect 1792 3590 1795 3612
tri 1795 3590 1817 3612 sw
tri 2453 3590 2475 3612 se
rect 2475 3590 2527 3612
rect 1792 3276 2527 3590
rect 2608 3612 2910 3618
rect 2608 3578 2620 3612
rect 2654 3578 2692 3612
rect 2726 3578 2764 3612
rect 2798 3578 2836 3612
rect 2870 3601 2910 3612
rect 2870 3589 2962 3601
rect 2870 3578 2910 3589
rect 2608 3572 2910 3578
tri 2882 3556 2898 3572 ne
rect 2898 3556 2910 3572
tri 2898 3548 2906 3556 ne
rect 2906 3548 2910 3556
tri 2906 3544 2910 3548 ne
rect 2910 3531 2962 3537
rect 3070 3654 3122 3697
rect 4418 3709 4470 3715
rect 4637 3830 4646 3844
rect 4680 3830 4689 3844
rect 4637 3829 4689 3830
rect 4637 3762 4646 3777
rect 4680 3762 4689 3777
rect 4749 3990 4801 3996
rect 4749 3924 4801 3938
rect 9214 3938 9329 3939
tri 9329 3938 9330 3939 nw
tri 9214 3926 9226 3938 ne
rect 9226 3926 9317 3938
tri 9317 3926 9329 3938 nw
rect 9459 3933 9511 3946
tri 9226 3909 9243 3926 ne
tri 4801 3872 4803 3874 sw
tri 9241 3872 9243 3874 se
rect 9243 3872 9300 3926
tri 9300 3909 9317 3926 nw
rect 4749 3858 4803 3872
rect 4801 3852 4803 3858
tri 4803 3852 4823 3872 sw
tri 9221 3852 9241 3872 se
rect 9241 3852 9300 3872
rect 4801 3840 4823 3852
tri 4823 3840 4835 3852 sw
tri 9209 3840 9221 3852 se
rect 9221 3840 9300 3852
rect 4801 3806 9300 3840
rect 4749 3791 9300 3806
rect 4801 3782 9300 3791
rect 9459 3872 9468 3881
rect 9502 3872 9511 3881
rect 9459 3868 9511 3872
rect 9459 3804 9468 3816
rect 9502 3804 9511 3816
rect 4801 3778 4831 3782
tri 4831 3778 4835 3782 nw
rect 4801 3777 4830 3778
tri 4830 3777 4831 3778 nw
rect 4801 3759 4812 3777
tri 4812 3759 4830 3777 nw
tri 9441 3759 9459 3777 se
rect 4801 3758 4811 3759
tri 4811 3758 4812 3759 nw
tri 9440 3758 9441 3759 se
rect 9441 3758 9459 3759
tri 4801 3748 4811 3758 nw
tri 9434 3752 9440 3758 se
rect 9440 3752 9459 3758
rect 4749 3733 4801 3739
rect 5037 3747 7393 3752
rect 5037 3746 5163 3747
rect 5215 3746 5230 3747
rect 5282 3746 5297 3747
rect 5349 3746 5364 3747
rect 5416 3746 5431 3747
rect 5483 3746 5498 3747
rect 5550 3746 5565 3747
rect 5617 3746 5632 3747
rect 5684 3746 5699 3747
rect 5751 3746 5766 3747
rect 5818 3746 5834 3747
rect 5886 3746 5902 3747
rect 5954 3746 5970 3747
rect 6022 3746 6142 3747
rect 6706 3746 6719 3747
rect 6771 3746 6784 3747
rect 6836 3746 6849 3747
rect 6901 3746 7393 3747
rect 7445 3746 7461 3752
rect 7513 3746 7529 3752
rect 7581 3746 7598 3752
rect 7650 3746 7667 3752
rect 7719 3746 7736 3752
rect 7788 3746 7805 3752
rect 7857 3746 7874 3752
rect 7926 3746 7943 3752
rect 7995 3746 8012 3752
rect 8064 3746 8187 3752
rect 8239 3746 8255 3752
rect 8307 3746 8323 3752
rect 8375 3746 8391 3752
rect 8443 3746 8459 3752
rect 8511 3746 8528 3752
rect 8580 3746 8597 3752
rect 8649 3746 8666 3752
rect 8718 3746 8735 3752
rect 8787 3746 8804 3752
rect 8856 3746 8873 3752
rect 8925 3746 8942 3752
rect 8994 3746 9011 3752
rect 4258 3654 4310 3697
tri 4070 3611 4098 3639 se
rect 4098 3638 4150 3644
tri 4064 3605 4070 3611 se
rect 4070 3605 4098 3611
rect 3070 3560 3122 3602
rect 4084 3586 4098 3605
rect 4084 3574 4150 3586
rect 4084 3559 4098 3574
tri 4064 3556 4067 3559 ne
rect 4067 3556 4098 3559
tri 4067 3548 4075 3556 ne
rect 4075 3548 4098 3556
tri 2829 3514 2830 3515 se
rect 2830 3514 2882 3515
tri 2817 3502 2829 3514 se
rect 2829 3509 2882 3514
rect 2829 3502 2830 3509
tri 2797 3482 2817 3502 se
rect 2817 3482 2830 3502
tri 2789 3474 2797 3482 se
rect 2797 3474 2830 3482
rect 2789 3457 2830 3474
tri 4075 3530 4093 3548 ne
rect 4093 3530 4098 3548
tri 3220 3520 3230 3530 ne
rect 3230 3520 3300 3530
tri 4093 3525 4098 3530 ne
rect 4098 3516 4150 3522
rect 4258 3560 4310 3602
rect 3070 3502 3122 3508
rect 4258 3502 4310 3508
rect 4637 3706 4689 3710
rect 4637 3695 4646 3706
rect 4680 3695 4689 3706
rect 4637 3628 4689 3643
tri 5018 3640 5037 3659 se
rect 5037 3640 5049 3746
rect 8994 3712 9010 3746
rect 8994 3700 9011 3712
rect 9063 3700 9080 3752
rect 9132 3746 9468 3752
rect 9132 3712 9156 3746
rect 9190 3712 9229 3746
rect 9263 3712 9302 3746
rect 9336 3712 9375 3746
rect 9409 3740 9468 3746
rect 9502 3740 9511 3752
rect 9409 3712 9459 3740
rect 9132 3700 9459 3712
rect 8971 3688 9459 3700
rect 8994 3674 9011 3688
rect 8994 3640 9010 3674
rect 5012 3631 5163 3640
rect 5215 3631 5230 3640
rect 5282 3631 5297 3640
rect 5349 3631 5364 3640
rect 5416 3631 5431 3640
rect 5483 3631 5498 3640
rect 5550 3631 5565 3640
rect 5617 3631 5632 3640
rect 5684 3631 5699 3640
rect 5751 3631 5766 3640
rect 5818 3631 5834 3640
rect 5886 3631 5902 3640
rect 5954 3631 5970 3640
rect 6022 3631 6142 3640
rect 6706 3631 6719 3640
rect 6771 3631 6784 3640
rect 6836 3631 6849 3640
rect 6901 3636 7393 3640
rect 7445 3636 7461 3640
rect 7513 3636 7529 3640
rect 7581 3636 7598 3640
rect 7650 3636 7667 3640
rect 7719 3636 7736 3640
rect 7788 3636 7805 3640
rect 7857 3636 7874 3640
rect 7926 3636 7943 3640
rect 7995 3636 8012 3640
rect 8064 3636 8187 3640
rect 8239 3636 8255 3640
rect 8307 3636 8323 3640
rect 8375 3636 8391 3640
rect 8443 3636 8459 3640
rect 8511 3636 8528 3640
rect 8580 3636 8597 3640
rect 8649 3636 8666 3640
rect 8718 3636 8735 3640
rect 8787 3636 8804 3640
rect 8856 3636 8873 3640
rect 8925 3636 8942 3640
rect 8994 3636 9011 3640
rect 9063 3636 9080 3688
rect 9132 3684 9511 3688
rect 9132 3676 9468 3684
rect 9502 3676 9511 3684
rect 9132 3674 9459 3676
rect 9132 3640 9156 3674
rect 9190 3640 9229 3674
rect 9263 3640 9302 3674
rect 9336 3640 9375 3674
rect 9409 3640 9459 3674
rect 9132 3636 9459 3640
rect 6901 3634 9459 3636
rect 6901 3631 7035 3634
rect 5012 3630 7035 3631
tri 7035 3630 7039 3634 nw
tri 9434 3630 9438 3634 ne
rect 9438 3630 9459 3634
rect 5012 3615 7020 3630
tri 7020 3615 7035 3630 nw
tri 9438 3615 9453 3630 ne
rect 9453 3624 9459 3630
rect 9453 3615 9511 3624
rect 5012 3610 7015 3615
tri 7015 3610 7020 3615 nw
tri 9453 3610 9458 3615 ne
rect 9458 3612 9511 3615
rect 9458 3610 9459 3612
rect 5012 3588 7014 3610
tri 7014 3609 7015 3610 nw
tri 9458 3609 9459 3610 ne
rect 5013 3586 7013 3587
rect 4637 3560 4689 3576
rect 4637 3502 4689 3508
rect 5013 3549 7013 3550
rect 7014 3548 7033 3550
rect 9459 3548 9511 3560
rect 5012 3496 6911 3548
rect 6963 3496 6975 3548
rect 7027 3496 7033 3548
rect 7203 3496 7209 3548
rect 7261 3496 7273 3548
rect 7325 3496 9282 3548
rect 9459 3490 9511 3496
tri 9540 4972 9548 4980 se
rect 9548 4972 9606 4980
tri 9606 4972 9614 4980 nw
tri 10263 4972 10271 4980 ne
rect 10271 4972 10323 4980
rect 9540 4961 9595 4972
tri 9595 4961 9606 4972 nw
rect 10143 4966 10195 4972
tri 10271 4966 10277 4972 ne
rect 9540 4958 9592 4961
tri 9592 4958 9595 4961 nw
tri 10140 4958 10143 4961 se
rect 2789 3445 2882 3457
tri 9518 3447 9540 3469 se
rect 9540 3447 9586 4958
tri 9586 4952 9592 4958 nw
tri 10134 4952 10140 4958 se
rect 10140 4952 10143 4958
tri 10109 4927 10134 4952 se
rect 10134 4927 10143 4952
rect 9694 4921 9824 4927
rect 9694 4887 9706 4921
rect 9740 4887 9778 4921
rect 9812 4887 9824 4921
rect 9694 4881 9824 4887
rect 9928 4921 10143 4927
rect 9928 4887 9942 4921
rect 9976 4887 10014 4921
rect 10048 4914 10143 4921
rect 10048 4902 10195 4914
rect 10048 4887 10143 4902
rect 9928 4881 10143 4887
tri 9698 4852 9727 4881 ne
rect 9727 4852 9789 4881
tri 9789 4852 9818 4881 nw
rect 2789 3428 2830 3445
tri 2789 3408 2809 3428 ne
rect 2809 3408 2830 3428
tri 2809 3399 2818 3408 ne
rect 2818 3399 2830 3408
tri 2818 3396 2821 3399 ne
rect 2821 3396 2830 3399
tri 2821 3388 2829 3396 ne
rect 2829 3393 2830 3396
tri 9514 3443 9518 3447 se
rect 9518 3443 9586 3447
rect 2829 3388 2882 3393
tri 2829 3387 2830 3388 ne
rect 2830 3387 2882 3388
rect 3070 3394 3122 3400
rect 4637 3394 4689 3400
tri 3238 3388 3241 3391 se
rect 3241 3388 3306 3391
tri 2905 3354 2910 3359 se
rect 2910 3354 2962 3359
tri 2901 3350 2905 3354 se
rect 2905 3353 2962 3354
rect 2905 3350 2910 3353
tri 2898 3347 2901 3350 se
rect 2901 3347 2910 3350
tri 2869 3318 2898 3347 se
rect 2898 3318 2910 3347
rect 1792 3272 1813 3276
tri 1813 3272 1817 3276 nw
tri 2453 3272 2457 3276 ne
rect 2457 3272 2527 3276
rect 2608 3312 2829 3318
rect 2608 3278 2620 3312
rect 2654 3278 2692 3312
rect 2726 3278 2764 3312
rect 2798 3278 2829 3312
rect 2608 3272 2829 3278
rect 2830 3273 2831 3317
rect 2867 3273 2868 3317
rect 2869 3301 2910 3318
rect 2869 3289 2962 3301
rect 2869 3272 2910 3289
rect 1792 3268 1809 3272
tri 1809 3268 1813 3272 nw
tri 2457 3268 2461 3272 ne
rect 2461 3268 2527 3272
tri 2869 3268 2873 3272 ne
rect 2873 3268 2910 3272
tri 1792 3251 1809 3268 nw
tri 2461 3251 2478 3268 ne
rect 1663 3208 1709 3247
rect 1663 3174 1669 3208
rect 1703 3174 1709 3208
rect 1820 3179 2032 3231
rect 2084 3179 2096 3231
rect 2148 3179 2160 3231
rect 2212 3179 2224 3231
rect 2276 3179 2288 3231
rect 2340 3179 2403 3231
rect 1663 3135 1709 3174
rect 1663 3101 1669 3135
rect 1703 3101 1709 3135
rect 1663 3062 1709 3101
rect 1663 3028 1669 3062
rect 1703 3028 1709 3062
rect 1663 2989 1709 3028
rect 1663 2955 1669 2989
rect 1703 2955 1709 2989
rect 1663 2943 1709 2955
tri 1792 3143 1808 3159 sw
tri 2462 3143 2478 3159 se
rect 2478 3143 2527 3268
tri 2873 3241 2900 3268 ne
rect 2900 3241 2910 3268
tri 2900 3239 2902 3241 ne
rect 2902 3239 2910 3241
tri 2902 3231 2910 3239 ne
rect 2910 3231 2962 3237
tri 3237 3387 3238 3388 se
rect 3238 3387 3306 3388
tri 3220 3370 3237 3387 se
rect 3237 3370 3306 3387
rect 3070 3323 3122 3342
rect 3070 3268 3079 3271
rect 3113 3268 3122 3271
rect 3070 3253 3122 3268
rect 3544 3347 3884 3359
rect 3544 3313 3550 3347
rect 3584 3313 3884 3347
rect 3544 3307 3884 3313
rect 3936 3307 3948 3359
rect 4000 3307 4012 3359
rect 4064 3307 4070 3359
rect 4637 3318 4689 3342
rect 3544 3275 3636 3307
tri 3636 3275 3668 3307 nw
rect 4258 3279 4310 3285
rect 3544 3241 3550 3275
rect 3584 3273 3634 3275
tri 3634 3273 3636 3275 nw
rect 3584 3260 3621 3273
tri 3621 3260 3634 3273 nw
rect 3584 3241 3600 3260
rect 3544 3239 3600 3241
tri 3600 3239 3621 3260 nw
rect 3544 3238 3599 3239
tri 3599 3238 3600 3239 nw
rect 3544 3231 3592 3238
tri 3592 3231 3599 3238 nw
rect 3544 3230 3591 3231
tri 3591 3230 3592 3231 nw
rect 3544 3229 3590 3230
tri 3590 3229 3591 3230 nw
tri 2809 3182 2830 3203 se
rect 2830 3197 2882 3203
tri 2806 3179 2809 3182 se
rect 2809 3179 2830 3182
tri 2793 3166 2806 3179 se
rect 2806 3166 2830 3179
rect 1792 3135 1808 3143
tri 1808 3135 1816 3143 sw
tri 2454 3135 2462 3143 se
rect 2462 3135 2527 3143
rect 1792 3134 1816 3135
tri 1816 3134 1817 3135 sw
tri 2453 3134 2454 3135 se
rect 2454 3134 2527 3135
rect 1792 3129 2527 3134
rect 1792 3077 2475 3129
tri 2789 3162 2793 3166 se
rect 2793 3162 2830 3166
rect 2789 3145 2830 3162
rect 2789 3133 2882 3145
rect 2789 3116 2830 3133
tri 2789 3097 2808 3116 ne
rect 2808 3097 2830 3116
tri 2808 3093 2812 3097 ne
rect 2812 3093 2830 3097
rect 1792 3065 2527 3077
tri 2812 3075 2830 3093 ne
rect 2830 3075 2882 3081
rect 3070 3183 3079 3201
rect 3113 3183 3122 3201
rect 4637 3242 4689 3266
rect 4258 3211 4310 3227
rect 3070 3113 3079 3131
rect 3113 3113 3122 3131
rect 3878 3103 3884 3155
rect 3936 3103 3948 3155
rect 4000 3103 4012 3155
rect 4064 3103 4084 3155
rect 4258 3143 4310 3159
rect 1792 3013 2475 3065
tri 4177 3093 4178 3094 se
rect 4178 3093 4230 3098
tri 4159 3075 4177 3093 se
rect 4177 3092 4230 3093
rect 4177 3075 4178 3092
tri 4154 3070 4159 3075 se
rect 4159 3070 4178 3075
rect 3070 3046 3122 3061
tri 4144 3060 4154 3070 se
rect 4154 3060 4178 3070
rect 3070 3043 3079 3046
rect 3113 3043 3122 3046
tri 2527 3014 2544 3031 sw
rect 2527 3013 2544 3014
rect 1792 3012 2544 3013
tri 2544 3012 2546 3014 sw
tri 3762 3036 3774 3048 se
rect 3774 3036 3820 3048
tri 3757 3031 3762 3036 se
rect 3762 3031 3780 3036
tri 3750 3024 3757 3031 se
rect 3757 3024 3780 3031
rect 1792 3006 2546 3012
tri 2546 3006 2552 3012 sw
rect 1792 3001 2608 3006
rect 1792 2949 2475 3001
rect 2527 2960 2608 3001
rect 3070 2973 3122 2991
rect 2527 2949 2532 2960
rect 1792 2943 2532 2949
tri 2532 2943 2549 2960 nw
rect 2910 2959 2962 2965
tri 557 2895 571 2909 ne
rect 571 2895 631 2909
tri 401 2885 411 2895 sw
tri 571 2885 581 2895 ne
rect 581 2885 631 2895
rect 329 2879 411 2885
tri 411 2879 417 2885 sw
tri 581 2879 587 2885 ne
rect 329 2866 417 2879
tri 417 2866 430 2879 sw
rect 329 2814 429 2866
rect 481 2814 493 2866
rect 545 2863 556 2866
tri 556 2863 559 2866 sw
rect 545 2857 559 2863
rect 547 2823 559 2857
rect 545 2817 559 2823
rect 545 2814 556 2817
tri 556 2814 559 2817 nw
rect 329 2804 490 2814
tri 490 2804 500 2814 nw
rect 329 2801 487 2804
tri 487 2801 490 2804 nw
rect 329 2799 485 2801
tri 485 2799 487 2801 nw
tri 585 2799 587 2801 se
rect 587 2799 631 2885
rect 958 2837 1010 2873
rect 1150 2870 1156 2922
rect 1208 2870 1220 2922
rect 1272 2870 1284 2922
rect 1336 2870 1352 2922
tri 2897 2927 2910 2940 se
tri 2892 2922 2897 2927 se
rect 2897 2922 2910 2927
tri 2885 2915 2892 2922 se
rect 2892 2915 2910 2922
rect 1471 2901 1523 2915
tri 1642 2904 1653 2915 se
rect 1653 2907 2910 2915
rect 1653 2904 2962 2907
tri 1613 2875 1642 2904 se
rect 1642 2895 2962 2904
rect 1642 2887 2910 2895
rect 1642 2875 1653 2887
tri 1653 2875 1665 2887 nw
tri 2885 2875 2897 2887 ne
rect 2897 2875 2910 2887
tri 1612 2874 1613 2875 se
rect 1613 2874 1652 2875
tri 1652 2874 1653 2875 nw
tri 2897 2874 2898 2875 ne
rect 2898 2874 2910 2875
tri 1608 2870 1612 2874 se
rect 1612 2870 1643 2874
tri 1603 2865 1608 2870 se
rect 1608 2865 1643 2870
tri 1643 2865 1652 2874 nw
tri 2898 2865 2907 2874 ne
rect 2907 2865 2910 2874
tri 1596 2858 1603 2865 se
rect 1603 2858 1636 2865
tri 1636 2858 1643 2865 nw
tri 2907 2862 2910 2865 ne
tri 1588 2850 1596 2858 se
rect 1596 2850 1628 2858
tri 1628 2850 1636 2858 nw
rect 1471 2843 1523 2849
tri 1581 2843 1588 2850 se
rect 1588 2843 1616 2850
tri 1576 2838 1581 2843 se
rect 1581 2838 1616 2843
tri 1616 2838 1628 2850 nw
rect 1746 2844 2527 2850
rect 1746 2838 2475 2844
tri 1575 2837 1576 2838 se
rect 1576 2837 1613 2838
tri 1573 2835 1575 2837 se
rect 1575 2835 1613 2837
tri 1613 2835 1616 2838 nw
tri 1547 2809 1573 2835 se
rect 1573 2809 1582 2835
rect 0 2787 273 2799
rect 0 2753 233 2787
rect 267 2753 273 2787
rect 0 2714 273 2753
rect 0 2680 233 2714
rect 267 2680 273 2714
rect 0 2641 273 2680
rect 0 2607 233 2641
rect 267 2607 273 2641
rect 0 2595 273 2607
rect 329 2797 483 2799
tri 483 2797 485 2799 nw
tri 583 2797 585 2799 se
rect 585 2797 631 2799
rect 329 2691 473 2797
tri 473 2787 483 2797 nw
tri 573 2787 583 2797 se
rect 583 2787 631 2797
tri 557 2771 573 2787 se
rect 573 2771 631 2787
rect 501 2765 631 2771
rect 501 2731 513 2765
rect 547 2731 585 2765
rect 619 2731 631 2765
rect 501 2725 631 2731
rect 687 2797 1150 2809
tri 1542 2804 1547 2809 se
rect 1547 2804 1582 2809
tri 1582 2804 1613 2835 nw
rect 1746 2804 1752 2838
rect 1786 2820 2475 2838
rect 1786 2804 1801 2820
tri 1801 2804 1817 2820 nw
tri 2450 2804 2466 2820 ne
rect 2466 2804 2475 2820
rect 2750 2844 2802 2850
tri 1539 2801 1542 2804 se
rect 1542 2801 1579 2804
tri 1579 2801 1582 2804 nw
rect 1746 2801 1798 2804
tri 1798 2801 1801 2804 nw
tri 2466 2801 2469 2804 ne
rect 2469 2801 2475 2804
rect 687 2763 693 2797
rect 727 2763 1052 2797
rect 1086 2763 1150 2797
tri 1533 2795 1539 2801 se
rect 1539 2795 1573 2801
tri 1573 2795 1579 2801 nw
tri 1525 2787 1533 2795 se
rect 1533 2787 1565 2795
tri 1565 2787 1573 2795 nw
tri 1504 2766 1525 2787 se
rect 1525 2766 1544 2787
tri 1544 2766 1565 2787 nw
rect 1746 2766 1792 2801
tri 1792 2795 1798 2801 nw
tri 2469 2795 2475 2801 ne
tri 2725 2801 2728 2804 ne
rect 2728 2801 2750 2804
rect 2475 2780 2527 2792
tri 2728 2787 2742 2801 ne
rect 2742 2792 2750 2801
rect 2910 2837 2962 2843
rect 2990 2940 3042 2946
rect 3590 3018 3780 3024
rect 3642 3002 3780 3018
rect 3814 3002 3820 3036
rect 4084 3040 4178 3060
rect 4084 3028 4230 3040
rect 4084 3014 4178 3028
rect 3642 2966 3820 3002
tri 4144 2994 4164 3014 ne
rect 4164 2994 4178 3014
tri 4164 2981 4177 2994 ne
rect 4177 2981 4178 2994
tri 4177 2980 4178 2981 ne
rect 4178 2970 4230 2976
rect 4418 3232 4470 3238
rect 4757 3399 9586 3443
rect 9617 4840 9663 4852
tri 9727 4850 9729 4852 ne
rect 9729 4850 9787 4852
tri 9787 4850 9789 4852 nw
tri 9729 4847 9732 4850 ne
rect 9617 4806 9623 4840
rect 9657 4806 9663 4840
rect 9617 4767 9663 4806
rect 9617 4733 9623 4767
rect 9657 4733 9663 4767
rect 9617 4694 9663 4733
rect 9732 4816 9784 4850
tri 9784 4847 9787 4850 nw
rect 9732 4752 9784 4764
rect 9732 4694 9784 4700
rect 9848 4840 9900 4852
rect 9848 4806 9859 4840
rect 9893 4806 9900 4840
rect 9848 4767 9900 4806
rect 9848 4733 9859 4767
rect 9893 4733 9900 4767
rect 9848 4694 9900 4733
rect 9617 4660 9623 4694
rect 9657 4660 9663 4694
rect 9617 4621 9663 4660
rect 9617 4587 9623 4621
rect 9657 4587 9663 4621
rect 9617 4548 9663 4587
rect 9617 4514 9623 4548
rect 9657 4514 9663 4548
rect 9617 4475 9663 4514
rect 9617 4441 9623 4475
rect 9657 4441 9663 4475
rect 9617 4402 9663 4441
rect 9617 4368 9623 4402
rect 9657 4368 9663 4402
rect 9617 4329 9663 4368
rect 9617 4295 9623 4329
rect 9657 4295 9663 4329
rect 9617 4256 9663 4295
rect 9617 4222 9623 4256
rect 9657 4222 9663 4256
rect 9617 4182 9663 4222
rect 9617 4148 9623 4182
rect 9657 4148 9663 4182
rect 9617 4108 9663 4148
rect 9617 4074 9623 4108
rect 9657 4074 9663 4108
rect 9617 4034 9663 4074
rect 9617 4000 9623 4034
rect 9657 4000 9663 4034
rect 9617 3960 9663 4000
rect 9617 3926 9623 3960
rect 9657 3926 9663 3960
rect 9617 3886 9663 3926
rect 9617 3852 9623 3886
rect 9657 3852 9663 3886
rect 9617 3812 9663 3852
rect 9617 3778 9623 3812
rect 9657 3778 9663 3812
rect 9617 3738 9663 3778
rect 9617 3704 9623 3738
rect 9657 3704 9663 3738
rect 9617 3664 9663 3704
rect 9617 3630 9623 3664
rect 9657 3630 9663 3664
rect 9617 3590 9663 3630
rect 9617 3556 9623 3590
rect 9657 3556 9663 3590
rect 9617 3516 9663 3556
rect 9617 3482 9623 3516
rect 9657 3482 9663 3516
rect 9617 3442 9663 3482
rect 9617 3408 9623 3442
rect 9657 3408 9663 3442
rect 4757 3396 4832 3399
tri 4832 3396 4835 3399 nw
rect 4757 3387 4823 3396
tri 4823 3387 4832 3396 nw
rect 4757 3373 4809 3387
tri 4809 3373 4823 3387 nw
rect 4757 3368 4804 3373
tri 4804 3368 4809 3373 nw
rect 9617 3368 9663 3408
rect 4637 3184 4689 3190
tri 4756 3189 4757 3190 se
rect 4757 3189 4801 3368
tri 4801 3365 4804 3368 nw
tri 9456 3359 9459 3362 se
rect 9459 3359 9511 3362
tri 9447 3350 9456 3359 se
rect 9456 3356 9511 3359
rect 9456 3350 9459 3356
tri 9442 3345 9447 3350 se
rect 9447 3345 9459 3350
tri 4755 3188 4756 3189 se
rect 4756 3188 4801 3189
tri 4753 3186 4755 3188 se
rect 4755 3186 4801 3188
tri 4751 3184 4753 3186 se
rect 4753 3184 4801 3186
tri 4750 3183 4751 3184 se
rect 4751 3183 4801 3184
tri 4748 3181 4750 3183 se
rect 4750 3181 4801 3183
rect 4418 3177 4470 3180
tri 4470 3177 4474 3181 sw
tri 4744 3177 4748 3181 se
rect 4748 3177 4801 3181
rect 4418 3168 4474 3177
rect 4470 3156 4474 3168
tri 4474 3156 4495 3177 sw
tri 4723 3156 4744 3177 se
rect 4744 3156 4801 3177
rect 4470 3116 4801 3156
rect 4418 3110 4801 3116
rect 4829 3339 4892 3345
tri 9440 3343 9442 3345 se
rect 9442 3343 9459 3345
rect 4829 3333 4840 3339
rect 4829 3299 4835 3333
tri 4892 3325 4910 3343 sw
tri 9422 3325 9440 3343 se
rect 9440 3325 9459 3343
rect 4892 3324 4910 3325
tri 4910 3324 4911 3325 sw
tri 9421 3324 9422 3325 se
rect 9422 3324 9459 3325
rect 4892 3316 4911 3324
tri 4911 3316 4919 3324 sw
tri 9413 3316 9421 3324 se
rect 9421 3316 9459 3324
rect 4892 3314 4919 3316
tri 4919 3314 4921 3316 sw
tri 9411 3314 9413 3316 se
rect 9413 3314 9459 3316
rect 4892 3312 4921 3314
tri 4921 3312 4923 3314 sw
rect 4829 3287 4840 3299
rect 4892 3287 6164 3312
rect 4829 3274 6164 3287
rect 4829 3255 4840 3274
rect 4892 3260 6164 3274
rect 6216 3260 6241 3312
rect 6293 3260 6318 3312
rect 6370 3260 6395 3312
rect 6447 3260 6471 3312
rect 6523 3260 7014 3312
rect 7280 3262 7400 3314
rect 7452 3262 7467 3314
rect 7519 3262 7534 3314
rect 7586 3262 7601 3314
rect 7653 3262 7668 3314
rect 7720 3262 7735 3314
rect 7787 3262 7802 3314
rect 7854 3262 7869 3314
rect 7921 3262 7936 3314
rect 7988 3262 8002 3314
rect 8054 3304 9459 3314
rect 8054 3272 9511 3304
rect 8054 3262 9459 3272
rect 7280 3260 9459 3262
rect 4829 3221 4835 3255
rect 4892 3238 4901 3260
tri 4901 3238 4923 3260 nw
tri 9413 3238 9435 3260 ne
rect 9435 3238 9459 3260
tri 4892 3229 4901 3238 nw
tri 9435 3229 9444 3238 ne
rect 9444 3229 9459 3238
tri 9444 3227 9446 3229 ne
rect 9446 3227 9459 3229
tri 9446 3225 9448 3227 ne
rect 9448 3225 9459 3227
rect 4869 3221 4892 3222
rect 4829 3209 4892 3221
tri 9448 3220 9453 3225 ne
rect 9453 3220 9459 3225
tri 9453 3214 9459 3220 ne
rect 9459 3214 9511 3220
rect 9617 3334 9623 3368
rect 9657 3334 9663 3368
rect 9617 3294 9663 3334
rect 9617 3260 9623 3294
rect 9657 3260 9663 3294
rect 9617 3220 9663 3260
rect 4829 3177 4840 3209
tri 5375 3186 5377 3188 se
rect 5377 3186 5383 3188
tri 5372 3183 5375 3186 se
rect 5375 3183 5383 3186
tri 5371 3182 5372 3183 se
rect 5372 3182 5383 3183
rect 4829 3143 4835 3177
rect 4869 3144 4892 3157
rect 4258 3075 4310 3091
rect 4829 3099 4840 3143
rect 5377 3136 5383 3182
rect 5435 3136 5447 3188
rect 5499 3186 5505 3188
tri 5505 3186 5507 3188 sw
rect 5499 3183 5507 3186
tri 5507 3183 5510 3186 sw
rect 5499 3182 5510 3183
tri 5510 3182 5511 3183 sw
rect 5499 3136 5505 3182
rect 7280 3137 8638 3189
rect 8690 3137 8702 3189
rect 8754 3137 9282 3189
rect 7280 3132 9282 3137
rect 9617 3186 9623 3220
rect 9657 3186 9663 3220
rect 9617 3154 9663 3186
rect 9848 4660 9859 4694
rect 9893 4660 9900 4694
rect 9848 4621 9900 4660
rect 9848 4587 9859 4621
rect 9893 4587 9900 4621
rect 9848 4548 9900 4587
rect 9848 4514 9859 4548
rect 9893 4514 9900 4548
rect 9848 4475 9900 4514
rect 9848 4441 9859 4475
rect 9893 4441 9900 4475
rect 9848 4402 9900 4441
rect 9848 4368 9859 4402
rect 9893 4368 9900 4402
rect 9928 4850 9983 4881
tri 9983 4850 10014 4881 nw
tri 10109 4850 10140 4881 ne
rect 10140 4850 10143 4881
rect 9928 4510 9980 4850
tri 9980 4847 9983 4850 nw
tri 10140 4847 10143 4850 ne
rect 10143 4844 10195 4850
rect 9928 4446 9980 4458
rect 9928 4388 9980 4394
rect 10089 4801 10135 4813
rect 10089 4767 10095 4801
rect 10129 4767 10135 4801
rect 10089 4729 10135 4767
rect 10089 4695 10095 4729
rect 10129 4695 10135 4729
rect 10089 4657 10135 4695
rect 10089 4623 10095 4657
rect 10129 4623 10135 4657
rect 10089 4585 10135 4623
rect 10089 4551 10095 4585
rect 10129 4551 10135 4585
rect 10089 4513 10135 4551
rect 10089 4479 10095 4513
rect 10129 4479 10135 4513
rect 10089 4441 10135 4479
rect 10089 4407 10095 4441
rect 10129 4407 10135 4441
rect 9848 4329 9900 4368
rect 9848 4295 9859 4329
rect 9893 4295 9900 4329
rect 9848 4256 9900 4295
rect 9848 4222 9859 4256
rect 9893 4222 9900 4256
rect 9848 4183 9900 4222
rect 9848 4149 9859 4183
rect 9893 4149 9900 4183
rect 9848 4110 9900 4149
rect 9848 4076 9859 4110
rect 9893 4076 9900 4110
rect 9848 4037 9900 4076
rect 9848 4003 9859 4037
rect 9893 4003 9900 4037
rect 9848 3964 9900 4003
rect 9848 3930 9859 3964
rect 9893 3930 9900 3964
rect 9848 3891 9900 3930
rect 9848 3857 9859 3891
rect 9893 3857 9900 3891
rect 9848 3817 9900 3857
rect 9848 3783 9859 3817
rect 9893 3783 9900 3817
rect 9848 3743 9900 3783
rect 9848 3709 9859 3743
rect 9893 3709 9900 3743
rect 9848 3669 9900 3709
rect 9848 3635 9859 3669
rect 9893 3635 9900 3669
rect 9848 3595 9900 3635
rect 9848 3561 9859 3595
rect 9893 3561 9900 3595
rect 9848 3521 9900 3561
rect 9848 3487 9859 3521
rect 9893 3487 9900 3521
rect 9848 3447 9900 3487
rect 9848 3413 9859 3447
rect 9893 3413 9900 3447
rect 9848 3407 9900 3413
rect 9848 3339 9859 3355
rect 9893 3339 9900 3355
rect 9848 3329 9900 3339
rect 9848 3265 9859 3277
rect 9893 3265 9900 3277
rect 9848 3250 9900 3265
rect 9848 3191 9859 3198
rect 9893 3191 9900 3198
rect 9848 3171 9900 3191
tri 9663 3154 9672 3163 sw
rect 9617 3148 9672 3154
rect 6958 3102 7092 3108
tri 6956 3100 6958 3102 se
rect 6958 3100 7040 3102
rect 4258 3020 4266 3023
rect 4300 3020 4310 3023
rect 4258 3008 4310 3020
rect 3590 2950 3820 2966
rect 3070 2915 3122 2921
tri 3220 2915 3227 2922 ne
rect 3227 2915 3306 2922
tri 3227 2907 3235 2915 ne
rect 3235 2907 3306 2915
tri 3235 2904 3238 2907 ne
rect 3238 2904 3306 2907
tri 3238 2901 3241 2904 ne
rect 3241 2901 3306 2904
rect 3642 2938 3820 2950
rect 3642 2904 3780 2938
rect 3814 2904 3820 2938
rect 3878 2907 3884 2959
rect 3936 2907 3948 2959
rect 4000 2907 4012 2959
rect 4064 2907 4070 2959
rect 4258 2947 4266 2956
rect 4300 2947 4310 2956
rect 4098 2940 4150 2946
rect 3642 2898 3820 2904
rect 3590 2892 3820 2898
rect 2990 2876 3042 2888
tri 3042 2874 3057 2889 sw
tri 4083 2874 4098 2889 se
rect 4098 2876 4150 2888
rect 3042 2865 3057 2874
tri 3057 2865 3066 2874 sw
tri 4074 2865 4083 2874 se
rect 4083 2865 4098 2874
rect 3042 2864 3066 2865
tri 3066 2864 3067 2865 sw
tri 4073 2864 4074 2865 se
rect 4074 2864 4098 2865
rect 3042 2858 4098 2864
rect 3042 2824 3894 2858
rect 3928 2824 3966 2858
rect 4000 2824 4098 2858
rect 2990 2818 4150 2824
rect 4258 2941 4310 2947
rect 4258 2874 4266 2889
rect 4300 2874 4310 2889
rect 4258 2807 4266 2822
rect 4300 2807 4310 2822
rect 2802 2801 2824 2804
tri 2824 2801 2827 2804 nw
rect 2802 2795 2818 2801
tri 2818 2795 2824 2801 nw
rect 2802 2792 2812 2795
rect 2742 2789 2812 2792
tri 2812 2789 2818 2795 nw
rect 2742 2787 2810 2789
tri 2810 2787 2812 2789 nw
tri 1501 2763 1504 2766 se
rect 1504 2763 1533 2766
rect 687 2725 733 2763
tri 733 2738 758 2763 nw
tri 1021 2738 1046 2763 ne
rect 1046 2749 1106 2763
tri 1106 2749 1120 2763 nw
tri 1493 2755 1501 2763 se
rect 1501 2755 1533 2763
tri 1533 2755 1544 2766 nw
tri 1487 2749 1493 2755 se
rect 1493 2749 1527 2755
tri 1527 2749 1533 2755 nw
rect 1046 2737 1094 2749
tri 1094 2737 1106 2749 nw
rect 1380 2737 1510 2749
tri 473 2691 491 2709 sw
rect 687 2691 693 2725
rect 727 2691 733 2725
rect 329 2682 491 2691
tri 491 2682 500 2691 sw
rect 329 2630 445 2682
rect 497 2630 509 2682
rect 561 2630 573 2682
rect 625 2630 631 2682
tri 313 2576 329 2592 se
rect 329 2576 473 2630
tri 473 2603 500 2630 nw
tri 686 2593 687 2594 se
rect 687 2593 733 2691
tri 669 2576 686 2593 se
rect 686 2576 733 2593
tri 306 2569 313 2576 se
rect 313 2569 473 2576
tri 662 2569 669 2576 se
rect 669 2569 733 2576
tri 304 2567 306 2569 se
rect 306 2567 473 2569
rect 0 2492 473 2567
rect 501 2563 733 2569
rect 501 2529 513 2563
rect 547 2529 585 2563
rect 619 2529 733 2563
rect 501 2523 733 2529
rect 772 2714 818 2726
rect 772 2680 778 2714
rect 812 2680 818 2714
rect 772 2637 818 2680
rect 772 2603 778 2637
rect 812 2603 818 2637
rect 772 2560 818 2603
rect 772 2526 778 2560
rect 812 2526 818 2560
tri 473 2492 476 2495 sw
rect 0 2489 476 2492
tri 476 2489 479 2492 sw
rect 0 2483 479 2489
tri 479 2483 485 2489 sw
rect 772 2483 818 2526
rect 0 2470 485 2483
tri 485 2470 498 2483 sw
rect 0 2416 631 2470
rect 0 2364 445 2416
rect 497 2364 509 2416
rect 561 2364 573 2416
rect 625 2364 631 2416
rect 772 2449 778 2483
rect 812 2449 818 2483
rect 772 2407 818 2449
rect 772 2373 778 2407
rect 812 2373 818 2407
tri 763 2355 772 2364 se
rect 772 2355 818 2373
tri 752 2344 763 2355 se
rect 763 2344 818 2355
tri 747 2339 752 2344 se
rect 752 2339 818 2344
tri 744 2336 747 2339 se
rect 747 2336 818 2339
rect 0 2331 818 2336
rect 0 2324 778 2331
rect 0 2290 233 2324
rect 267 2297 778 2324
rect 812 2297 818 2331
rect 267 2290 818 2297
rect 958 2720 1010 2726
rect 958 2646 1010 2668
rect 1046 2725 1092 2737
tri 1092 2735 1094 2737 nw
rect 1046 2691 1052 2725
rect 1086 2691 1092 2725
rect 1046 2681 1092 2691
tri 1092 2681 1097 2686 sw
rect 1046 2679 1097 2681
tri 1097 2679 1099 2681 sw
rect 1046 2668 1099 2679
tri 1099 2668 1110 2679 sw
rect 1150 2668 1156 2720
rect 1208 2668 1220 2720
rect 1272 2668 1284 2720
rect 1336 2668 1352 2720
rect 1380 2703 1386 2737
rect 1420 2732 1510 2737
tri 1510 2732 1527 2749 nw
rect 1746 2732 1752 2766
rect 1786 2732 1792 2766
rect 1420 2729 1507 2732
tri 1507 2729 1510 2732 nw
rect 1420 2721 1499 2729
tri 1499 2721 1507 2729 nw
rect 1420 2709 1439 2721
tri 1439 2709 1451 2721 nw
rect 1420 2703 1426 2709
rect 1046 2666 1110 2668
tri 1046 2665 1047 2666 ne
rect 1047 2665 1110 2666
tri 1110 2665 1113 2668 sw
rect 1380 2665 1426 2703
tri 1426 2696 1439 2709 nw
rect 1746 2694 1792 2732
rect 1820 2723 2032 2775
rect 2084 2723 2096 2775
rect 2148 2723 2160 2775
rect 2212 2723 2224 2775
rect 2276 2723 2288 2775
rect 2340 2723 2403 2775
tri 2742 2779 2750 2787 ne
rect 2750 2785 2808 2787
tri 2808 2785 2810 2787 nw
rect 2750 2780 2802 2785
tri 2462 2709 2475 2722 se
rect 2475 2709 2527 2728
tri 2802 2779 2808 2785 nw
rect 2910 2779 3287 2785
rect 2750 2722 2802 2728
rect 2962 2766 3287 2779
tri 3287 2766 3306 2785 sw
rect 2962 2763 3306 2766
tri 3306 2763 3309 2766 sw
rect 2962 2749 3309 2763
rect 2962 2746 2985 2749
tri 2985 2746 2988 2749 nw
tri 3257 2746 3260 2749 ne
rect 3260 2746 3309 2749
tri 3309 2746 3326 2763 sw
rect 2962 2729 2968 2746
tri 2968 2729 2985 2746 nw
tri 3260 2729 3277 2746 ne
rect 3277 2729 3326 2746
tri 3326 2729 3343 2746 sw
rect 4258 2740 4266 2755
rect 4300 2740 4310 2755
tri 2527 2709 2540 2722 sw
rect 2910 2715 2962 2727
tri 2962 2723 2968 2729 nw
tri 3277 2723 3283 2729 ne
rect 3283 2723 3343 2729
tri 3283 2719 3287 2723 ne
rect 3287 2719 3343 2723
tri 2456 2703 2462 2709 se
rect 2462 2703 2540 2709
tri 1792 2694 1801 2703 sw
tri 2447 2694 2456 2703 se
rect 2456 2694 2540 2703
tri 2540 2694 2555 2709 sw
tri 1047 2631 1081 2665 ne
rect 1081 2631 1113 2665
tri 1113 2631 1147 2665 sw
rect 1380 2631 1386 2665
rect 1420 2631 1426 2665
tri 1081 2630 1082 2631 ne
rect 1082 2630 1147 2631
tri 1147 2630 1148 2631 sw
tri 1082 2625 1087 2630 ne
rect 1087 2625 1148 2630
tri 1148 2625 1153 2630 sw
tri 1087 2620 1092 2625 ne
rect 1092 2620 1150 2625
tri 1092 2619 1093 2620 ne
rect 1093 2619 1150 2620
tri 1093 2594 1118 2619 ne
rect 1118 2594 1150 2619
rect 958 2572 1010 2594
tri 1118 2593 1119 2594 ne
rect 1119 2593 1150 2594
tri 1119 2579 1133 2593 ne
rect 1133 2579 1150 2593
rect 1380 2593 1426 2631
rect 958 2498 1010 2520
rect 1043 2570 1095 2576
rect 1380 2559 1386 2593
rect 1420 2559 1426 2593
rect 1380 2547 1426 2559
rect 1471 2687 1523 2693
rect 1746 2660 1752 2694
rect 1786 2678 1801 2694
tri 1801 2678 1817 2694 sw
tri 2431 2678 2447 2694 se
rect 2447 2678 2484 2694
rect 1786 2660 2484 2678
rect 2518 2660 2608 2694
rect 1746 2648 2608 2660
tri 3287 2711 3295 2719 ne
rect 3295 2711 3343 2719
tri 3343 2711 3361 2729 sw
rect 2910 2657 2962 2663
rect 2990 2705 3042 2711
tri 3295 2709 3297 2711 ne
rect 3297 2709 3361 2711
tri 3361 2709 3363 2711 sw
tri 3297 2691 3315 2709 ne
rect 3315 2691 3363 2709
tri 3363 2691 3381 2709 sw
tri 3315 2680 3326 2691 ne
rect 3326 2680 3381 2691
tri 3381 2680 3392 2691 sw
tri 3326 2657 3349 2680 ne
rect 3349 2674 4150 2680
rect 3349 2657 4098 2674
tri 3349 2656 3350 2657 ne
rect 3350 2656 4098 2657
rect 2990 2641 3042 2653
rect 1471 2580 1523 2635
tri 2984 2631 2990 2637 se
tri 2972 2619 2984 2631 se
rect 2984 2619 2990 2631
tri 2964 2611 2972 2619 se
rect 2972 2611 2990 2619
tri 1638 2594 1655 2611 se
rect 1655 2594 2990 2611
tri 1627 2583 1638 2594 se
rect 1638 2589 2990 2594
tri 3350 2634 3372 2656 ne
rect 3372 2634 4098 2656
tri 4073 2631 4076 2634 ne
rect 4076 2631 4098 2634
tri 4076 2619 4088 2631 ne
rect 4088 2622 4098 2631
rect 4088 2619 4150 2622
tri 4088 2609 4098 2619 ne
rect 4098 2610 4150 2619
rect 1638 2583 3042 2589
rect 3070 2600 3122 2606
tri 1615 2571 1627 2583 se
rect 1627 2571 1655 2583
tri 1655 2571 1667 2583 nw
rect 1043 2504 1095 2518
rect 1150 2484 1156 2536
rect 1208 2484 1220 2536
rect 1272 2484 1284 2536
rect 1336 2484 1352 2536
tri 1604 2560 1615 2571 se
rect 1615 2560 1644 2571
tri 1644 2560 1655 2571 nw
tri 3236 2591 3241 2596 se
rect 3241 2591 3306 2596
tri 3230 2585 3236 2591 se
rect 3236 2585 3306 2591
tri 3228 2583 3230 2585 se
rect 3230 2583 3306 2585
tri 3227 2582 3228 2583 se
rect 3228 2582 3306 2583
tri 3220 2575 3227 2582 se
rect 3227 2575 3306 2582
tri 1599 2555 1604 2560 se
rect 1604 2555 1639 2560
tri 1639 2555 1644 2560 nw
tri 1592 2548 1599 2555 se
rect 1599 2548 1632 2555
tri 1632 2548 1639 2555 nw
rect 1792 2549 2527 2555
tri 1591 2547 1592 2548 se
rect 1592 2547 1631 2548
tri 1631 2547 1632 2548 nw
tri 1589 2545 1591 2547 se
rect 1591 2545 1629 2547
tri 1629 2545 1631 2547 nw
tri 1580 2536 1589 2545 se
rect 1589 2536 1620 2545
tri 1620 2536 1629 2545 nw
tri 1575 2531 1580 2536 se
rect 1580 2531 1615 2536
tri 1615 2531 1620 2536 nw
rect 1471 2522 1523 2528
tri 1568 2524 1575 2531 se
rect 1575 2524 1608 2531
tri 1608 2524 1615 2531 nw
rect 1663 2524 1709 2536
tri 1566 2522 1568 2524 se
rect 1568 2522 1575 2524
tri 1535 2491 1566 2522 se
rect 1566 2491 1575 2522
tri 1575 2491 1608 2524 nw
tri 1534 2490 1535 2491 se
rect 1535 2490 1574 2491
tri 1574 2490 1575 2491 nw
rect 1663 2490 1669 2524
rect 1703 2490 1709 2524
tri 1529 2485 1534 2490 se
rect 1534 2485 1569 2490
tri 1569 2485 1574 2490 nw
tri 1528 2484 1529 2485 se
rect 1529 2484 1560 2485
tri 1520 2476 1528 2484 se
rect 1528 2476 1560 2484
tri 1560 2476 1569 2485 nw
tri 1519 2475 1520 2476 se
rect 1520 2475 1559 2476
tri 1559 2475 1560 2476 nw
tri 1517 2473 1519 2475 se
rect 1519 2473 1557 2475
tri 1557 2473 1559 2475 nw
rect 1043 2446 1095 2452
rect 1380 2461 1535 2473
rect 958 2424 1010 2446
tri 1119 2427 1133 2441 se
rect 1133 2427 1150 2441
tri 1109 2417 1119 2427 se
rect 1119 2417 1150 2427
tri 1108 2416 1109 2417 se
rect 1109 2416 1150 2417
tri 1102 2410 1108 2416 se
rect 1108 2410 1150 2416
tri 1095 2403 1102 2410 se
rect 1102 2403 1150 2410
tri 1085 2393 1095 2403 se
rect 1095 2395 1150 2403
rect 1380 2427 1386 2461
rect 1420 2451 1535 2461
tri 1535 2451 1557 2473 nw
rect 1663 2451 1709 2490
rect 1420 2445 1529 2451
tri 1529 2445 1535 2451 nw
rect 1420 2427 1426 2445
rect 1095 2393 1151 2395
tri 1151 2393 1153 2395 nw
tri 1081 2389 1085 2393 se
rect 1085 2389 1147 2393
tri 1147 2389 1151 2393 nw
rect 1380 2389 1426 2427
tri 1426 2420 1451 2445 nw
rect 1663 2417 1669 2451
rect 1703 2417 1709 2451
tri 1067 2375 1081 2389 se
rect 1081 2375 1133 2389
tri 1133 2375 1147 2389 nw
rect 958 2351 1010 2372
tri 1056 2364 1067 2375 se
rect 1067 2364 1113 2375
tri 1047 2355 1056 2364 se
rect 1056 2355 1113 2364
tri 1113 2355 1133 2375 nw
rect 1380 2355 1386 2389
rect 1420 2355 1426 2389
rect 958 2293 1010 2299
tri 1046 2354 1047 2355 se
rect 1047 2354 1112 2355
tri 1112 2354 1113 2355 nw
rect 1046 2352 1110 2354
tri 1110 2352 1112 2354 nw
rect 1046 2344 1102 2352
tri 1102 2344 1110 2352 nw
rect 1046 2335 1093 2344
tri 1093 2335 1102 2344 nw
rect 0 2285 818 2290
rect 0 2282 295 2285
tri 295 2282 298 2285 nw
rect 1046 2282 1092 2335
tri 1092 2334 1093 2335 nw
rect 1150 2300 1156 2352
rect 1208 2300 1220 2352
rect 1272 2300 1284 2352
rect 1336 2300 1352 2352
rect 1380 2343 1426 2355
rect 1471 2399 1523 2405
rect 1471 2334 1523 2347
tri 1092 2282 1095 2285 sw
rect 0 2271 284 2282
tri 284 2271 295 2282 nw
tri 1035 2271 1046 2282 se
rect 1046 2271 1095 2282
tri 1095 2271 1106 2282 sw
rect 0 2234 273 2271
tri 273 2260 284 2271 nw
tri 1024 2260 1035 2271 se
rect 1035 2260 1106 2271
tri 1106 2260 1117 2271 sw
rect 1471 2269 1523 2282
tri 1023 2259 1024 2260 se
rect 1024 2259 1117 2260
tri 1117 2259 1118 2260 sw
tri 1021 2257 1023 2259 se
rect 1023 2257 1118 2259
tri 1118 2257 1120 2259 sw
rect 0 2200 233 2234
rect 267 2200 273 2234
rect 631 2235 1150 2257
rect 631 2211 1043 2235
rect 0 2145 273 2200
tri 1018 2198 1031 2211 ne
rect 1031 2198 1043 2211
tri 1031 2186 1043 2198 ne
rect 1095 2211 1150 2235
rect 1471 2211 1480 2217
rect 1514 2211 1523 2217
rect 1095 2198 1107 2211
tri 1107 2198 1120 2211 nw
rect 1471 2204 1523 2211
tri 1095 2186 1107 2198 nw
rect 0 2111 233 2145
rect 267 2140 273 2145
tri 273 2140 298 2165 sw
tri 747 2140 772 2165 se
rect 772 2140 818 2183
rect 267 2134 818 2140
rect 267 2111 333 2134
rect 0 2100 333 2111
rect 367 2100 414 2134
rect 448 2100 495 2134
rect 529 2100 576 2134
rect 610 2100 658 2134
rect 692 2100 740 2134
rect 774 2100 818 2134
rect 0 2094 818 2100
rect 849 2177 901 2183
rect 1043 2169 1095 2183
tri 901 2137 919 2155 sw
rect 901 2125 919 2137
tri 919 2125 931 2137 sw
rect 849 2113 931 2125
rect 901 2111 931 2113
tri 931 2111 945 2125 sw
rect 1043 2111 1095 2117
rect 1150 2116 1156 2168
rect 1208 2116 1220 2168
rect 1272 2116 1284 2168
rect 1336 2116 1352 2168
rect 1471 2139 1480 2152
rect 1514 2139 1523 2152
rect 901 2110 945 2111
tri 945 2110 946 2111 sw
rect 901 2102 946 2110
tri 946 2102 954 2110 sw
rect 901 2099 954 2102
tri 954 2099 957 2102 sw
rect 901 2097 957 2099
tri 957 2097 959 2099 sw
rect 901 2072 959 2097
tri 959 2072 984 2097 sw
rect 1471 2074 1480 2087
rect 1514 2074 1523 2087
rect 901 2063 984 2072
tri 984 2063 993 2072 sw
rect 901 2061 993 2063
rect 849 2055 993 2061
tri 993 2055 1001 2063 sw
tri 947 2052 950 2055 ne
rect 950 2052 1001 2055
tri 1001 2052 1004 2055 sw
tri 950 2038 964 2052 ne
rect 964 2038 1004 2052
tri 1004 2038 1018 2052 sw
tri 232 2028 240 2036 se
rect 240 2030 292 2036
tri 228 2024 232 2028 se
rect 232 2024 240 2028
tri 227 2023 228 2024 se
rect 228 2023 240 2024
tri 224 2020 227 2023 se
rect 227 2020 240 2023
rect 0 1978 240 2020
rect 329 1986 335 2038
rect 387 1986 399 2038
rect 451 1986 463 2038
rect 515 2028 521 2038
tri 521 2028 531 2038 sw
tri 964 2028 974 2038 ne
rect 974 2028 1018 2038
tri 1018 2028 1028 2038 sw
rect 515 2027 531 2028
tri 531 2027 532 2028 sw
tri 974 2027 975 2028 ne
rect 975 2027 1028 2028
tri 1028 2027 1029 2028 sw
rect 515 2021 901 2027
tri 975 2024 978 2027 ne
rect 978 2024 1029 2027
tri 1029 2024 1032 2027 sw
tri 978 2023 979 2024 ne
rect 979 2023 1032 2024
tri 1032 2023 1033 2024 sw
rect 515 1986 849 2021
tri 824 1979 831 1986 ne
rect 831 1979 849 1986
rect 0 1966 292 1978
rect 0 1953 240 1966
tri 195 1950 198 1953 ne
rect 198 1950 240 1953
tri 198 1949 199 1950 ne
rect 199 1949 240 1950
tri 199 1946 202 1949 ne
rect 202 1946 240 1949
tri 202 1912 236 1946 ne
rect 236 1914 240 1946
tri 831 1961 849 1979 ne
tri 979 2018 984 2023 ne
rect 984 2018 1033 2023
tri 1033 2018 1038 2023 sw
tri 984 1989 1013 2018 ne
rect 1013 1989 1038 2018
tri 1038 1989 1067 2018 sw
rect 1471 2009 1480 2022
rect 1514 2009 1523 2022
tri 1013 1979 1023 1989 ne
rect 1023 1979 1067 1989
tri 1067 1979 1077 1989 sw
rect 849 1957 901 1969
tri 1023 1964 1038 1979 ne
rect 1038 1964 1077 1979
tri 1077 1964 1092 1979 sw
rect 236 1912 292 1914
tri 236 1908 240 1912 ne
rect 240 1908 292 1912
rect 333 1946 818 1952
rect 333 1912 345 1946
rect 379 1912 423 1946
rect 457 1912 501 1946
rect 535 1912 579 1946
rect 613 1912 657 1946
rect 691 1912 818 1946
rect 333 1908 818 1912
rect 333 1906 778 1908
tri 747 1881 772 1906 ne
rect 2 1874 317 1880
tri 317 1874 323 1880 sw
rect 772 1874 778 1906
rect 812 1886 818 1908
tri 1038 1956 1046 1964 ne
rect 849 1899 901 1905
rect 958 1944 1010 1950
tri 818 1886 820 1888 sw
tri 956 1886 958 1888 se
rect 958 1886 1010 1892
rect 812 1875 820 1886
tri 820 1875 831 1886 sw
tri 945 1875 956 1886 se
rect 956 1879 1010 1886
rect 956 1875 958 1879
rect 812 1874 831 1875
rect 2 1859 323 1874
tri 323 1859 338 1874 sw
rect 772 1863 831 1874
tri 831 1863 843 1875 sw
tri 933 1863 945 1875 se
rect 945 1863 958 1875
rect 2 1834 338 1859
tri 338 1834 363 1859 sw
rect 2 1825 228 1834
tri 228 1825 237 1834 nw
tri 292 1825 301 1834 ne
rect 301 1825 363 1834
tri 363 1825 372 1834 sw
rect 2 1810 213 1825
tri 213 1810 228 1825 nw
tri 301 1810 316 1825 ne
rect 316 1816 372 1825
tri 372 1816 381 1825 sw
rect 316 1810 389 1816
rect 2 1809 212 1810
tri 212 1809 213 1810 nw
tri 316 1809 317 1810 ne
rect 317 1809 389 1810
rect 2 1804 74 1809
tri 74 1804 79 1809 nw
tri 317 1804 322 1809 ne
rect 322 1804 389 1809
rect 2 1784 54 1804
tri 54 1784 74 1804 nw
tri 322 1784 342 1804 ne
rect 342 1784 349 1804
tri 342 1783 343 1784 ne
rect 343 1770 349 1784
rect 383 1770 389 1804
rect 619 1788 733 1834
tri 649 1780 657 1788 ne
rect 657 1780 733 1788
rect 241 1736 293 1742
rect 343 1732 389 1770
tri 657 1750 687 1780 ne
rect 343 1698 349 1732
rect 383 1698 389 1732
rect 343 1686 389 1698
rect 241 1663 293 1684
rect 241 1591 293 1611
rect 241 1519 293 1539
rect 241 1447 293 1467
rect 241 1375 293 1395
rect 241 1303 293 1323
rect 329 1612 417 1658
rect 329 1588 389 1612
tri 389 1588 413 1612 nw
rect 329 1579 380 1588
tri 380 1579 389 1588 nw
rect 329 1339 375 1579
tri 375 1574 380 1579 nw
tri 677 1510 687 1520 se
rect 687 1510 733 1780
rect 772 1827 958 1863
rect 772 1825 967 1827
rect 1001 1825 1010 1827
rect 772 1791 778 1825
rect 812 1814 1010 1825
rect 812 1791 958 1814
rect 772 1762 958 1791
rect 772 1749 967 1762
rect 1001 1749 1010 1762
rect 772 1743 958 1749
rect 772 1709 778 1743
rect 812 1709 958 1743
rect 772 1697 958 1709
rect 772 1684 967 1697
rect 1001 1684 1010 1697
rect 772 1661 958 1684
rect 772 1627 778 1661
rect 812 1632 958 1661
rect 812 1627 1010 1632
rect 772 1622 1010 1627
rect 772 1620 967 1622
rect 1001 1620 1010 1622
rect 772 1606 958 1620
rect 772 1588 825 1606
tri 825 1588 843 1606 nw
tri 933 1588 951 1606 ne
rect 951 1588 958 1606
rect 1046 1851 1092 1964
rect 1471 1949 1523 1957
rect 1471 1944 1480 1949
rect 1514 1944 1523 1949
rect 1150 1865 1156 1917
rect 1208 1865 1220 1917
rect 1272 1865 1284 1917
rect 1336 1865 1352 1917
rect 1471 1879 1523 1892
rect 1046 1817 1052 1851
rect 1086 1817 1092 1851
rect 1046 1779 1092 1817
rect 1150 1828 1426 1834
rect 1150 1794 1162 1828
rect 1196 1794 1234 1828
rect 1268 1794 1306 1828
rect 1340 1794 1426 1828
rect 1150 1788 1426 1794
rect 1046 1745 1052 1779
rect 1086 1745 1092 1779
tri 1352 1767 1373 1788 ne
rect 1373 1767 1426 1788
tri 1373 1760 1380 1767 ne
rect 1046 1707 1092 1745
rect 1046 1673 1052 1707
rect 1086 1673 1092 1707
rect 1150 1696 1156 1748
rect 1208 1696 1220 1748
rect 1272 1696 1284 1748
rect 1336 1696 1352 1748
tri 1377 1681 1380 1684 se
rect 1380 1681 1426 1767
rect 1046 1635 1092 1673
tri 1352 1656 1377 1681 se
rect 1377 1656 1426 1681
rect 1046 1601 1052 1635
rect 1086 1601 1092 1635
rect 1150 1650 1426 1656
rect 1150 1616 1162 1650
rect 1196 1616 1234 1650
rect 1268 1616 1306 1650
rect 1340 1616 1426 1650
rect 1150 1610 1426 1616
rect 1046 1589 1092 1601
tri 1352 1600 1362 1610 ne
rect 1362 1600 1426 1610
tri 1362 1590 1372 1600 ne
rect 1372 1590 1426 1600
tri 1372 1589 1373 1590 ne
rect 1373 1589 1426 1590
rect 772 1579 818 1588
tri 818 1581 825 1588 nw
tri 951 1581 958 1588 ne
rect 772 1545 778 1579
rect 812 1545 818 1579
rect 772 1533 818 1545
rect 849 1564 901 1570
tri 676 1509 677 1510 se
rect 677 1509 733 1510
tri 672 1505 676 1509 se
rect 676 1505 733 1509
tri 733 1505 737 1509 sw
tri 649 1482 672 1505 se
rect 672 1482 737 1505
rect 619 1471 737 1482
tri 737 1471 771 1505 sw
rect 849 1500 901 1512
rect 619 1470 771 1471
tri 771 1470 772 1471 sw
rect 619 1468 772 1470
tri 772 1468 774 1470 sw
rect 619 1442 774 1468
tri 774 1442 800 1468 sw
tri 1373 1582 1380 1589 ne
rect 958 1556 1010 1568
rect 1150 1518 1156 1570
rect 1208 1518 1220 1570
rect 1272 1518 1284 1570
rect 1336 1518 1352 1570
rect 958 1498 1010 1504
tri 901 1471 925 1495 sw
rect 901 1470 925 1471
tri 925 1470 926 1471 sw
rect 901 1448 1092 1470
rect 849 1442 1092 1448
tri 1358 1442 1380 1464 se
rect 1380 1442 1426 1589
rect 619 1440 800 1442
tri 800 1440 802 1442 sw
tri 1021 1440 1023 1442 ne
rect 1023 1440 1092 1442
tri 1356 1440 1358 1442 se
rect 1358 1440 1426 1442
rect 619 1439 802 1440
tri 802 1439 803 1440 sw
tri 1023 1439 1024 1440 ne
rect 1024 1439 1092 1440
tri 1355 1439 1356 1440 se
rect 1356 1439 1426 1440
rect 619 1436 803 1439
tri 750 1431 755 1436 ne
rect 755 1431 803 1436
tri 803 1431 811 1439 sw
tri 1024 1431 1032 1439 ne
rect 1032 1431 1092 1439
tri 755 1414 772 1431 ne
rect 772 1414 811 1431
tri 811 1414 828 1431 sw
tri 1032 1417 1046 1431 ne
tri 772 1400 786 1414 ne
rect 786 1400 901 1414
tri 786 1388 798 1400 ne
rect 798 1388 901 1400
rect 687 1382 739 1388
tri 798 1385 801 1388 ne
rect 801 1385 901 1388
tri 375 1339 380 1344 sw
rect 329 1323 380 1339
tri 380 1323 396 1339 sw
tri 679 1323 687 1331 se
tri 801 1366 820 1385 ne
rect 820 1366 901 1385
tri 820 1340 846 1366 ne
rect 687 1323 739 1330
rect 329 1322 396 1323
tri 396 1322 397 1323 sw
tri 678 1322 679 1323 se
rect 679 1322 739 1323
rect 329 1321 397 1322
tri 397 1321 398 1322 sw
tri 677 1321 678 1322 se
rect 678 1321 739 1322
rect 329 1315 398 1321
tri 398 1315 404 1321 sw
tri 671 1315 677 1321 se
rect 677 1318 739 1321
rect 677 1315 687 1318
rect 329 1306 404 1315
tri 404 1306 413 1315 sw
tri 662 1306 671 1315 se
rect 671 1306 687 1315
rect 329 1260 417 1306
rect 619 1266 687 1306
rect 619 1260 739 1266
rect 772 1315 818 1327
rect 772 1281 778 1315
rect 812 1281 818 1315
rect 241 1231 293 1251
rect 772 1250 818 1281
rect 846 1287 901 1366
rect 958 1406 1010 1412
rect 958 1333 1010 1354
tri 901 1287 903 1289 sw
rect 846 1274 903 1287
tri 846 1270 850 1274 ne
rect 850 1270 903 1274
tri 903 1270 920 1287 sw
rect 958 1275 1010 1281
rect 1046 1373 1092 1431
tri 1352 1436 1355 1439 se
rect 1355 1436 1426 1439
rect 1352 1390 1426 1436
tri 1352 1385 1357 1390 ne
rect 1357 1385 1426 1390
rect 1046 1339 1052 1373
rect 1086 1339 1092 1373
tri 1357 1366 1376 1385 ne
rect 1376 1366 1426 1385
tri 1376 1364 1378 1366 ne
rect 1378 1364 1426 1366
tri 1378 1362 1380 1364 ne
rect 1046 1301 1092 1339
tri 850 1267 853 1270 ne
rect 853 1267 920 1270
tri 920 1267 923 1270 sw
rect 1046 1267 1052 1301
rect 1086 1267 1092 1301
tri 853 1260 860 1267 ne
rect 860 1260 923 1267
tri 923 1260 930 1267 sw
tri 860 1258 862 1260 ne
rect 862 1258 930 1260
tri 818 1250 826 1258 sw
tri 862 1250 870 1258 ne
rect 870 1255 930 1258
tri 930 1255 935 1260 sw
rect 1046 1255 1092 1267
rect 870 1250 935 1255
tri 935 1250 940 1255 sw
rect 772 1249 826 1250
tri 826 1249 827 1250 sw
tri 870 1249 871 1250 ne
rect 871 1249 940 1250
tri 940 1249 941 1250 sw
rect 772 1230 827 1249
tri 827 1230 846 1249 sw
tri 871 1230 890 1249 ne
rect 890 1230 941 1249
tri 941 1230 960 1249 sw
rect 772 1225 846 1230
tri 846 1225 851 1230 sw
tri 890 1225 895 1230 ne
rect 895 1225 960 1230
tri 960 1225 965 1230 sw
rect 772 1219 851 1225
tri 851 1219 857 1225 sw
tri 895 1219 901 1225 ne
rect 901 1219 965 1225
rect 772 1211 857 1219
tri 857 1211 865 1219 sw
tri 901 1211 909 1219 ne
rect 909 1211 965 1219
tri 965 1211 979 1225 sw
rect 772 1200 865 1211
tri 865 1200 876 1211 sw
tri 909 1200 920 1211 ne
rect 920 1200 979 1211
tri 979 1200 990 1211 sw
rect 772 1199 876 1200
tri 876 1199 877 1200 sw
tri 920 1199 921 1200 ne
rect 921 1199 1227 1200
rect 241 1173 293 1179
rect 417 1147 445 1199
rect 497 1147 509 1199
rect 561 1147 573 1199
rect 625 1147 631 1199
rect 772 1177 877 1199
tri 877 1177 899 1199 sw
tri 921 1177 943 1199 ne
rect 943 1177 1227 1199
rect 772 1176 899 1177
tri 899 1176 900 1177 sw
tri 943 1176 944 1177 ne
rect 944 1176 1227 1177
rect 0 1133 389 1145
rect 0 1099 349 1133
rect 383 1099 389 1133
rect 772 1142 778 1176
rect 812 1170 900 1176
tri 900 1170 906 1176 sw
tri 944 1170 950 1176 ne
rect 950 1170 1227 1176
rect 812 1162 906 1170
tri 906 1162 914 1170 sw
tri 950 1162 958 1170 ne
rect 958 1162 1227 1170
rect 812 1154 914 1162
tri 914 1154 922 1162 sw
tri 958 1154 966 1162 ne
rect 966 1154 1227 1162
rect 812 1151 922 1154
tri 922 1151 925 1154 sw
tri 966 1151 969 1154 ne
rect 969 1151 1190 1154
rect 812 1147 925 1151
tri 925 1147 929 1151 sw
tri 1098 1147 1102 1151 ne
rect 1102 1147 1190 1151
tri 1190 1147 1197 1154 nw
rect 812 1145 929 1147
tri 929 1145 931 1147 sw
tri 1102 1145 1104 1147 ne
rect 1104 1145 1188 1147
tri 1188 1145 1190 1147 nw
rect 812 1142 931 1145
rect 772 1138 931 1142
tri 931 1138 938 1145 sw
tri 1104 1138 1111 1145 ne
rect 1111 1138 1181 1145
tri 1181 1138 1188 1145 nw
rect 772 1130 938 1138
tri 938 1130 946 1138 sw
tri 1111 1130 1119 1138 ne
rect 1119 1130 1169 1138
tri 834 1118 846 1130 ne
rect 846 1126 946 1130
tri 946 1126 950 1130 sw
tri 1119 1126 1123 1130 ne
rect 846 1118 950 1126
tri 950 1118 958 1126 sw
tri 846 1106 858 1118 ne
rect 858 1112 1010 1118
rect 858 1106 958 1112
tri 858 1102 862 1106 ne
rect 862 1102 958 1106
tri 318 1074 343 1099 ne
rect 343 1061 389 1099
rect 343 1027 349 1061
rect 383 1027 389 1061
rect 769 1096 821 1102
tri 755 1031 769 1045 se
tri 862 1072 892 1102 ne
rect 892 1072 958 1102
tri 892 1065 899 1072 ne
rect 899 1065 958 1072
rect 769 1032 821 1044
tri 754 1030 755 1031 se
rect 755 1030 769 1031
rect 343 1015 389 1027
tri 744 1020 754 1030 se
rect 754 1020 769 1030
rect 619 980 769 1020
tri 899 1031 933 1065 ne
rect 933 1060 958 1065
rect 933 1042 1010 1060
rect 933 1031 958 1042
tri 933 1030 934 1031 ne
rect 934 1030 958 1031
tri 934 1006 958 1030 ne
rect 958 984 1010 990
rect 1043 1042 1095 1048
rect 619 974 821 980
rect 1043 976 1095 990
rect 0 958 198 972
tri 198 958 212 972 sw
tri 1030 958 1043 971 se
rect 0 946 212 958
tri 212 946 224 958 sw
tri 1018 946 1030 958 se
rect 1030 946 1043 958
rect 0 944 1043 946
tri 186 924 206 944 ne
rect 206 924 1043 944
tri 206 919 211 924 ne
rect 211 919 1095 924
tri 211 918 212 919 ne
rect 212 918 1095 919
rect 241 878 293 890
rect 241 867 250 878
rect 284 867 293 878
rect 241 801 293 815
rect 241 735 293 749
rect 241 669 293 683
rect 241 610 250 617
rect 284 610 293 617
rect 241 602 293 610
rect 241 535 250 550
rect 284 535 293 550
rect 343 871 389 883
rect 343 837 349 871
rect 383 837 389 871
rect 777 876 1010 882
rect 343 799 389 837
rect 343 765 349 799
rect 383 765 389 799
rect 417 795 445 847
rect 497 795 509 847
rect 561 795 573 847
rect 625 795 631 847
rect 777 842 789 876
rect 823 842 861 876
rect 895 842 958 876
rect 777 836 958 842
tri 875 812 899 836 ne
rect 899 824 958 836
rect 899 812 1010 824
tri 899 811 900 812 ne
rect 900 811 1010 812
tri 900 802 909 811 ne
rect 909 808 1010 811
rect 909 802 958 808
tri 909 796 915 802 ne
rect 915 796 958 802
tri 915 795 916 796 ne
rect 916 795 958 796
tri 916 773 938 795 ne
rect 938 773 958 795
rect 343 727 389 765
tri 938 753 958 773 ne
rect 343 693 349 727
rect 383 693 389 727
rect 769 744 821 750
rect 343 655 389 693
tri 744 668 769 693 se
rect 769 680 821 692
rect 343 621 349 655
rect 383 621 389 655
rect 619 628 769 668
rect 619 622 821 628
rect 849 744 901 750
rect 958 740 1010 756
tri 901 694 903 696 sw
rect 901 692 903 694
rect 849 682 903 692
tri 903 682 915 694 sw
rect 958 682 1010 688
rect 1123 750 1169 1130
tri 1169 1126 1181 1138 nw
tri 1352 964 1380 992 se
rect 1380 964 1426 1364
rect 1197 958 1426 964
rect 1197 924 1209 958
rect 1243 924 1319 958
rect 1353 924 1426 958
rect 1197 918 1426 924
tri 1352 890 1380 918 ne
tri 1169 750 1175 756 sw
rect 1123 739 1175 750
tri 1175 739 1186 750 sw
rect 1123 738 1186 739
tri 1186 738 1187 739 sw
rect 1123 729 1187 738
tri 1187 729 1196 738 sw
rect 1123 728 1196 729
tri 1196 728 1197 729 sw
rect 1123 682 1227 728
rect 849 680 915 682
rect 901 666 915 680
tri 915 666 931 682 sw
rect 901 665 931 666
tri 931 665 932 666 sw
rect 901 661 932 665
tri 932 661 936 665 sw
rect 901 658 936 661
tri 936 658 939 661 sw
rect 901 656 939 658
tri 939 656 941 658 sw
rect 901 654 941 656
tri 941 654 943 656 sw
rect 901 642 1092 654
rect 901 628 1052 642
rect 343 583 389 621
rect 849 608 1052 628
rect 1086 608 1092 642
rect 343 549 349 583
rect 383 549 389 583
rect 343 537 389 549
rect 772 582 818 594
rect 772 548 778 582
rect 812 548 818 582
rect 849 571 1092 608
tri 849 570 850 571 ne
rect 850 570 1092 571
rect 772 520 818 548
tri 850 536 884 570 ne
rect 884 536 1052 570
rect 1086 536 1092 570
tri 884 524 896 536 ne
rect 896 524 1092 536
tri 818 520 819 521 sw
rect 772 519 819 520
tri 819 519 820 520 sw
tri 1379 519 1380 520 se
rect 1380 519 1426 918
rect 772 517 820 519
tri 820 517 822 519 sw
tri 1377 517 1379 519 se
rect 1379 517 1426 519
rect 772 506 822 517
tri 822 506 833 517 sw
tri 1366 506 1377 517 se
rect 1377 506 1426 517
rect 772 499 833 506
rect 241 468 250 483
rect 284 468 293 483
rect 417 443 433 495
rect 485 443 497 495
rect 549 443 561 495
rect 613 443 619 495
rect 772 465 778 499
rect 812 496 833 499
tri 833 496 843 506 sw
tri 1356 496 1366 506 se
rect 1366 496 1426 506
rect 812 484 1007 496
rect 812 465 967 484
rect 772 450 967 465
rect 1001 450 1007 484
rect 241 407 293 416
rect 241 401 250 407
rect 284 401 293 407
rect 772 407 1007 450
tri 1352 492 1356 496 se
rect 1356 492 1426 496
rect 1352 446 1426 492
rect 1471 1814 1523 1827
rect 1471 1749 1523 1762
rect 1471 1693 1480 1697
rect 1514 1693 1523 1697
rect 1471 1684 1523 1693
rect 1471 1620 1480 1632
rect 1514 1620 1523 1632
rect 1471 1556 1480 1568
rect 1514 1556 1523 1568
rect 1471 1492 1480 1504
rect 1514 1492 1523 1504
rect 1471 1431 1523 1440
rect 1471 1428 1480 1431
rect 1514 1428 1523 1431
rect 1471 1364 1523 1376
rect 1471 1300 1523 1312
rect 1471 1236 1523 1248
rect 1471 1177 1480 1184
rect 1514 1177 1523 1184
rect 1471 1172 1523 1177
rect 1471 1108 1480 1120
rect 1514 1108 1523 1120
rect 1471 1044 1480 1056
rect 1514 1044 1523 1056
rect 1471 980 1480 992
rect 1514 980 1523 992
rect 1471 919 1523 928
rect 1471 916 1480 919
rect 1514 916 1523 919
rect 1471 852 1523 864
rect 1471 788 1523 800
rect 1471 724 1523 736
rect 1471 666 1480 672
rect 1514 666 1523 672
rect 1471 660 1523 666
rect 1471 596 1480 608
rect 1514 596 1523 608
rect 1471 532 1480 544
rect 1514 532 1523 544
rect 1471 468 1480 480
rect 1514 468 1523 480
tri 293 375 318 400 sw
tri 747 375 772 400 se
rect 772 375 967 407
rect 293 373 967 375
rect 1001 375 1007 407
rect 1471 404 1523 416
tri 1007 375 1032 400 sw
tri 1446 375 1471 400 se
rect 1001 373 1471 375
rect 293 369 1471 373
rect 293 349 365 369
rect 241 335 365 349
rect 399 335 440 369
rect 474 335 515 369
rect 549 335 590 369
rect 624 335 665 369
rect 699 335 740 369
rect 774 335 1077 369
rect 1111 335 1150 369
rect 1184 335 1223 369
rect 1257 335 1296 369
rect 1330 335 1369 369
rect 1403 335 1442 369
rect 1476 335 1523 352
rect 241 329 1523 335
rect 1663 2378 1709 2417
rect 1663 2344 1669 2378
rect 1703 2344 1709 2378
rect 1663 2305 1709 2344
rect 1792 2497 2475 2549
rect 1792 2485 2527 2497
rect 1792 2433 2475 2485
rect 1792 2421 2527 2433
rect 2910 2545 3040 2551
rect 2962 2511 2994 2545
rect 3028 2511 3040 2545
rect 2962 2505 3040 2511
rect 3070 2526 3122 2548
rect 3878 2539 3884 2591
rect 3936 2539 3948 2591
rect 4000 2539 4012 2591
rect 4064 2539 4070 2591
rect 4098 2552 4150 2558
rect 4258 2673 4266 2688
rect 4300 2673 4310 2688
rect 4258 2619 4310 2621
rect 4258 2606 4266 2619
rect 4300 2606 4310 2619
rect 4258 2547 4310 2554
rect 4258 2539 4266 2547
rect 4300 2539 4310 2547
rect 2962 2498 2980 2505
tri 2980 2498 2987 2505 nw
rect 2962 2493 2967 2498
rect 2910 2485 2967 2493
tri 2967 2485 2980 2498 nw
rect 2910 2484 2966 2485
tri 2966 2484 2967 2485 nw
rect 2910 2481 2962 2484
tri 2962 2480 2966 2484 nw
rect 2910 2423 2962 2429
tri 4164 2484 4178 2498 se
rect 4178 2492 4230 2498
rect 3070 2452 3122 2474
rect 1792 2369 2475 2421
tri 2817 2410 2830 2423 se
rect 2830 2417 2882 2423
tri 2810 2403 2817 2410 se
rect 2817 2403 2830 2410
rect 1792 2364 2527 2369
rect 1792 2363 1816 2364
tri 1816 2363 1817 2364 nw
tri 2453 2363 2454 2364 ne
rect 2454 2363 2527 2364
tri 1792 2339 1816 2363 nw
tri 2454 2339 2478 2363 ne
rect 1663 2271 1669 2305
rect 1703 2271 1709 2305
rect 1663 2232 1709 2271
rect 1820 2267 2032 2319
rect 2084 2267 2096 2319
rect 2148 2267 2160 2319
rect 2212 2267 2224 2319
rect 2276 2267 2288 2319
rect 2340 2267 2403 2319
rect 1663 2198 1669 2232
rect 1703 2198 1709 2232
rect 1663 2159 1709 2198
rect 1663 2125 1669 2159
rect 1703 2125 1709 2159
rect 1663 2086 1709 2125
rect 1663 2052 1669 2086
rect 1703 2052 1709 2086
rect 1663 2013 1709 2052
rect 1663 1979 1669 2013
rect 1703 1979 1709 2013
rect 1663 1940 1709 1979
rect 1663 1906 1669 1940
rect 1703 1906 1709 1940
rect 1663 1867 1709 1906
tri 1792 2226 1813 2247 sw
tri 2457 2226 2478 2247 se
rect 2478 2226 2527 2363
tri 2789 2382 2810 2403 se
rect 2810 2382 2830 2403
rect 2789 2365 2830 2382
rect 2789 2353 2882 2365
rect 2789 2336 2830 2353
tri 2789 2335 2790 2336 ne
rect 2790 2335 2830 2336
tri 2790 2331 2794 2335 ne
rect 2794 2331 2830 2335
tri 2794 2297 2828 2331 ne
rect 2828 2301 2830 2331
rect 2828 2297 2882 2301
tri 2828 2295 2830 2297 ne
rect 2830 2295 2882 2297
rect 4084 2440 4178 2484
rect 4084 2438 4230 2440
tri 4144 2428 4154 2438 ne
rect 4154 2428 4230 2438
tri 4154 2423 4159 2428 ne
rect 4159 2423 4178 2428
tri 4159 2411 4171 2423 ne
rect 4171 2411 4178 2423
tri 4171 2404 4178 2411 ne
rect 3070 2378 3122 2400
rect 3878 2343 3884 2395
rect 3936 2343 3948 2395
rect 4000 2343 4012 2395
rect 4064 2343 4084 2395
rect 4178 2370 4230 2376
rect 4258 2475 4310 2487
rect 4258 2472 4266 2475
rect 4300 2472 4310 2475
rect 4258 2405 4310 2420
rect 4637 3076 4689 3082
rect 4637 3010 4689 3024
rect 4637 2943 4689 2958
rect 4637 2884 4646 2891
rect 4680 2884 4689 2891
rect 4637 2876 4689 2884
rect 4637 2809 4646 2824
rect 4680 2809 4689 2824
rect 4637 2742 4646 2757
rect 4680 2742 4689 2757
rect 4637 2675 4646 2690
rect 4680 2675 4689 2690
rect 4637 2614 4689 2623
rect 4637 2608 4646 2614
rect 4680 2608 4689 2614
rect 4637 2541 4689 2556
rect 4637 2474 4689 2489
rect 4829 3065 4835 3099
tri 6954 3098 6956 3100 se
rect 6956 3098 7040 3100
tri 6952 3096 6954 3098 se
rect 6954 3096 7040 3098
rect 4869 3079 4892 3092
rect 4829 3027 4840 3065
tri 6920 3064 6952 3096 se
rect 6952 3064 6970 3096
rect 4829 3021 4892 3027
rect 4829 2987 4835 3021
rect 4869 3014 4892 3021
rect 4946 3062 6970 3064
rect 7004 3062 7040 3096
rect 9617 3096 9620 3148
rect 9617 3084 9672 3096
rect 4946 3058 7040 3062
rect 4946 3024 4958 3058
rect 4992 3024 5030 3058
rect 5064 3050 7040 3058
rect 5064 3048 7092 3050
rect 5064 3031 6953 3048
tri 6953 3031 6970 3048 nw
tri 7014 3031 7031 3048 ne
rect 7031 3038 7092 3048
rect 7031 3031 7040 3038
rect 5064 3024 6946 3031
tri 6946 3024 6953 3031 nw
tri 7031 3024 7038 3031 ne
rect 7038 3024 7040 3031
rect 4946 3018 6940 3024
tri 6940 3018 6946 3024 nw
tri 7038 3022 7040 3024 ne
rect 4829 2962 4840 2987
rect 7126 3019 7132 3071
rect 7184 3019 7196 3071
rect 7248 3065 9326 3071
rect 7252 3031 7290 3065
rect 7324 3031 9208 3065
rect 9242 3031 9280 3065
rect 9314 3031 9326 3065
rect 7248 3025 9326 3031
rect 9617 3032 9620 3084
rect 9617 3026 9672 3032
rect 9848 3117 9859 3119
rect 9893 3117 9900 3119
rect 9848 3092 9900 3117
rect 9848 3031 9900 3040
rect 10089 4369 10135 4407
rect 10089 4335 10095 4369
rect 10129 4335 10135 4369
rect 10089 4297 10135 4335
rect 10089 4263 10095 4297
rect 10129 4263 10135 4297
rect 10089 4225 10135 4263
rect 10089 4191 10095 4225
rect 10129 4191 10135 4225
rect 10089 4153 10135 4191
rect 10089 4119 10095 4153
rect 10129 4119 10135 4153
rect 10089 4081 10135 4119
rect 10089 4047 10095 4081
rect 10129 4047 10135 4081
rect 10089 4009 10135 4047
rect 10089 3975 10095 4009
rect 10129 3975 10135 4009
rect 10089 3937 10135 3975
rect 10089 3903 10095 3937
rect 10129 3903 10135 3937
rect 10089 3865 10135 3903
rect 10089 3831 10095 3865
rect 10129 3831 10135 3865
rect 10089 3793 10135 3831
rect 10089 3759 10095 3793
rect 10129 3759 10135 3793
rect 10089 3721 10135 3759
rect 10089 3687 10095 3721
rect 10129 3687 10135 3721
rect 10089 3649 10135 3687
rect 10089 3615 10095 3649
rect 10129 3615 10135 3649
rect 10089 3577 10135 3615
rect 10089 3543 10095 3577
rect 10129 3543 10135 3577
rect 10089 3505 10135 3543
rect 10089 3471 10095 3505
rect 10129 3471 10135 3505
rect 10089 3433 10135 3471
rect 10089 3399 10095 3433
rect 10129 3399 10135 3433
rect 10089 3361 10135 3399
rect 10089 3327 10095 3361
rect 10129 3327 10135 3361
rect 10089 3289 10135 3327
rect 10089 3255 10095 3289
rect 10129 3255 10135 3289
rect 10089 3217 10135 3255
rect 10089 3183 10095 3217
rect 10129 3183 10135 3217
rect 10089 3145 10135 3183
rect 10089 3111 10095 3145
rect 10129 3111 10135 3145
rect 10277 3186 10323 4972
rect 10483 4859 10489 4911
rect 10541 4859 10553 4911
rect 10605 4859 10617 4911
rect 10669 4859 10682 4911
rect 10734 4859 10747 4911
rect 10799 4859 10812 4911
rect 10864 4859 10877 4911
rect 10929 4859 10942 4911
rect 10994 4859 11007 4911
rect 11059 4859 11965 4911
rect 12017 4859 12029 4911
rect 12081 4859 12093 4911
rect 12145 4859 12157 4911
rect 12209 4859 12221 4911
rect 12273 4859 12399 4911
rect 12451 4859 12493 4911
rect 12545 4859 12558 4911
tri 12559 4813 12587 4841 se
rect 12587 4819 12641 5251
tri 12641 5245 12647 5251 nw
tri 14704 5245 14710 5251 se
rect 14710 5245 14762 5251
tri 14696 5237 14704 5245 se
rect 14704 5237 14762 5245
tri 14762 5237 14823 5298 nw
tri 16424 5283 16439 5298 ne
rect 13046 5219 14744 5237
tri 14744 5219 14762 5237 nw
rect 13046 5190 14715 5219
tri 14715 5190 14744 5219 nw
rect 16439 5196 16491 5298
tri 16439 5190 16445 5196 ne
rect 16445 5190 16491 5196
rect 12587 4813 12632 4819
tri 12556 4810 12559 4813 se
rect 12559 4810 12632 4813
tri 12632 4810 12641 4819 nw
rect 12669 5112 12721 5118
rect 12669 5047 12721 5060
rect 12669 4982 12721 4995
rect 12669 4924 12675 4930
rect 12709 4924 12721 4930
rect 12669 4917 12721 4924
rect 12669 4851 12675 4865
rect 12709 4851 12721 4865
tri 12549 4803 12556 4810 se
rect 12556 4803 12610 4810
rect 10417 4797 12610 4803
rect 10417 4791 11121 4797
rect 10417 4765 10423 4791
rect 10457 4765 11121 4791
rect 10469 4745 11121 4765
rect 11173 4784 11851 4797
rect 11173 4750 11290 4784
rect 11324 4750 11372 4784
rect 11406 4750 11454 4784
rect 11488 4750 11536 4784
rect 11570 4750 11618 4784
rect 11652 4750 11700 4784
rect 11734 4750 11851 4784
rect 11173 4745 11851 4750
rect 11903 4745 12553 4797
rect 12605 4788 12610 4797
tri 12610 4788 12632 4810 nw
tri 12605 4783 12610 4788 nw
rect 12669 4785 12675 4799
rect 12709 4785 12721 4799
rect 10469 4727 12605 4745
rect 10469 4713 11121 4727
rect 10417 4711 11121 4713
rect 10417 4698 10423 4711
rect 10457 4698 11121 4711
rect 10469 4675 11121 4698
rect 11173 4708 11851 4727
rect 11173 4675 11290 4708
rect 10469 4674 11290 4675
rect 11324 4674 11372 4708
rect 11406 4674 11454 4708
rect 11488 4674 11536 4708
rect 11570 4674 11618 4708
rect 11652 4674 11700 4708
rect 11734 4675 11851 4708
rect 11903 4675 12553 4727
rect 11734 4674 12605 4675
rect 10469 4657 12605 4674
rect 10469 4646 11121 4657
rect 10417 4631 11121 4646
rect 11173 4632 11851 4657
rect 10469 4605 11121 4631
rect 11173 4605 11290 4632
rect 10469 4597 11130 4605
rect 11164 4598 11290 4605
rect 11324 4598 11372 4632
rect 11406 4598 11454 4632
rect 11488 4598 11536 4632
rect 11570 4598 11618 4632
rect 11652 4598 11700 4632
rect 11734 4605 11851 4632
rect 11903 4605 12553 4657
rect 11734 4598 11860 4605
rect 11164 4597 11860 4598
rect 11894 4597 12565 4605
rect 12599 4597 12605 4605
rect 10469 4587 12605 4597
rect 10469 4579 11121 4587
rect 10417 4565 11121 4579
rect 10469 4535 11121 4565
rect 11173 4555 11851 4587
rect 11173 4535 11290 4555
rect 10469 4518 11130 4535
rect 11164 4521 11290 4535
rect 11324 4521 11372 4555
rect 11406 4521 11454 4555
rect 11488 4521 11536 4555
rect 11570 4521 11618 4555
rect 11652 4521 11700 4555
rect 11734 4535 11851 4555
rect 11903 4535 12553 4587
rect 11734 4521 11860 4535
rect 11164 4518 11860 4521
rect 11894 4518 12565 4535
rect 12599 4518 12605 4535
rect 10469 4517 12605 4518
rect 10469 4513 11121 4517
rect 10417 4499 11121 4513
rect 10469 4465 11121 4499
rect 11173 4478 11851 4517
rect 11173 4465 11290 4478
rect 10469 4447 11130 4465
rect 11164 4447 11290 4465
rect 10417 4439 10423 4447
rect 10457 4439 11121 4447
rect 11173 4444 11290 4447
rect 11324 4444 11372 4478
rect 11406 4444 11454 4478
rect 11488 4444 11536 4478
rect 11570 4444 11618 4478
rect 11652 4444 11700 4478
rect 11734 4465 11851 4478
rect 11903 4465 12553 4517
rect 11734 4447 11860 4465
rect 11894 4447 12565 4465
rect 12599 4447 12605 4465
rect 11734 4444 11851 4447
rect 10417 4433 11121 4439
rect 10469 4395 11121 4433
rect 11173 4401 11851 4444
rect 11173 4395 11290 4401
rect 10469 4394 11290 4395
rect 10469 4381 11130 4394
rect 10417 4367 10423 4381
rect 10457 4377 11130 4381
rect 11164 4377 11290 4394
rect 10457 4367 11121 4377
rect 10469 4325 11121 4367
rect 11173 4367 11290 4377
rect 11324 4367 11372 4401
rect 11406 4367 11454 4401
rect 11488 4367 11536 4401
rect 11570 4367 11618 4401
rect 11652 4367 11700 4401
rect 11734 4395 11851 4401
rect 11903 4395 12553 4447
rect 11734 4394 12605 4395
rect 11734 4377 11860 4394
rect 11894 4377 12565 4394
rect 12599 4377 12605 4394
rect 11734 4367 11851 4377
rect 11173 4325 11851 4367
rect 11903 4325 12553 4377
rect 10469 4324 12605 4325
rect 10469 4315 11290 4324
rect 10417 4301 10423 4315
rect 10457 4307 11130 4315
rect 11164 4307 11290 4315
rect 10457 4301 11121 4307
rect 10469 4255 11121 4301
rect 11173 4290 11290 4307
rect 11324 4290 11372 4324
rect 11406 4290 11454 4324
rect 11488 4290 11536 4324
rect 11570 4290 11618 4324
rect 11652 4290 11700 4324
rect 11734 4315 12605 4324
rect 11734 4307 11860 4315
rect 11894 4307 12565 4315
rect 12599 4307 12605 4315
rect 11734 4290 11851 4307
rect 11173 4255 11851 4290
rect 11903 4255 12553 4307
rect 10469 4249 12605 4255
rect 10417 4247 12605 4249
rect 10417 4238 11290 4247
rect 10417 4236 11121 4238
rect 10417 4235 10423 4236
rect 10457 4235 11121 4236
rect 10469 4186 11121 4235
rect 11173 4213 11290 4238
rect 11324 4213 11372 4247
rect 11406 4213 11454 4247
rect 11488 4213 11536 4247
rect 11570 4213 11618 4247
rect 11652 4213 11700 4247
rect 11734 4238 12605 4247
rect 11734 4213 11851 4238
rect 11173 4186 11851 4213
rect 11903 4186 12553 4238
rect 10469 4183 12605 4186
rect 10417 4170 12605 4183
rect 10417 4169 11290 4170
rect 10469 4117 11121 4169
rect 11173 4136 11290 4169
rect 11324 4136 11372 4170
rect 11406 4136 11454 4170
rect 11488 4136 11536 4170
rect 11570 4136 11618 4170
rect 11652 4136 11700 4170
rect 11734 4169 12605 4170
rect 11734 4136 11851 4169
rect 11173 4117 11851 4136
rect 11903 4117 12553 4169
rect 10417 4111 12605 4117
rect 12669 4719 12675 4733
rect 12709 4719 12721 4733
rect 12669 4662 12721 4667
rect 12669 4653 12675 4662
rect 12709 4653 12721 4662
rect 12669 4588 12721 4601
rect 12669 4587 12675 4588
rect 12709 4587 12721 4588
rect 12669 4521 12721 4535
rect 12669 4455 12721 4469
rect 12669 4389 12721 4403
rect 12669 4331 12675 4337
rect 12709 4331 12721 4337
rect 12669 4323 12721 4331
rect 12669 4257 12675 4271
rect 12709 4257 12721 4271
rect 12669 4191 12675 4205
rect 12709 4191 12721 4205
rect 12669 4125 12675 4139
rect 12709 4125 12721 4139
rect 12669 4065 12721 4073
rect 12669 4059 12675 4065
rect 12709 4059 12721 4065
rect 10536 4003 10588 4055
rect 10640 4003 10657 4055
rect 10709 4003 10727 4055
rect 10779 4003 10797 4055
rect 10849 4003 10867 4055
rect 10919 4003 10937 4055
rect 10989 4003 11007 4055
rect 11059 4003 12399 4055
rect 12451 4003 12467 4055
rect 12519 4003 12558 4055
rect 12669 3993 12721 4007
rect 10391 3965 11254 3966
tri 11254 3965 11255 3966 sw
rect 10391 3959 11255 3965
rect 10443 3907 11121 3959
rect 11173 3956 11255 3959
tri 11255 3956 11264 3965 sw
rect 11173 3915 11264 3956
tri 11264 3915 11305 3956 sw
rect 11173 3907 11305 3915
rect 10391 3895 11305 3907
rect 10443 3874 11121 3895
tri 10443 3849 10468 3874 nw
tri 10532 3849 10557 3874 ne
rect 10557 3849 11121 3874
tri 10557 3848 10558 3849 ne
rect 10558 3848 11121 3849
rect 11173 3881 11305 3895
tri 11305 3881 11339 3915 sw
rect 11996 3905 12558 3966
rect 11173 3861 11339 3881
tri 11339 3861 11359 3881 sw
rect 10391 3836 10443 3843
tri 10558 3837 10569 3848 ne
rect 10569 3843 11121 3848
rect 11173 3843 11662 3861
rect 10569 3837 11662 3843
tri 11662 3837 11686 3861 sw
rect 11996 3853 12307 3905
rect 12359 3853 12558 3905
rect 12669 3927 12721 3941
rect 12669 3869 12721 3875
rect 10474 3836 10526 3837
tri 10526 3836 10527 3837 sw
tri 10569 3836 10570 3837 ne
rect 10570 3836 11686 3837
tri 11686 3836 11687 3837 sw
rect 10474 3831 10527 3836
rect 10526 3829 10527 3831
tri 10527 3829 10534 3836 sw
tri 11200 3829 11207 3836 ne
rect 11207 3829 11687 3836
tri 11687 3829 11694 3836 sw
rect 10526 3796 10534 3829
tri 10534 3796 10567 3829 sw
tri 11207 3796 11240 3829 ne
rect 11240 3796 11694 3829
tri 11694 3796 11727 3829 sw
rect 11996 3816 12558 3853
rect 10526 3790 11098 3796
tri 11240 3795 11241 3796 ne
rect 11241 3795 11532 3796
rect 10526 3779 10620 3790
rect 10474 3767 10620 3779
rect 10526 3756 10620 3767
rect 10654 3756 10692 3790
rect 10726 3756 10764 3790
rect 10798 3756 10836 3790
rect 10870 3756 10908 3790
rect 10942 3756 10980 3790
rect 11014 3756 11052 3790
rect 11086 3756 11098 3790
tri 11241 3756 11280 3795 ne
rect 11280 3756 11532 3795
rect 10526 3750 11098 3756
tri 11280 3750 11286 3756 ne
rect 11286 3750 11532 3756
rect 11996 3764 12307 3816
rect 12359 3764 12558 3816
rect 10526 3722 10539 3750
tri 10539 3722 10567 3750 nw
rect 11996 3727 12558 3764
rect 10526 3715 10527 3722
rect 10474 3710 10527 3715
tri 10527 3710 10539 3722 nw
rect 10391 3703 10443 3710
rect 10474 3709 10526 3710
tri 10526 3709 10527 3710 nw
tri 10569 3709 10570 3710 se
rect 10570 3709 11183 3710
tri 10558 3698 10569 3709 se
rect 10569 3703 11183 3709
rect 10569 3698 11121 3703
tri 10557 3697 10558 3698 se
rect 10558 3697 11121 3698
tri 10443 3672 10468 3697 sw
tri 10532 3672 10557 3697 se
rect 10557 3672 11121 3697
rect 10443 3651 11121 3672
rect 11173 3651 11183 3703
rect 10391 3639 11183 3651
rect 10443 3587 11121 3639
rect 11173 3587 11183 3639
rect 10391 3580 11183 3587
rect 11996 3675 12307 3727
rect 12359 3675 12558 3727
rect 12586 3835 12822 3841
rect 12586 3829 12770 3835
rect 12586 3795 12592 3829
rect 12626 3795 12770 3829
rect 12586 3783 12770 3795
rect 12586 3768 12822 3783
rect 12586 3756 12770 3768
rect 12586 3722 12592 3756
rect 12626 3722 12770 3756
rect 12586 3716 12770 3722
rect 12586 3710 12822 3716
rect 11996 3638 12558 3675
rect 11996 3586 12307 3638
rect 12359 3586 12558 3638
rect 11996 3580 12558 3586
rect 12661 3676 12715 3682
rect 12713 3624 12715 3676
rect 12661 3606 12715 3624
rect 12713 3554 12715 3606
rect 10536 3543 12558 3544
rect 10536 3491 10588 3543
rect 10640 3491 10657 3543
rect 10709 3491 10727 3543
rect 10779 3491 10797 3543
rect 10849 3491 10867 3543
rect 10919 3491 10937 3543
rect 10989 3491 11007 3543
rect 11059 3491 11207 3543
rect 11259 3491 11273 3543
rect 11325 3491 11339 3543
rect 11391 3491 11405 3543
rect 11457 3491 11471 3543
rect 11523 3491 11537 3543
rect 11589 3491 11603 3543
rect 11655 3491 11670 3543
rect 11722 3491 11737 3543
rect 11789 3491 12399 3543
rect 12451 3491 12467 3543
rect 12519 3491 12558 3543
rect 12661 3536 12715 3554
rect 12713 3484 12715 3536
rect 12661 3476 12675 3484
rect 12709 3476 12715 3484
rect 12661 3466 12715 3476
rect 10391 3447 12633 3454
rect 10443 3395 11121 3447
rect 11173 3395 11851 3447
rect 11903 3395 12581 3447
rect 10391 3383 12633 3395
rect 10443 3362 11121 3383
tri 10443 3337 10468 3362 nw
tri 10532 3337 10557 3362 ne
rect 10557 3337 11121 3362
tri 10557 3336 10558 3337 ne
rect 10558 3336 11121 3337
rect 10391 3324 10443 3331
tri 10558 3325 10569 3336 ne
rect 10569 3331 11121 3336
rect 11173 3331 11851 3383
rect 11903 3331 12581 3383
rect 10569 3325 12633 3331
rect 10474 3324 10526 3325
tri 10526 3324 10527 3325 sw
tri 10569 3324 10570 3325 ne
rect 10570 3324 12633 3325
rect 12713 3414 12715 3466
rect 12661 3396 12675 3414
rect 12709 3396 12715 3414
rect 12661 3395 12715 3396
rect 12713 3343 12715 3395
rect 12661 3324 12675 3343
rect 12709 3324 12715 3343
rect 10474 3319 10527 3324
rect 10526 3316 10527 3319
tri 10527 3316 10535 3324 sw
rect 10526 3284 10535 3316
tri 10535 3284 10567 3316 sw
rect 10526 3278 11266 3284
rect 10526 3267 10620 3278
rect 10474 3255 10620 3267
rect 10526 3244 10620 3255
rect 10654 3244 10692 3278
rect 10726 3244 10764 3278
rect 10798 3244 10836 3278
rect 10870 3244 10908 3278
rect 10942 3244 10980 3278
rect 11014 3244 11052 3278
rect 11086 3244 11266 3278
rect 10526 3238 11266 3244
rect 11828 3238 11880 3284
rect 11881 3239 11882 3283
rect 11918 3239 11919 3283
rect 11920 3278 12414 3284
rect 11920 3244 12008 3278
rect 12042 3244 12080 3278
rect 12114 3244 12152 3278
rect 12186 3244 12224 3278
rect 12258 3244 12296 3278
rect 12330 3244 12368 3278
rect 12402 3244 12414 3278
rect 11920 3238 12414 3244
rect 12448 3278 12525 3284
rect 12448 3238 12473 3278
rect 10526 3236 10565 3238
tri 10565 3236 10567 3238 nw
tri 12448 3236 12450 3238 ne
rect 12450 3236 12473 3238
rect 10474 3197 10526 3203
tri 10526 3197 10565 3236 nw
tri 12450 3213 12473 3236 ne
rect 12473 3214 12525 3226
tri 10323 3186 10326 3189 sw
rect 10277 3180 10326 3186
tri 10326 3180 10332 3186 sw
rect 10277 3162 10332 3180
tri 10332 3162 10350 3180 sw
tri 10531 3162 10549 3180 se
rect 10549 3179 12326 3180
tri 12326 3179 12327 3180 sw
rect 10549 3162 12327 3179
rect 10277 3156 12327 3162
tri 12327 3156 12350 3179 sw
tri 12450 3156 12473 3179 se
rect 12713 3272 12715 3324
rect 12661 3270 12715 3272
rect 12661 3253 12675 3270
rect 12709 3253 12715 3270
rect 12713 3201 12715 3253
rect 12473 3156 12525 3162
rect 10277 3154 12350 3156
tri 12350 3154 12352 3156 sw
tri 12448 3154 12450 3156 se
rect 12450 3154 12525 3156
rect 10277 3147 12525 3154
tri 10277 3134 10290 3147 ne
rect 10290 3134 12525 3147
tri 10290 3116 10308 3134 ne
rect 10308 3116 10551 3134
tri 10551 3116 10569 3134 nw
tri 12306 3116 12324 3134 ne
rect 12324 3116 12525 3134
tri 12324 3114 12326 3116 ne
rect 12326 3114 12525 3116
rect 10089 3072 10135 3111
tri 12326 3110 12330 3114 ne
rect 12330 3110 12525 3114
rect 12581 3191 12633 3198
rect 12581 3127 12633 3139
tri 10575 3100 10581 3106 se
rect 10581 3100 11894 3106
tri 10563 3088 10575 3100 se
rect 10575 3088 11046 3100
rect 10089 3038 10095 3072
rect 10129 3038 10135 3072
rect 7248 3024 7373 3025
tri 7373 3024 7374 3025 nw
rect 7248 3019 7368 3024
tri 7368 3019 7373 3024 nw
tri 10083 2999 10089 3005 se
rect 10089 2999 10135 3038
rect 7040 2980 7092 2986
tri 10064 2980 10083 2999 se
rect 10083 2980 10095 2999
tri 10055 2971 10064 2980 se
rect 10064 2971 10095 2980
tri 9602 2970 9603 2971 se
rect 9603 2970 10095 2971
tri 9597 2965 9602 2970 se
rect 9602 2965 10095 2970
rect 10129 2965 10135 2999
rect 4829 2949 4892 2962
tri 9591 2959 9597 2965 se
rect 9597 2959 10135 2965
tri 9585 2953 9591 2959 se
rect 9591 2953 10135 2959
tri 9584 2952 9585 2953 se
rect 9585 2952 10135 2953
rect 4829 2943 4840 2949
rect 4829 2909 4835 2943
rect 4829 2897 4840 2909
rect 5012 2944 7142 2952
tri 7142 2944 7150 2952 sw
rect 5012 2910 7150 2944
tri 7150 2910 7184 2944 sw
rect 5012 2900 7184 2910
tri 7184 2900 7194 2910 sw
rect 7280 2900 8783 2952
rect 8835 2900 8847 2952
rect 8899 2900 9282 2952
tri 9576 2944 9584 2952 se
rect 9584 2944 10135 2952
tri 9554 2922 9576 2944 se
rect 9576 2922 10135 2944
rect 10391 3066 11046 3088
rect 11080 3066 11118 3100
rect 11152 3066 11776 3100
rect 11810 3066 11848 3100
rect 11882 3066 11894 3100
rect 12581 3068 12633 3075
rect 12661 3190 12715 3201
rect 12661 3182 12675 3190
rect 12709 3182 12715 3190
rect 12713 3130 12715 3182
rect 12661 3111 12715 3130
rect 10391 3063 11894 3066
rect 10443 3060 11894 3063
tri 10443 3035 10468 3060 nw
rect 12713 3059 12715 3111
rect 12661 3040 12715 3059
rect 10391 2999 10443 3011
rect 10536 2979 10588 3031
rect 10640 2979 10657 3031
rect 10709 2979 10727 3031
rect 10779 2979 10797 3031
rect 10849 2979 10867 3031
rect 10919 2979 10937 3031
rect 10989 2979 11007 3031
rect 11059 2979 11207 3031
rect 11259 2979 11273 3031
rect 11325 2979 11339 3031
rect 11391 2979 11405 3031
rect 11457 2979 11471 3031
rect 11523 2979 11537 3031
rect 11589 2979 11603 3031
rect 11655 2979 11670 3031
rect 11722 2979 11737 3031
rect 11789 2979 11965 3031
rect 12017 2979 12029 3031
rect 12081 2979 12093 3031
rect 12145 2979 12157 3031
rect 12209 2979 12221 3031
rect 12273 2979 12558 3031
rect 12713 2988 12715 3040
rect 12661 2982 12715 2988
tri 10443 2950 10468 2975 sw
rect 10443 2947 11894 2950
rect 10391 2944 11894 2947
rect 10391 2922 11046 2944
tri 9551 2919 9554 2922 se
rect 9554 2919 10135 2922
tri 10563 2919 10566 2922 ne
rect 10566 2919 11046 2922
tri 9542 2910 9551 2919 se
rect 9551 2910 9616 2919
tri 9616 2910 9625 2919 nw
tri 10566 2910 10575 2919 ne
rect 10575 2910 11046 2919
rect 11080 2910 11118 2944
rect 11152 2910 11776 2944
rect 11810 2910 11848 2944
rect 11882 2910 11894 2944
tri 9532 2900 9542 2910 se
rect 9542 2904 9610 2910
tri 9610 2904 9616 2910 nw
tri 10575 2904 10581 2910 ne
rect 10581 2904 11894 2910
tri 13037 2904 13046 2913 se
rect 13046 2904 13093 5190
tri 13093 5165 13118 5190 nw
tri 16445 5165 16470 5190 ne
rect 16470 5165 16491 5190
tri 16470 5162 16473 5165 ne
rect 16473 5162 16491 5165
tri 16491 5162 16548 5219 sw
rect 13873 5046 13879 5162
rect 13995 5046 14001 5162
tri 16473 5159 16476 5162 ne
rect 16476 5157 16548 5162
tri 16548 5157 16553 5162 sw
rect 16476 5106 16553 5157
rect 9542 2900 9606 2904
tri 9606 2900 9610 2904 nw
tri 13033 2900 13037 2904 se
rect 13037 2900 13093 2904
rect 4829 2884 4892 2897
rect 4829 2865 4840 2884
tri 7120 2871 7149 2900 ne
rect 7149 2871 7194 2900
tri 7194 2871 7223 2900 sw
tri 9503 2871 9532 2900 se
rect 9532 2871 9551 2900
rect 4829 2831 4835 2865
rect 4869 2831 4892 2832
rect 4829 2818 4892 2831
tri 7149 2826 7194 2871 ne
rect 7194 2845 9551 2871
tri 9551 2845 9606 2900 nw
tri 13024 2891 13033 2900 se
rect 13033 2891 13093 2900
tri 9642 2866 9667 2891 se
rect 9667 2885 10551 2891
tri 10551 2885 10557 2891 sw
tri 13018 2885 13024 2891 se
rect 13024 2885 13093 2891
rect 9667 2866 10557 2885
tri 10557 2866 10576 2885 sw
tri 12385 2866 12404 2885 se
rect 12404 2866 13093 2885
tri 9621 2845 9642 2866 se
rect 9642 2859 13093 2866
rect 9642 2845 9667 2859
rect 7194 2826 9525 2845
tri 7194 2819 7201 2826 ne
rect 7201 2819 9525 2826
tri 9525 2819 9551 2845 nw
tri 9616 2840 9621 2845 se
rect 9621 2840 9667 2845
tri 9667 2840 9686 2859 nw
tri 10527 2840 10546 2859 ne
rect 10546 2842 13093 2859
rect 10546 2840 12405 2842
tri 9595 2819 9616 2840 se
rect 9616 2819 9641 2840
rect 4829 2787 4840 2818
tri 9590 2814 9595 2819 se
rect 9595 2814 9641 2819
tri 9641 2814 9667 2840 nw
tri 10546 2820 10566 2840 ne
rect 10566 2820 12405 2840
tri 12405 2820 12427 2842 nw
tri 9589 2813 9590 2814 se
rect 9590 2813 9640 2814
tri 9640 2813 9641 2814 nw
tri 9580 2804 9589 2813 se
rect 9589 2804 9631 2813
tri 9631 2804 9640 2813 nw
tri 10465 2804 10474 2813 se
rect 10474 2807 10526 2813
tri 9578 2802 9580 2804 se
rect 9580 2802 9629 2804
tri 9629 2802 9631 2804 nw
tri 10463 2802 10465 2804 se
rect 10465 2802 10474 2804
tri 9571 2795 9578 2802 se
rect 9578 2795 9622 2802
tri 9622 2795 9629 2802 nw
tri 10456 2795 10463 2802 se
rect 10463 2795 10474 2802
tri 6951 2789 6957 2795 se
rect 6957 2789 6963 2795
rect 4829 2753 4835 2787
rect 4869 2753 4892 2766
rect 4829 2752 4892 2753
rect 4829 2709 4840 2752
rect 4946 2783 6963 2789
rect 4946 2749 4958 2783
rect 4992 2749 5030 2783
rect 5064 2749 6963 2783
rect 4946 2743 6963 2749
rect 7015 2743 7027 2795
rect 7079 2743 7088 2795
tri 9567 2791 9571 2795 se
rect 9571 2791 9618 2795
tri 9618 2791 9622 2795 nw
tri 10452 2791 10456 2795 se
rect 10456 2791 10474 2795
rect 7126 2739 7132 2791
rect 7184 2739 7196 2791
rect 7248 2785 9599 2791
rect 7252 2751 7290 2785
rect 7324 2751 9147 2785
rect 9181 2751 9219 2785
rect 9253 2772 9599 2785
tri 9599 2772 9618 2791 nw
tri 10433 2772 10452 2791 se
rect 10452 2772 10474 2791
rect 9253 2768 9595 2772
tri 9595 2768 9599 2772 nw
tri 9677 2768 9681 2772 se
rect 9681 2768 10474 2772
rect 9253 2766 9593 2768
tri 9593 2766 9595 2768 nw
tri 9675 2766 9677 2768 se
rect 9677 2766 10474 2768
rect 9253 2751 9572 2766
rect 7248 2745 9572 2751
tri 9572 2745 9593 2766 nw
tri 9654 2745 9675 2766 se
rect 9675 2755 10474 2766
tri 12466 2806 12473 2813 se
rect 12473 2807 12525 2813
tri 10526 2802 10530 2806 sw
tri 12462 2802 12466 2806 se
rect 12466 2802 12473 2806
rect 10526 2772 10530 2802
tri 10530 2772 10560 2802 sw
tri 12432 2772 12462 2802 se
rect 12462 2772 12473 2802
rect 10526 2766 11266 2772
rect 10526 2755 10620 2766
rect 9675 2745 10620 2755
rect 7248 2739 7374 2745
tri 7374 2739 7380 2745 nw
tri 9648 2739 9654 2745 se
rect 9654 2743 10620 2745
rect 9654 2739 10474 2743
tri 9641 2732 9648 2739 se
rect 9648 2732 10474 2739
tri 9639 2730 9641 2732 se
rect 9641 2730 10474 2732
tri 9635 2726 9639 2730 se
rect 9639 2726 10474 2730
tri 9621 2712 9635 2726 se
rect 9635 2712 9687 2726
tri 9687 2712 9701 2726 nw
tri 10433 2712 10447 2726 ne
rect 10447 2712 10474 2726
rect 4829 2675 4835 2709
rect 4869 2686 4892 2700
rect 4829 2634 4840 2675
rect 5012 2660 5345 2712
rect 5397 2660 5409 2712
rect 5461 2660 7014 2712
tri 9619 2710 9621 2712 se
rect 9621 2710 9685 2712
tri 9685 2710 9687 2712 nw
tri 10447 2710 10449 2712 ne
rect 10449 2710 10474 2712
rect 7280 2658 8638 2710
rect 8690 2658 8702 2710
rect 8754 2658 9282 2710
tri 9605 2696 9619 2710 se
rect 9619 2696 9671 2710
tri 9671 2696 9685 2710 nw
tri 10449 2696 10463 2710 ne
rect 10463 2696 10474 2710
tri 9581 2672 9605 2696 se
rect 9605 2685 9660 2696
tri 9660 2685 9671 2696 nw
tri 10463 2685 10474 2696 ne
rect 10526 2732 10620 2743
rect 10654 2732 10692 2766
rect 10726 2732 10764 2766
rect 10798 2732 10836 2766
rect 10870 2732 10908 2766
rect 10942 2732 10980 2766
rect 11014 2732 11052 2766
rect 11086 2732 11266 2766
rect 10526 2726 11266 2732
rect 11996 2766 12473 2772
rect 11996 2732 12008 2766
rect 12042 2732 12080 2766
rect 12114 2732 12152 2766
rect 12186 2732 12224 2766
rect 12258 2732 12296 2766
rect 12330 2732 12368 2766
rect 12402 2732 12440 2766
rect 12474 2743 12525 2755
rect 11996 2726 12473 2732
rect 10526 2696 10530 2726
tri 10530 2696 10560 2726 nw
tri 12432 2696 12462 2726 ne
rect 12462 2696 12473 2726
tri 10526 2692 10530 2696 nw
tri 12462 2692 12466 2696 ne
rect 12466 2692 12473 2696
rect 10474 2685 10526 2691
tri 12466 2685 12473 2692 ne
rect 12473 2685 12525 2691
rect 12581 2807 12633 2814
rect 12581 2743 12633 2755
rect 9605 2684 9659 2685
tri 9659 2684 9660 2685 nw
rect 12581 2684 12633 2691
rect 12661 2796 12713 2802
rect 12661 2714 12713 2744
rect 9605 2672 9647 2684
tri 9647 2672 9659 2684 nw
tri 9569 2660 9581 2672 se
rect 9581 2660 9635 2672
tri 9635 2660 9647 2672 nw
tri 9567 2658 9569 2660 se
rect 9569 2658 9633 2660
tri 9633 2658 9635 2660 nw
rect 4829 2631 4892 2634
rect 4829 2597 4835 2631
rect 4869 2620 4892 2631
tri 9531 2622 9567 2658 se
rect 9567 2622 9597 2658
tri 9597 2622 9633 2658 nw
rect 12661 2632 12713 2662
tri 9513 2604 9531 2622 se
rect 9531 2604 9569 2622
rect 4829 2568 4840 2597
tri 9503 2594 9513 2604 se
rect 9513 2594 9569 2604
tri 9569 2594 9597 2622 nw
tri 9499 2590 9503 2594 se
rect 9503 2590 9565 2594
tri 9565 2590 9569 2594 nw
tri 10577 2590 10581 2594 se
rect 10581 2590 11894 2594
tri 7278 2588 7280 2590 se
rect 7280 2588 9334 2590
rect 9336 2589 9372 2590
tri 7277 2587 7278 2588 se
rect 7278 2587 9334 2588
rect 4829 2554 4892 2568
rect 4829 2553 4840 2554
rect 4829 2519 4835 2553
rect 5012 2535 6638 2587
rect 6690 2535 6702 2587
rect 6754 2535 6825 2587
tri 6825 2584 6828 2587 sw
tri 7274 2584 7277 2587 se
rect 7277 2584 9334 2587
rect 7014 2538 9334 2584
rect 9335 2539 9373 2589
rect 9374 2588 9563 2590
tri 9563 2588 9565 2590 nw
tri 10575 2588 10577 2590 se
rect 10577 2588 11894 2590
rect 9374 2576 9551 2588
tri 9551 2576 9563 2588 nw
tri 10563 2576 10575 2588 se
rect 10575 2576 11046 2588
rect 9374 2554 9529 2576
tri 9529 2554 9551 2576 nw
rect 10391 2554 11046 2576
rect 11080 2554 11118 2588
rect 11152 2554 11776 2588
rect 11810 2554 11848 2588
rect 11882 2554 11894 2588
rect 9374 2546 9521 2554
tri 9521 2546 9529 2554 nw
rect 10391 2551 11894 2554
rect 10443 2548 11894 2551
rect 12661 2549 12713 2580
rect 9336 2538 9372 2539
rect 9374 2538 9513 2546
tri 9513 2538 9521 2546 nw
tri 6825 2535 6828 2538 nw
rect 4829 2502 4840 2519
rect 10443 2538 10458 2548
tri 10458 2538 10468 2548 nw
tri 10443 2523 10458 2538 nw
rect 4829 2488 4892 2502
rect 4829 2476 4840 2488
rect 4829 2442 4835 2476
rect 7040 2458 7046 2510
rect 7098 2458 7110 2510
rect 7162 2504 7331 2510
tri 7331 2504 7337 2510 sw
rect 7162 2498 7337 2504
rect 7162 2464 7218 2498
rect 7252 2464 7290 2498
rect 7324 2474 7337 2498
tri 7337 2474 7367 2504 sw
rect 10391 2487 10443 2499
rect 7324 2466 7367 2474
tri 7367 2466 7375 2474 sw
rect 7324 2464 10360 2466
rect 7162 2460 10360 2464
rect 7162 2458 9208 2460
tri 7317 2451 7324 2458 ne
rect 7324 2451 9208 2458
rect 4829 2436 4840 2442
rect 4829 2430 4892 2436
rect 4946 2445 6919 2451
rect 4637 2416 4689 2422
rect 4946 2411 4958 2445
rect 4992 2411 5030 2445
rect 5064 2430 6919 2445
tri 6919 2430 6940 2451 sw
tri 7324 2430 7345 2451 ne
rect 7345 2430 9208 2451
rect 5064 2424 7132 2430
rect 5064 2411 6970 2424
rect 4946 2405 6970 2411
tri 6899 2390 6914 2405 ne
rect 6914 2390 6970 2405
rect 7004 2390 7042 2424
rect 7076 2390 7132 2424
tri 6914 2388 6916 2390 ne
rect 6916 2388 7132 2390
rect 3070 2304 3122 2326
tri 2983 2260 2990 2267 se
rect 2990 2261 3042 2267
tri 2982 2259 2983 2260 se
rect 2983 2259 2990 2260
tri 2980 2257 2982 2259 se
rect 2982 2257 2990 2259
tri 2949 2226 2980 2257 se
rect 2980 2226 2990 2257
rect 1792 2223 1813 2226
tri 1813 2223 1816 2226 sw
tri 2454 2223 2457 2226 se
rect 2457 2223 2527 2226
rect 1792 2222 1816 2223
tri 1816 2222 1817 2223 sw
tri 2453 2222 2454 2223 se
rect 2454 2222 2527 2223
rect 1792 1908 2527 2222
rect 2857 2180 2909 2226
rect 2910 2181 2911 2225
rect 2947 2181 2948 2225
rect 2949 2209 2990 2226
rect 2949 2197 3042 2209
rect 2949 2180 2990 2197
tri 2949 2151 2978 2180 ne
rect 2978 2151 2990 2180
tri 2978 2148 2981 2151 ne
rect 2981 2148 2990 2151
tri 2981 2144 2985 2148 ne
rect 2985 2145 2990 2148
rect 2985 2144 3042 2145
tri 2985 2139 2990 2144 ne
rect 2990 2139 3042 2144
rect 4258 2338 4310 2353
rect 4258 2271 4310 2286
rect 3070 2230 3122 2252
rect 3070 2156 3122 2178
tri 2829 2110 2830 2111 se
rect 2830 2110 2882 2111
tri 2821 2102 2829 2110 se
rect 2829 2105 2882 2110
rect 2829 2102 2830 2105
tri 2818 2099 2821 2102 se
rect 2821 2099 2830 2102
tri 2796 2077 2818 2099 se
rect 2818 2077 2830 2099
tri 2789 2070 2796 2077 se
rect 2796 2070 2830 2077
rect 2789 2053 2830 2070
rect 3544 2267 3590 2269
tri 3590 2267 3592 2269 sw
rect 3544 2260 3592 2267
tri 3592 2260 3599 2267 sw
rect 3544 2259 3599 2260
tri 3599 2259 3600 2260 sw
rect 4418 2384 4470 2388
tri 4470 2384 4474 2388 sw
tri 6916 2384 6920 2388 ne
rect 6920 2384 7132 2388
rect 4418 2382 4474 2384
rect 4470 2378 4474 2382
tri 4474 2378 4480 2384 sw
tri 6920 2378 6926 2384 ne
rect 6926 2378 7132 2384
rect 7184 2378 7196 2430
rect 7248 2378 7254 2430
tri 7345 2426 7349 2430 ne
rect 7349 2426 9208 2430
rect 9242 2426 9280 2460
rect 9314 2432 10360 2460
rect 9314 2426 9385 2432
tri 7349 2420 7355 2426 ne
rect 7355 2420 9385 2426
tri 9385 2420 9397 2432 nw
tri 10292 2420 10304 2432 ne
rect 10304 2420 10360 2432
tri 10304 2404 10320 2420 ne
rect 10320 2404 10360 2420
rect 10536 2467 10588 2519
rect 10640 2467 10657 2519
rect 10709 2467 10727 2519
rect 10779 2467 10797 2519
rect 10849 2467 10867 2519
rect 10919 2467 10937 2519
rect 10989 2467 11007 2519
rect 11059 2467 11207 2519
rect 11259 2467 11273 2519
rect 11325 2467 11339 2519
rect 11391 2467 11405 2519
rect 11457 2467 11471 2519
rect 11523 2467 11537 2519
rect 11589 2467 11603 2519
rect 11655 2467 11670 2519
rect 11722 2467 11737 2519
rect 11789 2467 11965 2519
rect 12017 2467 12029 2519
rect 12081 2467 12093 2519
rect 12145 2467 12157 2519
rect 12209 2467 12221 2519
rect 12273 2467 12558 2519
rect 12661 2491 12713 2497
rect 12910 2468 12950 2588
rect 12910 2467 12983 2468
tri 12983 2467 12984 2468 nw
rect 12910 2463 12979 2467
tri 12979 2463 12983 2467 nw
tri 10443 2438 10468 2463 sw
rect 12910 2457 12973 2463
tri 12973 2457 12979 2463 nw
tri 12891 2438 12910 2457 se
rect 12910 2438 12950 2457
rect 10443 2435 11894 2438
rect 10391 2432 11894 2435
rect 10391 2410 11046 2432
rect 9620 2397 9672 2404
tri 10320 2398 10326 2404 ne
tri 9616 2378 9620 2382 se
rect 4470 2357 4480 2378
tri 4480 2357 4501 2378 sw
tri 9595 2357 9616 2378 se
rect 9616 2357 9620 2378
rect 4470 2352 4803 2357
tri 4803 2352 4808 2357 sw
tri 9590 2352 9595 2357 se
rect 9595 2352 9620 2357
rect 4470 2332 4808 2352
tri 4808 2332 4828 2352 sw
rect 4470 2330 4828 2332
rect 4418 2318 4828 2330
rect 4470 2311 4828 2318
tri 4470 2277 4504 2311 nw
tri 4783 2277 4817 2311 ne
rect 4817 2300 4828 2311
tri 4828 2300 4860 2332 sw
rect 5012 2302 6637 2352
tri 6637 2348 6641 2352 sw
tri 9586 2348 9590 2352 se
rect 9590 2348 9620 2352
rect 7014 2342 7053 2348
tri 7053 2342 7059 2348 sw
rect 9282 2345 9620 2348
rect 10326 2392 10360 2404
tri 11016 2398 11028 2410 ne
rect 11028 2398 11046 2410
rect 11080 2398 11118 2432
rect 11152 2410 11776 2432
rect 11152 2398 11170 2410
tri 11170 2398 11182 2410 nw
tri 11746 2398 11758 2410 ne
rect 11758 2398 11776 2410
rect 11810 2398 11848 2432
rect 11882 2398 11894 2432
tri 12876 2423 12891 2438 se
rect 12891 2423 12950 2438
tri 12950 2434 12973 2457 nw
tri 10360 2392 10366 2398 sw
tri 11028 2392 11034 2398 ne
rect 11034 2392 11164 2398
tri 11164 2392 11170 2398 nw
tri 11758 2392 11764 2398 ne
rect 11764 2392 11894 2398
tri 12110 2392 12141 2423 se
rect 12141 2392 12950 2423
rect 7014 2302 7059 2342
tri 7059 2302 7099 2342 sw
rect 9282 2333 9672 2345
rect 10172 2367 10224 2373
rect 9282 2302 9620 2333
rect 5012 2301 6638 2302
tri 6638 2301 6639 2302 nw
tri 7033 2301 7034 2302 ne
rect 7034 2301 7099 2302
tri 7099 2301 7100 2302 sw
tri 9593 2301 9594 2302 ne
rect 9594 2301 9620 2302
rect 5012 2300 6637 2301
tri 6637 2300 6638 2301 nw
tri 7034 2300 7035 2301 ne
rect 7035 2300 7100 2301
rect 4817 2289 4860 2300
tri 4860 2289 4871 2300 sw
tri 7035 2289 7046 2300 ne
rect 7046 2289 7100 2300
tri 7100 2289 7112 2301 sw
tri 9594 2289 9606 2301 ne
rect 9606 2289 9620 2301
rect 4817 2277 4871 2289
tri 4871 2277 4883 2289 sw
tri 7046 2277 7058 2289 ne
rect 7058 2277 7112 2289
tri 7112 2277 7124 2289 sw
tri 9606 2277 9618 2289 ne
rect 9618 2281 9620 2289
tri 10160 2329 10172 2341 se
tri 10133 2302 10160 2329 se
rect 10160 2315 10172 2329
rect 10326 2364 10366 2392
tri 10366 2364 10394 2392 sw
tri 12083 2365 12110 2392 se
rect 12110 2383 12950 2392
rect 12110 2365 12141 2383
tri 12141 2365 12159 2383 nw
tri 12082 2364 12083 2365 se
rect 12083 2364 12140 2365
tri 12140 2364 12141 2365 nw
rect 10326 2342 12118 2364
tri 12118 2342 12140 2364 nw
rect 10326 2329 12105 2342
tri 12105 2329 12118 2342 nw
rect 12473 2336 12525 2342
rect 10160 2303 10224 2315
rect 10160 2302 10172 2303
tri 10132 2301 10133 2302 se
rect 10133 2301 10172 2302
tri 10122 2291 10132 2301 se
rect 10132 2291 10172 2301
tri 9903 2289 9905 2291 se
rect 9905 2289 10172 2291
rect 9618 2277 9672 2281
tri 9891 2277 9903 2289 se
rect 9903 2277 10172 2289
tri 4817 2266 4828 2277 ne
rect 4828 2266 4883 2277
tri 4883 2266 4894 2277 sw
tri 7058 2266 7069 2277 ne
rect 7069 2266 7124 2277
rect 4418 2260 4470 2266
tri 4828 2260 4834 2266 ne
rect 4834 2260 4894 2266
tri 4894 2260 4900 2266 sw
tri 7069 2260 7075 2266 ne
rect 7075 2262 7124 2266
tri 7124 2262 7139 2277 sw
tri 9618 2275 9620 2277 ne
rect 9620 2275 9672 2277
tri 9889 2275 9891 2277 se
rect 9891 2275 10172 2277
tri 9876 2262 9889 2275 se
rect 9889 2262 10172 2275
rect 7075 2260 9548 2262
rect 3544 2257 3600 2259
rect 3544 2223 3550 2257
rect 3584 2225 3600 2257
tri 3600 2225 3634 2259 sw
tri 4834 2243 4851 2260 ne
rect 4851 2243 4900 2260
tri 4900 2243 4917 2260 sw
tri 7075 2243 7092 2260 ne
rect 7092 2243 9548 2260
tri 9548 2243 9567 2262 sw
tri 9857 2243 9876 2262 se
rect 9876 2251 10172 2262
rect 10474 2295 10526 2301
rect 9876 2245 10224 2251
rect 10391 2283 10443 2289
rect 9876 2243 9923 2245
tri 9923 2243 9925 2245 nw
tri 4851 2227 4867 2243 ne
rect 4867 2236 4917 2243
tri 4917 2236 4924 2243 sw
tri 7092 2236 7099 2243 ne
rect 7099 2236 9567 2243
rect 4867 2227 4924 2236
tri 4924 2227 4933 2236 sw
tri 7099 2227 7108 2236 ne
rect 7108 2227 9567 2236
tri 9567 2227 9583 2243 sw
tri 9853 2239 9857 2243 se
rect 9857 2239 9919 2243
tri 9919 2239 9923 2243 nw
rect 9853 2227 9900 2239
rect 3584 2223 3634 2225
rect 3544 2207 3634 2223
tri 3634 2207 3652 2225 sw
rect 4258 2213 4310 2219
tri 4867 2213 4881 2227 ne
rect 4881 2216 4933 2227
tri 4933 2216 4944 2227 sw
tri 7108 2216 7119 2227 ne
rect 7119 2216 9583 2227
tri 9583 2216 9594 2227 sw
rect 4881 2213 4944 2216
tri 4944 2213 4947 2216 sw
tri 9528 2213 9531 2216 ne
rect 9531 2213 9594 2216
tri 4881 2207 4887 2213 ne
rect 4887 2207 4947 2213
tri 4947 2207 4953 2213 sw
rect 5055 2207 6940 2213
rect 3544 2200 3652 2207
tri 3652 2200 3659 2207 sw
tri 4887 2200 4894 2207 ne
rect 4894 2200 4953 2207
tri 4953 2200 4960 2207 sw
rect 3544 2191 3659 2200
tri 3659 2191 3668 2200 sw
tri 4894 2191 4903 2200 ne
rect 4903 2191 4960 2200
rect 3544 2185 3884 2191
rect 3544 2151 3550 2185
rect 3584 2151 3884 2185
rect 3544 2139 3884 2151
rect 3936 2139 3948 2191
rect 4000 2139 4012 2191
rect 4064 2139 4070 2191
tri 4903 2180 4914 2191 ne
tri 3220 2111 3236 2127 ne
rect 3236 2111 3306 2127
tri 3236 2106 3241 2111 ne
rect 3241 2106 3306 2111
rect 3070 2098 3122 2104
rect 2789 2041 2882 2053
rect 2789 2024 2830 2041
tri 2789 2002 2811 2024 ne
rect 2811 2002 2830 2024
tri 2811 1988 2825 2002 ne
rect 2825 1989 2830 2002
rect 2825 1988 2882 1989
tri 2825 1984 2829 1988 ne
rect 2829 1984 2882 1988
tri 2829 1983 2830 1984 ne
rect 2830 1983 2882 1984
rect 3070 1990 3122 1996
tri 2985 1950 2990 1955 se
rect 2990 1950 3042 1955
tri 2984 1949 2985 1950 se
rect 2985 1949 3042 1950
tri 2962 1927 2984 1949 se
rect 2984 1927 2990 1949
tri 2949 1914 2962 1927 se
rect 2962 1914 2990 1927
rect 1792 1886 1795 1908
tri 1795 1886 1817 1908 nw
tri 2453 1886 2475 1908 ne
rect 2475 1886 2527 1908
tri 1792 1883 1795 1886 nw
tri 2475 1883 2478 1886 ne
rect 1663 1833 1669 1867
rect 1703 1833 1709 1867
rect 1663 1794 1709 1833
rect 1820 1811 2032 1863
rect 2084 1811 2096 1863
rect 2148 1811 2160 1863
rect 2212 1811 2224 1863
rect 2276 1811 2288 1863
rect 2340 1811 2403 1863
rect 1663 1760 1669 1794
rect 1703 1760 1709 1794
rect 1663 1721 1709 1760
rect 1663 1687 1669 1721
rect 1703 1687 1709 1721
rect 1663 1648 1709 1687
rect 1663 1614 1669 1648
rect 1703 1614 1709 1648
rect 1663 1575 1709 1614
rect 1663 1541 1669 1575
rect 1703 1541 1709 1575
rect 1663 1502 1709 1541
rect 1663 1468 1669 1502
rect 1703 1468 1709 1502
rect 1663 1429 1709 1468
rect 1663 1395 1669 1429
rect 1703 1395 1709 1429
tri 1792 1789 1794 1791 sw
tri 2476 1789 2478 1791 se
rect 2478 1789 2527 1886
rect 2882 1897 2990 1914
rect 2882 1885 3042 1897
rect 2882 1868 2990 1885
tri 2949 1852 2965 1868 ne
rect 2965 1852 2990 1868
tri 2965 1840 2977 1852 ne
rect 2977 1840 2990 1852
rect 2830 1834 2882 1840
tri 2820 1789 2830 1799 se
rect 1792 1766 1794 1789
tri 1794 1766 1817 1789 sw
tri 2453 1766 2476 1789 se
rect 2476 1766 2527 1789
rect 1792 1708 2527 1766
tri 2789 1758 2820 1789 se
rect 2820 1782 2830 1789
tri 2977 1829 2988 1840 ne
rect 2988 1833 2990 1840
rect 2988 1829 3042 1833
tri 2988 1827 2990 1829 ne
rect 2990 1827 3042 1829
rect 4258 1990 4310 1996
rect 3932 1966 4150 1972
rect 3220 1952 3306 1953
rect 3070 1895 3122 1938
rect 2820 1770 2882 1782
rect 2820 1758 2830 1770
rect 3070 1801 3122 1843
rect 3932 1914 4098 1966
rect 3932 1902 4150 1914
rect 3932 1850 4098 1902
rect 3220 1823 3306 1824
rect 3932 1802 4150 1850
rect 4258 1875 4310 1938
rect 4914 1880 4960 2191
rect 5055 2173 5067 2207
rect 5101 2173 5139 2207
rect 5173 2193 6940 2207
tri 6940 2193 6960 2213 sw
tri 9531 2193 9551 2213 ne
rect 9551 2193 9594 2213
tri 9594 2193 9617 2216 sw
rect 9853 2193 9859 2227
rect 9893 2220 9900 2227
tri 9900 2220 9919 2239 nw
rect 9893 2193 9899 2220
tri 9899 2219 9900 2220 nw
rect 10391 2219 10443 2231
rect 5173 2192 6960 2193
tri 6960 2192 6961 2193 sw
tri 9551 2192 9552 2193 ne
rect 9552 2192 9617 2193
rect 5173 2186 7089 2192
tri 9552 2188 9556 2192 ne
rect 9556 2188 9617 2192
rect 5173 2173 6970 2186
rect 5055 2167 6970 2173
tri 6920 2152 6935 2167 ne
rect 6935 2152 6970 2167
rect 7004 2152 7042 2186
rect 7076 2152 7089 2186
tri 6935 2148 6939 2152 ne
rect 6939 2148 7089 2152
tri 6939 2146 6941 2148 ne
rect 6941 2146 7089 2148
tri 6941 2142 6945 2146 ne
rect 6945 2142 7089 2146
rect 7171 2182 9348 2188
rect 7171 2148 7218 2182
rect 7252 2148 7290 2182
rect 7324 2148 9230 2182
rect 9264 2148 9302 2182
rect 9336 2148 9348 2182
tri 9556 2171 9573 2188 ne
rect 9573 2171 9617 2188
tri 9617 2171 9639 2193 sw
tri 9573 2152 9592 2171 ne
rect 9592 2152 9639 2171
tri 9639 2152 9658 2171 sw
rect 9853 2152 9899 2193
tri 10526 2260 10567 2301 sw
rect 12473 2272 12525 2284
rect 10526 2254 11266 2260
rect 10526 2243 10620 2254
rect 10474 2231 10620 2243
rect 10526 2220 10620 2231
rect 10654 2220 10692 2254
rect 10726 2220 10764 2254
rect 10798 2220 10836 2254
rect 10870 2220 10908 2254
rect 10942 2220 10980 2254
rect 11014 2220 11052 2254
rect 11086 2220 11266 2254
rect 10526 2214 11266 2220
rect 11828 2214 11880 2260
rect 11881 2215 11882 2259
rect 11918 2215 11919 2259
rect 11920 2254 12414 2260
rect 11920 2220 12008 2254
rect 12042 2220 12080 2254
rect 12114 2220 12152 2254
rect 12186 2220 12224 2254
rect 12258 2220 12296 2254
rect 12330 2220 12368 2254
rect 12402 2220 12414 2254
rect 11920 2214 12414 2220
rect 10526 2179 10527 2214
rect 10474 2174 10527 2179
tri 10527 2174 10567 2214 nw
rect 10474 2173 10526 2174
tri 10526 2173 10527 2174 nw
rect 10391 2159 10443 2167
tri 9592 2150 9594 2152 ne
rect 9594 2150 9658 2152
tri 9658 2150 9660 2152 sw
tri 9594 2148 9596 2150 ne
rect 9596 2148 9660 2150
tri 9660 2148 9662 2150 sw
rect 7171 2142 9348 2148
tri 9596 2142 9602 2148 ne
rect 9602 2142 9663 2148
tri 6945 2140 6947 2142 ne
rect 6947 2140 7089 2142
tri 9602 2140 9604 2142 ne
rect 9604 2140 9663 2142
tri 9604 2136 9608 2140 ne
rect 9608 2136 9663 2140
tri 9608 2127 9617 2136 ne
rect 5012 2066 6634 2118
rect 6686 2066 6698 2118
rect 6750 2066 6756 2118
tri 6756 2112 6762 2118 sw
rect 7014 2066 7280 2112
rect 9617 2102 9623 2136
rect 9657 2102 9663 2136
rect 9617 2062 9663 2102
rect 9617 2028 9623 2062
rect 9657 2028 9663 2062
rect 5012 1940 6164 1992
rect 6216 1940 6243 1992
rect 6295 1940 6322 1992
rect 6374 1940 6401 1992
rect 6453 1940 7014 1992
rect 7280 1940 8946 1992
rect 8998 1940 9013 1992
rect 9065 1940 9080 1992
rect 9132 1940 9282 1992
rect 9617 1988 9663 2028
rect 9617 1954 9623 1988
rect 9657 1954 9663 1988
rect 9617 1914 9663 1954
tri 4960 1880 4988 1908 sw
rect 9617 1880 9623 1914
rect 9657 1880 9663 1914
rect 4914 1874 4988 1880
tri 4988 1874 4994 1880 sw
rect 4914 1872 9489 1874
tri 9489 1872 9491 1874 sw
rect 4914 1852 9491 1872
tri 9491 1852 9511 1872 sw
rect 4914 1845 9511 1852
tri 9511 1845 9518 1852 sw
tri 4378 1844 4379 1845 se
rect 4379 1844 4652 1845
tri 4652 1844 4653 1845 sw
rect 4914 1844 9518 1845
tri 9518 1844 9519 1845 sw
tri 4374 1840 4378 1844 se
rect 4378 1840 4653 1844
tri 4653 1840 4657 1844 sw
rect 4914 1840 9519 1844
tri 9519 1840 9523 1844 sw
rect 9617 1840 9663 1880
tri 4361 1827 4374 1840 se
rect 4374 1827 4657 1840
tri 4657 1827 4670 1840 sw
rect 4914 1828 9523 1840
tri 9523 1828 9535 1840 sw
tri 9469 1827 9470 1828 ne
rect 9470 1827 9535 1828
rect 4258 1817 4310 1823
tri 4351 1817 4361 1827 se
rect 4361 1817 4670 1827
tri 4340 1806 4351 1817 se
rect 4351 1806 4385 1817
tri 4385 1806 4396 1817 nw
tri 4622 1806 4633 1817 ne
rect 4633 1806 4670 1817
tri 4670 1806 4691 1827 sw
tri 9470 1806 9491 1827 ne
rect 9491 1806 9535 1827
tri 9535 1806 9557 1828 sw
rect 9617 1806 9623 1840
rect 9657 1806 9663 1840
tri 4336 1802 4340 1806 se
rect 4340 1802 4379 1806
tri 4334 1800 4336 1802 se
rect 4336 1800 4379 1802
tri 4379 1800 4385 1806 nw
tri 4633 1800 4639 1806 ne
rect 4639 1800 4691 1806
tri 4691 1800 4697 1806 sw
tri 9491 1800 9497 1806 ne
rect 9497 1800 9557 1806
tri 9557 1800 9563 1806 sw
tri 4333 1799 4334 1800 se
rect 4334 1799 4378 1800
tri 4378 1799 4379 1800 nw
tri 4639 1799 4640 1800 ne
rect 4640 1799 4697 1800
tri 4697 1799 4698 1800 sw
tri 9497 1799 9498 1800 ne
rect 9498 1799 9563 1800
tri 9563 1799 9564 1800 sw
tri 3122 1797 3124 1799 sw
tri 4331 1797 4333 1799 se
rect 4333 1797 4376 1799
tri 4376 1797 4378 1799 nw
tri 4640 1797 4642 1799 ne
rect 4642 1797 4698 1799
tri 4698 1797 4700 1799 sw
tri 9498 1797 9500 1799 ne
rect 9500 1797 9564 1799
rect 3122 1789 3124 1797
tri 3124 1789 3132 1797 sw
tri 4323 1789 4331 1797 se
rect 4331 1789 4368 1797
tri 4368 1789 4376 1797 nw
tri 4642 1789 4650 1797 ne
rect 4650 1789 4801 1797
tri 9500 1789 9508 1797 ne
rect 9508 1789 9564 1797
tri 9564 1789 9574 1799 sw
rect 3122 1777 3132 1789
tri 3132 1777 3144 1789 sw
tri 4311 1777 4323 1789 se
rect 4323 1777 4356 1789
tri 4356 1777 4368 1789 nw
rect 4418 1783 4470 1789
tri 4650 1788 4651 1789 ne
rect 4651 1788 4801 1789
tri 9508 1788 9509 1789 ne
rect 9509 1788 9574 1789
tri 9574 1788 9575 1789 sw
tri 4651 1787 4652 1788 ne
rect 4652 1787 4749 1788
rect 3122 1774 3144 1777
tri 3144 1774 3147 1777 sw
tri 4308 1774 4311 1777 se
rect 4311 1774 4353 1777
tri 4353 1774 4356 1777 nw
rect 3122 1766 4345 1774
tri 4345 1766 4353 1774 nw
rect 3122 1749 4322 1766
rect 3070 1743 4322 1749
tri 4322 1743 4345 1766 nw
tri 4410 1732 4418 1740 se
rect 2830 1712 2882 1718
tri 4393 1715 4410 1732 se
rect 4410 1731 4418 1732
tri 4652 1777 4662 1787 ne
rect 4662 1777 4749 1787
tri 4662 1769 4670 1777 ne
rect 4670 1769 4749 1777
tri 4715 1766 4718 1769 ne
rect 4718 1766 4749 1769
tri 4718 1738 4746 1766 ne
rect 4746 1738 4749 1766
tri 4746 1735 4749 1738 ne
tri 9509 1777 9520 1788 ne
rect 9520 1778 9575 1788
tri 9575 1778 9585 1788 sw
rect 9520 1777 9585 1778
tri 9520 1769 9528 1777 ne
rect 9528 1769 9585 1777
tri 9528 1766 9531 1769 ne
rect 9531 1766 9585 1769
tri 9531 1762 9535 1766 ne
rect 9535 1762 9585 1766
tri 9535 1758 9539 1762 ne
rect 6892 1738 6898 1752
rect 4410 1719 4470 1731
rect 4410 1715 4418 1719
tri 3099 1712 3102 1715 se
rect 3102 1712 4418 1715
tri 3096 1709 3099 1712 se
rect 3099 1709 4418 1712
tri 2527 1708 2528 1709 sw
tri 3095 1708 3096 1709 se
rect 3096 1708 4418 1709
rect 1792 1702 2528 1708
tri 2528 1702 2534 1708 sw
tri 3089 1702 3095 1708 se
rect 3095 1702 4418 1708
rect 1792 1692 2534 1702
tri 2534 1692 2544 1702 sw
tri 3079 1692 3089 1702 se
rect 3089 1692 4418 1702
rect 1792 1684 2544 1692
tri 2544 1684 2552 1692 sw
tri 3071 1684 3079 1692 se
rect 3079 1684 4418 1692
rect 1792 1667 4418 1684
rect 4749 1723 4801 1736
rect 1792 1661 4470 1667
rect 4637 1687 4689 1693
rect 1792 1648 3114 1661
tri 3114 1648 3127 1661 nw
rect 1792 1647 3113 1648
tri 3113 1647 3114 1648 nw
rect 1792 1630 3096 1647
tri 3096 1630 3113 1647 nw
rect 1792 1627 2549 1630
tri 2549 1627 2552 1630 nw
rect 1792 1618 2540 1627
tri 2540 1618 2549 1627 nw
rect 1792 1452 2527 1618
tri 2527 1605 2540 1618 nw
tri 3220 1605 3229 1614 se
rect 3229 1605 3300 1614
rect 4637 1609 4689 1635
rect 2882 1556 2965 1602
tri 2894 1538 2912 1556 ne
rect 2912 1538 2965 1556
tri 2912 1531 2919 1538 ne
tri 2823 1480 2830 1487 se
rect 2830 1481 2882 1487
tri 2811 1468 2823 1480 se
rect 2823 1468 2830 1480
rect 1792 1440 1805 1452
tri 1805 1440 1817 1452 nw
tri 2453 1440 2465 1452 ne
rect 2465 1440 2527 1452
rect 1792 1439 1804 1440
tri 1804 1439 1805 1440 nw
tri 2465 1439 2466 1440 ne
rect 2466 1439 2527 1440
tri 1792 1427 1804 1439 nw
tri 2466 1427 2478 1439 ne
rect 1663 1356 1709 1395
rect 1663 1322 1669 1356
rect 1703 1322 1709 1356
rect 1820 1355 2032 1407
rect 2084 1355 2096 1407
rect 2148 1355 2160 1407
rect 2212 1355 2224 1407
rect 2276 1355 2288 1407
rect 2340 1355 2403 1407
rect 1663 1283 1709 1322
rect 1663 1249 1669 1283
rect 1703 1249 1709 1283
rect 1663 1210 1709 1249
rect 1663 1176 1669 1210
rect 1703 1176 1709 1210
rect 1663 1137 1709 1176
rect 1663 1103 1669 1137
rect 1703 1103 1709 1137
rect 1663 1064 1709 1103
rect 1663 1030 1669 1064
rect 1703 1030 1709 1064
rect 1663 991 1709 1030
rect 1663 957 1669 991
rect 1703 957 1709 991
tri 1792 1330 1797 1335 sw
tri 2473 1330 2478 1335 se
rect 2478 1330 2527 1439
tri 2789 1446 2811 1468 se
rect 2811 1446 2830 1468
rect 2789 1429 2830 1446
rect 2789 1417 2882 1429
rect 2789 1400 2830 1417
tri 2789 1366 2823 1400 ne
rect 2823 1366 2830 1400
tri 2823 1364 2825 1366 ne
rect 2825 1365 2830 1366
rect 2825 1364 2882 1365
tri 2825 1359 2830 1364 ne
rect 2830 1359 2882 1364
rect 1792 1326 1797 1330
tri 1797 1326 1801 1330 sw
tri 2469 1326 2473 1330 se
rect 2473 1326 2527 1330
rect 1792 1320 1801 1326
tri 1801 1320 1807 1326 sw
tri 2463 1320 2469 1326 se
rect 2469 1320 2527 1326
rect 1792 1313 1807 1320
tri 1807 1313 1814 1320 sw
tri 2456 1313 2463 1320 se
rect 2463 1313 2527 1320
tri 2917 1313 2919 1315 se
rect 2919 1313 2965 1538
rect 3070 1596 3122 1602
rect 3070 1522 3122 1544
rect 3070 1449 3122 1470
rect 4637 1530 4689 1557
rect 4084 1414 4180 1460
tri 4100 1406 4108 1414 ne
rect 4108 1406 4180 1414
tri 4108 1400 4114 1406 ne
rect 4114 1400 4180 1406
rect 3070 1376 3122 1397
tri 4114 1380 4134 1400 ne
rect 4134 1366 4140 1400
rect 4174 1366 4180 1400
rect 4637 1451 4689 1478
rect 5012 1700 6898 1738
rect 6950 1700 6962 1752
rect 7014 1700 7020 1752
rect 7265 1700 7271 1752
rect 7323 1700 7335 1752
rect 7387 1700 9282 1752
rect 5012 1686 7020 1700
rect 5013 1684 7013 1685
rect 7014 1684 7020 1686
rect 4749 1658 4801 1671
rect 4749 1592 4801 1606
rect 5013 1647 7013 1648
rect 5012 1618 7014 1646
tri 9444 1627 9459 1642 se
rect 9459 1641 9511 1647
tri 9436 1619 9444 1627 se
rect 9444 1619 9459 1627
tri 7014 1618 7015 1619 sw
tri 9435 1618 9436 1619 se
rect 9436 1618 9459 1619
rect 5012 1615 7015 1618
tri 7015 1615 7018 1618 sw
tri 9432 1615 9435 1618 se
rect 9435 1615 9459 1618
rect 5012 1594 5043 1615
tri 5012 1584 5022 1594 ne
rect 5022 1584 5043 1594
tri 5022 1578 5028 1584 ne
rect 5028 1578 5043 1584
tri 5028 1572 5034 1578 ne
rect 5034 1572 5043 1578
tri 5034 1569 5037 1572 ne
rect 4749 1526 4801 1540
rect 5037 1563 5043 1572
rect 5095 1563 5113 1615
rect 5165 1563 5183 1615
rect 5235 1563 5253 1615
rect 5305 1572 5837 1615
rect 5305 1563 5337 1572
rect 5037 1551 5049 1563
rect 5083 1551 5121 1563
rect 5155 1551 5193 1563
rect 5227 1551 5265 1563
rect 5299 1551 5337 1563
rect 5037 1499 5043 1551
rect 5095 1499 5113 1551
rect 5165 1499 5183 1551
rect 5235 1499 5253 1551
rect 5305 1538 5337 1551
rect 5371 1538 5409 1572
rect 5443 1538 5481 1572
rect 5515 1538 5553 1572
rect 5587 1538 5625 1572
rect 5659 1538 5697 1572
rect 5731 1538 5769 1572
rect 5803 1563 5837 1572
rect 5889 1563 5903 1615
rect 5955 1563 5970 1615
rect 6022 1572 6142 1615
rect 6194 1572 6211 1615
rect 6263 1572 6281 1615
rect 6333 1572 6351 1615
rect 6403 1572 6421 1615
rect 6473 1589 9459 1615
rect 6473 1578 9511 1589
rect 6473 1572 7505 1578
rect 7557 1572 7578 1578
rect 7630 1572 7651 1578
rect 7703 1572 7724 1578
rect 7776 1572 7796 1578
rect 7848 1572 7868 1578
rect 7920 1572 7940 1578
rect 7992 1572 8012 1578
rect 8064 1572 8187 1578
rect 8239 1572 8289 1578
rect 8341 1572 8390 1578
rect 8442 1577 9511 1578
rect 8442 1572 8953 1577
rect 9005 1572 9080 1577
rect 9132 1575 9511 1577
rect 9132 1572 9459 1575
rect 6022 1563 6057 1572
rect 5803 1551 5841 1563
rect 5875 1551 5913 1563
rect 5947 1551 5985 1563
rect 6019 1551 6057 1563
rect 5803 1538 5837 1551
rect 5305 1499 5837 1538
rect 5889 1499 5903 1551
rect 5955 1499 5970 1551
rect 6022 1538 6057 1551
rect 6091 1538 6129 1572
rect 6194 1563 6201 1572
rect 6263 1563 6273 1572
rect 6333 1563 6345 1572
rect 6403 1563 6417 1572
rect 6473 1563 6489 1572
rect 6163 1551 6201 1563
rect 6235 1551 6273 1563
rect 6307 1551 6345 1563
rect 6379 1551 6417 1563
rect 6451 1551 6489 1563
rect 6194 1538 6201 1551
rect 6263 1538 6273 1551
rect 6333 1538 6345 1551
rect 6403 1538 6417 1551
rect 6473 1538 6489 1551
rect 6523 1538 6561 1572
rect 6595 1538 6633 1572
rect 6667 1538 6705 1572
rect 6739 1538 6777 1572
rect 6811 1538 6849 1572
rect 6883 1538 6921 1572
rect 6955 1538 6993 1572
rect 7027 1538 7065 1572
rect 7099 1538 7137 1572
rect 7171 1538 7209 1572
rect 7243 1538 7281 1572
rect 7315 1538 7353 1572
rect 7387 1538 7425 1572
rect 7459 1538 7497 1572
rect 7557 1538 7569 1572
rect 7630 1538 7641 1572
rect 7703 1538 7713 1572
rect 7776 1538 7785 1572
rect 7848 1538 7857 1572
rect 7920 1538 7929 1572
rect 7992 1538 8001 1572
rect 8064 1538 8073 1572
rect 8107 1538 8145 1572
rect 8179 1538 8187 1572
rect 8251 1538 8289 1572
rect 8341 1538 8361 1572
rect 8467 1538 8505 1572
rect 8539 1538 8577 1572
rect 8611 1538 8649 1572
rect 8683 1538 8721 1572
rect 8755 1538 8793 1572
rect 8827 1538 8865 1572
rect 8899 1538 8937 1572
rect 9005 1538 9010 1572
rect 9044 1538 9080 1572
rect 9132 1538 9156 1572
rect 9190 1538 9229 1572
rect 9263 1538 9302 1572
rect 9336 1538 9375 1572
rect 9409 1538 9459 1572
rect 6022 1499 6142 1538
rect 6194 1499 6211 1538
rect 6263 1499 6281 1538
rect 6333 1499 6351 1538
rect 6403 1499 6421 1538
rect 6473 1526 7505 1538
rect 7557 1526 7578 1538
rect 7630 1526 7651 1538
rect 7703 1526 7724 1538
rect 7776 1526 7796 1538
rect 7848 1526 7868 1538
rect 7920 1526 7940 1538
rect 7992 1526 8012 1538
rect 8064 1526 8187 1538
rect 8239 1526 8289 1538
rect 8341 1526 8390 1538
rect 8442 1526 8953 1538
rect 6473 1525 8953 1526
rect 9005 1525 9080 1538
rect 9132 1525 9459 1538
rect 6473 1523 9459 1525
rect 6473 1509 9511 1523
rect 6473 1499 9459 1509
tri 9428 1487 9440 1499 ne
rect 9440 1487 9459 1499
rect 4749 1468 4801 1474
tri 9440 1468 9459 1487 ne
rect 9459 1443 9511 1457
tri 3220 1340 3229 1349 ne
rect 3229 1340 3300 1349
rect 3070 1318 3122 1324
tri 2965 1313 2967 1315 sw
tri 3764 1313 3766 1315 se
rect 3766 1313 3812 1315
rect 1792 1310 1814 1313
tri 1814 1310 1817 1313 sw
tri 2453 1310 2456 1313 se
rect 2456 1310 2527 1313
rect 1792 996 2527 1310
tri 2894 1290 2917 1313 se
rect 2917 1308 2967 1313
tri 2967 1308 2972 1313 sw
tri 3759 1308 3764 1313 se
rect 3764 1308 3812 1313
rect 4134 1313 4180 1366
rect 2917 1290 2972 1308
tri 2972 1290 2990 1308 sw
tri 3741 1290 3759 1308 se
rect 3759 1290 3812 1308
rect 2608 1284 2854 1290
rect 2608 1250 2620 1284
rect 2654 1250 2692 1284
rect 2726 1250 2764 1284
rect 2798 1250 2854 1284
rect 2608 1244 2854 1250
rect 2855 1245 2856 1289
rect 2892 1245 2893 1289
rect 2894 1244 3812 1290
rect 3878 1256 3884 1308
rect 3936 1256 3948 1308
rect 4000 1256 4012 1308
rect 4064 1256 4084 1308
rect 4134 1279 4140 1313
rect 4174 1279 4180 1313
tri 3741 1225 3760 1244 ne
rect 3760 1225 3812 1244
tri 3760 1219 3766 1225 ne
rect 2830 1210 2882 1216
tri 2825 1170 2830 1175 se
tri 2792 1137 2825 1170 se
rect 2825 1158 2830 1170
rect 2825 1146 2882 1158
rect 2825 1137 2830 1146
tri 2789 1134 2792 1137 se
rect 2792 1134 2830 1137
rect 2830 1088 2882 1094
rect 3070 1210 3122 1216
tri 3228 1191 3230 1193 se
rect 3230 1191 3300 1193
tri 3220 1183 3228 1191 se
rect 3228 1183 3300 1191
rect 3070 1138 3122 1158
rect 1792 992 1813 996
tri 1813 992 1817 996 nw
tri 2453 992 2457 996 ne
rect 2457 992 2527 996
rect 1792 986 1807 992
tri 1807 986 1813 992 nw
tri 2457 986 2463 992 ne
rect 2463 986 2527 992
rect 1792 984 1805 986
tri 1805 984 1807 986 nw
tri 2463 984 2465 986 ne
rect 2465 984 2527 986
rect 1792 981 1802 984
tri 1802 981 1805 984 nw
tri 2465 981 2468 984 ne
rect 2468 981 2527 984
rect 3766 1172 3812 1225
rect 4134 1244 4180 1279
rect 4258 1370 4310 1376
rect 4258 1262 4310 1318
rect 4637 1372 4689 1399
tri 8529 1398 8554 1423 se
rect 8554 1417 8606 1423
tri 8525 1394 8529 1398 se
rect 8529 1394 8554 1398
tri 8524 1393 8525 1394 se
rect 8525 1393 8554 1394
tri 8606 1394 8635 1423 sw
rect 8606 1393 8635 1394
tri 8635 1393 8636 1394 sw
rect 8554 1353 8606 1365
tri 8520 1320 8551 1351 ne
rect 8551 1320 8554 1351
rect 4637 1314 4689 1320
tri 8551 1317 8554 1320 ne
rect 9459 1377 9511 1391
rect 8606 1320 8609 1351
tri 8609 1320 8640 1351 nw
rect 9459 1320 9468 1325
rect 9502 1320 9511 1325
tri 8606 1317 8609 1320 nw
rect 9459 1311 9511 1320
rect 8554 1295 8606 1301
tri 9261 1295 9268 1302 se
tri 9252 1286 9261 1295 se
rect 9261 1286 9268 1295
tri 9246 1280 9252 1286 se
rect 9252 1280 9268 1286
tri 9241 1275 9246 1280 se
rect 9246 1275 9268 1280
tri 4180 1244 4186 1250 sw
rect 4134 1225 4186 1244
rect 4134 1191 4140 1225
rect 4174 1216 4186 1225
tri 4186 1216 4214 1244 sw
rect 9459 1246 9468 1259
rect 9502 1246 9511 1259
rect 9459 1244 9511 1246
tri 9237 1216 9238 1217 ne
rect 9238 1216 9268 1217
rect 4174 1210 4230 1216
rect 4174 1191 4178 1210
tri 3812 1172 3822 1182 sw
tri 4124 1172 4134 1182 se
rect 4134 1172 4178 1191
rect 3766 1170 3822 1172
tri 3822 1170 3824 1172 sw
tri 4122 1170 4124 1172 se
rect 4124 1170 4178 1172
rect 3766 1148 3824 1170
tri 3824 1148 3846 1170 sw
tri 4100 1148 4122 1170 se
rect 4122 1158 4178 1170
tri 9238 1211 9243 1216 ne
rect 9243 1211 9268 1216
rect 4258 1204 4310 1210
tri 9243 1206 9248 1211 ne
rect 9248 1206 9268 1211
tri 9248 1204 9250 1206 ne
rect 9250 1204 9268 1206
tri 9250 1186 9268 1204 ne
rect 4122 1148 4230 1158
rect 3766 1146 4230 1148
rect 3766 1137 4178 1146
rect 3766 1103 4140 1137
rect 4174 1103 4178 1137
rect 3766 1094 4178 1103
rect 3766 1088 4230 1094
rect 9459 1177 9468 1192
rect 9502 1177 9511 1192
rect 9459 1110 9468 1125
rect 9502 1110 9511 1125
rect 3070 1067 3122 1086
rect 9459 1043 9468 1058
rect 9502 1043 9511 1058
rect 3070 996 3122 1015
rect 6830 1019 6964 1023
tri 1792 971 1802 981 nw
tri 2468 971 2478 981 ne
rect 1663 918 1709 957
rect 1663 884 1669 918
rect 1703 884 1709 918
rect 1820 899 2032 951
rect 2084 899 2096 951
rect 2148 899 2160 951
rect 2212 899 2224 951
rect 2276 899 2288 951
rect 2340 899 2424 951
rect 1663 845 1709 884
rect 1663 811 1669 845
rect 1703 811 1709 845
rect 1663 772 1709 811
rect 1663 738 1669 772
rect 1703 738 1709 772
rect 1663 699 1709 738
rect 1663 665 1669 699
rect 1703 665 1709 699
rect 1663 626 1709 665
rect 1663 592 1669 626
rect 1703 592 1709 626
rect 1663 553 1709 592
rect 1663 519 1669 553
rect 1703 519 1709 553
rect 1663 480 1709 519
tri 1792 876 1795 879 sw
tri 2475 876 2478 879 se
rect 2478 876 2527 981
rect 2566 929 2572 981
rect 2624 929 2636 981
rect 2688 929 2882 981
rect 3070 938 3122 944
rect 3878 940 3884 992
rect 3936 940 3948 992
rect 4000 940 4012 992
rect 4064 940 4084 992
rect 6830 967 6842 1019
rect 6894 967 6906 1019
rect 6958 967 6964 1019
rect 6830 965 6964 967
rect 9459 984 9511 991
rect 9459 976 9468 984
rect 9502 976 9511 984
rect 9459 910 9511 924
tri 2976 901 2985 910 se
rect 2985 901 4408 910
tri 4408 901 4417 910 sw
rect 9459 909 9468 910
rect 9502 909 9511 910
rect 1792 872 1795 876
tri 1795 872 1799 876 sw
tri 2471 872 2475 876 se
rect 2475 872 2527 876
rect 1792 870 1799 872
tri 1799 870 1801 872 sw
tri 2469 870 2471 872 se
rect 2471 870 2527 872
rect 1792 854 1801 870
tri 1801 854 1817 870 sw
tri 2453 854 2469 870 se
rect 2469 854 2527 870
rect 1792 540 2527 854
rect 2750 895 4417 901
rect 2802 843 2814 895
rect 2866 890 4417 895
tri 4417 890 4428 901 sw
rect 2866 876 4428 890
tri 4428 876 4442 890 sw
rect 2866 872 4442 876
tri 4442 872 4446 876 sw
rect 2866 870 4446 872
tri 4446 870 4448 872 sw
rect 2866 864 4448 870
rect 2750 837 2866 843
tri 2866 837 2893 864 nw
tri 4370 837 4397 864 ne
rect 4397 837 4448 864
tri 4448 837 4481 870 sw
rect 9459 842 9511 857
tri 4397 836 4398 837 ne
rect 4398 836 4481 837
tri 4481 836 4482 837 sw
rect 2940 828 3738 834
rect 2992 810 3738 828
tri 3738 810 3762 834 sw
rect 4084 830 4164 836
rect 2992 806 3762 810
tri 3762 806 3766 810 sw
rect 2992 802 3766 806
tri 3766 802 3770 806 sw
rect 2992 796 3770 802
tri 3770 796 3776 802 sw
rect 2992 795 3776 796
tri 3776 795 3777 796 sw
rect 2992 787 3777 795
tri 3777 787 3785 795 sw
rect 4084 790 4112 830
tri 4078 787 4081 790 ne
rect 4081 787 4112 790
rect 2992 780 3026 787
tri 3026 780 3033 787 nw
tri 3721 780 3728 787 ne
rect 3728 780 3785 787
tri 3785 780 3792 787 sw
tri 4081 780 4088 787 ne
rect 4088 780 4112 787
rect 2992 776 3009 780
rect 2940 764 3009 776
rect 2992 763 3009 764
tri 3009 763 3026 780 nw
tri 3728 763 3745 780 ne
rect 3745 763 3792 780
tri 3792 763 3809 780 sw
tri 4088 763 4105 780 ne
rect 4105 778 4112 780
tri 4398 806 4428 836 ne
rect 4428 806 4482 836
tri 4482 806 4512 836 sw
tri 4428 802 4432 806 ne
rect 4432 802 4512 806
tri 4432 796 4438 802 ne
rect 4438 796 4512 802
tri 4438 795 4439 796 ne
rect 4439 795 4512 796
tri 4439 780 4454 795 ne
rect 4105 763 4164 778
tri 2992 746 3009 763 nw
tri 3745 746 3762 763 ne
rect 3762 758 3809 763
tri 3809 758 3814 763 sw
rect 2940 706 2992 712
rect 1792 525 1802 540
tri 1802 525 1817 540 nw
tri 2453 525 2468 540 ne
rect 2468 525 2527 540
rect 3070 701 3122 707
rect 3070 628 3122 649
rect 3070 555 3122 576
rect 1792 517 1794 525
tri 1794 517 1802 525 nw
tri 2468 517 2476 525 ne
rect 2476 517 2527 525
tri 1792 515 1794 517 nw
tri 2476 515 2478 517 ne
rect 1663 446 1669 480
rect 1703 446 1709 480
rect 1663 407 1709 446
rect 1820 443 2032 495
rect 2084 443 2096 495
rect 2148 443 2160 495
rect 2212 443 2224 495
rect 2276 443 2288 495
rect 2340 443 2403 495
rect 2478 481 2527 517
rect 2566 473 2572 525
rect 2624 473 2636 525
rect 2688 473 2882 525
rect 3070 482 3122 503
rect 3762 495 3814 758
tri 4105 756 4112 763 ne
rect 4112 756 4164 763
rect 4112 682 4164 704
rect 3878 630 3884 682
rect 3936 630 3948 682
rect 4000 630 4012 682
rect 4064 630 4084 682
rect 4112 609 4164 630
tri 4098 544 4112 558 se
rect 4112 544 4164 557
tri 4094 540 4098 544 se
rect 4098 540 4164 544
tri 4078 524 4094 540 se
rect 4094 536 4164 540
rect 4094 524 4112 536
tri 3814 495 3823 504 sw
rect 3762 489 3823 495
tri 3823 489 3829 495 sw
rect 3762 486 3829 489
tri 3829 486 3832 489 sw
rect 3762 482 3832 486
tri 3832 482 3836 486 sw
rect 4084 484 4112 524
tri 3762 471 3773 482 ne
rect 3773 471 3836 482
tri 3836 471 3847 482 sw
rect 4084 478 4164 484
rect 4258 698 4310 704
rect 4454 690 4512 795
rect 9459 775 9511 790
rect 9459 708 9511 723
tri 4512 690 4517 695 sw
rect 4454 682 4517 690
tri 4517 682 4525 690 sw
rect 4454 671 4525 682
tri 4525 671 4536 682 sw
tri 4454 656 4469 671 ne
rect 4469 656 4536 671
tri 4536 656 4551 671 sw
rect 4258 624 4310 646
tri 4469 643 4482 656 ne
rect 4482 643 4551 656
tri 4551 643 4564 656 sw
tri 4482 630 4495 643 ne
rect 4495 630 4564 643
tri 4564 630 4577 643 sw
rect 9459 641 9511 656
tri 4495 617 4508 630 ne
rect 4508 617 4577 630
tri 4577 617 4590 630 sw
tri 4508 589 4536 617 ne
rect 4536 589 4590 617
tri 4590 589 4618 617 sw
tri 4536 583 4542 589 ne
rect 4542 583 4870 589
tri 4870 583 4876 589 sw
rect 9459 583 9468 589
rect 9502 583 9511 589
rect 4258 550 4310 572
tri 4542 570 4555 583 ne
rect 4555 570 4876 583
tri 4876 570 4889 583 sw
rect 9459 574 9511 583
tri 4555 569 4556 570 ne
rect 4556 569 4889 570
tri 4889 569 4890 570 sw
tri 4556 544 4581 569 ne
rect 4581 544 4890 569
tri 4890 544 4915 569 sw
tri 4581 531 4594 544 ne
rect 4594 531 4915 544
tri 4846 519 4858 531 ne
rect 4858 519 4915 531
tri 4915 519 4940 544 sw
tri 4858 510 4867 519 ne
rect 4867 510 4980 519
tri 4867 507 4870 510 ne
rect 4870 507 4980 510
rect 4258 477 4310 498
tri 4870 495 4882 507 ne
rect 4882 495 4980 507
tri 4882 489 4888 495 ne
rect 4888 489 4980 495
tri 3773 470 3774 471 ne
rect 3774 470 3847 471
tri 3847 470 3848 471 sw
tri 3774 465 3779 470 ne
rect 3779 465 3848 470
tri 3848 465 3853 470 sw
tri 4888 471 4906 489 ne
rect 4906 471 4980 489
tri 4906 470 4907 471 ne
rect 4907 470 4980 471
tri 4907 469 4908 470 ne
rect 4908 469 4980 470
tri 3779 464 3780 465 ne
rect 3780 464 3853 465
tri 3853 464 3854 465 sw
tri 3780 461 3783 464 ne
rect 3783 461 3854 464
tri 3854 461 3857 464 sw
tri 3783 449 3795 461 ne
rect 3795 450 3857 461
tri 3857 450 3868 461 sw
rect 3795 449 4184 450
tri 4184 449 4185 450 sw
rect 1663 373 1669 407
rect 1703 402 1709 407
tri 3795 431 3813 449 ne
rect 3813 447 4185 449
tri 4185 447 4187 449 sw
rect 3813 431 4187 447
tri 4187 431 4203 447 sw
tri 1709 402 1710 403 sw
tri 3069 402 3070 403 se
rect 3070 402 3122 430
tri 3813 414 3830 431 ne
rect 3830 414 4203 431
tri 4203 414 4220 431 sw
rect 4258 419 4310 425
rect 4637 463 4689 469
tri 4908 464 4913 469 ne
rect 4913 464 4980 469
tri 4913 461 4916 464 ne
rect 4916 461 4980 464
rect 9459 510 9468 522
rect 9502 510 9511 522
rect 9459 507 9511 510
rect 9539 548 9585 1762
rect 9617 1766 9663 1806
rect 9617 1732 9623 1766
rect 9657 1732 9663 1766
rect 9617 1692 9663 1732
rect 9617 1658 9623 1692
rect 9657 1658 9663 1692
rect 9617 1618 9663 1658
rect 9617 1584 9623 1618
rect 9657 1584 9663 1618
rect 9617 1544 9663 1584
rect 9617 1510 9623 1544
rect 9657 1510 9663 1544
rect 9617 1470 9663 1510
rect 9617 1436 9623 1470
rect 9657 1436 9663 1470
rect 9617 1395 9663 1436
rect 9617 1361 9623 1395
rect 9657 1361 9663 1395
rect 9617 1320 9663 1361
rect 9617 1286 9623 1320
rect 9657 1286 9663 1320
rect 9617 1245 9663 1286
rect 9617 1211 9623 1245
rect 9657 1211 9663 1245
rect 9617 1170 9663 1211
rect 9617 1136 9623 1170
rect 9657 1136 9663 1170
rect 9617 1095 9663 1136
rect 9617 1061 9623 1095
rect 9657 1061 9663 1095
rect 9617 1020 9663 1061
rect 9617 986 9623 1020
rect 9657 986 9663 1020
rect 9617 945 9663 986
rect 9617 911 9623 945
rect 9657 911 9663 945
rect 9617 870 9663 911
rect 9617 836 9623 870
rect 9657 836 9663 870
rect 9853 2118 9859 2152
rect 9893 2118 9899 2152
tri 12457 2142 12473 2158 se
rect 12473 2142 12525 2220
tri 12455 2140 12457 2142 se
rect 12457 2140 12525 2142
tri 12454 2139 12455 2140 se
rect 12455 2139 12525 2140
tri 12448 2133 12454 2139 se
rect 12454 2133 12525 2139
rect 9853 2077 9899 2118
tri 10483 2111 10505 2133 se
rect 10505 2111 12525 2133
tri 10471 2099 10483 2111 se
rect 10483 2099 12525 2111
rect 9853 2043 9859 2077
rect 9893 2043 9899 2077
tri 10447 2075 10471 2099 se
rect 10471 2087 12525 2099
rect 12661 2254 12715 2261
rect 12713 2202 12715 2254
rect 12661 2190 12715 2202
rect 12713 2138 12715 2190
rect 12661 2126 12715 2138
rect 10471 2075 10505 2087
rect 9853 2002 9899 2043
rect 9853 1968 9859 2002
rect 9893 1968 9899 2002
rect 9853 1927 9899 1968
rect 9853 1893 9859 1927
rect 9893 1893 9899 1927
rect 9853 1852 9899 1893
rect 9853 1818 9859 1852
rect 9893 1818 9899 1852
rect 9853 1777 9899 1818
rect 9853 1743 9859 1777
rect 9893 1743 9899 1777
rect 9853 1702 9899 1743
rect 9853 1668 9859 1702
rect 9893 1668 9899 1702
rect 9853 1627 9899 1668
rect 9853 1593 9859 1627
rect 9893 1593 9899 1627
rect 9853 1552 9899 1593
rect 9853 1518 9859 1552
rect 9893 1518 9899 1552
rect 9853 1477 9899 1518
rect 9853 1443 9859 1477
rect 9893 1443 9899 1477
rect 9853 1402 9899 1443
rect 10089 2063 10135 2075
tri 10439 2067 10447 2075 se
rect 10447 2067 10505 2075
tri 10505 2067 10525 2087 nw
rect 12713 2074 12715 2126
tri 10437 2065 10439 2067 se
rect 10439 2065 10503 2067
tri 10503 2065 10505 2067 nw
rect 12661 2065 12675 2074
rect 12709 2065 12715 2074
rect 10089 2029 10095 2063
rect 10129 2029 10135 2063
rect 10089 1989 10135 2029
tri 10396 2024 10437 2065 se
rect 10437 2024 10462 2065
tri 10462 2024 10503 2065 nw
rect 12661 2062 12715 2065
tri 10385 2013 10396 2024 se
rect 10396 2013 10451 2024
tri 10451 2013 10462 2024 nw
tri 10343 1992 10364 2013 se
rect 10364 1992 10428 2013
tri 10341 1990 10343 1992 se
rect 10343 1990 10428 1992
tri 10428 1990 10451 2013 nw
rect 12713 2010 12715 2062
rect 10536 2007 12558 2008
rect 10089 1955 10095 1989
rect 10129 1955 10135 1989
tri 10322 1971 10341 1990 se
rect 10341 1983 10421 1990
tri 10421 1983 10428 1990 nw
rect 10341 1972 10410 1983
tri 10410 1972 10421 1983 nw
rect 10341 1971 10409 1972
tri 10409 1971 10410 1972 nw
rect 10089 1915 10135 1955
tri 10300 1949 10322 1971 se
rect 10322 1949 10366 1971
tri 10366 1949 10388 1971 nw
rect 10536 1955 10588 2007
rect 10640 1955 10657 2007
rect 10709 1955 10727 2007
rect 10779 1955 10797 2007
rect 10849 1955 10867 2007
rect 10919 1955 10937 2007
rect 10989 1955 11007 2007
rect 11059 1955 11207 2007
rect 11259 1955 11274 2007
rect 11326 1955 11341 2007
rect 11393 1955 11600 2007
rect 11652 1955 11668 2007
rect 11720 1955 11737 2007
rect 11789 1955 12399 2007
rect 12451 1955 12467 2007
rect 12519 1955 12558 2007
rect 12661 1998 12675 2010
rect 12709 1998 12715 2010
tri 10291 1940 10300 1949 se
rect 10300 1940 10357 1949
tri 10357 1940 10366 1949 nw
rect 12713 1946 12715 1998
rect 10089 1881 10095 1915
rect 10129 1881 10135 1915
rect 10089 1841 10135 1881
rect 10089 1807 10095 1841
rect 10129 1807 10135 1841
rect 10089 1767 10135 1807
rect 10089 1733 10095 1767
rect 10129 1733 10135 1767
rect 10089 1693 10135 1733
rect 10089 1659 10095 1693
rect 10129 1659 10135 1693
rect 10089 1619 10135 1659
rect 10089 1585 10095 1619
rect 10129 1585 10135 1619
rect 10089 1545 10135 1585
rect 10089 1511 10095 1545
rect 10129 1511 10135 1545
rect 10089 1470 10135 1511
rect 10089 1436 10095 1470
rect 10129 1436 10135 1470
rect 9853 1368 9859 1402
rect 9893 1368 9899 1402
rect 9853 1327 9899 1368
rect 9853 1293 9859 1327
rect 9893 1293 9899 1327
rect 9853 1252 9899 1293
rect 9853 1218 9859 1252
rect 9893 1218 9899 1252
rect 9853 1176 9899 1218
rect 9853 1142 9859 1176
rect 9893 1142 9899 1176
rect 9853 1100 9899 1142
rect 9853 1066 9859 1100
rect 9893 1066 9899 1100
rect 9853 1024 9899 1066
rect 9853 990 9859 1024
rect 9893 990 9899 1024
rect 9853 948 9899 990
rect 9853 914 9859 948
rect 9893 914 9899 948
rect 9853 872 9899 914
rect 9617 795 9663 836
rect 9617 761 9623 795
rect 9657 761 9663 795
rect 9617 720 9663 761
rect 9617 686 9623 720
rect 9657 686 9663 720
rect 9617 674 9663 686
rect 9732 834 9784 840
rect 9732 770 9784 782
tri 9728 643 9732 647 se
rect 9732 643 9784 718
rect 9853 838 9859 872
rect 9893 838 9899 872
rect 9853 796 9899 838
rect 9853 762 9859 796
rect 9893 762 9899 796
rect 9853 720 9899 762
rect 9853 686 9859 720
rect 9893 686 9899 720
rect 9853 674 9899 686
rect 10008 1399 10060 1405
rect 10008 1335 10060 1347
tri 10007 647 10008 648 se
rect 10008 647 10060 1283
rect 10089 1395 10135 1436
rect 10089 1361 10095 1395
rect 10129 1361 10135 1395
rect 10089 1320 10135 1361
rect 10089 1286 10095 1320
rect 10129 1286 10135 1320
rect 10089 1245 10135 1286
rect 10089 1211 10095 1245
rect 10129 1211 10135 1245
rect 10089 1170 10135 1211
rect 10089 1136 10095 1170
rect 10129 1136 10135 1170
rect 10089 1095 10135 1136
rect 10089 1061 10095 1095
rect 10129 1061 10135 1095
rect 10089 1020 10135 1061
rect 10089 986 10095 1020
rect 10129 986 10135 1020
rect 10089 945 10135 986
rect 10089 911 10095 945
rect 10129 911 10135 945
rect 10089 870 10135 911
rect 10089 836 10095 870
rect 10129 836 10135 870
rect 10089 802 10135 836
tri 10276 1925 10291 1940 se
rect 10291 1925 10335 1940
rect 10276 1918 10335 1925
tri 10335 1918 10357 1940 nw
rect 12661 1934 12675 1946
rect 12709 1934 12715 1946
rect 10276 1917 10334 1918
tri 10334 1917 10335 1918 nw
rect 10276 1915 10332 1917
tri 10332 1915 10334 1917 nw
rect 10276 1906 10323 1915
tri 10323 1906 10332 1915 nw
rect 10391 1911 11173 1918
tri 10135 802 10141 808 sw
rect 10089 796 10141 802
rect 10089 732 10141 744
rect 10089 674 10141 680
tri 9784 643 9788 647 sw
tri 10003 643 10007 647 se
rect 10007 643 10060 647
tri 9699 614 9728 643 se
rect 9728 614 9788 643
tri 9788 614 9817 643 sw
tri 9974 614 10003 643 se
rect 10003 614 10060 643
tri 9698 613 9699 614 se
rect 9699 613 9817 614
tri 9817 613 9818 614 sw
rect 9694 604 9824 613
rect 9694 570 9706 604
rect 9740 570 9778 604
rect 9812 570 9824 604
rect 9694 561 9824 570
rect 9930 605 10060 614
rect 9930 571 9942 605
rect 9976 571 10014 605
rect 10048 571 10060 605
rect 9930 562 10060 571
tri 9585 548 9593 556 sw
rect 9539 536 9593 548
tri 9593 536 9605 548 sw
tri 10264 536 10276 548 se
rect 10276 536 10322 1906
tri 10322 1905 10323 1906 nw
rect 10443 1859 11121 1911
rect 10391 1847 11173 1859
rect 10443 1826 11121 1847
tri 10443 1801 10468 1826 nw
tri 10532 1801 10557 1826 ne
rect 10557 1801 11121 1826
tri 10557 1800 10558 1801 ne
rect 10558 1800 11121 1801
tri 10558 1799 10559 1800 ne
rect 10559 1799 11121 1800
rect 10391 1788 10443 1795
tri 10559 1789 10569 1799 ne
rect 10569 1795 11121 1799
rect 10569 1789 11173 1795
rect 10474 1788 10526 1789
tri 10526 1788 10527 1789 sw
tri 10569 1788 10570 1789 ne
rect 10570 1788 11173 1789
rect 11996 1912 12633 1918
rect 11996 1860 12307 1912
rect 12359 1906 12633 1912
rect 12359 1872 12590 1906
rect 12624 1872 12633 1906
rect 12359 1860 12633 1872
rect 11996 1834 12633 1860
rect 11996 1833 12590 1834
rect 10474 1783 10527 1788
rect 10526 1765 10527 1783
tri 10527 1765 10550 1788 sw
rect 11996 1781 12307 1833
rect 12359 1800 12590 1833
rect 12624 1800 12633 1834
rect 12359 1781 12633 1800
rect 10526 1748 10550 1765
tri 10550 1748 10567 1765 sw
rect 11996 1753 12633 1781
rect 10526 1742 11098 1748
rect 10526 1731 10620 1742
rect 10474 1719 10620 1731
rect 10526 1708 10620 1719
rect 10654 1708 10692 1742
rect 10726 1708 10764 1742
rect 10798 1708 10836 1742
rect 10870 1708 10908 1742
rect 10942 1708 10980 1742
rect 11014 1708 11052 1742
rect 11086 1708 11098 1742
rect 10526 1702 11098 1708
rect 10526 1690 10555 1702
tri 10555 1690 10567 1702 nw
rect 11996 1701 12307 1753
rect 12359 1701 12633 1753
rect 10526 1667 10527 1690
rect 10474 1662 10527 1667
tri 10527 1662 10555 1690 nw
rect 11996 1673 12633 1701
rect 10391 1655 10443 1662
rect 10474 1661 10526 1662
tri 10526 1661 10527 1662 nw
tri 10569 1661 10570 1662 se
rect 10570 1661 11173 1662
tri 10558 1650 10569 1661 se
rect 10569 1655 11173 1661
rect 10569 1650 11121 1655
tri 10557 1649 10558 1650 se
rect 10558 1649 11121 1650
tri 10443 1624 10468 1649 sw
tri 10532 1624 10557 1649 se
rect 10557 1624 11121 1649
rect 10443 1603 11121 1624
rect 10391 1591 11173 1603
rect 10443 1539 11121 1591
rect 10391 1532 11173 1539
rect 11996 1621 12307 1673
rect 12359 1650 12633 1673
rect 12359 1621 12590 1650
rect 11996 1616 12590 1621
rect 12624 1616 12633 1650
rect 11996 1593 12633 1616
rect 11996 1541 12307 1593
rect 12359 1578 12633 1593
rect 12359 1544 12590 1578
rect 12624 1544 12633 1578
rect 12359 1541 12633 1544
rect 11996 1532 12633 1541
rect 12713 1882 12715 1934
rect 12661 1874 12715 1882
rect 12661 1870 12675 1874
rect 12709 1870 12715 1874
rect 12713 1818 12715 1870
rect 12661 1806 12715 1818
rect 12713 1754 12715 1806
rect 12661 1742 12715 1754
rect 12713 1690 12715 1742
rect 12661 1678 12715 1690
rect 12713 1626 12715 1678
rect 12661 1615 12675 1626
rect 12709 1615 12715 1626
rect 12661 1614 12715 1615
rect 12713 1562 12715 1614
rect 12661 1550 12675 1562
rect 12709 1550 12715 1562
rect 12713 1498 12715 1550
rect 10536 1495 12558 1496
rect 10536 1443 10588 1495
rect 10640 1443 10657 1495
rect 10709 1443 10727 1495
rect 10779 1443 10797 1495
rect 10849 1443 10867 1495
rect 10919 1443 10937 1495
rect 10989 1443 11007 1495
rect 11059 1443 12399 1495
rect 12451 1443 12467 1495
rect 12519 1443 12558 1495
rect 12661 1486 12675 1498
rect 12709 1486 12715 1498
rect 12713 1434 12715 1486
rect 12661 1424 12715 1434
rect 12661 1422 12675 1424
rect 12709 1422 12715 1424
rect 10416 1381 12605 1387
rect 10468 1329 11121 1381
rect 11173 1329 11851 1381
rect 11903 1329 12553 1381
rect 10416 1311 12605 1329
rect 10468 1259 11121 1311
rect 11173 1259 11851 1311
rect 11903 1259 12553 1311
rect 10416 1241 12605 1259
rect 10468 1189 11121 1241
rect 11173 1189 11851 1241
rect 11903 1189 12553 1241
rect 10416 1181 10423 1189
rect 10457 1181 11130 1189
rect 11164 1181 11860 1189
rect 11894 1181 12565 1189
rect 12599 1181 12605 1189
rect 10416 1171 12605 1181
rect 10468 1119 11121 1171
rect 11173 1119 11851 1171
rect 11903 1119 12553 1171
rect 10416 1102 10423 1119
rect 10457 1102 11130 1119
rect 11164 1102 11860 1119
rect 11894 1102 12565 1119
rect 12599 1102 12605 1119
rect 10416 1101 12605 1102
rect 10468 1049 11121 1101
rect 11173 1049 11851 1101
rect 11903 1049 12553 1101
rect 10416 1031 10423 1049
rect 10457 1031 11130 1049
rect 11164 1031 11860 1049
rect 11894 1031 12565 1049
rect 12599 1031 12605 1049
rect 10468 979 11121 1031
rect 11173 979 11851 1031
rect 11903 979 12553 1031
rect 10416 978 12605 979
rect 10416 961 10423 978
rect 10457 961 11130 978
rect 11164 961 11860 978
rect 11894 961 12565 978
rect 12599 961 12605 978
rect 10468 909 11121 961
rect 11173 909 11851 961
rect 11903 909 12553 961
rect 10416 899 12605 909
rect 10416 891 10423 899
rect 10457 891 11130 899
rect 11164 891 11860 899
rect 11894 891 12565 899
rect 12599 891 12605 899
rect 10468 839 11121 891
rect 11173 839 11851 891
rect 11903 839 12553 891
rect 10416 822 12605 839
rect 10468 770 11121 822
rect 11173 770 11851 822
rect 11903 770 12553 822
rect 10416 753 12605 770
rect 10468 701 11121 753
rect 11173 701 11851 753
rect 11903 701 12553 753
rect 10416 695 12605 701
rect 12713 1370 12715 1422
rect 12661 1357 12715 1370
rect 12713 1305 12715 1357
rect 12661 1292 12715 1305
rect 12713 1240 12715 1292
rect 12661 1227 12715 1240
rect 12713 1175 12715 1227
rect 12661 1165 12675 1175
rect 12709 1165 12715 1175
rect 12661 1162 12715 1165
rect 12713 1110 12715 1162
rect 12661 1097 12675 1110
rect 12709 1097 12715 1110
rect 12713 1045 12715 1097
rect 12661 1032 12675 1045
rect 12709 1032 12715 1045
rect 12713 980 12715 1032
rect 12661 974 12715 980
rect 12661 967 12675 974
rect 12709 967 12715 974
rect 12713 915 12715 967
rect 12661 902 12715 915
rect 12713 850 12715 902
rect 12661 837 12715 850
rect 12713 785 12715 837
rect 12661 772 12715 785
rect 12713 720 12715 772
rect 12661 717 12675 720
rect 12709 717 12715 720
rect 12661 707 12715 717
rect 12713 655 12715 707
rect 12661 643 12675 655
rect 12709 643 12715 655
rect 12661 642 12715 643
rect 10499 587 10505 639
rect 10557 587 10576 639
rect 10628 587 10647 639
rect 10699 587 10719 639
rect 10771 587 10791 639
rect 10843 587 10863 639
rect 10915 587 10935 639
rect 10987 587 11007 639
rect 11059 587 11965 639
rect 12017 587 12029 639
rect 12081 587 12093 639
rect 12145 587 12157 639
rect 12209 587 12221 639
rect 12273 587 12399 639
rect 12451 587 12500 639
rect 12552 587 12558 639
rect 12713 590 12715 642
tri 9539 495 9580 536 ne
rect 9580 528 9605 536
tri 9605 528 9613 536 sw
tri 10256 528 10264 536 se
rect 10264 528 10322 536
rect 9580 510 9613 528
tri 9613 510 9631 528 sw
tri 10238 510 10256 528 se
rect 10256 510 10289 528
rect 9580 495 10289 510
tri 10289 495 10322 528 nw
rect 12661 569 12675 590
rect 12709 569 12715 590
tri 12636 498 12661 523 se
rect 12661 498 12715 569
tri 9580 489 9586 495 ne
rect 9586 489 10283 495
tri 10283 489 10289 495 nw
tri 9586 470 9605 489 ne
rect 9605 470 10264 489
tri 10264 470 10283 489 nw
tri 9605 464 9611 470 ne
rect 9611 464 10258 470
tri 10258 464 10264 470 nw
tri 3830 412 3832 414 ne
rect 3832 412 4220 414
tri 4220 412 4222 414 sw
tri 4158 409 4161 412 ne
rect 4161 409 4222 412
rect 1703 398 1710 402
tri 1710 398 1714 402 sw
tri 3065 398 3069 402 se
rect 3069 398 3122 402
rect 1703 378 1714 398
tri 1714 378 1734 398 sw
tri 3045 378 3065 398 se
rect 3065 383 3122 398
tri 3706 402 3713 409 sw
tri 4161 402 4168 409 ne
rect 4168 402 4222 409
tri 4222 402 4232 412 sw
rect 3706 398 3713 402
tri 3713 398 3717 402 sw
tri 4168 398 4172 402 ne
rect 4172 398 4232 402
tri 4232 398 4236 402 sw
rect 3706 392 3717 398
tri 3717 392 3723 398 sw
tri 4172 392 4178 398 ne
rect 4178 395 4236 398
tri 4236 395 4239 398 sw
rect 4178 392 4239 395
tri 3122 383 3131 392 sw
rect 3706 383 3723 392
tri 3723 383 3732 392 sw
tri 4178 383 4187 392 ne
rect 3065 378 3131 383
rect 1703 373 2032 378
rect 1663 369 2032 373
rect 2084 369 2096 378
rect 2148 369 2160 378
rect 1663 335 1783 369
rect 1817 335 1857 369
rect 1891 335 1931 369
rect 1965 335 2005 369
rect 2148 335 2153 369
rect 1663 326 2032 335
rect 2084 326 2096 335
rect 2148 326 2160 335
rect 2212 326 2224 378
rect 2276 326 2288 378
rect 2340 369 2380 378
rect 2340 335 2375 369
rect 2340 326 2380 335
rect 2432 326 2444 378
rect 2496 326 2508 378
rect 2560 326 2572 378
rect 2624 369 2636 378
rect 2688 369 2700 378
rect 2752 369 2769 378
rect 2821 369 2838 378
rect 2890 369 2907 378
rect 2959 369 2977 378
rect 3029 369 3047 378
rect 3099 377 3131 378
tri 3131 377 3137 383 sw
rect 3706 377 4144 383
rect 3099 375 3137 377
tri 3137 375 3139 377 sw
rect 2631 335 2636 369
rect 2890 335 2893 369
rect 2959 335 2967 369
rect 3029 335 3041 369
rect 3099 343 3139 375
tri 3139 343 3171 375 sw
tri 3220 343 3248 371 ne
rect 3248 343 3300 371
rect 3099 337 3171 343
tri 3171 337 3177 343 sw
tri 3248 337 3254 343 ne
rect 3254 337 3300 343
rect 3706 343 3738 377
rect 3772 343 3810 377
rect 3844 343 3882 377
rect 3916 343 3954 377
rect 3988 343 4026 377
rect 4060 343 4098 377
rect 4132 343 4144 377
rect 3706 337 4144 343
rect 2624 326 2636 335
rect 2688 326 2700 335
rect 2752 326 2769 335
rect 2821 326 2838 335
rect 2890 326 2907 335
rect 2959 326 2977 335
rect 3029 326 3047 335
rect 3099 330 3177 337
tri 3177 330 3184 337 sw
rect 3099 326 3184 330
tri 3184 326 3188 330 sw
tri 3131 318 3139 326 ne
rect 3139 318 3188 326
tri 3188 318 3196 326 sw
tri 3139 296 3161 318 ne
rect 3161 315 3196 318
tri 3196 315 3199 318 sw
rect 3161 296 3199 315
tri 3199 296 3218 315 sw
tri 3161 294 3163 296 ne
rect 3163 294 3218 296
tri 3218 294 3220 296 sw
tri 3163 291 3166 294 ne
rect 3166 291 3220 294
tri 3220 291 3223 294 sw
tri 3166 281 3176 291 ne
rect 3176 281 3223 291
tri 3223 281 3233 291 sw
tri 3176 261 3196 281 ne
rect 3196 272 3233 281
tri 3233 272 3242 281 sw
rect 3196 261 3242 272
tri 3242 261 3253 272 sw
tri 3196 247 3210 261 ne
rect 3210 247 3926 261
tri 3926 247 3940 261 sw
tri 3210 245 3212 247 ne
rect 3212 245 3940 247
tri 3940 245 3942 247 sw
tri 3212 227 3230 245 ne
rect 3230 227 3942 245
tri 3942 227 3960 245 sw
tri 3230 218 3239 227 ne
rect 3239 218 3960 227
tri 3891 211 3898 218 ne
rect 3898 211 3960 218
tri 3960 211 3976 227 sw
tri 3898 208 3901 211 ne
rect 3901 208 3976 211
tri 3976 208 3979 211 sw
tri 3901 149 3960 208 ne
rect 3960 205 3979 208
tri 3979 205 3982 208 sw
rect 3960 169 3982 205
tri 3982 169 4018 205 sw
rect 4187 177 4239 392
rect 4637 351 4689 411
rect 4637 296 4646 299
rect 4680 296 4689 299
rect 4637 281 4689 296
rect 4829 436 4881 448
rect 4829 411 4835 436
rect 4869 411 4881 436
rect 4829 328 4881 359
rect 4829 309 4835 328
rect 4869 309 4881 328
rect 9459 440 9468 455
rect 9502 440 9511 455
rect 10493 446 10501 498
rect 10553 446 10573 498
rect 10625 446 10645 498
rect 10697 446 10717 498
rect 10769 446 10789 498
rect 10841 446 10861 498
rect 10913 446 10934 498
rect 10986 446 11007 498
rect 11059 446 11207 498
rect 11259 446 11273 498
rect 11325 446 11339 498
rect 11391 489 11405 498
rect 11457 489 11471 498
rect 11523 489 11537 498
rect 11589 489 11603 498
rect 11655 489 11670 498
rect 11396 455 11405 489
rect 11655 455 11662 489
rect 11391 446 11405 455
rect 11457 446 11471 455
rect 11523 446 11537 455
rect 11589 446 11603 455
rect 11655 446 11670 455
rect 11722 446 11737 498
rect 11789 489 11965 498
rect 11789 455 11812 489
rect 11846 455 11887 489
rect 11921 455 11962 489
rect 11789 446 11965 455
rect 12017 446 12029 498
rect 12081 446 12093 498
rect 12145 489 12157 498
rect 12209 489 12221 498
rect 12273 489 12399 498
rect 12451 489 12500 498
rect 12552 489 12715 498
rect 12146 455 12157 489
rect 12296 455 12337 489
rect 12371 455 12399 489
rect 12451 455 12487 489
rect 12552 455 12562 489
rect 12596 455 12637 489
rect 12671 455 12715 489
rect 12145 446 12157 455
rect 12209 446 12221 455
rect 12273 446 12399 455
rect 12451 446 12500 455
rect 12552 446 12715 455
rect 9459 373 9468 388
rect 9502 373 9511 388
rect 9459 291 9468 321
rect 9502 291 9511 321
tri 4881 281 4887 287 sw
tri 4992 281 4998 287 se
rect 4881 272 4887 281
tri 4887 272 4896 281 sw
tri 4983 272 4992 281 se
rect 4992 272 4998 281
rect 4881 257 4896 272
rect 4829 253 4896 257
tri 4896 253 4915 272 sw
tri 4964 253 4983 272 se
rect 4983 253 4998 272
tri 5116 281 5122 287 sw
tri 9204 281 9210 287 se
rect 5116 272 5122 281
tri 5122 272 5131 281 sw
tri 9195 272 9204 281 se
rect 9204 272 9210 281
rect 5116 253 5131 272
tri 5131 253 5150 272 sw
tri 9176 253 9195 272 se
rect 9195 253 9210 272
tri 9328 281 9334 287 sw
tri 9453 281 9459 287 se
rect 9459 281 9511 291
rect 11294 314 11340 326
rect 9328 253 9334 281
tri 9334 253 9362 281 sw
tri 9425 253 9453 281 se
rect 9453 253 9511 281
rect 9638 281 9910 287
rect 9912 286 9948 287
rect 4829 245 5034 253
rect 5086 245 5107 253
rect 5159 245 5180 253
rect 5232 245 5253 253
rect 5305 245 5838 253
rect 5890 245 5902 253
rect 5954 245 5966 253
rect 6018 245 6142 253
rect 4829 211 4844 245
rect 4878 211 4917 245
rect 4951 211 4990 245
rect 5024 211 5034 245
rect 5097 211 5107 245
rect 5170 211 5180 245
rect 5243 211 5253 245
rect 5316 211 5355 245
rect 5389 211 5428 245
rect 5462 211 5501 245
rect 5535 211 5574 245
rect 5608 211 5646 245
rect 5680 211 5718 245
rect 5752 211 5790 245
rect 5824 211 5838 245
rect 5896 211 5902 245
rect 6040 211 6078 245
rect 6112 211 6142 245
rect 4829 201 5034 211
rect 5086 201 5107 211
rect 5159 201 5180 211
rect 5232 201 5253 211
rect 5305 201 5838 211
rect 5890 201 5902 211
rect 5954 201 5966 211
rect 6018 201 6142 211
rect 6194 201 6211 253
rect 6263 201 6281 253
rect 6333 201 6351 253
rect 6403 201 6421 253
rect 6473 245 7505 253
rect 6473 211 6510 245
rect 6544 211 6582 245
rect 6616 211 6654 245
rect 6688 211 6726 245
rect 6760 211 6798 245
rect 6832 211 6870 245
rect 6904 211 6942 245
rect 6976 211 7014 245
rect 7048 211 7086 245
rect 7120 211 7158 245
rect 7192 211 7230 245
rect 7264 211 7302 245
rect 7336 211 7374 245
rect 7408 211 7446 245
rect 7480 211 7505 245
rect 6473 201 7505 211
rect 7557 201 7577 253
rect 7629 201 7649 253
rect 7701 201 7721 253
rect 7773 201 7793 253
rect 7845 201 7866 253
rect 7918 201 7939 253
rect 7991 201 8012 253
rect 8064 245 8187 253
rect 8239 245 8254 253
rect 8306 245 8322 253
rect 8374 245 8390 253
rect 8442 245 8953 253
rect 9005 245 9033 253
rect 9085 245 9114 253
rect 9166 245 9511 253
tri 9607 247 9638 278 se
rect 9638 247 9650 281
rect 9684 247 9722 281
rect 9756 247 9910 281
rect 8064 211 8094 245
rect 8128 211 8166 245
rect 8306 211 8310 245
rect 8374 211 8382 245
rect 8442 211 8454 245
rect 8488 211 8526 245
rect 8560 211 8598 245
rect 8632 211 8670 245
rect 8704 211 8742 245
rect 8776 211 8814 245
rect 8848 211 8886 245
rect 8920 211 8953 245
rect 9005 211 9030 245
rect 9085 211 9102 245
rect 9166 211 9174 245
rect 9208 211 9246 245
rect 9280 211 9318 245
rect 9352 211 9390 245
rect 9424 211 9462 245
rect 9496 211 9511 245
tri 9602 242 9607 247 se
rect 9607 242 9910 247
tri 9601 241 9602 242 se
rect 9602 241 9910 242
tri 9595 235 9601 241 se
rect 9601 235 9910 241
rect 9911 236 9949 286
rect 9912 235 9948 236
rect 9950 235 10086 287
rect 10138 235 10150 287
rect 10202 235 10208 287
rect 10431 235 10461 287
rect 10513 235 10525 287
rect 10577 235 10718 287
rect 10720 286 10756 287
rect 10719 236 10757 286
rect 10758 281 11011 287
rect 10758 247 10893 281
rect 10927 247 10965 281
rect 10999 247 11011 281
rect 10720 235 10756 236
rect 10758 235 11011 247
rect 8064 201 8187 211
rect 8239 201 8254 211
rect 8306 201 8322 211
rect 8374 201 8390 211
rect 8442 201 8953 211
rect 9005 201 9033 211
rect 9085 201 9114 211
rect 9166 201 9511 211
tri 9568 208 9595 235 se
rect 9595 208 9648 235
tri 9648 208 9675 235 nw
tri 10931 208 10958 235 ne
rect 10958 208 11011 235
tri 9567 207 9568 208 se
rect 9568 207 9647 208
tri 9647 207 9648 208 nw
tri 10958 207 10959 208 ne
tri 9565 205 9567 207 se
rect 9567 205 9609 207
tri 9561 201 9565 205 se
rect 9565 201 9609 205
tri 9559 199 9561 201 se
rect 9561 199 9609 201
tri 4239 177 4261 199 sw
tri 9537 177 9559 199 se
rect 9559 177 9609 199
tri 4187 169 4195 177 ne
rect 4195 169 4261 177
tri 4261 169 4269 177 sw
tri 9529 169 9537 177 se
rect 9537 169 9609 177
tri 9609 169 9647 207 nw
rect 3960 149 4018 169
tri 4018 149 4038 169 sw
tri 4195 149 4215 169 ne
rect 4215 149 4269 169
tri 3960 71 4038 149 ne
tri 4038 117 4070 149 sw
tri 4215 117 4247 149 ne
rect 4247 117 4269 149
tri 4269 117 4321 169 sw
rect 4749 117 4755 169
rect 4807 117 4819 169
rect 4871 117 8484 169
rect 8536 117 8548 169
rect 8600 117 8606 169
rect 8670 117 8676 169
rect 8728 117 8740 169
rect 8792 117 9557 169
tri 9557 117 9609 169 nw
rect 4038 85 4070 117
tri 4070 85 4102 117 sw
tri 4247 103 4261 117 ne
rect 4261 103 4321 117
tri 4321 103 4335 117 sw
tri 10949 103 10959 113 se
rect 10959 103 11011 208
tri 4261 85 4279 103 ne
rect 4279 85 4335 103
tri 4335 85 4353 103 sw
tri 10931 85 10949 103 se
rect 10949 85 11011 103
rect 4038 71 4102 85
tri 4102 71 4116 85 sw
tri 4279 71 4293 85 ne
rect 4293 76 4353 85
tri 4353 76 4362 85 sw
rect 4293 71 5246 76
tri 4038 -7 4116 71 ne
tri 4116 33 4154 71 sw
tri 4293 33 4331 71 ne
rect 4331 33 5246 71
tri 5246 33 5289 76 sw
rect 5377 33 5383 85
rect 5435 33 5447 85
rect 5499 33 11011 85
rect 11294 280 11300 314
rect 11334 280 11340 314
rect 12568 314 12614 326
tri 11340 280 11368 308 sw
tri 12540 280 12568 308 se
rect 12568 280 12574 314
rect 12608 280 12614 314
rect 11294 276 11368 280
tri 11368 276 11372 280 sw
tri 12536 276 12540 280 se
rect 12540 276 12614 280
rect 11294 242 11689 276
rect 11294 208 11300 242
rect 11334 224 11689 242
rect 11690 225 11691 275
rect 11727 225 11728 275
rect 11729 224 11840 276
rect 11892 224 11917 276
rect 11969 224 11994 276
rect 12046 224 12070 276
rect 12122 224 12206 276
rect 12207 225 12208 275
rect 12244 225 12245 275
rect 12246 242 12614 276
rect 12246 224 12574 242
rect 11334 208 11356 224
tri 11356 208 11372 224 nw
tri 12536 208 12552 224 ne
rect 12552 208 12574 224
rect 12608 208 12614 242
rect 4116 1 4154 33
tri 4154 1 4186 33 sw
tri 4331 29 4335 33 ne
rect 4335 29 5289 33
tri 5289 29 5293 33 sw
tri 4335 24 4340 29 ne
rect 4340 24 5293 29
tri 5293 24 5298 29 sw
tri 5224 1 5247 24 ne
rect 5247 1 5298 24
tri 5298 1 5321 24 sw
rect 4116 -2 4186 1
tri 4186 -2 4189 1 sw
tri 5247 -2 5250 1 ne
rect 5250 -2 5321 1
tri 5321 -2 5324 1 sw
tri 10077 -2 10080 1 se
rect 10080 -2 10086 1
rect 4116 -7 4189 -2
tri 4189 -7 4194 -2 sw
tri 4116 -8 4117 -7 ne
rect 4117 -8 4194 -7
tri 5250 -8 5256 -2 ne
rect 5256 -8 5324 -2
tri 5324 -8 5330 -2 sw
rect 8295 -8 10086 -2
tri 4117 -33 4142 -8 ne
rect 4142 -50 4194 -8
tri 5256 -42 5290 -8 ne
rect 5290 -32 5330 -8
tri 5330 -32 5354 -8 sw
rect 5290 -42 5354 -32
tri 5354 -42 5364 -32 sw
rect 8295 -42 8307 -8
rect 8341 -42 8379 -8
rect 8413 -42 10086 -8
tri 5290 -48 5296 -42 ne
rect 5296 -48 5364 -42
tri 5364 -48 5370 -42 sw
rect 8295 -48 10086 -42
tri 5296 -49 5297 -48 ne
rect 5297 -49 5370 -48
tri 4194 -50 4195 -49 sw
tri 5297 -50 5298 -49 ne
rect 5298 -50 5370 -49
tri 5370 -50 5372 -48 sw
tri 10077 -50 10079 -48 ne
rect 10079 -50 10086 -48
rect 4142 -51 4195 -50
tri 4195 -51 4196 -50 sw
tri 5298 -51 5299 -50 ne
rect 5299 -51 5372 -50
tri 5372 -51 5373 -50 sw
tri 10079 -51 10080 -50 ne
rect 10080 -51 10086 -50
rect 10138 -51 10150 1
rect 10202 -51 10208 1
rect 4142 -62 4196 -51
tri 4196 -62 4207 -51 sw
tri 5299 -62 5310 -51 ne
rect 5310 -54 5373 -51
tri 5373 -54 5376 -51 sw
rect 5310 -62 6842 -54
rect 4142 -83 4207 -62
tri 4207 -83 4228 -62 sw
tri 5310 -83 5331 -62 ne
rect 5331 -83 6842 -62
rect 4142 -135 4667 -83
rect 4719 -135 4743 -83
rect 4795 -135 4801 -83
tri 5331 -86 5334 -83 ne
rect 5334 -86 6842 -83
tri 5334 -92 5340 -86 ne
rect 5340 -92 6842 -86
tri 5340 -106 5354 -92 ne
rect 5354 -106 6842 -92
rect 6894 -106 6906 -54
rect 6958 -106 7974 -54
rect 8026 -106 8038 -54
rect 8090 -106 8096 -54
tri 10452 -86 10455 -83 se
rect 10455 -86 10461 -83
rect 9225 -132 10461 -86
tri 10452 -134 10454 -132 ne
rect 10454 -134 10461 -132
tri 10454 -135 10455 -134 ne
rect 10455 -135 10461 -134
rect 10513 -135 10525 -83
rect 10577 -85 10583 -83
tri 10583 -85 10585 -83 sw
rect 10577 -86 10585 -85
tri 10585 -86 10586 -85 sw
tri 11293 -86 11294 -85 se
rect 11294 -86 11340 208
tri 11340 192 11356 208 nw
tri 12552 192 12568 208 ne
rect 10577 -92 10907 -86
rect 10577 -126 10789 -92
rect 10823 -126 10861 -92
rect 10895 -126 10907 -92
tri 11279 -100 11293 -86 se
rect 11293 -100 11340 -86
rect 10577 -132 10907 -126
tri 11247 -132 11279 -100 se
rect 11279 -105 11340 -100
rect 11279 -132 11311 -105
rect 10577 -134 10584 -132
tri 10584 -134 10586 -132 nw
tri 11245 -134 11247 -132 se
rect 11247 -134 11311 -132
tri 11311 -134 11340 -105 nw
rect 12568 -28 12614 208
rect 12568 -62 12574 -28
rect 12608 -62 12614 -28
rect 12568 -100 12614 -62
rect 12568 -134 12574 -100
rect 12608 -134 12614 -100
rect 10577 -135 10583 -134
tri 10583 -135 10584 -134 nw
tri 11244 -135 11245 -134 se
rect 11245 -135 11299 -134
tri 11233 -146 11244 -135 se
rect 11244 -146 11299 -135
tri 11299 -146 11311 -134 nw
rect 12568 -146 12614 -134
tri 11228 -151 11233 -146 se
rect 11233 -151 11294 -146
tri 11294 -151 11299 -146 nw
tri 11213 -166 11228 -151 se
rect 11228 -166 11279 -151
tri 11279 -166 11294 -151 nw
rect 6496 -172 11233 -166
rect 6496 -206 6508 -172
rect 6542 -206 6580 -172
rect 6614 -206 11233 -172
rect 6496 -212 11233 -206
tri 11233 -212 11279 -166 nw
<< rmetal1 >>
rect 2842 3941 2844 3942
rect 2842 3897 2843 3941
rect 2842 3896 2844 3897
rect 2880 3941 2882 3942
rect 2881 3897 2882 3941
rect 2880 3896 2882 3897
rect 5012 3587 7014 3588
rect 5012 3586 5013 3587
rect 7013 3586 7014 3587
rect 5012 3549 5013 3550
rect 7013 3549 7014 3550
rect 5012 3548 7014 3549
rect 2829 3317 2831 3318
rect 2829 3273 2830 3317
rect 2829 3272 2831 3273
rect 2867 3317 2869 3318
rect 2868 3273 2869 3317
rect 2867 3272 2869 3273
rect 11880 3283 11882 3284
rect 11880 3239 11881 3283
rect 11880 3238 11882 3239
rect 11918 3283 11920 3284
rect 11919 3239 11920 3283
rect 11918 3238 11920 3239
rect 9334 2589 9336 2590
rect 9372 2589 9374 2590
rect 9334 2539 9335 2589
rect 9373 2539 9374 2589
rect 9334 2538 9336 2539
rect 9372 2538 9374 2539
rect 2909 2225 2911 2226
rect 2909 2181 2910 2225
rect 2909 2180 2911 2181
rect 2947 2225 2949 2226
rect 2948 2181 2949 2225
rect 2947 2180 2949 2181
rect 11880 2259 11882 2260
rect 11880 2215 11881 2259
rect 11880 2214 11882 2215
rect 11918 2259 11920 2260
rect 11919 2215 11920 2259
rect 11918 2214 11920 2215
rect 5012 1685 7014 1686
rect 5012 1684 5013 1685
rect 7013 1684 7014 1685
rect 5012 1647 5013 1648
rect 7013 1647 7014 1648
rect 5012 1646 7014 1647
rect 2854 1289 2856 1290
rect 2854 1245 2855 1289
rect 2854 1244 2856 1245
rect 2892 1289 2894 1290
rect 2893 1245 2894 1289
rect 2892 1244 2894 1245
rect 9910 286 9912 287
rect 9948 286 9950 287
rect 9910 236 9911 286
rect 9949 236 9950 286
rect 9910 235 9912 236
rect 9948 235 9950 236
rect 10718 286 10720 287
rect 10756 286 10758 287
rect 10718 236 10719 286
rect 10757 236 10758 286
rect 10718 235 10720 236
rect 10756 235 10758 236
rect 11689 275 11691 276
rect 11689 225 11690 275
rect 11689 224 11691 225
rect 11727 275 11729 276
rect 11728 225 11729 275
rect 11727 224 11729 225
rect 12206 275 12208 276
rect 12206 225 12207 275
rect 12206 224 12208 225
rect 12244 275 12246 276
rect 12245 225 12246 275
rect 12244 224 12246 225
<< via1 >>
rect 2379 13136 2431 13188
rect 2379 13072 2431 13124
rect 2471 13136 2523 13188
rect 10102 13172 10154 13224
rect 2471 13072 2523 13124
rect 10102 13108 10154 13160
rect 6152 13061 6204 13067
rect 6152 13027 6161 13061
rect 6161 13027 6195 13061
rect 6195 13027 6204 13061
rect 6152 13015 6204 13027
rect 6152 12989 6204 13001
rect 6152 12955 6161 12989
rect 6161 12955 6195 12989
rect 6195 12955 6204 12989
rect 6152 12949 6204 12955
rect 6152 12917 6204 12935
rect 6152 12883 6161 12917
rect 6161 12883 6195 12917
rect 6195 12883 6204 12917
rect 6152 12845 6204 12869
rect 6152 12817 6161 12845
rect 6161 12817 6195 12845
rect 6195 12817 6204 12845
rect 6152 12773 6204 12803
rect 6152 12751 6161 12773
rect 6161 12751 6195 12773
rect 6195 12751 6204 12773
rect 6152 12701 6204 12737
rect 6152 12685 6161 12701
rect 6161 12685 6195 12701
rect 6195 12685 6204 12701
rect 6152 12667 6161 12671
rect 6161 12667 6195 12671
rect 6195 12667 6204 12671
rect 6152 12629 6204 12667
rect 6152 12619 6161 12629
rect 6161 12619 6195 12629
rect 6195 12619 6204 12629
rect 6152 12595 6161 12605
rect 6161 12595 6195 12605
rect 6195 12595 6204 12605
rect 6152 12557 6204 12595
rect 6152 12553 6161 12557
rect 6161 12553 6195 12557
rect 6195 12553 6204 12557
rect 6152 12523 6161 12539
rect 6161 12523 6195 12539
rect 6195 12523 6204 12539
rect 6152 12487 6204 12523
rect 6152 12451 6161 12473
rect 6161 12451 6195 12473
rect 6195 12451 6204 12473
rect 6152 12421 6204 12451
rect 6152 12379 6161 12407
rect 6161 12379 6195 12407
rect 6195 12379 6204 12407
rect 6152 12355 6204 12379
rect 6152 12307 6161 12341
rect 6161 12307 6195 12341
rect 6195 12307 6204 12341
rect 6152 12289 6204 12307
rect 6152 12269 6204 12275
rect 6152 12235 6161 12269
rect 6161 12235 6195 12269
rect 6195 12235 6204 12269
rect 6152 12223 6204 12235
rect 6152 12197 6204 12209
rect 6152 12163 6161 12197
rect 6161 12163 6195 12197
rect 6195 12163 6204 12197
rect 6152 12157 6204 12163
rect 6152 12125 6204 12143
rect 6152 12091 6161 12125
rect 6161 12091 6195 12125
rect 6195 12091 6204 12125
rect 6152 12053 6204 12077
rect 6152 12025 6161 12053
rect 6161 12025 6195 12053
rect 6195 12025 6204 12053
rect 6152 11981 6204 12011
rect 6152 11959 6161 11981
rect 6161 11959 6195 11981
rect 6195 11959 6204 11981
rect 6152 11909 6204 11945
rect 6152 11893 6161 11909
rect 6161 11893 6195 11909
rect 6195 11893 6204 11909
rect 6152 11875 6161 11879
rect 6161 11875 6195 11879
rect 6195 11875 6204 11879
rect 6152 11837 6204 11875
rect 6152 11827 6161 11837
rect 6161 11827 6195 11837
rect 6195 11827 6204 11837
rect 6152 11803 6161 11813
rect 6161 11803 6195 11813
rect 6195 11803 6204 11813
rect 6152 11765 6204 11803
rect 6152 11761 6161 11765
rect 6161 11761 6195 11765
rect 6195 11761 6204 11765
rect 6152 11731 6161 11747
rect 6161 11731 6195 11747
rect 6195 11731 6204 11747
rect 6152 11695 6204 11731
rect 2471 11627 2523 11679
rect 6152 11659 6161 11681
rect 6161 11659 6195 11681
rect 6195 11659 6204 11681
rect 6152 11629 6204 11659
rect 2471 11563 2523 11615
rect 6152 11587 6161 11615
rect 6161 11587 6195 11615
rect 6195 11587 6204 11615
rect 6152 11563 6204 11587
rect 6152 11515 6161 11549
rect 6161 11515 6195 11549
rect 6195 11515 6204 11549
rect 6152 11497 6204 11515
rect 6152 11477 6204 11483
rect 6152 11443 6161 11477
rect 6161 11443 6195 11477
rect 6195 11443 6204 11477
rect 6152 11431 6204 11443
rect 6152 11405 6204 11417
rect 6152 11371 6161 11405
rect 6161 11371 6195 11405
rect 6195 11371 6204 11405
rect 6152 11365 6204 11371
rect 6152 11333 6204 11351
rect 6152 11299 6161 11333
rect 6161 11299 6195 11333
rect 6195 11299 6204 11333
rect 11266 11319 11318 11325
rect 11330 11319 11382 11325
rect 11266 11285 11290 11319
rect 11290 11285 11318 11319
rect 11330 11285 11365 11319
rect 11365 11285 11382 11319
rect 6152 11232 6204 11284
rect 6152 11199 6204 11217
rect 11266 11273 11318 11285
rect 11330 11273 11382 11285
rect 6152 11165 6167 11199
rect 6167 11165 6201 11199
rect 6201 11165 6204 11199
rect 2350 11061 2402 11113
rect 2414 11061 2466 11113
rect 7068 11014 7120 11017
rect 7068 10980 7070 11014
rect 7070 10980 7104 11014
rect 7104 10980 7120 11014
rect 7068 10965 7120 10980
rect 7144 11014 7196 11017
rect 7144 10980 7149 11014
rect 7149 10980 7183 11014
rect 7183 10980 7196 11014
rect 7144 10965 7196 10980
rect 7220 11014 7272 11017
rect 7220 10980 7228 11014
rect 7228 10980 7262 11014
rect 7262 10980 7272 11014
rect 7220 10965 7272 10980
rect 7296 11014 7348 11017
rect 7296 10980 7306 11014
rect 7306 10980 7340 11014
rect 7340 10980 7348 11014
rect 7296 10965 7348 10980
rect 7372 11014 7424 11017
rect 7372 10980 7384 11014
rect 7384 10980 7418 11014
rect 7418 10980 7424 11014
rect 7372 10965 7424 10980
rect 7447 11014 7499 11017
rect 7447 10980 7462 11014
rect 7462 10980 7496 11014
rect 7496 10980 7499 11014
rect 7447 10965 7499 10980
rect 7068 10936 7120 10953
rect 7068 10902 7070 10936
rect 7070 10902 7104 10936
rect 7104 10902 7120 10936
rect 7068 10901 7120 10902
rect 7144 10936 7196 10953
rect 7144 10902 7149 10936
rect 7149 10902 7183 10936
rect 7183 10902 7196 10936
rect 7144 10901 7196 10902
rect 7220 10936 7272 10953
rect 7220 10902 7228 10936
rect 7228 10902 7262 10936
rect 7262 10902 7272 10936
rect 7220 10901 7272 10902
rect 7296 10936 7348 10953
rect 7296 10902 7306 10936
rect 7306 10902 7340 10936
rect 7340 10902 7348 10936
rect 7296 10901 7348 10902
rect 7372 10936 7424 10953
rect 7372 10902 7384 10936
rect 7384 10902 7418 10936
rect 7418 10902 7424 10936
rect 7372 10901 7424 10902
rect 7447 10936 7499 10953
rect 7447 10902 7462 10936
rect 7462 10902 7496 10936
rect 7496 10902 7499 10936
rect 7447 10901 7499 10902
rect 326 10666 378 10672
rect 326 10632 332 10666
rect 332 10632 366 10666
rect 366 10632 378 10666
rect 326 10620 378 10632
rect 326 10594 378 10608
rect 326 10560 332 10594
rect 332 10560 366 10594
rect 366 10560 378 10594
rect 326 10556 378 10560
rect 11266 10437 11318 10443
rect 11330 10437 11382 10443
rect 11266 10403 11302 10437
rect 11302 10403 11318 10437
rect 11330 10403 11336 10437
rect 11336 10403 11374 10437
rect 11374 10403 11382 10437
rect 11266 10391 11318 10403
rect 11330 10391 11382 10403
rect 7067 10098 7069 10132
rect 7069 10098 7103 10132
rect 7103 10098 7119 10132
rect 7067 10080 7119 10098
rect 7131 10098 7147 10132
rect 7147 10098 7181 10132
rect 7181 10098 7183 10132
rect 7131 10080 7183 10098
rect 7195 10098 7225 10132
rect 7225 10098 7247 10132
rect 7195 10080 7247 10098
rect 7259 10080 7311 10132
rect 7323 10098 7372 10132
rect 7372 10098 7375 10132
rect 7387 10098 7406 10132
rect 7406 10098 7439 10132
rect 7451 10098 7478 10132
rect 7478 10098 7503 10132
rect 7323 10080 7375 10098
rect 7387 10080 7439 10098
rect 7451 10080 7503 10098
rect 7067 10051 7119 10065
rect 7067 10017 7069 10051
rect 7069 10017 7103 10051
rect 7103 10017 7119 10051
rect 7067 10013 7119 10017
rect 7131 10051 7183 10065
rect 7131 10017 7147 10051
rect 7147 10017 7181 10051
rect 7181 10017 7183 10051
rect 7131 10013 7183 10017
rect 7195 10051 7247 10065
rect 7195 10017 7225 10051
rect 7225 10017 7247 10051
rect 7195 10013 7247 10017
rect 7259 10013 7311 10065
rect 7323 10051 7375 10065
rect 7387 10051 7439 10065
rect 7451 10051 7503 10065
rect 7323 10017 7372 10051
rect 7372 10017 7375 10051
rect 7387 10017 7406 10051
rect 7406 10017 7439 10051
rect 7451 10017 7478 10051
rect 7478 10017 7503 10051
rect 7323 10013 7375 10017
rect 7387 10013 7439 10017
rect 7451 10013 7503 10017
rect 7067 9970 7119 9998
rect 7067 9946 7069 9970
rect 7069 9946 7103 9970
rect 7103 9946 7119 9970
rect 7131 9970 7183 9998
rect 7131 9946 7147 9970
rect 7147 9946 7181 9970
rect 7181 9946 7183 9970
rect 7195 9970 7247 9998
rect 7195 9946 7225 9970
rect 7225 9946 7247 9970
rect 7259 9946 7311 9998
rect 7323 9970 7375 9998
rect 7387 9970 7439 9998
rect 7451 9970 7503 9998
rect 7323 9946 7372 9970
rect 7372 9946 7375 9970
rect 7387 9946 7406 9970
rect 7406 9946 7439 9970
rect 7451 9946 7478 9970
rect 7478 9946 7503 9970
rect 7067 9889 7119 9930
rect 7067 9878 7069 9889
rect 7069 9878 7103 9889
rect 7103 9878 7119 9889
rect 7131 9889 7183 9930
rect 7131 9878 7147 9889
rect 7147 9878 7181 9889
rect 7181 9878 7183 9889
rect 7195 9889 7247 9930
rect 7195 9878 7225 9889
rect 7225 9878 7247 9889
rect 7259 9878 7311 9930
rect 7323 9889 7375 9930
rect 7387 9889 7439 9930
rect 7451 9889 7503 9930
rect 7323 9878 7372 9889
rect 7372 9878 7375 9889
rect 7387 9878 7406 9889
rect 7406 9878 7439 9889
rect 7451 9878 7478 9889
rect 7478 9878 7503 9889
rect 7067 9855 7069 9862
rect 7069 9855 7103 9862
rect 7103 9855 7119 9862
rect 7067 9810 7119 9855
rect 7131 9855 7147 9862
rect 7147 9855 7181 9862
rect 7181 9855 7183 9862
rect 7131 9810 7183 9855
rect 7195 9855 7225 9862
rect 7225 9855 7247 9862
rect 7195 9810 7247 9855
rect 7259 9810 7311 9862
rect 7323 9855 7372 9862
rect 7372 9855 7375 9862
rect 7387 9855 7406 9862
rect 7406 9855 7439 9862
rect 7451 9855 7478 9862
rect 7478 9855 7503 9862
rect 7323 9810 7375 9855
rect 7387 9810 7439 9855
rect 7451 9810 7503 9855
rect 7067 9773 7069 9794
rect 7069 9773 7103 9794
rect 7103 9773 7119 9794
rect 7067 9742 7119 9773
rect 7131 9773 7147 9794
rect 7147 9773 7181 9794
rect 7181 9773 7183 9794
rect 7131 9742 7183 9773
rect 7195 9773 7225 9794
rect 7225 9773 7247 9794
rect 7195 9742 7247 9773
rect 7259 9742 7311 9794
rect 7323 9773 7372 9794
rect 7372 9773 7375 9794
rect 7387 9773 7406 9794
rect 7406 9773 7439 9794
rect 7451 9773 7478 9794
rect 7478 9773 7503 9794
rect 7323 9742 7375 9773
rect 7387 9742 7439 9773
rect 7451 9742 7503 9773
rect 7067 9725 7119 9726
rect 7067 9691 7069 9725
rect 7069 9691 7103 9725
rect 7103 9691 7119 9725
rect 7067 9674 7119 9691
rect 7131 9725 7183 9726
rect 7131 9691 7147 9725
rect 7147 9691 7181 9725
rect 7181 9691 7183 9725
rect 7131 9674 7183 9691
rect 7195 9725 7247 9726
rect 7195 9691 7225 9725
rect 7225 9691 7247 9725
rect 7195 9674 7247 9691
rect 7259 9674 7311 9726
rect 7323 9725 7375 9726
rect 7387 9725 7439 9726
rect 7451 9725 7503 9726
rect 7323 9691 7372 9725
rect 7372 9691 7375 9725
rect 7387 9691 7406 9725
rect 7406 9691 7439 9725
rect 7451 9691 7478 9725
rect 7478 9691 7503 9725
rect 7323 9674 7375 9691
rect 7387 9674 7439 9691
rect 7451 9674 7503 9691
rect 7067 9643 7119 9658
rect 7067 9609 7069 9643
rect 7069 9609 7103 9643
rect 7103 9609 7119 9643
rect 7067 9606 7119 9609
rect 7131 9643 7183 9658
rect 7131 9609 7147 9643
rect 7147 9609 7181 9643
rect 7181 9609 7183 9643
rect 7131 9606 7183 9609
rect 7195 9643 7247 9658
rect 7195 9609 7225 9643
rect 7225 9609 7247 9643
rect 7195 9606 7247 9609
rect 7259 9606 7311 9658
rect 7323 9643 7375 9658
rect 7387 9643 7439 9658
rect 7451 9643 7503 9658
rect 7323 9609 7372 9643
rect 7372 9609 7375 9643
rect 7387 9609 7406 9643
rect 7406 9609 7439 9643
rect 7451 9609 7478 9643
rect 7478 9609 7503 9643
rect 7323 9606 7375 9609
rect 7387 9606 7439 9609
rect 7451 9606 7503 9609
rect 10331 9507 10383 9559
rect 10395 9507 10447 9559
rect 11266 9507 11318 9559
rect 11330 9507 11382 9559
rect 7067 9368 7069 9402
rect 7069 9368 7103 9402
rect 7103 9368 7119 9402
rect 7067 9350 7119 9368
rect 7131 9368 7147 9402
rect 7147 9368 7181 9402
rect 7181 9368 7183 9402
rect 7131 9350 7183 9368
rect 7195 9368 7225 9402
rect 7225 9368 7247 9402
rect 7195 9350 7247 9368
rect 7259 9350 7311 9402
rect 7323 9368 7372 9402
rect 7372 9368 7375 9402
rect 7387 9368 7406 9402
rect 7406 9368 7439 9402
rect 7451 9368 7478 9402
rect 7478 9368 7503 9402
rect 7323 9350 7375 9368
rect 7387 9350 7439 9368
rect 7451 9350 7503 9368
rect 7067 9321 7119 9335
rect 7067 9287 7069 9321
rect 7069 9287 7103 9321
rect 7103 9287 7119 9321
rect 7067 9283 7119 9287
rect 7131 9321 7183 9335
rect 7131 9287 7147 9321
rect 7147 9287 7181 9321
rect 7181 9287 7183 9321
rect 7131 9283 7183 9287
rect 7195 9321 7247 9335
rect 7195 9287 7225 9321
rect 7225 9287 7247 9321
rect 7195 9283 7247 9287
rect 7259 9283 7311 9335
rect 7323 9321 7375 9335
rect 7387 9321 7439 9335
rect 7451 9321 7503 9335
rect 7323 9287 7372 9321
rect 7372 9287 7375 9321
rect 7387 9287 7406 9321
rect 7406 9287 7439 9321
rect 7451 9287 7478 9321
rect 7478 9287 7503 9321
rect 7323 9283 7375 9287
rect 7387 9283 7439 9287
rect 7451 9283 7503 9287
rect 7067 9240 7119 9268
rect 7067 9216 7069 9240
rect 7069 9216 7103 9240
rect 7103 9216 7119 9240
rect 7131 9240 7183 9268
rect 7131 9216 7147 9240
rect 7147 9216 7181 9240
rect 7181 9216 7183 9240
rect 7195 9240 7247 9268
rect 7195 9216 7225 9240
rect 7225 9216 7247 9240
rect 7259 9216 7311 9268
rect 7323 9240 7375 9268
rect 7387 9240 7439 9268
rect 7451 9240 7503 9268
rect 7323 9216 7372 9240
rect 7372 9216 7375 9240
rect 7387 9216 7406 9240
rect 7406 9216 7439 9240
rect 7451 9216 7478 9240
rect 7478 9216 7503 9240
rect 7067 9159 7119 9200
rect 7067 9148 7069 9159
rect 7069 9148 7103 9159
rect 7103 9148 7119 9159
rect 7131 9159 7183 9200
rect 7131 9148 7147 9159
rect 7147 9148 7181 9159
rect 7181 9148 7183 9159
rect 7195 9159 7247 9200
rect 7195 9148 7225 9159
rect 7225 9148 7247 9159
rect 7259 9148 7311 9200
rect 7323 9159 7375 9200
rect 7387 9159 7439 9200
rect 7451 9159 7503 9200
rect 7323 9148 7372 9159
rect 7372 9148 7375 9159
rect 7387 9148 7406 9159
rect 7406 9148 7439 9159
rect 7451 9148 7478 9159
rect 7478 9148 7503 9159
rect 7067 9125 7069 9132
rect 7069 9125 7103 9132
rect 7103 9125 7119 9132
rect 7067 9080 7119 9125
rect 7131 9125 7147 9132
rect 7147 9125 7181 9132
rect 7181 9125 7183 9132
rect 7131 9080 7183 9125
rect 7195 9125 7225 9132
rect 7225 9125 7247 9132
rect 7195 9080 7247 9125
rect 7259 9080 7311 9132
rect 7323 9125 7372 9132
rect 7372 9125 7375 9132
rect 7387 9125 7406 9132
rect 7406 9125 7439 9132
rect 7451 9125 7478 9132
rect 7478 9125 7503 9132
rect 7323 9080 7375 9125
rect 7387 9080 7439 9125
rect 7451 9080 7503 9125
rect 7067 9043 7069 9064
rect 7069 9043 7103 9064
rect 7103 9043 7119 9064
rect 7067 9012 7119 9043
rect 7131 9043 7147 9064
rect 7147 9043 7181 9064
rect 7181 9043 7183 9064
rect 7131 9012 7183 9043
rect 7195 9043 7225 9064
rect 7225 9043 7247 9064
rect 7195 9012 7247 9043
rect 7259 9012 7311 9064
rect 7323 9043 7372 9064
rect 7372 9043 7375 9064
rect 7387 9043 7406 9064
rect 7406 9043 7439 9064
rect 7451 9043 7478 9064
rect 7478 9043 7503 9064
rect 7323 9012 7375 9043
rect 7387 9012 7439 9043
rect 7451 9012 7503 9043
rect 7067 8995 7119 8996
rect 7067 8961 7069 8995
rect 7069 8961 7103 8995
rect 7103 8961 7119 8995
rect 7067 8944 7119 8961
rect 7131 8995 7183 8996
rect 7131 8961 7147 8995
rect 7147 8961 7181 8995
rect 7181 8961 7183 8995
rect 7131 8944 7183 8961
rect 7195 8995 7247 8996
rect 7195 8961 7225 8995
rect 7225 8961 7247 8995
rect 7195 8944 7247 8961
rect 7259 8944 7311 8996
rect 7323 8995 7375 8996
rect 7387 8995 7439 8996
rect 7451 8995 7503 8996
rect 7323 8961 7372 8995
rect 7372 8961 7375 8995
rect 7387 8961 7406 8995
rect 7406 8961 7439 8995
rect 7451 8961 7478 8995
rect 7478 8961 7503 8995
rect 7323 8944 7375 8961
rect 7387 8944 7439 8961
rect 7451 8944 7503 8961
rect 7067 8913 7119 8928
rect 7067 8879 7069 8913
rect 7069 8879 7103 8913
rect 7103 8879 7119 8913
rect 7067 8876 7119 8879
rect 7131 8913 7183 8928
rect 7131 8879 7147 8913
rect 7147 8879 7181 8913
rect 7181 8879 7183 8913
rect 7131 8876 7183 8879
rect 7195 8913 7247 8928
rect 7195 8879 7225 8913
rect 7225 8879 7247 8913
rect 7195 8876 7247 8879
rect 7259 8876 7311 8928
rect 7323 8913 7375 8928
rect 7387 8913 7439 8928
rect 7451 8913 7503 8928
rect 7323 8879 7372 8913
rect 7372 8879 7375 8913
rect 7387 8879 7406 8913
rect 7406 8879 7439 8913
rect 7451 8879 7478 8913
rect 7478 8879 7503 8913
rect 7323 8876 7375 8879
rect 7387 8876 7439 8879
rect 7451 8876 7503 8879
rect 4831 8517 4883 8569
rect 4895 8517 4947 8569
rect 13697 8273 13749 8325
rect 13761 8273 13813 8325
rect 153 7797 205 7849
rect 217 7797 269 7849
rect 884 7797 936 7849
rect 948 7797 1000 7849
rect 12649 7194 12701 7246
rect 12733 7194 12785 7246
rect 12818 7194 12870 7246
rect 12903 7194 12955 7246
rect 12997 7194 13049 7246
rect 13069 7194 13121 7246
rect 13141 7194 13193 7246
rect 13213 7194 13265 7246
rect 13286 7194 13338 7246
rect 13879 6791 13995 6907
rect 13767 6695 13819 6747
rect 13767 6631 13819 6683
rect -87 6181 -35 6233
rect 2931 6237 2983 6289
rect -87 6117 -35 6169
rect 244 6147 296 6153
rect 244 6113 250 6147
rect 250 6113 284 6147
rect 284 6113 296 6147
rect 766 6147 818 6153
rect 244 6101 296 6113
rect 445 6094 497 6146
rect 509 6094 561 6146
rect 573 6094 625 6146
rect 766 6113 778 6147
rect 778 6113 812 6147
rect 812 6113 818 6147
rect 766 6101 818 6113
rect 244 6041 296 6086
rect 244 6034 250 6041
rect 250 6034 284 6041
rect 284 6034 296 6041
rect 244 6007 250 6019
rect 250 6007 284 6019
rect 284 6007 296 6019
rect 766 6061 818 6073
rect 766 6027 778 6061
rect 778 6027 812 6061
rect 812 6027 818 6061
rect 958 6144 1010 6150
rect 958 6110 967 6144
rect 967 6110 1001 6144
rect 1001 6110 1010 6144
rect 958 6098 1010 6110
rect 1156 6094 1208 6146
rect 1225 6094 1277 6146
rect 1294 6094 1346 6146
rect 1471 6144 1523 6150
rect 2931 6169 2983 6221
rect 4637 6163 4689 6215
rect 1471 6110 1480 6144
rect 1480 6110 1514 6144
rect 1514 6110 1523 6144
rect 1471 6098 1523 6110
rect 958 6056 1010 6068
rect 766 6021 818 6027
rect 244 5969 296 6007
rect 878 5992 930 6044
rect 958 6022 967 6056
rect 967 6022 1001 6056
rect 1001 6022 1010 6056
rect 958 6016 1010 6022
rect 1471 6069 1523 6085
rect 1471 6035 1480 6069
rect 1480 6035 1514 6069
rect 1514 6035 1523 6069
rect 1471 6033 1523 6035
rect 1471 5994 1523 6020
rect 244 5967 250 5969
rect 250 5967 284 5969
rect 284 5967 296 5969
rect 244 5935 250 5952
rect 250 5935 284 5952
rect 284 5935 296 5952
rect 244 5900 296 5935
rect 244 5853 250 5885
rect 250 5853 284 5885
rect 284 5853 296 5885
rect 244 5833 296 5853
rect 244 5804 296 5818
rect 244 5770 250 5804
rect 250 5770 284 5804
rect 284 5770 296 5804
rect 244 5766 296 5770
rect 244 5721 296 5751
rect 244 5699 250 5721
rect 250 5699 284 5721
rect 284 5699 296 5721
rect 244 5638 296 5684
rect 244 5632 250 5638
rect 250 5632 284 5638
rect 284 5632 296 5638
rect 244 5604 250 5617
rect 250 5604 284 5617
rect 284 5604 296 5617
rect 244 5565 296 5604
rect 244 5521 250 5550
rect 250 5521 284 5550
rect 284 5521 296 5550
rect 244 5498 296 5521
rect 244 5472 296 5484
rect 244 5438 250 5472
rect 250 5438 284 5472
rect 284 5438 296 5472
rect 244 5432 296 5438
rect 878 5927 930 5979
rect 1471 5968 1480 5994
rect 1480 5968 1514 5994
rect 1514 5968 1523 5994
rect 1471 5919 1523 5955
rect 1471 5903 1480 5919
rect 1480 5903 1514 5919
rect 1514 5903 1523 5919
rect 445 5742 497 5794
rect 509 5742 561 5794
rect 573 5742 625 5794
rect 769 5881 821 5887
rect 769 5847 778 5881
rect 778 5847 812 5881
rect 812 5847 821 5881
rect 769 5835 821 5847
rect 769 5786 821 5795
rect 769 5752 778 5786
rect 778 5752 812 5786
rect 812 5752 821 5786
rect 769 5743 821 5752
rect 769 5691 821 5703
rect 769 5657 778 5691
rect 778 5657 812 5691
rect 812 5657 821 5691
rect 769 5651 821 5657
rect 958 5881 1010 5887
rect 958 5847 967 5881
rect 967 5847 1001 5881
rect 1001 5847 1010 5881
rect 958 5835 1010 5847
rect 958 5786 1010 5795
rect 958 5752 967 5786
rect 967 5752 1001 5786
rect 1001 5752 1010 5786
rect 958 5743 1010 5752
rect 958 5691 1010 5703
rect 958 5657 967 5691
rect 967 5657 1001 5691
rect 1001 5657 1010 5691
rect 958 5651 1010 5657
rect 1471 5885 1480 5890
rect 1480 5885 1514 5890
rect 1514 5885 1523 5890
rect 3023 6065 3075 6117
rect 3023 5997 3075 6049
rect 4637 6094 4689 6146
rect 4637 6025 4689 6077
rect 4637 5956 4689 6008
rect 4637 5887 4689 5939
rect 1471 5843 1523 5885
rect 1471 5838 1480 5843
rect 1480 5838 1514 5843
rect 1514 5838 1523 5843
rect 1471 5809 1480 5825
rect 1480 5809 1514 5825
rect 1514 5809 1523 5825
rect 1156 5742 1208 5794
rect 1225 5742 1277 5794
rect 1294 5742 1346 5794
rect 1471 5773 1523 5809
rect 1471 5733 1480 5759
rect 1480 5733 1514 5759
rect 1514 5733 1523 5759
rect 4637 5818 4689 5870
rect 4637 5749 4689 5801
rect 1471 5707 1523 5733
rect 1471 5691 1523 5693
rect 1471 5657 1480 5691
rect 1480 5657 1514 5691
rect 1514 5657 1523 5691
rect 4637 5679 4689 5731
rect 1471 5641 1523 5657
rect 1471 5615 1523 5627
rect 1471 5581 1480 5615
rect 1480 5581 1514 5615
rect 1514 5581 1523 5615
rect 3023 5604 3075 5656
rect 1471 5575 1523 5581
rect 160 5350 212 5402
rect 445 5390 497 5442
rect 509 5390 561 5442
rect 573 5390 625 5442
rect 160 5286 212 5338
rect 769 5526 821 5532
rect 769 5492 778 5526
rect 778 5492 812 5526
rect 812 5492 821 5526
rect 769 5480 821 5492
rect 769 5420 821 5467
rect 769 5415 778 5420
rect 778 5415 812 5420
rect 812 5415 821 5420
rect 769 5386 778 5403
rect 778 5386 812 5403
rect 812 5386 821 5403
rect 769 5351 821 5386
rect 769 5315 821 5339
rect 769 5287 778 5315
rect 778 5287 812 5315
rect 812 5287 821 5315
rect 769 5223 821 5275
rect 1043 5483 1095 5535
rect 3023 5540 3075 5592
rect 11859 5534 11911 5586
rect 11923 5534 11975 5586
rect 958 5447 1010 5453
rect 958 5413 967 5447
rect 967 5413 1001 5447
rect 1001 5413 1010 5447
rect 1043 5419 1095 5471
rect 1471 5451 1523 5458
rect 1471 5417 1480 5451
rect 1480 5417 1514 5451
rect 1514 5417 1523 5451
rect 958 5401 1010 5413
rect 958 5357 1010 5382
rect 1471 5406 1523 5417
rect 1471 5378 1523 5393
rect 958 5330 967 5357
rect 967 5330 1001 5357
rect 1001 5330 1010 5357
rect 1471 5344 1480 5378
rect 1480 5344 1514 5378
rect 1514 5344 1523 5378
rect 958 5267 1010 5311
rect 958 5259 967 5267
rect 967 5259 1001 5267
rect 1001 5259 1010 5267
rect 958 5233 967 5241
rect 967 5233 1001 5241
rect 1001 5233 1010 5241
rect 958 5189 1010 5233
rect 958 5144 967 5171
rect 967 5144 1001 5171
rect 1001 5144 1010 5171
rect 958 5119 1010 5144
rect 244 5095 296 5101
rect 244 5061 250 5095
rect 250 5061 284 5095
rect 284 5061 296 5095
rect 244 5049 296 5061
rect 244 5017 296 5033
rect 244 4983 250 5017
rect 250 4983 284 5017
rect 284 4983 296 5017
rect 244 4981 296 4983
rect 244 4939 296 4965
rect 244 4913 250 4939
rect 250 4913 284 4939
rect 284 4913 296 4939
rect 244 4861 296 4897
rect 244 4845 250 4861
rect 250 4845 284 4861
rect 284 4845 296 4861
rect 244 4827 250 4829
rect 250 4827 284 4829
rect 284 4827 296 4829
rect 244 4782 296 4827
rect 244 4777 250 4782
rect 250 4777 284 4782
rect 284 4777 296 4782
rect 244 4748 250 4761
rect 250 4748 284 4761
rect 284 4748 296 4761
rect 244 4709 296 4748
rect 244 4669 250 4693
rect 250 4669 284 4693
rect 284 4669 296 4693
rect 244 4641 296 4669
rect 244 4624 296 4625
rect 244 4590 250 4624
rect 250 4590 284 4624
rect 284 4590 296 4624
rect 244 4573 296 4590
rect 244 4545 296 4557
rect 244 4511 250 4545
rect 250 4511 284 4545
rect 284 4511 296 4545
rect 244 4505 296 4511
rect 445 5038 497 5090
rect 509 5038 561 5090
rect 573 5038 625 5090
rect 958 5089 1010 5101
rect 958 5055 967 5089
rect 967 5055 1001 5089
rect 1001 5055 1010 5089
rect 958 5049 1010 5055
rect 1471 5341 1523 5344
rect 1471 5305 1523 5328
rect 1471 5276 1480 5305
rect 1480 5276 1514 5305
rect 1514 5276 1523 5305
rect 1221 5200 1273 5252
rect 1285 5200 1337 5252
rect 1471 5232 1523 5263
rect 1471 5211 1480 5232
rect 1480 5211 1514 5232
rect 1514 5211 1523 5232
rect 1769 5330 1885 5510
rect 2750 5464 2802 5516
rect 2750 5400 2802 5452
rect 2937 5378 2989 5430
rect 3005 5378 3057 5430
rect 4831 5359 4883 5411
rect 4895 5359 4947 5411
rect 2836 5295 2888 5347
rect 2900 5295 2952 5347
rect 3590 5208 3642 5260
rect 1471 5159 1523 5198
rect 1471 5146 1480 5159
rect 1480 5146 1514 5159
rect 1514 5146 1523 5159
rect 1471 5125 1480 5133
rect 1480 5125 1514 5133
rect 1514 5125 1523 5133
rect 1471 5086 1523 5125
rect 1471 5081 1480 5086
rect 1480 5081 1514 5086
rect 1514 5081 1523 5086
rect 1471 5052 1480 5068
rect 1480 5052 1514 5068
rect 1514 5052 1523 5068
rect 1471 5016 1523 5052
rect 699 4931 751 4983
rect 763 4931 815 4983
rect 1471 4979 1480 5003
rect 1480 4979 1514 5003
rect 1514 4979 1523 5003
rect 1471 4951 1523 4979
rect 1471 4906 1480 4938
rect 1480 4906 1514 4938
rect 1514 4906 1523 4938
rect 1471 4886 1523 4906
rect 445 4772 497 4824
rect 509 4772 561 4824
rect 573 4772 625 4824
rect 687 4689 739 4741
rect 687 4625 739 4677
rect 849 4747 901 4799
rect 849 4683 901 4735
rect 409 4542 461 4551
rect 409 4508 415 4542
rect 415 4508 449 4542
rect 449 4508 461 4542
rect 409 4499 461 4508
rect 495 4542 547 4551
rect 582 4542 634 4551
rect 495 4508 496 4542
rect 496 4508 530 4542
rect 530 4508 547 4542
rect 582 4508 611 4542
rect 611 4508 634 4542
rect 495 4499 547 4508
rect 582 4499 634 4508
rect 958 4635 1010 4641
rect 958 4601 967 4635
rect 967 4601 1001 4635
rect 1001 4601 1010 4635
rect 958 4589 1010 4601
rect 958 4558 1010 4565
rect 958 4524 967 4558
rect 967 4524 1001 4558
rect 1001 4524 1010 4558
rect 958 4513 1010 4524
rect 958 4481 1010 4490
rect 958 4447 967 4481
rect 967 4447 1001 4481
rect 1001 4447 1010 4481
rect 958 4438 1010 4447
rect 958 4405 1010 4415
rect 958 4371 967 4405
rect 967 4371 1001 4405
rect 1001 4371 1010 4405
rect 958 4363 1010 4371
rect 958 4329 1010 4340
rect 958 4295 967 4329
rect 967 4295 1001 4329
rect 1001 4295 1010 4329
rect 958 4288 1010 4295
rect 958 4253 1010 4265
rect 958 4219 967 4253
rect 967 4219 1001 4253
rect 1001 4219 1010 4253
rect 958 4213 1010 4219
rect 849 4043 901 4095
rect 849 3979 901 4031
rect 849 3915 901 3967
rect 958 3859 1010 3865
rect 958 3825 967 3859
rect 967 3825 1001 3859
rect 1001 3825 1010 3859
rect 958 3813 1010 3825
rect 958 3785 1010 3792
rect 958 3751 967 3785
rect 967 3751 1001 3785
rect 1001 3751 1010 3785
rect 1156 3759 1208 3811
rect 1220 3759 1272 3811
rect 1284 3759 1336 3811
rect 958 3740 1010 3751
rect 958 3711 1010 3720
rect 958 3677 967 3711
rect 967 3677 1001 3711
rect 1001 3677 1010 3711
rect 769 3614 821 3666
rect 769 3550 821 3602
rect 958 3668 1010 3677
rect 958 3638 1010 3648
rect 958 3604 967 3638
rect 967 3604 1001 3638
rect 1001 3604 1010 3638
rect 958 3596 1010 3604
rect 958 3565 1010 3576
rect 958 3531 967 3565
rect 967 3531 1001 3565
rect 1001 3531 1010 3565
rect 958 3524 1010 3531
rect 240 3442 292 3494
rect 958 3492 1010 3504
rect 958 3458 967 3492
rect 967 3458 1001 3492
rect 1001 3458 1010 3492
rect 958 3452 1010 3458
rect 1156 3581 1208 3633
rect 1220 3581 1272 3633
rect 1284 3581 1336 3633
rect 1471 4867 1523 4873
rect 1471 4833 1480 4867
rect 1480 4833 1514 4867
rect 1514 4833 1523 4867
rect 1471 4821 1523 4833
rect 1471 4794 1523 4808
rect 1471 4760 1480 4794
rect 1480 4760 1514 4794
rect 1514 4760 1523 4794
rect 1471 4756 1523 4760
rect 1471 4721 1523 4743
rect 1471 4691 1480 4721
rect 1480 4691 1514 4721
rect 1514 4691 1523 4721
rect 1471 4648 1523 4678
rect 1471 4626 1480 4648
rect 1480 4626 1514 4648
rect 1514 4626 1523 4648
rect 1471 4575 1523 4613
rect 1471 4561 1480 4575
rect 1480 4561 1514 4575
rect 1514 4561 1523 4575
rect 1471 4541 1480 4548
rect 1480 4541 1514 4548
rect 1514 4541 1523 4548
rect 1471 4502 1523 4541
rect 1471 4496 1480 4502
rect 1480 4496 1514 4502
rect 1514 4496 1523 4502
rect 1471 4468 1480 4483
rect 1480 4468 1514 4483
rect 1514 4468 1523 4483
rect 1471 4431 1523 4468
rect 1471 4395 1480 4418
rect 1480 4395 1514 4418
rect 1514 4395 1523 4418
rect 1471 4366 1523 4395
rect 1471 4322 1480 4353
rect 1480 4322 1514 4353
rect 1514 4322 1523 4353
rect 1471 4301 1523 4322
rect 1471 4283 1523 4287
rect 1471 4249 1480 4283
rect 1480 4249 1514 4283
rect 1514 4249 1523 4283
rect 1471 4235 1523 4249
rect 1471 4210 1523 4221
rect 1471 4176 1480 4210
rect 1480 4176 1514 4210
rect 1514 4176 1523 4210
rect 1471 4169 1523 4176
rect 1471 4137 1523 4155
rect 1471 4103 1480 4137
rect 1480 4103 1514 4137
rect 1514 4103 1523 4137
rect 1471 4064 1523 4089
rect 1471 4037 1480 4064
rect 1480 4037 1514 4064
rect 1514 4037 1523 4064
rect 1471 3991 1523 4023
rect 1471 3971 1480 3991
rect 1480 3971 1514 3991
rect 1514 3971 1523 3991
rect 1471 3918 1523 3957
rect 1471 3905 1480 3918
rect 1480 3905 1514 3918
rect 1514 3905 1523 3918
rect 1471 3884 1480 3891
rect 1480 3884 1514 3891
rect 1514 3884 1523 3891
rect 1471 3845 1523 3884
rect 1471 3839 1480 3845
rect 1480 3839 1514 3845
rect 1514 3839 1523 3845
rect 1471 3811 1480 3825
rect 1480 3811 1514 3825
rect 1514 3811 1523 3825
rect 1471 3773 1523 3811
rect 1471 3738 1480 3759
rect 1480 3738 1514 3759
rect 1514 3738 1523 3759
rect 1471 3707 1523 3738
rect 1471 3665 1480 3693
rect 1480 3665 1514 3693
rect 1514 3665 1523 3693
rect 1471 3641 1523 3665
rect 1471 3626 1523 3627
rect 1471 3592 1480 3626
rect 1480 3592 1514 3626
rect 1514 3592 1523 3626
rect 1471 3575 1523 3592
rect 1471 3553 1523 3561
rect 1471 3519 1480 3553
rect 1480 3519 1514 3553
rect 1514 3519 1523 3553
rect 1471 3509 1523 3519
rect 240 3378 292 3430
rect 849 3273 901 3325
rect 445 3200 497 3252
rect 509 3200 561 3252
rect 573 3200 625 3252
rect 849 3209 901 3261
rect 240 2973 292 2977
rect 240 2939 249 2973
rect 249 2939 283 2973
rect 283 2939 292 2973
rect 240 2925 292 2939
rect 240 2901 292 2913
rect 240 2867 249 2901
rect 249 2867 283 2901
rect 283 2867 292 2901
rect 240 2861 292 2867
rect 1471 3480 1523 3495
rect 1156 3412 1208 3464
rect 1220 3412 1272 3464
rect 1284 3412 1336 3464
rect 1471 3446 1480 3480
rect 1480 3446 1514 3480
rect 1514 3446 1523 3480
rect 1471 3443 1523 3446
rect 1471 3407 1523 3429
rect 1471 3377 1480 3407
rect 1480 3377 1514 3407
rect 1514 3377 1523 3407
rect 1471 3333 1523 3363
rect 1471 3311 1480 3333
rect 1480 3311 1514 3333
rect 1514 3311 1523 3333
rect 1156 3164 1208 3216
rect 1220 3164 1272 3216
rect 1284 3164 1336 3216
rect 849 2989 901 3041
rect 849 2925 901 2977
rect 1471 3259 1523 3297
rect 1471 3245 1480 3259
rect 1480 3245 1514 3259
rect 1514 3245 1523 3259
rect 1471 3225 1480 3231
rect 1480 3225 1514 3231
rect 1514 3225 1523 3231
rect 1471 3185 1523 3225
rect 1471 3179 1480 3185
rect 1480 3179 1514 3185
rect 1514 3179 1523 3185
rect 1471 3151 1480 3165
rect 1480 3151 1514 3165
rect 1514 3151 1523 3165
rect 1471 3113 1523 3151
rect 1471 3077 1480 3099
rect 1480 3077 1514 3099
rect 1514 3077 1523 3099
rect 1471 3047 1523 3077
rect 1471 3003 1480 3033
rect 1480 3003 1514 3033
rect 1514 3003 1523 3033
rect 1471 2981 1523 3003
rect 1471 2963 1523 2967
rect 958 2919 1010 2925
rect 1471 2929 1480 2963
rect 1480 2929 1514 2963
rect 1514 2929 1523 2963
rect 3020 5163 3072 5172
rect 3020 5129 3026 5163
rect 3026 5129 3068 5163
rect 3068 5129 3072 5163
rect 3590 5140 3642 5192
rect 4124 5244 4176 5252
rect 4124 5210 4138 5244
rect 4138 5210 4176 5244
rect 4124 5200 4176 5210
rect 4188 5200 4240 5252
rect 6780 5231 6832 5283
rect 6844 5231 6896 5283
rect 10267 5247 10319 5299
rect 11859 5278 11911 5330
rect 11926 5278 11978 5330
rect 12407 5278 12459 5330
rect 12474 5278 12526 5330
rect 10267 5183 10319 5235
rect 11455 5193 11507 5245
rect 3020 5120 3072 5129
rect 11455 5126 11507 5178
rect 12234 5175 12286 5227
rect 12301 5175 12353 5227
rect 3070 5057 3079 5079
rect 3079 5057 3113 5079
rect 3113 5057 3122 5079
rect 2032 5003 2084 5055
rect 2096 5003 2148 5055
rect 2160 5003 2212 5055
rect 2224 5003 2276 5055
rect 2288 5003 2340 5055
rect 3070 5027 3122 5057
rect 2572 4973 2624 5025
rect 2636 4973 2688 5025
rect 3070 4981 3079 5012
rect 3079 4981 3113 5012
rect 3113 4981 3122 5012
rect 1946 4900 1998 4952
rect 1946 4816 1998 4868
rect 1946 4733 1998 4785
rect 1946 4650 1998 4702
rect 2032 4547 2084 4599
rect 2096 4547 2148 4599
rect 2160 4547 2212 4599
rect 2224 4547 2276 4599
rect 2288 4547 2340 4599
rect 3070 4960 3122 4981
rect 4098 5027 4150 5079
rect 4098 4963 4150 5015
rect 4258 5058 4310 5108
rect 4258 5056 4266 5058
rect 4266 5056 4300 5058
rect 4300 5056 4310 5058
rect 4258 5024 4266 5026
rect 4266 5024 4300 5026
rect 4300 5024 4310 5026
rect 4258 4974 4310 5024
rect 3070 4939 3122 4945
rect 3070 4905 3079 4939
rect 3079 4905 3113 4939
rect 3113 4905 3122 4939
rect 3070 4893 3122 4905
rect 3070 4863 3122 4878
rect 3070 4829 3079 4863
rect 3079 4829 3113 4863
rect 3113 4829 3122 4863
rect 3070 4826 3122 4829
rect 3070 4787 3122 4811
rect 4258 4920 4266 4944
rect 4266 4920 4300 4944
rect 4300 4920 4310 4944
rect 4258 4892 4310 4920
rect 4258 4850 4310 4862
rect 4258 4816 4266 4850
rect 4266 4816 4300 4850
rect 4300 4816 4310 4850
rect 4258 4810 4310 4816
rect 4637 5066 4689 5118
rect 4637 4997 4689 5049
rect 4637 4928 4689 4980
rect 4637 4859 4689 4911
rect 5034 5120 5086 5124
rect 5100 5120 5152 5124
rect 5166 5120 5218 5124
rect 5232 5120 5284 5124
rect 5298 5120 5350 5124
rect 5364 5120 5416 5124
rect 5430 5120 5482 5124
rect 5496 5120 5548 5124
rect 5562 5120 5614 5124
rect 5034 5086 5057 5120
rect 5057 5086 5086 5120
rect 5100 5086 5129 5120
rect 5129 5086 5152 5120
rect 5166 5086 5201 5120
rect 5201 5086 5218 5120
rect 5232 5086 5235 5120
rect 5235 5086 5273 5120
rect 5273 5086 5284 5120
rect 5298 5086 5307 5120
rect 5307 5086 5345 5120
rect 5345 5086 5350 5120
rect 5364 5086 5379 5120
rect 5379 5086 5416 5120
rect 5430 5086 5451 5120
rect 5451 5086 5482 5120
rect 5496 5086 5523 5120
rect 5523 5086 5548 5120
rect 5562 5086 5595 5120
rect 5595 5086 5614 5120
rect 5034 5072 5086 5086
rect 5100 5072 5152 5086
rect 5166 5072 5218 5086
rect 5232 5072 5284 5086
rect 5298 5072 5350 5086
rect 5364 5072 5416 5086
rect 5430 5072 5482 5086
rect 5496 5072 5548 5086
rect 5562 5072 5614 5086
rect 5628 5120 5680 5124
rect 5628 5086 5633 5120
rect 5633 5086 5667 5120
rect 5667 5086 5680 5120
rect 5628 5072 5680 5086
rect 5694 5120 5746 5124
rect 5694 5086 5705 5120
rect 5705 5086 5739 5120
rect 5739 5086 5746 5120
rect 5694 5072 5746 5086
rect 5760 5120 5812 5124
rect 5760 5086 5777 5120
rect 5777 5086 5811 5120
rect 5811 5086 5812 5120
rect 5760 5072 5812 5086
rect 5826 5120 5878 5124
rect 5892 5120 5944 5124
rect 5959 5120 6011 5124
rect 6142 5120 6194 5124
rect 5826 5086 5849 5120
rect 5849 5086 5878 5120
rect 5892 5086 5921 5120
rect 5921 5086 5944 5120
rect 5959 5086 5993 5120
rect 5993 5086 6011 5120
rect 6142 5086 6171 5120
rect 6171 5086 6194 5120
rect 5826 5072 5878 5086
rect 5892 5072 5944 5086
rect 5959 5072 6011 5086
rect 6142 5072 6194 5086
rect 6206 5120 6258 5124
rect 6206 5086 6209 5120
rect 6209 5086 6243 5120
rect 6243 5086 6258 5120
rect 6206 5072 6258 5086
rect 6270 5120 6322 5124
rect 6270 5086 6281 5120
rect 6281 5086 6315 5120
rect 6315 5086 6322 5120
rect 6270 5072 6322 5086
rect 6334 5120 6386 5124
rect 6399 5120 6451 5124
rect 6464 5120 6516 5124
rect 6529 5120 6581 5124
rect 6594 5120 6646 5124
rect 6969 5120 7021 5124
rect 7045 5120 7097 5124
rect 7121 5120 7173 5124
rect 7197 5120 7249 5124
rect 7273 5120 7325 5124
rect 7393 5120 7445 5124
rect 7461 5120 7513 5124
rect 7529 5120 7581 5124
rect 7598 5120 7650 5124
rect 7667 5120 7719 5124
rect 7736 5120 7788 5124
rect 6334 5086 6353 5120
rect 6353 5086 6386 5120
rect 6399 5086 6425 5120
rect 6425 5086 6451 5120
rect 6464 5086 6497 5120
rect 6497 5086 6516 5120
rect 6529 5086 6531 5120
rect 6531 5086 6569 5120
rect 6569 5086 6581 5120
rect 6594 5086 6603 5120
rect 6603 5086 6641 5120
rect 6641 5086 6646 5120
rect 6969 5086 7004 5120
rect 7004 5086 7021 5120
rect 7045 5086 7077 5120
rect 7077 5086 7097 5120
rect 7121 5086 7150 5120
rect 7150 5086 7173 5120
rect 7197 5086 7223 5120
rect 7223 5086 7249 5120
rect 7273 5086 7296 5120
rect 7296 5086 7325 5120
rect 7393 5086 7403 5120
rect 7403 5086 7442 5120
rect 7442 5086 7445 5120
rect 7461 5086 7476 5120
rect 7476 5086 7513 5120
rect 7529 5086 7549 5120
rect 7549 5086 7581 5120
rect 7598 5086 7622 5120
rect 7622 5086 7650 5120
rect 7667 5086 7695 5120
rect 7695 5086 7719 5120
rect 7736 5086 7768 5120
rect 7768 5086 7788 5120
rect 6334 5072 6386 5086
rect 6399 5072 6451 5086
rect 6464 5072 6516 5086
rect 6529 5072 6581 5086
rect 6594 5072 6646 5086
rect 6969 5072 7021 5086
rect 7045 5072 7097 5086
rect 7121 5072 7173 5086
rect 7197 5072 7249 5086
rect 7273 5072 7325 5086
rect 7393 5072 7445 5086
rect 7461 5072 7513 5086
rect 7529 5072 7581 5086
rect 7598 5072 7650 5086
rect 7667 5072 7719 5086
rect 7736 5072 7788 5086
rect 7805 5120 7857 5124
rect 7805 5086 7807 5120
rect 7807 5086 7841 5120
rect 7841 5086 7857 5120
rect 7805 5072 7857 5086
rect 7874 5120 7926 5124
rect 7874 5086 7880 5120
rect 7880 5086 7914 5120
rect 7914 5086 7926 5120
rect 7874 5072 7926 5086
rect 7943 5120 7995 5124
rect 7943 5086 7953 5120
rect 7953 5086 7987 5120
rect 7987 5086 7995 5120
rect 7943 5072 7995 5086
rect 8012 5120 8064 5124
rect 8187 5120 8239 5124
rect 8255 5120 8307 5124
rect 8323 5120 8375 5124
rect 8012 5086 8026 5120
rect 8026 5086 8060 5120
rect 8060 5086 8064 5120
rect 8187 5086 8206 5120
rect 8206 5086 8239 5120
rect 8255 5086 8279 5120
rect 8279 5086 8307 5120
rect 8323 5086 8352 5120
rect 8352 5086 8375 5120
rect 8012 5072 8064 5086
rect 8187 5072 8239 5086
rect 8255 5072 8307 5086
rect 8323 5072 8375 5086
rect 8391 5120 8443 5124
rect 8391 5086 8425 5120
rect 8425 5086 8443 5120
rect 8391 5072 8443 5086
rect 8459 5120 8511 5124
rect 8459 5086 8464 5120
rect 8464 5086 8498 5120
rect 8498 5086 8511 5120
rect 8459 5072 8511 5086
rect 8528 5120 8580 5124
rect 8528 5086 8537 5120
rect 8537 5086 8571 5120
rect 8571 5086 8580 5120
rect 8528 5072 8580 5086
rect 8597 5120 8649 5124
rect 8597 5086 8610 5120
rect 8610 5086 8644 5120
rect 8644 5086 8649 5120
rect 8597 5072 8649 5086
rect 8666 5120 8718 5124
rect 8666 5086 8683 5120
rect 8683 5086 8717 5120
rect 8717 5086 8718 5120
rect 8666 5072 8718 5086
rect 8735 5120 8787 5124
rect 8804 5120 8856 5124
rect 8873 5120 8925 5124
rect 8942 5120 8994 5124
rect 9011 5120 9063 5124
rect 9080 5120 9132 5124
rect 8735 5086 8756 5120
rect 8756 5086 8787 5120
rect 8804 5086 8829 5120
rect 8829 5086 8856 5120
rect 8873 5086 8902 5120
rect 8902 5086 8925 5120
rect 8942 5086 8975 5120
rect 8975 5086 8994 5120
rect 9011 5086 9048 5120
rect 9048 5086 9063 5120
rect 9080 5086 9082 5120
rect 9082 5086 9121 5120
rect 9121 5086 9132 5120
rect 9554 5117 9606 5126
rect 9622 5117 9674 5126
rect 9690 5117 9742 5126
rect 9759 5117 9811 5126
rect 9828 5117 9880 5126
rect 9897 5117 9949 5126
rect 9966 5117 10018 5126
rect 10490 5117 10542 5126
rect 10554 5117 10606 5126
rect 10618 5117 10670 5126
rect 8735 5072 8787 5086
rect 8804 5072 8856 5086
rect 8873 5072 8925 5086
rect 8942 5072 8994 5086
rect 9011 5072 9063 5086
rect 9080 5072 9132 5086
rect 9459 5083 9506 5103
rect 9506 5083 9511 5103
rect 9554 5083 9580 5117
rect 9580 5083 9606 5117
rect 9622 5083 9654 5117
rect 9654 5083 9674 5117
rect 9690 5083 9728 5117
rect 9728 5083 9742 5117
rect 9759 5083 9762 5117
rect 9762 5083 9802 5117
rect 9802 5083 9811 5117
rect 9828 5083 9836 5117
rect 9836 5083 9876 5117
rect 9876 5083 9880 5117
rect 9897 5083 9910 5117
rect 9910 5083 9949 5117
rect 9966 5083 9984 5117
rect 9984 5083 10018 5117
rect 10490 5083 10502 5117
rect 10502 5083 10542 5117
rect 10554 5083 10576 5117
rect 10576 5083 10606 5117
rect 10618 5083 10650 5117
rect 10650 5083 10670 5117
rect 4840 5024 4892 5066
rect 9459 5051 9511 5083
rect 9554 5074 9606 5083
rect 9622 5074 9674 5083
rect 9690 5074 9742 5083
rect 9759 5074 9811 5083
rect 9828 5074 9880 5083
rect 9897 5074 9949 5083
rect 9966 5074 10018 5083
rect 10490 5074 10542 5083
rect 10554 5074 10606 5083
rect 10618 5074 10670 5083
rect 10682 5117 10734 5126
rect 10682 5083 10690 5117
rect 10690 5083 10724 5117
rect 10724 5083 10734 5117
rect 10682 5074 10734 5083
rect 10747 5117 10799 5126
rect 10747 5083 10764 5117
rect 10764 5083 10798 5117
rect 10798 5083 10799 5117
rect 10747 5074 10799 5083
rect 10812 5117 10864 5126
rect 10877 5117 10929 5126
rect 10942 5117 10994 5126
rect 11007 5117 11059 5126
rect 11207 5117 11259 5126
rect 10812 5083 10838 5117
rect 10838 5083 10864 5117
rect 10877 5083 10912 5117
rect 10912 5083 10929 5117
rect 10942 5083 10946 5117
rect 10946 5083 10986 5117
rect 10986 5083 10994 5117
rect 11007 5083 11020 5117
rect 11020 5083 11059 5117
rect 11207 5083 11241 5117
rect 11241 5083 11259 5117
rect 10812 5074 10864 5083
rect 10877 5074 10929 5083
rect 10942 5074 10994 5083
rect 11007 5074 11059 5083
rect 11207 5074 11259 5083
rect 11274 5117 11326 5126
rect 11274 5083 11280 5117
rect 11280 5083 11314 5117
rect 11314 5083 11326 5117
rect 11274 5074 11326 5083
rect 11341 5117 11393 5126
rect 11341 5083 11353 5117
rect 11353 5083 11387 5117
rect 11387 5083 11393 5117
rect 11341 5074 11393 5083
rect 11603 5117 11655 5126
rect 11603 5083 11609 5117
rect 11609 5083 11643 5117
rect 11643 5083 11655 5117
rect 11603 5074 11655 5083
rect 11670 5117 11722 5126
rect 11670 5083 11683 5117
rect 11683 5083 11717 5117
rect 11717 5083 11722 5117
rect 11670 5074 11722 5083
rect 11737 5117 11789 5126
rect 11965 5117 12017 5126
rect 11737 5083 11757 5117
rect 11757 5083 11789 5117
rect 11965 5083 11982 5117
rect 11982 5083 12016 5117
rect 12016 5083 12017 5117
rect 11737 5074 11789 5083
rect 11965 5074 12017 5083
rect 12029 5117 12081 5126
rect 12093 5117 12145 5126
rect 12157 5117 12209 5126
rect 12221 5117 12273 5126
rect 12399 5117 12451 5126
rect 12495 5117 12547 5126
rect 12029 5083 12057 5117
rect 12057 5083 12081 5117
rect 12093 5083 12132 5117
rect 12132 5083 12145 5117
rect 12157 5083 12166 5117
rect 12166 5083 12207 5117
rect 12207 5083 12209 5117
rect 12221 5083 12241 5117
rect 12241 5083 12273 5117
rect 12399 5083 12432 5117
rect 12432 5083 12451 5117
rect 12495 5083 12507 5117
rect 12507 5083 12541 5117
rect 12541 5083 12547 5117
rect 12029 5074 12081 5083
rect 12093 5074 12145 5083
rect 12157 5074 12209 5083
rect 12221 5074 12273 5083
rect 12399 5074 12451 5083
rect 12495 5074 12547 5083
rect 4840 5014 4869 5024
rect 4869 5014 4892 5024
rect 4840 4952 4892 4964
rect 4840 4918 4869 4952
rect 4869 4918 4892 4952
rect 4840 4912 4892 4918
rect 9459 5005 9511 5038
rect 9459 4986 9468 5005
rect 9468 4986 9502 5005
rect 9502 4986 9511 5005
rect 9459 4971 9468 4973
rect 9468 4971 9502 4973
rect 9502 4971 9511 4973
rect 9459 4932 9511 4971
rect 9459 4921 9468 4932
rect 9468 4921 9502 4932
rect 9502 4921 9511 4932
rect 9459 4898 9468 4908
rect 9468 4898 9502 4908
rect 9502 4898 9511 4908
rect 4637 4790 4689 4842
rect 3070 4759 3079 4787
rect 3079 4759 3113 4787
rect 3113 4759 3122 4787
rect 3070 4711 3122 4744
rect 3884 4738 3936 4790
rect 3948 4738 4000 4790
rect 4012 4738 4064 4790
rect 4637 4721 4689 4773
rect 4749 4812 4801 4864
rect 9459 4859 9511 4898
rect 9459 4856 9468 4859
rect 9468 4856 9502 4859
rect 9502 4856 9511 4859
rect 9459 4825 9468 4843
rect 9468 4825 9502 4843
rect 9502 4825 9511 4843
rect 9459 4791 9511 4825
rect 4749 4727 4801 4779
rect 3070 4692 3079 4711
rect 3079 4692 3113 4711
rect 3113 4692 3122 4711
rect 3070 4635 3122 4677
rect 4749 4641 4801 4693
rect 4840 4771 4892 4777
rect 4840 4737 4869 4771
rect 4869 4737 4892 4771
rect 4840 4725 4892 4737
rect 4840 4690 4892 4708
rect 4840 4656 4869 4690
rect 4869 4656 4892 4690
rect 3070 4625 3079 4635
rect 3079 4625 3113 4635
rect 3113 4625 3122 4635
rect 4840 4610 4892 4639
rect 3070 4601 3079 4610
rect 3079 4601 3113 4610
rect 3113 4601 3122 4610
rect 2572 4517 2624 4569
rect 2636 4517 2688 4569
rect 3070 4559 3122 4601
rect 3070 4558 3079 4559
rect 3079 4558 3113 4559
rect 3113 4558 3122 4559
rect 3070 4525 3079 4543
rect 3079 4525 3113 4543
rect 3113 4525 3122 4543
rect 4565 4561 4574 4586
rect 4574 4561 4608 4586
rect 4608 4561 4617 4586
rect 4565 4534 4617 4561
rect 4637 4561 4646 4586
rect 4646 4561 4680 4586
rect 4680 4561 4689 4586
rect 4637 4534 4689 4561
rect 4840 4587 4869 4610
rect 4869 4587 4892 4610
rect 4840 4530 4892 4570
rect 3070 4491 3122 4525
rect 3070 4448 3079 4476
rect 3079 4448 3113 4476
rect 3113 4448 3122 4476
rect 4840 4518 4869 4530
rect 4869 4518 4892 4530
rect 4840 4496 4869 4501
rect 4869 4496 4892 4501
rect 3070 4424 3122 4448
rect 2830 4352 2882 4404
rect 2830 4288 2882 4340
rect 3070 4405 3122 4408
rect 3070 4371 3079 4405
rect 3079 4371 3113 4405
rect 3113 4371 3122 4405
rect 3070 4356 3122 4371
rect 3070 4328 3122 4340
rect 3070 4294 3079 4328
rect 3079 4294 3113 4328
rect 3113 4294 3122 4328
rect 4840 4450 4892 4496
rect 4840 4449 4869 4450
rect 4869 4449 4892 4450
rect 4840 4416 4869 4432
rect 4869 4416 4892 4432
rect 3070 4288 3122 4294
rect 3884 4337 3936 4389
rect 3948 4337 4000 4389
rect 4012 4337 4064 4389
rect 4637 4402 4689 4408
rect 4637 4368 4646 4402
rect 4646 4368 4680 4402
rect 4680 4368 4689 4402
rect 4637 4356 4689 4368
rect 2032 4091 2084 4143
rect 2096 4091 2148 4143
rect 2160 4091 2212 4143
rect 2224 4091 2276 4143
rect 2288 4091 2340 4143
rect 2830 4081 2882 4133
rect 2830 4017 2882 4069
rect 3070 4168 3122 4174
rect 3070 4134 3079 4168
rect 3079 4134 3113 4168
rect 3113 4134 3122 4168
rect 4258 4330 4310 4336
rect 4258 4296 4266 4330
rect 4266 4296 4300 4330
rect 4300 4296 4310 4330
rect 4258 4284 4310 4296
rect 4258 4222 4310 4234
rect 4258 4188 4266 4222
rect 4266 4188 4300 4222
rect 4300 4188 4310 4222
rect 4258 4182 4310 4188
rect 4637 4299 4689 4342
rect 4637 4290 4646 4299
rect 4646 4290 4680 4299
rect 4680 4290 4689 4299
rect 4637 4265 4646 4275
rect 4646 4265 4680 4275
rect 4680 4265 4689 4275
rect 4637 4223 4689 4265
rect 4637 4196 4689 4208
rect 4637 4162 4646 4196
rect 4646 4162 4680 4196
rect 4680 4162 4689 4196
rect 4840 4380 4892 4416
rect 9459 4752 9468 4778
rect 9468 4752 9502 4778
rect 9502 4752 9511 4778
rect 9459 4726 9511 4752
rect 9459 4679 9468 4713
rect 9468 4679 9502 4713
rect 9502 4679 9511 4713
rect 9459 4661 9511 4679
rect 9459 4640 9511 4648
rect 9459 4606 9468 4640
rect 9468 4606 9502 4640
rect 9502 4606 9511 4640
rect 9459 4596 9511 4606
rect 9459 4567 9511 4583
rect 9459 4533 9468 4567
rect 9468 4533 9502 4567
rect 9502 4533 9511 4567
rect 9459 4531 9511 4533
rect 9459 4494 9511 4518
rect 9459 4466 9468 4494
rect 9468 4466 9502 4494
rect 9502 4466 9511 4494
rect 9459 4421 9511 4453
rect 9459 4401 9468 4421
rect 9468 4401 9502 4421
rect 9502 4401 9511 4421
rect 9459 4387 9468 4388
rect 9468 4387 9502 4388
rect 9502 4387 9511 4388
rect 4840 4336 4869 4362
rect 4869 4336 4892 4362
rect 4840 4310 4892 4336
rect 6780 4321 6832 4373
rect 6844 4321 6896 4373
rect 9459 4348 9511 4387
rect 9459 4336 9468 4348
rect 9468 4336 9502 4348
rect 9502 4336 9511 4348
rect 4840 4290 4892 4292
rect 4840 4256 4869 4290
rect 4869 4256 4892 4290
rect 4840 4240 4892 4256
rect 4840 4210 4892 4222
rect 4840 4176 4869 4210
rect 4869 4176 4892 4210
rect 4840 4170 4892 4176
rect 9459 4314 9468 4323
rect 9468 4314 9502 4323
rect 9502 4314 9511 4323
rect 9459 4275 9511 4314
rect 9459 4271 9468 4275
rect 9468 4271 9502 4275
rect 9502 4271 9511 4275
rect 9459 4241 9468 4258
rect 9468 4241 9502 4258
rect 9502 4241 9511 4258
rect 9459 4206 9511 4241
rect 9459 4168 9468 4193
rect 9468 4168 9502 4193
rect 9502 4168 9511 4193
rect 4637 4156 4689 4162
rect 3070 4122 3122 4134
rect 3070 4092 3122 4100
rect 3070 4058 3079 4092
rect 3079 4058 3113 4092
rect 3113 4058 3122 4092
rect 9459 4141 9511 4168
rect 3070 4048 3122 4058
rect 3070 4017 3122 4027
rect 3884 4021 3936 4073
rect 3948 4021 4000 4073
rect 4012 4021 4064 4073
rect 4178 4064 4230 4116
rect 9459 4094 9468 4128
rect 9468 4094 9502 4128
rect 9502 4094 9511 4128
rect 9459 4076 9511 4094
rect 3070 3983 3079 4017
rect 3079 3983 3113 4017
rect 3113 3983 3122 4017
rect 4178 4000 4230 4052
rect 9459 4054 9511 4063
rect 4637 4024 4689 4030
rect 3070 3975 3122 3983
rect 3070 3942 3122 3954
rect 3070 3908 3079 3942
rect 3079 3908 3113 3942
rect 3113 3908 3122 3942
rect 4637 3990 4646 4024
rect 4646 3990 4680 4024
rect 4680 3990 4689 4024
rect 9459 4020 9468 4054
rect 9468 4020 9502 4054
rect 9502 4020 9511 4054
rect 9459 4011 9511 4020
rect 4637 3978 4689 3990
rect 4637 3944 4689 3963
rect 3070 3902 3122 3908
rect 4098 3871 4150 3923
rect 4637 3911 4646 3944
rect 4646 3911 4680 3944
rect 4680 3911 4689 3944
rect 4637 3864 4689 3896
rect 4637 3844 4646 3864
rect 4646 3844 4680 3864
rect 4680 3844 4689 3864
rect 2830 3728 2882 3780
rect 4418 3779 4470 3831
rect 2032 3635 2084 3687
rect 2096 3635 2148 3687
rect 2160 3635 2212 3687
rect 2224 3635 2276 3687
rect 2288 3635 2340 3687
rect 2830 3664 2882 3716
rect 3070 3743 3122 3749
rect 3070 3709 3079 3743
rect 3079 3709 3113 3743
rect 3113 3709 3122 3743
rect 3884 3711 3936 3763
rect 3948 3711 4000 3763
rect 4012 3711 4064 3763
rect 4258 3743 4310 3749
rect 3070 3697 3122 3709
rect 2910 3601 2962 3653
rect 2910 3537 2962 3589
rect 3070 3645 3122 3654
rect 3070 3611 3079 3645
rect 3079 3611 3113 3645
rect 3113 3611 3122 3645
rect 4258 3709 4266 3743
rect 4266 3709 4300 3743
rect 4300 3709 4310 3743
rect 4418 3715 4470 3767
rect 4637 3785 4689 3829
rect 4637 3777 4646 3785
rect 4646 3777 4680 3785
rect 4680 3777 4689 3785
rect 4637 3751 4646 3762
rect 4646 3751 4680 3762
rect 4680 3751 4689 3762
rect 4637 3710 4689 3751
rect 4749 3938 4801 3990
rect 9459 3980 9511 3998
rect 9459 3946 9468 3980
rect 9468 3946 9502 3980
rect 9502 3946 9511 3980
rect 4749 3872 4801 3924
rect 4749 3806 4801 3858
rect 4749 3739 4801 3791
rect 9459 3906 9511 3933
rect 9459 3881 9468 3906
rect 9468 3881 9502 3906
rect 9502 3881 9511 3906
rect 9459 3832 9511 3868
rect 9459 3816 9468 3832
rect 9468 3816 9502 3832
rect 9502 3816 9511 3832
rect 9459 3798 9468 3804
rect 9468 3798 9502 3804
rect 9502 3798 9511 3804
rect 9459 3758 9511 3798
rect 9459 3752 9468 3758
rect 9468 3752 9502 3758
rect 9502 3752 9511 3758
rect 5163 3746 5215 3747
rect 5230 3746 5282 3747
rect 5297 3746 5349 3747
rect 5364 3746 5416 3747
rect 5431 3746 5483 3747
rect 5498 3746 5550 3747
rect 5565 3746 5617 3747
rect 5632 3746 5684 3747
rect 5699 3746 5751 3747
rect 5766 3746 5818 3747
rect 5834 3746 5886 3747
rect 5902 3746 5954 3747
rect 5970 3746 6022 3747
rect 6142 3746 6706 3747
rect 6719 3746 6771 3747
rect 6784 3746 6836 3747
rect 6849 3746 6901 3747
rect 7393 3746 7445 3752
rect 7461 3746 7513 3752
rect 7529 3746 7581 3752
rect 7598 3746 7650 3752
rect 7667 3746 7719 3752
rect 7736 3746 7788 3752
rect 7805 3746 7857 3752
rect 7874 3746 7926 3752
rect 7943 3746 7995 3752
rect 8012 3746 8064 3752
rect 8187 3746 8239 3752
rect 8255 3746 8307 3752
rect 8323 3746 8375 3752
rect 8391 3746 8443 3752
rect 8459 3746 8511 3752
rect 8528 3746 8580 3752
rect 8597 3746 8649 3752
rect 8666 3746 8718 3752
rect 8735 3746 8787 3752
rect 8804 3746 8856 3752
rect 8873 3746 8925 3752
rect 8942 3746 8994 3752
rect 9011 3746 9063 3752
rect 4258 3697 4310 3709
rect 4258 3645 4310 3654
rect 3070 3602 3122 3611
rect 3070 3548 3122 3560
rect 4098 3586 4150 3638
rect 2830 3457 2882 3509
rect 3070 3514 3079 3548
rect 3079 3514 3113 3548
rect 3113 3514 3122 3548
rect 4098 3522 4150 3574
rect 4258 3611 4266 3645
rect 4266 3611 4300 3645
rect 4300 3611 4310 3645
rect 4258 3602 4310 3611
rect 4258 3548 4310 3560
rect 3070 3508 3122 3514
rect 4258 3514 4266 3548
rect 4266 3514 4300 3548
rect 4300 3514 4310 3548
rect 4258 3508 4310 3514
rect 4637 3672 4646 3695
rect 4646 3672 4680 3695
rect 4680 3672 4689 3695
rect 4637 3643 4689 3672
rect 5163 3695 5215 3746
rect 5230 3695 5282 3746
rect 5297 3695 5349 3746
rect 5364 3695 5416 3746
rect 5431 3695 5483 3746
rect 5498 3695 5550 3746
rect 5565 3695 5617 3746
rect 5632 3695 5684 3746
rect 5699 3695 5751 3746
rect 5766 3695 5818 3746
rect 5834 3695 5886 3746
rect 5902 3695 5954 3746
rect 5970 3695 6022 3746
rect 5163 3640 5215 3683
rect 5230 3640 5282 3683
rect 5297 3640 5349 3683
rect 5364 3640 5416 3683
rect 5431 3640 5483 3683
rect 5498 3640 5550 3683
rect 5565 3640 5617 3683
rect 5632 3640 5684 3683
rect 5699 3640 5751 3683
rect 5766 3640 5818 3683
rect 5834 3640 5886 3683
rect 5902 3640 5954 3683
rect 5970 3640 6022 3683
rect 6142 3640 6706 3746
rect 6719 3695 6771 3746
rect 6784 3695 6836 3746
rect 6849 3695 6901 3746
rect 7393 3700 7445 3746
rect 7461 3700 7513 3746
rect 7529 3700 7581 3746
rect 7598 3700 7650 3746
rect 7667 3700 7719 3746
rect 7736 3700 7788 3746
rect 7805 3700 7857 3746
rect 7874 3700 7926 3746
rect 7943 3700 7995 3746
rect 8012 3700 8064 3746
rect 8187 3700 8239 3746
rect 8255 3700 8307 3746
rect 8323 3700 8375 3746
rect 8391 3700 8443 3746
rect 8459 3700 8511 3746
rect 8528 3700 8580 3746
rect 8597 3700 8649 3746
rect 8666 3700 8718 3746
rect 8735 3700 8787 3746
rect 8804 3700 8856 3746
rect 8873 3700 8925 3746
rect 8942 3700 8971 3746
rect 8971 3700 8994 3746
rect 9011 3712 9044 3746
rect 9044 3712 9063 3746
rect 9011 3700 9063 3712
rect 9080 3746 9132 3752
rect 9080 3712 9083 3746
rect 9083 3712 9117 3746
rect 9117 3712 9132 3746
rect 9459 3724 9468 3740
rect 9468 3724 9502 3740
rect 9502 3724 9511 3740
rect 9080 3700 9132 3712
rect 9459 3688 9511 3724
rect 6719 3640 6771 3683
rect 6784 3640 6836 3683
rect 6849 3640 6901 3683
rect 7393 3640 7445 3688
rect 7461 3640 7513 3688
rect 7529 3640 7581 3688
rect 7598 3640 7650 3688
rect 7667 3640 7719 3688
rect 7736 3640 7788 3688
rect 7805 3640 7857 3688
rect 7874 3640 7926 3688
rect 7943 3640 7995 3688
rect 8012 3640 8064 3688
rect 8187 3640 8239 3688
rect 8255 3640 8307 3688
rect 8323 3640 8375 3688
rect 8391 3640 8443 3688
rect 8459 3640 8511 3688
rect 8528 3640 8580 3688
rect 8597 3640 8649 3688
rect 8666 3640 8718 3688
rect 8735 3640 8787 3688
rect 8804 3640 8856 3688
rect 8873 3640 8925 3688
rect 8942 3640 8971 3688
rect 8971 3640 8994 3688
rect 9011 3674 9063 3688
rect 9011 3640 9044 3674
rect 9044 3640 9063 3674
rect 4637 3627 4689 3628
rect 4637 3593 4646 3627
rect 4646 3593 4680 3627
rect 4680 3593 4689 3627
rect 4637 3576 4689 3593
rect 5163 3631 5215 3640
rect 5230 3631 5282 3640
rect 5297 3631 5349 3640
rect 5364 3631 5416 3640
rect 5431 3631 5483 3640
rect 5498 3631 5550 3640
rect 5565 3631 5617 3640
rect 5632 3631 5684 3640
rect 5699 3631 5751 3640
rect 5766 3631 5818 3640
rect 5834 3631 5886 3640
rect 5902 3631 5954 3640
rect 5970 3631 6022 3640
rect 6142 3631 6706 3640
rect 6719 3631 6771 3640
rect 6784 3631 6836 3640
rect 6849 3631 6901 3640
rect 7393 3636 7445 3640
rect 7461 3636 7513 3640
rect 7529 3636 7581 3640
rect 7598 3636 7650 3640
rect 7667 3636 7719 3640
rect 7736 3636 7788 3640
rect 7805 3636 7857 3640
rect 7874 3636 7926 3640
rect 7943 3636 7995 3640
rect 8012 3636 8064 3640
rect 8187 3636 8239 3640
rect 8255 3636 8307 3640
rect 8323 3636 8375 3640
rect 8391 3636 8443 3640
rect 8459 3636 8511 3640
rect 8528 3636 8580 3640
rect 8597 3636 8649 3640
rect 8666 3636 8718 3640
rect 8735 3636 8787 3640
rect 8804 3636 8856 3640
rect 8873 3636 8925 3640
rect 8942 3636 8994 3640
rect 9011 3636 9063 3640
rect 9080 3674 9132 3688
rect 9080 3640 9083 3674
rect 9083 3640 9117 3674
rect 9117 3640 9132 3674
rect 9459 3650 9468 3676
rect 9468 3650 9502 3676
rect 9502 3650 9511 3676
rect 9080 3636 9132 3640
rect 9459 3624 9511 3650
rect 9459 3610 9511 3612
rect 4637 3548 4689 3560
rect 9459 3576 9468 3610
rect 9468 3576 9502 3610
rect 9502 3576 9511 3610
rect 9459 3560 9511 3576
rect 4637 3514 4646 3548
rect 4646 3514 4680 3548
rect 4680 3514 4689 3548
rect 4637 3508 4689 3514
rect 6911 3496 6963 3548
rect 6975 3496 7027 3548
rect 7209 3496 7261 3548
rect 7273 3496 7325 3548
rect 9459 3536 9511 3548
rect 9459 3502 9468 3536
rect 9468 3502 9502 3536
rect 9502 3502 9511 3536
rect 9459 3496 9511 3502
rect 10143 4914 10195 4966
rect 2830 3393 2882 3445
rect 3070 3388 3122 3394
rect 2910 3301 2962 3353
rect 2032 3179 2084 3231
rect 2096 3179 2148 3231
rect 2160 3179 2212 3231
rect 2224 3179 2276 3231
rect 2288 3179 2340 3231
rect 2910 3237 2962 3289
rect 3070 3354 3079 3388
rect 3079 3354 3113 3388
rect 3113 3354 3122 3388
rect 4637 3388 4689 3394
rect 3070 3342 3122 3354
rect 3070 3302 3122 3323
rect 3070 3271 3079 3302
rect 3079 3271 3113 3302
rect 3113 3271 3122 3302
rect 3070 3216 3122 3253
rect 3884 3307 3936 3359
rect 3948 3307 4000 3359
rect 4012 3307 4064 3359
rect 4637 3354 4646 3388
rect 4646 3354 4680 3388
rect 4680 3354 4689 3388
rect 4637 3342 4689 3354
rect 4637 3309 4689 3318
rect 4258 3273 4310 3279
rect 4258 3239 4266 3273
rect 4266 3239 4300 3273
rect 4300 3239 4310 3273
rect 2475 3077 2527 3129
rect 2830 3145 2882 3197
rect 2830 3081 2882 3133
rect 3070 3201 3079 3216
rect 3079 3201 3113 3216
rect 3113 3201 3122 3216
rect 3070 3182 3079 3183
rect 3079 3182 3113 3183
rect 3113 3182 3122 3183
rect 3070 3131 3122 3182
rect 4258 3227 4310 3239
rect 4637 3275 4646 3309
rect 4646 3275 4680 3309
rect 4680 3275 4689 3309
rect 4637 3266 4689 3275
rect 4258 3200 4310 3211
rect 4258 3166 4266 3200
rect 4266 3166 4300 3200
rect 4300 3166 4310 3200
rect 4258 3159 4310 3166
rect 3070 3097 3079 3113
rect 3079 3097 3113 3113
rect 3113 3097 3122 3113
rect 3884 3103 3936 3155
rect 3948 3103 4000 3155
rect 4012 3103 4064 3155
rect 4258 3127 4310 3143
rect 2475 3013 2527 3065
rect 3070 3061 3122 3097
rect 3070 3012 3079 3043
rect 3079 3012 3113 3043
rect 3113 3012 3122 3043
rect 2475 2949 2527 3001
rect 3070 2991 3122 3012
rect 429 2857 481 2866
rect 429 2823 441 2857
rect 441 2823 475 2857
rect 475 2823 481 2857
rect 429 2814 481 2823
rect 493 2857 545 2866
rect 493 2823 513 2857
rect 513 2823 545 2857
rect 493 2814 545 2823
rect 958 2885 967 2919
rect 967 2885 1001 2919
rect 1001 2885 1010 2919
rect 958 2873 1010 2885
rect 1156 2870 1208 2922
rect 1220 2870 1272 2922
rect 1284 2870 1336 2922
rect 1471 2915 1523 2929
rect 2910 2907 2962 2959
rect 3070 2961 3122 2973
rect 1471 2889 1523 2901
rect 1471 2855 1480 2889
rect 1480 2855 1514 2889
rect 1514 2855 1523 2889
rect 1471 2849 1523 2855
rect 2475 2838 2527 2844
rect 2475 2804 2484 2838
rect 2484 2804 2518 2838
rect 2518 2804 2527 2838
rect 2475 2792 2527 2804
rect 2750 2792 2802 2844
rect 2910 2843 2962 2895
rect 2990 2888 3042 2940
rect 3070 2927 3079 2961
rect 3079 2927 3113 2961
rect 3113 2927 3122 2961
rect 3070 2921 3122 2927
rect 3590 2966 3642 3018
rect 4178 3040 4230 3092
rect 4178 2976 4230 3028
rect 4258 3093 4266 3127
rect 4266 3093 4300 3127
rect 4300 3093 4310 3127
rect 4418 3180 4470 3232
rect 4637 3230 4689 3242
rect 4637 3196 4646 3230
rect 4646 3196 4680 3230
rect 4680 3196 4689 3230
rect 4637 3190 4689 3196
rect 9732 4764 9784 4816
rect 9732 4700 9784 4752
rect 9459 3350 9511 3356
rect 4418 3116 4470 3168
rect 4840 3333 4892 3339
rect 4840 3299 4869 3333
rect 4869 3299 4892 3333
rect 9459 3316 9468 3350
rect 9468 3316 9502 3350
rect 9502 3316 9511 3350
rect 4840 3287 4892 3299
rect 4840 3255 4892 3274
rect 6164 3260 6216 3312
rect 6241 3260 6293 3312
rect 6318 3260 6370 3312
rect 6395 3260 6447 3312
rect 6471 3260 6523 3312
rect 7400 3262 7452 3314
rect 7467 3262 7519 3314
rect 7534 3262 7586 3314
rect 7601 3262 7653 3314
rect 7668 3262 7720 3314
rect 7735 3262 7787 3314
rect 7802 3262 7854 3314
rect 7869 3262 7921 3314
rect 7936 3262 7988 3314
rect 8002 3262 8054 3314
rect 9459 3304 9511 3316
rect 9459 3261 9511 3272
rect 4840 3222 4869 3255
rect 4869 3222 4892 3255
rect 9459 3227 9468 3261
rect 9468 3227 9502 3261
rect 9502 3227 9511 3261
rect 9459 3220 9511 3227
rect 4840 3177 4892 3209
rect 4840 3157 4869 3177
rect 4869 3157 4892 3177
rect 4840 3143 4869 3144
rect 4869 3143 4892 3144
rect 4258 3091 4310 3093
rect 4840 3099 4892 3143
rect 5383 3136 5435 3188
rect 5447 3136 5499 3188
rect 8638 3137 8690 3189
rect 8702 3137 8754 3189
rect 10143 4850 10195 4902
rect 9928 4458 9980 4510
rect 9928 4394 9980 4446
rect 9848 3373 9900 3407
rect 9848 3355 9859 3373
rect 9859 3355 9893 3373
rect 9893 3355 9900 3373
rect 9848 3299 9900 3329
rect 9848 3277 9859 3299
rect 9859 3277 9893 3299
rect 9893 3277 9900 3299
rect 9848 3225 9900 3250
rect 9848 3198 9859 3225
rect 9859 3198 9893 3225
rect 9893 3198 9900 3225
rect 4258 3054 4310 3075
rect 4258 3023 4266 3054
rect 4266 3023 4300 3054
rect 4300 3023 4310 3054
rect 4258 2981 4310 3008
rect 3590 2898 3642 2950
rect 3884 2950 3936 2959
rect 3884 2916 3894 2950
rect 3894 2916 3928 2950
rect 3928 2916 3936 2950
rect 3884 2907 3936 2916
rect 3948 2950 4000 2959
rect 3948 2916 3966 2950
rect 3966 2916 4000 2950
rect 3948 2907 4000 2916
rect 4012 2907 4064 2959
rect 4258 2956 4266 2981
rect 4266 2956 4300 2981
rect 4300 2956 4310 2981
rect 2990 2824 3042 2876
rect 4098 2888 4150 2940
rect 4098 2824 4150 2876
rect 4258 2908 4310 2941
rect 4258 2889 4266 2908
rect 4266 2889 4300 2908
rect 4300 2889 4310 2908
rect 4258 2835 4310 2874
rect 4258 2822 4266 2835
rect 4266 2822 4300 2835
rect 4300 2822 4310 2835
rect 4258 2801 4266 2807
rect 4266 2801 4300 2807
rect 4300 2801 4310 2807
rect 445 2630 497 2682
rect 509 2630 561 2682
rect 573 2630 625 2682
rect 445 2364 497 2416
rect 509 2364 561 2416
rect 573 2364 625 2416
rect 958 2714 1010 2720
rect 958 2680 967 2714
rect 967 2680 1001 2714
rect 1001 2680 1010 2714
rect 958 2668 1010 2680
rect 1156 2668 1208 2720
rect 1220 2668 1272 2720
rect 1284 2668 1336 2720
rect 2032 2723 2084 2775
rect 2096 2723 2148 2775
rect 2160 2723 2212 2775
rect 2224 2723 2276 2775
rect 2288 2723 2340 2775
rect 2475 2766 2527 2780
rect 2475 2732 2484 2766
rect 2484 2732 2518 2766
rect 2518 2732 2527 2766
rect 2475 2728 2527 2732
rect 2750 2728 2802 2780
rect 2910 2727 2962 2779
rect 4258 2763 4310 2801
rect 4258 2755 4266 2763
rect 4266 2755 4300 2763
rect 4300 2755 4310 2763
rect 4258 2729 4266 2740
rect 4266 2729 4300 2740
rect 4300 2729 4310 2740
rect 958 2639 1010 2646
rect 958 2605 967 2639
rect 967 2605 1001 2639
rect 1001 2605 1010 2639
rect 958 2594 1010 2605
rect 958 2564 1010 2572
rect 958 2530 967 2564
rect 967 2530 1001 2564
rect 1001 2530 1010 2564
rect 958 2520 1010 2530
rect 958 2489 1010 2498
rect 958 2455 967 2489
rect 967 2455 1001 2489
rect 1001 2455 1010 2489
rect 958 2446 1010 2455
rect 1043 2564 1095 2570
rect 1043 2530 1052 2564
rect 1052 2530 1086 2564
rect 1086 2530 1095 2564
rect 1471 2681 1523 2687
rect 1471 2647 1480 2681
rect 1480 2647 1514 2681
rect 1514 2647 1523 2681
rect 2910 2663 2962 2715
rect 2990 2653 3042 2705
rect 4258 2691 4310 2729
rect 4258 2688 4266 2691
rect 4266 2688 4300 2691
rect 4300 2688 4310 2691
rect 1471 2635 1523 2647
rect 2990 2589 3042 2641
rect 4098 2622 4150 2674
rect 3070 2594 3122 2600
rect 1471 2568 1523 2580
rect 1043 2518 1095 2530
rect 1043 2492 1095 2504
rect 1043 2458 1052 2492
rect 1052 2458 1086 2492
rect 1086 2458 1095 2492
rect 1156 2484 1208 2536
rect 1220 2484 1272 2536
rect 1284 2484 1336 2536
rect 1471 2534 1480 2568
rect 1480 2534 1514 2568
rect 1514 2534 1523 2568
rect 3070 2560 3079 2594
rect 3079 2560 3113 2594
rect 3113 2560 3122 2594
rect 1471 2528 1523 2534
rect 1043 2452 1095 2458
rect 958 2414 1010 2424
rect 958 2380 967 2414
rect 967 2380 1001 2414
rect 1001 2380 1010 2414
rect 958 2372 1010 2380
rect 958 2339 1010 2351
rect 958 2305 967 2339
rect 967 2305 1001 2339
rect 1001 2305 1010 2339
rect 958 2299 1010 2305
rect 1156 2300 1208 2352
rect 1220 2300 1272 2352
rect 1284 2300 1336 2352
rect 1471 2393 1523 2399
rect 1471 2359 1480 2393
rect 1480 2359 1514 2393
rect 1514 2359 1523 2393
rect 1471 2347 1523 2359
rect 1471 2319 1523 2334
rect 1471 2285 1480 2319
rect 1480 2285 1514 2319
rect 1514 2285 1523 2319
rect 1471 2282 1523 2285
rect 1043 2183 1095 2235
rect 1471 2245 1523 2269
rect 1471 2217 1480 2245
rect 1480 2217 1514 2245
rect 1514 2217 1523 2245
rect 849 2125 901 2177
rect 849 2061 901 2113
rect 1043 2117 1095 2169
rect 1471 2171 1523 2204
rect 1156 2116 1208 2168
rect 1220 2116 1272 2168
rect 1284 2116 1336 2168
rect 1471 2152 1480 2171
rect 1480 2152 1514 2171
rect 1514 2152 1523 2171
rect 1471 2137 1480 2139
rect 1480 2137 1514 2139
rect 1514 2137 1523 2139
rect 1471 2097 1523 2137
rect 1471 2087 1480 2097
rect 1480 2087 1514 2097
rect 1514 2087 1523 2097
rect 1471 2063 1480 2074
rect 1480 2063 1514 2074
rect 1514 2063 1523 2074
rect 240 1978 292 2030
rect 335 1986 387 2038
rect 399 1986 451 2038
rect 463 1986 515 2038
rect 1471 2023 1523 2063
rect 240 1914 292 1966
rect 849 1969 901 2021
rect 1471 2022 1480 2023
rect 1480 2022 1514 2023
rect 1514 2022 1523 2023
rect 1471 1989 1480 2009
rect 1480 1989 1514 2009
rect 1514 1989 1523 2009
rect 849 1905 901 1957
rect 958 1938 1010 1944
rect 958 1904 967 1938
rect 967 1904 1001 1938
rect 1001 1904 1010 1938
rect 958 1892 1010 1904
rect 241 1730 293 1736
rect 241 1696 250 1730
rect 250 1696 284 1730
rect 284 1696 293 1730
rect 241 1684 293 1696
rect 241 1657 293 1663
rect 241 1623 250 1657
rect 250 1623 284 1657
rect 284 1623 293 1657
rect 241 1611 293 1623
rect 241 1584 293 1591
rect 241 1550 250 1584
rect 250 1550 284 1584
rect 284 1550 293 1584
rect 241 1539 293 1550
rect 241 1511 293 1519
rect 241 1477 250 1511
rect 250 1477 284 1511
rect 284 1477 293 1511
rect 241 1467 293 1477
rect 241 1438 293 1447
rect 241 1404 250 1438
rect 250 1404 284 1438
rect 284 1404 293 1438
rect 241 1395 293 1404
rect 241 1365 293 1375
rect 241 1331 250 1365
rect 250 1331 284 1365
rect 284 1331 293 1365
rect 241 1323 293 1331
rect 241 1292 293 1303
rect 241 1258 250 1292
rect 250 1258 284 1292
rect 284 1258 293 1292
rect 958 1859 1010 1879
rect 958 1827 967 1859
rect 967 1827 1001 1859
rect 1001 1827 1010 1859
rect 958 1780 1010 1814
rect 958 1762 967 1780
rect 967 1762 1001 1780
rect 1001 1762 1010 1780
rect 958 1746 967 1749
rect 967 1746 1001 1749
rect 1001 1746 1010 1749
rect 958 1701 1010 1746
rect 958 1697 967 1701
rect 967 1697 1001 1701
rect 1001 1697 1010 1701
rect 958 1667 967 1684
rect 967 1667 1001 1684
rect 1001 1667 1010 1684
rect 958 1632 1010 1667
rect 958 1588 967 1620
rect 967 1588 1001 1620
rect 1001 1588 1010 1620
rect 1471 1957 1523 1989
rect 1156 1865 1208 1917
rect 1220 1865 1272 1917
rect 1284 1865 1336 1917
rect 1471 1915 1480 1944
rect 1480 1915 1514 1944
rect 1514 1915 1523 1944
rect 1471 1892 1523 1915
rect 1471 1875 1523 1879
rect 1471 1841 1480 1875
rect 1480 1841 1514 1875
rect 1514 1841 1523 1875
rect 1156 1696 1208 1748
rect 1220 1696 1272 1748
rect 1284 1696 1336 1748
rect 849 1512 901 1564
rect 849 1448 901 1500
rect 958 1568 1010 1588
rect 958 1544 1010 1556
rect 958 1510 967 1544
rect 967 1510 1001 1544
rect 1001 1510 1010 1544
rect 1156 1518 1208 1570
rect 1220 1518 1272 1570
rect 1284 1518 1336 1570
rect 958 1504 1010 1510
rect 687 1330 739 1382
rect 687 1266 739 1318
rect 241 1251 293 1258
rect 241 1219 293 1231
rect 241 1185 250 1219
rect 250 1185 284 1219
rect 284 1185 293 1219
rect 958 1400 1010 1406
rect 958 1366 967 1400
rect 967 1366 1001 1400
rect 1001 1366 1010 1400
rect 958 1354 1010 1366
rect 958 1321 1010 1333
rect 958 1287 967 1321
rect 967 1287 1001 1321
rect 1001 1287 1010 1321
rect 958 1281 1010 1287
rect 241 1179 293 1185
rect 445 1147 497 1199
rect 509 1147 561 1199
rect 573 1147 625 1199
rect 958 1106 1010 1112
rect 769 1044 821 1096
rect 958 1072 967 1106
rect 967 1072 1001 1106
rect 1001 1072 1010 1106
rect 769 980 821 1032
rect 958 1060 1010 1072
rect 958 1030 1010 1042
rect 958 996 967 1030
rect 967 996 1001 1030
rect 1001 996 1010 1030
rect 958 990 1010 996
rect 1043 990 1095 1042
rect 1043 924 1095 976
rect 241 844 250 867
rect 250 844 284 867
rect 284 844 293 867
rect 241 815 293 844
rect 241 800 293 801
rect 241 766 250 800
rect 250 766 284 800
rect 284 766 293 800
rect 241 749 293 766
rect 241 722 293 735
rect 241 688 250 722
rect 250 688 284 722
rect 284 688 293 722
rect 241 683 293 688
rect 241 644 293 669
rect 241 617 250 644
rect 250 617 284 644
rect 284 617 293 644
rect 241 565 293 602
rect 241 550 250 565
rect 250 550 284 565
rect 284 550 293 565
rect 445 795 497 847
rect 509 795 561 847
rect 573 795 625 847
rect 958 870 1010 876
rect 958 836 967 870
rect 967 836 1001 870
rect 1001 836 1010 870
rect 958 824 1010 836
rect 958 756 1010 808
rect 769 692 821 744
rect 769 628 821 680
rect 849 692 901 744
rect 958 728 1010 740
rect 958 694 967 728
rect 967 694 1001 728
rect 1001 694 1010 728
rect 958 688 1010 694
rect 849 628 901 680
rect 241 531 250 535
rect 250 531 284 535
rect 284 531 293 535
rect 241 486 293 531
rect 241 483 250 486
rect 250 483 284 486
rect 284 483 293 486
rect 241 452 250 468
rect 250 452 284 468
rect 284 452 293 468
rect 241 416 293 452
rect 433 443 485 495
rect 497 443 549 495
rect 561 443 613 495
rect 241 373 250 401
rect 250 373 284 401
rect 284 373 293 401
rect 1471 1827 1523 1841
rect 1471 1801 1523 1814
rect 1471 1767 1480 1801
rect 1480 1767 1514 1801
rect 1514 1767 1523 1801
rect 1471 1762 1523 1767
rect 1471 1727 1523 1749
rect 1471 1697 1480 1727
rect 1480 1697 1514 1727
rect 1514 1697 1523 1727
rect 1471 1653 1523 1684
rect 1471 1632 1480 1653
rect 1480 1632 1514 1653
rect 1514 1632 1523 1653
rect 1471 1619 1480 1620
rect 1480 1619 1514 1620
rect 1514 1619 1523 1620
rect 1471 1579 1523 1619
rect 1471 1568 1480 1579
rect 1480 1568 1514 1579
rect 1514 1568 1523 1579
rect 1471 1545 1480 1556
rect 1480 1545 1514 1556
rect 1514 1545 1523 1556
rect 1471 1505 1523 1545
rect 1471 1504 1480 1505
rect 1480 1504 1514 1505
rect 1514 1504 1523 1505
rect 1471 1471 1480 1492
rect 1480 1471 1514 1492
rect 1514 1471 1523 1492
rect 1471 1440 1523 1471
rect 1471 1397 1480 1428
rect 1480 1397 1514 1428
rect 1514 1397 1523 1428
rect 1471 1376 1523 1397
rect 1471 1357 1523 1364
rect 1471 1323 1480 1357
rect 1480 1323 1514 1357
rect 1514 1323 1523 1357
rect 1471 1312 1523 1323
rect 1471 1284 1523 1300
rect 1471 1250 1480 1284
rect 1480 1250 1514 1284
rect 1514 1250 1523 1284
rect 1471 1248 1523 1250
rect 1471 1211 1523 1236
rect 1471 1184 1480 1211
rect 1480 1184 1514 1211
rect 1514 1184 1523 1211
rect 1471 1138 1523 1172
rect 1471 1120 1480 1138
rect 1480 1120 1514 1138
rect 1514 1120 1523 1138
rect 1471 1104 1480 1108
rect 1480 1104 1514 1108
rect 1514 1104 1523 1108
rect 1471 1065 1523 1104
rect 1471 1056 1480 1065
rect 1480 1056 1514 1065
rect 1514 1056 1523 1065
rect 1471 1031 1480 1044
rect 1480 1031 1514 1044
rect 1514 1031 1523 1044
rect 1471 992 1523 1031
rect 1471 958 1480 980
rect 1480 958 1514 980
rect 1514 958 1523 980
rect 1471 928 1523 958
rect 1471 885 1480 916
rect 1480 885 1514 916
rect 1514 885 1523 916
rect 1471 864 1523 885
rect 1471 846 1523 852
rect 1471 812 1480 846
rect 1480 812 1514 846
rect 1514 812 1523 846
rect 1471 800 1523 812
rect 1471 773 1523 788
rect 1471 739 1480 773
rect 1480 739 1514 773
rect 1514 739 1523 773
rect 1471 736 1523 739
rect 1471 700 1523 724
rect 1471 672 1480 700
rect 1480 672 1514 700
rect 1514 672 1523 700
rect 1471 627 1523 660
rect 1471 608 1480 627
rect 1480 608 1514 627
rect 1514 608 1523 627
rect 1471 593 1480 596
rect 1480 593 1514 596
rect 1514 593 1523 596
rect 1471 554 1523 593
rect 1471 544 1480 554
rect 1480 544 1514 554
rect 1514 544 1523 554
rect 1471 520 1480 532
rect 1480 520 1514 532
rect 1514 520 1523 532
rect 1471 481 1523 520
rect 1471 480 1480 481
rect 1480 480 1514 481
rect 1514 480 1523 481
rect 1471 447 1480 468
rect 1480 447 1514 468
rect 1514 447 1523 468
rect 1471 416 1523 447
rect 241 349 293 373
rect 1471 369 1523 404
rect 1471 352 1476 369
rect 1476 352 1523 369
rect 2475 2497 2527 2549
rect 2475 2433 2527 2485
rect 2910 2511 2922 2545
rect 2922 2511 2956 2545
rect 2956 2511 2962 2545
rect 2910 2493 2962 2511
rect 3070 2548 3122 2560
rect 3884 2582 3936 2591
rect 3884 2548 3894 2582
rect 3894 2548 3928 2582
rect 3928 2548 3936 2582
rect 3884 2539 3936 2548
rect 3948 2582 4000 2591
rect 3948 2548 3966 2582
rect 3966 2548 4000 2582
rect 3948 2539 4000 2548
rect 4012 2539 4064 2591
rect 4098 2558 4150 2610
rect 4258 2657 4266 2673
rect 4266 2657 4300 2673
rect 4300 2657 4310 2673
rect 4258 2621 4310 2657
rect 4258 2585 4266 2606
rect 4266 2585 4300 2606
rect 4300 2585 4310 2606
rect 4258 2554 4310 2585
rect 3070 2519 3122 2526
rect 3070 2485 3079 2519
rect 3079 2485 3113 2519
rect 3113 2485 3122 2519
rect 4258 2513 4266 2539
rect 4266 2513 4300 2539
rect 4300 2513 4310 2539
rect 2910 2429 2962 2481
rect 3070 2474 3122 2485
rect 3070 2444 3122 2452
rect 2475 2369 2527 2421
rect 2032 2267 2084 2319
rect 2096 2267 2148 2319
rect 2160 2267 2212 2319
rect 2224 2267 2276 2319
rect 2288 2267 2340 2319
rect 2830 2365 2882 2417
rect 2830 2301 2882 2353
rect 3070 2410 3079 2444
rect 3079 2410 3113 2444
rect 3113 2410 3122 2444
rect 4178 2440 4230 2492
rect 3070 2400 3122 2410
rect 3070 2369 3122 2378
rect 3070 2335 3079 2369
rect 3079 2335 3113 2369
rect 3113 2335 3122 2369
rect 3884 2343 3936 2395
rect 3948 2343 4000 2395
rect 4012 2343 4064 2395
rect 4178 2376 4230 2428
rect 4258 2487 4310 2513
rect 4258 2441 4266 2472
rect 4266 2441 4300 2472
rect 4300 2441 4310 2472
rect 4258 2420 4310 2441
rect 4637 3070 4689 3076
rect 4637 3036 4646 3070
rect 4646 3036 4680 3070
rect 4680 3036 4689 3070
rect 4637 3024 4689 3036
rect 4637 2994 4689 3010
rect 4637 2960 4646 2994
rect 4646 2960 4680 2994
rect 4680 2960 4689 2994
rect 4637 2958 4689 2960
rect 4637 2918 4689 2943
rect 4637 2891 4646 2918
rect 4646 2891 4680 2918
rect 4680 2891 4689 2918
rect 4637 2842 4689 2876
rect 4637 2824 4646 2842
rect 4646 2824 4680 2842
rect 4680 2824 4689 2842
rect 4637 2808 4646 2809
rect 4646 2808 4680 2809
rect 4680 2808 4689 2809
rect 4637 2766 4689 2808
rect 4637 2757 4646 2766
rect 4646 2757 4680 2766
rect 4680 2757 4689 2766
rect 4637 2732 4646 2742
rect 4646 2732 4680 2742
rect 4680 2732 4689 2742
rect 4637 2690 4689 2732
rect 4637 2656 4646 2675
rect 4646 2656 4680 2675
rect 4680 2656 4689 2675
rect 4637 2623 4689 2656
rect 4637 2580 4646 2608
rect 4646 2580 4680 2608
rect 4680 2580 4689 2608
rect 4637 2556 4689 2580
rect 4637 2538 4689 2541
rect 4637 2504 4646 2538
rect 4646 2504 4680 2538
rect 4680 2504 4689 2538
rect 4637 2489 4689 2504
rect 4637 2462 4689 2474
rect 4637 2428 4646 2462
rect 4646 2428 4680 2462
rect 4680 2428 4689 2462
rect 4840 3092 4869 3099
rect 4869 3092 4892 3099
rect 7040 3096 7092 3102
rect 4840 3065 4869 3079
rect 4869 3065 4892 3079
rect 4840 3027 4892 3065
rect 7040 3062 7042 3096
rect 7042 3062 7076 3096
rect 7076 3062 7092 3096
rect 9620 3146 9672 3148
rect 9620 3112 9623 3146
rect 9623 3112 9657 3146
rect 9657 3112 9672 3146
rect 9620 3096 9672 3112
rect 7040 3050 7092 3062
rect 4840 2987 4869 3014
rect 4869 2987 4892 3014
rect 4840 2962 4892 2987
rect 7040 2986 7092 3038
rect 7132 3019 7184 3071
rect 7196 3065 7248 3071
rect 7196 3031 7218 3065
rect 7218 3031 7248 3065
rect 7196 3019 7248 3031
rect 9620 3072 9672 3084
rect 9620 3038 9623 3072
rect 9623 3038 9657 3072
rect 9657 3038 9672 3072
rect 9620 3032 9672 3038
rect 9848 3151 9900 3171
rect 9848 3119 9859 3151
rect 9859 3119 9893 3151
rect 9893 3119 9900 3151
rect 9848 3077 9900 3092
rect 9848 3043 9859 3077
rect 9859 3043 9893 3077
rect 9893 3043 9900 3077
rect 9848 3040 9900 3043
rect 10489 4859 10541 4911
rect 10553 4859 10605 4911
rect 10617 4859 10669 4911
rect 10682 4859 10734 4911
rect 10747 4859 10799 4911
rect 10812 4859 10864 4911
rect 10877 4859 10929 4911
rect 10942 4859 10994 4911
rect 11007 4859 11059 4911
rect 11965 4859 12017 4911
rect 12029 4859 12081 4911
rect 12093 4859 12145 4911
rect 12157 4859 12209 4911
rect 12221 4859 12273 4911
rect 12399 4859 12451 4911
rect 12493 4859 12545 4911
rect 12669 5106 12721 5112
rect 12669 5072 12675 5106
rect 12675 5072 12709 5106
rect 12709 5072 12721 5106
rect 12669 5060 12721 5072
rect 12669 5032 12721 5047
rect 12669 4998 12675 5032
rect 12675 4998 12709 5032
rect 12709 4998 12721 5032
rect 12669 4995 12721 4998
rect 12669 4958 12721 4982
rect 12669 4930 12675 4958
rect 12675 4930 12709 4958
rect 12709 4930 12721 4958
rect 12669 4884 12721 4917
rect 12669 4865 12675 4884
rect 12675 4865 12709 4884
rect 12709 4865 12721 4884
rect 12669 4850 12675 4851
rect 12675 4850 12709 4851
rect 12709 4850 12721 4851
rect 12669 4810 12721 4850
rect 11121 4791 11173 4797
rect 10417 4757 10423 4765
rect 10423 4757 10457 4765
rect 10457 4757 10469 4765
rect 10417 4713 10469 4757
rect 11121 4757 11130 4791
rect 11130 4757 11164 4791
rect 11164 4757 11173 4791
rect 11851 4791 11903 4797
rect 11121 4745 11173 4757
rect 11851 4757 11860 4791
rect 11860 4757 11894 4791
rect 11894 4757 11903 4791
rect 11851 4745 11903 4757
rect 12553 4791 12605 4797
rect 12553 4757 12565 4791
rect 12565 4757 12599 4791
rect 12599 4757 12605 4791
rect 12669 4799 12675 4810
rect 12675 4799 12709 4810
rect 12709 4799 12721 4810
rect 12553 4745 12605 4757
rect 11121 4711 11173 4727
rect 10417 4677 10423 4698
rect 10423 4677 10457 4698
rect 10457 4677 10469 4698
rect 10417 4646 10469 4677
rect 11121 4677 11130 4711
rect 11130 4677 11164 4711
rect 11164 4677 11173 4711
rect 11851 4711 11903 4727
rect 11121 4675 11173 4677
rect 11851 4677 11860 4711
rect 11860 4677 11894 4711
rect 11894 4677 11903 4711
rect 11851 4675 11903 4677
rect 12553 4711 12605 4727
rect 12553 4677 12565 4711
rect 12565 4677 12599 4711
rect 12599 4677 12605 4711
rect 12553 4675 12605 4677
rect 11121 4631 11173 4657
rect 10417 4597 10423 4631
rect 10423 4597 10457 4631
rect 10457 4597 10469 4631
rect 11121 4605 11130 4631
rect 11130 4605 11164 4631
rect 11164 4605 11173 4631
rect 11851 4631 11903 4657
rect 11851 4605 11860 4631
rect 11860 4605 11894 4631
rect 11894 4605 11903 4631
rect 12553 4631 12605 4657
rect 12553 4605 12565 4631
rect 12565 4605 12599 4631
rect 12599 4605 12605 4631
rect 10417 4579 10469 4597
rect 10417 4552 10469 4565
rect 10417 4518 10423 4552
rect 10423 4518 10457 4552
rect 10457 4518 10469 4552
rect 11121 4552 11173 4587
rect 11121 4535 11130 4552
rect 11130 4535 11164 4552
rect 11164 4535 11173 4552
rect 11851 4552 11903 4587
rect 11851 4535 11860 4552
rect 11860 4535 11894 4552
rect 11894 4535 11903 4552
rect 12553 4552 12605 4587
rect 12553 4535 12565 4552
rect 12565 4535 12599 4552
rect 12599 4535 12605 4552
rect 10417 4513 10469 4518
rect 10417 4473 10469 4499
rect 10417 4447 10423 4473
rect 10423 4447 10457 4473
rect 10457 4447 10469 4473
rect 11121 4473 11173 4517
rect 11121 4465 11130 4473
rect 11130 4465 11164 4473
rect 11164 4465 11173 4473
rect 11121 4439 11130 4447
rect 11130 4439 11164 4447
rect 11164 4439 11173 4447
rect 11851 4473 11903 4517
rect 11851 4465 11860 4473
rect 11860 4465 11894 4473
rect 11894 4465 11903 4473
rect 12553 4473 12605 4517
rect 12553 4465 12565 4473
rect 12565 4465 12599 4473
rect 12599 4465 12605 4473
rect 10417 4394 10469 4433
rect 11121 4395 11173 4439
rect 11851 4439 11860 4447
rect 11860 4439 11894 4447
rect 11894 4439 11903 4447
rect 10417 4381 10423 4394
rect 10423 4381 10457 4394
rect 10457 4381 10469 4394
rect 10417 4360 10423 4367
rect 10423 4360 10457 4367
rect 10457 4360 10469 4367
rect 10417 4315 10469 4360
rect 11121 4360 11130 4377
rect 11130 4360 11164 4377
rect 11164 4360 11173 4377
rect 11851 4395 11903 4439
rect 12553 4439 12565 4447
rect 12565 4439 12599 4447
rect 12599 4439 12605 4447
rect 12553 4395 12605 4439
rect 11121 4325 11173 4360
rect 11851 4360 11860 4377
rect 11860 4360 11894 4377
rect 11894 4360 11903 4377
rect 11851 4325 11903 4360
rect 12553 4360 12565 4377
rect 12565 4360 12599 4377
rect 12599 4360 12605 4377
rect 12553 4325 12605 4360
rect 10417 4281 10423 4301
rect 10423 4281 10457 4301
rect 10457 4281 10469 4301
rect 10417 4249 10469 4281
rect 11121 4281 11130 4307
rect 11130 4281 11164 4307
rect 11164 4281 11173 4307
rect 11121 4255 11173 4281
rect 11851 4281 11860 4307
rect 11860 4281 11894 4307
rect 11894 4281 11903 4307
rect 11851 4255 11903 4281
rect 12553 4281 12565 4307
rect 12565 4281 12599 4307
rect 12599 4281 12605 4307
rect 12553 4255 12605 4281
rect 11121 4236 11173 4238
rect 10417 4202 10423 4235
rect 10423 4202 10457 4235
rect 10457 4202 10469 4235
rect 10417 4183 10469 4202
rect 11121 4202 11130 4236
rect 11130 4202 11164 4236
rect 11164 4202 11173 4236
rect 11851 4236 11903 4238
rect 11121 4186 11173 4202
rect 11851 4202 11860 4236
rect 11860 4202 11894 4236
rect 11894 4202 11903 4236
rect 11851 4186 11903 4202
rect 12553 4236 12605 4238
rect 12553 4202 12565 4236
rect 12565 4202 12599 4236
rect 12599 4202 12605 4236
rect 12553 4186 12605 4202
rect 10417 4157 10469 4169
rect 10417 4123 10423 4157
rect 10423 4123 10457 4157
rect 10457 4123 10469 4157
rect 10417 4117 10469 4123
rect 11121 4157 11173 4169
rect 11121 4123 11130 4157
rect 11130 4123 11164 4157
rect 11164 4123 11173 4157
rect 11851 4157 11903 4169
rect 11121 4117 11173 4123
rect 11851 4123 11860 4157
rect 11860 4123 11894 4157
rect 11894 4123 11903 4157
rect 11851 4117 11903 4123
rect 12553 4157 12605 4169
rect 12553 4123 12565 4157
rect 12565 4123 12599 4157
rect 12599 4123 12605 4157
rect 12553 4117 12605 4123
rect 12669 4776 12675 4785
rect 12675 4776 12709 4785
rect 12709 4776 12721 4785
rect 12669 4736 12721 4776
rect 12669 4733 12675 4736
rect 12675 4733 12709 4736
rect 12709 4733 12721 4736
rect 12669 4702 12675 4719
rect 12675 4702 12709 4719
rect 12709 4702 12721 4719
rect 12669 4667 12721 4702
rect 12669 4628 12675 4653
rect 12675 4628 12709 4653
rect 12709 4628 12721 4653
rect 12669 4601 12721 4628
rect 12669 4554 12675 4587
rect 12675 4554 12709 4587
rect 12709 4554 12721 4587
rect 12669 4535 12721 4554
rect 12669 4514 12721 4521
rect 12669 4480 12675 4514
rect 12675 4480 12709 4514
rect 12709 4480 12721 4514
rect 12669 4469 12721 4480
rect 12669 4440 12721 4455
rect 12669 4406 12675 4440
rect 12675 4406 12709 4440
rect 12709 4406 12721 4440
rect 12669 4403 12721 4406
rect 12669 4365 12721 4389
rect 12669 4337 12675 4365
rect 12675 4337 12709 4365
rect 12709 4337 12721 4365
rect 12669 4290 12721 4323
rect 12669 4271 12675 4290
rect 12675 4271 12709 4290
rect 12709 4271 12721 4290
rect 12669 4256 12675 4257
rect 12675 4256 12709 4257
rect 12709 4256 12721 4257
rect 12669 4215 12721 4256
rect 12669 4205 12675 4215
rect 12675 4205 12709 4215
rect 12709 4205 12721 4215
rect 12669 4181 12675 4191
rect 12675 4181 12709 4191
rect 12709 4181 12721 4191
rect 12669 4140 12721 4181
rect 12669 4139 12675 4140
rect 12675 4139 12709 4140
rect 12709 4139 12721 4140
rect 12669 4106 12675 4125
rect 12675 4106 12709 4125
rect 12709 4106 12721 4125
rect 12669 4073 12721 4106
rect 10588 4003 10640 4055
rect 10657 4003 10709 4055
rect 10727 4003 10779 4055
rect 10797 4003 10849 4055
rect 10867 4003 10919 4055
rect 10937 4003 10989 4055
rect 11007 4003 11059 4055
rect 12399 4003 12451 4055
rect 12467 4003 12519 4055
rect 12669 4031 12675 4059
rect 12675 4031 12709 4059
rect 12709 4031 12721 4059
rect 12669 4007 12721 4031
rect 12669 3990 12721 3993
rect 10391 3954 10443 3959
rect 10391 3920 10400 3954
rect 10400 3920 10434 3954
rect 10434 3920 10443 3954
rect 10391 3907 10443 3920
rect 11121 3954 11173 3959
rect 11121 3920 11130 3954
rect 11130 3920 11164 3954
rect 11164 3920 11173 3954
rect 11121 3907 11173 3920
rect 10391 3882 10443 3895
rect 10391 3848 10400 3882
rect 10400 3848 10434 3882
rect 10434 3848 10443 3882
rect 11121 3882 11173 3895
rect 11121 3848 11130 3882
rect 11130 3848 11164 3882
rect 11164 3848 11173 3882
rect 10391 3843 10443 3848
rect 11121 3843 11173 3848
rect 12307 3853 12359 3905
rect 12669 3956 12675 3990
rect 12675 3956 12709 3990
rect 12709 3956 12721 3990
rect 12669 3941 12721 3956
rect 12669 3915 12721 3927
rect 12669 3881 12675 3915
rect 12675 3881 12709 3915
rect 12709 3881 12721 3915
rect 12669 3875 12721 3881
rect 10474 3779 10526 3831
rect 10474 3715 10526 3767
rect 12307 3764 12359 3816
rect 10391 3698 10443 3703
rect 11121 3698 11173 3703
rect 10391 3664 10400 3698
rect 10400 3664 10434 3698
rect 10434 3664 10443 3698
rect 10391 3651 10443 3664
rect 11121 3664 11130 3698
rect 11130 3664 11164 3698
rect 11164 3664 11173 3698
rect 11121 3651 11173 3664
rect 10391 3626 10443 3639
rect 10391 3592 10400 3626
rect 10400 3592 10434 3626
rect 10434 3592 10443 3626
rect 10391 3587 10443 3592
rect 11121 3626 11173 3639
rect 11121 3592 11130 3626
rect 11130 3592 11164 3626
rect 11164 3592 11173 3626
rect 11121 3587 11173 3592
rect 12307 3675 12359 3727
rect 12770 3783 12822 3835
rect 12770 3716 12822 3768
rect 12307 3586 12359 3638
rect 12661 3670 12713 3676
rect 12661 3636 12675 3670
rect 12675 3636 12709 3670
rect 12709 3636 12713 3670
rect 12661 3624 12713 3636
rect 12661 3590 12713 3606
rect 12661 3556 12675 3590
rect 12675 3556 12709 3590
rect 12709 3556 12713 3590
rect 12661 3554 12713 3556
rect 10588 3491 10640 3543
rect 10657 3491 10709 3543
rect 10727 3491 10779 3543
rect 10797 3491 10849 3543
rect 10867 3491 10919 3543
rect 10937 3491 10989 3543
rect 11007 3491 11059 3543
rect 11207 3491 11259 3543
rect 11273 3491 11325 3543
rect 11339 3491 11391 3543
rect 11405 3491 11457 3543
rect 11471 3491 11523 3543
rect 11537 3491 11589 3543
rect 11603 3491 11655 3543
rect 11670 3491 11722 3543
rect 11737 3491 11789 3543
rect 12399 3491 12451 3543
rect 12467 3491 12519 3543
rect 12661 3510 12713 3536
rect 12661 3484 12675 3510
rect 12675 3484 12709 3510
rect 12709 3484 12713 3510
rect 10391 3442 10443 3447
rect 10391 3408 10400 3442
rect 10400 3408 10434 3442
rect 10434 3408 10443 3442
rect 10391 3395 10443 3408
rect 11121 3442 11173 3447
rect 11121 3408 11130 3442
rect 11130 3408 11164 3442
rect 11164 3408 11173 3442
rect 11121 3395 11173 3408
rect 11851 3442 11903 3447
rect 11851 3408 11860 3442
rect 11860 3408 11894 3442
rect 11894 3408 11903 3442
rect 11851 3395 11903 3408
rect 12581 3442 12633 3447
rect 12581 3408 12590 3442
rect 12590 3408 12624 3442
rect 12624 3408 12633 3442
rect 12581 3395 12633 3408
rect 10391 3370 10443 3383
rect 10391 3336 10400 3370
rect 10400 3336 10434 3370
rect 10434 3336 10443 3370
rect 11121 3370 11173 3383
rect 11121 3336 11130 3370
rect 11130 3336 11164 3370
rect 11164 3336 11173 3370
rect 10391 3331 10443 3336
rect 11121 3331 11173 3336
rect 11851 3370 11903 3383
rect 11851 3336 11860 3370
rect 11860 3336 11894 3370
rect 11894 3336 11903 3370
rect 11851 3331 11903 3336
rect 12581 3370 12633 3383
rect 12581 3336 12590 3370
rect 12590 3336 12624 3370
rect 12624 3336 12633 3370
rect 12581 3331 12633 3336
rect 12661 3430 12713 3466
rect 12661 3414 12675 3430
rect 12675 3414 12709 3430
rect 12709 3414 12713 3430
rect 12661 3350 12713 3395
rect 12661 3343 12675 3350
rect 12675 3343 12709 3350
rect 12709 3343 12713 3350
rect 10474 3267 10526 3319
rect 12661 3316 12675 3324
rect 12675 3316 12709 3324
rect 12709 3316 12713 3324
rect 10474 3203 10526 3255
rect 12473 3226 12525 3278
rect 12473 3162 12525 3214
rect 12661 3272 12713 3316
rect 12661 3236 12675 3253
rect 12675 3236 12709 3253
rect 12709 3236 12713 3253
rect 12661 3201 12713 3236
rect 12581 3186 12633 3191
rect 12581 3152 12590 3186
rect 12590 3152 12624 3186
rect 12624 3152 12633 3186
rect 12581 3139 12633 3152
rect 12581 3114 12633 3127
rect 4840 2943 4892 2949
rect 4840 2909 4869 2943
rect 4869 2909 4892 2943
rect 4840 2897 4892 2909
rect 8783 2900 8835 2952
rect 8847 2900 8899 2952
rect 12581 3080 12590 3114
rect 12590 3080 12624 3114
rect 12624 3080 12633 3114
rect 12581 3075 12633 3080
rect 12661 3156 12675 3182
rect 12675 3156 12709 3182
rect 12709 3156 12713 3182
rect 12661 3130 12713 3156
rect 12661 3109 12713 3111
rect 12661 3075 12675 3109
rect 12675 3075 12709 3109
rect 12709 3075 12713 3109
rect 10391 3058 10443 3063
rect 10391 3024 10400 3058
rect 10400 3024 10434 3058
rect 10434 3024 10443 3058
rect 12661 3059 12713 3075
rect 10391 3011 10443 3024
rect 10391 2986 10443 2999
rect 10391 2952 10400 2986
rect 10400 2952 10434 2986
rect 10434 2952 10443 2986
rect 10588 2979 10640 3031
rect 10657 2979 10709 3031
rect 10727 2979 10779 3031
rect 10797 2979 10849 3031
rect 10867 2979 10919 3031
rect 10937 2979 10989 3031
rect 11007 2979 11059 3031
rect 11207 2979 11259 3031
rect 11273 2979 11325 3031
rect 11339 2979 11391 3031
rect 11405 2979 11457 3031
rect 11471 2979 11523 3031
rect 11537 2979 11589 3031
rect 11603 2979 11655 3031
rect 11670 2979 11722 3031
rect 11737 2979 11789 3031
rect 11965 2979 12017 3031
rect 12029 2979 12081 3031
rect 12093 2979 12145 3031
rect 12157 2979 12209 3031
rect 12221 2979 12273 3031
rect 12661 3028 12713 3040
rect 12661 2994 12675 3028
rect 12675 2994 12709 3028
rect 12709 2994 12713 3028
rect 12661 2988 12713 2994
rect 10391 2947 10443 2952
rect 13879 5046 13995 5162
rect 4840 2865 4892 2884
rect 4840 2832 4869 2865
rect 4869 2832 4892 2865
rect 4840 2787 4892 2818
rect 4840 2766 4869 2787
rect 4869 2766 4892 2787
rect 4840 2709 4892 2752
rect 6963 2783 7015 2795
rect 6963 2749 6970 2783
rect 6970 2749 7004 2783
rect 7004 2749 7015 2783
rect 6963 2743 7015 2749
rect 7027 2783 7079 2795
rect 7027 2749 7042 2783
rect 7042 2749 7076 2783
rect 7076 2749 7079 2783
rect 7027 2743 7079 2749
rect 7132 2739 7184 2791
rect 7196 2785 7248 2791
rect 7196 2751 7218 2785
rect 7218 2751 7248 2785
rect 7196 2739 7248 2751
rect 10474 2755 10526 2807
rect 4840 2700 4869 2709
rect 4869 2700 4892 2709
rect 4840 2675 4869 2686
rect 4869 2675 4892 2686
rect 4840 2634 4892 2675
rect 5345 2660 5397 2712
rect 5409 2660 5461 2712
rect 8638 2658 8690 2710
rect 8702 2658 8754 2710
rect 10474 2691 10526 2743
rect 12473 2766 12525 2807
rect 12473 2755 12474 2766
rect 12474 2755 12525 2766
rect 12473 2732 12474 2743
rect 12474 2732 12525 2743
rect 12473 2691 12525 2732
rect 12581 2802 12633 2807
rect 12581 2768 12590 2802
rect 12590 2768 12624 2802
rect 12624 2768 12633 2802
rect 12581 2755 12633 2768
rect 12581 2730 12633 2743
rect 12581 2696 12590 2730
rect 12590 2696 12624 2730
rect 12624 2696 12633 2730
rect 12581 2691 12633 2696
rect 12661 2789 12713 2796
rect 12661 2755 12670 2789
rect 12670 2755 12704 2789
rect 12704 2755 12713 2789
rect 12661 2744 12713 2755
rect 12661 2706 12713 2714
rect 12661 2672 12670 2706
rect 12670 2672 12704 2706
rect 12704 2672 12713 2706
rect 12661 2662 12713 2672
rect 12661 2622 12713 2632
rect 4840 2597 4869 2620
rect 4869 2597 4892 2620
rect 4840 2568 4892 2597
rect 4840 2553 4892 2554
rect 4840 2519 4869 2553
rect 4869 2519 4892 2553
rect 6638 2535 6690 2587
rect 6702 2535 6754 2587
rect 10391 2546 10443 2551
rect 12661 2588 12670 2622
rect 12670 2588 12704 2622
rect 12704 2588 12713 2622
rect 12661 2580 12713 2588
rect 4840 2502 4892 2519
rect 10391 2512 10400 2546
rect 10400 2512 10434 2546
rect 10434 2512 10443 2546
rect 12661 2538 12713 2549
rect 4840 2476 4892 2488
rect 4840 2442 4869 2476
rect 4869 2442 4892 2476
rect 7046 2458 7098 2510
rect 7110 2458 7162 2510
rect 10391 2499 10443 2512
rect 10391 2474 10443 2487
rect 4840 2436 4892 2442
rect 4637 2422 4689 2428
rect 4258 2403 4310 2405
rect 4258 2369 4266 2403
rect 4266 2369 4300 2403
rect 4300 2369 4310 2403
rect 4258 2353 4310 2369
rect 3070 2326 3122 2335
rect 3070 2294 3122 2304
rect 2990 2209 3042 2261
rect 2990 2145 3042 2197
rect 3070 2260 3079 2294
rect 3079 2260 3113 2294
rect 3113 2260 3122 2294
rect 4258 2331 4310 2338
rect 4258 2297 4266 2331
rect 4266 2297 4300 2331
rect 4300 2297 4310 2331
rect 4258 2286 4310 2297
rect 3070 2252 3122 2260
rect 3070 2219 3122 2230
rect 3070 2185 3079 2219
rect 3079 2185 3113 2219
rect 3113 2185 3122 2219
rect 3070 2178 3122 2185
rect 3070 2144 3122 2156
rect 2830 2053 2882 2105
rect 3070 2110 3079 2144
rect 3079 2110 3113 2144
rect 3113 2110 3122 2144
rect 4258 2259 4310 2271
rect 4418 2330 4470 2382
rect 7132 2378 7184 2430
rect 7196 2378 7248 2430
rect 10391 2440 10400 2474
rect 10400 2440 10434 2474
rect 10434 2440 10443 2474
rect 10588 2467 10640 2519
rect 10657 2467 10709 2519
rect 10727 2467 10779 2519
rect 10797 2467 10849 2519
rect 10867 2467 10919 2519
rect 10937 2467 10989 2519
rect 11007 2467 11059 2519
rect 11207 2467 11259 2519
rect 11273 2467 11325 2519
rect 11339 2467 11391 2519
rect 11405 2467 11457 2519
rect 11471 2467 11523 2519
rect 11537 2467 11589 2519
rect 11603 2467 11655 2519
rect 11670 2467 11722 2519
rect 11737 2467 11789 2519
rect 11965 2467 12017 2519
rect 12029 2467 12081 2519
rect 12093 2467 12145 2519
rect 12157 2467 12209 2519
rect 12221 2467 12273 2519
rect 12661 2504 12670 2538
rect 12670 2504 12704 2538
rect 12704 2504 12713 2538
rect 12661 2497 12713 2504
rect 10391 2435 10443 2440
rect 4418 2266 4470 2318
rect 9620 2345 9672 2397
rect 9620 2281 9672 2333
rect 10172 2315 10224 2367
rect 4258 2225 4266 2259
rect 4266 2225 4300 2259
rect 4300 2225 4310 2259
rect 10172 2251 10224 2303
rect 10391 2277 10443 2283
rect 10391 2243 10400 2277
rect 10400 2243 10434 2277
rect 10434 2243 10443 2277
rect 4258 2219 4310 2225
rect 3884 2139 3936 2191
rect 3948 2139 4000 2191
rect 4012 2139 4064 2191
rect 3070 2104 3122 2110
rect 2830 1989 2882 2041
rect 3070 1984 3122 1990
rect 2032 1811 2084 1863
rect 2096 1811 2148 1863
rect 2160 1811 2212 1863
rect 2224 1811 2276 1863
rect 2288 1811 2340 1863
rect 2990 1897 3042 1949
rect 2830 1782 2882 1834
rect 2990 1833 3042 1885
rect 3070 1950 3079 1984
rect 3079 1950 3113 1984
rect 3113 1950 3122 1984
rect 4258 1984 4310 1990
rect 3070 1938 3122 1950
rect 3070 1886 3122 1895
rect 3070 1852 3079 1886
rect 3079 1852 3113 1886
rect 3113 1852 3122 1886
rect 3070 1843 3122 1852
rect 2830 1718 2882 1770
rect 4098 1914 4150 1966
rect 4098 1850 4150 1902
rect 4258 1950 4266 1984
rect 4266 1950 4300 1984
rect 4300 1950 4310 1984
rect 4258 1938 4310 1950
rect 4258 1863 4310 1875
rect 4258 1829 4266 1863
rect 4266 1829 4300 1863
rect 4300 1829 4310 1863
rect 10391 2231 10443 2243
rect 10391 2205 10443 2219
rect 10391 2171 10400 2205
rect 10400 2171 10434 2205
rect 10434 2171 10443 2205
rect 10474 2243 10526 2295
rect 12473 2284 12525 2336
rect 10474 2179 10526 2231
rect 12473 2220 12525 2272
rect 10391 2167 10443 2171
rect 6634 2066 6686 2118
rect 6698 2066 6750 2118
rect 6164 1940 6216 1992
rect 6243 1940 6295 1992
rect 6322 1940 6374 1992
rect 6401 1940 6453 1992
rect 8946 1940 8998 1992
rect 9013 1940 9065 1992
rect 9080 1940 9132 1992
rect 4258 1823 4310 1829
rect 3070 1789 3122 1801
rect 3070 1755 3079 1789
rect 3079 1755 3113 1789
rect 3113 1755 3122 1789
rect 3070 1749 3122 1755
rect 4418 1731 4470 1783
rect 4749 1736 4801 1788
rect 4418 1667 4470 1719
rect 4637 1681 4689 1687
rect 4637 1647 4646 1681
rect 4646 1647 4680 1681
rect 4680 1647 4689 1681
rect 4637 1635 4689 1647
rect 2032 1355 2084 1407
rect 2096 1355 2148 1407
rect 2160 1355 2212 1407
rect 2224 1355 2276 1407
rect 2288 1355 2340 1407
rect 2830 1429 2882 1481
rect 2830 1365 2882 1417
rect 3070 1590 3122 1596
rect 3070 1556 3079 1590
rect 3079 1556 3113 1590
rect 3113 1556 3122 1590
rect 3070 1544 3122 1556
rect 3070 1514 3122 1522
rect 3070 1480 3079 1514
rect 3079 1480 3113 1514
rect 3113 1480 3122 1514
rect 3070 1470 3122 1480
rect 4637 1600 4689 1609
rect 4637 1566 4646 1600
rect 4646 1566 4680 1600
rect 4680 1566 4689 1600
rect 4637 1557 4689 1566
rect 4637 1520 4689 1530
rect 4637 1486 4646 1520
rect 4646 1486 4680 1520
rect 4680 1486 4689 1520
rect 4637 1478 4689 1486
rect 3070 1439 3122 1449
rect 3070 1405 3079 1439
rect 3079 1405 3113 1439
rect 3113 1405 3122 1439
rect 3070 1397 3122 1405
rect 3070 1364 3122 1376
rect 3070 1330 3079 1364
rect 3079 1330 3113 1364
rect 3113 1330 3122 1364
rect 4749 1671 4801 1723
rect 6898 1700 6950 1752
rect 6962 1700 7014 1752
rect 7271 1700 7323 1752
rect 7335 1700 7387 1752
rect 4749 1606 4801 1658
rect 4749 1540 4801 1592
rect 5043 1572 5095 1615
rect 4749 1474 4801 1526
rect 5043 1563 5049 1572
rect 5049 1563 5083 1572
rect 5083 1563 5095 1572
rect 5113 1572 5165 1615
rect 5113 1563 5121 1572
rect 5121 1563 5155 1572
rect 5155 1563 5165 1572
rect 5183 1572 5235 1615
rect 5183 1563 5193 1572
rect 5193 1563 5227 1572
rect 5227 1563 5235 1572
rect 5253 1572 5305 1615
rect 5837 1572 5889 1615
rect 5253 1563 5265 1572
rect 5265 1563 5299 1572
rect 5299 1563 5305 1572
rect 5043 1538 5049 1551
rect 5049 1538 5083 1551
rect 5083 1538 5095 1551
rect 5043 1499 5095 1538
rect 5113 1538 5121 1551
rect 5121 1538 5155 1551
rect 5155 1538 5165 1551
rect 5113 1499 5165 1538
rect 5183 1538 5193 1551
rect 5193 1538 5227 1551
rect 5227 1538 5235 1551
rect 5183 1499 5235 1538
rect 5253 1538 5265 1551
rect 5265 1538 5299 1551
rect 5299 1538 5305 1551
rect 5837 1563 5841 1572
rect 5841 1563 5875 1572
rect 5875 1563 5889 1572
rect 5903 1572 5955 1615
rect 5903 1563 5913 1572
rect 5913 1563 5947 1572
rect 5947 1563 5955 1572
rect 5970 1572 6022 1615
rect 6142 1572 6194 1615
rect 6211 1572 6263 1615
rect 6281 1572 6333 1615
rect 6351 1572 6403 1615
rect 6421 1572 6473 1615
rect 9459 1589 9511 1641
rect 7505 1572 7557 1578
rect 7578 1572 7630 1578
rect 7651 1572 7703 1578
rect 7724 1572 7776 1578
rect 7796 1572 7848 1578
rect 7868 1572 7920 1578
rect 7940 1572 7992 1578
rect 8012 1572 8064 1578
rect 8187 1572 8239 1578
rect 8289 1572 8341 1578
rect 8390 1572 8442 1578
rect 8953 1572 9005 1577
rect 9080 1572 9132 1577
rect 5970 1563 5985 1572
rect 5985 1563 6019 1572
rect 6019 1563 6022 1572
rect 5837 1538 5841 1551
rect 5841 1538 5875 1551
rect 5875 1538 5889 1551
rect 5253 1499 5305 1538
rect 5837 1499 5889 1538
rect 5903 1538 5913 1551
rect 5913 1538 5947 1551
rect 5947 1538 5955 1551
rect 5903 1499 5955 1538
rect 5970 1538 5985 1551
rect 5985 1538 6019 1551
rect 6019 1538 6022 1551
rect 6142 1563 6163 1572
rect 6163 1563 6194 1572
rect 6211 1563 6235 1572
rect 6235 1563 6263 1572
rect 6281 1563 6307 1572
rect 6307 1563 6333 1572
rect 6351 1563 6379 1572
rect 6379 1563 6403 1572
rect 6421 1563 6451 1572
rect 6451 1563 6473 1572
rect 6142 1538 6163 1551
rect 6163 1538 6194 1551
rect 6211 1538 6235 1551
rect 6235 1538 6263 1551
rect 6281 1538 6307 1551
rect 6307 1538 6333 1551
rect 6351 1538 6379 1551
rect 6379 1538 6403 1551
rect 6421 1538 6451 1551
rect 6451 1538 6473 1551
rect 7505 1538 7531 1572
rect 7531 1538 7557 1572
rect 7578 1538 7603 1572
rect 7603 1538 7630 1572
rect 7651 1538 7675 1572
rect 7675 1538 7703 1572
rect 7724 1538 7747 1572
rect 7747 1538 7776 1572
rect 7796 1538 7819 1572
rect 7819 1538 7848 1572
rect 7868 1538 7891 1572
rect 7891 1538 7920 1572
rect 7940 1538 7963 1572
rect 7963 1538 7992 1572
rect 8012 1538 8035 1572
rect 8035 1538 8064 1572
rect 8187 1538 8217 1572
rect 8217 1538 8239 1572
rect 8289 1538 8323 1572
rect 8323 1538 8341 1572
rect 8390 1538 8395 1572
rect 8395 1538 8433 1572
rect 8433 1538 8442 1572
rect 8953 1538 8971 1572
rect 8971 1538 9005 1572
rect 9080 1538 9083 1572
rect 9083 1538 9117 1572
rect 9117 1538 9132 1572
rect 5970 1499 6022 1538
rect 6142 1499 6194 1538
rect 6211 1499 6263 1538
rect 6281 1499 6333 1538
rect 6351 1499 6403 1538
rect 6421 1499 6473 1538
rect 7505 1526 7557 1538
rect 7578 1526 7630 1538
rect 7651 1526 7703 1538
rect 7724 1526 7776 1538
rect 7796 1526 7848 1538
rect 7868 1526 7920 1538
rect 7940 1526 7992 1538
rect 8012 1526 8064 1538
rect 8187 1526 8239 1538
rect 8289 1526 8341 1538
rect 8390 1526 8442 1538
rect 8953 1525 9005 1538
rect 9080 1525 9132 1538
rect 9459 1523 9511 1575
rect 9459 1502 9511 1509
rect 9459 1468 9468 1502
rect 9468 1468 9502 1502
rect 9502 1468 9511 1502
rect 4637 1440 4689 1451
rect 4637 1406 4646 1440
rect 4646 1406 4680 1440
rect 4680 1406 4689 1440
rect 9459 1457 9511 1468
rect 9459 1428 9511 1443
rect 4637 1399 4689 1406
rect 3070 1324 3122 1330
rect 3884 1256 3936 1308
rect 3948 1256 4000 1308
rect 4012 1256 4064 1308
rect 2830 1158 2882 1210
rect 2830 1094 2882 1146
rect 3070 1204 3122 1210
rect 3070 1170 3079 1204
rect 3079 1170 3113 1204
rect 3113 1170 3122 1204
rect 3070 1158 3122 1170
rect 3070 1130 3122 1138
rect 3070 1096 3079 1130
rect 3079 1096 3113 1130
rect 3113 1096 3122 1130
rect 3070 1086 3122 1096
rect 4258 1364 4310 1370
rect 4258 1330 4266 1364
rect 4266 1330 4300 1364
rect 4300 1330 4310 1364
rect 4258 1318 4310 1330
rect 4637 1360 4689 1372
rect 4637 1326 4646 1360
rect 4646 1326 4680 1360
rect 4680 1326 4689 1360
rect 8554 1365 8606 1417
rect 9459 1394 9468 1428
rect 9468 1394 9502 1428
rect 9502 1394 9511 1428
rect 4637 1320 4689 1326
rect 8554 1301 8606 1353
rect 9459 1391 9511 1394
rect 9459 1354 9511 1377
rect 9459 1325 9468 1354
rect 9468 1325 9502 1354
rect 9502 1325 9511 1354
rect 9459 1280 9511 1311
rect 4258 1250 4310 1262
rect 4258 1216 4266 1250
rect 4266 1216 4300 1250
rect 4300 1216 4310 1250
rect 9459 1259 9468 1280
rect 9468 1259 9502 1280
rect 9502 1259 9511 1280
rect 4178 1158 4230 1210
rect 4258 1210 4310 1216
rect 9459 1206 9511 1244
rect 9459 1192 9468 1206
rect 9468 1192 9502 1206
rect 9502 1192 9511 1206
rect 4178 1094 4230 1146
rect 9459 1172 9468 1177
rect 9468 1172 9502 1177
rect 9502 1172 9511 1177
rect 9459 1132 9511 1172
rect 9459 1125 9468 1132
rect 9468 1125 9502 1132
rect 9502 1125 9511 1132
rect 9459 1098 9468 1110
rect 9468 1098 9502 1110
rect 9502 1098 9511 1110
rect 3070 1057 3122 1067
rect 3070 1023 3079 1057
rect 3079 1023 3113 1057
rect 3113 1023 3122 1057
rect 9459 1058 9511 1098
rect 9459 1024 9468 1043
rect 9468 1024 9502 1043
rect 9502 1024 9511 1043
rect 3070 1015 3122 1023
rect 3070 984 3122 996
rect 2032 899 2084 951
rect 2096 899 2148 951
rect 2160 899 2212 951
rect 2224 899 2276 951
rect 2288 899 2340 951
rect 2572 929 2624 981
rect 2636 929 2688 981
rect 3070 950 3079 984
rect 3079 950 3113 984
rect 3113 950 3122 984
rect 3070 944 3122 950
rect 3884 940 3936 992
rect 3948 940 4000 992
rect 4012 940 4064 992
rect 6842 967 6894 1019
rect 6906 967 6958 1019
rect 9459 991 9511 1024
rect 9459 950 9468 976
rect 9468 950 9502 976
rect 9502 950 9511 976
rect 9459 924 9511 950
rect 2750 843 2802 895
rect 2814 843 2866 895
rect 9459 876 9468 909
rect 9468 876 9502 909
rect 9502 876 9511 909
rect 9459 857 9511 876
rect 9459 836 9511 842
rect 2940 776 2992 828
rect 2940 712 2992 764
rect 4112 778 4164 830
rect 3070 695 3122 701
rect 3070 661 3079 695
rect 3079 661 3113 695
rect 3113 661 3122 695
rect 3070 649 3122 661
rect 3070 623 3122 628
rect 3070 589 3079 623
rect 3079 589 3113 623
rect 3113 589 3122 623
rect 3070 576 3122 589
rect 3070 551 3122 555
rect 2032 443 2084 495
rect 2096 443 2148 495
rect 2160 443 2212 495
rect 2224 443 2276 495
rect 2288 443 2340 495
rect 2572 473 2624 525
rect 2636 473 2688 525
rect 3070 517 3079 551
rect 3079 517 3113 551
rect 3113 517 3122 551
rect 3070 503 3122 517
rect 3070 479 3122 482
rect 3070 445 3079 479
rect 3079 445 3113 479
rect 3113 445 3122 479
rect 4112 704 4164 756
rect 3884 630 3936 682
rect 3948 630 4000 682
rect 4012 630 4064 682
rect 4112 630 4164 682
rect 4112 557 4164 609
rect 4112 484 4164 536
rect 4258 692 4310 698
rect 4258 658 4266 692
rect 4266 658 4300 692
rect 4300 658 4310 692
rect 4258 646 4310 658
rect 9459 802 9468 836
rect 9468 802 9502 836
rect 9502 802 9511 836
rect 9459 790 9511 802
rect 9459 763 9511 775
rect 9459 729 9468 763
rect 9468 729 9502 763
rect 9502 729 9511 763
rect 9459 723 9511 729
rect 9459 690 9511 708
rect 9459 656 9468 690
rect 9468 656 9502 690
rect 9502 656 9511 690
rect 4258 616 4310 624
rect 9459 617 9511 641
rect 4258 582 4266 616
rect 4266 582 4300 616
rect 4300 582 4310 616
rect 9459 589 9468 617
rect 9468 589 9502 617
rect 9502 589 9511 617
rect 4258 572 4310 582
rect 4258 540 4310 550
rect 9459 544 9511 574
rect 4258 506 4266 540
rect 4266 506 4300 540
rect 4300 506 4310 540
rect 9459 522 9468 544
rect 9468 522 9502 544
rect 9502 522 9511 544
rect 4258 498 4310 506
rect 4258 465 4310 477
rect 3070 430 3122 445
rect 4258 431 4266 465
rect 4266 431 4300 465
rect 4300 431 4310 465
rect 4258 425 4310 431
rect 4637 448 4689 463
rect 9459 471 9511 507
rect 12661 2249 12713 2254
rect 12661 2215 12675 2249
rect 12675 2215 12709 2249
rect 12709 2215 12713 2249
rect 12661 2202 12713 2215
rect 12661 2174 12713 2190
rect 12661 2140 12675 2174
rect 12675 2140 12709 2174
rect 12709 2140 12713 2174
rect 12661 2138 12713 2140
rect 12661 2099 12713 2126
rect 12661 2074 12675 2099
rect 12675 2074 12709 2099
rect 12709 2074 12713 2099
rect 12661 2024 12713 2062
rect 12661 2010 12675 2024
rect 12675 2010 12709 2024
rect 12709 2010 12713 2024
rect 10588 1955 10640 2007
rect 10657 1955 10709 2007
rect 10727 1955 10779 2007
rect 10797 1955 10849 2007
rect 10867 1955 10919 2007
rect 10937 1955 10989 2007
rect 11007 1955 11059 2007
rect 11207 1955 11259 2007
rect 11274 1955 11326 2007
rect 11341 1955 11393 2007
rect 11600 1955 11652 2007
rect 11668 1955 11720 2007
rect 11737 1955 11789 2007
rect 12399 1955 12451 2007
rect 12467 1955 12519 2007
rect 12661 1990 12675 1998
rect 12675 1990 12709 1998
rect 12709 1990 12713 1998
rect 12661 1949 12713 1990
rect 12661 1946 12675 1949
rect 12675 1946 12709 1949
rect 12709 1946 12713 1949
rect 9732 782 9784 834
rect 9732 718 9784 770
rect 10008 1347 10060 1399
rect 10008 1283 10060 1335
rect 10391 1906 10443 1911
rect 10089 795 10141 796
rect 10089 761 10095 795
rect 10095 761 10129 795
rect 10129 761 10141 795
rect 10089 744 10141 761
rect 10089 720 10141 732
rect 10089 686 10095 720
rect 10095 686 10129 720
rect 10129 686 10141 720
rect 10089 680 10141 686
rect 10391 1872 10400 1906
rect 10400 1872 10434 1906
rect 10434 1872 10443 1906
rect 10391 1859 10443 1872
rect 11121 1906 11173 1911
rect 11121 1872 11130 1906
rect 11130 1872 11164 1906
rect 11164 1872 11173 1906
rect 11121 1859 11173 1872
rect 10391 1834 10443 1847
rect 10391 1800 10400 1834
rect 10400 1800 10434 1834
rect 10434 1800 10443 1834
rect 11121 1834 11173 1847
rect 11121 1800 11130 1834
rect 11130 1800 11164 1834
rect 11164 1800 11173 1834
rect 10391 1795 10443 1800
rect 11121 1795 11173 1800
rect 12307 1860 12359 1912
rect 10474 1731 10526 1783
rect 12307 1781 12359 1833
rect 10474 1667 10526 1719
rect 12307 1701 12359 1753
rect 10391 1650 10443 1655
rect 11121 1650 11173 1655
rect 10391 1616 10400 1650
rect 10400 1616 10434 1650
rect 10434 1616 10443 1650
rect 10391 1603 10443 1616
rect 11121 1616 11130 1650
rect 11130 1616 11164 1650
rect 11164 1616 11173 1650
rect 11121 1603 11173 1616
rect 10391 1578 10443 1591
rect 10391 1544 10400 1578
rect 10400 1544 10434 1578
rect 10434 1544 10443 1578
rect 10391 1539 10443 1544
rect 11121 1578 11173 1591
rect 11121 1544 11130 1578
rect 11130 1544 11164 1578
rect 11164 1544 11173 1578
rect 11121 1539 11173 1544
rect 12307 1621 12359 1673
rect 12307 1541 12359 1593
rect 12661 1915 12675 1934
rect 12675 1915 12709 1934
rect 12709 1915 12713 1934
rect 12661 1882 12713 1915
rect 12661 1840 12675 1870
rect 12675 1840 12709 1870
rect 12709 1840 12713 1870
rect 12661 1818 12713 1840
rect 12661 1799 12713 1806
rect 12661 1765 12675 1799
rect 12675 1765 12709 1799
rect 12709 1765 12713 1799
rect 12661 1754 12713 1765
rect 12661 1724 12713 1742
rect 12661 1690 12675 1724
rect 12675 1690 12709 1724
rect 12709 1690 12713 1724
rect 12661 1649 12713 1678
rect 12661 1626 12675 1649
rect 12675 1626 12709 1649
rect 12709 1626 12713 1649
rect 12661 1574 12713 1614
rect 12661 1562 12675 1574
rect 12675 1562 12709 1574
rect 12709 1562 12713 1574
rect 12661 1540 12675 1550
rect 12675 1540 12709 1550
rect 12709 1540 12713 1550
rect 12661 1499 12713 1540
rect 12661 1498 12675 1499
rect 12675 1498 12709 1499
rect 12709 1498 12713 1499
rect 10588 1443 10640 1495
rect 10657 1443 10709 1495
rect 10727 1443 10779 1495
rect 10797 1443 10849 1495
rect 10867 1443 10919 1495
rect 10937 1443 10989 1495
rect 11007 1443 11059 1495
rect 12399 1443 12451 1495
rect 12467 1443 12519 1495
rect 12661 1465 12675 1486
rect 12675 1465 12709 1486
rect 12709 1465 12713 1486
rect 12661 1434 12713 1465
rect 12661 1390 12675 1422
rect 12675 1390 12709 1422
rect 12709 1390 12713 1422
rect 10416 1375 10468 1381
rect 10416 1341 10423 1375
rect 10423 1341 10457 1375
rect 10457 1341 10468 1375
rect 10416 1329 10468 1341
rect 11121 1375 11173 1381
rect 11121 1341 11130 1375
rect 11130 1341 11164 1375
rect 11164 1341 11173 1375
rect 11121 1329 11173 1341
rect 11851 1375 11903 1381
rect 11851 1341 11860 1375
rect 11860 1341 11894 1375
rect 11894 1341 11903 1375
rect 11851 1329 11903 1341
rect 12553 1375 12605 1381
rect 12553 1341 12565 1375
rect 12565 1341 12599 1375
rect 12599 1341 12605 1375
rect 12553 1329 12605 1341
rect 10416 1295 10468 1311
rect 10416 1261 10423 1295
rect 10423 1261 10457 1295
rect 10457 1261 10468 1295
rect 10416 1259 10468 1261
rect 11121 1295 11173 1311
rect 11121 1261 11130 1295
rect 11130 1261 11164 1295
rect 11164 1261 11173 1295
rect 11121 1259 11173 1261
rect 11851 1295 11903 1311
rect 11851 1261 11860 1295
rect 11860 1261 11894 1295
rect 11894 1261 11903 1295
rect 11851 1259 11903 1261
rect 12553 1295 12605 1311
rect 12553 1261 12565 1295
rect 12565 1261 12599 1295
rect 12599 1261 12605 1295
rect 12553 1259 12605 1261
rect 10416 1215 10468 1241
rect 10416 1189 10423 1215
rect 10423 1189 10457 1215
rect 10457 1189 10468 1215
rect 11121 1215 11173 1241
rect 11121 1189 11130 1215
rect 11130 1189 11164 1215
rect 11164 1189 11173 1215
rect 11851 1215 11903 1241
rect 11851 1189 11860 1215
rect 11860 1189 11894 1215
rect 11894 1189 11903 1215
rect 12553 1215 12605 1241
rect 12553 1189 12565 1215
rect 12565 1189 12599 1215
rect 12599 1189 12605 1215
rect 10416 1136 10468 1171
rect 10416 1119 10423 1136
rect 10423 1119 10457 1136
rect 10457 1119 10468 1136
rect 11121 1136 11173 1171
rect 11121 1119 11130 1136
rect 11130 1119 11164 1136
rect 11164 1119 11173 1136
rect 11851 1136 11903 1171
rect 11851 1119 11860 1136
rect 11860 1119 11894 1136
rect 11894 1119 11903 1136
rect 12553 1136 12605 1171
rect 12553 1119 12565 1136
rect 12565 1119 12599 1136
rect 12599 1119 12605 1136
rect 10416 1057 10468 1101
rect 10416 1049 10423 1057
rect 10423 1049 10457 1057
rect 10457 1049 10468 1057
rect 11121 1057 11173 1101
rect 11121 1049 11130 1057
rect 11130 1049 11164 1057
rect 11164 1049 11173 1057
rect 11851 1057 11903 1101
rect 11851 1049 11860 1057
rect 11860 1049 11894 1057
rect 11894 1049 11903 1057
rect 12553 1057 12605 1101
rect 12553 1049 12565 1057
rect 12565 1049 12599 1057
rect 12599 1049 12605 1057
rect 10416 1023 10423 1031
rect 10423 1023 10457 1031
rect 10457 1023 10468 1031
rect 10416 979 10468 1023
rect 11121 1023 11130 1031
rect 11130 1023 11164 1031
rect 11164 1023 11173 1031
rect 11121 979 11173 1023
rect 11851 1023 11860 1031
rect 11860 1023 11894 1031
rect 11894 1023 11903 1031
rect 11851 979 11903 1023
rect 12553 1023 12565 1031
rect 12565 1023 12599 1031
rect 12599 1023 12605 1031
rect 12553 979 12605 1023
rect 10416 944 10423 961
rect 10423 944 10457 961
rect 10457 944 10468 961
rect 10416 909 10468 944
rect 11121 944 11130 961
rect 11130 944 11164 961
rect 11164 944 11173 961
rect 11121 909 11173 944
rect 11851 944 11860 961
rect 11860 944 11894 961
rect 11894 944 11903 961
rect 11851 909 11903 944
rect 12553 944 12565 961
rect 12565 944 12599 961
rect 12599 944 12605 961
rect 12553 909 12605 944
rect 10416 865 10423 891
rect 10423 865 10457 891
rect 10457 865 10468 891
rect 10416 839 10468 865
rect 11121 865 11130 891
rect 11130 865 11164 891
rect 11164 865 11173 891
rect 11121 839 11173 865
rect 11851 865 11860 891
rect 11860 865 11894 891
rect 11894 865 11903 891
rect 11851 839 11903 865
rect 12553 865 12565 891
rect 12565 865 12599 891
rect 12599 865 12605 891
rect 12553 839 12605 865
rect 10416 820 10468 822
rect 10416 786 10423 820
rect 10423 786 10457 820
rect 10457 786 10468 820
rect 10416 770 10468 786
rect 11121 820 11173 822
rect 11121 786 11130 820
rect 11130 786 11164 820
rect 11164 786 11173 820
rect 11121 770 11173 786
rect 11851 820 11903 822
rect 11851 786 11860 820
rect 11860 786 11894 820
rect 11894 786 11903 820
rect 11851 770 11903 786
rect 12553 820 12605 822
rect 12553 786 12565 820
rect 12565 786 12599 820
rect 12599 786 12605 820
rect 12553 770 12605 786
rect 10416 741 10468 753
rect 10416 707 10423 741
rect 10423 707 10457 741
rect 10457 707 10468 741
rect 10416 701 10468 707
rect 11121 741 11173 753
rect 11121 707 11130 741
rect 11130 707 11164 741
rect 11164 707 11173 741
rect 11121 701 11173 707
rect 11851 741 11903 753
rect 11851 707 11860 741
rect 11860 707 11894 741
rect 11894 707 11903 741
rect 11851 701 11903 707
rect 12553 741 12605 753
rect 12553 707 12565 741
rect 12565 707 12599 741
rect 12599 707 12605 741
rect 12553 701 12605 707
rect 12661 1370 12713 1390
rect 12661 1349 12713 1357
rect 12661 1315 12675 1349
rect 12675 1315 12709 1349
rect 12709 1315 12713 1349
rect 12661 1305 12713 1315
rect 12661 1274 12713 1292
rect 12661 1240 12675 1274
rect 12675 1240 12709 1274
rect 12709 1240 12713 1274
rect 12661 1199 12713 1227
rect 12661 1175 12675 1199
rect 12675 1175 12709 1199
rect 12709 1175 12713 1199
rect 12661 1124 12713 1162
rect 12661 1110 12675 1124
rect 12675 1110 12709 1124
rect 12709 1110 12713 1124
rect 12661 1090 12675 1097
rect 12675 1090 12709 1097
rect 12709 1090 12713 1097
rect 12661 1049 12713 1090
rect 12661 1045 12675 1049
rect 12675 1045 12709 1049
rect 12709 1045 12713 1049
rect 12661 1015 12675 1032
rect 12675 1015 12709 1032
rect 12709 1015 12713 1032
rect 12661 980 12713 1015
rect 12661 940 12675 967
rect 12675 940 12709 967
rect 12709 940 12713 967
rect 12661 915 12713 940
rect 12661 899 12713 902
rect 12661 865 12675 899
rect 12675 865 12709 899
rect 12709 865 12713 899
rect 12661 850 12713 865
rect 12661 825 12713 837
rect 12661 791 12675 825
rect 12675 791 12709 825
rect 12709 791 12713 825
rect 12661 785 12713 791
rect 12661 751 12713 772
rect 12661 720 12675 751
rect 12675 720 12709 751
rect 12709 720 12713 751
rect 12661 677 12713 707
rect 12661 655 12675 677
rect 12675 655 12709 677
rect 12709 655 12713 677
rect 10505 587 10557 639
rect 10576 587 10628 639
rect 10647 587 10699 639
rect 10719 587 10771 639
rect 10791 587 10843 639
rect 10863 587 10915 639
rect 10935 587 10987 639
rect 11007 587 11059 639
rect 11965 587 12017 639
rect 12029 587 12081 639
rect 12093 587 12145 639
rect 12157 587 12209 639
rect 12221 587 12273 639
rect 12399 587 12451 639
rect 12500 587 12552 639
rect 12661 603 12713 642
rect 12661 590 12675 603
rect 12675 590 12709 603
rect 12709 590 12713 603
rect 9459 455 9468 471
rect 9468 455 9502 471
rect 9502 455 9511 471
rect 4637 414 4646 448
rect 4646 414 4680 448
rect 4680 414 4689 448
rect 4637 411 4689 414
rect 2032 369 2084 378
rect 2096 369 2148 378
rect 2160 369 2212 378
rect 2032 335 2039 369
rect 2039 335 2079 369
rect 2079 335 2084 369
rect 2096 335 2113 369
rect 2113 335 2148 369
rect 2160 335 2187 369
rect 2187 335 2212 369
rect 2032 326 2084 335
rect 2096 326 2148 335
rect 2160 326 2212 335
rect 2224 369 2276 378
rect 2224 335 2227 369
rect 2227 335 2261 369
rect 2261 335 2276 369
rect 2224 326 2276 335
rect 2288 369 2340 378
rect 2380 369 2432 378
rect 2288 335 2301 369
rect 2301 335 2335 369
rect 2335 335 2340 369
rect 2380 335 2409 369
rect 2409 335 2432 369
rect 2288 326 2340 335
rect 2380 326 2432 335
rect 2444 369 2496 378
rect 2444 335 2449 369
rect 2449 335 2483 369
rect 2483 335 2496 369
rect 2444 326 2496 335
rect 2508 369 2560 378
rect 2508 335 2523 369
rect 2523 335 2557 369
rect 2557 335 2560 369
rect 2508 326 2560 335
rect 2572 369 2624 378
rect 2636 369 2688 378
rect 2700 369 2752 378
rect 2769 369 2821 378
rect 2838 369 2890 378
rect 2907 369 2959 378
rect 2977 369 3029 378
rect 3047 369 3099 378
rect 2572 335 2597 369
rect 2597 335 2624 369
rect 2636 335 2671 369
rect 2671 335 2688 369
rect 2700 335 2705 369
rect 2705 335 2745 369
rect 2745 335 2752 369
rect 2769 335 2779 369
rect 2779 335 2819 369
rect 2819 335 2821 369
rect 2838 335 2853 369
rect 2853 335 2890 369
rect 2907 335 2927 369
rect 2927 335 2959 369
rect 2977 335 3001 369
rect 3001 335 3029 369
rect 3047 335 3075 369
rect 3075 335 3099 369
rect 2572 326 2624 335
rect 2636 326 2688 335
rect 2700 326 2752 335
rect 2769 326 2821 335
rect 2838 326 2890 335
rect 2907 326 2959 335
rect 2977 326 3029 335
rect 3047 326 3099 335
rect 4637 330 4689 351
rect 4637 299 4646 330
rect 4646 299 4680 330
rect 4680 299 4689 330
rect 4829 402 4835 411
rect 4835 402 4869 411
rect 4869 402 4881 411
rect 4829 359 4881 402
rect 4829 294 4835 309
rect 4835 294 4869 309
rect 4869 294 4881 309
rect 4829 257 4881 294
rect 10501 446 10553 498
rect 10573 446 10625 498
rect 10645 446 10697 498
rect 10717 446 10769 498
rect 10789 446 10841 498
rect 10861 446 10913 498
rect 10934 446 10986 498
rect 11007 446 11059 498
rect 11207 489 11259 498
rect 11207 455 11212 489
rect 11212 455 11246 489
rect 11246 455 11259 489
rect 11207 446 11259 455
rect 11273 489 11325 498
rect 11273 455 11287 489
rect 11287 455 11321 489
rect 11321 455 11325 489
rect 11273 446 11325 455
rect 11339 489 11391 498
rect 11405 489 11457 498
rect 11471 489 11523 498
rect 11537 489 11589 498
rect 11603 489 11655 498
rect 11670 489 11722 498
rect 11339 455 11362 489
rect 11362 455 11391 489
rect 11405 455 11437 489
rect 11437 455 11457 489
rect 11471 455 11512 489
rect 11512 455 11523 489
rect 11537 455 11546 489
rect 11546 455 11587 489
rect 11587 455 11589 489
rect 11603 455 11621 489
rect 11621 455 11655 489
rect 11670 455 11696 489
rect 11696 455 11722 489
rect 11339 446 11391 455
rect 11405 446 11457 455
rect 11471 446 11523 455
rect 11537 446 11589 455
rect 11603 446 11655 455
rect 11670 446 11722 455
rect 11737 489 11789 498
rect 11965 489 12017 498
rect 11737 455 11771 489
rect 11771 455 11789 489
rect 11965 455 11996 489
rect 11996 455 12017 489
rect 11737 446 11789 455
rect 11965 446 12017 455
rect 12029 489 12081 498
rect 12029 455 12037 489
rect 12037 455 12071 489
rect 12071 455 12081 489
rect 12029 446 12081 455
rect 12093 489 12145 498
rect 12157 489 12209 498
rect 12221 489 12273 498
rect 12399 489 12451 498
rect 12500 489 12552 498
rect 12093 455 12112 489
rect 12112 455 12145 489
rect 12157 455 12187 489
rect 12187 455 12209 489
rect 12221 455 12262 489
rect 12262 455 12273 489
rect 12399 455 12412 489
rect 12412 455 12446 489
rect 12446 455 12451 489
rect 12500 455 12521 489
rect 12521 455 12552 489
rect 12093 446 12145 455
rect 12157 446 12209 455
rect 12221 446 12273 455
rect 12399 446 12451 455
rect 12500 446 12552 455
rect 9459 437 9468 440
rect 9468 437 9502 440
rect 9502 437 9511 440
rect 9459 398 9511 437
rect 9459 388 9468 398
rect 9468 388 9502 398
rect 9502 388 9511 398
rect 9459 364 9468 373
rect 9468 364 9502 373
rect 9502 364 9511 373
rect 9459 325 9511 364
rect 9459 321 9468 325
rect 9468 321 9502 325
rect 9502 321 9511 325
rect 5034 245 5086 253
rect 5107 245 5159 253
rect 5180 245 5232 253
rect 5253 245 5305 253
rect 5838 245 5890 253
rect 5902 245 5954 253
rect 5966 245 6018 253
rect 6142 245 6194 253
rect 5034 211 5063 245
rect 5063 211 5086 245
rect 5107 211 5136 245
rect 5136 211 5159 245
rect 5180 211 5209 245
rect 5209 211 5232 245
rect 5253 211 5282 245
rect 5282 211 5305 245
rect 5838 211 5862 245
rect 5862 211 5890 245
rect 5902 211 5934 245
rect 5934 211 5954 245
rect 5966 211 5968 245
rect 5968 211 6006 245
rect 6006 211 6018 245
rect 6142 211 6150 245
rect 6150 211 6184 245
rect 6184 211 6194 245
rect 5034 201 5086 211
rect 5107 201 5159 211
rect 5180 201 5232 211
rect 5253 201 5305 211
rect 5838 201 5890 211
rect 5902 201 5954 211
rect 5966 201 6018 211
rect 6142 201 6194 211
rect 6211 245 6263 253
rect 6211 211 6222 245
rect 6222 211 6256 245
rect 6256 211 6263 245
rect 6211 201 6263 211
rect 6281 245 6333 253
rect 6281 211 6294 245
rect 6294 211 6328 245
rect 6328 211 6333 245
rect 6281 201 6333 211
rect 6351 245 6403 253
rect 6351 211 6366 245
rect 6366 211 6400 245
rect 6400 211 6403 245
rect 6351 201 6403 211
rect 6421 245 6473 253
rect 7505 245 7557 253
rect 6421 211 6438 245
rect 6438 211 6472 245
rect 6472 211 6473 245
rect 7505 211 7518 245
rect 7518 211 7552 245
rect 7552 211 7557 245
rect 6421 201 6473 211
rect 7505 201 7557 211
rect 7577 245 7629 253
rect 7577 211 7590 245
rect 7590 211 7624 245
rect 7624 211 7629 245
rect 7577 201 7629 211
rect 7649 245 7701 253
rect 7649 211 7662 245
rect 7662 211 7696 245
rect 7696 211 7701 245
rect 7649 201 7701 211
rect 7721 245 7773 253
rect 7721 211 7734 245
rect 7734 211 7768 245
rect 7768 211 7773 245
rect 7721 201 7773 211
rect 7793 245 7845 253
rect 7793 211 7806 245
rect 7806 211 7840 245
rect 7840 211 7845 245
rect 7793 201 7845 211
rect 7866 245 7918 253
rect 7866 211 7878 245
rect 7878 211 7912 245
rect 7912 211 7918 245
rect 7866 201 7918 211
rect 7939 245 7991 253
rect 7939 211 7950 245
rect 7950 211 7984 245
rect 7984 211 7991 245
rect 7939 201 7991 211
rect 8012 245 8064 253
rect 8187 245 8239 253
rect 8254 245 8306 253
rect 8322 245 8374 253
rect 8390 245 8442 253
rect 8953 245 9005 253
rect 9033 245 9085 253
rect 9114 245 9166 253
rect 8012 211 8022 245
rect 8022 211 8056 245
rect 8056 211 8064 245
rect 8187 211 8200 245
rect 8200 211 8238 245
rect 8238 211 8239 245
rect 8254 211 8272 245
rect 8272 211 8306 245
rect 8322 211 8344 245
rect 8344 211 8374 245
rect 8390 211 8416 245
rect 8416 211 8442 245
rect 8953 211 8958 245
rect 8958 211 8992 245
rect 8992 211 9005 245
rect 9033 211 9064 245
rect 9064 211 9085 245
rect 9114 211 9136 245
rect 9136 211 9166 245
rect 10086 281 10138 287
rect 10086 247 10090 281
rect 10090 247 10124 281
rect 10124 247 10138 281
rect 10086 235 10138 247
rect 10150 281 10202 287
rect 10150 247 10162 281
rect 10162 247 10196 281
rect 10196 247 10202 281
rect 10150 235 10202 247
rect 10461 281 10513 287
rect 10461 247 10467 281
rect 10467 247 10501 281
rect 10501 247 10513 281
rect 10461 235 10513 247
rect 10525 281 10577 287
rect 10525 247 10539 281
rect 10539 247 10573 281
rect 10573 247 10577 281
rect 10525 235 10577 247
rect 8012 201 8064 211
rect 8187 201 8239 211
rect 8254 201 8306 211
rect 8322 201 8374 211
rect 8390 201 8442 211
rect 8953 201 9005 211
rect 9033 201 9085 211
rect 9114 201 9166 211
rect 4755 117 4807 169
rect 4819 117 4871 169
rect 8484 117 8536 169
rect 8548 117 8600 169
rect 8676 117 8728 169
rect 8740 117 8792 169
rect 5383 33 5435 85
rect 5447 33 5499 85
rect 11840 267 11892 276
rect 11840 233 11846 267
rect 11846 233 11880 267
rect 11880 233 11892 267
rect 11840 224 11892 233
rect 11917 267 11969 276
rect 11917 233 11925 267
rect 11925 233 11959 267
rect 11959 233 11969 267
rect 11917 224 11969 233
rect 11994 267 12046 276
rect 11994 233 12004 267
rect 12004 233 12038 267
rect 12038 233 12046 267
rect 11994 224 12046 233
rect 12070 267 12122 276
rect 12070 233 12082 267
rect 12082 233 12116 267
rect 12116 233 12122 267
rect 12070 224 12122 233
rect 10086 -51 10138 1
rect 10150 -51 10202 1
rect 4667 -135 4719 -83
rect 4743 -135 4795 -83
rect 6842 -106 6894 -54
rect 6906 -106 6958 -54
rect 7974 -106 8026 -54
rect 8038 -106 8090 -54
rect 10461 -135 10513 -83
rect 10525 -135 10577 -83
<< metal2 >>
rect 10102 13224 10154 13230
rect 2379 13188 2431 13194
rect 2379 13124 2431 13136
tri 2344 11113 2379 11148 se
rect 2379 11113 2431 13072
rect 2471 13188 2523 13194
rect 2471 13124 2523 13136
rect 10102 13160 10154 13172
rect 2471 11679 2523 13072
rect 2471 11615 2523 11627
rect 2471 11557 2523 11563
rect 6152 13067 6204 13073
rect 6152 13001 6204 13015
rect 6152 12935 6204 12949
rect 6152 12869 6204 12883
rect 6152 12803 6204 12817
rect 6152 12737 6204 12751
rect 6152 12671 6204 12685
rect 6152 12605 6204 12619
rect 6152 12539 6204 12553
rect 6152 12473 6204 12487
rect 6152 12407 6204 12421
rect 6152 12341 6204 12355
rect 6152 12275 6204 12289
rect 6152 12209 6204 12223
rect 6152 12143 6204 12157
rect 6152 12077 6204 12091
rect 6152 12011 6204 12025
rect 6152 11945 6204 11959
rect 6152 11879 6204 11893
rect 6152 11813 6204 11827
rect 6152 11747 6204 11761
rect 6152 11681 6204 11695
rect 6152 11615 6204 11629
rect 6152 11549 6204 11563
rect 6152 11483 6204 11497
rect 6152 11417 6204 11431
tri 10081 12780 10102 12801 se
rect 10102 12780 10154 13108
rect 10081 12779 10154 12780
rect 10081 11385 10133 12779
tri 10133 12758 10154 12779 nw
tri 10081 11383 10083 11385 ne
rect 10083 11383 10133 11385
tri 10133 11383 10157 11407 sw
rect 6152 11351 6204 11365
tri 10083 11333 10133 11383 ne
rect 10133 11333 10157 11383
tri 10133 11325 10141 11333 ne
rect 10141 11325 10157 11333
tri 10157 11325 10215 11383 sw
tri 10141 11309 10157 11325 ne
rect 10157 11309 10215 11325
tri 10215 11309 10231 11325 sw
rect 6152 11284 6204 11299
tri 10157 11273 10193 11309 ne
rect 10193 11273 10231 11309
tri 10231 11273 10267 11309 sw
rect 11260 11273 11266 11325
rect 11318 11273 11330 11325
rect 11382 11273 11388 11325
tri 10193 11235 10231 11273 ne
rect 10231 11235 10267 11273
tri 10267 11235 10305 11273 sw
tri 11260 11236 11297 11273 ne
rect 6152 11217 6204 11232
rect 6152 11159 6204 11165
tri 10231 11161 10305 11235 ne
tri 10305 11161 10379 11235 sw
tri 10305 11159 10307 11161 ne
rect 10307 11159 10379 11161
tri 10307 11148 10318 11159 ne
rect 10318 11148 10379 11159
tri 2431 11113 2466 11148 sw
tri 10318 11142 10324 11148 ne
rect 10324 11142 10379 11148
rect 2344 11061 2350 11113
rect 2402 11061 2414 11113
rect 2466 11061 2472 11113
rect 7062 10965 7068 11017
rect 7120 10965 7144 11017
rect 7196 10965 7220 11017
rect 7272 10965 7296 11017
rect 7348 10965 7372 11017
rect 7424 10965 7447 11017
rect 7499 10965 7505 11017
rect 7062 10953 7505 10965
rect 4983 10809 5175 10916
rect 7062 10901 7068 10953
rect 7120 10901 7144 10953
rect 7196 10901 7220 10953
rect 7272 10901 7296 10953
rect 7348 10901 7372 10953
rect 7424 10901 7447 10953
rect 7499 10901 7505 10953
tri 4983 10724 5068 10809 ne
rect 5068 10724 5175 10809
tri 5175 10724 5339 10888 sw
tri 5068 10678 5114 10724 ne
rect 5114 10678 5339 10724
rect 326 10672 378 10678
rect 326 10608 378 10620
tri 5114 10617 5175 10678 ne
rect 5175 10617 5339 10678
tri 320 8928 326 8934 se
rect 326 8928 378 10556
tri 5175 10512 5280 10617 ne
rect 5280 10512 5339 10617
tri 5339 10512 5551 10724 sw
tri 304 8912 320 8928 se
rect 320 8912 378 8928
tri 268 8876 304 8912 se
rect 304 8876 342 8912
tri 342 8876 378 8912 nw
tri 264 8872 268 8876 se
rect 268 8872 338 8876
tri 338 8872 342 8876 nw
tri 212 8820 264 8872 se
tri 178 7849 212 7883 se
rect 212 7849 264 8820
tri 264 8798 338 8872 nw
tri 264 7849 275 7860 sw
rect 147 7797 153 7849
rect 205 7797 217 7849
rect 269 7797 275 7849
rect 878 7797 884 7849
rect 936 7797 948 7849
rect 1000 7797 1006 7849
rect -87 6233 -35 6239
tri 306 6221 321 6236 se
rect 321 6221 821 6315
rect -87 6169 -35 6181
tri 254 6169 306 6221 se
rect 306 6169 821 6221
tri 248 6163 254 6169 se
rect 254 6163 821 6169
rect -87 6111 -35 6117
tri 244 6159 248 6163 se
rect 248 6159 821 6163
rect 244 6153 821 6159
rect 296 6146 766 6153
rect 296 6101 445 6146
rect 244 6094 445 6101
rect 497 6094 509 6146
rect 561 6094 573 6146
rect 625 6101 766 6146
rect 818 6101 821 6153
rect 625 6094 821 6101
rect 244 6086 821 6094
rect 296 6073 821 6086
rect 296 6034 766 6073
rect 244 6021 766 6034
rect 818 6021 821 6073
rect 244 6019 821 6021
rect 296 5967 821 6019
rect 244 5952 821 5967
rect 296 5900 821 5952
rect 878 6044 930 7797
tri 930 7763 964 7797 nw
rect 878 5979 930 5992
rect 878 5921 930 5927
rect 958 6150 1010 6315
rect 958 6068 1010 6098
rect 244 5887 821 5900
rect 244 5885 769 5887
rect 296 5835 769 5885
rect 296 5833 821 5835
rect 244 5818 821 5833
rect 296 5795 821 5818
rect 296 5794 769 5795
rect 296 5766 445 5794
rect 244 5751 445 5766
rect 296 5742 445 5751
rect 497 5742 509 5794
rect 561 5742 573 5794
rect 625 5743 769 5794
rect 625 5742 821 5743
rect 296 5703 821 5742
rect 296 5699 769 5703
rect 244 5684 769 5699
rect 296 5651 769 5684
rect 296 5632 821 5651
rect 244 5617 821 5632
rect 296 5565 821 5617
rect 244 5550 821 5565
rect 296 5532 821 5550
rect 296 5498 769 5532
rect 244 5484 769 5498
rect 296 5480 769 5484
rect 296 5467 821 5480
rect 296 5442 769 5467
rect 296 5432 445 5442
rect 160 5402 212 5408
rect 160 5338 212 5350
rect 160 215 212 5286
rect 244 5390 445 5432
rect 497 5390 509 5442
rect 561 5390 573 5442
rect 625 5415 769 5442
rect 625 5403 821 5415
rect 625 5390 769 5403
rect 244 5351 769 5390
rect 244 5339 821 5351
rect 244 5287 769 5339
rect 244 5275 821 5287
rect 244 5223 769 5275
rect 244 5196 821 5223
rect 244 5189 814 5196
tri 814 5189 821 5196 nw
rect 958 5887 1010 6016
rect 958 5795 1010 5835
rect 958 5703 1010 5743
rect 958 5453 1010 5651
rect 1124 6146 1443 6315
rect 1124 6094 1156 6146
rect 1208 6094 1225 6146
rect 1277 6094 1294 6146
rect 1346 6094 1443 6146
rect 1124 5794 1443 6094
rect 1124 5742 1156 5794
rect 1208 5742 1225 5794
rect 1277 5742 1294 5794
rect 1346 5742 1443 5794
rect 958 5382 1010 5401
rect 958 5311 1010 5330
rect 958 5241 1010 5259
rect 244 5171 796 5189
tri 796 5171 814 5189 nw
rect 958 5171 1010 5189
rect 244 5119 744 5171
tri 744 5119 796 5171 nw
rect 244 5107 732 5119
tri 732 5107 744 5119 nw
rect 244 5101 726 5107
tri 726 5101 732 5107 nw
rect 958 5101 1010 5119
rect 296 5090 715 5101
tri 715 5090 726 5101 nw
rect 296 5049 445 5090
rect 244 5038 445 5049
rect 497 5038 509 5090
rect 561 5038 573 5090
rect 625 5049 674 5090
tri 674 5049 715 5090 nw
rect 625 5043 668 5049
tri 668 5043 674 5049 nw
rect 625 5038 663 5043
tri 663 5038 668 5043 nw
rect 244 5033 641 5038
rect 296 5016 641 5033
tri 641 5016 663 5038 nw
rect 296 4981 640 5016
tri 640 5015 641 5016 nw
rect 244 4965 640 4981
rect 296 4913 640 4965
rect 693 4931 699 4983
rect 751 4931 763 4983
rect 815 4931 821 4983
rect 244 4897 640 4913
tri 744 4906 769 4931 ne
rect 296 4845 640 4897
rect 244 4829 640 4845
rect 296 4824 640 4829
rect 296 4777 445 4824
rect 244 4772 445 4777
rect 497 4772 509 4824
rect 561 4772 573 4824
rect 625 4772 640 4824
rect 244 4761 640 4772
rect 296 4709 640 4761
rect 244 4693 640 4709
rect 296 4641 640 4693
rect 244 4625 640 4641
rect 296 4573 640 4625
rect 244 4557 640 4573
rect 296 4551 640 4557
rect 296 4505 409 4551
rect 244 4499 409 4505
rect 461 4499 495 4551
rect 547 4499 582 4551
rect 634 4499 640 4551
rect 687 4741 739 4747
rect 687 4677 739 4689
rect 240 3494 292 3500
rect 240 3430 292 3442
rect 240 2977 292 3378
rect 240 2913 292 2925
rect 240 2030 292 2861
rect 240 1966 292 1978
rect 240 1908 292 1914
rect 321 3200 445 3252
rect 497 3200 509 3252
rect 561 3200 573 3252
rect 625 3200 640 3252
rect 321 2866 640 3200
rect 321 2814 429 2866
rect 481 2814 493 2866
rect 545 2814 640 2866
rect 321 2682 640 2814
rect 321 2630 445 2682
rect 497 2630 509 2682
rect 561 2630 573 2682
rect 625 2630 640 2682
rect 321 2416 640 2630
rect 321 2364 445 2416
rect 497 2364 509 2416
rect 561 2364 573 2416
rect 625 2364 640 2416
rect 321 2038 640 2364
rect 321 1986 335 2038
rect 387 1986 399 2038
rect 451 1986 463 2038
rect 515 1986 640 2038
rect 241 1736 293 1742
rect 241 1663 293 1684
rect 241 1591 293 1611
rect 241 1519 293 1539
rect 241 1447 293 1467
rect 241 1375 293 1395
rect 241 1303 293 1323
rect 321 1255 640 1986
rect 687 1382 739 4625
rect 687 1318 739 1330
rect 687 1260 739 1266
rect 769 3666 821 4931
rect 769 3602 821 3614
rect 241 1231 293 1251
rect 241 867 293 1179
rect 241 801 293 815
rect 241 735 293 749
rect 241 669 293 683
rect 241 602 293 617
rect 241 535 293 550
rect 241 468 293 483
rect 241 401 293 416
rect 241 329 293 349
rect 321 1147 445 1199
rect 497 1147 509 1199
rect 561 1147 573 1199
rect 625 1147 640 1199
rect 321 847 640 1147
rect 321 795 445 847
rect 497 795 509 847
rect 561 795 573 847
rect 625 795 640 847
rect 321 628 640 795
rect 769 1096 821 3550
rect 849 4799 901 4805
rect 849 4735 901 4747
rect 849 4095 901 4683
rect 849 4031 901 4043
rect 849 3967 901 3979
rect 849 3325 901 3915
rect 849 3261 901 3273
rect 849 3203 901 3209
rect 958 4641 1010 5049
rect 958 4565 1010 4589
rect 958 4490 1010 4513
rect 958 4415 1010 4438
rect 958 4340 1010 4363
rect 958 4265 1010 4288
rect 958 3865 1010 4213
rect 958 3792 1010 3813
rect 958 3720 1010 3740
rect 958 3648 1010 3668
rect 958 3576 1010 3596
rect 958 3504 1010 3524
rect 849 3041 901 3047
rect 849 2977 901 2989
rect 849 2177 901 2925
rect 849 2113 901 2125
rect 849 2055 901 2061
rect 958 2925 1010 3452
rect 958 2720 1010 2873
rect 958 2646 1010 2668
rect 958 2572 1010 2594
rect 958 2498 1010 2520
rect 1043 5535 1095 5541
rect 1043 5471 1095 5483
rect 1043 2570 1095 5419
rect 1043 2504 1095 2518
rect 1043 2446 1095 2452
rect 1124 5252 1443 5742
rect 1124 5200 1221 5252
rect 1273 5200 1285 5252
rect 1337 5200 1443 5252
rect 1124 3811 1443 5200
rect 1124 3759 1156 3811
rect 1208 3759 1220 3811
rect 1272 3759 1284 3811
rect 1336 3759 1443 3811
rect 1124 3633 1443 3759
rect 1124 3581 1156 3633
rect 1208 3581 1220 3633
rect 1272 3581 1284 3633
rect 1336 3581 1443 3633
rect 1124 3464 1443 3581
rect 1124 3412 1156 3464
rect 1208 3412 1220 3464
rect 1272 3412 1284 3464
rect 1336 3412 1443 3464
rect 1124 3216 1443 3412
rect 1124 3164 1156 3216
rect 1208 3164 1220 3216
rect 1272 3164 1284 3216
rect 1336 3164 1443 3216
rect 1124 2922 1443 3164
rect 1124 2870 1156 2922
rect 1208 2870 1220 2922
rect 1272 2870 1284 2922
rect 1336 2870 1443 2922
rect 1124 2720 1443 2870
rect 1124 2668 1156 2720
rect 1208 2668 1220 2720
rect 1272 2668 1284 2720
rect 1336 2668 1443 2720
rect 1124 2536 1443 2668
rect 1124 2484 1156 2536
rect 1208 2484 1220 2536
rect 1272 2484 1284 2536
rect 1336 2484 1443 2536
rect 958 2424 1010 2446
rect 958 2351 1010 2372
rect 769 1032 821 1044
rect 769 744 821 980
rect 769 680 821 692
tri 640 628 680 668 sw
rect 321 622 680 628
tri 680 622 686 628 sw
rect 769 622 821 628
rect 849 2021 901 2027
rect 849 1957 901 1969
rect 849 1564 901 1905
rect 849 1500 901 1512
rect 849 744 901 1448
rect 849 680 901 692
rect 958 1944 1010 2299
rect 1124 2352 1443 2484
rect 1124 2300 1156 2352
rect 1208 2300 1220 2352
rect 1272 2300 1284 2352
rect 1336 2300 1443 2352
rect 958 1879 1010 1892
rect 958 1814 1010 1827
rect 958 1749 1010 1762
rect 958 1684 1010 1697
rect 958 1620 1010 1632
rect 958 1556 1010 1568
rect 958 1406 1010 1504
rect 958 1333 1010 1354
rect 958 1112 1010 1281
rect 958 1042 1010 1060
rect 958 876 1010 990
rect 1043 2235 1095 2241
rect 1043 2169 1095 2183
rect 1043 1042 1095 2117
rect 1043 976 1095 990
rect 1043 915 1095 924
rect 1124 2168 1443 2300
rect 1124 2116 1156 2168
rect 1208 2116 1220 2168
rect 1272 2116 1284 2168
rect 1336 2116 1443 2168
rect 1124 1917 1443 2116
rect 1124 1865 1156 1917
rect 1208 1865 1220 1917
rect 1272 1865 1284 1917
rect 1336 1865 1443 1917
rect 1124 1748 1443 1865
rect 1124 1696 1156 1748
rect 1208 1696 1220 1748
rect 1272 1696 1284 1748
rect 1336 1696 1443 1748
rect 1124 1570 1443 1696
rect 1124 1518 1156 1570
rect 1208 1518 1220 1570
rect 1272 1518 1284 1570
rect 1336 1518 1443 1570
rect 958 808 1010 824
rect 958 740 1010 756
rect 958 682 1010 688
tri 1116 660 1124 668 se
rect 1124 660 1443 1518
rect 849 622 901 628
tri 1078 622 1116 660 se
rect 1116 622 1443 660
rect 321 608 686 622
tri 686 608 700 622 sw
tri 1064 608 1078 622 se
rect 1078 608 1443 622
rect 321 596 700 608
tri 700 596 712 608 sw
tri 1052 596 1064 608 se
rect 1064 596 1443 608
rect 321 544 712 596
tri 712 544 764 596 sw
tri 1000 544 1052 596 se
rect 1052 544 1443 596
rect 321 532 764 544
tri 764 532 776 544 sw
tri 988 532 1000 544 se
rect 1000 532 1443 544
rect 321 526 776 532
tri 776 526 782 532 sw
tri 982 526 988 532 se
rect 988 526 1443 532
rect 321 495 1443 526
rect 321 443 433 495
rect 485 443 497 495
rect 549 443 561 495
rect 613 443 1443 495
rect 321 326 1443 443
rect 1471 6150 1523 6315
rect 1471 6085 1523 6098
rect 1471 6020 1523 6033
rect 1471 5955 1523 5968
rect 1471 5890 1523 5903
rect 1471 5825 1523 5838
rect 1471 5759 1523 5773
rect 1471 5693 1523 5707
rect 1471 5627 1523 5641
rect 1471 5458 1523 5575
rect 1471 5393 1523 5406
rect 1471 5328 1523 5341
rect 1471 5263 1523 5276
rect 1471 5198 1523 5211
rect 1471 5133 1523 5146
rect 1471 5068 1523 5081
rect 1471 5003 1523 5016
rect 1471 4938 1523 4951
rect 1471 4873 1523 4886
rect 1471 4808 1523 4821
rect 1471 4743 1523 4756
rect 1471 4678 1523 4691
rect 1471 4613 1523 4626
rect 1471 4548 1523 4561
rect 1471 4483 1523 4496
rect 1471 4418 1523 4431
rect 1471 4353 1523 4366
rect 1471 4287 1523 4301
rect 1471 4221 1523 4235
rect 1471 4155 1523 4169
rect 1471 4089 1523 4103
rect 1471 4023 1523 4037
rect 1471 3957 1523 3971
rect 1471 3891 1523 3905
rect 1471 3825 1523 3839
rect 1471 3759 1523 3773
rect 1471 3693 1523 3707
rect 1471 3627 1523 3641
rect 1471 3561 1523 3575
rect 1471 3495 1523 3509
rect 1471 3429 1523 3443
rect 1471 3363 1523 3377
rect 1471 3297 1523 3311
rect 1471 3231 1523 3245
rect 1471 3165 1523 3179
rect 1471 3099 1523 3113
rect 1471 3033 1523 3047
rect 1471 2967 1523 2981
rect 1471 2901 1523 2915
rect 1471 2687 1523 2849
rect 1471 2580 1523 2635
rect 1471 2399 1523 2528
rect 1471 2334 1523 2347
rect 1471 2269 1523 2282
rect 1471 2204 1523 2217
rect 1471 2139 1523 2152
rect 1471 2074 1523 2087
rect 1471 2009 1523 2022
rect 1471 1944 1523 1957
rect 1471 1879 1523 1892
rect 1471 1814 1523 1827
rect 1471 1749 1523 1762
rect 1471 1684 1523 1697
rect 1471 1620 1523 1632
rect 1471 1556 1523 1568
rect 1471 1492 1523 1504
rect 1471 1428 1523 1440
rect 1471 1364 1523 1376
rect 1471 1300 1523 1312
rect 1471 1236 1523 1248
rect 1471 1172 1523 1184
rect 1471 1108 1523 1120
rect 1471 1044 1523 1056
rect 1471 980 1523 992
rect 1471 916 1523 928
rect 1471 852 1523 864
rect 1471 788 1523 800
rect 1471 724 1523 736
rect 1471 660 1523 672
rect 1471 596 1523 608
rect 1471 532 1523 544
rect 1471 468 1523 480
rect 1471 404 1523 416
rect 1471 329 1523 352
rect 1551 -139 1721 6054
rect 1749 5510 1918 5516
rect 1749 5330 1769 5510
rect 1885 5330 1918 5510
rect 1749 -139 1918 5330
rect 1946 4952 1998 6315
rect 2750 5516 2802 6298
rect 1946 4868 1998 4900
rect 1946 4785 1998 4816
rect 1946 4702 1998 4733
rect 1946 4644 1998 4650
rect 2026 5055 2346 5505
rect 2026 5003 2032 5055
rect 2084 5003 2096 5055
rect 2148 5003 2160 5055
rect 2212 5003 2224 5055
rect 2276 5003 2288 5055
rect 2340 5003 2346 5055
rect 2026 4599 2346 5003
rect 2026 4547 2032 4599
rect 2084 4547 2096 4599
rect 2148 4547 2160 4599
rect 2212 4547 2224 4599
rect 2276 4547 2288 4599
rect 2340 4547 2346 4599
rect 2026 4143 2346 4547
rect 2026 4091 2032 4143
rect 2084 4091 2096 4143
rect 2148 4091 2160 4143
rect 2212 4091 2224 4143
rect 2276 4091 2288 4143
rect 2340 4091 2346 4143
rect 2026 3687 2346 4091
rect 2026 3635 2032 3687
rect 2084 3635 2096 3687
rect 2148 3635 2160 3687
rect 2212 3635 2224 3687
rect 2276 3635 2288 3687
rect 2340 3635 2346 3687
rect 2026 3231 2346 3635
rect 2026 3179 2032 3231
rect 2084 3179 2096 3231
rect 2148 3179 2160 3231
rect 2212 3179 2224 3231
rect 2276 3179 2288 3231
rect 2340 3179 2346 3231
rect 2026 2775 2346 3179
rect 2026 2723 2032 2775
rect 2084 2723 2096 2775
rect 2148 2723 2160 2775
rect 2212 2723 2224 2775
rect 2276 2723 2288 2775
rect 2340 2723 2346 2775
rect 2026 2319 2346 2723
rect 2026 2267 2032 2319
rect 2084 2267 2096 2319
rect 2148 2267 2160 2319
rect 2212 2267 2224 2319
rect 2276 2267 2288 2319
rect 2340 2267 2346 2319
rect 2026 1863 2346 2267
rect 2026 1811 2032 1863
rect 2084 1811 2096 1863
rect 2148 1811 2160 1863
rect 2212 1811 2224 1863
rect 2276 1811 2288 1863
rect 2340 1811 2346 1863
rect 2026 1407 2346 1811
rect 2026 1355 2032 1407
rect 2084 1355 2096 1407
rect 2148 1355 2160 1407
rect 2212 1355 2224 1407
rect 2276 1355 2288 1407
rect 2340 1355 2346 1407
rect 2026 951 2346 1355
rect 2026 899 2032 951
rect 2084 899 2096 951
rect 2148 899 2160 951
rect 2212 899 2224 951
rect 2276 899 2288 951
rect 2340 899 2346 951
rect 2026 495 2346 899
rect 2026 443 2032 495
rect 2084 443 2096 495
rect 2148 443 2160 495
rect 2212 443 2224 495
rect 2276 443 2288 495
rect 2340 443 2346 495
rect 2026 378 2346 443
rect 2026 326 2032 378
rect 2084 326 2096 378
rect 2148 326 2160 378
rect 2212 326 2224 378
rect 2276 326 2288 378
rect 2340 326 2346 378
rect 2374 5025 2694 5505
rect 2374 4973 2572 5025
rect 2624 4973 2636 5025
rect 2688 4973 2694 5025
rect 2374 4569 2694 4973
rect 2374 4517 2572 4569
rect 2624 4517 2636 4569
rect 2688 4517 2694 4569
rect 2374 3229 2694 4517
rect 2374 2307 2427 3229
tri 2427 3204 2452 3229 nw
tri 2541 3204 2566 3229 ne
rect 2475 3129 2527 3135
rect 2475 3065 2527 3077
rect 2475 3001 2527 3013
rect 2475 2844 2527 2949
rect 2475 2780 2527 2792
rect 2475 2549 2527 2728
rect 2475 2485 2527 2497
rect 2475 2421 2527 2433
rect 2475 2363 2527 2369
tri 2427 2307 2452 2332 sw
tri 2541 2307 2566 2332 se
rect 2566 2307 2694 3229
rect 2750 5452 2802 5464
rect 2750 3051 2802 5400
rect 2931 6289 2983 6295
rect 2931 6221 2983 6237
rect 2931 5430 2983 6169
rect 3023 6117 3075 6123
rect 3023 6049 3075 6065
rect 3023 5656 3075 5997
rect 3023 5592 3075 5604
rect 3023 5534 3075 5540
tri 2983 5430 3008 5455 sw
rect 2931 5378 2937 5430
rect 2989 5378 3005 5430
rect 3057 5378 3063 5430
rect 2830 5295 2836 5347
rect 2888 5295 2900 5347
rect 2952 5295 2958 5347
rect 2830 5283 2920 5295
tri 2920 5283 2932 5295 nw
rect 2830 5260 2897 5283
tri 2897 5260 2920 5283 nw
rect 2830 5252 2889 5260
tri 2889 5252 2897 5260 nw
rect 2830 4404 2886 5252
tri 2886 5249 2889 5252 nw
rect 2987 5120 3020 5172
rect 3072 5120 3122 5172
tri 3045 5118 3047 5120 ne
rect 3047 5118 3122 5120
tri 3047 5108 3057 5118 ne
rect 3057 5108 3122 5118
tri 3057 5095 3070 5108 ne
rect 2882 4352 2886 4404
rect 2830 4340 2886 4352
rect 2882 4310 2886 4340
tri 2882 4306 2886 4310 nw
rect 3070 5079 3122 5108
rect 3070 5012 3122 5027
rect 3070 4945 3122 4960
rect 3070 4878 3122 4893
rect 3070 4811 3122 4826
rect 3070 4744 3122 4759
rect 3070 4677 3122 4692
rect 3070 4610 3122 4625
rect 3070 4543 3122 4558
rect 3070 4476 3122 4491
rect 3070 4408 3122 4424
rect 3070 4340 3122 4356
rect 2830 4133 2882 4288
rect 2830 4069 2882 4081
rect 2830 3780 2882 4017
rect 2830 3716 2882 3728
rect 2830 3509 2882 3664
rect 3070 4174 3122 4288
rect 3070 4100 3122 4122
rect 3070 4027 3122 4048
rect 3070 3954 3122 3975
rect 3070 3749 3122 3902
rect 2830 3445 2882 3457
rect 2830 3197 2882 3393
rect 2830 3133 2882 3145
rect 2830 3075 2882 3081
rect 2910 3653 2962 3659
rect 2910 3589 2962 3601
rect 2910 3353 2962 3537
rect 2910 3289 2962 3301
tri 2802 3051 2808 3057 sw
rect 2750 3043 2808 3051
tri 2808 3043 2816 3051 sw
rect 2750 3035 2816 3043
tri 2750 2991 2794 3035 ne
rect 2794 2991 2816 3035
tri 2816 2991 2868 3043 sw
tri 2794 2977 2808 2991 ne
rect 2808 2977 2868 2991
tri 2868 2977 2882 2991 sw
tri 2808 2973 2812 2977 ne
rect 2812 2973 2882 2977
tri 2812 2965 2820 2973 ne
rect 2820 2965 2882 2973
tri 2820 2959 2826 2965 ne
rect 2826 2959 2882 2965
tri 2826 2955 2830 2959 ne
rect 2374 981 2694 2307
rect 2374 929 2572 981
rect 2624 929 2636 981
rect 2688 929 2694 981
rect 2374 525 2694 929
rect 2750 2844 2802 2850
rect 2750 2780 2802 2792
rect 2750 924 2802 2728
rect 2830 2557 2882 2959
rect 2910 2959 2962 3237
rect 3070 3654 3122 3697
rect 3070 3560 3122 3602
rect 3070 3394 3122 3508
rect 3070 3323 3122 3342
rect 3070 3253 3122 3271
rect 3070 3183 3122 3201
rect 3070 3113 3122 3131
rect 3070 3043 3122 3061
rect 3070 2973 3122 2991
rect 2910 2895 2962 2907
rect 2910 2779 2962 2843
rect 2910 2715 2962 2727
rect 2910 2657 2962 2663
rect 2990 2940 3042 2946
rect 2990 2876 3042 2888
rect 2990 2705 3042 2824
rect 2990 2641 3042 2653
tri 2830 2551 2836 2557 ne
rect 2836 2551 2882 2557
tri 2882 2551 2910 2579 sw
tri 2836 2548 2839 2551 ne
rect 2839 2548 2962 2551
tri 2839 2545 2842 2548 ne
rect 2842 2545 2962 2548
tri 2842 2505 2882 2545 ne
rect 2882 2505 2910 2545
tri 2882 2493 2894 2505 ne
rect 2894 2493 2910 2505
tri 2894 2481 2906 2493 ne
rect 2906 2481 2962 2493
tri 2906 2477 2910 2481 ne
rect 2910 2423 2962 2429
rect 2830 2417 2882 2423
rect 2830 2353 2882 2365
rect 2830 2105 2882 2301
rect 2830 2041 2882 2053
rect 2830 1834 2882 1989
rect 2990 2261 3042 2589
rect 2990 2197 3042 2209
rect 2990 1949 3042 2145
rect 2990 1885 3042 1897
rect 2990 1827 3042 1833
rect 3070 2600 3122 2921
rect 3070 2526 3122 2548
rect 3070 2452 3122 2474
rect 3070 2378 3122 2400
rect 3070 2304 3122 2326
rect 3070 2230 3122 2252
rect 3070 2156 3122 2178
rect 3070 1990 3122 2104
rect 3070 1895 3122 1938
rect 2830 1770 2882 1782
rect 2830 1481 2882 1718
rect 2830 1417 2882 1429
rect 2830 1210 2882 1365
rect 2830 1146 2882 1158
rect 2830 996 2882 1094
rect 3070 1801 3122 1843
rect 3070 1596 3122 1749
rect 3070 1522 3122 1544
rect 3070 1449 3122 1470
rect 3070 1376 3122 1397
rect 3070 1210 3122 1324
rect 3070 1138 3122 1158
rect 3070 1067 3122 1086
tri 2882 996 2897 1011 sw
rect 3070 996 3122 1015
rect 2830 985 2897 996
tri 2897 985 2908 996 sw
tri 2830 944 2871 985 ne
rect 2871 953 2908 985
tri 2908 953 2940 985 sw
rect 2871 944 2940 953
tri 2940 944 2949 953 sw
tri 2871 940 2875 944 ne
rect 2875 940 2949 944
tri 2949 940 2953 944 sw
tri 2875 926 2889 940 ne
rect 2889 926 2953 940
tri 2802 924 2804 926 sw
tri 2889 924 2891 926 ne
rect 2891 924 2953 926
tri 2953 924 2969 940 sw
rect 2750 909 2804 924
tri 2804 909 2819 924 sw
tri 2891 909 2906 924 ne
rect 2906 909 2969 924
tri 2969 909 2984 924 sw
rect 2750 901 2819 909
tri 2819 901 2827 909 sw
tri 2906 907 2908 909 ne
rect 2908 907 2984 909
tri 2984 907 2986 909 sw
tri 2908 901 2914 907 ne
rect 2914 901 2986 907
tri 2986 901 2992 907 sw
rect 2750 895 2866 901
rect 2802 843 2814 895
tri 2914 875 2940 901 ne
rect 2750 837 2866 843
rect 2940 828 2992 901
rect 2940 764 2992 776
rect 2940 706 2992 712
rect 2374 473 2572 525
rect 2624 473 2636 525
rect 2688 503 2694 525
rect 3070 701 3122 944
rect 3070 628 3122 649
rect 3070 555 3122 576
tri 2694 503 2712 521 sw
rect 2688 484 2712 503
tri 2712 484 2731 503 sw
rect 2688 482 2731 484
tri 2731 482 2733 484 sw
rect 3070 482 3122 503
rect 2688 473 2733 482
tri 2733 473 2742 482 sw
rect 2374 430 2742 473
tri 2742 430 2785 473 sw
rect 2374 425 2785 430
tri 2785 425 2790 430 sw
rect 2374 411 2790 425
tri 2790 411 2804 425 sw
rect 2374 403 2804 411
tri 2804 403 2812 411 sw
rect 2374 378 2812 403
tri 2812 378 2837 403 sw
tri 3045 378 3070 403 se
rect 3070 378 3122 430
rect 2374 326 2380 378
rect 2432 326 2444 378
rect 2496 326 2508 378
rect 2560 326 2572 378
rect 2624 326 2636 378
rect 2688 326 2700 378
rect 2752 326 2769 378
rect 2821 326 2838 378
rect 2890 326 2907 378
rect 2959 326 2977 378
rect 3029 326 3047 378
rect 3099 326 3122 378
rect 3178 2824 3534 6315
rect 3590 6108 4415 10512
tri 3590 6094 3604 6108 ne
rect 3604 6094 4401 6108
tri 4401 6094 4415 6108 nw
rect 4471 6215 4773 10512
tri 5280 10453 5339 10512 ne
rect 5339 10453 5551 10512
tri 5551 10453 5610 10512 sw
tri 5339 10443 5349 10453 ne
rect 5349 10443 5610 10453
tri 5349 10391 5401 10443 ne
rect 5401 10391 5610 10443
tri 5401 10374 5418 10391 ne
rect 4471 6163 4637 6215
rect 4689 6163 4773 6215
rect 4471 6146 4773 6163
rect 4471 6094 4637 6146
rect 4689 6094 4773 6146
tri 3604 6077 3621 6094 ne
rect 3621 6077 4384 6094
tri 4384 6077 4401 6094 nw
rect 4471 6077 4773 6094
tri 3621 6025 3673 6077 ne
rect 3673 6025 4332 6077
tri 4332 6025 4384 6077 nw
rect 4471 6025 4637 6077
rect 4689 6025 4773 6077
tri 3673 6008 3690 6025 ne
rect 3690 6008 4315 6025
tri 4315 6008 4332 6025 nw
rect 4471 6008 4773 6025
tri 3690 5956 3742 6008 ne
rect 3742 5956 4263 6008
tri 4263 5956 4315 6008 nw
rect 4471 5956 4637 6008
rect 4689 5956 4773 6008
tri 3742 5948 3750 5956 ne
rect 3750 5948 4255 5956
tri 4255 5948 4263 5956 nw
rect 3750 5939 4246 5948
tri 4246 5939 4255 5948 nw
rect 4471 5939 4773 5956
rect 3750 5935 4242 5939
tri 4242 5935 4246 5939 nw
rect 3750 5887 4194 5935
tri 4194 5887 4242 5935 nw
tri 4423 5887 4471 5935 se
rect 4471 5887 4637 5939
rect 4689 5887 4773 5939
rect 3750 5870 4177 5887
tri 4177 5870 4194 5887 nw
tri 4418 5882 4423 5887 se
rect 4423 5882 4773 5887
rect 4418 5870 4773 5882
rect 3750 5818 4125 5870
tri 4125 5818 4177 5870 nw
rect 4418 5818 4637 5870
rect 4689 5818 4773 5870
rect 3750 5801 4108 5818
tri 4108 5801 4125 5818 nw
rect 4418 5809 4773 5818
rect 4418 5801 4717 5809
rect 3590 5260 3642 5266
rect 3590 5192 3642 5208
rect 3590 3018 3642 5140
rect 3590 2950 3642 2966
rect 3590 2892 3642 2898
rect 3750 4790 4070 5801
tri 4070 5763 4108 5801 nw
rect 4418 5749 4637 5801
rect 4689 5749 4717 5801
tri 4717 5753 4773 5809 nw
rect 4825 8517 4831 8569
rect 4883 8517 4895 8569
rect 4947 8517 4953 8569
rect 4418 5731 4717 5749
rect 4418 5679 4637 5731
rect 4689 5679 4717 5731
rect 4118 5200 4124 5252
rect 4176 5200 4188 5252
rect 4240 5200 4310 5252
tri 4233 5183 4250 5200 ne
rect 4250 5183 4310 5200
tri 4250 5178 4255 5183 ne
rect 4255 5178 4310 5183
tri 4255 5175 4258 5178 ne
rect 4258 5108 4310 5178
rect 3750 4738 3884 4790
rect 3936 4738 3948 4790
rect 4000 4738 4012 4790
rect 4064 4738 4070 4790
rect 3750 4389 4070 4738
rect 3750 4337 3884 4389
rect 3936 4337 3948 4389
rect 4000 4337 4012 4389
rect 4064 4337 4070 4389
rect 3750 4073 4070 4337
rect 3750 4021 3884 4073
rect 3936 4021 3948 4073
rect 4000 4021 4012 4073
rect 4064 4021 4070 4073
rect 3750 3763 4070 4021
rect 3750 3711 3884 3763
rect 3936 3711 3948 3763
rect 4000 3711 4012 3763
rect 4064 3711 4070 3763
rect 3750 3359 4070 3711
rect 3750 3307 3884 3359
rect 3936 3307 3948 3359
rect 4000 3307 4012 3359
rect 4064 3307 4070 3359
rect 3750 3155 4070 3307
rect 3750 3103 3884 3155
rect 3936 3103 3948 3155
rect 4000 3103 4012 3155
rect 4064 3103 4070 3155
rect 3750 2959 4070 3103
rect 3750 2907 3884 2959
rect 3936 2907 3948 2959
rect 4000 2907 4012 2959
rect 4064 2907 4070 2959
tri 3534 2824 3580 2870 sw
rect 3178 2822 3580 2824
tri 3580 2822 3582 2824 sw
rect 3178 2818 3582 2822
tri 3582 2818 3586 2822 sw
rect 3178 2809 3586 2818
tri 3586 2809 3595 2818 sw
rect 3178 2807 3595 2809
tri 3595 2807 3597 2809 sw
rect 3178 2795 3597 2807
tri 3597 2795 3609 2807 sw
rect 3178 2755 3609 2795
tri 3609 2755 3649 2795 sw
rect 3178 2752 3649 2755
tri 3649 2752 3652 2755 sw
rect 3178 2748 3652 2752
tri 3652 2748 3656 2752 sw
rect 3178 448 3656 2748
rect 3750 2591 4070 2907
rect 4098 5079 4150 5085
rect 4098 5015 4150 5027
rect 4098 3923 4150 4963
rect 4258 5026 4310 5056
rect 4258 4944 4310 4974
rect 4258 4862 4310 4892
rect 4258 4336 4310 4810
rect 4258 4234 4310 4284
rect 4098 3638 4150 3871
rect 4098 3574 4150 3586
rect 4098 2940 4150 3522
rect 4178 4116 4230 4122
rect 4178 4052 4230 4064
rect 4178 3092 4230 4000
rect 4178 3028 4230 3040
rect 4178 2970 4230 2976
rect 4258 3749 4310 4182
rect 4418 5118 4717 5679
rect 4825 5411 4877 8517
tri 4877 8483 4911 8517 nw
rect 5418 7302 5610 10391
tri 5610 7302 5682 7374 sw
rect 5869 7302 6280 10512
tri 6377 7302 6418 7343 se
rect 6418 7302 6610 10512
rect 7058 10132 7509 10512
rect 7058 10080 7067 10132
rect 7119 10080 7131 10132
rect 7183 10080 7195 10132
rect 7247 10080 7259 10132
rect 7311 10080 7323 10132
rect 7375 10080 7387 10132
rect 7439 10080 7451 10132
rect 7503 10080 7509 10132
rect 7058 10065 7509 10080
rect 7058 10013 7067 10065
rect 7119 10013 7131 10065
rect 7183 10013 7195 10065
rect 7247 10013 7259 10065
rect 7311 10013 7323 10065
rect 7375 10013 7387 10065
rect 7439 10013 7451 10065
rect 7503 10013 7509 10065
rect 7058 9998 7509 10013
rect 7058 9946 7067 9998
rect 7119 9946 7131 9998
rect 7183 9946 7195 9998
rect 7247 9946 7259 9998
rect 7311 9946 7323 9998
rect 7375 9946 7387 9998
rect 7439 9946 7451 9998
rect 7503 9946 7509 9998
rect 7058 9930 7509 9946
rect 7058 9878 7067 9930
rect 7119 9878 7131 9930
rect 7183 9878 7195 9930
rect 7247 9878 7259 9930
rect 7311 9878 7323 9930
rect 7375 9878 7387 9930
rect 7439 9878 7451 9930
rect 7503 9878 7509 9930
rect 7058 9862 7509 9878
rect 7058 9810 7067 9862
rect 7119 9810 7131 9862
rect 7183 9810 7195 9862
rect 7247 9810 7259 9862
rect 7311 9810 7323 9862
rect 7375 9810 7387 9862
rect 7439 9810 7451 9862
rect 7503 9810 7509 9862
rect 7058 9794 7509 9810
rect 7058 9742 7067 9794
rect 7119 9742 7131 9794
rect 7183 9742 7195 9794
rect 7247 9742 7259 9794
rect 7311 9742 7323 9794
rect 7375 9742 7387 9794
rect 7439 9742 7451 9794
rect 7503 9742 7509 9794
rect 7058 9726 7509 9742
rect 7058 9674 7067 9726
rect 7119 9674 7131 9726
rect 7183 9674 7195 9726
rect 7247 9674 7259 9726
rect 7311 9674 7323 9726
rect 7375 9674 7387 9726
rect 7439 9674 7451 9726
rect 7503 9674 7509 9726
rect 7058 9658 7509 9674
rect 7058 9606 7067 9658
rect 7119 9606 7131 9658
rect 7183 9606 7195 9658
rect 7247 9606 7259 9658
rect 7311 9606 7323 9658
rect 7375 9606 7387 9658
rect 7439 9606 7451 9658
rect 7503 9606 7509 9658
rect 7058 9402 7509 9606
rect 7058 9350 7067 9402
rect 7119 9350 7131 9402
rect 7183 9350 7195 9402
rect 7247 9350 7259 9402
rect 7311 9350 7323 9402
rect 7375 9350 7387 9402
rect 7439 9350 7451 9402
rect 7503 9350 7509 9402
rect 7058 9335 7509 9350
rect 7058 9283 7067 9335
rect 7119 9283 7131 9335
rect 7183 9283 7195 9335
rect 7247 9283 7259 9335
rect 7311 9283 7323 9335
rect 7375 9283 7387 9335
rect 7439 9283 7451 9335
rect 7503 9283 7509 9335
rect 7058 9268 7509 9283
rect 7058 9216 7067 9268
rect 7119 9216 7131 9268
rect 7183 9216 7195 9268
rect 7247 9216 7259 9268
rect 7311 9216 7323 9268
rect 7375 9216 7387 9268
rect 7439 9216 7451 9268
rect 7503 9216 7509 9268
rect 7058 9200 7509 9216
rect 7058 9148 7067 9200
rect 7119 9148 7131 9200
rect 7183 9148 7195 9200
rect 7247 9148 7259 9200
rect 7311 9148 7323 9200
rect 7375 9148 7387 9200
rect 7439 9148 7451 9200
rect 7503 9148 7509 9200
rect 7058 9132 7509 9148
rect 7058 9080 7067 9132
rect 7119 9080 7131 9132
rect 7183 9080 7195 9132
rect 7247 9080 7259 9132
rect 7311 9080 7323 9132
rect 7375 9080 7387 9132
rect 7439 9080 7451 9132
rect 7503 9080 7509 9132
rect 7058 9064 7509 9080
rect 7058 9012 7067 9064
rect 7119 9012 7131 9064
rect 7183 9012 7195 9064
rect 7247 9012 7259 9064
rect 7311 9012 7323 9064
rect 7375 9012 7387 9064
rect 7439 9012 7451 9064
rect 7503 9012 7509 9064
rect 7058 8996 7509 9012
rect 7058 8944 7067 8996
rect 7119 8944 7131 8996
rect 7183 8944 7195 8996
rect 7247 8944 7259 8996
rect 7311 8944 7323 8996
rect 7375 8944 7387 8996
rect 7439 8944 7451 8996
rect 7503 8944 7509 8996
rect 7058 8928 7509 8944
rect 7058 8876 7067 8928
rect 7119 8876 7131 8928
rect 7183 8876 7195 8928
rect 7247 8876 7259 8928
rect 7311 8876 7323 8928
rect 7375 8876 7387 8928
rect 7439 8876 7451 8928
rect 7503 8876 7509 8928
tri 7011 8273 7058 8320 se
rect 7058 8273 7509 8876
rect 5418 7253 5682 7302
tri 5682 7253 5731 7302 sw
tri 6328 7253 6377 7302 se
rect 6377 7253 6610 7302
tri 6734 7996 7011 8273 se
rect 7011 7996 7509 8273
rect 6734 7295 7509 7996
tri 6734 7293 6736 7295 ne
rect 6736 7293 7507 7295
tri 7507 7293 7509 7295 nw
tri 6736 7253 6776 7293 ne
rect 6776 7253 7467 7293
tri 7467 7253 7507 7293 nw
tri 7559 7253 7599 7293 se
rect 7599 7253 7791 10512
rect 8181 7618 8363 10512
rect 8419 7760 9126 10512
tri 8419 7674 8505 7760 ne
rect 8505 7674 9126 7760
tri 8363 7618 8419 7674 sw
tri 8505 7618 8561 7674 ne
rect 8561 7618 9126 7674
rect 8181 7527 8419 7618
tri 8181 7499 8209 7527 ne
rect 5418 7246 5731 7253
tri 5731 7246 5738 7253 sw
tri 6321 7246 6328 7253 se
rect 6328 7246 6610 7253
tri 6610 7246 6617 7253 sw
tri 6776 7246 6783 7253 ne
rect 6783 7246 7460 7253
tri 7460 7246 7467 7253 nw
tri 7552 7246 7559 7253 se
rect 7559 7246 7791 7253
rect 5418 7194 5738 7246
tri 5738 7194 5790 7246 sw
tri 6269 7194 6321 7246 se
rect 6321 7194 6617 7246
tri 6617 7194 6669 7246 sw
tri 6783 7235 6794 7246 ne
rect 6794 7235 7449 7246
tri 7449 7235 7460 7246 nw
tri 7541 7235 7552 7246 se
rect 7552 7235 7791 7246
rect 8209 7476 8419 7527
tri 8419 7476 8561 7618 sw
tri 8561 7476 8703 7618 ne
rect 8703 7476 9126 7618
rect 8209 7444 8561 7476
tri 8561 7444 8593 7476 sw
tri 8703 7444 8735 7476 ne
rect 8735 7444 9126 7476
rect 8209 7302 8593 7444
tri 8593 7302 8735 7444 sw
tri 8735 7302 8877 7444 ne
rect 8877 7302 9126 7444
rect 8209 7253 8735 7302
tri 8735 7253 8784 7302 sw
rect 8209 7246 8784 7253
tri 8784 7246 8791 7253 sw
tri 6794 7194 6835 7235 ne
rect 6835 7203 7417 7235
tri 7417 7203 7449 7235 nw
tri 7509 7203 7541 7235 se
rect 7541 7203 7791 7235
rect 6835 7194 7408 7203
tri 7408 7194 7417 7203 nw
tri 7500 7194 7509 7203 se
rect 7509 7194 7791 7203
tri 7791 7194 7832 7235 sw
rect 8209 7194 8791 7246
tri 8791 7194 8843 7246 sw
rect 5418 6956 5790 7194
tri 5790 6956 6028 7194 sw
tri 5397 5586 5418 5607 se
rect 5418 5586 6028 6956
tri 5345 5534 5397 5586 se
rect 5397 5534 6028 5586
tri 5316 5505 5345 5534 se
rect 5345 5505 6028 5534
tri 5256 5445 5316 5505 se
rect 5316 5445 6028 5505
tri 4877 5411 4911 5445 sw
tri 5222 5411 5256 5445 se
rect 5256 5411 6028 5445
rect 4825 5359 4831 5411
rect 4883 5359 4895 5411
rect 4947 5359 4953 5411
tri 5170 5359 5222 5411 se
rect 5222 5359 6028 5411
tri 5141 5330 5170 5359 se
rect 5170 5330 6028 5359
tri 5110 5299 5141 5330 se
rect 5141 5299 6028 5330
tri 5094 5283 5110 5299 se
rect 5110 5283 6028 5299
tri 5063 5252 5094 5283 se
rect 5094 5252 6028 5283
tri 5042 5231 5063 5252 se
rect 5063 5231 6028 5252
tri 5024 5213 5042 5231 se
rect 5042 5213 6028 5231
rect 5024 5124 6028 5213
rect 4418 5066 4637 5118
rect 4689 5066 4717 5118
rect 4418 5049 4717 5066
rect 4418 4997 4637 5049
rect 4689 4997 4717 5049
rect 4418 4980 4717 4997
rect 4418 4928 4637 4980
rect 4689 4928 4717 4980
rect 4418 4911 4717 4928
rect 4418 4859 4637 4911
rect 4689 4859 4717 4911
rect 4829 5066 4892 5124
rect 4829 5014 4840 5066
rect 4829 4964 4892 5014
rect 4829 4912 4840 4964
rect 4418 4842 4717 4859
rect 4418 4790 4637 4842
rect 4689 4790 4717 4842
rect 4418 4773 4717 4790
rect 4418 4721 4637 4773
rect 4689 4721 4717 4773
rect 4418 4586 4717 4721
rect 4418 4534 4565 4586
rect 4617 4534 4637 4586
rect 4689 4534 4717 4586
rect 4418 4408 4717 4534
rect 4418 4356 4637 4408
rect 4689 4356 4717 4408
rect 4418 4342 4717 4356
rect 4418 4290 4637 4342
rect 4689 4290 4717 4342
rect 4418 4275 4717 4290
rect 4418 4223 4637 4275
rect 4689 4223 4717 4275
rect 4418 4208 4717 4223
rect 4418 4156 4637 4208
rect 4689 4156 4717 4208
rect 4418 4030 4717 4156
rect 4418 3978 4637 4030
rect 4689 3978 4717 4030
rect 4418 3963 4717 3978
rect 4418 3937 4637 3963
tri 4418 3911 4444 3937 ne
rect 4444 3911 4637 3937
rect 4689 3911 4717 3963
tri 4444 3896 4459 3911 ne
rect 4459 3896 4717 3911
tri 4459 3857 4498 3896 ne
rect 4498 3844 4637 3896
rect 4689 3844 4717 3896
rect 4258 3654 4310 3697
rect 4258 3560 4310 3602
rect 4258 3279 4310 3508
rect 4258 3211 4310 3227
rect 4258 3143 4310 3159
rect 4258 3075 4310 3091
rect 4258 3008 4310 3023
rect 4098 2876 4150 2888
rect 4098 2818 4150 2824
rect 4258 2941 4310 2956
rect 4258 2874 4310 2889
rect 4258 2807 4310 2822
rect 4258 2740 4310 2755
rect 3750 2539 3884 2591
rect 3936 2539 3948 2591
rect 4000 2539 4012 2591
rect 4064 2539 4070 2591
rect 3750 2395 4070 2539
rect 3750 2343 3884 2395
rect 3936 2343 3948 2395
rect 4000 2343 4012 2395
rect 4064 2343 4070 2395
rect 3750 2191 4070 2343
rect 3750 2139 3884 2191
rect 3936 2139 3948 2191
rect 4000 2139 4012 2191
rect 4064 2139 4070 2191
rect 3750 1308 4070 2139
rect 3750 1256 3884 1308
rect 3936 1256 3948 1308
rect 4000 1256 4012 1308
rect 4064 1256 4070 1308
rect 3750 992 4070 1256
rect 3750 940 3884 992
rect 3936 940 3948 992
rect 4000 940 4012 992
rect 4064 940 4070 992
rect 3750 682 4070 940
rect 3750 630 3884 682
rect 3936 630 3948 682
rect 4000 630 4012 682
rect 4064 630 4070 682
tri 3656 448 3676 468 sw
rect 3750 454 4070 630
rect 4098 2674 4150 2680
rect 4098 2610 4150 2622
rect 4098 1966 4150 2558
rect 4258 2673 4310 2688
rect 4258 2606 4310 2621
rect 4258 2539 4310 2554
rect 4098 1902 4150 1914
rect 4098 842 4150 1850
rect 4178 2492 4230 2498
rect 4178 2428 4230 2440
rect 4178 1210 4230 2376
rect 4178 1146 4230 1158
rect 4178 1088 4230 1094
rect 4258 2472 4310 2487
rect 4258 2405 4310 2420
rect 4258 2338 4310 2353
rect 4258 2271 4310 2286
rect 4258 1990 4310 2219
rect 4258 1875 4310 1938
rect 4258 1370 4310 1823
rect 4418 3831 4470 3837
rect 4418 3767 4470 3779
rect 4418 3232 4470 3715
rect 4418 3168 4470 3180
rect 4418 2382 4470 3116
rect 4418 2318 4470 2330
rect 4418 1783 4470 2266
rect 4418 1719 4470 1731
rect 4418 1661 4470 1667
rect 4498 3829 4717 3844
rect 4498 3777 4637 3829
rect 4689 3777 4717 3829
rect 4498 3762 4717 3777
rect 4498 3710 4637 3762
rect 4689 3710 4717 3762
rect 4498 3695 4717 3710
rect 4498 3643 4637 3695
rect 4689 3643 4717 3695
rect 4498 3628 4717 3643
rect 4498 3576 4637 3628
rect 4689 3576 4717 3628
rect 4498 3560 4717 3576
rect 4498 3508 4637 3560
rect 4689 3508 4717 3560
rect 4498 3394 4717 3508
rect 4498 3342 4637 3394
rect 4689 3342 4717 3394
rect 4498 3318 4717 3342
rect 4498 3266 4637 3318
rect 4689 3266 4717 3318
rect 4498 3242 4717 3266
rect 4498 3190 4637 3242
rect 4689 3190 4717 3242
rect 4498 3076 4717 3190
rect 4498 3024 4637 3076
rect 4689 3024 4717 3076
rect 4498 3010 4717 3024
rect 4498 2958 4637 3010
rect 4689 2958 4717 3010
rect 4498 2943 4717 2958
rect 4498 2891 4637 2943
rect 4689 2891 4717 2943
rect 4498 2876 4717 2891
rect 4498 2824 4637 2876
rect 4689 2824 4717 2876
rect 4498 2809 4717 2824
rect 4498 2757 4637 2809
rect 4689 2757 4717 2809
rect 4498 2742 4717 2757
rect 4498 2690 4637 2742
rect 4689 2690 4717 2742
rect 4498 2675 4717 2690
rect 4498 2623 4637 2675
rect 4689 2623 4717 2675
rect 4498 2608 4717 2623
rect 4498 2556 4637 2608
rect 4689 2556 4717 2608
rect 4498 2541 4717 2556
rect 4498 2489 4637 2541
rect 4689 2489 4717 2541
rect 4498 2474 4717 2489
rect 4498 2422 4637 2474
rect 4689 2422 4717 2474
rect 4498 1687 4717 2422
tri 4492 1635 4498 1641 se
rect 4498 1635 4637 1687
rect 4689 1635 4717 1687
rect 4258 1262 4310 1318
tri 4150 842 4158 850 sw
rect 4098 836 4158 842
tri 4158 836 4164 842 sw
rect 4098 830 4164 836
rect 4098 778 4112 830
rect 4098 756 4164 778
rect 4098 704 4112 756
rect 4098 682 4164 704
rect 4098 630 4112 682
rect 4098 609 4164 630
rect 4098 557 4112 609
rect 4098 536 4164 557
rect 4098 484 4112 536
rect 4098 478 4164 484
rect 4258 698 4310 1210
rect 4258 624 4310 646
rect 4258 550 4310 572
rect 4258 477 4310 498
rect 3178 446 3676 448
tri 3676 446 3678 448 sw
rect 3178 425 3678 446
tri 3678 425 3699 446 sw
rect 3178 411 3699 425
tri 3699 411 3713 425 sw
rect 3178 409 3713 411
tri 3713 409 3715 411 sw
rect 3178 384 3715 409
tri 3715 384 3740 409 sw
tri 4233 384 4258 409 se
rect 4258 384 4310 425
rect 3178 332 4310 384
tri 4468 1611 4492 1635 se
rect 4492 1611 4717 1635
rect 4468 1609 4717 1611
rect 4468 1557 4637 1609
rect 4689 1557 4717 1609
rect 4468 1530 4717 1557
rect 4468 1478 4637 1530
rect 4689 1478 4717 1530
rect 4468 1451 4717 1478
rect 4468 1399 4637 1451
rect 4689 1399 4717 1451
rect 4468 1372 4717 1399
rect 4468 1320 4637 1372
rect 4689 1320 4717 1372
rect 4468 463 4717 1320
rect 4468 411 4637 463
rect 4689 411 4717 463
rect 4468 351 4717 411
rect 3178 326 3744 332
tri 3744 326 3750 332 nw
rect 3178 299 3717 326
tri 3717 299 3744 326 nw
rect 4468 299 4637 351
rect 4689 299 4717 351
rect 3178 -139 3716 299
tri 3716 298 3717 299 nw
rect 4468 293 4717 299
rect 4749 4864 4801 4870
rect 4749 4779 4801 4812
rect 4749 4693 4801 4727
rect 4749 3990 4801 4641
rect 4749 3924 4801 3938
rect 4749 3858 4801 3872
rect 4749 3791 4801 3806
rect 4749 1788 4801 3739
rect 4749 1723 4801 1736
rect 4749 1658 4801 1671
rect 4749 1592 4801 1606
rect 4749 1526 4801 1540
rect 4749 201 4801 1474
rect 4829 4777 4892 4912
rect 4829 4725 4840 4777
rect 4829 4708 4892 4725
rect 4829 4656 4840 4708
rect 4829 4639 4892 4656
rect 4829 4587 4840 4639
rect 4829 4570 4892 4587
rect 4829 4518 4840 4570
rect 4829 4501 4892 4518
rect 4829 4449 4840 4501
rect 4829 4432 4892 4449
rect 4829 4380 4840 4432
rect 4829 4362 4892 4380
rect 4829 4310 4840 4362
rect 4829 4292 4892 4310
rect 4829 4240 4840 4292
rect 4829 4222 4892 4240
rect 4829 4170 4840 4222
rect 4829 3339 4892 4170
rect 4829 3287 4840 3339
rect 4829 3274 4892 3287
rect 4829 3222 4840 3274
rect 4829 3209 4892 3222
rect 4829 3157 4840 3209
rect 4829 3144 4892 3157
rect 4829 3092 4840 3144
rect 4829 3079 4892 3092
rect 4829 3027 4840 3079
rect 4829 3014 4892 3027
rect 4829 2962 4840 3014
rect 4829 2949 4892 2962
rect 4829 2897 4840 2949
rect 4829 2884 4892 2897
rect 4829 2832 4840 2884
rect 4829 2818 4892 2832
rect 4829 2766 4840 2818
rect 4829 2752 4892 2766
rect 4829 2700 4840 2752
rect 4829 2686 4892 2700
rect 4829 2634 4840 2686
rect 4829 2620 4892 2634
rect 4829 2568 4840 2620
rect 4829 2554 4892 2568
rect 4829 2502 4840 2554
rect 4829 2488 4892 2502
rect 4829 2436 4840 2488
rect 4829 1536 4892 2436
rect 4829 1533 4889 1536
tri 4889 1533 4892 1536 nw
rect 5024 5072 5034 5124
rect 5086 5072 5100 5124
rect 5152 5072 5166 5124
rect 5218 5072 5232 5124
rect 5284 5072 5298 5124
rect 5350 5072 5364 5124
rect 5416 5072 5430 5124
rect 5482 5072 5496 5124
rect 5548 5072 5562 5124
rect 5614 5072 5628 5124
rect 5680 5072 5694 5124
rect 5746 5072 5760 5124
rect 5812 5072 5826 5124
rect 5878 5072 5892 5124
rect 5944 5072 5959 5124
rect 6011 5072 6028 5124
rect 5024 3747 6028 5072
rect 5024 3695 5163 3747
rect 5215 3695 5230 3747
rect 5282 3695 5297 3747
rect 5349 3695 5364 3747
rect 5416 3695 5431 3747
rect 5483 3695 5498 3747
rect 5550 3695 5565 3747
rect 5617 3695 5632 3747
rect 5684 3695 5699 3747
rect 5751 3695 5766 3747
rect 5818 3695 5834 3747
rect 5886 3695 5902 3747
rect 5954 3695 5970 3747
rect 6022 3695 6028 3747
rect 5024 3683 6028 3695
rect 5024 3631 5163 3683
rect 5215 3631 5230 3683
rect 5282 3631 5297 3683
rect 5349 3631 5364 3683
rect 5416 3631 5431 3683
rect 5483 3631 5498 3683
rect 5550 3631 5565 3683
rect 5617 3631 5632 3683
rect 5684 3631 5699 3683
rect 5751 3631 5766 3683
rect 5818 3631 5834 3683
rect 5886 3631 5902 3683
rect 5954 3631 5970 3683
rect 6022 3631 6028 3683
rect 5024 3350 6028 3631
rect 5024 3314 5452 3350
tri 5452 3314 5488 3350 nw
tri 5689 3314 5725 3350 ne
rect 5725 3314 6028 3350
rect 5024 3312 5450 3314
tri 5450 3312 5452 3314 nw
tri 5725 3312 5727 3314 ne
rect 5727 3312 6028 3314
rect 5024 3260 5398 3312
tri 5398 3260 5450 3312 nw
tri 5727 3260 5779 3312 ne
rect 5779 3260 6028 3312
rect 5024 3220 5358 3260
tri 5358 3220 5398 3260 nw
tri 5779 3220 5819 3260 ne
rect 5819 3220 6028 3260
rect 5024 3198 5336 3220
tri 5336 3198 5358 3220 nw
tri 5819 3208 5831 3220 ne
rect 5024 3189 5327 3198
tri 5327 3189 5336 3198 nw
rect 5024 3188 5326 3189
tri 5326 3188 5327 3189 nw
rect 5024 1615 5311 3188
tri 5311 3173 5326 3188 nw
rect 5377 3136 5383 3188
rect 5435 3136 5447 3188
rect 5499 3136 5505 3188
rect 5377 3108 5436 3136
tri 5436 3108 5464 3136 nw
rect 5377 3102 5430 3108
tri 5430 3102 5436 3108 nw
tri 5374 2743 5377 2746 se
rect 5377 2743 5429 3102
tri 5429 3101 5430 3102 nw
tri 5429 2743 5432 2746 sw
tri 5370 2739 5374 2743 se
rect 5374 2739 5432 2743
tri 5432 2739 5436 2743 sw
tri 5343 2712 5370 2739 se
rect 5370 2712 5436 2739
tri 5436 2712 5463 2739 sw
rect 5339 2660 5345 2712
rect 5397 2660 5409 2712
rect 5461 2660 5467 2712
tri 5347 2658 5349 2660 ne
rect 5349 2658 5457 2660
tri 5457 2658 5459 2660 nw
tri 5349 2632 5375 2658 ne
rect 5375 2632 5431 2658
tri 5431 2632 5457 2658 nw
tri 5375 2630 5377 2632 ne
rect 5024 1563 5043 1615
rect 5095 1563 5113 1615
rect 5165 1563 5183 1615
rect 5235 1563 5253 1615
rect 5305 1563 5311 1615
rect 5024 1551 5311 1563
rect 4829 411 4883 1533
tri 4883 1527 4889 1533 nw
rect 4881 359 4883 411
rect 4829 309 4883 359
rect 4881 257 4883 309
rect 4829 238 4883 257
rect 5024 1499 5043 1551
rect 5095 1499 5113 1551
rect 5165 1499 5183 1551
rect 5235 1499 5253 1551
rect 5305 1499 5311 1551
rect 5024 253 5311 1499
tri 4801 201 4803 203 sw
rect 5024 201 5034 253
rect 5086 201 5107 253
rect 5159 201 5180 253
rect 5232 201 5253 253
rect 5305 201 5311 253
rect 4749 169 4803 201
tri 4803 169 4835 201 sw
rect 4749 117 4755 169
rect 4807 117 4819 169
rect 4871 117 4877 169
rect 5377 117 5429 2632
tri 5429 2630 5431 2632 nw
rect 5831 1615 6028 3220
rect 5831 1563 5837 1615
rect 5889 1563 5903 1615
rect 5955 1563 5970 1615
rect 6022 1563 6028 1615
rect 5831 1551 6028 1563
rect 5831 1499 5837 1551
rect 5889 1499 5903 1551
rect 5955 1499 5970 1551
rect 6022 1499 6028 1551
rect 5831 253 6028 1499
rect 5831 201 5838 253
rect 5890 201 5902 253
rect 5954 201 5966 253
rect 6018 201 6028 253
tri 6136 7061 6269 7194 se
rect 6269 7141 6669 7194
tri 6669 7141 6722 7194 sw
tri 6835 7141 6888 7194 ne
rect 6888 7141 7355 7194
tri 7355 7141 7408 7194 nw
tri 7447 7141 7500 7194 se
rect 7500 7141 7832 7194
rect 6269 7061 6722 7141
rect 6136 6956 6722 7061
tri 6722 6956 6907 7141 sw
rect 6136 5486 6907 6956
tri 7387 7081 7447 7141 se
rect 7447 7081 7832 7141
rect 7387 6981 7832 7081
tri 7832 6981 8045 7194 sw
rect 6136 5414 6731 5486
tri 6731 5414 6803 5486 nw
rect 6136 5411 6728 5414
tri 6728 5411 6731 5414 nw
rect 6136 5124 6652 5411
tri 6652 5335 6728 5411 nw
rect 6774 5231 6780 5283
rect 6832 5231 6844 5283
rect 6896 5231 6902 5283
tri 6784 5203 6812 5231 ne
rect 6136 5072 6142 5124
rect 6194 5072 6206 5124
rect 6258 5072 6270 5124
rect 6322 5072 6334 5124
rect 6386 5072 6399 5124
rect 6451 5072 6464 5124
rect 6516 5072 6529 5124
rect 6581 5072 6594 5124
rect 6646 5072 6652 5124
rect 6136 4206 6652 5072
tri 6805 4394 6812 4401 se
rect 6812 4394 6864 5231
tri 6864 5203 6892 5231 nw
rect 6963 5124 7331 6918
rect 6963 5072 6969 5124
rect 7021 5072 7045 5124
rect 7097 5072 7121 5124
rect 7173 5072 7197 5124
rect 7249 5072 7273 5124
rect 7325 5072 7331 5124
tri 6864 4394 6871 4401 sw
tri 6799 4388 6805 4394 se
rect 6805 4388 6871 4394
tri 6871 4388 6877 4394 sw
tri 6784 4373 6799 4388 se
rect 6799 4373 6877 4388
tri 6877 4373 6892 4388 sw
rect 6774 4321 6780 4373
rect 6832 4321 6844 4373
rect 6896 4321 6902 4373
tri 6652 4206 6694 4248 sw
rect 6963 4212 7331 5072
rect 7387 5505 8045 6981
rect 8209 7001 8843 7194
tri 8843 7001 9036 7194 sw
rect 8209 5941 9036 7001
tri 9036 5941 9128 6033 sw
tri 8206 5530 8209 5533 se
rect 8209 5530 9128 5941
rect 9184 5601 9323 10512
rect 9497 7317 9566 10490
rect 9612 7555 10025 10512
tri 9612 7459 9708 7555 ne
rect 9708 7459 10025 7555
tri 9566 7317 9708 7459 sw
tri 9708 7317 9850 7459 ne
rect 9850 7317 10025 7459
rect 9497 7302 9708 7317
tri 9708 7302 9723 7317 sw
tri 9850 7302 9865 7317 ne
rect 9865 7302 10025 7317
rect 9497 7246 9723 7302
tri 9723 7246 9779 7302 sw
rect 9497 7194 9779 7246
tri 9779 7194 9831 7246 sw
rect 9497 7048 9831 7194
tri 9497 7001 9544 7048 ne
rect 9544 7001 9831 7048
tri 9831 7001 10024 7194 sw
tri 9541 5627 9544 5630 se
rect 9544 5627 10024 7001
tri 9323 5601 9349 5627 sw
tri 9515 5601 9541 5627 se
rect 9541 5601 10024 5627
rect 9184 5593 10024 5601
tri 9184 5586 9191 5593 ne
rect 9191 5586 10024 5593
tri 9191 5534 9243 5586 ne
rect 9243 5534 10024 5586
tri 9243 5533 9244 5534 ne
rect 9244 5533 10024 5534
tri 8045 5505 8070 5530 sw
rect 7387 5124 8070 5505
rect 7387 5072 7393 5124
rect 7445 5072 7461 5124
rect 7513 5072 7529 5124
rect 7581 5072 7598 5124
rect 7650 5072 7667 5124
rect 7719 5072 7736 5124
rect 7788 5072 7805 5124
rect 7857 5072 7874 5124
rect 7926 5072 7943 5124
rect 7995 5072 8012 5124
rect 8064 5072 8070 5124
rect 6136 4193 6694 4206
tri 6694 4193 6707 4206 sw
rect 6136 4141 6707 4193
tri 6707 4141 6759 4193 sw
rect 6136 4128 6759 4141
tri 6759 4128 6772 4141 sw
rect 6136 4099 6772 4128
tri 6772 4099 6801 4128 sw
rect 6136 3747 6907 4099
rect 6136 3631 6142 3747
rect 6706 3695 6719 3747
rect 6771 3695 6784 3747
rect 6836 3695 6849 3747
rect 6901 3695 6907 3747
rect 6706 3683 6907 3695
rect 6706 3631 6719 3683
rect 6771 3631 6784 3683
rect 6836 3631 6849 3683
rect 6901 3631 6907 3683
rect 6136 3624 6900 3631
tri 6900 3624 6907 3631 nw
rect 7387 3752 8070 5072
rect 7387 3700 7393 3752
rect 7445 3700 7461 3752
rect 7513 3700 7529 3752
rect 7581 3700 7598 3752
rect 7650 3700 7667 3752
rect 7719 3700 7736 3752
rect 7788 3700 7805 3752
rect 7857 3700 7874 3752
rect 7926 3700 7943 3752
rect 7995 3700 8012 3752
rect 8064 3700 8070 3752
rect 7387 3688 8070 3700
rect 7387 3636 7393 3688
rect 7445 3636 7461 3688
rect 7513 3636 7529 3688
rect 7581 3636 7598 3688
rect 7650 3636 7667 3688
rect 7719 3636 7736 3688
rect 7788 3636 7805 3688
rect 7857 3636 7874 3688
rect 7926 3636 7943 3688
rect 7995 3636 8012 3688
rect 8064 3636 8070 3688
rect 6136 3612 6888 3624
tri 6888 3612 6900 3624 nw
rect 6136 3560 6836 3612
tri 6836 3560 6888 3612 nw
rect 6136 3554 6830 3560
tri 6830 3554 6836 3560 nw
rect 6136 3548 6824 3554
tri 6824 3548 6830 3554 nw
rect 6136 3496 6772 3548
tri 6772 3496 6824 3548 nw
rect 6905 3496 6911 3548
rect 6963 3496 6975 3548
rect 7027 3496 7209 3548
rect 7261 3496 7273 3548
rect 7325 3496 7331 3548
rect 6136 3491 6767 3496
tri 6767 3491 6772 3496 nw
rect 6136 3484 6760 3491
tri 6760 3484 6767 3491 nw
rect 6136 3466 6742 3484
tri 6742 3466 6760 3484 nw
rect 6136 3447 6723 3466
tri 6723 3447 6742 3466 nw
rect 6136 3407 6683 3447
tri 6683 3407 6723 3447 nw
rect 6136 3356 6632 3407
tri 6632 3356 6683 3407 nw
rect 6136 3314 6590 3356
tri 6590 3314 6632 3356 nw
rect 7387 3314 8070 3636
rect 6136 3312 6588 3314
tri 6588 3312 6590 3314 nw
rect 6136 3260 6164 3312
rect 6216 3260 6241 3312
rect 6293 3260 6318 3312
rect 6370 3260 6395 3312
rect 6447 3260 6471 3312
rect 6523 3262 6538 3312
tri 6538 3262 6588 3312 nw
rect 7387 3262 7400 3314
rect 7452 3262 7467 3314
rect 7519 3262 7534 3314
rect 7586 3262 7601 3314
rect 7653 3262 7668 3314
rect 7720 3262 7735 3314
rect 7787 3262 7802 3314
rect 7854 3262 7869 3314
rect 7921 3262 7936 3314
rect 7988 3262 8002 3314
rect 8054 3262 8070 3314
rect 6523 3260 6536 3262
tri 6536 3260 6538 3262 nw
rect 6136 3220 6496 3260
tri 6496 3220 6536 3260 nw
rect 7387 3225 8070 3262
tri 7387 3220 7392 3225 ne
rect 7392 3220 8070 3225
rect 6136 1992 6479 3220
tri 6479 3203 6496 3220 nw
tri 7392 3203 7409 3220 ne
rect 7409 3203 8070 3220
tri 7409 3198 7414 3203 ne
rect 7414 3198 8070 3203
tri 7414 3189 7423 3198 ne
rect 7423 3189 8070 3198
tri 7423 3137 7475 3189 ne
rect 7475 3137 8070 3189
tri 7475 3113 7499 3137 ne
rect 7040 3102 7092 3108
rect 7040 3038 7092 3050
rect 7126 3019 7132 3071
rect 7184 3019 7196 3071
rect 7248 3019 7254 3071
tri 7146 3011 7154 3019 ne
rect 7154 3011 7254 3019
tri 7154 2999 7166 3011 ne
rect 7166 2999 7254 3011
rect 7040 2980 7092 2986
tri 7018 2807 7040 2829 se
rect 7040 2807 7085 2980
tri 7085 2973 7092 2980 nw
tri 7166 2973 7192 2999 ne
rect 7192 2973 7254 2999
tri 7192 2956 7209 2973 ne
tri 7199 2807 7209 2817 se
rect 7209 2807 7254 2973
tri 7006 2795 7018 2807 se
rect 7018 2795 7085 2807
rect 6957 2743 6963 2795
rect 7015 2743 7027 2795
rect 7079 2743 7085 2795
tri 7183 2791 7199 2807 se
rect 7199 2791 7254 2807
tri 7006 2739 7010 2743 ne
rect 7010 2739 7085 2743
rect 7126 2739 7132 2791
rect 7184 2739 7196 2791
rect 7248 2739 7254 2791
tri 7010 2710 7039 2739 ne
rect 7039 2710 7085 2739
tri 7165 2710 7194 2739 ne
rect 7194 2710 7254 2739
tri 7039 2709 7040 2710 ne
rect 6632 2535 6638 2587
rect 6690 2535 6702 2587
rect 6754 2586 6760 2587
rect 6754 2535 6760 2540
tri 6637 2510 6662 2535 ne
rect 6662 2510 6722 2535
tri 6722 2510 6747 2535 nw
rect 7040 2510 7085 2710
tri 7194 2697 7207 2710 ne
tri 7085 2510 7110 2535 sw
tri 6662 2506 6666 2510 ne
tri 6652 2138 6666 2152 se
rect 6666 2138 6718 2510
tri 6718 2506 6722 2510 nw
rect 7040 2458 7046 2510
rect 7098 2458 7110 2510
rect 7162 2458 7168 2510
tri 7187 2435 7207 2455 se
rect 7207 2435 7254 2710
tri 7182 2430 7187 2435 se
rect 7187 2430 7254 2435
rect 7126 2378 7132 2430
rect 7184 2378 7196 2430
rect 7248 2378 7254 2430
tri 6718 2138 6732 2152 sw
tri 6640 2126 6652 2138 se
rect 6652 2126 6732 2138
tri 6732 2126 6744 2138 sw
tri 6632 2118 6640 2126 se
rect 6640 2118 6744 2126
tri 6744 2118 6752 2126 sw
rect 6628 2066 6634 2118
rect 6686 2066 6698 2118
rect 6750 2066 6756 2118
tri 6632 2062 6636 2066 ne
rect 6636 2062 6748 2066
tri 6748 2062 6752 2066 nw
tri 6636 2032 6666 2062 ne
rect 6136 1940 6164 1992
rect 6216 1940 6243 1992
rect 6295 1940 6322 1992
rect 6374 1940 6401 1992
rect 6453 1940 6479 1992
rect 6136 1615 6479 1940
rect 6136 1563 6142 1615
rect 6194 1563 6211 1615
rect 6263 1563 6281 1615
rect 6333 1563 6351 1615
rect 6403 1563 6421 1615
rect 6473 1563 6479 1615
rect 6136 1551 6479 1563
rect 6136 1499 6142 1551
rect 6194 1499 6211 1551
rect 6263 1499 6281 1551
rect 6333 1499 6351 1551
rect 6403 1499 6421 1551
rect 6473 1499 6479 1551
rect 6666 1526 6718 2062
tri 6718 2032 6748 2062 nw
rect 6892 1700 6898 1752
rect 6950 1700 6962 1752
rect 7014 1700 7271 1752
rect 7323 1700 7335 1752
rect 7387 1700 7393 1752
rect 7499 1578 8070 3137
tri 6718 1526 6728 1536 sw
rect 7499 1526 7505 1578
rect 7557 1526 7578 1578
rect 7630 1526 7651 1578
rect 7703 1526 7724 1578
rect 7776 1526 7796 1578
rect 7848 1526 7868 1578
rect 7920 1526 7940 1578
rect 7992 1526 8012 1578
rect 8064 1526 8070 1578
rect 6666 1525 6728 1526
tri 6728 1525 6729 1526 sw
rect 6666 1523 6729 1525
tri 6729 1523 6731 1525 sw
rect 6666 1514 6731 1523
tri 6731 1514 6740 1523 sw
tri 6666 1509 6671 1514 ne
rect 6671 1509 6740 1514
tri 6740 1509 6745 1514 sw
rect 6136 253 6479 1499
tri 6671 1457 6723 1509 ne
rect 6723 1457 6745 1509
tri 6745 1457 6797 1509 sw
tri 6723 1443 6737 1457 ne
rect 6737 1443 6797 1457
tri 6797 1443 6811 1457 sw
tri 6737 1440 6740 1443 ne
rect 6740 1440 6811 1443
tri 6811 1440 6814 1443 sw
tri 6740 1417 6763 1440 ne
rect 6763 1417 6814 1440
tri 6814 1417 6837 1440 sw
tri 6763 1366 6814 1417 ne
rect 6814 1366 6837 1417
tri 6837 1366 6888 1417 sw
tri 6814 1365 6815 1366 ne
rect 6815 1365 6888 1366
tri 6888 1365 6889 1366 sw
tri 6815 1353 6827 1365 ne
rect 6827 1353 6889 1365
tri 6889 1353 6901 1365 sw
tri 6827 1301 6879 1353 ne
rect 6879 1301 6901 1353
tri 6901 1301 6953 1353 sw
tri 6879 1292 6888 1301 ne
rect 6888 1292 6953 1301
tri 6953 1292 6962 1301 sw
tri 6888 1259 6921 1292 ne
rect 6921 1259 6962 1292
tri 6962 1259 6995 1292 sw
tri 6921 1244 6936 1259 ne
rect 6936 1244 6995 1259
tri 6995 1244 7010 1259 sw
tri 6936 1218 6962 1244 ne
rect 6962 1218 7010 1244
tri 7010 1218 7036 1244 sw
tri 6962 1192 6988 1218 ne
rect 6988 1192 7036 1218
tri 7036 1192 7062 1218 sw
tri 6988 1189 6991 1192 ne
rect 6991 1189 7062 1192
tri 7062 1189 7065 1192 sw
tri 6991 1177 7003 1189 ne
rect 7003 1177 7065 1189
tri 7065 1177 7077 1189 sw
tri 7003 1144 7036 1177 ne
rect 7036 1144 7077 1177
tri 7077 1144 7110 1177 sw
tri 7036 1125 7055 1144 ne
rect 7055 1125 7110 1144
tri 7110 1125 7129 1144 sw
tri 7055 1119 7061 1125 ne
rect 7061 1119 7129 1125
tri 7129 1119 7135 1125 sw
tri 7061 1110 7070 1119 ne
rect 7070 1110 7135 1119
tri 7135 1110 7144 1119 sw
tri 7070 1070 7110 1110 ne
rect 7110 1070 7144 1110
tri 7144 1070 7184 1110 sw
tri 7110 1058 7122 1070 ne
rect 7122 1058 7184 1070
tri 7184 1058 7196 1070 sw
tri 7122 1049 7131 1058 ne
rect 7131 1049 7196 1058
tri 7196 1049 7205 1058 sw
tri 7131 1045 7135 1049 ne
rect 7135 1045 7205 1049
tri 7205 1045 7209 1049 sw
tri 7135 1043 7137 1045 ne
rect 7137 1043 7209 1045
tri 7209 1043 7211 1045 sw
tri 7137 1019 7161 1043 ne
rect 7161 1022 7211 1043
tri 7211 1022 7232 1043 sw
rect 7161 1019 7232 1022
rect 6836 967 6842 1019
rect 6894 967 6906 1019
rect 6958 967 6964 1019
tri 7161 996 7184 1019 ne
rect 7184 996 7232 1019
tri 7232 996 7258 1022 sw
tri 7184 991 7189 996 ne
rect 7189 991 7258 996
tri 7258 991 7263 996 sw
tri 7189 979 7201 991 ne
rect 7201 979 7263 991
tri 7263 979 7275 991 sw
tri 7201 976 7204 979 ne
rect 7204 976 7275 979
tri 7275 976 7278 979 sw
tri 7204 967 7213 976 ne
rect 7213 970 7278 976
tri 7278 970 7284 976 sw
rect 7213 967 7284 970
tri 6836 929 6874 967 ne
rect 6136 201 6142 253
rect 6194 201 6211 253
rect 6263 201 6281 253
rect 6333 201 6351 253
rect 6403 201 6421 253
rect 6473 201 6479 253
tri 5429 117 5434 122 sw
rect 4749 85 4803 117
tri 4803 85 4835 117 nw
rect 5377 85 5434 117
tri 5434 85 5466 117 sw
tri 4724 -83 4749 -58 se
rect 4749 -83 4801 85
tri 4801 83 4803 85 nw
rect 5377 33 5383 85
rect 5435 33 5447 85
rect 5499 33 5505 85
tri 6839 -51 6874 -16 se
rect 6874 -41 6926 967
tri 6926 929 6964 967 nw
tri 7213 948 7232 967 ne
rect 7232 33 7284 967
rect 7499 253 8070 1526
rect 7499 201 7505 253
rect 7557 201 7577 253
rect 7629 201 7649 253
rect 7701 201 7721 253
rect 7773 201 7793 253
rect 7845 201 7866 253
rect 7918 201 7939 253
rect 7991 201 8012 253
rect 8064 201 8070 253
tri 8181 5505 8206 5530 se
rect 8206 5505 9128 5530
tri 9244 5515 9262 5533 ne
rect 9262 5515 10024 5533
tri 9128 5505 9138 5515 sw
tri 9262 5505 9272 5515 ne
rect 9272 5505 10024 5515
rect 8181 5124 9138 5505
tri 9272 5486 9291 5505 ne
rect 9291 5486 10024 5505
tri 9291 5414 9363 5486 ne
rect 9363 5414 10024 5486
tri 9363 5411 9366 5414 ne
rect 9366 5411 10024 5414
tri 9410 5377 9444 5411 ne
rect 8181 5072 8187 5124
rect 8239 5072 8255 5124
rect 8307 5072 8323 5124
rect 8375 5072 8391 5124
rect 8443 5072 8459 5124
rect 8511 5072 8528 5124
rect 8580 5072 8597 5124
rect 8649 5072 8666 5124
rect 8718 5072 8735 5124
rect 8787 5072 8804 5124
rect 8856 5072 8873 5124
rect 8925 5072 8942 5124
rect 8994 5072 9011 5124
rect 9063 5072 9080 5124
rect 9132 5072 9138 5124
rect 8181 3752 9138 5072
rect 8181 3700 8187 3752
rect 8239 3700 8255 3752
rect 8307 3700 8323 3752
rect 8375 3700 8391 3752
rect 8443 3700 8459 3752
rect 8511 3700 8528 3752
rect 8580 3700 8597 3752
rect 8649 3700 8666 3752
rect 8718 3700 8735 3752
rect 8787 3700 8804 3752
rect 8856 3700 8873 3752
rect 8925 3700 8942 3752
rect 8994 3700 9011 3752
rect 9063 3700 9080 3752
rect 9132 3700 9138 3752
rect 8181 3688 9138 3700
rect 8181 3636 8187 3688
rect 8239 3636 8255 3688
rect 8307 3636 8323 3688
rect 8375 3636 8391 3688
rect 8443 3636 8459 3688
rect 8511 3636 8528 3688
rect 8580 3636 8597 3688
rect 8649 3636 8666 3688
rect 8718 3636 8735 3688
rect 8787 3636 8804 3688
rect 8856 3636 8873 3688
rect 8925 3636 8942 3688
rect 8994 3636 9011 3688
rect 9063 3636 9080 3688
rect 9132 3636 9138 3688
rect 8181 3346 9138 3636
rect 8181 3304 8548 3346
tri 8548 3304 8590 3346 nw
tri 8802 3304 8844 3346 ne
rect 8844 3304 9138 3346
rect 8181 3277 8521 3304
tri 8521 3277 8548 3304 nw
tri 8844 3277 8871 3304 ne
rect 8871 3277 9138 3304
rect 8181 3272 8516 3277
tri 8516 3272 8521 3277 nw
tri 8871 3272 8876 3277 ne
rect 8876 3272 9138 3277
rect 8181 3220 8464 3272
tri 8464 3220 8516 3272 nw
tri 8876 3220 8928 3272 ne
rect 8928 3220 9138 3272
rect 8181 1578 8448 3220
tri 8448 3204 8464 3220 nw
tri 8928 3204 8944 3220 ne
rect 8944 3204 9138 3220
tri 8944 3201 8947 3204 ne
rect 8632 3137 8638 3189
rect 8690 3137 8702 3189
rect 8754 3137 8760 3189
tri 8636 3103 8670 3137 ne
tri 8638 2710 8670 2742 se
rect 8670 2710 8722 3137
tri 8722 3103 8756 3137 nw
rect 8777 2900 8783 2952
rect 8835 2900 8847 2952
rect 8899 2900 8905 2952
tri 8782 2865 8817 2900 ne
tri 8722 2710 8754 2742 sw
rect 8632 2658 8638 2710
rect 8690 2658 8702 2710
rect 8754 2658 8760 2710
tri 8636 2632 8662 2658 ne
rect 8662 2632 8730 2658
tri 8730 2632 8756 2658 nw
tri 8662 2624 8670 2632 ne
rect 8181 1526 8187 1578
rect 8239 1526 8289 1578
rect 8341 1526 8390 1578
rect 8442 1526 8448 1578
rect 8181 253 8448 1526
rect 8181 201 8187 253
rect 8239 201 8254 253
rect 8306 201 8322 253
rect 8374 201 8390 253
rect 8442 201 8448 253
rect 8554 1417 8606 1423
rect 8554 1353 8606 1365
tri 8552 201 8554 203 se
rect 8554 201 8606 1301
tri 8520 169 8552 201 se
rect 8552 169 8606 201
rect 8478 117 8484 169
rect 8536 117 8548 169
rect 8600 117 8606 169
rect 8670 201 8722 2632
tri 8722 2624 8730 2632 nw
rect 8817 203 8869 2900
tri 8869 2865 8904 2900 nw
tri 8940 1992 8947 1999 se
rect 8947 1992 9138 3204
rect 8940 1940 8946 1992
rect 8998 1940 9013 1992
rect 9065 1940 9080 1992
rect 9132 1940 9138 1992
tri 8940 1934 8946 1940 ne
rect 8946 1934 9138 1940
tri 8946 1933 8947 1934 ne
rect 8947 1577 9138 1934
rect 8947 1525 8953 1577
rect 9005 1525 9080 1577
rect 9132 1525 9138 1577
rect 8947 1513 9138 1525
rect 9444 5126 10024 5411
rect 9444 5103 9554 5126
rect 9444 5051 9459 5103
rect 9511 5074 9554 5103
rect 9606 5074 9622 5126
rect 9674 5074 9690 5126
rect 9742 5074 9759 5126
rect 9811 5074 9828 5126
rect 9880 5074 9897 5126
rect 9949 5074 9966 5126
rect 10018 5074 10024 5126
rect 9511 5051 10024 5074
rect 9444 5038 10024 5051
rect 9444 4986 9459 5038
rect 9511 4986 10024 5038
rect 9444 4973 10024 4986
rect 9444 4921 9459 4973
rect 9511 4921 10024 4973
rect 9444 4908 10024 4921
rect 9444 4856 9459 4908
rect 9511 4859 10024 4908
rect 9511 4856 9662 4859
rect 9444 4850 9662 4856
tri 9662 4850 9671 4859 nw
rect 9444 4843 9634 4850
rect 9444 4791 9459 4843
rect 9511 4822 9634 4843
tri 9634 4822 9662 4850 nw
rect 9511 4816 9628 4822
tri 9628 4816 9634 4822 nw
rect 9732 4816 9784 4822
rect 9511 4791 9592 4816
rect 9444 4778 9592 4791
tri 9592 4780 9628 4816 nw
rect 9444 4726 9459 4778
rect 9511 4726 9592 4778
rect 9444 4713 9592 4726
rect 9444 4661 9459 4713
rect 9511 4661 9592 4713
rect 9444 4648 9592 4661
rect 9444 4596 9459 4648
rect 9511 4596 9592 4648
rect 9732 4752 9784 4764
rect 9732 4698 9784 4700
tri 9784 4698 9795 4709 sw
tri 10052 4698 10063 4709 se
rect 10063 4698 10115 11142
tri 10324 11087 10379 11142 ne
tri 10379 11087 10453 11161 sw
tri 10379 11065 10401 11087 ne
rect 10143 4966 10195 11055
tri 10350 9559 10401 9610 se
rect 10401 9559 10453 11087
rect 10325 9507 10331 9559
rect 10383 9507 10395 9559
rect 10447 9507 10453 9559
tri 10350 9456 10401 9507 ne
rect 10143 4902 10195 4914
rect 10143 4844 10195 4850
rect 10267 5299 10319 5305
rect 10267 5235 10319 5247
rect 9732 4694 9795 4698
tri 9795 4694 9799 4698 sw
tri 10048 4694 10052 4698 se
rect 10052 4694 10115 4698
rect 9732 4675 9799 4694
tri 9799 4675 9818 4694 sw
tri 10029 4675 10048 4694 se
rect 10048 4675 10115 4694
rect 9732 4623 10115 4675
tri 10261 4631 10267 4637 se
rect 10267 4631 10319 5183
rect 10401 4799 10453 9507
rect 10483 7001 10932 10512
tri 11260 10443 11297 10480 se
rect 11297 10443 11356 11273
tri 11356 11241 11388 11273 nw
tri 11356 10443 11388 10475 sw
rect 11260 10391 11266 10443
rect 11318 10391 11330 10443
rect 11382 10391 11388 10443
tri 11260 10354 11297 10391 ne
tri 11292 9591 11297 9596 se
rect 11297 9591 11356 10391
tri 11356 10359 11388 10391 nw
tri 11260 9559 11292 9591 se
rect 11292 9559 11356 9591
tri 11356 9559 11388 9591 sw
rect 11260 9507 11266 9559
rect 11318 9507 11330 9559
rect 11382 9507 11388 9559
tri 10932 7001 11012 7081 sw
rect 10483 6070 11012 7001
tri 11422 6791 11436 6805 se
rect 11436 6791 11488 10753
rect 14045 10446 14365 10494
rect 13691 8273 13697 8325
rect 13749 8273 13761 8325
rect 13813 8273 13819 8325
tri 13724 8230 13767 8273 ne
rect 10483 5991 10933 6070
tri 10933 5991 11012 6070 nw
tri 11390 6759 11422 6791 se
rect 11422 6783 11488 6791
rect 11422 6759 11464 6783
tri 11464 6759 11488 6783 nw
rect 11390 6747 11452 6759
tri 11452 6747 11464 6759 nw
rect 10483 5394 10879 5991
tri 10879 5937 10933 5991 nw
tri 10879 5394 10899 5414 sw
rect 10483 5330 10899 5394
tri 10899 5330 10963 5394 sw
rect 10483 5324 10963 5330
tri 10963 5324 10969 5330 sw
rect 10483 5278 10969 5324
tri 10969 5278 11015 5324 sw
rect 11120 5278 11318 5505
rect 11390 5317 11442 6747
tri 11442 6737 11452 6747 nw
tri 11477 5759 11516 5798 se
rect 11516 5759 11825 6923
rect 12056 6204 12530 7917
tri 12056 6159 12101 6204 ne
rect 12101 6159 12530 6204
tri 12101 6145 12115 6159 ne
rect 12115 6145 12530 6159
tri 12115 6048 12212 6145 ne
rect 12212 6048 12530 6145
rect 12643 7246 12963 7917
rect 12991 7437 13344 7917
rect 12643 7194 12649 7246
rect 12701 7194 12733 7246
rect 12785 7194 12818 7246
rect 12870 7194 12903 7246
rect 12955 7194 12963 7246
rect 12643 6145 12963 7194
rect 12991 7194 12997 7246
rect 13049 7194 13069 7246
rect 13121 7194 13141 7246
rect 13193 7194 13213 7246
rect 13265 7194 13286 7246
rect 13338 7194 13344 7246
rect 12991 6266 13344 7194
rect 13767 6747 13819 8273
rect 16182 7126 16474 7936
tri 15264 6946 15298 6980 sw
rect 13767 6683 13819 6695
rect 13767 6625 13819 6631
rect 13873 6791 13879 6907
rect 13995 6791 14001 6907
tri 16029 6860 16063 6894 ne
tri 13129 6232 13163 6266 ne
rect 13163 6193 13344 6266
tri 13163 6159 13197 6193 ne
rect 13197 6159 13344 6193
tri 12963 6145 12977 6159 sw
tri 13197 6145 13211 6159 ne
rect 13211 6145 13344 6159
tri 13344 6145 13469 6270 sw
rect 12643 6113 12977 6145
tri 12977 6113 13009 6145 sw
tri 13211 6113 13243 6145 ne
rect 13243 6113 13469 6145
tri 12643 6048 12708 6113 ne
rect 12708 6048 13009 6113
tri 13009 6048 13074 6113 sw
tri 13243 6048 13308 6113 ne
rect 13308 6048 13469 6113
tri 13469 6048 13566 6145 sw
tri 12212 5991 12269 6048 ne
rect 12269 5991 12530 6048
tri 12530 5991 12587 6048 sw
tri 12708 6028 12728 6048 ne
rect 12728 6044 13074 6048
tri 13074 6044 13078 6048 sw
tri 13308 6044 13312 6048 ne
rect 13312 6044 13566 6048
rect 12728 6028 13078 6044
tri 13078 6028 13094 6044 sw
tri 13312 6028 13328 6044 ne
rect 13328 6028 13566 6044
tri 13566 6028 13586 6048 sw
tri 12728 6012 12744 6028 ne
rect 12744 6012 13094 6028
tri 13094 6012 13110 6028 sw
tri 13328 6012 13344 6028 ne
rect 13344 6012 13586 6028
tri 12744 5991 12765 6012 ne
rect 12765 5991 13110 6012
tri 13110 5991 13131 6012 sw
tri 13344 5991 13365 6012 ne
rect 13365 5991 13586 6012
tri 13586 5991 13623 6028 sw
tri 12269 5957 12303 5991 ne
rect 12303 5957 12587 5991
tri 12587 5957 12621 5991 sw
tri 12765 5957 12799 5991 ne
rect 12799 5957 13131 5991
tri 13131 5957 13165 5991 sw
tri 13365 5957 13399 5991 ne
rect 13399 5957 13623 5991
tri 13623 5957 13657 5991 sw
tri 12303 5937 12323 5957 ne
rect 12323 5937 12621 5957
tri 12621 5937 12641 5957 sw
tri 12799 5937 12819 5957 ne
rect 12819 5937 13165 5957
tri 13165 5937 13185 5957 sw
tri 13399 5937 13419 5957 ne
rect 13419 5937 13657 5957
tri 13657 5937 13677 5957 sw
rect 11477 5654 11825 5759
tri 12323 5730 12530 5937 ne
rect 12530 5935 12641 5937
tri 12641 5935 12643 5937 sw
tri 12819 5935 12821 5937 ne
rect 12821 5935 13185 5937
rect 12530 5925 12643 5935
tri 12643 5925 12653 5935 sw
tri 12821 5925 12831 5935 ne
rect 12831 5925 13185 5935
rect 12530 5747 12653 5925
tri 12653 5747 12831 5925 sw
tri 12831 5770 12986 5925 ne
rect 12986 5810 13185 5925
tri 13185 5810 13312 5937 sw
tri 13419 5810 13546 5937 ne
rect 13546 5810 13677 5937
rect 12986 5770 13312 5810
tri 13312 5770 13352 5810 sw
tri 13546 5770 13586 5810 ne
rect 13586 5770 13677 5810
tri 13677 5770 13844 5937 sw
tri 12986 5747 13009 5770 ne
rect 13009 5747 13352 5770
tri 13352 5747 13375 5770 sw
tri 13586 5747 13609 5770 ne
rect 13609 5747 13844 5770
rect 12530 5730 12831 5747
rect 11477 5639 11810 5654
tri 11810 5639 11825 5654 nw
tri 12530 5639 12621 5730 ne
rect 12621 5639 12831 5730
tri 12831 5639 12939 5747 sw
tri 13009 5695 13061 5747 ne
rect 13061 5724 13375 5747
tri 13375 5724 13398 5747 sw
tri 13609 5724 13632 5747 ne
rect 13632 5724 13844 5747
rect 13061 5695 13398 5724
tri 13398 5695 13427 5724 sw
tri 13632 5695 13661 5724 ne
tri 13061 5639 13117 5695 ne
rect 13117 5639 13427 5695
rect 11477 5367 11797 5639
tri 11797 5626 11810 5639 nw
tri 12621 5626 12634 5639 ne
rect 12634 5626 12939 5639
tri 12634 5620 12640 5626 ne
rect 12640 5620 12939 5626
tri 11905 5586 11939 5620 sw
tri 12640 5586 12674 5620 ne
rect 12674 5586 12939 5620
tri 11477 5343 11501 5367 ne
rect 11501 5343 11797 5367
tri 11501 5330 11514 5343 ne
rect 11514 5330 11797 5343
tri 11442 5317 11455 5330 sw
tri 11514 5317 11527 5330 ne
rect 11527 5317 11797 5330
rect 11390 5308 11455 5317
tri 11455 5308 11464 5317 sw
tri 11527 5308 11536 5317 ne
rect 11536 5308 11797 5317
tri 11390 5289 11409 5308 ne
rect 11409 5295 11464 5308
tri 11464 5295 11477 5308 sw
tri 11536 5295 11549 5308 ne
rect 11549 5295 11797 5308
rect 11409 5289 11477 5295
tri 11318 5278 11329 5289 sw
tri 11409 5278 11420 5289 ne
rect 11420 5278 11477 5289
tri 11477 5278 11494 5295 sw
tri 11549 5278 11566 5295 ne
rect 11566 5278 11797 5295
rect 11853 5534 11859 5586
rect 11911 5534 11923 5586
rect 11975 5534 11981 5586
tri 12674 5534 12726 5586 ne
rect 12726 5569 12939 5586
tri 12939 5569 13009 5639 sw
tri 13117 5569 13187 5639 ne
rect 13187 5569 13427 5639
rect 12726 5534 13009 5569
rect 11853 5505 11910 5534
tri 11910 5505 11939 5534 nw
tri 12726 5505 12755 5534 ne
rect 12755 5505 13009 5534
tri 13009 5505 13073 5569 sw
tri 13187 5505 13251 5569 ne
rect 13251 5505 13427 5569
tri 13427 5505 13617 5695 sw
rect 13661 5505 13844 5724
rect 11853 5330 11905 5505
tri 11905 5500 11910 5505 nw
tri 12755 5500 12760 5505 ne
rect 12760 5500 13073 5505
tri 12760 5343 12917 5500 ne
rect 12917 5444 13073 5500
tri 13073 5444 13134 5505 sw
tri 13251 5444 13312 5505 ne
rect 13312 5490 13617 5505
tri 13617 5490 13632 5505 sw
rect 12917 5389 13134 5444
tri 13134 5389 13189 5444 sw
rect 12917 5343 13189 5389
tri 13189 5343 13235 5389 sw
rect 13312 5371 13632 5490
tri 12917 5330 12930 5343 ne
rect 12930 5330 13235 5343
tri 13235 5330 13248 5343 sw
rect 11853 5278 11859 5330
rect 11911 5278 11926 5330
rect 11978 5278 11984 5330
rect 12401 5278 12407 5330
rect 12459 5278 12474 5330
rect 12526 5321 12738 5330
tri 12738 5321 12747 5330 sw
tri 12930 5321 12939 5330 ne
rect 12939 5321 13248 5330
tri 13248 5321 13257 5330 sw
rect 12526 5320 12747 5321
tri 12747 5320 12748 5321 sw
tri 12939 5320 12940 5321 ne
rect 12940 5320 13257 5321
rect 12526 5317 12748 5320
tri 12748 5317 12751 5320 sw
tri 12940 5317 12943 5320 ne
rect 12943 5317 13257 5320
rect 12526 5308 12751 5317
tri 12751 5308 12760 5317 sw
tri 12943 5308 12952 5317 ne
rect 12952 5308 13257 5317
rect 12526 5278 12760 5308
rect 10483 5252 11015 5278
tri 11015 5252 11041 5278 sw
rect 11120 5265 11329 5278
tri 11329 5265 11342 5278 sw
tri 11420 5265 11433 5278 ne
rect 11433 5265 11494 5278
tri 11494 5265 11507 5278 sw
rect 11120 5252 11342 5265
tri 11342 5252 11355 5265 sw
tri 11433 5252 11446 5265 ne
rect 11446 5252 11507 5265
rect 10483 5245 11041 5252
tri 11041 5245 11048 5252 sw
rect 11120 5245 11355 5252
tri 11355 5245 11362 5252 sw
tri 11446 5245 11453 5252 ne
rect 11453 5245 11507 5252
tri 11566 5247 11597 5278 ne
rect 10483 5228 11048 5245
tri 11048 5228 11065 5245 sw
rect 10483 5126 11065 5228
rect 11120 5243 11362 5245
tri 11362 5243 11364 5245 sw
tri 11453 5243 11455 5245 ne
rect 11120 5208 11364 5243
tri 11364 5208 11399 5243 sw
rect 11120 5207 11399 5208
tri 11120 5193 11134 5207 ne
rect 11134 5193 11399 5207
tri 11134 5178 11149 5193 ne
rect 11149 5178 11399 5193
tri 11149 5162 11165 5178 ne
rect 11165 5162 11399 5178
tri 11165 5126 11201 5162 ne
rect 11201 5126 11399 5162
rect 10483 5074 10490 5126
rect 10542 5074 10554 5126
rect 10606 5074 10618 5126
rect 10670 5074 10682 5126
rect 10734 5074 10747 5126
rect 10799 5074 10812 5126
rect 10864 5074 10877 5126
rect 10929 5074 10942 5126
rect 10994 5074 11007 5126
rect 11059 5074 11065 5126
rect 10483 4911 11065 5074
rect 10483 4859 10489 4911
rect 10541 4859 10553 4911
rect 10605 4859 10617 4911
rect 10669 4859 10682 4911
rect 10734 4859 10747 4911
rect 10799 4859 10812 4911
rect 10864 4859 10877 4911
rect 10929 4859 10942 4911
rect 10994 4859 11007 4911
rect 11059 4859 11065 4911
tri 10483 4851 10491 4859 ne
rect 10491 4851 11065 4859
tri 10491 4813 10529 4851 ne
rect 10529 4813 11065 4851
tri 10453 4799 10467 4813 sw
tri 10529 4799 10543 4813 ne
rect 10543 4799 11065 4813
rect 11201 5074 11207 5126
rect 11259 5074 11274 5126
rect 11326 5074 11341 5126
rect 11393 5074 11399 5126
rect 11455 5178 11507 5193
rect 11455 5120 11507 5126
rect 11597 5126 11797 5278
tri 12716 5246 12748 5278 ne
rect 12748 5265 12760 5278
tri 12760 5265 12803 5308 sw
tri 12952 5296 12964 5308 ne
rect 12748 5246 12803 5265
tri 12803 5246 12822 5265 sw
tri 12748 5227 12767 5246 ne
rect 12767 5227 12822 5246
rect 12228 5175 12234 5227
rect 12286 5175 12301 5227
rect 12353 5175 12359 5227
tri 12767 5224 12770 5227 ne
rect 10401 4797 10467 4799
tri 10467 4797 10469 4799 sw
tri 10543 4797 10545 4799 ne
rect 10545 4797 11065 4799
rect 10401 4791 10469 4797
tri 10401 4775 10417 4791 ne
tri 10253 4623 10261 4631 se
rect 10261 4623 10319 4631
rect 9444 4583 9592 4596
tri 9974 4589 10008 4623 ne
rect 9444 4531 9459 4583
rect 9511 4531 9592 4583
rect 9444 4518 9592 4531
rect 9444 4466 9459 4518
rect 9511 4466 9592 4518
rect 9444 4453 9592 4466
rect 9444 4401 9459 4453
rect 9511 4401 9592 4453
rect 9444 4388 9592 4401
rect 9444 4336 9459 4388
rect 9511 4336 9592 4388
rect 9444 4323 9592 4336
rect 9444 4271 9459 4323
rect 9511 4271 9592 4323
rect 9444 4258 9592 4271
rect 9444 4206 9459 4258
rect 9511 4206 9592 4258
rect 9928 4510 9980 4516
rect 9928 4446 9980 4458
rect 9444 4193 9592 4206
rect 9444 4141 9459 4193
rect 9511 4141 9592 4193
tri 9876 4183 9928 4235 se
rect 9928 4213 9980 4394
rect 9928 4183 9950 4213
tri 9950 4183 9980 4213 nw
tri 9862 4169 9876 4183 se
rect 9876 4169 9936 4183
tri 9936 4169 9950 4183 nw
tri 9854 4161 9862 4169 se
rect 9862 4161 9928 4169
tri 9928 4161 9936 4169 nw
rect 9444 4128 9592 4141
rect 9444 4076 9459 4128
rect 9511 4076 9592 4128
tri 9810 4117 9854 4161 se
rect 9854 4117 9884 4161
tri 9884 4117 9928 4161 nw
tri 9780 4087 9810 4117 se
rect 9810 4087 9854 4117
tri 9854 4087 9884 4117 nw
rect 9444 4063 9592 4076
tri 9766 4073 9780 4087 se
rect 9780 4073 9840 4087
tri 9840 4073 9854 4087 nw
rect 9444 4011 9459 4063
rect 9511 4011 9592 4063
tri 9752 4059 9766 4073 se
rect 9766 4059 9826 4073
tri 9826 4059 9840 4073 nw
tri 9748 4055 9752 4059 se
rect 9752 4055 9822 4059
tri 9822 4055 9826 4059 nw
rect 9444 3998 9592 4011
rect 9444 3946 9459 3998
rect 9511 3946 9592 3998
rect 9444 3933 9592 3946
rect 9444 3881 9459 3933
rect 9511 3881 9592 3933
rect 9444 3868 9592 3881
rect 9444 3816 9459 3868
rect 9511 3816 9592 3868
rect 9444 3804 9592 3816
rect 9444 3752 9459 3804
rect 9511 3752 9592 3804
rect 9444 3740 9592 3752
rect 9444 3688 9459 3740
rect 9511 3688 9592 3740
rect 9444 3676 9592 3688
rect 9444 3624 9459 3676
rect 9511 3624 9592 3676
rect 9444 3612 9592 3624
rect 9444 3560 9459 3612
rect 9511 3560 9592 3612
rect 9444 3548 9592 3560
rect 9444 3496 9459 3548
rect 9511 3496 9592 3548
rect 9444 3356 9592 3496
rect 9444 3304 9459 3356
rect 9511 3304 9592 3356
rect 9444 3272 9592 3304
rect 9444 3220 9459 3272
rect 9511 3220 9592 3272
rect 9444 1641 9592 3220
tri 9732 4039 9748 4055 se
rect 9748 4039 9806 4055
tri 9806 4039 9822 4055 nw
rect 9620 3148 9672 3154
rect 9620 3084 9672 3096
rect 9620 2397 9672 3032
rect 9620 2333 9672 2345
rect 9620 2275 9672 2281
rect 9444 1589 9459 1641
rect 9511 1589 9592 1641
rect 9444 1575 9592 1589
rect 9444 1523 9459 1575
rect 9511 1523 9592 1575
rect 8947 1509 9091 1513
tri 9091 1509 9095 1513 nw
rect 9444 1509 9592 1523
rect 8947 1457 9039 1509
tri 9039 1457 9091 1509 nw
rect 9444 1457 9459 1509
rect 9511 1457 9592 1509
rect 8947 1058 9026 1457
tri 9026 1444 9039 1457 nw
rect 9444 1443 9592 1457
rect 9444 1391 9459 1443
rect 9511 1391 9592 1443
rect 9444 1377 9592 1391
rect 9444 1325 9459 1377
rect 9511 1325 9592 1377
rect 9444 1311 9592 1325
rect 9444 1259 9459 1311
rect 9511 1259 9592 1311
rect 9444 1244 9592 1259
rect 9444 1192 9459 1244
rect 9511 1192 9592 1244
rect 9444 1177 9592 1192
rect 9444 1125 9459 1177
rect 9511 1125 9592 1177
rect 9444 1110 9592 1125
tri 9026 1058 9064 1096 sw
rect 9444 1058 9459 1110
rect 9511 1058 9592 1110
rect 8947 1049 9064 1058
tri 9064 1049 9073 1058 sw
rect 8947 1045 9073 1049
tri 9073 1045 9077 1049 sw
rect 8947 1043 9077 1045
tri 9077 1043 9079 1045 sw
rect 9444 1043 9592 1058
rect 8947 1027 9079 1043
tri 9079 1027 9095 1043 sw
rect 8947 253 9138 1027
rect 9444 991 9459 1043
rect 9511 991 9592 1043
rect 9444 976 9592 991
rect 9444 924 9459 976
rect 9511 924 9592 976
rect 9444 909 9592 924
rect 9444 857 9459 909
rect 9511 857 9592 909
rect 9444 842 9592 857
rect 9444 790 9459 842
rect 9511 790 9592 842
rect 9444 775 9592 790
rect 9444 723 9459 775
rect 9511 723 9592 775
rect 9444 708 9592 723
rect 9732 834 9784 4039
tri 9784 4017 9806 4039 nw
rect 9845 3407 9901 3414
rect 9845 3355 9848 3407
rect 9900 3355 9901 3407
rect 9845 3329 9901 3355
rect 9845 3277 9848 3329
rect 9900 3277 9901 3329
rect 9845 3250 9901 3277
rect 9845 3198 9848 3250
rect 9900 3198 9901 3250
rect 9845 3171 9901 3198
rect 9845 3119 9848 3171
rect 9900 3119 9901 3171
rect 9845 3092 9901 3119
rect 9845 3040 9848 3092
rect 9900 3040 9901 3092
rect 9845 1259 9901 3040
rect 10008 1399 10060 4623
tri 10060 4589 10094 4623 nw
tri 10219 4589 10253 4623 se
rect 10253 4611 10319 4623
rect 10253 4589 10287 4611
tri 10209 4579 10219 4589 se
rect 10219 4579 10287 4589
tri 10287 4579 10319 4611 nw
rect 10417 4765 10469 4791
tri 10545 4760 10582 4797 ne
rect 10417 4698 10469 4713
rect 10417 4631 10469 4646
tri 10195 4565 10209 4579 se
rect 10209 4565 10273 4579
tri 10273 4565 10287 4579 nw
rect 10417 4565 10469 4579
tri 10189 4559 10195 4565 se
rect 10195 4559 10267 4565
tri 10267 4559 10273 4565 nw
tri 10172 4542 10189 4559 se
rect 10189 4542 10250 4559
tri 10250 4542 10267 4559 nw
rect 10172 2367 10228 4542
tri 10228 4520 10250 4542 nw
rect 10417 4499 10469 4513
rect 10417 4433 10469 4447
rect 10417 4367 10469 4381
rect 10417 4301 10469 4315
rect 10417 4235 10469 4249
rect 10417 4169 10469 4183
rect 10417 4111 10469 4117
rect 10582 4055 11065 4797
rect 10582 4003 10588 4055
rect 10640 4003 10657 4055
rect 10709 4003 10727 4055
rect 10779 4003 10797 4055
rect 10849 4003 10867 4055
rect 10919 4003 10937 4055
rect 10989 4003 11007 4055
rect 11059 4003 11065 4055
rect 10391 3959 10443 3965
rect 10391 3895 10443 3907
rect 10391 3837 10443 3843
rect 10474 3831 10526 3837
rect 10474 3767 10526 3779
rect 10391 3703 10443 3709
rect 10391 3639 10443 3651
rect 10391 3581 10443 3587
rect 10391 3447 10443 3453
rect 10391 3383 10443 3395
rect 10391 3325 10443 3331
rect 10474 3319 10526 3715
rect 10474 3255 10526 3267
rect 10391 3063 10443 3069
rect 10391 2999 10443 3011
rect 10391 2941 10443 2947
rect 10474 2807 10526 3203
rect 10474 2743 10526 2755
rect 10391 2551 10443 2557
rect 10391 2487 10443 2499
rect 10391 2429 10443 2435
rect 10224 2315 10228 2367
rect 10172 2303 10228 2315
rect 10224 2251 10228 2303
rect 10474 2295 10526 2691
rect 10172 2245 10228 2251
rect 10391 2283 10443 2289
rect 10391 2219 10443 2231
rect 10391 2161 10443 2167
rect 10474 2231 10526 2243
rect 10391 1911 10443 1917
rect 10391 1847 10443 1859
rect 10391 1789 10443 1795
rect 10474 1783 10526 2179
rect 10474 1719 10526 1731
rect 10474 1661 10526 1667
rect 10582 3543 11065 4003
rect 10582 3491 10588 3543
rect 10640 3491 10657 3543
rect 10709 3491 10727 3543
rect 10779 3491 10797 3543
rect 10849 3491 10867 3543
rect 10919 3491 10937 3543
rect 10989 3491 11007 3543
rect 11059 3491 11065 3543
rect 10582 3031 11065 3491
rect 10582 2979 10588 3031
rect 10640 2979 10657 3031
rect 10709 2979 10727 3031
rect 10779 2979 10797 3031
rect 10849 2979 10867 3031
rect 10919 2979 10937 3031
rect 10989 2979 11007 3031
rect 11059 2979 11065 3031
rect 10582 2519 11065 2979
rect 10582 2467 10588 2519
rect 10640 2467 10657 2519
rect 10709 2467 10727 2519
rect 10779 2467 10797 2519
rect 10849 2467 10867 2519
rect 10919 2467 10937 2519
rect 10989 2467 11007 2519
rect 11059 2467 11065 2519
rect 10582 2007 11065 2467
rect 10582 1955 10588 2007
rect 10640 1955 10657 2007
rect 10709 1955 10727 2007
rect 10779 1955 10797 2007
rect 10849 1955 10867 2007
rect 10919 1955 10937 2007
rect 10989 1955 11007 2007
rect 11059 1955 11065 2007
rect 10391 1655 10443 1661
rect 10391 1591 10443 1603
rect 10391 1533 10443 1539
rect 10582 1495 11065 1955
rect 10582 1443 10588 1495
rect 10640 1443 10657 1495
rect 10709 1443 10727 1495
rect 10779 1443 10797 1495
rect 10849 1443 10867 1495
rect 10919 1443 10937 1495
rect 10989 1443 11007 1495
rect 11059 1443 11065 1495
rect 10008 1335 10060 1347
rect 10008 1277 10060 1283
rect 10416 1381 10468 1387
rect 10416 1311 10468 1329
tri 9901 1259 9902 1260 sw
rect 9845 1241 9902 1259
tri 9902 1241 9920 1259 sw
rect 10416 1241 10468 1259
rect 9845 1238 9920 1241
tri 9845 1232 9851 1238 ne
rect 9851 1232 9920 1238
tri 9920 1232 9929 1241 sw
tri 9851 1189 9894 1232 ne
rect 9894 1189 9929 1232
tri 9929 1189 9972 1232 sw
tri 9894 1182 9901 1189 ne
rect 9901 1182 9972 1189
tri 9901 1175 9908 1182 ne
rect 9908 1175 9972 1182
tri 9972 1175 9986 1189 sw
tri 9908 1171 9912 1175 ne
rect 9912 1171 9986 1175
tri 9986 1171 9990 1175 sw
rect 10416 1171 10468 1189
tri 9912 1154 9929 1171 ne
rect 9929 1154 9990 1171
tri 9990 1154 10007 1171 sw
tri 9929 1119 9964 1154 ne
rect 9964 1119 10007 1154
tri 10007 1119 10042 1154 sw
tri 9964 1110 9973 1119 ne
rect 9973 1110 10042 1119
tri 10042 1110 10051 1119 sw
tri 9973 1101 9982 1110 ne
rect 9982 1101 10051 1110
tri 10051 1101 10060 1110 sw
rect 10416 1101 10468 1119
tri 9982 1076 10007 1101 ne
rect 10007 1076 10060 1101
tri 10060 1076 10085 1101 sw
tri 10007 1049 10034 1076 ne
rect 10034 1049 10085 1076
tri 10085 1049 10112 1076 sw
tri 10034 1045 10038 1049 ne
rect 10038 1045 10112 1049
tri 10112 1045 10116 1049 sw
tri 10038 1032 10051 1045 ne
rect 10051 1032 10116 1045
tri 10116 1032 10129 1045 sw
tri 10051 1031 10052 1032 ne
rect 10052 1031 10129 1032
tri 10129 1031 10130 1032 sw
rect 10416 1031 10468 1049
tri 10052 998 10085 1031 ne
rect 10085 998 10130 1031
tri 10130 998 10163 1031 sw
tri 10085 979 10104 998 ne
rect 10104 979 10163 998
tri 10163 979 10182 998 sw
tri 10104 967 10116 979 ne
rect 10116 967 10182 979
tri 10182 967 10194 979 sw
tri 10116 961 10122 967 ne
rect 10122 961 10194 967
tri 10194 961 10200 967 sw
rect 10416 961 10468 979
tri 10122 920 10163 961 ne
rect 10163 920 10200 961
tri 10200 920 10241 961 sw
tri 10163 909 10174 920 ne
rect 10174 909 10241 920
tri 10174 902 10181 909 ne
rect 10181 902 10241 909
tri 10181 898 10185 902 ne
rect 9732 770 9784 782
rect 9732 712 9784 718
rect 10089 796 10141 802
rect 10089 732 10141 744
rect 9444 656 9459 708
rect 9511 656 9592 708
rect 9444 641 9592 656
rect 9444 589 9459 641
rect 9511 589 9592 641
rect 9444 574 9592 589
tri 10040 587 10089 636 se
rect 10089 614 10141 680
rect 10089 587 10114 614
tri 10114 587 10141 614 nw
rect 9444 522 9459 574
rect 9511 522 9592 574
tri 10015 562 10040 587 se
rect 10040 566 10093 587
tri 10093 566 10114 587 nw
rect 10040 562 10089 566
tri 10089 562 10093 566 nw
tri 10181 562 10185 566 se
rect 10185 562 10241 902
rect 10416 891 10468 909
rect 10416 822 10468 839
rect 10416 753 10468 770
tri 10569 753 10582 766 se
rect 10582 753 11065 1443
tri 10517 701 10569 753 se
rect 10569 701 11065 753
rect 10416 695 10468 701
tri 10511 695 10517 701 se
rect 10517 695 11065 701
rect 11121 4797 11173 4803
rect 11121 4727 11173 4745
rect 11121 4657 11173 4675
rect 11121 4587 11173 4605
rect 11121 4517 11173 4535
rect 11121 4447 11173 4465
rect 11121 4377 11173 4395
rect 11121 4307 11173 4325
rect 11121 4238 11173 4255
rect 11121 4169 11173 4186
rect 11121 3959 11173 4117
rect 11121 3895 11173 3907
rect 11121 3703 11173 3843
rect 11121 3639 11173 3651
rect 11121 3447 11173 3587
rect 11121 3383 11173 3395
rect 11121 1911 11173 3331
rect 11121 1847 11173 1859
rect 11121 1655 11173 1795
rect 11121 1591 11173 1603
rect 11121 1381 11173 1539
rect 11121 1311 11173 1329
rect 11121 1241 11173 1259
rect 11121 1171 11173 1189
rect 11121 1101 11173 1119
rect 11121 1031 11173 1049
rect 11121 961 11173 979
rect 11121 891 11173 909
rect 11121 822 11173 839
rect 11121 753 11173 770
rect 11121 695 11173 701
rect 11201 3727 11399 5074
rect 11597 5074 11603 5126
rect 11655 5074 11670 5126
rect 11722 5074 11737 5126
rect 11789 5074 11797 5126
tri 11399 3727 11422 3750 sw
tri 11574 3727 11597 3750 se
rect 11597 3727 11797 5074
rect 11959 5074 11965 5126
rect 12017 5074 12029 5126
rect 12081 5074 12093 5126
rect 12145 5074 12157 5126
rect 12209 5074 12221 5126
rect 12273 5074 12279 5126
rect 11959 4911 12279 5074
rect 11959 4859 11965 4911
rect 12017 4859 12029 4911
rect 12081 4859 12093 4911
rect 12145 4859 12157 4911
rect 12209 4859 12221 4911
rect 12273 4859 12279 4911
rect 11201 3694 11422 3727
tri 11422 3694 11455 3727 sw
tri 11541 3694 11574 3727 se
rect 11574 3694 11797 3727
rect 11201 3543 11797 3694
rect 11201 3491 11207 3543
rect 11259 3491 11273 3543
rect 11325 3491 11339 3543
rect 11391 3491 11405 3543
rect 11457 3491 11471 3543
rect 11523 3491 11537 3543
rect 11589 3491 11603 3543
rect 11655 3491 11670 3543
rect 11722 3491 11737 3543
rect 11789 3491 11797 3543
rect 11201 3031 11797 3491
rect 11201 2979 11207 3031
rect 11259 2979 11273 3031
rect 11325 2979 11339 3031
rect 11391 2979 11405 3031
rect 11457 2979 11471 3031
rect 11523 2979 11537 3031
rect 11589 2979 11603 3031
rect 11655 2979 11670 3031
rect 11722 2979 11737 3031
rect 11789 2979 11797 3031
rect 11201 2519 11797 2979
rect 11201 2467 11207 2519
rect 11259 2467 11273 2519
rect 11325 2467 11339 2519
rect 11391 2467 11405 2519
rect 11457 2467 11471 2519
rect 11523 2467 11537 2519
rect 11589 2467 11603 2519
rect 11655 2467 11670 2519
rect 11722 2467 11737 2519
rect 11789 2467 11797 2519
rect 11201 2007 11797 2467
rect 11201 1955 11207 2007
rect 11259 1955 11274 2007
rect 11326 1955 11341 2007
rect 11393 1955 11600 2007
rect 11652 1955 11668 2007
rect 11720 1955 11737 2007
rect 11789 1955 11797 2007
rect 9444 507 9592 522
rect 9444 455 9459 507
rect 9511 455 9592 507
tri 9951 498 10015 562 se
rect 10015 498 10025 562
tri 10025 498 10089 562 nw
tri 10117 498 10181 562 se
rect 10181 544 10241 562
rect 10181 498 10195 544
tri 10195 498 10241 544 nw
tri 10495 679 10511 695 se
rect 10511 679 11065 695
rect 10495 639 11065 679
rect 10495 587 10505 639
rect 10557 587 10576 639
rect 10628 587 10647 639
rect 10699 587 10719 639
rect 10771 587 10791 639
rect 10843 587 10863 639
rect 10915 587 10935 639
rect 10987 587 11007 639
rect 11059 587 11065 639
rect 10495 498 11065 587
tri 9941 488 9951 498 se
rect 9951 488 10015 498
tri 10015 488 10025 498 nw
tri 10107 488 10117 498 se
rect 10117 488 10185 498
tri 10185 488 10195 498 nw
rect 9444 440 9592 455
tri 9901 448 9941 488 se
rect 9941 448 9975 488
tri 9975 448 10015 488 nw
tri 10067 448 10107 488 se
rect 10107 448 10145 488
tri 10145 448 10185 488 nw
tri 9899 446 9901 448 se
rect 9901 446 9973 448
tri 9973 446 9975 448 nw
tri 10065 446 10067 448 se
rect 10067 446 10143 448
tri 10143 446 10145 448 nw
rect 10495 446 10501 498
rect 10553 446 10573 498
rect 10625 446 10645 498
rect 10697 446 10717 498
rect 10769 446 10789 498
rect 10841 446 10861 498
rect 10913 446 10934 498
rect 10986 446 11007 498
rect 11059 446 11065 498
rect 11201 498 11797 1955
rect 11851 4797 11903 4803
rect 11851 4727 11903 4745
rect 11851 4657 11903 4675
rect 11851 4587 11903 4605
rect 11851 4517 11903 4535
rect 11851 4447 11903 4465
rect 11851 4377 11903 4395
rect 11851 4307 11903 4325
rect 11851 4238 11903 4255
rect 11851 4169 11903 4186
rect 11851 3447 11903 4117
rect 11851 3383 11903 3395
rect 11851 1381 11903 3331
rect 11851 1311 11903 1329
rect 11851 1241 11903 1259
rect 11851 1171 11903 1189
rect 11851 1101 11903 1119
rect 11851 1031 11903 1049
rect 11851 961 11903 979
rect 11851 891 11903 909
rect 11851 822 11903 839
rect 11851 753 11903 770
rect 11851 695 11903 701
rect 11959 3031 12279 4859
rect 11959 2979 11965 3031
rect 12017 2979 12029 3031
rect 12081 2979 12093 3031
rect 12145 2979 12157 3031
rect 12209 2979 12221 3031
rect 12273 2979 12279 3031
rect 11959 2519 12279 2979
rect 11959 2467 11965 2519
rect 12017 2467 12029 2519
rect 12081 2467 12093 2519
rect 12145 2467 12157 2519
rect 12209 2467 12221 2519
rect 12273 2467 12279 2519
rect 11201 446 11207 498
rect 11259 446 11273 498
rect 11325 446 11339 498
rect 11391 446 11405 498
rect 11457 446 11471 498
rect 11523 446 11537 498
rect 11589 446 11603 498
rect 11655 446 11670 498
rect 11722 446 11737 498
rect 11789 446 11797 498
rect 11959 639 12279 2467
rect 12307 3905 12359 5175
rect 12307 3816 12359 3853
rect 12307 3727 12359 3764
rect 12307 3638 12359 3675
rect 12307 1912 12359 3586
rect 12307 1833 12359 1860
rect 12307 1753 12359 1781
rect 12307 1673 12359 1701
rect 12307 1593 12359 1621
rect 12307 1535 12359 1541
rect 12393 5126 12721 5221
rect 12393 5074 12399 5126
rect 12451 5074 12495 5126
rect 12547 5112 12721 5126
rect 12547 5074 12669 5112
rect 12393 5060 12669 5074
rect 12393 5047 12721 5060
rect 12393 4995 12669 5047
rect 12393 4982 12721 4995
rect 12393 4930 12669 4982
rect 12393 4917 12721 4930
rect 12393 4911 12669 4917
rect 12393 4859 12399 4911
rect 12451 4859 12493 4911
rect 12545 4865 12669 4911
rect 12545 4859 12721 4865
rect 12393 4851 12721 4859
rect 12393 4847 12669 4851
rect 12393 4055 12525 4847
tri 12525 4815 12557 4847 nw
tri 12636 4822 12661 4847 ne
rect 12553 4797 12633 4803
rect 12605 4745 12633 4797
rect 12553 4727 12633 4745
rect 12605 4675 12633 4727
rect 12553 4657 12633 4675
rect 12605 4605 12633 4657
rect 12553 4587 12633 4605
rect 12605 4535 12633 4587
rect 12553 4517 12633 4535
rect 12605 4465 12633 4517
rect 12553 4447 12633 4465
rect 12605 4395 12633 4447
rect 12553 4377 12633 4395
rect 12605 4325 12633 4377
rect 12553 4307 12633 4325
rect 12605 4255 12633 4307
rect 12553 4238 12633 4255
rect 12605 4186 12633 4238
rect 12553 4169 12633 4186
rect 12605 4117 12633 4169
rect 12553 4111 12633 4117
tri 12556 4086 12581 4111 ne
rect 12393 4003 12399 4055
rect 12451 4003 12467 4055
rect 12519 4003 12525 4055
rect 12393 3543 12525 4003
rect 12393 3491 12399 3543
rect 12451 3491 12467 3543
rect 12519 3491 12525 3543
rect 12393 3417 12525 3491
rect 12393 3395 12503 3417
tri 12503 3395 12525 3417 nw
rect 12581 3447 12633 4111
rect 12393 3383 12491 3395
tri 12491 3383 12503 3395 nw
rect 12581 3383 12633 3395
rect 12393 2138 12445 3383
tri 12445 3337 12491 3383 nw
rect 12473 3278 12525 3284
rect 12473 3214 12525 3226
rect 12473 2807 12525 3162
rect 12473 2743 12525 2755
rect 12473 2336 12525 2691
rect 12473 2272 12525 2284
rect 12473 2214 12525 2220
rect 12581 3191 12633 3331
rect 12581 3127 12633 3139
rect 12581 2807 12633 3075
rect 12581 2743 12633 2755
tri 12445 2138 12469 2162 sw
rect 12393 2126 12469 2138
tri 12469 2126 12481 2138 sw
rect 12393 2082 12481 2126
tri 12481 2082 12525 2126 sw
rect 12393 2007 12525 2082
rect 12393 1955 12399 2007
rect 12451 1955 12467 2007
rect 12519 1955 12525 2007
rect 11959 587 11965 639
rect 12017 587 12029 639
rect 12081 587 12093 639
rect 12145 587 12157 639
rect 12209 587 12221 639
rect 12273 587 12279 639
rect 11959 498 12279 587
rect 11959 446 11965 498
rect 12017 446 12029 498
rect 12081 446 12093 498
rect 12145 446 12157 498
rect 12209 446 12221 498
rect 12273 446 12279 498
rect 12393 1495 12525 1955
rect 12393 1443 12399 1495
rect 12451 1443 12467 1495
rect 12519 1443 12525 1495
rect 12393 676 12525 1443
tri 12556 1387 12581 1412 se
rect 12581 1387 12633 2691
rect 12553 1381 12633 1387
rect 12605 1329 12633 1381
rect 12553 1311 12633 1329
rect 12605 1259 12633 1311
rect 12553 1241 12633 1259
rect 12605 1189 12633 1241
rect 12553 1171 12633 1189
rect 12605 1119 12633 1171
rect 12553 1101 12633 1119
rect 12605 1049 12633 1101
rect 12553 1031 12633 1049
rect 12605 979 12633 1031
rect 12553 961 12633 979
rect 12605 909 12633 961
rect 12553 891 12633 909
rect 12605 839 12633 891
rect 12553 822 12633 839
rect 12605 770 12633 822
rect 12553 753 12633 770
rect 12605 701 12633 753
rect 12553 695 12633 701
rect 12661 4799 12669 4847
rect 12661 4785 12721 4799
rect 12661 4733 12669 4785
rect 12661 4719 12721 4733
rect 12661 4667 12669 4719
rect 12661 4653 12721 4667
rect 12661 4601 12669 4653
rect 12661 4587 12721 4601
rect 12661 4535 12669 4587
rect 12661 4521 12721 4535
rect 12661 4469 12669 4521
rect 12661 4455 12721 4469
rect 12661 4403 12669 4455
rect 12661 4389 12721 4403
rect 12661 4337 12669 4389
rect 12661 4323 12721 4337
rect 12661 4271 12669 4323
rect 12661 4257 12721 4271
rect 12661 4205 12669 4257
rect 12661 4191 12721 4205
rect 12661 4139 12669 4191
rect 12661 4125 12721 4139
rect 12661 4073 12669 4125
rect 12661 4059 12721 4073
rect 12661 4007 12669 4059
rect 12661 3993 12721 4007
rect 12661 3941 12669 3993
rect 12661 3927 12721 3941
rect 12661 3875 12669 3927
rect 12661 3676 12721 3875
rect 12770 3835 12822 5227
rect 12964 5158 13257 5308
rect 13873 5162 14001 6791
tri 14365 5324 14430 5389 sw
rect 14365 5265 14430 5324
tri 14430 5265 14489 5324 sw
rect 13873 5046 13879 5162
rect 13995 5046 14001 5162
tri 15676 5162 15723 5209 sw
tri 15250 5075 15281 5106 ne
rect 15281 5075 15394 5106
rect 15676 5075 15723 5162
tri 15723 5075 15810 5162 sw
tri 15281 5046 15310 5075 ne
rect 15310 5046 15394 5075
tri 15647 5046 15676 5075 se
rect 15676 5046 15810 5075
tri 15310 5041 15315 5046 ne
rect 15315 5041 15394 5046
tri 15642 5041 15647 5046 se
rect 15647 5041 15810 5046
tri 15810 5041 15844 5075 sw
tri 15315 4962 15394 5041 ne
rect 15394 4945 15747 5041
tri 14813 4697 14890 4774 ne
rect 12770 3768 12822 3783
rect 12770 3710 12822 3716
rect 12713 3624 12721 3676
rect 12661 3606 12721 3624
rect 12713 3554 12721 3606
rect 12661 3536 12721 3554
rect 12713 3484 12721 3536
rect 12661 3466 12721 3484
rect 12713 3414 12721 3466
rect 12661 3395 12721 3414
rect 12713 3343 12721 3395
rect 12661 3324 12721 3343
rect 12713 3272 12721 3324
rect 12661 3253 12721 3272
rect 12713 3201 12721 3253
rect 12661 3182 12721 3201
rect 12713 3130 12721 3182
rect 12661 3111 12721 3130
rect 12713 3059 12721 3111
rect 12661 3040 12721 3059
rect 12713 2988 12721 3040
rect 12661 2796 12721 2988
rect 12713 2744 12721 2796
rect 12661 2714 12721 2744
rect 12713 2662 12721 2714
rect 12661 2632 12721 2662
rect 12713 2580 12721 2632
rect 12661 2549 12721 2580
rect 12713 2497 12721 2549
rect 12661 2254 12721 2497
rect 12713 2202 12721 2254
rect 12661 2190 12721 2202
rect 12713 2138 12721 2190
rect 12661 2126 12721 2138
rect 12713 2074 12721 2126
rect 12661 2062 12721 2074
rect 12713 2010 12721 2062
rect 12661 1998 12721 2010
rect 12713 1946 12721 1998
rect 12661 1934 12721 1946
rect 12713 1882 12721 1934
rect 12661 1870 12721 1882
rect 12713 1818 12721 1870
rect 12661 1806 12721 1818
rect 12713 1754 12721 1806
rect 12661 1742 12721 1754
rect 12713 1690 12721 1742
rect 12661 1678 12721 1690
rect 12713 1626 12721 1678
rect 12661 1614 12721 1626
rect 12713 1562 12721 1614
rect 12661 1550 12721 1562
rect 12713 1498 12721 1550
rect 12661 1486 12721 1498
rect 12713 1434 12721 1486
rect 12661 1422 12721 1434
rect 12713 1370 12721 1422
rect 12661 1357 12721 1370
rect 12713 1305 12721 1357
rect 12661 1292 12721 1305
rect 12713 1240 12721 1292
rect 12661 1227 12721 1240
rect 12713 1175 12721 1227
rect 12661 1162 12721 1175
rect 12713 1110 12721 1162
rect 12661 1097 12721 1110
rect 12713 1045 12721 1097
rect 12661 1032 12721 1045
rect 12713 980 12721 1032
rect 12661 967 12721 980
rect 12713 915 12721 967
rect 12661 902 12721 915
rect 12713 850 12721 902
rect 12661 837 12721 850
rect 12713 785 12721 837
rect 12661 772 12721 785
rect 12713 720 12721 772
rect 12661 707 12721 720
tri 12525 676 12532 683 sw
rect 12393 655 12532 676
tri 12532 655 12553 676 sw
tri 12640 655 12661 676 se
rect 12713 655 12721 707
rect 12393 651 12553 655
tri 12553 651 12557 655 sw
tri 12636 651 12640 655 se
rect 12640 651 12721 655
rect 12393 642 12721 651
rect 12393 639 12661 642
rect 12393 587 12399 639
rect 12451 587 12500 639
rect 12552 590 12661 639
rect 12713 590 12721 642
rect 12552 587 12721 590
rect 12393 498 12721 587
rect 12393 446 12399 498
rect 12451 446 12500 498
rect 12552 446 12721 498
rect 9444 388 9459 440
rect 9511 388 9592 440
tri 9867 414 9899 446 se
rect 9899 414 9941 446
tri 9941 414 9973 446 nw
tri 10033 414 10065 446 se
rect 10065 414 10107 446
rect 9444 373 9592 388
rect 9444 321 9459 373
rect 9511 321 9592 373
tri 9793 340 9867 414 se
tri 9867 340 9941 414 nw
tri 10029 410 10033 414 se
rect 10033 410 10107 414
tri 10107 410 10143 446 nw
tri 9959 340 10029 410 se
tri 9138 253 9172 287 sw
tri 8869 203 8883 217 sw
tri 8722 201 8724 203 sw
rect 8817 201 8883 203
tri 8883 201 8885 203 sw
rect 8947 201 8953 253
rect 9005 201 9033 253
rect 9085 201 9114 253
rect 9166 201 9172 253
rect 8670 169 8724 201
tri 8724 169 8756 201 sw
rect 8817 195 8885 201
tri 8817 169 8843 195 ne
rect 8843 194 8885 195
tri 8885 194 8892 201 sw
rect 9444 194 9592 321
tri 9740 287 9793 340 se
rect 9793 287 9814 340
tri 9814 287 9867 340 nw
tri 9951 332 9959 340 se
rect 9959 332 10029 340
tri 10029 332 10107 410 nw
tri 9906 287 9951 332 se
rect 9951 287 9984 332
tri 9984 287 10029 332 nw
tri 9719 266 9740 287 se
rect 9740 266 9793 287
tri 9793 266 9814 287 nw
tri 9885 266 9906 287 se
rect 9906 266 9951 287
tri 9688 235 9719 266 se
rect 9719 235 9762 266
tri 9762 235 9793 266 nw
tri 9873 254 9885 266 se
rect 9885 254 9951 266
tri 9951 254 9984 287 nw
tri 9854 235 9873 254 se
rect 9873 235 9932 254
tri 9932 235 9951 254 nw
rect 10080 235 10086 287
rect 10138 235 10150 287
rect 10202 235 10208 287
tri 9677 224 9688 235 se
rect 9688 224 9751 235
tri 9751 224 9762 235 nw
tri 9843 224 9854 235 se
rect 9854 224 9921 235
tri 9921 224 9932 235 nw
tri 10080 224 10091 235 ne
rect 10091 224 10197 235
tri 10197 224 10208 235 nw
rect 10455 235 10461 287
rect 10513 235 10525 287
rect 10577 235 10583 287
tri 11394 235 11435 276 se
rect 11435 235 11840 276
tri 10455 224 10466 235 ne
rect 10466 224 10572 235
tri 10572 224 10583 235 nw
tri 11383 224 11394 235 se
rect 11394 224 11840 235
rect 11892 224 11917 276
rect 11969 224 11994 276
rect 12046 224 12070 276
rect 12122 224 12128 276
tri 9650 197 9677 224 se
rect 9677 197 9724 224
tri 9724 197 9751 224 nw
tri 9816 197 9843 224 se
rect 9843 197 9894 224
tri 9894 197 9921 224 nw
tri 10091 197 10118 224 ne
tri 9647 194 9650 197 se
rect 9650 194 9719 197
rect 8843 192 8892 194
tri 8892 192 8894 194 sw
tri 9645 192 9647 194 se
rect 9647 192 9719 194
tri 9719 192 9724 197 nw
tri 9811 192 9816 197 se
rect 9816 192 9873 197
rect 8843 169 8894 192
tri 8894 169 8917 192 sw
tri 9622 169 9645 192 se
rect 9645 176 9703 192
tri 9703 176 9719 192 nw
tri 9795 176 9811 192 se
rect 9811 176 9873 192
tri 9873 176 9894 197 nw
rect 9645 169 9656 176
rect 8670 117 8676 169
rect 8728 117 8740 169
rect 8792 117 8798 169
tri 8843 129 8883 169 ne
rect 8883 129 8917 169
tri 8917 129 8957 169 sw
tri 9582 129 9622 169 se
rect 9622 129 9656 169
tri 9656 129 9703 176 nw
tri 9748 129 9795 176 se
tri 8883 117 8895 129 ne
rect 8895 117 9625 129
tri 8895 77 8935 117 ne
rect 8935 98 9625 117
tri 9625 98 9656 129 nw
tri 9717 98 9748 129 se
rect 9748 98 9795 129
tri 9795 98 9873 176 nw
rect 8935 77 9604 98
tri 9604 77 9625 98 nw
tri 9696 77 9717 98 se
rect 9717 77 9736 98
tri 9674 55 9696 77 se
rect 9696 55 9736 77
tri 7284 33 7306 55 sw
tri 9658 39 9674 55 se
rect 9674 39 9736 55
tri 9736 39 9795 98 nw
tri 9652 33 9658 39 se
rect 9658 33 9730 39
tri 9730 33 9736 39 nw
tri 10112 33 10118 39 se
rect 10118 33 10170 224
tri 10170 197 10197 224 nw
tri 10466 197 10493 224 ne
tri 7232 1 7264 33 ne
rect 7264 3 7306 33
tri 7306 3 7336 33 sw
tri 9639 20 9652 33 se
rect 9652 20 9717 33
tri 9717 20 9730 33 nw
tri 10099 20 10112 33 se
rect 10112 20 10170 33
tri 9622 3 9639 20 se
rect 9639 3 9700 20
tri 9700 3 9717 20 nw
tri 10082 3 10099 20 se
rect 10099 3 10170 20
rect 7264 1 7336 3
tri 7336 1 7338 3 sw
tri 9620 1 9622 3 se
rect 9622 1 9698 3
tri 9698 1 9700 3 nw
tri 10080 1 10082 3 se
rect 10082 1 10170 3
tri 10170 1 10208 39 sw
tri 7264 -16 7281 1 ne
rect 7281 -16 7338 1
tri 6926 -41 6951 -16 sw
tri 7281 -41 7306 -16 ne
rect 7306 -41 7338 -16
tri 7338 -41 7380 1 sw
tri 9578 -41 9620 1 se
rect 9620 -41 9646 1
rect 6874 -45 6951 -41
tri 6951 -45 6955 -41 sw
tri 7306 -45 7310 -41 ne
rect 7310 -45 7380 -41
tri 7380 -45 7384 -41 sw
tri 9574 -45 9578 -41 se
rect 9578 -45 9646 -41
rect 6874 -51 6955 -45
tri 6955 -51 6961 -45 sw
tri 7310 -51 7316 -45 ne
rect 7316 -51 7384 -45
tri 7384 -51 7390 -45 sw
tri 9568 -51 9574 -45 se
rect 9574 -51 9646 -45
tri 9646 -51 9698 1 nw
rect 10080 -51 10086 1
rect 10138 -51 10150 1
rect 10202 -51 10208 1
tri 10487 -51 10493 -45 se
rect 10493 -51 10545 224
tri 10545 197 10572 224 nw
tri 11356 197 11383 224 se
rect 11383 197 11427 224
tri 11353 194 11356 197 se
rect 11356 194 11427 197
tri 11427 194 11457 224 nw
tri 11328 169 11353 194 se
rect 11353 169 11402 194
tri 11402 169 11427 194 nw
tri 11310 151 11328 169 se
rect 11328 151 11384 169
tri 11384 151 11402 169 nw
tri 11276 117 11310 151 se
rect 11310 117 11350 151
tri 11350 117 11384 151 nw
tri 11244 85 11276 117 se
rect 11276 85 11318 117
tri 11318 85 11350 117 nw
tri 11236 77 11244 85 se
rect 11244 77 11310 85
tri 11310 77 11318 85 nw
tri 11192 33 11236 77 se
rect 11236 33 11266 77
tri 11266 33 11310 77 nw
tri 11162 3 11192 33 se
rect 11192 3 11236 33
tri 11236 3 11266 33 nw
tri 11118 -41 11162 3 se
rect 11162 -41 11192 3
tri 11192 -41 11236 3 nw
tri 11114 -45 11118 -41 se
rect 11118 -45 11188 -41
tri 11188 -45 11192 -41 nw
rect 4661 -135 4667 -83
rect 4719 -135 4743 -83
rect 4795 -135 4801 -83
tri 6836 -54 6839 -51 se
rect 6839 -54 6961 -51
tri 6961 -54 6964 -51 sw
tri 7316 -54 7319 -51 ne
rect 7319 -54 7390 -51
tri 7390 -54 7393 -51 sw
tri 9565 -54 9568 -51 se
rect 9568 -54 9643 -51
tri 9643 -54 9646 -51 nw
tri 10484 -54 10487 -51 se
rect 10487 -54 10545 -51
tri 10545 -54 10554 -45 sw
tri 11105 -54 11114 -45 se
rect 11114 -54 11179 -45
tri 11179 -54 11188 -45 nw
rect 6836 -106 6842 -54
rect 6894 -106 6906 -54
rect 6958 -106 6964 -54
tri 7319 -106 7371 -54 ne
rect 7371 -106 7393 -54
tri 7393 -106 7445 -54 sw
rect 7968 -106 7974 -54
rect 8026 -106 8038 -54
rect 8090 -83 9614 -54
tri 9614 -83 9643 -54 nw
tri 10455 -83 10484 -54 se
rect 10484 -83 10554 -54
tri 10554 -83 10583 -54 sw
tri 11088 -71 11105 -54 se
rect 11105 -71 11162 -54
tri 11162 -71 11179 -54 nw
tri 11076 -83 11088 -71 se
rect 11088 -83 11150 -71
tri 11150 -83 11162 -71 nw
rect 8090 -106 9591 -83
tri 9591 -106 9614 -83 nw
tri 7371 -115 7380 -106 ne
rect 7380 -115 7445 -106
tri 7445 -115 7454 -106 sw
tri 7380 -135 7400 -115 ne
rect 7400 -135 7454 -115
tri 7454 -135 7474 -115 sw
rect 10455 -135 10461 -83
rect 10513 -135 10525 -83
rect 10577 -135 10583 -83
tri 11053 -106 11076 -83 se
rect 11076 -106 11127 -83
tri 11127 -106 11150 -83 nw
tri 11044 -115 11053 -106 se
rect 11053 -115 11118 -106
tri 11118 -115 11127 -106 nw
tri 11024 -135 11044 -115 se
rect 11044 -135 11088 -115
tri 7400 -139 7404 -135 ne
rect 7404 -139 7474 -135
tri 7404 -189 7454 -139 ne
rect 7454 -145 7474 -139
tri 7474 -145 7484 -135 sw
tri 11014 -145 11024 -135 se
rect 11024 -145 11088 -135
tri 11088 -145 11118 -115 nw
rect 7454 -167 7484 -145
tri 7484 -167 7506 -145 sw
tri 10992 -167 11014 -145 se
rect 11014 -167 11044 -145
rect 7454 -189 11044 -167
tri 11044 -189 11088 -145 nw
tri 7454 -219 7484 -189 ne
rect 7484 -219 11014 -189
tri 11014 -219 11044 -189 nw
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_0
timestamp 1701704242
transform 1 0 10836 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_1
timestamp 1701704242
transform 1 0 9649 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_2
timestamp 1701704242
transform 1 0 12566 0 1 -142
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_3
timestamp 1701704242
transform 1 0 11187 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_4
timestamp 1701704242
transform 1 0 6516 0 1 -142
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_5
timestamp 1701704242
transform 1 0 8299 0 1 -142
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_6
timestamp 1701704242
transform 1 0 10428 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_7
timestamp 1701704242
transform 1 0 10783 0 1 -142
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_8
timestamp 1701704242
transform 1 0 10057 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_9
timestamp 1701704242
transform 1 0 12562 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_10
timestamp 1701704242
transform 1 0 12154 0 1 196
box 0 0 1 1
use DFL1_CDNS_524688791851239  DFL1_CDNS_524688791851239_11
timestamp 1701704242
transform 1 0 11595 0 1 196
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform 0 -1 1420 -1 0 2461
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform 0 -1 727 -1 0 2797
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform 0 -1 1086 -1 0 2797
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform 0 -1 283 -1 0 2973
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform 0 -1 1012 -1 0 3314
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 0 -1 1086 -1 0 2564
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 0 -1 369 -1 0 4756
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1701704242
transform 0 -1 1086 -1 0 5151
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1701704242
transform 0 -1 1160 -1 0 5290
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1701704242
transform 0 -1 1086 -1 0 4793
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1701704242
transform 0 -1 1086 -1 0 1373
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1701704242
transform 0 -1 383 -1 0 1804
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1701704242
transform 0 -1 383 -1 0 1133
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1701704242
transform 0 -1 48 -1 0 3728
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1701704242
transform 0 1 693 -1 0 4887
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1701704242
transform -1 0 3028 0 1 2511
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1701704242
transform -1 0 619 0 1 2731
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1701704242
transform -1 0 619 0 1 2529
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1701704242
transform -1 0 547 0 1 2823
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1701704242
transform -1 0 895 0 1 842
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1701704242
transform -1 0 1326 0 1 5427
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1701704242
transform -1 0 5173 0 1 2173
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1701704242
transform -1 0 5064 0 1 2411
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1701704242
transform -1 0 10048 0 -1 4921
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1701704242
transform -1 0 9812 0 -1 4921
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1701704242
transform -1 0 5064 0 -1 3058
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1701704242
transform -1 0 9314 0 -1 2460
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1701704242
transform -1 0 7324 0 -1 2498
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1701704242
transform -1 0 5064 0 -1 2783
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1701704242
transform -1 0 9314 0 -1 3065
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1701704242
transform -1 0 7324 0 -1 2182
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1701704242
transform -1 0 9812 0 -1 604
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1701704242
transform -1 0 10048 0 -1 605
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1701704242
transform 0 1 1052 1 0 5775
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1701704242
transform 0 -1 12624 1 0 2696
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1701704242
transform 0 -1 10434 1 0 2171
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1701704242
transform 0 -1 12624 1 0 1800
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1701704242
transform 0 -1 11164 1 0 1800
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1701704242
transform 0 -1 10434 1 0 1800
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1701704242
transform 0 -1 10434 1 0 1544
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1701704242
transform 0 -1 12624 1 0 1544
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1701704242
transform 0 -1 10434 1 0 3592
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1701704242
transform 0 -1 11164 1 0 3592
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1701704242
transform 0 -1 10434 1 0 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1701704242
transform 0 -1 12624 1 0 3080
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_45
timestamp 1701704242
transform 0 -1 11164 1 0 3848
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_46
timestamp 1701704242
transform 0 -1 10434 1 0 3848
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_47
timestamp 1701704242
transform 0 -1 11164 1 0 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_48
timestamp 1701704242
transform 0 -1 11894 1 0 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_49
timestamp 1701704242
transform 0 -1 12624 1 0 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_50
timestamp 1701704242
transform 0 -1 10434 1 0 2440
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_51
timestamp 1701704242
transform 0 -1 11164 1 0 1544
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_52
timestamp 1701704242
transform 0 -1 10434 1 0 2952
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_53
timestamp 1701704242
transform 0 -1 369 1 0 5001
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_54
timestamp 1701704242
transform 0 -1 1086 1 0 536
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_55
timestamp 1701704242
transform 1 0 11776 0 -1 3100
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_56
timestamp 1701704242
transform 1 0 11046 0 -1 3100
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_57
timestamp 1701704242
transform 1 0 11776 0 -1 2588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_58
timestamp 1701704242
transform 1 0 11046 0 -1 2588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_59
timestamp 1701704242
transform 1 0 14513 0 -1 5305
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_60
timestamp 1701704242
transform 1 0 13740 0 -1 5500
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_61
timestamp 1701704242
transform 1 0 13740 0 -1 5574
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_62
timestamp 1701704242
transform 1 0 14355 0 -1 5305
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_63
timestamp 1701704242
transform 1 0 7218 0 -1 2785
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_64
timestamp 1701704242
transform 1 0 6970 0 -1 2783
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_65
timestamp 1701704242
transform 1 0 9230 0 -1 2182
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_66
timestamp 1701704242
transform 1 0 6970 0 -1 3096
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_67
timestamp 1701704242
transform 1 0 3894 0 1 2916
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_68
timestamp 1701704242
transform 1 0 11776 0 1 2910
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_69
timestamp 1701704242
transform 1 0 11046 0 1 2910
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_70
timestamp 1701704242
transform 1 0 11046 0 1 2398
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_71
timestamp 1701704242
transform 1 0 11776 0 1 2398
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_72
timestamp 1701704242
transform 1 0 3894 0 1 2548
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_73
timestamp 1701704242
transform 1 0 6508 0 1 -206
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_74
timestamp 1701704242
transform 1 0 9147 0 1 2751
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_75
timestamp 1701704242
transform 1 0 6970 0 1 2390
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_76
timestamp 1701704242
transform 1 0 6970 0 1 2152
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_77
timestamp 1701704242
transform 1 0 7218 0 1 3031
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 1 2484 -1 0 2838
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 1 1752 -1 0 2838
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform -1 0 1340 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1701704242
transform -1 0 1340 0 1 1794
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1701704242
transform -1 0 1340 0 1 3679
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1701704242
transform -1 0 1340 0 1 3501
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1701704242
transform 0 -1 1420 1 0 2559
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1701704242
transform 1 0 2620 0 1 3278
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1701704242
transform 1 0 2620 0 1 1250
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1701704242
transform 1 0 2620 0 1 3902
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1701704242
transform 0 -1 383 -1 0 871
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1701704242
transform 0 -1 1086 -1 0 1851
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1701704242
transform 0 -1 1086 1 0 3478
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_2
timestamp 1701704242
transform 1 0 2620 0 1 3578
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1701704242
transform 0 1 693 1 0 5487
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_1
timestamp 1701704242
transform 1 0 3738 0 -1 377
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_2
timestamp 1701704242
transform 1 0 3744 0 -1 5244
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_3
timestamp 1701704242
transform 1 0 12008 0 1 2220
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_4
timestamp 1701704242
transform 1 0 12008 0 1 3244
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1701704242
transform 1 0 12008 0 1 2732
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_1
timestamp 1701704242
transform 1 0 10620 0 1 3756
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_2
timestamp 1701704242
transform 1 0 10620 0 1 3244
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_3
timestamp 1701704242
transform 1 0 10620 0 1 2732
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_4
timestamp 1701704242
transform 1 0 10620 0 1 2220
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_5
timestamp 1701704242
transform 1 0 10620 0 1 1708
box 0 0 1 1
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_0
timestamp 1701704242
transform 0 1 2484 -1 0 2543
box -12 -6 2062 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_1
timestamp 1701704242
transform 0 1 1752 -1 0 2543
box -12 -6 2062 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_2
timestamp 1701704242
transform 0 1 2484 1 0 2955
box -12 -6 2062 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_3
timestamp 1701704242
transform 0 1 1752 1 0 2955
box -12 -6 2062 40
use L1M1_CDNS_524688791851240  L1M1_CDNS_524688791851240_0
timestamp 1701704242
transform 0 -1 3700 -1 0 743
box -12 -6 406 400
use L1M1_CDNS_524688791851241  L1M1_CDNS_524688791851241_0
timestamp 1701704242
transform 0 -1 3700 1 0 4322
box -12 -6 262 400
use L1M1_CDNS_524688791851241  L1M1_CDNS_524688791851241_1
timestamp 1701704242
transform 0 -1 3700 1 0 3897
box -12 -6 262 400
use L1M1_CDNS_524688791851241  L1M1_CDNS_524688791851241_2
timestamp 1701704242
transform 0 -1 3700 1 0 1352
box -12 -6 262 400
use L1M1_CDNS_524688791851242  L1M1_CDNS_524688791851242_0
timestamp 1701704242
transform 0 -1 3700 1 0 4755
box -12 -6 334 400
use L1M1_CDNS_524688791851243  L1M1_CDNS_524688791851243_0
timestamp 1701704242
transform 0 -1 3706 1 0 1835
box -12 -6 118 400
use L1M1_CDNS_524688791851244  L1M1_CDNS_524688791851244_0
timestamp 1701704242
transform 0 1 3312 1 0 2913
box -12 -6 478 112
use L1M1_CDNS_524688791851244  L1M1_CDNS_524688791851244_1
timestamp 1701704242
transform 0 1 3312 1 0 2118
box -12 -6 478 112
use L1M1_CDNS_524688791851245  L1M1_CDNS_524688791851245_0
timestamp 1701704242
transform 0 -1 3700 1 0 3532
box -12 -6 190 400
use L1M1_CDNS_524688791851245  L1M1_CDNS_524688791851245_1
timestamp 1701704242
transform 0 -1 3700 1 0 1003
box -12 -6 190 400
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 901 -1 0 3331
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 901 -1 0 750
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 2962 -1 0 2965
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 -1 -35 -1 0 6239
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 1 4098 -1 0 5085
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 1 4178 -1 0 3098
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 1 4098 -1 0 2946
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 1 12581 -1 0 3197
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 1 12581 -1 0 2813
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 0 1 10391 -1 0 3965
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 0 1 11121 -1 0 3965
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 0 1 10391 -1 0 3709
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1701704242
transform 0 1 11121 -1 0 3709
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1701704242
transform 0 1 10391 -1 0 3453
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1701704242
transform 0 1 11121 -1 0 3453
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1701704242
transform 0 1 11851 -1 0 3453
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1701704242
transform 0 1 12581 -1 0 3453
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1701704242
transform 0 1 11121 -1 0 1661
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1701704242
transform 0 1 11121 -1 0 1917
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1701704242
transform 0 1 10391 -1 0 2289
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1701704242
transform 0 1 10391 -1 0 1661
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1701704242
transform 0 1 12473 -1 0 3284
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1701704242
transform 0 1 12473 -1 0 2813
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1701704242
transform 0 1 10391 -1 0 2557
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1701704242
transform 0 1 10391 -1 0 1917
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1701704242
transform 0 1 10474 -1 0 1789
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1701704242
transform 0 1 10474 -1 0 3837
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1701704242
transform 0 1 10474 -1 0 3325
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1701704242
transform 0 1 10474 -1 0 2301
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1701704242
transform 0 1 10474 -1 0 2813
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1701704242
transform 0 1 4418 -1 0 3837
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1701704242
transform 0 1 4418 -1 0 3238
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1701704242
transform 0 1 4178 -1 0 4122
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_33
timestamp 1701704242
transform 0 1 240 -1 0 3500
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_34
timestamp 1701704242
transform 0 1 687 -1 0 1388
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_35
timestamp 1701704242
transform 0 1 687 -1 0 4747
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_36
timestamp 1701704242
transform 0 1 769 -1 0 3672
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_37
timestamp 1701704242
transform 0 1 769 -1 0 1102
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_38
timestamp 1701704242
transform 0 1 769 -1 0 750
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_39
timestamp 1701704242
transform -1 0 2694 0 1 4973
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_40
timestamp 1701704242
transform -1 0 2694 0 1 4517
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_41
timestamp 1701704242
transform -1 0 2694 0 1 929
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_42
timestamp 1701704242
transform -1 0 2694 0 1 473
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_43
timestamp 1701704242
transform -1 0 1343 0 -1 5252
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_44
timestamp 1701704242
transform -1 0 821 0 -1 4983
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_45
timestamp 1701704242
transform -1 0 7168 0 -1 2510
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_46
timestamp 1701704242
transform -1 0 7085 0 -1 2795
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_47
timestamp 1701704242
transform 0 1 2830 1 0 3658
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_48
timestamp 1701704242
transform 0 1 2830 1 0 4011
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_49
timestamp 1701704242
transform 0 1 2830 1 0 4282
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_50
timestamp 1701704242
transform 0 1 4098 1 0 1844
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_51
timestamp 1701704242
transform 0 1 2910 1 0 3231
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_52
timestamp 1701704242
transform 0 1 2910 1 0 2657
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_53
timestamp 1701704242
transform 0 1 2990 1 0 2139
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_54
timestamp 1701704242
transform 0 1 2990 1 0 1827
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_55
timestamp 1701704242
transform 0 1 2990 1 0 2818
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_56
timestamp 1701704242
transform 0 1 4418 1 0 1661
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_57
timestamp 1701704242
transform 0 1 2475 1 0 2722
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_58
timestamp 1701704242
transform 0 1 2830 1 0 2295
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_59
timestamp 1701704242
transform 0 1 2830 1 0 1983
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_60
timestamp 1701704242
transform 0 1 2830 1 0 1712
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_61
timestamp 1701704242
transform 0 1 2830 1 0 1359
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_62
timestamp 1701704242
transform 0 1 2830 1 0 1088
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_63
timestamp 1701704242
transform 0 1 2910 1 0 3531
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_64
timestamp 1701704242
transform 0 1 4178 1 0 1088
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_65
timestamp 1701704242
transform 0 1 12473 1 0 2214
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_66
timestamp 1701704242
transform 0 1 10391 1 0 2941
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_67
timestamp 1701704242
transform 0 1 2830 1 0 3387
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_68
timestamp 1701704242
transform 0 1 2830 1 0 3075
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_69
timestamp 1701704242
transform 0 1 4418 1 0 2260
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_70
timestamp 1701704242
transform 0 1 2910 1 0 2423
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_71
timestamp 1701704242
transform 0 1 4098 1 0 2552
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_72
timestamp 1701704242
transform 0 1 2750 1 0 2722
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_73
timestamp 1701704242
transform 0 1 240 1 0 2855
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_74
timestamp 1701704242
transform 0 1 849 1 0 2055
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_75
timestamp 1701704242
transform 0 1 2990 1 0 2583
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_76
timestamp 1701704242
transform 0 1 4178 1 0 2370
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_77
timestamp 1701704242
transform 0 1 240 1 0 1908
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_78
timestamp 1701704242
transform 0 -1 2802 1 0 5394
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_79
timestamp 1701704242
transform 0 -1 901 1 0 2919
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_80
timestamp 1701704242
transform 0 -1 901 1 0 4677
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_81
timestamp 1701704242
transform 0 -1 901 1 0 1442
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_82
timestamp 1701704242
transform 0 -1 901 1 0 1899
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_83
timestamp 1701704242
transform 0 -1 1095 1 0 5413
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_84
timestamp 1701704242
transform 0 -1 7092 1 0 2980
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_85
timestamp 1701704242
transform 1 0 4118 0 -1 5252
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_86
timestamp 1701704242
transform 1 0 7126 0 -1 3071
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_87
timestamp 1701704242
transform 1 0 7126 0 -1 2791
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_88
timestamp 1701704242
transform 1 0 7126 0 -1 2430
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_89
timestamp 1701704242
transform 1 0 423 0 1 2814
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1701704242
transform 0 1 1769 1 0 5324
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1701704242
transform -1 0 14001 0 -1 5162
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1701704242
transform -1 0 14001 0 -1 6907
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1701704242
transform 0 1 2475 -1 0 2555
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1701704242
transform -1 0 4070 0 1 2539
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1701704242
transform -1 0 4070 0 1 2139
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1701704242
transform -1 0 4070 0 1 4738
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_4
timestamp 1701704242
transform -1 0 521 0 1 1986
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_5
timestamp 1701704242
transform -1 0 4070 0 1 2343
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_6
timestamp 1701704242
transform -1 0 4070 0 1 3103
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_7
timestamp 1701704242
transform -1 0 4070 0 1 2907
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_8
timestamp 1701704242
transform -1 0 1342 0 1 2484
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_9
timestamp 1701704242
transform -1 0 1342 0 1 2300
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_10
timestamp 1701704242
transform -1 0 1342 0 1 2668
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_11
timestamp 1701704242
transform -1 0 1342 0 1 2116
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_12
timestamp 1701704242
transform -1 0 619 0 1 443
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_13
timestamp 1701704242
transform -1 0 631 0 1 795
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_14
timestamp 1701704242
transform -1 0 631 0 1 4772
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_15
timestamp 1701704242
transform -1 0 631 0 1 1147
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_16
timestamp 1701704242
transform -1 0 631 0 1 5742
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_17
timestamp 1701704242
transform -1 0 631 0 1 5390
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_18
timestamp 1701704242
transform -1 0 631 0 1 6094
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_19
timestamp 1701704242
transform -1 0 631 0 1 5038
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_20
timestamp 1701704242
transform -1 0 4070 0 1 3307
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_21
timestamp 1701704242
transform -1 0 4070 0 1 4337
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_22
timestamp 1701704242
transform -1 0 4070 0 1 4021
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_23
timestamp 1701704242
transform -1 0 4070 0 1 3711
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_24
timestamp 1701704242
transform -1 0 4070 0 1 630
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_25
timestamp 1701704242
transform -1 0 4070 0 1 940
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_26
timestamp 1701704242
transform -1 0 4070 0 1 1256
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_27
timestamp 1701704242
transform -1 0 631 0 1 2630
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_28
timestamp 1701704242
transform -1 0 631 0 1 2364
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_29
timestamp 1701704242
transform -1 0 631 0 1 3200
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_30
timestamp 1701704242
transform -1 0 1342 0 -1 2922
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_31
timestamp 1701704242
transform -1 0 1342 0 -1 3216
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_32
timestamp 1701704242
transform -1 0 1342 0 -1 3464
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_33
timestamp 1701704242
transform -1 0 1342 0 -1 3633
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_34
timestamp 1701704242
transform -1 0 1342 0 -1 3811
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_35
timestamp 1701704242
transform -1 0 1342 0 -1 1570
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_36
timestamp 1701704242
transform -1 0 1342 0 -1 1748
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_37
timestamp 1701704242
transform -1 0 1342 0 -1 1917
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_38
timestamp 1701704242
transform 0 1 2475 1 0 2943
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 0 1 2750 1 0 837
box 0 0 1 1
use M1M2_CDNS_52468879185958  M1M2_CDNS_52468879185958_0
timestamp 1701704242
transform 0 1 3220 1 0 991
box 0 0 192 436
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_0
timestamp 1701704242
transform 0 -1 4067 1 0 5124
box 0 0 128 308
use M1M2_CDNS_524688791851176  M1M2_CDNS_524688791851176_0
timestamp 1701704242
transform 0 -1 3528 1 0 4319
box 0 0 256 308
use M1M2_CDNS_524688791851176  M1M2_CDNS_524688791851176_1
timestamp 1701704242
transform 0 -1 3528 1 0 3894
box 0 0 256 308
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1701704242
transform 0 1 1570 1 0 5670
box 0 0 384 116
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_0
timestamp 1701704242
transform 0 -1 3528 1 0 3530
box 0 0 192 308
use M1M2_CDNS_524688791851246  M1M2_CDNS_524688791851246_0
timestamp 1701704242
transform 0 -1 3528 1 0 4752
box 0 0 320 308
use M1M2_CDNS_524688791851247  M1M2_CDNS_524688791851247_0
timestamp 1701704242
transform 0 1 3220 1 0 1349
box 0 0 256 436
use M1M2_CDNS_524688791851248  M1M2_CDNS_524688791851248_0
timestamp 1701704242
transform 0 1 3220 1 0 371
box 0 0 384 436
use M1M2_CDNS_524688791851249  M1M2_CDNS_524688791851249_0
timestamp 1701704242
transform 0 1 3220 1 0 1824
box 0 0 128 436
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_0
timestamp 1701704242
transform 0 -1 3400 1 0 2922
box 0 0 448 180
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_1
timestamp 1701704242
transform 0 -1 3400 1 0 2127
box 0 0 448 180
use nDFres_CDNS_524688791851251  nDFres_CDNS_524688791851251_0
timestamp 1701704242
transform -1 0 10844 0 1 191
box -68 -26 374 162
use nDFres_CDNS_524688791851251  nDFres_CDNS_524688791851251_1
timestamp 1701704242
transform -1 0 10065 0 1 191
box -68 -26 374 162
use nDFres_CDNS_524688791851251  nDFres_CDNS_524688791851251_2
timestamp 1701704242
transform -1 0 12570 0 1 191
box -68 -26 374 162
use nDFres_CDNS_524688791851251  nDFres_CDNS_524688791851251_3
timestamp 1701704242
transform -1 0 11603 0 1 191
box -68 -26 374 162
use nDFres_CDNS_524688791851253  nDFres_CDNS_524688791851253_0
timestamp 1701704242
transform -1 0 8307 0 1 -147
box -68 -26 1749 162
use nDFres_CDNS_524688791851253  nDFres_CDNS_524688791851253_1
timestamp 1701704242
transform -1 0 12574 0 1 -147
box -68 -26 1749 162
use nfet_CDNS_524688791851308  nfet_CDNS_524688791851308_0
timestamp 1701704242
transform 1 0 10205 0 1 11370
box -79 -26 1735 626
use nfet_CDNS_524688791851309  nfet_CDNS_524688791851309_0
timestamp 1701704242
transform 1 0 6488 0 1 9602
box -79 -26 3447 626
use nfet_CDNS_524688791851310  nfet_CDNS_524688791851310_0
timestamp 1701704242
transform 1 0 6488 0 1 8872
box -79 -26 3447 626
use nfet_CDNS_524688791851311  nfet_CDNS_524688791851311_0
timestamp 1701704242
transform 1 0 6488 0 1 10479
box -79 -26 5159 626
use nfet_CDNS_524688791851312  nfet_CDNS_524688791851312_0
timestamp 1701704242
transform 0 -1 11812 -1 0 4001
box -79 -26 279 626
use nfet_CDNS_524688791851312  nfet_CDNS_524688791851312_1
timestamp 1701704242
transform 0 -1 11812 1 0 1497
box -79 -26 279 626
use nfet_CDNS_524688791851313  nfet_CDNS_524688791851313_0
timestamp 1701704242
transform 0 -1 11812 1 0 641
box -79 -26 879 626
use nfet_CDNS_524688791851313  nfet_CDNS_524688791851313_1
timestamp 1701704242
transform 0 -1 11812 1 0 4057
box -79 -26 879 626
use nfet_CDNS_524688791851314  nfet_CDNS_524688791851314_0
timestamp 1701704242
transform 0 -1 11812 -1 0 1953
box -79 -26 279 626
use nfet_CDNS_524688791851314  nfet_CDNS_524688791851314_1
timestamp 1701704242
transform 0 -1 11812 1 0 3545
box -79 -26 279 626
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_0
timestamp 1701704242
transform 0 -1 9266 -1 0 2533
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_1
timestamp 1701704242
transform 0 -1 9266 -1 0 3131
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_2
timestamp 1701704242
transform 0 -1 9266 -1 0 3491
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_3
timestamp 1701704242
transform 0 -1 9266 -1 0 1937
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_4
timestamp 1701704242
transform 0 1 5028 -1 0 3131
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_5
timestamp 1701704242
transform 0 1 5028 -1 0 2533
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_6
timestamp 1701704242
transform 0 1 5028 -1 0 3491
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_7
timestamp 1701704242
transform 0 1 5028 -1 0 1937
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_8
timestamp 1701704242
transform 0 1 5028 1 0 2117
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_9
timestamp 1701704242
transform 0 1 5028 1 0 2715
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_10
timestamp 1701704242
transform 0 -1 9266 1 0 2715
box -79 -52 259 2052
use nfet_CDNS_524688791851315  nfet_CDNS_524688791851315_11
timestamp 1701704242
transform 0 -1 9266 1 0 2117
box -79 -52 259 2052
use nfet_CDNS_524688791851316  nfet_CDNS_524688791851316_0
timestamp 1701704242
transform -1 0 9848 0 1 679
box -82 -52 262 2052
use nfet_CDNS_524688791851316  nfet_CDNS_524688791851316_1
timestamp 1701704242
transform -1 0 10084 0 1 679
box -82 -52 262 2052
use nfet_CDNS_524688791851316  nfet_CDNS_524688791851316_2
timestamp 1701704242
transform -1 0 10084 0 1 2879
box -82 -52 262 2052
use nfet_CDNS_524688791851316  nfet_CDNS_524688791851316_3
timestamp 1701704242
transform -1 0 9848 0 1 2879
box -82 -52 262 2052
use nfet_CDNS_524688791851317  nfet_CDNS_524688791851317_0
timestamp 1701704242
transform 0 1 3898 -1 0 4022
box -79 -26 491 226
use nfet_CDNS_524688791851317  nfet_CDNS_524688791851317_1
timestamp 1701704242
transform 0 1 3898 1 0 997
box -79 -26 491 226
use nfet_CDNS_524688791851318  nfet_CDNS_524688791851318_0
timestamp 1701704242
transform 0 1 3898 -1 0 941
box -79 -26 491 226
use nfet_CDNS_524688791851318  nfet_CDNS_524688791851318_1
timestamp 1701704242
transform 0 1 3898 1 0 4078
box -79 -26 491 226
use nfet_CDNS_524688791851319  nfet_CDNS_524688791851319_0
timestamp 1701704242
transform 0 1 3898 -1 0 3101
box -79 -26 115 226
use nfet_CDNS_524688791851320  nfet_CDNS_524688791851320_0
timestamp 1701704242
transform 0 -1 11812 1 0 2009
box -79 -26 1559 626
use nfet_CDNS_524688791851321  nfet_CDNS_524688791851321_0
timestamp 1701704242
transform 0 -1 12542 1 0 641
box -79 -26 879 626
use nfet_CDNS_524688791851321  nfet_CDNS_524688791851321_1
timestamp 1701704242
transform 0 -1 11082 1 0 4057
box -79 -26 879 626
use nfet_CDNS_524688791851321  nfet_CDNS_524688791851321_2
timestamp 1701704242
transform 0 -1 11082 1 0 641
box -79 -26 879 626
use nfet_CDNS_524688791851321  nfet_CDNS_524688791851321_3
timestamp 1701704242
transform 0 -1 12542 1 0 4057
box -79 -26 879 626
use nfet_CDNS_524688791851322  nfet_CDNS_524688791851322_0
timestamp 1701704242
transform 0 -1 11082 1 0 1497
box -79 -26 2583 626
use nfet_CDNS_524688791851323  nfet_CDNS_524688791851323_0
timestamp 1701704242
transform 0 -1 12542 1 0 3033
box -79 -26 535 626
use nfet_CDNS_524688791851324  nfet_CDNS_524688791851324_0
timestamp 1701704242
transform 0 -1 12542 1 0 2009
box -79 -26 535 626
use nfet_CDNS_524688791851324  nfet_CDNS_524688791851324_1
timestamp 1701704242
transform 0 -1 12542 1 0 2521
box -79 -26 535 626
use nfet_CDNS_524688791851325  nfet_CDNS_524688791851325_0
timestamp 1701704242
transform 0 -1 1336 -1 0 3162
box -79 -26 115 226
use nfet_CDNS_524688791851325  nfet_CDNS_524688791851325_1
timestamp 1701704242
transform 0 1 3898 1 0 2397
box -79 -26 115 226
use nfet_CDNS_524688791851325  nfet_CDNS_524688791851325_2
timestamp 1701704242
transform 0 -1 1336 1 0 2924
box -79 -26 115 226
use nfet_CDNS_524688791851326  nfet_CDNS_524688791851326_0
timestamp 1701704242
transform 0 1 3948 -1 0 2137
box -79 -26 239 176
use nfet_CDNS_524688791851326  nfet_CDNS_524688791851326_1
timestamp 1701704242
transform 0 1 3948 1 0 4792
box -79 -26 239 176
use nfet_CDNS_524688791851327  nfet_CDNS_524688791851327_0
timestamp 1701704242
transform 0 1 433 -1 0 1145
box -79 -26 727 226
use nfet_CDNS_524688791851328  nfet_CDNS_524688791851328_0
timestamp 1701704242
transform 0 -1 1336 1 0 3218
box -79 -26 115 226
use nfet_CDNS_524688791851328  nfet_CDNS_524688791851328_1
timestamp 1701704242
transform 0 -1 1336 1 0 2170
box -79 -26 115 226
use nfet_CDNS_524688791851329  nfet_CDNS_524688791851329_0
timestamp 1701704242
transform 0 -1 1336 -1 0 5740
box -79 -26 199 226
use nfet_CDNS_524688791851330  nfet_CDNS_524688791851330_0
timestamp 1701704242
transform 0 -1 1336 1 0 5796
box -79 -26 375 226
use nfet_CDNS_524688791851331  nfet_CDNS_524688791851331_0
timestamp 1701704242
transform 0 -1 1336 -1 0 4832
box -79 -26 967 226
use nfet_CDNS_524688791851332  nfet_CDNS_524688791851332_0
timestamp 1701704242
transform 0 1 433 -1 0 4149
box -79 -26 551 226
use nfet_CDNS_524688791851332  nfet_CDNS_524688791851332_1
timestamp 1701704242
transform 0 1 433 -1 0 1783
box -79 -26 551 226
use nfet_CDNS_524688791851333  nfet_CDNS_524688791851333_0
timestamp 1701704242
transform 0 -1 1336 -1 0 2482
box -79 -26 299 226
use nfet_CDNS_524688791851333  nfet_CDNS_524688791851333_1
timestamp 1701704242
transform 0 -1 1336 1 0 2538
box -79 -26 299 226
use nfet_CDNS_524688791851334  nfet_CDNS_524688791851334_0
timestamp 1701704242
transform 0 1 3898 1 0 2593
box -79 -26 115 226
use nfet_CDNS_524688791851335  nfet_CDNS_524688791851335_0
timestamp 1701704242
transform 0 1 3898 -1 0 2905
box -79 -26 115 226
use nfet_CDNS_524688791851336  nfet_CDNS_524688791851336_0
timestamp 1701704242
transform 0 -1 1336 -1 0 1863
box -79 -26 367 226
use nfet_CDNS_524688791851336  nfet_CDNS_524688791851336_1
timestamp 1701704242
transform 0 -1 1336 -1 0 3754
box -79 -26 367 226
use nfet_CDNS_524688791851337  nfet_CDNS_524688791851337_0
timestamp 1701704242
transform 0 -1 1336 -1 0 5198
box -79 -26 279 176
use nfet_CDNS_524688791851338  nfet_CDNS_524688791851338_0
timestamp 1701704242
transform 0 -1 1336 1 0 5254
box -79 -26 279 176
use nfet_CDNS_524688791851339  nfet_CDNS_524688791851339_0
timestamp 1701704242
transform 0 -1 1336 -1 0 1385
box -79 -26 967 226
use pfet_CDNS_524688791851340  pfet_CDNS_524688791851340_0
timestamp 1701704242
transform 0 1 1836 1 0 497
box -119 -66 4623 666
use pfet_CDNS_524688791851341  pfet_CDNS_524688791851341_0
timestamp 1701704242
transform 0 -1 2866 -1 0 4515
box -119 -66 219 366
use pfet_CDNS_524688791851341  pfet_CDNS_524688791851341_1
timestamp 1701704242
transform 0 -1 2866 -1 0 2487
box -119 -66 219 366
use pfet_CDNS_524688791851341  pfet_CDNS_524688791851341_2
timestamp 1701704242
transform 0 -1 2866 1 0 2543
box -119 -66 219 366
use pfet_CDNS_524688791851341  pfet_CDNS_524688791851341_3
timestamp 1701704242
transform 0 -1 2866 1 0 3011
box -119 -66 219 366
use pfet_CDNS_524688791851341  pfet_CDNS_524688791851341_4
timestamp 1701704242
transform 0 -1 2866 1 0 983
box -119 -66 219 366
use pfet_CDNS_524688791851342  pfet_CDNS_524688791851342_0
timestamp 1701704242
transform 0 -1 2866 1 0 2699
box -119 -66 375 366
use pfet_CDNS_524688791851342  pfet_CDNS_524688791851342_1
timestamp 1701704242
transform 0 -1 2866 1 0 1451
box -119 -66 375 366
use pfet_CDNS_524688791851342  pfet_CDNS_524688791851342_2
timestamp 1701704242
transform 0 -1 2866 1 0 1763
box -119 -66 375 366
use pfet_CDNS_524688791851342  pfet_CDNS_524688791851342_3
timestamp 1701704242
transform 0 -1 2866 1 0 2075
box -119 -66 375 366
use pfet_CDNS_524688791851342  pfet_CDNS_524688791851342_4
timestamp 1701704242
transform 0 -1 2866 1 0 4103
box -119 -66 375 366
use pfet_CDNS_524688791851343  pfet_CDNS_524688791851343_0
timestamp 1701704242
transform 0 -1 2866 1 0 4571
box -119 -66 519 366
use pfet_CDNS_524688791851343  pfet_CDNS_524688791851343_1
timestamp 1701704242
transform 0 -1 2866 1 0 527
box -119 -66 519 366
use pfet_CDNS_524688791851344  pfet_CDNS_524688791851344_0
timestamp 1701704242
transform 0 -1 2866 1 0 1139
box -119 -66 375 366
use pfet_CDNS_524688791851344  pfet_CDNS_524688791851344_1
timestamp 1701704242
transform 0 -1 2866 1 0 3479
box -119 -66 375 366
use pfet_CDNS_524688791851344  pfet_CDNS_524688791851344_2
timestamp 1701704242
transform 0 -1 2866 1 0 3167
box -119 -66 375 366
use pfet_CDNS_524688791851344  pfet_CDNS_524688791851344_3
timestamp 1701704242
transform 0 -1 2866 1 0 3791
box -119 -66 375 366
use pfet_CDNS_524688791851345  pfet_CDNS_524688791851345_0
timestamp 1701704242
transform 0 1 433 1 0 5092
box -119 -66 415 266
use pfet_CDNS_524688791851346  pfet_CDNS_524688791851346_0
timestamp 1701704242
transform 0 1 433 1 0 5444
box -119 -66 767 266
use pfet_CDNS_524688791851347  pfet_CDNS_524688791851347_0
timestamp 1701704242
transform 0 1 445 -1 0 2362
box -89 -36 189 236
use pfet_CDNS_524688791851348  pfet_CDNS_524688791851348_0
timestamp 1701704242
transform 0 -1 583 -1 0 4770
box -119 -66 219 216
use pfet_CDNS_524688791851348  pfet_CDNS_524688791851348_1
timestamp 1701704242
transform 0 -1 583 1 0 4826
box -119 -66 219 216
use pfet_CDNS_524688791851349  pfet_CDNS_524688791851349_0
timestamp 1701704242
transform 0 1 445 -1 0 3198
box -89 -36 125 236
use pfet_CDNS_524688791851349  pfet_CDNS_524688791851349_1
timestamp 1701704242
transform 0 1 445 1 0 2960
box -89 -36 125 236
use pfet_CDNS_524688791851350  pfet_CDNS_524688791851350_0
timestamp 1701704242
transform 0 1 445 1 0 2684
box -89 -36 309 236
use pfet_CDNS_524688791851351  pfet_CDNS_524688791851351_0
timestamp 1701704242
transform 0 1 445 -1 0 2518
box -89 -36 189 236
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform 0 -1 3600 -1 0 2171
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1701704242
transform 0 -1 3600 1 0 3276
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1701704242
transform 1 0 2898 0 1 4432
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1701704242
transform 1 0 2898 0 1 3028
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1701704242
transform 1 0 2898 0 1 2566
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1701704242
transform 1 0 2898 0 1 1000
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1701704242
transform 0 1 9928 -1 0 5003
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1701704242
transform 0 1 9692 -1 0 5003
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1701704242
transform 0 1 9692 -1 0 620
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1701704242
transform 0 1 9928 -1 0 621
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1701704242
transform -1 0 1102 0 1 2924
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1701704242
transform -1 0 1102 0 1 2072
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1701704242
transform -1 0 11180 0 -1 1664
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1701704242
transform -1 0 12640 0 -1 1664
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1701704242
transform -1 0 11180 0 -1 1920
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1701704242
transform -1 0 12640 0 -1 1920
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1701704242
transform -1 0 11180 0 -1 2176
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_11
timestamp 1701704242
transform -1 0 11910 0 -1 2176
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_12
timestamp 1701704242
transform -1 0 12640 0 -1 2176
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_13
timestamp 1701704242
transform -1 0 11180 0 -1 2432
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_14
timestamp 1701704242
transform -1 0 11910 0 -1 2432
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_15
timestamp 1701704242
transform -1 0 11180 0 -1 2688
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_16
timestamp 1701704242
transform -1 0 11910 0 -1 2688
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_17
timestamp 1701704242
transform -1 0 12640 0 -1 2688
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_18
timestamp 1701704242
transform -1 0 11180 0 -1 2944
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_19
timestamp 1701704242
transform -1 0 11910 0 -1 2944
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_20
timestamp 1701704242
transform -1 0 12640 0 -1 2944
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_21
timestamp 1701704242
transform -1 0 11180 0 -1 3200
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_22
timestamp 1701704242
transform -1 0 11910 0 -1 3200
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_23
timestamp 1701704242
transform -1 0 11180 0 -1 3456
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_24
timestamp 1701704242
transform -1 0 11910 0 -1 3456
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_25
timestamp 1701704242
transform -1 0 12640 0 -1 3456
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_26
timestamp 1701704242
transform -1 0 11180 0 -1 3712
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_27
timestamp 1701704242
transform -1 0 11180 0 -1 3968
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_28
timestamp 1701704242
transform -1 0 12640 0 -1 3200
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_29
timestamp 1701704242
transform -1 0 413 0 -1 2362
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_30
timestamp 1701704242
transform -1 0 1102 0 -1 3352
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_31
timestamp 1701704242
transform -1 0 399 0 -1 3198
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_32
timestamp 1701704242
transform -1 0 9364 0 -1 2872
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_33
timestamp 1701704242
transform -1 0 9364 0 -1 2510
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_34
timestamp 1701704242
transform -1 0 9364 0 -1 3108
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_35
timestamp 1701704242
transform -1 0 9364 0 -1 2274
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_36
timestamp 1701704242
transform -1 0 7126 0 -1 2510
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_37
timestamp 1701704242
transform -1 0 7126 0 -1 2872
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_38
timestamp 1701704242
transform -1 0 9364 0 -1 1914
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_39
timestamp 1701704242
transform -1 0 9364 0 -1 3468
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_40
timestamp 1701704242
transform -1 0 7126 0 -1 2274
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_41
timestamp 1701704242
transform -1 0 7126 0 -1 3108
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_42
timestamp 1701704242
transform 0 -1 3032 1 0 2420
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_43
timestamp 1701704242
transform 1 0 10384 0 -1 1664
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_44
timestamp 1701704242
transform 1 0 10384 0 -1 1920
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_45
timestamp 1701704242
transform 1 0 10384 0 -1 2176
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_46
timestamp 1701704242
transform 1 0 10384 0 -1 2432
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_47
timestamp 1701704242
transform 1 0 10384 0 -1 2688
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_48
timestamp 1701704242
transform 1 0 10384 0 -1 2944
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_49
timestamp 1701704242
transform 1 0 10384 0 -1 3200
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_50
timestamp 1701704242
transform 1 0 10384 0 -1 3456
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_51
timestamp 1701704242
transform 1 0 10384 0 -1 3712
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_52
timestamp 1701704242
transform 1 0 10384 0 -1 3968
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_53
timestamp 1701704242
transform 1 0 4930 0 -1 2877
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_54
timestamp 1701704242
transform 1 0 677 0 -1 3094
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_55
timestamp 1701704242
transform 1 0 4930 0 -1 3113
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_56
timestamp 1701704242
transform 1 0 7168 0 -1 2510
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_57
timestamp 1701704242
transform 1 0 4930 0 -1 3468
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_58
timestamp 1701704242
transform 1 0 4930 0 -1 2510
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_59
timestamp 1701704242
transform 1 0 4930 0 -1 2274
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_60
timestamp 1701704242
transform 1 0 7168 0 -1 2872
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_61
timestamp 1701704242
transform 1 0 7168 0 -1 2274
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_62
timestamp 1701704242
transform 1 0 7168 0 -1 3108
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_63
timestamp 1701704242
transform 1 0 4930 0 -1 1914
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_64
timestamp 1701704242
transform 1 0 677 0 1 2418
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_65
timestamp 1701704242
transform 1 0 1370 0 1 3028
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1701704242
transform -1 0 12640 0 -1 3908
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1701704242
transform -1 0 12640 0 -1 1414
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_1
timestamp 1701704242
transform -1 0 11180 0 -1 1414
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_2
timestamp 1701704242
transform -1 0 11910 0 -1 1414
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_3
timestamp 1701704242
transform -1 0 11180 0 -1 4830
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_4
timestamp 1701704242
transform -1 0 11910 0 -1 4830
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_5
timestamp 1701704242
transform -1 0 12640 0 -1 4830
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_6
timestamp 1701704242
transform 1 0 10384 0 -1 1414
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_7
timestamp 1701704242
transform 1 0 10384 0 -1 4830
box 0 0 66 746
use PYres_CDNS_524688791851352  PYres_CDNS_524688791851352_0
timestamp 1701704242
transform 0 1 3534 1 0 2155
box -50 0 1187 66
use sky130_fd_io__sio_biasgen  sky130_fd_io__sio_biasgen_0
timestamp 1701704242
transform 1 0 751 0 1 -1274
box -631 681 14756 14857
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1701704242
transform 1 0 1702 0 1 10579
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_0
timestamp 1701704242
transform 1 0 1996 0 1 10579
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_inv_x4  sky130_fd_io__sio_hvsbt_inv_x4_0
timestamp 1701704242
transform 1 0 2572 0 1 10579
box -107 21 811 1369
use sky130_fd_io__sio_in_diff_iclmp  sky130_fd_io__sio_in_diff_iclmp_0
timestamp 1701704242
transform 1 0 14148 0 1 5419
box -2092 -378 2348 5075
use sky130_fd_io__sio_in_diff_localesd  sky130_fd_io__sio_in_diff_localesd_0
timestamp 1701704242
transform -1 0 16429 0 1 0
box -429 -66 3479 5505
use sky130_fd_io__sio_in_diff_res_9k  sky130_fd_io__sio_in_diff_res_9k_0
timestamp 1701704242
transform -1 0 9386 0 1 1313
box 14 -378 4446 118
use sky130_fd_io__sio_in_diff_res_9k  sky130_fd_io__sio_in_diff_res_9k_1
timestamp 1701704242
transform -1 0 9386 0 -1 4026
box 14 -378 4446 118
use sky130_fd_io__sio_in_diff_res_40k  sky130_fd_io__sio_in_diff_res_40k_0
timestamp 1701704242
transform -1 0 9372 0 1 402
box 0 -159 4432 4742
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_0
timestamp 1701704242
transform -1 0 12298 0 1 224
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_1
timestamp 1701704242
transform 1 0 11637 0 1 224
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_0
timestamp 1701704242
transform -1 0 11972 0 1 3238
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_1
timestamp 1701704242
transform -1 0 11972 0 1 2214
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_2
timestamp 1701704242
transform -1 0 2934 0 1 3896
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_3
timestamp 1701704242
transform 1 0 2802 0 -1 1290
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_4
timestamp 1701704242
transform 1 0 2777 0 1 3272
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_5
timestamp 1701704242
transform 1 0 2857 0 1 2180
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851307  sky130_fd_io__sio_tk_em1o_CDNS_524688791851307_0
timestamp 1701704242
transform 0 -1 7014 -1 0 3640
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851307  sky130_fd_io__sio_tk_em1o_CDNS_524688791851307_1
timestamp 1701704242
transform 0 -1 7014 1 0 1594
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1701704242
transform -1 0 10810 0 1 235
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1701704242
transform 1 0 9282 0 -1 2590
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_2
timestamp 1701704242
transform 1 0 9858 0 1 235
box 0 0 1 1
<< labels >>
flabel comment s 8184 2327 8184 2327 0 FreeSans 1000 0 0 0 I1735
flabel comment s 8171 2947 8171 2947 0 FreeSans 1000 0 0 0 ndiffref
flabel comment s 6065 2345 6065 2345 0 FreeSans 1000 0 0 0 I1736
flabel comment s 6011 2936 6011 2936 0 FreeSans 1000 0 0 0 ndiffin
flabel comment s 4661 5250 4661 5250 0 FreeSans 400 90 0 0 lv_net
flabel comment s 5409 5178 5409 5178 0 FreeSans 400 0 0 0 condiode
flabel comment s 6930 10413 6930 10413 3 FreeSans 200 90 0 0 od_h
flabel comment s 3622 8334 3622 8334 3 FreeSans 200 0 0 0 od_h
flabel comment s 1687 -63 1687 -63 3 FreeSans 200 90 0 0 pad_a_noesd_h
flabel comment s 1788 -63 1788 -63 3 FreeSans 200 90 0 0 pad_a_esd_h
flabel comment s 2556 5552 2556 5552 3 FreeSans 200 180 0 0 pad_a_esd_h
flabel comment s 2572 6053 2572 6053 3 FreeSans 200 180 0 0 pad_a_noesd_h
flabel comment s 1386 6093 1386 6093 0 FreeSans 200 0 0 0 vgnd
flabel comment s 1226 6224 1226 6224 0 FreeSans 200 0 0 0 vnb
flabel comment s 595 6263 595 6263 0 FreeSans 200 0 0 0 vcc_ioq
flabel comment s 2926 2556 2926 2556 0 FreeSans 200 0 0 0 ie_diff_sel_h
flabel comment s 2778 5266 2778 5266 0 FreeSans 200 90 0 0 ie_diff_sel_h
flabel comment s 6011 2941 6011 2941 0 FreeSans 1000 0 0 0 ndiffin
flabel comment s 12313 4031 12313 4031 0 FreeSans 400 0 0 0 vgnd
flabel comment s 13359 11250 13359 11250 0 FreeSans 400 90 0 0 lv_net
flabel comment s 12618 3476 12618 3476 0 FreeSans 400 90 0 0 ngate
flabel comment s 12273 3516 12273 3516 0 FreeSans 400 0 0 0 vgnd
flabel metal1 s 7125 2089 7125 2089 0 FreeSans 100 0 0 0 ndiffcom
flabel metal1 s 0 2595 42 2799 0 FreeSans 200 90 0 0 vpb
port 6 nsew
flabel metal1 s 9586 8742 9678 8788 3 FreeSans 520 0 0 0 vgnd
port 2 nsew
flabel metal1 s 2931 6241 2983 6300 3 FreeSans 520 0 0 0 ie_diff_sel_n
port 3 nsew
flabel metal1 s 7927 5624 8019 5670 3 FreeSans 520 0 0 0 vgnd
port 2 nsew
flabel metal1 s 1754 10892 2074 10940 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 10715 8983 10775 9029 3 FreeSans 520 0 0 0 vpwr
port 4 nsew
flabel metal1 s 212 12980 272 13026 3 FreeSans 520 0 0 0 vpwr
port 4 nsew
flabel metal1 s 15265 13446 15325 13492 3 FreeSans 520 0 0 0 vpwr
port 4 nsew
flabel metal1 s 5786 11457 5878 11563 3 FreeSans 520 0 0 0 vgnd
port 2 nsew
flabel metal1 s 1782 11337 2102 11385 0 FreeSans 400 180 0 0 vcc_io
port 5 nsew
flabel metal1 s 0 2364 42 2567 0 FreeSans 200 90 0 0 vpwr
port 4 nsew
flabel metal1 s 0 3018 59 3344 3 FreeSans 200 0 0 0 vpb
port 6 nsew
flabel metal1 s 0 1953 56 2020 3 FreeSans 200 0 0 0 ie_diff_dly_n
port 12 nsew
flabel metal1 s 16501 5106 16553 5157 0 FreeSans 400 180 0 0 vinref
port 7 nsew
flabel metal1 s 0 1099 54 1145 3 FreeSans 200 0 0 0 ie_diff_sel_h_n
port 11 nsew
flabel metal1 s 0 5147 53 5189 3 FreeSans 200 0 0 0 ie_diff_n
port 8 nsew
flabel metal1 s 8 3610 51 3664 3 FreeSans 200 0 0 0 ie_diff_sel_h
port 9 nsew
flabel metal1 s 2 1809 28 1880 3 FreeSans 200 0 0 0 ie_diff_sel_h
port 9 nsew
flabel metal1 s 0 944 28 972 3 FreeSans 200 0 0 0 out
port 10 nsew
flabel metal1 s 0 2094 42 2336 0 FreeSans 200 90 0 0 vpb
port 6 nsew
flabel locali s 9982 11539 10016 11645 3 FreeSans 520 0 0 0 vgnd
port 2 nsew
flabel metal2 s -81 6117 -42 6227 0 FreeSans 200 0 0 0 ie_diff_sel_h_n
port 11 nsew
flabel metal2 s 15394 4945 15747 5041 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 12964 5158 13257 5253 0 FreeSans 400 180 0 0 vcc_io
port 5 nsew
flabel metal2 s 1471 6267 1523 6315 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 2939 2911 2939 2911 0 FreeSans 100 0 0 0 n2b
flabel metal2 s 1946 6267 1998 6315 3 FreeSans 400 90 0 0 pcasc
port 13 nsew
flabel metal2 s 11477 5411 11797 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 321 1255 640 1306 0 FreeSans 200 180 0 0 vpwr
port 4 nsew
flabel metal2 s 878 6267 930 6315 3 FreeSans 400 90 0 0 out_h
port 14 nsew
flabel metal2 s 1124 6267 1443 6315 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 321 6267 821 6315 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 11120 5411 11318 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 10483 5411 10879 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 9366 5411 10024 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 8181 5411 9138 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 7387 5411 8070 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 6963 5411 7331 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 6136 5411 6708 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 5338 5411 6028 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 3750 5443 4070 5505 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 13873 5409 14001 5505 0 FreeSans 400 180 0 0 pad_esd
port 16 nsew
flabel metal2 s 2374 5457 2694 5505 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 2750 6260 2802 6298 7 FreeSans 200 90 0 0 ie_diff_sel_h
port 9 nsew
flabel metal2 s 12991 6266 13344 6362 0 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal2 s 16182 7126 16474 7936 0 FreeSans 200 0 0 0 vpwr
port 4 nsew
flabel metal2 s 4418 5411 4717 5506 0 FreeSans 400 180 0 0 vcc_io
port 5 nsew
flabel metal2 s 2026 5457 2346 5505 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
flabel metal2 s 14045 10446 14365 10494 0 FreeSans 400 180 0 0 vcc_ioq
port 15 nsew
<< properties >>
string GDS_END 87458466
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86923478
string path 58.650 125.725 50.650 125.725 
<< end >>
