magic
tech sky130B
timestamp 1701704242
<< metal1 >>
rect 0 0 3 186
rect 157 0 160 186
<< via1 >>
rect 3 0 157 186
<< metal2 >>
rect 0 0 3 186
rect 157 0 160 186
<< properties >>
string GDS_END 85776914
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85774862
<< end >>
