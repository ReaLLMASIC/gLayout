magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< locali >>
rect 191 470 199 504
rect 233 470 271 504
rect 305 470 343 504
rect 377 470 415 504
rect 449 470 487 504
rect 521 470 529 504
rect 191 30 199 64
rect 233 30 271 64
rect 305 30 343 64
rect 377 30 415 64
rect 449 30 487 64
rect 521 30 529 64
<< viali >>
rect 199 470 233 504
rect 271 470 305 504
rect 343 470 377 504
rect 415 470 449 504
rect 487 470 521 504
rect 199 30 233 64
rect 271 30 305 64
rect 343 30 377 64
rect 415 30 449 64
rect 487 30 521 64
<< obsli1 >>
rect 48 392 82 402
rect 48 320 82 358
rect 48 248 82 286
rect 48 176 82 214
rect 48 132 82 142
rect 159 98 193 436
rect 251 98 285 436
rect 343 98 377 436
rect 435 98 469 436
rect 527 98 561 436
rect 638 392 672 402
rect 638 320 672 358
rect 638 248 672 286
rect 638 176 672 214
rect 638 132 672 142
<< obsli1c >>
rect 48 358 82 392
rect 48 286 82 320
rect 48 214 82 248
rect 48 142 82 176
rect 638 358 672 392
rect 638 286 672 320
rect 638 214 672 248
rect 638 142 672 176
<< metal1 >>
rect 187 504 533 524
rect 187 470 199 504
rect 233 470 271 504
rect 305 470 343 504
rect 377 470 415 504
rect 449 470 487 504
rect 521 470 533 504
rect 187 458 533 470
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 626 392 684 420
rect 626 358 638 392
rect 672 358 684 392
rect 626 320 684 358
rect 626 286 638 320
rect 672 286 684 320
rect 626 248 684 286
rect 626 214 638 248
rect 672 214 684 248
rect 626 176 684 214
rect 626 142 638 176
rect 672 142 684 176
rect 626 114 684 142
rect 187 64 533 76
rect 187 30 199 64
rect 233 30 271 64
rect 305 30 343 64
rect 377 30 415 64
rect 449 30 487 64
rect 521 30 533 64
rect 187 10 533 30
<< obsm1 >>
rect 150 114 202 420
rect 242 114 294 420
rect 334 114 386 420
rect 426 114 478 420
rect 518 114 570 420
<< metal2 >>
rect 10 292 710 420
rect 10 114 710 242
<< labels >>
rlabel metal2 s 10 292 710 420 6 DRAIN
port 1 nsew
rlabel viali s 487 470 521 504 6 GATE
port 2 nsew
rlabel viali s 487 30 521 64 6 GATE
port 2 nsew
rlabel viali s 415 470 449 504 6 GATE
port 2 nsew
rlabel viali s 415 30 449 64 6 GATE
port 2 nsew
rlabel viali s 343 470 377 504 6 GATE
port 2 nsew
rlabel viali s 343 30 377 64 6 GATE
port 2 nsew
rlabel viali s 271 470 305 504 6 GATE
port 2 nsew
rlabel viali s 271 30 305 64 6 GATE
port 2 nsew
rlabel viali s 199 470 233 504 6 GATE
port 2 nsew
rlabel viali s 199 30 233 64 6 GATE
port 2 nsew
rlabel locali s 191 470 529 504 6 GATE
port 2 nsew
rlabel locali s 191 30 529 64 6 GATE
port 2 nsew
rlabel metal1 s 187 458 533 524 6 GATE
port 2 nsew
rlabel metal1 s 187 10 533 76 6 GATE
port 2 nsew
rlabel metal2 s 10 114 710 242 6 SOURCE
port 3 nsew
rlabel metal1 s 36 114 94 420 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 626 114 684 420 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 10 10 710 524
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4984682
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4974286
<< end >>
