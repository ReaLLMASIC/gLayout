magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 978 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 614 47 644 177
rect 698 47 728 177
rect 782 47 812 177
rect 866 47 896 177
<< scpmoshvt >>
rect 79 297 109 497
rect 267 309 297 497
rect 351 309 381 497
rect 435 309 465 497
rect 519 309 549 497
rect 614 297 644 497
rect 698 297 728 497
rect 782 297 812 497
rect 866 297 896 497
<< ndiff >>
rect 27 106 79 177
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 163 177
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 124 251 177
rect 193 90 207 124
rect 241 90 251 124
rect 193 47 251 90
rect 281 89 335 177
rect 281 55 291 89
rect 325 55 335 89
rect 281 47 335 55
rect 365 124 419 177
rect 365 90 375 124
rect 409 90 419 124
rect 365 47 419 90
rect 449 89 505 177
rect 449 55 459 89
rect 493 55 505 89
rect 449 47 505 55
rect 562 124 614 177
rect 562 90 570 124
rect 604 90 614 124
rect 562 47 614 90
rect 644 169 698 177
rect 644 135 654 169
rect 688 135 698 169
rect 644 47 698 135
rect 728 89 782 177
rect 728 55 738 89
rect 772 55 782 89
rect 728 47 782 55
rect 812 169 866 177
rect 812 135 822 169
rect 856 135 866 169
rect 812 47 866 135
rect 896 89 952 177
rect 896 55 906 89
rect 940 55 952 89
rect 896 47 952 55
<< pdiff >>
rect 27 450 79 497
rect 27 416 35 450
rect 69 416 79 450
rect 27 297 79 416
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 297 161 451
rect 215 465 267 497
rect 215 431 223 465
rect 257 431 267 465
rect 215 309 267 431
rect 297 489 351 497
rect 297 455 307 489
rect 341 455 351 489
rect 297 421 351 455
rect 297 387 307 421
rect 341 387 351 421
rect 297 309 351 387
rect 381 477 435 497
rect 381 443 391 477
rect 425 443 435 477
rect 381 409 435 443
rect 381 375 391 409
rect 425 375 435 409
rect 381 309 435 375
rect 465 489 519 497
rect 465 455 475 489
rect 509 455 519 489
rect 465 421 519 455
rect 465 387 475 421
rect 509 387 519 421
rect 465 309 519 387
rect 549 477 614 497
rect 549 443 565 477
rect 599 443 614 477
rect 549 409 614 443
rect 549 375 565 409
rect 599 375 614 409
rect 549 309 614 375
rect 564 297 614 309
rect 644 407 698 497
rect 644 373 654 407
rect 688 373 698 407
rect 644 339 698 373
rect 644 305 654 339
rect 688 305 698 339
rect 644 297 698 305
rect 728 477 782 497
rect 728 443 738 477
rect 772 443 782 477
rect 728 409 782 443
rect 728 375 738 409
rect 772 375 782 409
rect 728 297 782 375
rect 812 407 866 497
rect 812 373 822 407
rect 856 373 866 407
rect 812 339 866 373
rect 812 305 822 339
rect 856 305 866 339
rect 812 297 866 305
rect 896 477 948 497
rect 896 443 906 477
rect 940 443 948 477
rect 896 409 948 443
rect 896 375 906 409
rect 940 375 948 409
rect 896 297 948 375
<< ndiffc >>
rect 35 72 69 106
rect 119 55 153 89
rect 207 90 241 124
rect 291 55 325 89
rect 375 90 409 124
rect 459 55 493 89
rect 570 90 604 124
rect 654 135 688 169
rect 738 55 772 89
rect 822 135 856 169
rect 906 55 940 89
<< pdiffc >>
rect 35 416 69 450
rect 119 451 153 485
rect 223 431 257 465
rect 307 455 341 489
rect 307 387 341 421
rect 391 443 425 477
rect 391 375 425 409
rect 475 455 509 489
rect 475 387 509 421
rect 565 443 599 477
rect 565 375 599 409
rect 654 373 688 407
rect 654 305 688 339
rect 738 443 772 477
rect 738 375 772 409
rect 822 373 856 407
rect 822 305 856 339
rect 906 443 940 477
rect 906 375 940 409
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 614 497 644 523
rect 698 497 728 523
rect 782 497 812 523
rect 866 497 896 523
rect 79 265 109 297
rect 21 249 109 265
rect 267 294 297 309
rect 351 294 381 309
rect 435 294 465 309
rect 519 294 549 309
rect 267 264 549 294
rect 21 215 32 249
rect 66 222 109 249
rect 495 249 549 264
rect 66 215 449 222
rect 21 199 449 215
rect 495 215 505 249
rect 539 215 549 249
rect 495 199 549 215
rect 614 265 644 297
rect 698 265 728 297
rect 614 259 728 265
rect 782 259 812 297
rect 866 261 896 297
rect 866 259 950 261
rect 614 249 950 259
rect 614 215 764 249
rect 798 215 832 249
rect 866 215 900 249
rect 934 215 950 249
rect 614 205 950 215
rect 614 199 728 205
rect 79 192 449 199
rect 79 177 109 192
rect 163 177 193 192
rect 251 177 281 192
rect 335 177 365 192
rect 419 177 449 192
rect 614 177 644 199
rect 698 177 728 199
rect 782 177 812 205
rect 866 203 950 205
rect 866 177 896 203
rect 79 21 109 47
rect 163 21 193 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 614 21 644 47
rect 698 21 728 47
rect 782 21 812 47
rect 866 21 896 47
<< polycont >>
rect 32 215 66 249
rect 505 215 539 249
rect 764 215 798 249
rect 832 215 866 249
rect 900 215 934 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 450 69 493
rect 17 416 35 450
rect 103 485 175 527
rect 103 451 119 485
rect 153 451 175 485
rect 103 425 175 451
rect 215 465 257 493
rect 215 431 223 465
rect 17 391 69 416
rect 17 357 175 391
rect 17 249 66 323
rect 17 215 32 249
rect 17 199 66 215
rect 100 265 175 357
rect 215 345 257 431
rect 291 489 357 527
rect 291 455 307 489
rect 341 455 357 489
rect 291 421 357 455
rect 291 387 307 421
rect 341 387 357 421
rect 291 379 357 387
rect 391 477 425 493
rect 391 409 425 443
rect 459 489 531 527
rect 459 455 475 489
rect 509 455 531 489
rect 459 421 531 455
rect 459 387 475 421
rect 509 387 531 421
rect 459 379 531 387
rect 565 477 995 493
rect 599 459 738 477
rect 565 409 599 443
rect 772 459 906 477
rect 391 345 425 375
rect 565 345 599 375
rect 215 311 599 345
rect 638 407 704 425
rect 638 373 654 407
rect 688 373 704 407
rect 638 339 704 373
rect 738 409 772 443
rect 940 443 995 477
rect 738 357 772 375
rect 806 407 872 425
rect 806 373 822 407
rect 856 373 872 407
rect 638 305 654 339
rect 688 323 704 339
rect 806 339 872 373
rect 806 323 822 339
rect 688 305 822 323
rect 856 305 872 339
rect 638 289 872 305
rect 906 409 995 443
rect 940 375 995 409
rect 906 289 995 375
rect 100 249 604 265
rect 100 215 505 249
rect 539 215 604 249
rect 100 199 604 215
rect 100 165 139 199
rect 638 170 714 289
rect 748 249 995 255
rect 748 215 764 249
rect 798 215 832 249
rect 866 215 900 249
rect 934 215 995 249
rect 748 204 995 215
rect 638 169 995 170
rect 17 131 139 165
rect 207 131 604 165
rect 17 106 69 131
rect 17 72 35 106
rect 207 124 241 131
rect 17 51 69 72
rect 103 89 169 97
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 375 124 409 131
rect 207 51 241 90
rect 275 89 341 97
rect 275 55 291 89
rect 325 55 341 89
rect 275 17 341 55
rect 547 124 604 131
rect 638 135 654 169
rect 688 135 822 169
rect 856 135 995 169
rect 638 127 995 135
rect 375 51 409 90
rect 443 89 511 97
rect 443 55 459 89
rect 493 55 511 89
rect 443 17 511 55
rect 547 90 570 124
rect 604 90 995 93
rect 547 89 995 90
rect 547 55 738 89
rect 772 55 906 89
rect 940 55 995 89
rect 547 51 995 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 TE
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 TE
port 2 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 770 289 804 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 678 289 712 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 678 153 712 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 678 221 712 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 einvp_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 2038900
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2030936
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 25.300 13.600 
<< end >>
