magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect 811 1782 831 2514
rect 4464 1464 4504 2596
<< poly >>
rect 322 1472 463 1536
rect 322 1438 338 1472
rect 372 1438 406 1472
rect 440 1438 463 1472
rect 322 1405 463 1438
rect 526 1475 639 1536
rect 526 1455 660 1475
rect 526 1421 542 1455
rect 576 1421 610 1455
rect 644 1421 660 1455
rect 526 1405 660 1421
rect 704 1472 838 1536
rect 704 1438 720 1472
rect 754 1438 788 1472
rect 822 1438 838 1472
rect 704 1405 838 1438
rect 5059 1386 5113 1462
rect 4857 1012 5313 1034
rect 4857 978 4893 1012
rect 4927 978 4961 1012
rect 4995 978 5029 1012
rect 5063 978 5097 1012
rect 5131 978 5165 1012
rect 5199 978 5233 1012
rect 5267 978 5313 1012
rect 4857 958 5313 978
rect 5059 530 5113 606
<< polycont >>
rect 338 1438 372 1472
rect 406 1438 440 1472
rect 542 1421 576 1455
rect 610 1421 644 1455
rect 720 1438 754 1472
rect 788 1438 822 1472
rect 4893 978 4927 1012
rect 4961 978 4995 1012
rect 5029 978 5063 1012
rect 5097 978 5131 1012
rect 5165 978 5199 1012
rect 5233 978 5267 1012
<< locali >>
rect 542 2100 564 2134
rect 598 2100 616 2134
rect 542 2062 616 2100
rect 542 2028 564 2062
rect 598 2028 616 2062
rect 298 1688 332 1726
rect 298 1616 332 1654
rect 368 1502 406 1536
rect 334 1472 440 1502
rect 334 1438 338 1472
rect 372 1438 406 1472
rect 334 1422 440 1438
rect 474 1386 508 1624
rect 542 1471 616 2028
rect 856 1988 890 2166
rect 860 1954 890 1988
rect 1121 1954 1159 1988
rect 826 1916 890 1954
rect 860 1882 890 1916
rect 650 1688 684 1726
rect 650 1616 684 1654
rect 720 1472 822 1488
rect 542 1455 644 1471
rect 576 1421 610 1455
rect 754 1438 788 1472
rect 720 1422 822 1438
rect 542 1405 644 1421
rect 318 1352 474 1383
rect 318 1314 508 1352
rect 318 1280 474 1314
rect 738 1386 812 1422
rect 738 1352 750 1386
rect 784 1352 812 1386
rect 738 1314 812 1352
rect 738 1280 750 1314
rect 784 1280 812 1314
rect 670 1162 704 1200
rect 856 1181 890 1882
rect 4869 1432 5034 1433
rect 5059 1432 5113 1442
rect 4869 1398 4895 1432
rect 4929 1398 4967 1432
rect 5001 1398 5039 1432
rect 5073 1398 5111 1432
rect 5145 1398 5183 1432
rect 5217 1398 5255 1432
rect 5289 1398 5315 1408
rect 4869 1342 5034 1398
rect 4869 1308 4901 1342
rect 4935 1308 4973 1342
rect 5007 1308 5034 1342
rect 670 1090 704 1128
rect 4869 1012 5034 1308
rect 5136 1342 5315 1398
rect 5136 1308 5167 1342
rect 5201 1308 5239 1342
rect 5273 1308 5315 1342
rect 6311 1357 6417 1408
rect 6345 1323 6383 1357
rect 6567 1357 6673 1408
rect 6601 1323 6639 1357
rect 5136 1012 5315 1308
rect 4869 978 4893 1012
rect 4927 978 4961 1012
rect 4995 978 5029 1012
rect 5063 978 5097 1012
rect 5131 978 5165 1012
rect 5199 978 5233 1012
rect 5267 978 5315 1012
rect 4869 924 5034 978
rect 4869 890 4895 924
rect 4929 890 4967 924
rect 5001 890 5034 924
rect 4869 584 5034 890
rect 5136 924 5315 978
rect 5136 890 5169 924
rect 5203 890 5241 924
rect 5275 890 5315 924
rect 5136 584 5315 890
rect 5059 550 5113 584
rect 6311 527 6349 561
rect 6567 527 6605 561
rect 3184 305 3222 339
<< viali >>
rect 564 2100 598 2134
rect 564 2028 598 2062
rect 298 1726 332 1760
rect 298 1654 332 1688
rect 298 1582 332 1616
rect 334 1502 368 1536
rect 406 1502 440 1536
rect 826 1954 860 1988
rect 1087 1954 1121 1988
rect 1159 1954 1193 1988
rect 826 1882 860 1916
rect 650 1726 684 1760
rect 650 1654 684 1688
rect 650 1582 684 1616
rect 474 1352 508 1386
rect 474 1280 508 1314
rect 750 1352 784 1386
rect 750 1280 784 1314
rect 670 1200 704 1234
rect 4895 1398 4929 1432
rect 4967 1398 5001 1432
rect 5039 1398 5073 1432
rect 5111 1398 5145 1432
rect 5183 1398 5217 1432
rect 5255 1398 5289 1432
rect 4901 1308 4935 1342
rect 4973 1308 5007 1342
rect 670 1128 704 1162
rect 670 1056 704 1090
rect 5167 1308 5201 1342
rect 5239 1308 5273 1342
rect 6311 1323 6345 1357
rect 6383 1323 6417 1357
rect 6567 1323 6601 1357
rect 6639 1323 6673 1357
rect 4895 890 4929 924
rect 4967 890 5001 924
rect 5169 890 5203 924
rect 5241 890 5275 924
rect 6277 527 6311 561
rect 6349 527 6383 561
rect 6533 527 6567 561
rect 6605 527 6639 561
rect 3150 305 3184 339
rect 3222 305 3256 339
<< metal1 >>
rect -66 2284 7072 2430
rect 4464 2250 7072 2256
rect 4464 2228 4715 2250
tri 4690 2203 4715 2228 ne
rect 4464 2172 4562 2200
tri 4562 2172 4590 2200 sw
rect 4767 2228 6809 2250
tri 4767 2203 4792 2228 nw
tri 6784 2203 6809 2228 ne
rect 4715 2186 4767 2198
tri 4550 2140 4582 2172 ne
rect 4582 2140 4590 2172
rect 552 2134 610 2140
rect 552 2100 564 2134
rect 598 2100 610 2134
tri 4582 2132 4590 2140 ne
tri 4590 2132 4630 2172 sw
tri 4590 2128 4594 2132 ne
rect 4594 2128 4630 2132
tri 4630 2128 4634 2132 sw
rect 4715 2128 4767 2134
rect 5437 2194 5489 2200
rect 5437 2130 5489 2142
tri 4594 2105 4617 2128 ne
rect 4617 2105 4634 2128
tri 527 2068 552 2093 se
rect 552 2068 610 2100
tri 610 2068 635 2093 sw
tri 1295 2068 1320 2093 se
rect 1320 2068 1366 2105
tri 4617 2092 4630 2105 ne
rect 4630 2100 4634 2105
tri 4634 2100 4662 2128 sw
tri 5412 2100 5437 2125 se
rect 4630 2092 5437 2100
tri 4630 2072 4650 2092 ne
rect 4650 2078 5437 2092
rect 6087 2194 6139 2200
rect 6087 2130 6139 2142
tri 5489 2100 5514 2125 sw
tri 6062 2100 6087 2125 se
rect 5489 2078 6087 2100
rect 6861 2228 7072 2250
tri 6861 2203 6886 2228 nw
rect 6809 2186 6861 2198
rect 6809 2128 6861 2134
tri 6139 2100 6164 2125 sw
rect 6139 2078 7072 2100
rect 4650 2072 7072 2078
rect 0 2062 1366 2068
rect 0 2028 564 2062
rect 598 2028 1366 2062
rect 0 2022 1366 2028
rect 691 1988 1205 1994
rect 743 1954 826 1988
rect 860 1954 1087 1988
rect 1121 1954 1159 1988
rect 1193 1954 1205 1988
rect 743 1948 1205 1954
rect 743 1936 878 1948
rect 691 1924 878 1936
rect 743 1916 878 1924
tri 878 1923 903 1948 nw
rect 743 1882 826 1916
rect 860 1882 878 1916
rect 743 1872 878 1882
rect 691 1866 878 1872
rect 4464 1800 4560 1846
rect 5700 1800 5740 1846
rect 5836 1800 5877 1846
rect 7016 1800 7072 1846
rect -66 1760 7072 1772
rect -66 1726 298 1760
rect 332 1726 650 1760
rect 684 1726 7072 1760
rect -66 1688 7072 1726
rect -66 1654 298 1688
rect 332 1654 650 1688
rect 684 1654 7072 1688
rect -66 1616 7072 1654
rect -66 1582 298 1616
rect 332 1582 650 1616
rect 684 1606 7072 1616
rect 684 1582 1445 1606
rect -66 1570 1445 1582
tri 1445 1570 1481 1606 nw
tri 1595 1570 1631 1606 ne
rect 1631 1570 7072 1606
rect 0 1536 452 1542
rect 0 1502 334 1536
rect 368 1502 406 1536
rect 440 1502 452 1536
rect 0 1496 452 1502
tri 4467 1468 4492 1493 se
rect 4492 1490 4569 1542
rect 4571 1541 4607 1542
rect 4570 1491 4608 1541
rect 4609 1514 5301 1542
rect 4571 1490 4607 1491
rect 4609 1490 4687 1514
rect 4492 1468 4544 1490
rect 4464 1416 4544 1468
tri 4544 1465 4569 1490 nw
tri 4610 1465 4635 1490 ne
rect 4635 1465 4687 1490
tri 4687 1489 4712 1514 nw
tri 4858 1489 4883 1514 ne
rect 4636 1463 4686 1464
rect 4883 1432 5301 1514
tri 4467 1398 4485 1416 ne
rect 4485 1402 4544 1416
tri 4544 1402 4569 1427 sw
rect 4636 1426 4686 1427
rect 4485 1398 4607 1402
tri 4485 1392 4491 1398 ne
rect 4491 1396 4607 1398
rect 4491 1392 4555 1396
rect 462 1386 525 1392
rect 462 1352 474 1386
rect 508 1352 525 1386
rect 462 1340 525 1352
rect 577 1386 796 1392
tri 4491 1391 4492 1392 ne
rect 577 1352 750 1386
rect 784 1352 796 1386
rect 577 1340 796 1352
rect 462 1328 796 1340
rect 462 1314 525 1328
rect 462 1280 474 1314
rect 508 1280 525 1314
rect 462 1276 525 1280
rect 577 1314 796 1328
rect 577 1280 750 1314
rect 784 1280 796 1314
rect 577 1276 796 1280
rect 462 1274 796 1276
rect 4492 1344 4555 1392
rect 4492 1332 4607 1344
rect 4492 1280 4555 1332
rect 4492 1274 4607 1280
rect 4635 1396 4687 1425
rect 4635 1332 4687 1344
rect 4635 1274 4687 1280
rect 4883 1398 4895 1432
rect 4929 1398 4967 1432
rect 5001 1398 5039 1432
rect 5073 1398 5111 1432
rect 5145 1398 5183 1432
rect 5217 1398 5255 1432
rect 5289 1398 5301 1432
rect 4883 1342 5301 1398
rect 5786 1475 6685 1481
rect 5838 1429 6685 1475
rect 5786 1411 5838 1423
tri 5838 1404 5863 1429 nw
tri 6274 1404 6299 1429 ne
rect 6299 1404 6429 1429
tri 6429 1404 6454 1429 nw
tri 6530 1404 6555 1429 ne
rect 6555 1404 6685 1429
rect 5786 1353 5838 1359
rect 6300 1402 6428 1403
rect 6299 1366 6429 1402
rect 6300 1365 6428 1366
rect 6299 1357 6429 1364
rect 4883 1308 4901 1342
rect 4935 1308 4973 1342
rect 5007 1308 5167 1342
rect 5201 1308 5239 1342
rect 5273 1308 5301 1342
rect 6299 1323 6311 1357
rect 6345 1323 6383 1357
rect 6417 1323 6429 1357
rect 6299 1311 6429 1323
rect 6300 1309 6428 1310
rect 6556 1402 6684 1403
rect 6555 1366 6685 1402
rect 6556 1365 6684 1366
rect 6555 1357 6685 1364
rect 6555 1323 6567 1357
rect 6601 1323 6639 1357
rect 6673 1323 6685 1357
rect 6555 1311 6685 1323
rect 6556 1309 6684 1310
rect 4883 1274 5301 1308
rect 6300 1272 6428 1273
rect 6556 1272 6684 1273
tri 6274 1246 6299 1271 se
rect 6299 1246 6429 1271
tri 6429 1246 6454 1271 sw
tri 6530 1246 6555 1271 se
rect 6555 1246 6685 1271
tri 6685 1246 6710 1271 sw
rect -66 1234 7006 1246
rect -66 1200 670 1234
rect 704 1200 7006 1234
rect -66 1162 7006 1200
rect -66 1128 670 1162
rect 704 1128 7006 1162
rect -66 1090 7006 1128
rect -66 1056 670 1090
rect 704 1056 7006 1090
rect -66 1044 7006 1056
rect 7036 1044 7072 1246
rect 4889 924 5007 936
rect 4889 890 4895 924
rect 4929 890 4967 924
rect 5001 890 5007 924
rect 4889 878 5007 890
rect 5163 924 5281 936
rect 5163 890 5169 924
rect 5203 890 5241 924
rect 5275 890 5281 924
rect 5163 878 5281 890
rect -66 632 7072 762
tri 6240 607 6265 632 ne
rect 6265 607 6395 632
tri 6395 607 6420 632 nw
rect 6266 605 6394 606
rect 5786 598 5838 604
tri 5774 573 5786 585 se
rect 691 567 743 573
tri 5762 561 5774 573 se
rect 5774 561 5786 573
tri 5761 560 5762 561 se
rect 5762 560 5786 561
tri 4526 527 4559 560 se
rect 4559 554 5721 560
rect 4559 527 4635 554
tri 4515 516 4526 527 se
rect 4526 516 4635 527
rect 691 503 743 515
tri 494 417 519 442 se
rect 519 435 525 487
rect 577 435 583 487
tri 743 491 768 516 sw
tri 4490 491 4515 516 se
rect 4515 502 4635 516
rect 4687 508 5721 554
rect 5722 509 5723 559
rect 5759 509 5760 559
rect 5761 546 5786 560
rect 6266 568 6394 569
rect 6265 561 6395 567
rect 5761 534 5838 546
rect 5761 508 5786 534
rect 4515 491 4687 502
rect 743 490 4687 491
rect 743 451 4635 490
rect 691 445 4635 451
tri 4622 442 4625 445 ne
rect 4625 442 4635 445
rect 519 432 583 435
tri 583 432 593 442 sw
tri 4625 432 4635 442 ne
tri 4687 483 4712 508 nw
tri 5761 483 5786 508 ne
rect 4635 432 4687 438
tri 5838 527 5860 549 sw
rect 6265 527 6277 561
rect 6311 527 6349 561
rect 6383 527 6395 561
rect 5838 524 5860 527
tri 5860 524 5863 527 sw
rect 5838 508 5987 524
tri 5987 508 6003 524 sw
rect 6265 515 6395 527
rect 6266 513 6394 514
rect 5838 484 6003 508
tri 6003 484 6027 508 sw
rect 5786 459 5838 482
tri 5838 459 5863 484 nw
tri 5969 459 5994 484 ne
rect 5994 475 6027 484
tri 6027 475 6036 484 sw
rect 6265 477 6395 513
rect 6266 476 6394 477
rect 6521 561 6653 567
rect 6521 527 6533 561
rect 6567 527 6605 561
rect 6639 527 6653 561
rect 5994 459 6036 475
tri 6036 459 6052 475 sw
tri 6249 459 6265 475 se
rect 6265 459 6395 475
tri 5994 458 5995 459 ne
rect 5995 458 6052 459
rect 5787 457 5837 458
tri 5995 457 5996 458 ne
rect 5996 457 6052 458
rect 519 423 593 432
rect 519 417 525 423
rect 462 371 525 417
rect 577 417 593 423
tri 593 417 608 432 sw
tri 5335 417 5350 432 se
rect 5350 419 5603 432
tri 5603 419 5616 432 sw
rect 5786 421 5838 457
tri 5996 450 6003 457 ne
rect 6003 450 6052 457
tri 6052 450 6061 459 sw
tri 6240 450 6249 459 se
rect 6249 450 6395 459
tri 6395 450 6420 475 sw
tri 6496 450 6521 475 se
rect 6521 450 6653 527
tri 6003 423 6030 450 ne
rect 6030 423 6653 450
tri 6030 421 6032 423 ne
rect 6032 421 6653 423
rect 5787 420 5837 421
tri 6032 420 6033 421 ne
rect 6033 420 6653 421
tri 6033 419 6034 420 ne
rect 6034 419 6653 420
rect 5350 417 5616 419
tri 5616 417 5618 419 sw
tri 5784 417 5786 419 se
rect 5786 417 5838 419
rect 577 371 3268 417
tri 3113 346 3138 371 ne
rect 3138 339 3268 371
rect 3138 305 3150 339
rect 3184 305 3222 339
rect 3256 305 3268 339
rect 3138 299 3268 305
rect 4555 411 4607 417
tri 5312 394 5335 417 se
rect 5335 394 5618 417
tri 5618 394 5641 417 sw
tri 5761 394 5784 417 se
rect 5784 394 5838 417
tri 6034 409 6044 419 ne
rect 6044 409 6653 419
tri 5285 367 5312 394 se
rect 5312 380 5838 394
rect 5312 367 5359 380
tri 5359 367 5372 380 nw
tri 5581 367 5594 380 ne
rect 5594 367 5838 380
tri 5284 366 5285 367 se
rect 5285 366 5350 367
rect 4555 347 4607 359
tri 4607 341 4632 366 sw
tri 5276 358 5284 366 se
rect 5284 358 5350 366
tri 5350 358 5359 367 nw
tri 5594 358 5603 367 ne
rect 5603 358 5838 367
tri 5259 341 5276 358 se
rect 5276 341 5333 358
tri 5333 341 5350 358 nw
tri 5603 342 5619 358 ne
rect 5619 342 5838 358
rect 4607 295 5281 341
rect 4555 289 5281 295
tri 5281 289 5333 341 nw
<< rmetal1 >>
rect 4569 1541 4571 1542
rect 4607 1541 4609 1542
rect 4569 1491 4570 1541
rect 4608 1491 4609 1541
rect 4569 1490 4571 1491
rect 4607 1490 4609 1491
rect 4635 1464 4687 1465
rect 4635 1463 4636 1464
rect 4686 1463 4687 1464
rect 4635 1426 4636 1427
rect 4686 1426 4687 1427
rect 4635 1425 4687 1426
rect 6299 1403 6429 1404
rect 6299 1402 6300 1403
rect 6428 1402 6429 1403
rect 6299 1365 6300 1366
rect 6428 1365 6429 1366
rect 6299 1364 6429 1365
rect 6299 1310 6429 1311
rect 6299 1309 6300 1310
rect 6428 1309 6429 1310
rect 6555 1403 6685 1404
rect 6555 1402 6556 1403
rect 6684 1402 6685 1403
rect 6555 1365 6556 1366
rect 6684 1365 6685 1366
rect 6555 1364 6685 1365
rect 6555 1310 6685 1311
rect 6555 1309 6556 1310
rect 6684 1309 6685 1310
rect 6299 1272 6300 1273
rect 6428 1272 6429 1273
rect 6299 1271 6429 1272
rect 6555 1272 6556 1273
rect 6684 1272 6685 1273
rect 6555 1271 6685 1272
rect 6265 606 6395 607
rect 6265 605 6266 606
rect 6394 605 6395 606
rect 5721 559 5723 560
rect 5721 509 5722 559
rect 5721 508 5723 509
rect 5759 559 5761 560
rect 5760 509 5761 559
rect 6265 568 6266 569
rect 6394 568 6395 569
rect 6265 567 6395 568
rect 5759 508 5761 509
rect 6265 514 6395 515
rect 6265 513 6266 514
rect 6394 513 6395 514
rect 6265 476 6266 477
rect 6394 476 6395 477
rect 6265 475 6395 476
rect 5786 458 5838 459
rect 5786 457 5787 458
rect 5837 457 5838 458
rect 5786 420 5787 421
rect 5837 420 5838 421
rect 5786 419 5838 420
<< via1 >>
rect 4715 2198 4767 2250
rect 4715 2134 4767 2186
rect 5437 2142 5489 2194
rect 5437 2078 5489 2130
rect 6087 2142 6139 2194
rect 6087 2078 6139 2130
rect 6809 2198 6861 2250
rect 6809 2134 6861 2186
rect 691 1936 743 1988
rect 691 1872 743 1924
rect 525 1340 577 1392
rect 525 1276 577 1328
rect 4555 1344 4607 1396
rect 4555 1280 4607 1332
rect 4635 1344 4687 1396
rect 4635 1280 4687 1332
rect 5786 1423 5838 1475
rect 5786 1359 5838 1411
rect 691 515 743 567
rect 525 435 577 487
rect 691 451 743 503
rect 4635 502 4687 554
rect 5786 546 5838 598
rect 4635 438 4687 490
rect 5786 482 5838 534
rect 525 371 577 423
rect 4555 359 4607 411
rect 4555 295 4607 347
<< metal2 >>
rect 4715 2250 4767 2256
rect 6809 2250 6861 2256
rect 4715 2186 4767 2198
rect 4715 2128 4767 2134
rect 5437 2194 5489 2200
rect 5437 2130 5489 2142
rect 5437 2072 5489 2078
rect 6087 2194 6139 2200
rect 6087 2130 6139 2142
rect 6809 2186 6861 2198
rect 6809 2128 6861 2134
rect 6087 2072 6139 2078
rect 691 1988 743 1994
rect 691 1924 743 1936
rect 519 1340 525 1392
rect 577 1340 583 1392
rect 519 1328 583 1340
rect 519 1276 525 1328
rect 577 1276 583 1328
rect 519 487 583 1276
rect 519 435 525 487
rect 577 435 583 487
rect 691 567 743 1872
rect 5786 1475 5838 1481
rect 5786 1411 5838 1423
rect 691 503 743 515
rect 691 445 743 451
rect 4555 1396 4607 1402
rect 4555 1332 4607 1344
rect 519 423 583 435
rect 519 371 525 423
rect 577 371 583 423
rect 4555 411 4607 1280
rect 4635 1396 4687 1402
rect 4635 1332 4687 1344
rect 4635 554 4687 1280
rect 4635 490 4687 502
rect 5786 598 5838 1359
rect 5786 534 5838 546
rect 5786 476 5838 482
rect 4635 432 4687 438
rect 4555 347 4607 359
rect 4555 289 4607 295
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_0
timestamp 1701704242
transform -1 0 659 0 -1 1379
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_1
timestamp 1701704242
transform 1 0 363 0 -1 1379
box -79 -26 196 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_0
timestamp 1701704242
transform 1 0 715 0 -1 1379
box -79 -26 199 226
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_0
timestamp 1701704242
transform 1 0 343 0 -1 2162
box -119 -66 415 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_0
timestamp 1701704242
transform 1 0 695 0 -1 2162
box -119 -66 239 666
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1701704242
transform -1 0 598 0 1 2028
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1701704242
transform -1 0 860 0 1 1882
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1701704242
transform -1 0 508 0 1 1280
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1701704242
transform -1 0 784 0 1 1280
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1701704242
transform 0 1 4895 1 0 890
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1701704242
transform 0 1 5169 1 0 890
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1701704242
transform 0 1 4901 1 0 1308
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1701704242
transform 0 1 5167 1 0 1308
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1701704242
transform -1 0 6417 0 1 1323
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1701704242
transform -1 0 6673 0 1 1323
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1701704242
transform -1 0 1193 0 1 1954
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1701704242
transform -1 0 3256 0 1 305
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1701704242
transform -1 0 440 0 -1 1536
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1701704242
transform 1 0 6277 0 1 527
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1701704242
transform 1 0 6533 0 1 527
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1701704242
transform 0 -1 684 -1 0 1760
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1701704242
transform 0 -1 704 -1 0 1234
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1701704242
transform 0 -1 332 -1 0 1760
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1701704242
transform 1 0 4895 0 1 1398
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1701704242
transform 0 -1 4607 -1 0 1402
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1701704242
transform 0 -1 5838 -1 0 604
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1701704242
transform 0 -1 4687 -1 0 1402
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1701704242
transform 0 1 691 -1 0 1994
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1701704242
transform 0 1 5786 -1 0 1481
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1701704242
transform 0 1 4555 1 0 289
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1701704242
transform 0 1 6809 1 0 2128
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1701704242
transform 0 1 5437 1 0 2072
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1701704242
transform 0 1 6087 1 0 2072
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1701704242
transform 0 1 4715 1 0 2128
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1701704242
transform 0 -1 743 1 0 445
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1701704242
transform 0 -1 4687 1 0 432
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1701704242
transform 1 0 519 0 -1 1392
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1701704242
transform 1 0 519 0 1 371
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1701704242
transform 1 0 526 0 -1 1471
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1701704242
transform 1 0 322 0 -1 1488
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1701704242
transform 1 0 704 0 1 1422
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1701704242
transform 0 1 4877 1 0 962
box 0 0 1 1
use sky130_fd_io__sio_com_pupredrvr_nbias  sky130_fd_io__sio_com_pupredrvr_nbias_0
timestamp 1701704242
transform 1 0 831 0 1 165
box 0 10 3633 2349
use sky130_fd_io__sio_com_pupredrvr_strong_nd2  sky130_fd_io__sio_com_pupredrvr_strong_nd2_0
timestamp 1701704242
transform -1 0 7072 0 1 0
box 0 10 1284 2632
use sky130_fd_io__sio_com_pupredrvr_strong_nd2  sky130_fd_io__sio_com_pupredrvr_strong_nd2_1
timestamp 1701704242
transform 1 0 4504 0 1 0
box 0 10 1284 2632
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_0
timestamp 1701704242
transform 0 -1 4687 1 0 1373
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_1
timestamp 1701704242
transform 1 0 5669 0 1 508
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851421  sky130_fd_io__sio_tk_em1o_CDNS_524688791851421_0
timestamp 1701704242
transform 0 -1 6685 1 0 1219
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851421  sky130_fd_io__sio_tk_em1o_CDNS_524688791851421_1
timestamp 1701704242
transform 0 -1 6429 1 0 1219
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851421  sky130_fd_io__sio_tk_em1o_CDNS_524688791851421_2
timestamp 1701704242
transform 0 -1 6395 1 0 515
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1701704242
transform 0 1 5786 -1 0 511
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1701704242
transform -1 0 4661 0 1 1490
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851418  sky130_fd_io__sio_tk_em1s_CDNS_524688791851418_0
timestamp 1701704242
transform 0 1 6265 -1 0 567
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851418  sky130_fd_io__sio_tk_em1s_CDNS_524688791851418_1
timestamp 1701704242
transform 0 -1 6685 1 0 1312
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851418  sky130_fd_io__sio_tk_em1s_CDNS_524688791851418_2
timestamp 1701704242
transform 0 -1 6429 1 0 1312
box 0 0 1 1
<< labels >>
flabel comment s 633 397 633 397 0 FreeSans 300 0 0 0 en_fast_h_n
flabel comment s 839 1978 839 1978 0 FreeSans 300 0 0 0 en_fast_h
flabel comment s 902 469 902 469 0 FreeSans 300 0 0 0 en_fast_h
flabel comment s 5108 521 5108 521 0 FreeSans 300 180 0 0 en_fast_h
flabel metal1 s 7036 2228 7072 2256 7 FreeSans 300 180 0 0 drvhi_h
port 6 nsew
flabel metal1 s 7036 2072 7072 2100 7 FreeSans 300 180 0 0 puen_h
port 5 nsew
flabel metal1 s 0 1496 37 1542 3 FreeSans 300 180 0 0 slow_h_n
port 7 nsew
flabel metal1 s 7036 2284 7072 2430 7 FreeSans 300 180 0 0 vcc_io
port 1 nsew
flabel metal1 s -66 1570 -24 1772 3 FreeSans 300 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 5700 1800 5740 1846 2 FreeSans 300 180 0 0 pu_h_n<2>
port 2 nsew
flabel metal1 s -66 2284 -29 2430 3 FreeSans 300 0 0 0 vcc_io
port 1 nsew
flabel metal1 s -66 1044 -24 1246 3 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel metal1 s -66 632 -24 762 3 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel metal1 s 7036 1570 7072 1772 7 FreeSans 300 180 0 0 vcc_io
port 1 nsew
flabel metal1 s 7036 1044 7072 1246 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 7036 632 7072 762 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 7036 1800 7072 1846 7 FreeSans 300 180 0 0 pu_h_n<3>
port 4 nsew
flabel metal1 s 4504 1800 4540 1846 1 FreeSans 300 0 0 0 pu_h_n<2>
port 2 nsew
flabel metal1 s 5836 1800 5877 1846 2 FreeSans 300 0 0 0 pu_h_n<3>
port 4 nsew
flabel metal1 s 0 2022 36 2068 3 FreeSans 300 180 0 0 puen_h
port 5 nsew
flabel metal1 s 7055 2242 7055 2242 7 FreeSans 300 180 0 0 drvhi_h
flabel metal1 s 7054 2086 7054 2086 7 FreeSans 300 180 0 0 puen_h
flabel metal1 s 19 1519 19 1519 3 FreeSans 300 180 0 0 slow_h_n
flabel metal1 s 6402 1342 6402 1342 3 FreeSans 400 0 0 0 en_fast_h_3<1>
flabel metal1 s 6659 1339 6659 1339 3 FreeSans 400 0 0 0 en_fast_h_3<0>
flabel metal1 s 999 1979 999 1979 3 FreeSans 400 0 0 0 en_fast_h
flabel metal1 s 6367 547 6367 547 3 FreeSans 400 0 0 0 en_fast_h_3<2>
flabel metal1 s 866 393 866 393 3 FreeSans 400 0 0 0 en_fast_h_n
flabel metal1 s 6618 558 6618 558 3 FreeSans 400 0 0 0 en_fast_h_3<3>
flabel metal1 s 4319 1449 4319 1449 3 FreeSans 400 0 0 0 nbias_out
<< properties >>
string GDS_END 87821206
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87808002
<< end >>
