magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect -1298 -1522 1448 7522
<< nwell >>
rect -898 6600 1048 7122
rect -898 6026 -500 6600
rect 650 6026 1048 6600
rect -898 -26 -526 6026
rect 676 -26 1048 6026
rect -898 -600 -500 -26
rect 650 -600 1048 -26
rect -898 -1122 1048 -600
<< pwell >>
rect -1606 7696 1756 7830
rect -1606 -1696 -1472 7696
rect -526 -26 -274 6026
tri -26 5996 4 6026 se
rect 4 5996 146 6026
tri 146 5996 176 6026 sw
rect -26 4 176 5996
tri -26 -26 4 4 ne
rect 4 -26 146 4
tri 146 -26 176 4 nw
rect 424 -26 676 6026
rect 1622 -1696 1756 7696
rect -1606 -1830 1756 -1696
<< mvpmos >>
rect -600 0 -500 6000
rect 650 0 750 6000
<< mvpdiff >>
rect -658 5971 -600 6000
rect -658 5937 -646 5971
rect -612 5937 -600 5971
rect -658 5903 -600 5937
rect -658 5869 -646 5903
rect -612 5869 -600 5903
rect -658 5835 -600 5869
rect -658 5801 -646 5835
rect -612 5801 -600 5835
rect -658 5767 -600 5801
rect -658 5733 -646 5767
rect -612 5733 -600 5767
rect -658 5699 -600 5733
rect -658 5665 -646 5699
rect -612 5665 -600 5699
rect -658 5631 -600 5665
rect -658 5597 -646 5631
rect -612 5597 -600 5631
rect -658 5563 -600 5597
rect -658 5529 -646 5563
rect -612 5529 -600 5563
rect -658 5495 -600 5529
rect -658 5461 -646 5495
rect -612 5461 -600 5495
rect -658 5427 -600 5461
rect -658 5393 -646 5427
rect -612 5393 -600 5427
rect -658 5359 -600 5393
rect -658 5325 -646 5359
rect -612 5325 -600 5359
rect -658 5291 -600 5325
rect -658 5257 -646 5291
rect -612 5257 -600 5291
rect -658 5223 -600 5257
rect -658 5189 -646 5223
rect -612 5189 -600 5223
rect -658 5155 -600 5189
rect -658 5121 -646 5155
rect -612 5121 -600 5155
rect -658 5087 -600 5121
rect -658 5053 -646 5087
rect -612 5053 -600 5087
rect -658 5019 -600 5053
rect -658 4985 -646 5019
rect -612 4985 -600 5019
rect -658 4951 -600 4985
rect -658 4917 -646 4951
rect -612 4917 -600 4951
rect -658 4883 -600 4917
rect -658 4849 -646 4883
rect -612 4849 -600 4883
rect -658 4815 -600 4849
rect -658 4781 -646 4815
rect -612 4781 -600 4815
rect -658 4747 -600 4781
rect -658 4713 -646 4747
rect -612 4713 -600 4747
rect -658 4679 -600 4713
rect -658 4645 -646 4679
rect -612 4645 -600 4679
rect -658 4611 -600 4645
rect -658 4577 -646 4611
rect -612 4577 -600 4611
rect -658 4543 -600 4577
rect -658 4509 -646 4543
rect -612 4509 -600 4543
rect -658 4475 -600 4509
rect -658 4441 -646 4475
rect -612 4441 -600 4475
rect -658 4407 -600 4441
rect -658 4373 -646 4407
rect -612 4373 -600 4407
rect -658 4339 -600 4373
rect -658 4305 -646 4339
rect -612 4305 -600 4339
rect -658 4271 -600 4305
rect -658 4237 -646 4271
rect -612 4237 -600 4271
rect -658 4203 -600 4237
rect -658 4169 -646 4203
rect -612 4169 -600 4203
rect -658 4135 -600 4169
rect -658 4101 -646 4135
rect -612 4101 -600 4135
rect -658 4067 -600 4101
rect -658 4033 -646 4067
rect -612 4033 -600 4067
rect -658 3999 -600 4033
rect -658 3965 -646 3999
rect -612 3965 -600 3999
rect -658 3931 -600 3965
rect -658 3897 -646 3931
rect -612 3897 -600 3931
rect -658 3863 -600 3897
rect -658 3829 -646 3863
rect -612 3829 -600 3863
rect -658 3795 -600 3829
rect -658 3761 -646 3795
rect -612 3761 -600 3795
rect -658 3727 -600 3761
rect -658 3693 -646 3727
rect -612 3693 -600 3727
rect -658 3659 -600 3693
rect -658 3625 -646 3659
rect -612 3625 -600 3659
rect -658 3591 -600 3625
rect -658 3557 -646 3591
rect -612 3557 -600 3591
rect -658 3523 -600 3557
rect -658 3489 -646 3523
rect -612 3489 -600 3523
rect -658 3455 -600 3489
rect -658 3421 -646 3455
rect -612 3421 -600 3455
rect -658 3387 -600 3421
rect -658 3353 -646 3387
rect -612 3353 -600 3387
rect -658 3319 -600 3353
rect -658 3285 -646 3319
rect -612 3285 -600 3319
rect -658 3251 -600 3285
rect -658 3217 -646 3251
rect -612 3217 -600 3251
rect -658 3183 -600 3217
rect -658 3149 -646 3183
rect -612 3149 -600 3183
rect -658 3115 -600 3149
rect -658 3081 -646 3115
rect -612 3081 -600 3115
rect -658 3047 -600 3081
rect -658 3013 -646 3047
rect -612 3013 -600 3047
rect -658 2979 -600 3013
rect -658 2945 -646 2979
rect -612 2945 -600 2979
rect -658 2911 -600 2945
rect -658 2877 -646 2911
rect -612 2877 -600 2911
rect -658 2843 -600 2877
rect -658 2809 -646 2843
rect -612 2809 -600 2843
rect -658 2775 -600 2809
rect -658 2741 -646 2775
rect -612 2741 -600 2775
rect -658 2707 -600 2741
rect -658 2673 -646 2707
rect -612 2673 -600 2707
rect -658 2639 -600 2673
rect -658 2605 -646 2639
rect -612 2605 -600 2639
rect -658 2571 -600 2605
rect -658 2537 -646 2571
rect -612 2537 -600 2571
rect -658 2503 -600 2537
rect -658 2469 -646 2503
rect -612 2469 -600 2503
rect -658 2435 -600 2469
rect -658 2401 -646 2435
rect -612 2401 -600 2435
rect -658 2367 -600 2401
rect -658 2333 -646 2367
rect -612 2333 -600 2367
rect -658 2299 -600 2333
rect -658 2265 -646 2299
rect -612 2265 -600 2299
rect -658 2231 -600 2265
rect -658 2197 -646 2231
rect -612 2197 -600 2231
rect -658 2163 -600 2197
rect -658 2129 -646 2163
rect -612 2129 -600 2163
rect -658 2095 -600 2129
rect -658 2061 -646 2095
rect -612 2061 -600 2095
rect -658 2027 -600 2061
rect -658 1993 -646 2027
rect -612 1993 -600 2027
rect -658 1959 -600 1993
rect -658 1925 -646 1959
rect -612 1925 -600 1959
rect -658 1891 -600 1925
rect -658 1857 -646 1891
rect -612 1857 -600 1891
rect -658 1823 -600 1857
rect -658 1789 -646 1823
rect -612 1789 -600 1823
rect -658 1755 -600 1789
rect -658 1721 -646 1755
rect -612 1721 -600 1755
rect -658 1687 -600 1721
rect -658 1653 -646 1687
rect -612 1653 -600 1687
rect -658 1619 -600 1653
rect -658 1585 -646 1619
rect -612 1585 -600 1619
rect -658 1551 -600 1585
rect -658 1517 -646 1551
rect -612 1517 -600 1551
rect -658 1483 -600 1517
rect -658 1449 -646 1483
rect -612 1449 -600 1483
rect -658 1415 -600 1449
rect -658 1381 -646 1415
rect -612 1381 -600 1415
rect -658 1347 -600 1381
rect -658 1313 -646 1347
rect -612 1313 -600 1347
rect -658 1279 -600 1313
rect -658 1245 -646 1279
rect -612 1245 -600 1279
rect -658 1211 -600 1245
rect -658 1177 -646 1211
rect -612 1177 -600 1211
rect -658 1143 -600 1177
rect -658 1109 -646 1143
rect -612 1109 -600 1143
rect -658 1075 -600 1109
rect -658 1041 -646 1075
rect -612 1041 -600 1075
rect -658 1007 -600 1041
rect -658 973 -646 1007
rect -612 973 -600 1007
rect -658 939 -600 973
rect -658 905 -646 939
rect -612 905 -600 939
rect -658 871 -600 905
rect -658 837 -646 871
rect -612 837 -600 871
rect -658 803 -600 837
rect -658 769 -646 803
rect -612 769 -600 803
rect -658 735 -600 769
rect -658 701 -646 735
rect -612 701 -600 735
rect -658 667 -600 701
rect -658 633 -646 667
rect -612 633 -600 667
rect -658 599 -600 633
rect -658 565 -646 599
rect -612 565 -600 599
rect -658 531 -600 565
rect -658 497 -646 531
rect -612 497 -600 531
rect -658 463 -600 497
rect -658 429 -646 463
rect -612 429 -600 463
rect -658 395 -600 429
rect -658 361 -646 395
rect -612 361 -600 395
rect -658 327 -600 361
rect -658 293 -646 327
rect -612 293 -600 327
rect -658 259 -600 293
rect -658 225 -646 259
rect -612 225 -600 259
rect -658 191 -600 225
rect -658 157 -646 191
rect -612 157 -600 191
rect -658 123 -600 157
rect -658 89 -646 123
rect -612 89 -600 123
rect -658 55 -600 89
rect -658 21 -646 55
rect -612 21 -600 55
rect -658 0 -600 21
rect 750 5971 808 6000
rect 750 5937 762 5971
rect 796 5937 808 5971
rect 750 5903 808 5937
rect 750 5869 762 5903
rect 796 5869 808 5903
rect 750 5835 808 5869
rect 750 5801 762 5835
rect 796 5801 808 5835
rect 750 5767 808 5801
rect 750 5733 762 5767
rect 796 5733 808 5767
rect 750 5699 808 5733
rect 750 5665 762 5699
rect 796 5665 808 5699
rect 750 5631 808 5665
rect 750 5597 762 5631
rect 796 5597 808 5631
rect 750 5563 808 5597
rect 750 5529 762 5563
rect 796 5529 808 5563
rect 750 5495 808 5529
rect 750 5461 762 5495
rect 796 5461 808 5495
rect 750 5427 808 5461
rect 750 5393 762 5427
rect 796 5393 808 5427
rect 750 5359 808 5393
rect 750 5325 762 5359
rect 796 5325 808 5359
rect 750 5291 808 5325
rect 750 5257 762 5291
rect 796 5257 808 5291
rect 750 5223 808 5257
rect 750 5189 762 5223
rect 796 5189 808 5223
rect 750 5155 808 5189
rect 750 5121 762 5155
rect 796 5121 808 5155
rect 750 5087 808 5121
rect 750 5053 762 5087
rect 796 5053 808 5087
rect 750 5019 808 5053
rect 750 4985 762 5019
rect 796 4985 808 5019
rect 750 4951 808 4985
rect 750 4917 762 4951
rect 796 4917 808 4951
rect 750 4883 808 4917
rect 750 4849 762 4883
rect 796 4849 808 4883
rect 750 4815 808 4849
rect 750 4781 762 4815
rect 796 4781 808 4815
rect 750 4747 808 4781
rect 750 4713 762 4747
rect 796 4713 808 4747
rect 750 4679 808 4713
rect 750 4645 762 4679
rect 796 4645 808 4679
rect 750 4611 808 4645
rect 750 4577 762 4611
rect 796 4577 808 4611
rect 750 4543 808 4577
rect 750 4509 762 4543
rect 796 4509 808 4543
rect 750 4475 808 4509
rect 750 4441 762 4475
rect 796 4441 808 4475
rect 750 4407 808 4441
rect 750 4373 762 4407
rect 796 4373 808 4407
rect 750 4339 808 4373
rect 750 4305 762 4339
rect 796 4305 808 4339
rect 750 4271 808 4305
rect 750 4237 762 4271
rect 796 4237 808 4271
rect 750 4203 808 4237
rect 750 4169 762 4203
rect 796 4169 808 4203
rect 750 4135 808 4169
rect 750 4101 762 4135
rect 796 4101 808 4135
rect 750 4067 808 4101
rect 750 4033 762 4067
rect 796 4033 808 4067
rect 750 3999 808 4033
rect 750 3965 762 3999
rect 796 3965 808 3999
rect 750 3931 808 3965
rect 750 3897 762 3931
rect 796 3897 808 3931
rect 750 3863 808 3897
rect 750 3829 762 3863
rect 796 3829 808 3863
rect 750 3795 808 3829
rect 750 3761 762 3795
rect 796 3761 808 3795
rect 750 3727 808 3761
rect 750 3693 762 3727
rect 796 3693 808 3727
rect 750 3659 808 3693
rect 750 3625 762 3659
rect 796 3625 808 3659
rect 750 3591 808 3625
rect 750 3557 762 3591
rect 796 3557 808 3591
rect 750 3523 808 3557
rect 750 3489 762 3523
rect 796 3489 808 3523
rect 750 3455 808 3489
rect 750 3421 762 3455
rect 796 3421 808 3455
rect 750 3387 808 3421
rect 750 3353 762 3387
rect 796 3353 808 3387
rect 750 3319 808 3353
rect 750 3285 762 3319
rect 796 3285 808 3319
rect 750 3251 808 3285
rect 750 3217 762 3251
rect 796 3217 808 3251
rect 750 3183 808 3217
rect 750 3149 762 3183
rect 796 3149 808 3183
rect 750 3115 808 3149
rect 750 3081 762 3115
rect 796 3081 808 3115
rect 750 3047 808 3081
rect 750 3013 762 3047
rect 796 3013 808 3047
rect 750 2979 808 3013
rect 750 2945 762 2979
rect 796 2945 808 2979
rect 750 2911 808 2945
rect 750 2877 762 2911
rect 796 2877 808 2911
rect 750 2843 808 2877
rect 750 2809 762 2843
rect 796 2809 808 2843
rect 750 2775 808 2809
rect 750 2741 762 2775
rect 796 2741 808 2775
rect 750 2707 808 2741
rect 750 2673 762 2707
rect 796 2673 808 2707
rect 750 2639 808 2673
rect 750 2605 762 2639
rect 796 2605 808 2639
rect 750 2571 808 2605
rect 750 2537 762 2571
rect 796 2537 808 2571
rect 750 2503 808 2537
rect 750 2469 762 2503
rect 796 2469 808 2503
rect 750 2435 808 2469
rect 750 2401 762 2435
rect 796 2401 808 2435
rect 750 2367 808 2401
rect 750 2333 762 2367
rect 796 2333 808 2367
rect 750 2299 808 2333
rect 750 2265 762 2299
rect 796 2265 808 2299
rect 750 2231 808 2265
rect 750 2197 762 2231
rect 796 2197 808 2231
rect 750 2163 808 2197
rect 750 2129 762 2163
rect 796 2129 808 2163
rect 750 2095 808 2129
rect 750 2061 762 2095
rect 796 2061 808 2095
rect 750 2027 808 2061
rect 750 1993 762 2027
rect 796 1993 808 2027
rect 750 1959 808 1993
rect 750 1925 762 1959
rect 796 1925 808 1959
rect 750 1891 808 1925
rect 750 1857 762 1891
rect 796 1857 808 1891
rect 750 1823 808 1857
rect 750 1789 762 1823
rect 796 1789 808 1823
rect 750 1755 808 1789
rect 750 1721 762 1755
rect 796 1721 808 1755
rect 750 1687 808 1721
rect 750 1653 762 1687
rect 796 1653 808 1687
rect 750 1619 808 1653
rect 750 1585 762 1619
rect 796 1585 808 1619
rect 750 1551 808 1585
rect 750 1517 762 1551
rect 796 1517 808 1551
rect 750 1483 808 1517
rect 750 1449 762 1483
rect 796 1449 808 1483
rect 750 1415 808 1449
rect 750 1381 762 1415
rect 796 1381 808 1415
rect 750 1347 808 1381
rect 750 1313 762 1347
rect 796 1313 808 1347
rect 750 1279 808 1313
rect 750 1245 762 1279
rect 796 1245 808 1279
rect 750 1211 808 1245
rect 750 1177 762 1211
rect 796 1177 808 1211
rect 750 1143 808 1177
rect 750 1109 762 1143
rect 796 1109 808 1143
rect 750 1075 808 1109
rect 750 1041 762 1075
rect 796 1041 808 1075
rect 750 1007 808 1041
rect 750 973 762 1007
rect 796 973 808 1007
rect 750 939 808 973
rect 750 905 762 939
rect 796 905 808 939
rect 750 871 808 905
rect 750 837 762 871
rect 796 837 808 871
rect 750 803 808 837
rect 750 769 762 803
rect 796 769 808 803
rect 750 735 808 769
rect 750 701 762 735
rect 796 701 808 735
rect 750 667 808 701
rect 750 633 762 667
rect 796 633 808 667
rect 750 599 808 633
rect 750 565 762 599
rect 796 565 808 599
rect 750 531 808 565
rect 750 497 762 531
rect 796 497 808 531
rect 750 463 808 497
rect 750 429 762 463
rect 796 429 808 463
rect 750 395 808 429
rect 750 361 762 395
rect 796 361 808 395
rect 750 327 808 361
rect 750 293 762 327
rect 796 293 808 327
rect 750 259 808 293
rect 750 225 762 259
rect 796 225 808 259
rect 750 191 808 225
rect 750 157 762 191
rect 796 157 808 191
rect 750 123 808 157
rect 750 89 762 123
rect 796 89 808 123
rect 750 55 808 89
rect 750 21 762 55
rect 796 21 808 55
rect 750 0 808 21
<< mvpdiffc >>
rect -646 5937 -612 5971
rect -646 5869 -612 5903
rect -646 5801 -612 5835
rect -646 5733 -612 5767
rect -646 5665 -612 5699
rect -646 5597 -612 5631
rect -646 5529 -612 5563
rect -646 5461 -612 5495
rect -646 5393 -612 5427
rect -646 5325 -612 5359
rect -646 5257 -612 5291
rect -646 5189 -612 5223
rect -646 5121 -612 5155
rect -646 5053 -612 5087
rect -646 4985 -612 5019
rect -646 4917 -612 4951
rect -646 4849 -612 4883
rect -646 4781 -612 4815
rect -646 4713 -612 4747
rect -646 4645 -612 4679
rect -646 4577 -612 4611
rect -646 4509 -612 4543
rect -646 4441 -612 4475
rect -646 4373 -612 4407
rect -646 4305 -612 4339
rect -646 4237 -612 4271
rect -646 4169 -612 4203
rect -646 4101 -612 4135
rect -646 4033 -612 4067
rect -646 3965 -612 3999
rect -646 3897 -612 3931
rect -646 3829 -612 3863
rect -646 3761 -612 3795
rect -646 3693 -612 3727
rect -646 3625 -612 3659
rect -646 3557 -612 3591
rect -646 3489 -612 3523
rect -646 3421 -612 3455
rect -646 3353 -612 3387
rect -646 3285 -612 3319
rect -646 3217 -612 3251
rect -646 3149 -612 3183
rect -646 3081 -612 3115
rect -646 3013 -612 3047
rect -646 2945 -612 2979
rect -646 2877 -612 2911
rect -646 2809 -612 2843
rect -646 2741 -612 2775
rect -646 2673 -612 2707
rect -646 2605 -612 2639
rect -646 2537 -612 2571
rect -646 2469 -612 2503
rect -646 2401 -612 2435
rect -646 2333 -612 2367
rect -646 2265 -612 2299
rect -646 2197 -612 2231
rect -646 2129 -612 2163
rect -646 2061 -612 2095
rect -646 1993 -612 2027
rect -646 1925 -612 1959
rect -646 1857 -612 1891
rect -646 1789 -612 1823
rect -646 1721 -612 1755
rect -646 1653 -612 1687
rect -646 1585 -612 1619
rect -646 1517 -612 1551
rect -646 1449 -612 1483
rect -646 1381 -612 1415
rect -646 1313 -612 1347
rect -646 1245 -612 1279
rect -646 1177 -612 1211
rect -646 1109 -612 1143
rect -646 1041 -612 1075
rect -646 973 -612 1007
rect -646 905 -612 939
rect -646 837 -612 871
rect -646 769 -612 803
rect -646 701 -612 735
rect -646 633 -612 667
rect -646 565 -612 599
rect -646 497 -612 531
rect -646 429 -612 463
rect -646 361 -612 395
rect -646 293 -612 327
rect -646 225 -612 259
rect -646 157 -612 191
rect -646 89 -612 123
rect -646 21 -612 55
rect 762 5937 796 5971
rect 762 5869 796 5903
rect 762 5801 796 5835
rect 762 5733 796 5767
rect 762 5665 796 5699
rect 762 5597 796 5631
rect 762 5529 796 5563
rect 762 5461 796 5495
rect 762 5393 796 5427
rect 762 5325 796 5359
rect 762 5257 796 5291
rect 762 5189 796 5223
rect 762 5121 796 5155
rect 762 5053 796 5087
rect 762 4985 796 5019
rect 762 4917 796 4951
rect 762 4849 796 4883
rect 762 4781 796 4815
rect 762 4713 796 4747
rect 762 4645 796 4679
rect 762 4577 796 4611
rect 762 4509 796 4543
rect 762 4441 796 4475
rect 762 4373 796 4407
rect 762 4305 796 4339
rect 762 4237 796 4271
rect 762 4169 796 4203
rect 762 4101 796 4135
rect 762 4033 796 4067
rect 762 3965 796 3999
rect 762 3897 796 3931
rect 762 3829 796 3863
rect 762 3761 796 3795
rect 762 3693 796 3727
rect 762 3625 796 3659
rect 762 3557 796 3591
rect 762 3489 796 3523
rect 762 3421 796 3455
rect 762 3353 796 3387
rect 762 3285 796 3319
rect 762 3217 796 3251
rect 762 3149 796 3183
rect 762 3081 796 3115
rect 762 3013 796 3047
rect 762 2945 796 2979
rect 762 2877 796 2911
rect 762 2809 796 2843
rect 762 2741 796 2775
rect 762 2673 796 2707
rect 762 2605 796 2639
rect 762 2537 796 2571
rect 762 2469 796 2503
rect 762 2401 796 2435
rect 762 2333 796 2367
rect 762 2265 796 2299
rect 762 2197 796 2231
rect 762 2129 796 2163
rect 762 2061 796 2095
rect 762 1993 796 2027
rect 762 1925 796 1959
rect 762 1857 796 1891
rect 762 1789 796 1823
rect 762 1721 796 1755
rect 762 1653 796 1687
rect 762 1585 796 1619
rect 762 1517 796 1551
rect 762 1449 796 1483
rect 762 1381 796 1415
rect 762 1313 796 1347
rect 762 1245 796 1279
rect 762 1177 796 1211
rect 762 1109 796 1143
rect 762 1041 796 1075
rect 762 973 796 1007
rect 762 905 796 939
rect 762 837 796 871
rect 762 769 796 803
rect 762 701 796 735
rect 762 633 796 667
rect 762 565 796 599
rect 762 497 796 531
rect 762 429 796 463
rect 762 361 796 395
rect 762 293 796 327
rect 762 225 796 259
rect 762 157 796 191
rect 762 89 796 123
rect 762 21 796 55
<< mvpsubdiff >>
rect -1580 7780 1730 7804
rect -1580 7746 -1472 7780
rect -1438 7746 -1404 7780
rect -1370 7746 -1336 7780
rect -1302 7746 -1268 7780
rect -1234 7746 -1200 7780
rect -1166 7746 -1132 7780
rect -1098 7746 -1064 7780
rect -1030 7746 -996 7780
rect -962 7746 -928 7780
rect -894 7746 -860 7780
rect -826 7746 -792 7780
rect -758 7746 -724 7780
rect -690 7746 -656 7780
rect -622 7746 -588 7780
rect -554 7746 -520 7780
rect -486 7746 -452 7780
rect -418 7746 -384 7780
rect -350 7746 -316 7780
rect -282 7746 -248 7780
rect -214 7746 -180 7780
rect -146 7746 -112 7780
rect -78 7746 -44 7780
rect -10 7746 24 7780
rect 58 7746 92 7780
rect 126 7746 160 7780
rect 194 7746 228 7780
rect 262 7746 296 7780
rect 330 7746 364 7780
rect 398 7746 432 7780
rect 466 7746 500 7780
rect 534 7746 568 7780
rect 602 7746 636 7780
rect 670 7746 704 7780
rect 738 7746 772 7780
rect 806 7746 840 7780
rect 874 7746 908 7780
rect 942 7746 976 7780
rect 1010 7746 1044 7780
rect 1078 7746 1112 7780
rect 1146 7746 1180 7780
rect 1214 7746 1248 7780
rect 1282 7746 1316 7780
rect 1350 7746 1384 7780
rect 1418 7746 1452 7780
rect 1486 7746 1520 7780
rect 1554 7746 1588 7780
rect 1622 7746 1730 7780
rect -1580 7722 1730 7746
rect -1580 7672 -1498 7722
rect -1580 7638 -1556 7672
rect -1522 7638 -1498 7672
rect -1580 7604 -1498 7638
rect -1580 7570 -1556 7604
rect -1522 7570 -1498 7604
rect -1580 7536 -1498 7570
rect -1580 7502 -1556 7536
rect -1522 7502 -1498 7536
rect -1580 7468 -1498 7502
rect -1580 7434 -1556 7468
rect -1522 7434 -1498 7468
rect -1580 7400 -1498 7434
rect -1580 7366 -1556 7400
rect -1522 7366 -1498 7400
rect -1580 7332 -1498 7366
rect -1580 7298 -1556 7332
rect -1522 7298 -1498 7332
rect -1580 7264 -1498 7298
rect -1580 7230 -1556 7264
rect -1522 7230 -1498 7264
rect -1580 7196 -1498 7230
rect -1580 7162 -1556 7196
rect -1522 7162 -1498 7196
rect -1580 7128 -1498 7162
rect -1580 7094 -1556 7128
rect -1522 7094 -1498 7128
rect -1580 7060 -1498 7094
rect -1580 7026 -1556 7060
rect -1522 7026 -1498 7060
rect -1580 6992 -1498 7026
rect 1648 7672 1730 7722
rect 1648 7638 1672 7672
rect 1706 7638 1730 7672
rect 1648 7604 1730 7638
rect 1648 7570 1672 7604
rect 1706 7570 1730 7604
rect 1648 7536 1730 7570
rect 1648 7502 1672 7536
rect 1706 7502 1730 7536
rect 1648 7468 1730 7502
rect 1648 7434 1672 7468
rect 1706 7434 1730 7468
rect 1648 7400 1730 7434
rect 1648 7366 1672 7400
rect 1706 7366 1730 7400
rect 1648 7332 1730 7366
rect 1648 7298 1672 7332
rect 1706 7298 1730 7332
rect 1648 7264 1730 7298
rect 1648 7230 1672 7264
rect 1706 7230 1730 7264
rect 1648 7196 1730 7230
rect 1648 7162 1672 7196
rect 1706 7162 1730 7196
rect 1648 7128 1730 7162
rect 1648 7094 1672 7128
rect 1706 7094 1730 7128
rect 1648 7060 1730 7094
rect 1648 7026 1672 7060
rect 1706 7026 1730 7060
rect -1580 6958 -1556 6992
rect -1522 6958 -1498 6992
rect -1580 6924 -1498 6958
rect -1580 6890 -1556 6924
rect -1522 6890 -1498 6924
rect -1580 6856 -1498 6890
rect -1580 6822 -1556 6856
rect -1522 6822 -1498 6856
rect -1580 6788 -1498 6822
rect -1580 6754 -1556 6788
rect -1522 6754 -1498 6788
rect -1580 6720 -1498 6754
rect -1580 6686 -1556 6720
rect -1522 6686 -1498 6720
rect -1580 6652 -1498 6686
rect -1580 6618 -1556 6652
rect -1522 6618 -1498 6652
rect -1580 6584 -1498 6618
rect -1580 6550 -1556 6584
rect -1522 6550 -1498 6584
rect -1580 6516 -1498 6550
rect -1580 6482 -1556 6516
rect -1522 6482 -1498 6516
rect -1580 6448 -1498 6482
rect -1580 6414 -1556 6448
rect -1522 6414 -1498 6448
rect -1580 6380 -1498 6414
rect -1580 6346 -1556 6380
rect -1522 6346 -1498 6380
rect -1580 6312 -1498 6346
rect -1580 6278 -1556 6312
rect -1522 6278 -1498 6312
rect -1580 6244 -1498 6278
rect -1580 6210 -1556 6244
rect -1522 6210 -1498 6244
rect -1580 6176 -1498 6210
rect -1580 6142 -1556 6176
rect -1522 6142 -1498 6176
rect -1580 6108 -1498 6142
rect -1580 6074 -1556 6108
rect -1522 6074 -1498 6108
rect -1580 6040 -1498 6074
rect -1580 6006 -1556 6040
rect -1522 6006 -1498 6040
rect -1580 5972 -1498 6006
rect -1580 5938 -1556 5972
rect -1522 5938 -1498 5972
rect -1580 5904 -1498 5938
rect -1580 5870 -1556 5904
rect -1522 5870 -1498 5904
rect -1580 5836 -1498 5870
rect -1580 5802 -1556 5836
rect -1522 5802 -1498 5836
rect -1580 5768 -1498 5802
rect -1580 5734 -1556 5768
rect -1522 5734 -1498 5768
rect -1580 5700 -1498 5734
rect -1580 5666 -1556 5700
rect -1522 5666 -1498 5700
rect -1580 5632 -1498 5666
rect -1580 5598 -1556 5632
rect -1522 5598 -1498 5632
rect -1580 5564 -1498 5598
rect -1580 5530 -1556 5564
rect -1522 5530 -1498 5564
rect -1580 5496 -1498 5530
rect -1580 5462 -1556 5496
rect -1522 5462 -1498 5496
rect -1580 5428 -1498 5462
rect -1580 5394 -1556 5428
rect -1522 5394 -1498 5428
rect -1580 5360 -1498 5394
rect -1580 5326 -1556 5360
rect -1522 5326 -1498 5360
rect -1580 5292 -1498 5326
rect -1580 5258 -1556 5292
rect -1522 5258 -1498 5292
rect -1580 5224 -1498 5258
rect -1580 5190 -1556 5224
rect -1522 5190 -1498 5224
rect -1580 5156 -1498 5190
rect -1580 5122 -1556 5156
rect -1522 5122 -1498 5156
rect -1580 5088 -1498 5122
rect -1580 5054 -1556 5088
rect -1522 5054 -1498 5088
rect -1580 5020 -1498 5054
rect -1580 4986 -1556 5020
rect -1522 4986 -1498 5020
rect -1580 4952 -1498 4986
rect -1580 4918 -1556 4952
rect -1522 4918 -1498 4952
rect -1580 4884 -1498 4918
rect -1580 4850 -1556 4884
rect -1522 4850 -1498 4884
rect -1580 4816 -1498 4850
rect -1580 4782 -1556 4816
rect -1522 4782 -1498 4816
rect -1580 4748 -1498 4782
rect -1580 4714 -1556 4748
rect -1522 4714 -1498 4748
rect -1580 4680 -1498 4714
rect -1580 4646 -1556 4680
rect -1522 4646 -1498 4680
rect -1580 4612 -1498 4646
rect -1580 4578 -1556 4612
rect -1522 4578 -1498 4612
rect -1580 4544 -1498 4578
rect -1580 4510 -1556 4544
rect -1522 4510 -1498 4544
rect -1580 4476 -1498 4510
rect -1580 4442 -1556 4476
rect -1522 4442 -1498 4476
rect -1580 4408 -1498 4442
rect -1580 4374 -1556 4408
rect -1522 4374 -1498 4408
rect -1580 4340 -1498 4374
rect -1580 4306 -1556 4340
rect -1522 4306 -1498 4340
rect -1580 4272 -1498 4306
rect -1580 4238 -1556 4272
rect -1522 4238 -1498 4272
rect -1580 4204 -1498 4238
rect -1580 4170 -1556 4204
rect -1522 4170 -1498 4204
rect -1580 4136 -1498 4170
rect -1580 4102 -1556 4136
rect -1522 4102 -1498 4136
rect -1580 4068 -1498 4102
rect -1580 4034 -1556 4068
rect -1522 4034 -1498 4068
rect -1580 4000 -1498 4034
rect -1580 3966 -1556 4000
rect -1522 3966 -1498 4000
rect -1580 3932 -1498 3966
rect -1580 3898 -1556 3932
rect -1522 3898 -1498 3932
rect -1580 3864 -1498 3898
rect -1580 3830 -1556 3864
rect -1522 3830 -1498 3864
rect -1580 3796 -1498 3830
rect -1580 3762 -1556 3796
rect -1522 3762 -1498 3796
rect -1580 3728 -1498 3762
rect -1580 3694 -1556 3728
rect -1522 3694 -1498 3728
rect -1580 3660 -1498 3694
rect -1580 3626 -1556 3660
rect -1522 3626 -1498 3660
rect -1580 3592 -1498 3626
rect -1580 3558 -1556 3592
rect -1522 3558 -1498 3592
rect -1580 3524 -1498 3558
rect -1580 3490 -1556 3524
rect -1522 3490 -1498 3524
rect -1580 3456 -1498 3490
rect -1580 3422 -1556 3456
rect -1522 3422 -1498 3456
rect -1580 3388 -1498 3422
rect -1580 3354 -1556 3388
rect -1522 3354 -1498 3388
rect -1580 3320 -1498 3354
rect -1580 3286 -1556 3320
rect -1522 3286 -1498 3320
rect -1580 3252 -1498 3286
rect -1580 3218 -1556 3252
rect -1522 3218 -1498 3252
rect -1580 3184 -1498 3218
rect -1580 3150 -1556 3184
rect -1522 3150 -1498 3184
rect -1580 3116 -1498 3150
rect -1580 3082 -1556 3116
rect -1522 3082 -1498 3116
rect -1580 3048 -1498 3082
rect -1580 3014 -1556 3048
rect -1522 3014 -1498 3048
rect -1580 2980 -1498 3014
rect -1580 2946 -1556 2980
rect -1522 2946 -1498 2980
rect -1580 2912 -1498 2946
rect -1580 2878 -1556 2912
rect -1522 2878 -1498 2912
rect -1580 2844 -1498 2878
rect -1580 2810 -1556 2844
rect -1522 2810 -1498 2844
rect -1580 2776 -1498 2810
rect -1580 2742 -1556 2776
rect -1522 2742 -1498 2776
rect -1580 2708 -1498 2742
rect -1580 2674 -1556 2708
rect -1522 2674 -1498 2708
rect -1580 2640 -1498 2674
rect -1580 2606 -1556 2640
rect -1522 2606 -1498 2640
rect -1580 2572 -1498 2606
rect -1580 2538 -1556 2572
rect -1522 2538 -1498 2572
rect -1580 2504 -1498 2538
rect -1580 2470 -1556 2504
rect -1522 2470 -1498 2504
rect -1580 2436 -1498 2470
rect -1580 2402 -1556 2436
rect -1522 2402 -1498 2436
rect -1580 2368 -1498 2402
rect -1580 2334 -1556 2368
rect -1522 2334 -1498 2368
rect -1580 2300 -1498 2334
rect -1580 2266 -1556 2300
rect -1522 2266 -1498 2300
rect -1580 2232 -1498 2266
rect -1580 2198 -1556 2232
rect -1522 2198 -1498 2232
rect -1580 2164 -1498 2198
rect -1580 2130 -1556 2164
rect -1522 2130 -1498 2164
rect -1580 2096 -1498 2130
rect -1580 2062 -1556 2096
rect -1522 2062 -1498 2096
rect -1580 2028 -1498 2062
rect -1580 1994 -1556 2028
rect -1522 1994 -1498 2028
rect -1580 1960 -1498 1994
rect -1580 1926 -1556 1960
rect -1522 1926 -1498 1960
rect -1580 1892 -1498 1926
rect -1580 1858 -1556 1892
rect -1522 1858 -1498 1892
rect -1580 1824 -1498 1858
rect -1580 1790 -1556 1824
rect -1522 1790 -1498 1824
rect -1580 1756 -1498 1790
rect -1580 1722 -1556 1756
rect -1522 1722 -1498 1756
rect -1580 1688 -1498 1722
rect -1580 1654 -1556 1688
rect -1522 1654 -1498 1688
rect -1580 1620 -1498 1654
rect -1580 1586 -1556 1620
rect -1522 1586 -1498 1620
rect -1580 1552 -1498 1586
rect -1580 1518 -1556 1552
rect -1522 1518 -1498 1552
rect -1580 1484 -1498 1518
rect -1580 1450 -1556 1484
rect -1522 1450 -1498 1484
rect -1580 1416 -1498 1450
rect -1580 1382 -1556 1416
rect -1522 1382 -1498 1416
rect -1580 1348 -1498 1382
rect -1580 1314 -1556 1348
rect -1522 1314 -1498 1348
rect -1580 1280 -1498 1314
rect -1580 1246 -1556 1280
rect -1522 1246 -1498 1280
rect -1580 1212 -1498 1246
rect -1580 1178 -1556 1212
rect -1522 1178 -1498 1212
rect -1580 1144 -1498 1178
rect -1580 1110 -1556 1144
rect -1522 1110 -1498 1144
rect -1580 1076 -1498 1110
rect -1580 1042 -1556 1076
rect -1522 1042 -1498 1076
rect -1580 1008 -1498 1042
rect -1580 974 -1556 1008
rect -1522 974 -1498 1008
rect -1580 940 -1498 974
rect -1580 906 -1556 940
rect -1522 906 -1498 940
rect -1580 872 -1498 906
rect -1580 838 -1556 872
rect -1522 838 -1498 872
rect -1580 804 -1498 838
rect -1580 770 -1556 804
rect -1522 770 -1498 804
rect -1580 736 -1498 770
rect -1580 702 -1556 736
rect -1522 702 -1498 736
rect -1580 668 -1498 702
rect -1580 634 -1556 668
rect -1522 634 -1498 668
rect -1580 600 -1498 634
rect -1580 566 -1556 600
rect -1522 566 -1498 600
rect -1580 532 -1498 566
rect -1580 498 -1556 532
rect -1522 498 -1498 532
rect -1580 464 -1498 498
rect -1580 430 -1556 464
rect -1522 430 -1498 464
rect -1580 396 -1498 430
rect -1580 362 -1556 396
rect -1522 362 -1498 396
rect -1580 328 -1498 362
rect -1580 294 -1556 328
rect -1522 294 -1498 328
rect -1580 260 -1498 294
rect -1580 226 -1556 260
rect -1522 226 -1498 260
rect -1580 192 -1498 226
rect -1580 158 -1556 192
rect -1522 158 -1498 192
rect -1580 124 -1498 158
rect -1580 90 -1556 124
rect -1522 90 -1498 124
rect -1580 56 -1498 90
rect -1580 22 -1556 56
rect -1522 22 -1498 56
rect -1580 -12 -1498 22
rect -1580 -46 -1556 -12
rect -1522 -46 -1498 -12
rect -1580 -80 -1498 -46
rect -1580 -114 -1556 -80
rect -1522 -114 -1498 -80
rect -1580 -148 -1498 -114
rect -1580 -182 -1556 -148
rect -1522 -182 -1498 -148
rect -1580 -216 -1498 -182
rect -1580 -250 -1556 -216
rect -1522 -250 -1498 -216
rect -1580 -284 -1498 -250
rect -1580 -318 -1556 -284
rect -1522 -318 -1498 -284
rect -1580 -352 -1498 -318
rect -1580 -386 -1556 -352
rect -1522 -386 -1498 -352
rect -1580 -420 -1498 -386
rect -1580 -454 -1556 -420
rect -1522 -454 -1498 -420
rect -1580 -488 -1498 -454
rect -1580 -522 -1556 -488
rect -1522 -522 -1498 -488
rect -1580 -556 -1498 -522
rect -1580 -590 -1556 -556
rect -1522 -590 -1498 -556
rect -1580 -624 -1498 -590
rect -1580 -658 -1556 -624
rect -1522 -658 -1498 -624
rect -1580 -692 -1498 -658
rect -1580 -726 -1556 -692
rect -1522 -726 -1498 -692
rect -1580 -760 -1498 -726
rect -1580 -794 -1556 -760
rect -1522 -794 -1498 -760
rect -1580 -828 -1498 -794
rect -1580 -862 -1556 -828
rect -1522 -862 -1498 -828
rect -1580 -896 -1498 -862
rect -1580 -930 -1556 -896
rect -1522 -930 -1498 -896
rect -1580 -964 -1498 -930
rect -1580 -998 -1556 -964
rect -1522 -998 -1498 -964
rect -1580 -1032 -1498 -998
rect -500 0 -300 6000
tri 0 5970 30 6000 se
rect 30 5970 120 6000
tri 120 5970 150 6000 sw
rect 0 5939 150 5970
rect 0 57 24 5939
rect 126 57 150 5939
rect 0 30 150 57
tri 0 0 30 30 ne
rect 30 0 120 30
tri 120 0 150 30 nw
rect 450 0 650 6000
rect 1648 6992 1730 7026
rect 1648 6958 1672 6992
rect 1706 6958 1730 6992
rect 1648 6924 1730 6958
rect 1648 6890 1672 6924
rect 1706 6890 1730 6924
rect 1648 6856 1730 6890
rect 1648 6822 1672 6856
rect 1706 6822 1730 6856
rect 1648 6788 1730 6822
rect 1648 6754 1672 6788
rect 1706 6754 1730 6788
rect 1648 6720 1730 6754
rect 1648 6686 1672 6720
rect 1706 6686 1730 6720
rect 1648 6652 1730 6686
rect 1648 6618 1672 6652
rect 1706 6618 1730 6652
rect 1648 6584 1730 6618
rect 1648 6550 1672 6584
rect 1706 6550 1730 6584
rect 1648 6516 1730 6550
rect 1648 6482 1672 6516
rect 1706 6482 1730 6516
rect 1648 6448 1730 6482
rect 1648 6414 1672 6448
rect 1706 6414 1730 6448
rect 1648 6380 1730 6414
rect 1648 6346 1672 6380
rect 1706 6346 1730 6380
rect 1648 6312 1730 6346
rect 1648 6278 1672 6312
rect 1706 6278 1730 6312
rect 1648 6244 1730 6278
rect 1648 6210 1672 6244
rect 1706 6210 1730 6244
rect 1648 6176 1730 6210
rect 1648 6142 1672 6176
rect 1706 6142 1730 6176
rect 1648 6108 1730 6142
rect 1648 6074 1672 6108
rect 1706 6074 1730 6108
rect 1648 6040 1730 6074
rect 1648 6006 1672 6040
rect 1706 6006 1730 6040
rect 1648 5972 1730 6006
rect 1648 5938 1672 5972
rect 1706 5938 1730 5972
rect 1648 5904 1730 5938
rect 1648 5870 1672 5904
rect 1706 5870 1730 5904
rect 1648 5836 1730 5870
rect 1648 5802 1672 5836
rect 1706 5802 1730 5836
rect 1648 5768 1730 5802
rect 1648 5734 1672 5768
rect 1706 5734 1730 5768
rect 1648 5700 1730 5734
rect 1648 5666 1672 5700
rect 1706 5666 1730 5700
rect 1648 5632 1730 5666
rect 1648 5598 1672 5632
rect 1706 5598 1730 5632
rect 1648 5564 1730 5598
rect 1648 5530 1672 5564
rect 1706 5530 1730 5564
rect 1648 5496 1730 5530
rect 1648 5462 1672 5496
rect 1706 5462 1730 5496
rect 1648 5428 1730 5462
rect 1648 5394 1672 5428
rect 1706 5394 1730 5428
rect 1648 5360 1730 5394
rect 1648 5326 1672 5360
rect 1706 5326 1730 5360
rect 1648 5292 1730 5326
rect 1648 5258 1672 5292
rect 1706 5258 1730 5292
rect 1648 5224 1730 5258
rect 1648 5190 1672 5224
rect 1706 5190 1730 5224
rect 1648 5156 1730 5190
rect 1648 5122 1672 5156
rect 1706 5122 1730 5156
rect 1648 5088 1730 5122
rect 1648 5054 1672 5088
rect 1706 5054 1730 5088
rect 1648 5020 1730 5054
rect 1648 4986 1672 5020
rect 1706 4986 1730 5020
rect 1648 4952 1730 4986
rect 1648 4918 1672 4952
rect 1706 4918 1730 4952
rect 1648 4884 1730 4918
rect 1648 4850 1672 4884
rect 1706 4850 1730 4884
rect 1648 4816 1730 4850
rect 1648 4782 1672 4816
rect 1706 4782 1730 4816
rect 1648 4748 1730 4782
rect 1648 4714 1672 4748
rect 1706 4714 1730 4748
rect 1648 4680 1730 4714
rect 1648 4646 1672 4680
rect 1706 4646 1730 4680
rect 1648 4612 1730 4646
rect 1648 4578 1672 4612
rect 1706 4578 1730 4612
rect 1648 4544 1730 4578
rect 1648 4510 1672 4544
rect 1706 4510 1730 4544
rect 1648 4476 1730 4510
rect 1648 4442 1672 4476
rect 1706 4442 1730 4476
rect 1648 4408 1730 4442
rect 1648 4374 1672 4408
rect 1706 4374 1730 4408
rect 1648 4340 1730 4374
rect 1648 4306 1672 4340
rect 1706 4306 1730 4340
rect 1648 4272 1730 4306
rect 1648 4238 1672 4272
rect 1706 4238 1730 4272
rect 1648 4204 1730 4238
rect 1648 4170 1672 4204
rect 1706 4170 1730 4204
rect 1648 4136 1730 4170
rect 1648 4102 1672 4136
rect 1706 4102 1730 4136
rect 1648 4068 1730 4102
rect 1648 4034 1672 4068
rect 1706 4034 1730 4068
rect 1648 4000 1730 4034
rect 1648 3966 1672 4000
rect 1706 3966 1730 4000
rect 1648 3932 1730 3966
rect 1648 3898 1672 3932
rect 1706 3898 1730 3932
rect 1648 3864 1730 3898
rect 1648 3830 1672 3864
rect 1706 3830 1730 3864
rect 1648 3796 1730 3830
rect 1648 3762 1672 3796
rect 1706 3762 1730 3796
rect 1648 3728 1730 3762
rect 1648 3694 1672 3728
rect 1706 3694 1730 3728
rect 1648 3660 1730 3694
rect 1648 3626 1672 3660
rect 1706 3626 1730 3660
rect 1648 3592 1730 3626
rect 1648 3558 1672 3592
rect 1706 3558 1730 3592
rect 1648 3524 1730 3558
rect 1648 3490 1672 3524
rect 1706 3490 1730 3524
rect 1648 3456 1730 3490
rect 1648 3422 1672 3456
rect 1706 3422 1730 3456
rect 1648 3388 1730 3422
rect 1648 3354 1672 3388
rect 1706 3354 1730 3388
rect 1648 3320 1730 3354
rect 1648 3286 1672 3320
rect 1706 3286 1730 3320
rect 1648 3252 1730 3286
rect 1648 3218 1672 3252
rect 1706 3218 1730 3252
rect 1648 3184 1730 3218
rect 1648 3150 1672 3184
rect 1706 3150 1730 3184
rect 1648 3116 1730 3150
rect 1648 3082 1672 3116
rect 1706 3082 1730 3116
rect 1648 3048 1730 3082
rect 1648 3014 1672 3048
rect 1706 3014 1730 3048
rect 1648 2980 1730 3014
rect 1648 2946 1672 2980
rect 1706 2946 1730 2980
rect 1648 2912 1730 2946
rect 1648 2878 1672 2912
rect 1706 2878 1730 2912
rect 1648 2844 1730 2878
rect 1648 2810 1672 2844
rect 1706 2810 1730 2844
rect 1648 2776 1730 2810
rect 1648 2742 1672 2776
rect 1706 2742 1730 2776
rect 1648 2708 1730 2742
rect 1648 2674 1672 2708
rect 1706 2674 1730 2708
rect 1648 2640 1730 2674
rect 1648 2606 1672 2640
rect 1706 2606 1730 2640
rect 1648 2572 1730 2606
rect 1648 2538 1672 2572
rect 1706 2538 1730 2572
rect 1648 2504 1730 2538
rect 1648 2470 1672 2504
rect 1706 2470 1730 2504
rect 1648 2436 1730 2470
rect 1648 2402 1672 2436
rect 1706 2402 1730 2436
rect 1648 2368 1730 2402
rect 1648 2334 1672 2368
rect 1706 2334 1730 2368
rect 1648 2300 1730 2334
rect 1648 2266 1672 2300
rect 1706 2266 1730 2300
rect 1648 2232 1730 2266
rect 1648 2198 1672 2232
rect 1706 2198 1730 2232
rect 1648 2164 1730 2198
rect 1648 2130 1672 2164
rect 1706 2130 1730 2164
rect 1648 2096 1730 2130
rect 1648 2062 1672 2096
rect 1706 2062 1730 2096
rect 1648 2028 1730 2062
rect 1648 1994 1672 2028
rect 1706 1994 1730 2028
rect 1648 1960 1730 1994
rect 1648 1926 1672 1960
rect 1706 1926 1730 1960
rect 1648 1892 1730 1926
rect 1648 1858 1672 1892
rect 1706 1858 1730 1892
rect 1648 1824 1730 1858
rect 1648 1790 1672 1824
rect 1706 1790 1730 1824
rect 1648 1756 1730 1790
rect 1648 1722 1672 1756
rect 1706 1722 1730 1756
rect 1648 1688 1730 1722
rect 1648 1654 1672 1688
rect 1706 1654 1730 1688
rect 1648 1620 1730 1654
rect 1648 1586 1672 1620
rect 1706 1586 1730 1620
rect 1648 1552 1730 1586
rect 1648 1518 1672 1552
rect 1706 1518 1730 1552
rect 1648 1484 1730 1518
rect 1648 1450 1672 1484
rect 1706 1450 1730 1484
rect 1648 1416 1730 1450
rect 1648 1382 1672 1416
rect 1706 1382 1730 1416
rect 1648 1348 1730 1382
rect 1648 1314 1672 1348
rect 1706 1314 1730 1348
rect 1648 1280 1730 1314
rect 1648 1246 1672 1280
rect 1706 1246 1730 1280
rect 1648 1212 1730 1246
rect 1648 1178 1672 1212
rect 1706 1178 1730 1212
rect 1648 1144 1730 1178
rect 1648 1110 1672 1144
rect 1706 1110 1730 1144
rect 1648 1076 1730 1110
rect 1648 1042 1672 1076
rect 1706 1042 1730 1076
rect 1648 1008 1730 1042
rect 1648 974 1672 1008
rect 1706 974 1730 1008
rect 1648 940 1730 974
rect 1648 906 1672 940
rect 1706 906 1730 940
rect 1648 872 1730 906
rect 1648 838 1672 872
rect 1706 838 1730 872
rect 1648 804 1730 838
rect 1648 770 1672 804
rect 1706 770 1730 804
rect 1648 736 1730 770
rect 1648 702 1672 736
rect 1706 702 1730 736
rect 1648 668 1730 702
rect 1648 634 1672 668
rect 1706 634 1730 668
rect 1648 600 1730 634
rect 1648 566 1672 600
rect 1706 566 1730 600
rect 1648 532 1730 566
rect 1648 498 1672 532
rect 1706 498 1730 532
rect 1648 464 1730 498
rect 1648 430 1672 464
rect 1706 430 1730 464
rect 1648 396 1730 430
rect 1648 362 1672 396
rect 1706 362 1730 396
rect 1648 328 1730 362
rect 1648 294 1672 328
rect 1706 294 1730 328
rect 1648 260 1730 294
rect 1648 226 1672 260
rect 1706 226 1730 260
rect 1648 192 1730 226
rect 1648 158 1672 192
rect 1706 158 1730 192
rect 1648 124 1730 158
rect 1648 90 1672 124
rect 1706 90 1730 124
rect 1648 56 1730 90
rect 1648 22 1672 56
rect 1706 22 1730 56
rect 1648 -12 1730 22
rect 1648 -46 1672 -12
rect 1706 -46 1730 -12
rect 1648 -80 1730 -46
rect 1648 -114 1672 -80
rect 1706 -114 1730 -80
rect 1648 -148 1730 -114
rect 1648 -182 1672 -148
rect 1706 -182 1730 -148
rect 1648 -216 1730 -182
rect 1648 -250 1672 -216
rect 1706 -250 1730 -216
rect 1648 -284 1730 -250
rect 1648 -318 1672 -284
rect 1706 -318 1730 -284
rect 1648 -352 1730 -318
rect 1648 -386 1672 -352
rect 1706 -386 1730 -352
rect 1648 -420 1730 -386
rect 1648 -454 1672 -420
rect 1706 -454 1730 -420
rect 1648 -488 1730 -454
rect 1648 -522 1672 -488
rect 1706 -522 1730 -488
rect 1648 -556 1730 -522
rect 1648 -590 1672 -556
rect 1706 -590 1730 -556
rect 1648 -624 1730 -590
rect 1648 -658 1672 -624
rect 1706 -658 1730 -624
rect 1648 -692 1730 -658
rect 1648 -726 1672 -692
rect 1706 -726 1730 -692
rect 1648 -760 1730 -726
rect 1648 -794 1672 -760
rect 1706 -794 1730 -760
rect 1648 -828 1730 -794
rect 1648 -862 1672 -828
rect 1706 -862 1730 -828
rect 1648 -896 1730 -862
rect 1648 -930 1672 -896
rect 1706 -930 1730 -896
rect 1648 -964 1730 -930
rect 1648 -998 1672 -964
rect 1706 -998 1730 -964
rect -1580 -1066 -1556 -1032
rect -1522 -1066 -1498 -1032
rect -1580 -1100 -1498 -1066
rect -1580 -1134 -1556 -1100
rect -1522 -1134 -1498 -1100
rect -1580 -1168 -1498 -1134
rect -1580 -1202 -1556 -1168
rect -1522 -1202 -1498 -1168
rect -1580 -1236 -1498 -1202
rect -1580 -1270 -1556 -1236
rect -1522 -1270 -1498 -1236
rect -1580 -1304 -1498 -1270
rect -1580 -1338 -1556 -1304
rect -1522 -1338 -1498 -1304
rect -1580 -1372 -1498 -1338
rect -1580 -1406 -1556 -1372
rect -1522 -1406 -1498 -1372
rect -1580 -1440 -1498 -1406
rect -1580 -1474 -1556 -1440
rect -1522 -1474 -1498 -1440
rect -1580 -1508 -1498 -1474
rect -1580 -1542 -1556 -1508
rect -1522 -1542 -1498 -1508
rect -1580 -1576 -1498 -1542
rect -1580 -1610 -1556 -1576
rect -1522 -1610 -1498 -1576
rect -1580 -1644 -1498 -1610
rect -1580 -1678 -1556 -1644
rect -1522 -1678 -1498 -1644
rect -1580 -1722 -1498 -1678
rect 1648 -1032 1730 -998
rect 1648 -1066 1672 -1032
rect 1706 -1066 1730 -1032
rect 1648 -1100 1730 -1066
rect 1648 -1134 1672 -1100
rect 1706 -1134 1730 -1100
rect 1648 -1168 1730 -1134
rect 1648 -1202 1672 -1168
rect 1706 -1202 1730 -1168
rect 1648 -1236 1730 -1202
rect 1648 -1270 1672 -1236
rect 1706 -1270 1730 -1236
rect 1648 -1304 1730 -1270
rect 1648 -1338 1672 -1304
rect 1706 -1338 1730 -1304
rect 1648 -1372 1730 -1338
rect 1648 -1406 1672 -1372
rect 1706 -1406 1730 -1372
rect 1648 -1440 1730 -1406
rect 1648 -1474 1672 -1440
rect 1706 -1474 1730 -1440
rect 1648 -1508 1730 -1474
rect 1648 -1542 1672 -1508
rect 1706 -1542 1730 -1508
rect 1648 -1576 1730 -1542
rect 1648 -1610 1672 -1576
rect 1706 -1610 1730 -1576
rect 1648 -1644 1730 -1610
rect 1648 -1678 1672 -1644
rect 1706 -1678 1730 -1644
rect 1648 -1722 1730 -1678
rect -1580 -1746 1730 -1722
rect -1580 -1780 -1472 -1746
rect -1438 -1780 -1404 -1746
rect -1370 -1780 -1336 -1746
rect -1302 -1780 -1268 -1746
rect -1234 -1780 -1200 -1746
rect -1166 -1780 -1132 -1746
rect -1098 -1780 -1064 -1746
rect -1030 -1780 -996 -1746
rect -962 -1780 -928 -1746
rect -894 -1780 -860 -1746
rect -826 -1780 -792 -1746
rect -758 -1780 -724 -1746
rect -690 -1780 -656 -1746
rect -622 -1780 -588 -1746
rect -554 -1780 -520 -1746
rect -486 -1780 -452 -1746
rect -418 -1780 -384 -1746
rect -350 -1780 -316 -1746
rect -282 -1780 -248 -1746
rect -214 -1780 -180 -1746
rect -146 -1780 -112 -1746
rect -78 -1780 -44 -1746
rect -10 -1780 24 -1746
rect 58 -1780 92 -1746
rect 126 -1780 160 -1746
rect 194 -1780 228 -1746
rect 262 -1780 296 -1746
rect 330 -1780 364 -1746
rect 398 -1780 432 -1746
rect 466 -1780 500 -1746
rect 534 -1780 568 -1746
rect 602 -1780 636 -1746
rect 670 -1780 704 -1746
rect 738 -1780 772 -1746
rect 806 -1780 840 -1746
rect 874 -1780 908 -1746
rect 942 -1780 976 -1746
rect 1010 -1780 1044 -1746
rect 1078 -1780 1112 -1746
rect 1146 -1780 1180 -1746
rect 1214 -1780 1248 -1746
rect 1282 -1780 1316 -1746
rect 1350 -1780 1384 -1746
rect 1418 -1780 1452 -1746
rect 1486 -1780 1520 -1746
rect 1554 -1780 1588 -1746
rect 1622 -1780 1730 -1746
rect -1580 -1804 1730 -1780
<< mvnsubdiff >>
rect -798 6998 948 7022
rect -798 6964 -520 6998
rect -486 6964 -452 6998
rect -418 6964 -384 6998
rect -350 6964 -316 6998
rect -282 6964 -248 6998
rect -214 6964 -180 6998
rect -146 6964 -112 6998
rect -78 6964 -44 6998
rect -10 6964 24 6998
rect 58 6964 92 6998
rect 126 6964 160 6998
rect 194 6964 228 6998
rect 262 6964 296 6998
rect 330 6964 364 6998
rect 398 6964 432 6998
rect 466 6964 500 6998
rect 534 6964 568 6998
rect 602 6964 636 6998
rect 670 6964 948 6998
rect -798 6940 948 6964
rect -798 6856 -716 6940
rect -798 6822 -774 6856
rect -740 6822 -716 6856
rect -798 6788 -716 6822
rect 866 6856 948 6940
rect 866 6822 890 6856
rect 924 6822 948 6856
rect -798 6754 -774 6788
rect -740 6754 -716 6788
rect -798 6720 -716 6754
rect -798 6686 -774 6720
rect -740 6686 -716 6720
rect -798 6652 -716 6686
rect -798 6618 -774 6652
rect -740 6618 -716 6652
rect -798 6584 -716 6618
rect -798 6550 -774 6584
rect -740 6550 -716 6584
rect -798 6516 -716 6550
rect -798 6482 -774 6516
rect -740 6482 -716 6516
rect -798 6448 -716 6482
rect -798 6414 -774 6448
rect -740 6414 -716 6448
rect -798 6380 -716 6414
rect -798 6346 -774 6380
rect -740 6346 -716 6380
rect -798 6312 -716 6346
rect -798 6278 -774 6312
rect -740 6278 -716 6312
rect -798 6244 -716 6278
rect -798 6210 -774 6244
rect -740 6210 -716 6244
rect -798 6176 -716 6210
rect -798 6142 -774 6176
rect -740 6142 -716 6176
rect -798 6108 -716 6142
rect -798 6074 -774 6108
rect -740 6074 -716 6108
rect -798 6040 -716 6074
rect -798 6006 -774 6040
rect -740 6006 -716 6040
rect -798 5972 -716 6006
rect 866 6788 948 6822
rect 866 6754 890 6788
rect 924 6754 948 6788
rect 866 6720 948 6754
rect 866 6686 890 6720
rect 924 6686 948 6720
rect 866 6652 948 6686
rect 866 6618 890 6652
rect 924 6618 948 6652
rect 866 6584 948 6618
rect 866 6550 890 6584
rect 924 6550 948 6584
rect 866 6516 948 6550
rect 866 6482 890 6516
rect 924 6482 948 6516
rect 866 6448 948 6482
rect 866 6414 890 6448
rect 924 6414 948 6448
rect 866 6380 948 6414
rect 866 6346 890 6380
rect 924 6346 948 6380
rect 866 6312 948 6346
rect 866 6278 890 6312
rect 924 6278 948 6312
rect 866 6244 948 6278
rect 866 6210 890 6244
rect 924 6210 948 6244
rect 866 6176 948 6210
rect 866 6142 890 6176
rect 924 6142 948 6176
rect 866 6108 948 6142
rect 866 6074 890 6108
rect 924 6074 948 6108
rect 866 6040 948 6074
rect 866 6006 890 6040
rect 924 6006 948 6040
rect -798 5938 -774 5972
rect -740 5938 -716 5972
rect -798 5904 -716 5938
rect -798 5870 -774 5904
rect -740 5870 -716 5904
rect -798 5836 -716 5870
rect -798 5802 -774 5836
rect -740 5802 -716 5836
rect -798 5768 -716 5802
rect -798 5734 -774 5768
rect -740 5734 -716 5768
rect -798 5700 -716 5734
rect -798 5666 -774 5700
rect -740 5666 -716 5700
rect -798 5632 -716 5666
rect -798 5598 -774 5632
rect -740 5598 -716 5632
rect -798 5564 -716 5598
rect -798 5530 -774 5564
rect -740 5530 -716 5564
rect -798 5496 -716 5530
rect -798 5462 -774 5496
rect -740 5462 -716 5496
rect -798 5428 -716 5462
rect -798 5394 -774 5428
rect -740 5394 -716 5428
rect -798 5360 -716 5394
rect -798 5326 -774 5360
rect -740 5326 -716 5360
rect -798 5292 -716 5326
rect -798 5258 -774 5292
rect -740 5258 -716 5292
rect -798 5224 -716 5258
rect -798 5190 -774 5224
rect -740 5190 -716 5224
rect -798 5156 -716 5190
rect -798 5122 -774 5156
rect -740 5122 -716 5156
rect -798 5088 -716 5122
rect -798 5054 -774 5088
rect -740 5054 -716 5088
rect -798 5020 -716 5054
rect -798 4986 -774 5020
rect -740 4986 -716 5020
rect -798 4952 -716 4986
rect -798 4918 -774 4952
rect -740 4918 -716 4952
rect -798 4884 -716 4918
rect -798 4850 -774 4884
rect -740 4850 -716 4884
rect -798 4816 -716 4850
rect -798 4782 -774 4816
rect -740 4782 -716 4816
rect -798 4748 -716 4782
rect -798 4714 -774 4748
rect -740 4714 -716 4748
rect -798 4680 -716 4714
rect -798 4646 -774 4680
rect -740 4646 -716 4680
rect -798 4612 -716 4646
rect -798 4578 -774 4612
rect -740 4578 -716 4612
rect -798 4544 -716 4578
rect -798 4510 -774 4544
rect -740 4510 -716 4544
rect -798 4476 -716 4510
rect -798 4442 -774 4476
rect -740 4442 -716 4476
rect -798 4408 -716 4442
rect -798 4374 -774 4408
rect -740 4374 -716 4408
rect -798 4340 -716 4374
rect -798 4306 -774 4340
rect -740 4306 -716 4340
rect -798 4272 -716 4306
rect -798 4238 -774 4272
rect -740 4238 -716 4272
rect -798 4204 -716 4238
rect -798 4170 -774 4204
rect -740 4170 -716 4204
rect -798 4136 -716 4170
rect -798 4102 -774 4136
rect -740 4102 -716 4136
rect -798 4068 -716 4102
rect -798 4034 -774 4068
rect -740 4034 -716 4068
rect -798 4000 -716 4034
rect -798 3966 -774 4000
rect -740 3966 -716 4000
rect -798 3932 -716 3966
rect -798 3898 -774 3932
rect -740 3898 -716 3932
rect -798 3864 -716 3898
rect -798 3830 -774 3864
rect -740 3830 -716 3864
rect -798 3796 -716 3830
rect -798 3762 -774 3796
rect -740 3762 -716 3796
rect -798 3728 -716 3762
rect -798 3694 -774 3728
rect -740 3694 -716 3728
rect -798 3660 -716 3694
rect -798 3626 -774 3660
rect -740 3626 -716 3660
rect -798 3592 -716 3626
rect -798 3558 -774 3592
rect -740 3558 -716 3592
rect -798 3524 -716 3558
rect -798 3490 -774 3524
rect -740 3490 -716 3524
rect -798 3456 -716 3490
rect -798 3422 -774 3456
rect -740 3422 -716 3456
rect -798 3388 -716 3422
rect -798 3354 -774 3388
rect -740 3354 -716 3388
rect -798 3320 -716 3354
rect -798 3286 -774 3320
rect -740 3286 -716 3320
rect -798 3252 -716 3286
rect -798 3218 -774 3252
rect -740 3218 -716 3252
rect -798 3184 -716 3218
rect -798 3150 -774 3184
rect -740 3150 -716 3184
rect -798 3116 -716 3150
rect -798 3082 -774 3116
rect -740 3082 -716 3116
rect -798 3048 -716 3082
rect -798 3014 -774 3048
rect -740 3014 -716 3048
rect -798 2980 -716 3014
rect -798 2946 -774 2980
rect -740 2946 -716 2980
rect -798 2912 -716 2946
rect -798 2878 -774 2912
rect -740 2878 -716 2912
rect -798 2844 -716 2878
rect -798 2810 -774 2844
rect -740 2810 -716 2844
rect -798 2776 -716 2810
rect -798 2742 -774 2776
rect -740 2742 -716 2776
rect -798 2708 -716 2742
rect -798 2674 -774 2708
rect -740 2674 -716 2708
rect -798 2640 -716 2674
rect -798 2606 -774 2640
rect -740 2606 -716 2640
rect -798 2572 -716 2606
rect -798 2538 -774 2572
rect -740 2538 -716 2572
rect -798 2504 -716 2538
rect -798 2470 -774 2504
rect -740 2470 -716 2504
rect -798 2436 -716 2470
rect -798 2402 -774 2436
rect -740 2402 -716 2436
rect -798 2368 -716 2402
rect -798 2334 -774 2368
rect -740 2334 -716 2368
rect -798 2300 -716 2334
rect -798 2266 -774 2300
rect -740 2266 -716 2300
rect -798 2232 -716 2266
rect -798 2198 -774 2232
rect -740 2198 -716 2232
rect -798 2164 -716 2198
rect -798 2130 -774 2164
rect -740 2130 -716 2164
rect -798 2096 -716 2130
rect -798 2062 -774 2096
rect -740 2062 -716 2096
rect -798 2028 -716 2062
rect -798 1994 -774 2028
rect -740 1994 -716 2028
rect -798 1960 -716 1994
rect -798 1926 -774 1960
rect -740 1926 -716 1960
rect -798 1892 -716 1926
rect -798 1858 -774 1892
rect -740 1858 -716 1892
rect -798 1824 -716 1858
rect -798 1790 -774 1824
rect -740 1790 -716 1824
rect -798 1756 -716 1790
rect -798 1722 -774 1756
rect -740 1722 -716 1756
rect -798 1688 -716 1722
rect -798 1654 -774 1688
rect -740 1654 -716 1688
rect -798 1620 -716 1654
rect -798 1586 -774 1620
rect -740 1586 -716 1620
rect -798 1552 -716 1586
rect -798 1518 -774 1552
rect -740 1518 -716 1552
rect -798 1484 -716 1518
rect -798 1450 -774 1484
rect -740 1450 -716 1484
rect -798 1416 -716 1450
rect -798 1382 -774 1416
rect -740 1382 -716 1416
rect -798 1348 -716 1382
rect -798 1314 -774 1348
rect -740 1314 -716 1348
rect -798 1280 -716 1314
rect -798 1246 -774 1280
rect -740 1246 -716 1280
rect -798 1212 -716 1246
rect -798 1178 -774 1212
rect -740 1178 -716 1212
rect -798 1144 -716 1178
rect -798 1110 -774 1144
rect -740 1110 -716 1144
rect -798 1076 -716 1110
rect -798 1042 -774 1076
rect -740 1042 -716 1076
rect -798 1008 -716 1042
rect -798 974 -774 1008
rect -740 974 -716 1008
rect -798 940 -716 974
rect -798 906 -774 940
rect -740 906 -716 940
rect -798 872 -716 906
rect -798 838 -774 872
rect -740 838 -716 872
rect -798 804 -716 838
rect -798 770 -774 804
rect -740 770 -716 804
rect -798 736 -716 770
rect -798 702 -774 736
rect -740 702 -716 736
rect -798 668 -716 702
rect -798 634 -774 668
rect -740 634 -716 668
rect -798 600 -716 634
rect -798 566 -774 600
rect -740 566 -716 600
rect -798 532 -716 566
rect -798 498 -774 532
rect -740 498 -716 532
rect -798 464 -716 498
rect -798 430 -774 464
rect -740 430 -716 464
rect -798 396 -716 430
rect -798 362 -774 396
rect -740 362 -716 396
rect -798 328 -716 362
rect -798 294 -774 328
rect -740 294 -716 328
rect -798 260 -716 294
rect -798 226 -774 260
rect -740 226 -716 260
rect -798 192 -716 226
rect -798 158 -774 192
rect -740 158 -716 192
rect -798 124 -716 158
rect -798 90 -774 124
rect -740 90 -716 124
rect -798 56 -716 90
rect -798 22 -774 56
rect -740 22 -716 56
rect -798 -12 -716 22
rect 866 5972 948 6006
rect 866 5938 890 5972
rect 924 5938 948 5972
rect 866 5904 948 5938
rect 866 5870 890 5904
rect 924 5870 948 5904
rect 866 5836 948 5870
rect 866 5802 890 5836
rect 924 5802 948 5836
rect 866 5768 948 5802
rect 866 5734 890 5768
rect 924 5734 948 5768
rect 866 5700 948 5734
rect 866 5666 890 5700
rect 924 5666 948 5700
rect 866 5632 948 5666
rect 866 5598 890 5632
rect 924 5598 948 5632
rect 866 5564 948 5598
rect 866 5530 890 5564
rect 924 5530 948 5564
rect 866 5496 948 5530
rect 866 5462 890 5496
rect 924 5462 948 5496
rect 866 5428 948 5462
rect 866 5394 890 5428
rect 924 5394 948 5428
rect 866 5360 948 5394
rect 866 5326 890 5360
rect 924 5326 948 5360
rect 866 5292 948 5326
rect 866 5258 890 5292
rect 924 5258 948 5292
rect 866 5224 948 5258
rect 866 5190 890 5224
rect 924 5190 948 5224
rect 866 5156 948 5190
rect 866 5122 890 5156
rect 924 5122 948 5156
rect 866 5088 948 5122
rect 866 5054 890 5088
rect 924 5054 948 5088
rect 866 5020 948 5054
rect 866 4986 890 5020
rect 924 4986 948 5020
rect 866 4952 948 4986
rect 866 4918 890 4952
rect 924 4918 948 4952
rect 866 4884 948 4918
rect 866 4850 890 4884
rect 924 4850 948 4884
rect 866 4816 948 4850
rect 866 4782 890 4816
rect 924 4782 948 4816
rect 866 4748 948 4782
rect 866 4714 890 4748
rect 924 4714 948 4748
rect 866 4680 948 4714
rect 866 4646 890 4680
rect 924 4646 948 4680
rect 866 4612 948 4646
rect 866 4578 890 4612
rect 924 4578 948 4612
rect 866 4544 948 4578
rect 866 4510 890 4544
rect 924 4510 948 4544
rect 866 4476 948 4510
rect 866 4442 890 4476
rect 924 4442 948 4476
rect 866 4408 948 4442
rect 866 4374 890 4408
rect 924 4374 948 4408
rect 866 4340 948 4374
rect 866 4306 890 4340
rect 924 4306 948 4340
rect 866 4272 948 4306
rect 866 4238 890 4272
rect 924 4238 948 4272
rect 866 4204 948 4238
rect 866 4170 890 4204
rect 924 4170 948 4204
rect 866 4136 948 4170
rect 866 4102 890 4136
rect 924 4102 948 4136
rect 866 4068 948 4102
rect 866 4034 890 4068
rect 924 4034 948 4068
rect 866 4000 948 4034
rect 866 3966 890 4000
rect 924 3966 948 4000
rect 866 3932 948 3966
rect 866 3898 890 3932
rect 924 3898 948 3932
rect 866 3864 948 3898
rect 866 3830 890 3864
rect 924 3830 948 3864
rect 866 3796 948 3830
rect 866 3762 890 3796
rect 924 3762 948 3796
rect 866 3728 948 3762
rect 866 3694 890 3728
rect 924 3694 948 3728
rect 866 3660 948 3694
rect 866 3626 890 3660
rect 924 3626 948 3660
rect 866 3592 948 3626
rect 866 3558 890 3592
rect 924 3558 948 3592
rect 866 3524 948 3558
rect 866 3490 890 3524
rect 924 3490 948 3524
rect 866 3456 948 3490
rect 866 3422 890 3456
rect 924 3422 948 3456
rect 866 3388 948 3422
rect 866 3354 890 3388
rect 924 3354 948 3388
rect 866 3320 948 3354
rect 866 3286 890 3320
rect 924 3286 948 3320
rect 866 3252 948 3286
rect 866 3218 890 3252
rect 924 3218 948 3252
rect 866 3184 948 3218
rect 866 3150 890 3184
rect 924 3150 948 3184
rect 866 3116 948 3150
rect 866 3082 890 3116
rect 924 3082 948 3116
rect 866 3048 948 3082
rect 866 3014 890 3048
rect 924 3014 948 3048
rect 866 2980 948 3014
rect 866 2946 890 2980
rect 924 2946 948 2980
rect 866 2912 948 2946
rect 866 2878 890 2912
rect 924 2878 948 2912
rect 866 2844 948 2878
rect 866 2810 890 2844
rect 924 2810 948 2844
rect 866 2776 948 2810
rect 866 2742 890 2776
rect 924 2742 948 2776
rect 866 2708 948 2742
rect 866 2674 890 2708
rect 924 2674 948 2708
rect 866 2640 948 2674
rect 866 2606 890 2640
rect 924 2606 948 2640
rect 866 2572 948 2606
rect 866 2538 890 2572
rect 924 2538 948 2572
rect 866 2504 948 2538
rect 866 2470 890 2504
rect 924 2470 948 2504
rect 866 2436 948 2470
rect 866 2402 890 2436
rect 924 2402 948 2436
rect 866 2368 948 2402
rect 866 2334 890 2368
rect 924 2334 948 2368
rect 866 2300 948 2334
rect 866 2266 890 2300
rect 924 2266 948 2300
rect 866 2232 948 2266
rect 866 2198 890 2232
rect 924 2198 948 2232
rect 866 2164 948 2198
rect 866 2130 890 2164
rect 924 2130 948 2164
rect 866 2096 948 2130
rect 866 2062 890 2096
rect 924 2062 948 2096
rect 866 2028 948 2062
rect 866 1994 890 2028
rect 924 1994 948 2028
rect 866 1960 948 1994
rect 866 1926 890 1960
rect 924 1926 948 1960
rect 866 1892 948 1926
rect 866 1858 890 1892
rect 924 1858 948 1892
rect 866 1824 948 1858
rect 866 1790 890 1824
rect 924 1790 948 1824
rect 866 1756 948 1790
rect 866 1722 890 1756
rect 924 1722 948 1756
rect 866 1688 948 1722
rect 866 1654 890 1688
rect 924 1654 948 1688
rect 866 1620 948 1654
rect 866 1586 890 1620
rect 924 1586 948 1620
rect 866 1552 948 1586
rect 866 1518 890 1552
rect 924 1518 948 1552
rect 866 1484 948 1518
rect 866 1450 890 1484
rect 924 1450 948 1484
rect 866 1416 948 1450
rect 866 1382 890 1416
rect 924 1382 948 1416
rect 866 1348 948 1382
rect 866 1314 890 1348
rect 924 1314 948 1348
rect 866 1280 948 1314
rect 866 1246 890 1280
rect 924 1246 948 1280
rect 866 1212 948 1246
rect 866 1178 890 1212
rect 924 1178 948 1212
rect 866 1144 948 1178
rect 866 1110 890 1144
rect 924 1110 948 1144
rect 866 1076 948 1110
rect 866 1042 890 1076
rect 924 1042 948 1076
rect 866 1008 948 1042
rect 866 974 890 1008
rect 924 974 948 1008
rect 866 940 948 974
rect 866 906 890 940
rect 924 906 948 940
rect 866 872 948 906
rect 866 838 890 872
rect 924 838 948 872
rect 866 804 948 838
rect 866 770 890 804
rect 924 770 948 804
rect 866 736 948 770
rect 866 702 890 736
rect 924 702 948 736
rect 866 668 948 702
rect 866 634 890 668
rect 924 634 948 668
rect 866 600 948 634
rect 866 566 890 600
rect 924 566 948 600
rect 866 532 948 566
rect 866 498 890 532
rect 924 498 948 532
rect 866 464 948 498
rect 866 430 890 464
rect 924 430 948 464
rect 866 396 948 430
rect 866 362 890 396
rect 924 362 948 396
rect 866 328 948 362
rect 866 294 890 328
rect 924 294 948 328
rect 866 260 948 294
rect 866 226 890 260
rect 924 226 948 260
rect 866 192 948 226
rect 866 158 890 192
rect 924 158 948 192
rect 866 124 948 158
rect 866 90 890 124
rect 924 90 948 124
rect 866 56 948 90
rect 866 22 890 56
rect 924 22 948 56
rect -798 -46 -774 -12
rect -740 -46 -716 -12
rect -798 -80 -716 -46
rect -798 -114 -774 -80
rect -740 -114 -716 -80
rect -798 -148 -716 -114
rect -798 -182 -774 -148
rect -740 -182 -716 -148
rect -798 -216 -716 -182
rect -798 -250 -774 -216
rect -740 -250 -716 -216
rect -798 -284 -716 -250
rect -798 -318 -774 -284
rect -740 -318 -716 -284
rect -798 -352 -716 -318
rect -798 -386 -774 -352
rect -740 -386 -716 -352
rect -798 -420 -716 -386
rect -798 -454 -774 -420
rect -740 -454 -716 -420
rect -798 -488 -716 -454
rect -798 -522 -774 -488
rect -740 -522 -716 -488
rect -798 -556 -716 -522
rect -798 -590 -774 -556
rect -740 -590 -716 -556
rect -798 -624 -716 -590
rect -798 -658 -774 -624
rect -740 -658 -716 -624
rect -798 -692 -716 -658
rect -798 -726 -774 -692
rect -740 -726 -716 -692
rect -798 -760 -716 -726
rect -798 -794 -774 -760
rect -740 -794 -716 -760
rect -798 -828 -716 -794
rect 866 -12 948 22
rect 866 -46 890 -12
rect 924 -46 948 -12
rect 866 -80 948 -46
rect 866 -114 890 -80
rect 924 -114 948 -80
rect 866 -148 948 -114
rect 866 -182 890 -148
rect 924 -182 948 -148
rect 866 -216 948 -182
rect 866 -250 890 -216
rect 924 -250 948 -216
rect 866 -284 948 -250
rect 866 -318 890 -284
rect 924 -318 948 -284
rect 866 -352 948 -318
rect 866 -386 890 -352
rect 924 -386 948 -352
rect 866 -420 948 -386
rect 866 -454 890 -420
rect 924 -454 948 -420
rect 866 -488 948 -454
rect 866 -522 890 -488
rect 924 -522 948 -488
rect 866 -556 948 -522
rect 866 -590 890 -556
rect 924 -590 948 -556
rect 866 -624 948 -590
rect 866 -658 890 -624
rect 924 -658 948 -624
rect 866 -692 948 -658
rect 866 -726 890 -692
rect 924 -726 948 -692
rect 866 -760 948 -726
rect 866 -794 890 -760
rect 924 -794 948 -760
rect -798 -862 -774 -828
rect -740 -862 -716 -828
rect -798 -896 -716 -862
rect -798 -930 -774 -896
rect -740 -930 -716 -896
rect -798 -940 -716 -930
rect 866 -828 948 -794
rect 866 -862 890 -828
rect 924 -862 948 -828
rect 866 -896 948 -862
rect 866 -930 890 -896
rect 924 -930 948 -896
rect 866 -940 948 -930
rect -798 -964 948 -940
rect -798 -998 -774 -964
rect -740 -998 -520 -964
rect -486 -998 -452 -964
rect -418 -998 -384 -964
rect -350 -998 -316 -964
rect -282 -998 -248 -964
rect -214 -998 -180 -964
rect -146 -998 -112 -964
rect -78 -998 -44 -964
rect -10 -998 24 -964
rect 58 -998 92 -964
rect 126 -998 160 -964
rect 194 -998 228 -964
rect 262 -998 296 -964
rect 330 -998 364 -964
rect 398 -998 432 -964
rect 466 -998 500 -964
rect 534 -998 568 -964
rect 602 -998 636 -964
rect 670 -998 890 -964
rect 924 -998 948 -964
rect -798 -1022 948 -998
<< mvpsubdiffcont >>
rect -1472 7746 -1438 7780
rect -1404 7746 -1370 7780
rect -1336 7746 -1302 7780
rect -1268 7746 -1234 7780
rect -1200 7746 -1166 7780
rect -1132 7746 -1098 7780
rect -1064 7746 -1030 7780
rect -996 7746 -962 7780
rect -928 7746 -894 7780
rect -860 7746 -826 7780
rect -792 7746 -758 7780
rect -724 7746 -690 7780
rect -656 7746 -622 7780
rect -588 7746 -554 7780
rect -520 7746 -486 7780
rect -452 7746 -418 7780
rect -384 7746 -350 7780
rect -316 7746 -282 7780
rect -248 7746 -214 7780
rect -180 7746 -146 7780
rect -112 7746 -78 7780
rect -44 7746 -10 7780
rect 24 7746 58 7780
rect 92 7746 126 7780
rect 160 7746 194 7780
rect 228 7746 262 7780
rect 296 7746 330 7780
rect 364 7746 398 7780
rect 432 7746 466 7780
rect 500 7746 534 7780
rect 568 7746 602 7780
rect 636 7746 670 7780
rect 704 7746 738 7780
rect 772 7746 806 7780
rect 840 7746 874 7780
rect 908 7746 942 7780
rect 976 7746 1010 7780
rect 1044 7746 1078 7780
rect 1112 7746 1146 7780
rect 1180 7746 1214 7780
rect 1248 7746 1282 7780
rect 1316 7746 1350 7780
rect 1384 7746 1418 7780
rect 1452 7746 1486 7780
rect 1520 7746 1554 7780
rect 1588 7746 1622 7780
rect -1556 7638 -1522 7672
rect -1556 7570 -1522 7604
rect -1556 7502 -1522 7536
rect -1556 7434 -1522 7468
rect -1556 7366 -1522 7400
rect -1556 7298 -1522 7332
rect -1556 7230 -1522 7264
rect -1556 7162 -1522 7196
rect -1556 7094 -1522 7128
rect -1556 7026 -1522 7060
rect 1672 7638 1706 7672
rect 1672 7570 1706 7604
rect 1672 7502 1706 7536
rect 1672 7434 1706 7468
rect 1672 7366 1706 7400
rect 1672 7298 1706 7332
rect 1672 7230 1706 7264
rect 1672 7162 1706 7196
rect 1672 7094 1706 7128
rect 1672 7026 1706 7060
rect -1556 6958 -1522 6992
rect -1556 6890 -1522 6924
rect -1556 6822 -1522 6856
rect -1556 6754 -1522 6788
rect -1556 6686 -1522 6720
rect -1556 6618 -1522 6652
rect -1556 6550 -1522 6584
rect -1556 6482 -1522 6516
rect -1556 6414 -1522 6448
rect -1556 6346 -1522 6380
rect -1556 6278 -1522 6312
rect -1556 6210 -1522 6244
rect -1556 6142 -1522 6176
rect -1556 6074 -1522 6108
rect -1556 6006 -1522 6040
rect -1556 5938 -1522 5972
rect -1556 5870 -1522 5904
rect -1556 5802 -1522 5836
rect -1556 5734 -1522 5768
rect -1556 5666 -1522 5700
rect -1556 5598 -1522 5632
rect -1556 5530 -1522 5564
rect -1556 5462 -1522 5496
rect -1556 5394 -1522 5428
rect -1556 5326 -1522 5360
rect -1556 5258 -1522 5292
rect -1556 5190 -1522 5224
rect -1556 5122 -1522 5156
rect -1556 5054 -1522 5088
rect -1556 4986 -1522 5020
rect -1556 4918 -1522 4952
rect -1556 4850 -1522 4884
rect -1556 4782 -1522 4816
rect -1556 4714 -1522 4748
rect -1556 4646 -1522 4680
rect -1556 4578 -1522 4612
rect -1556 4510 -1522 4544
rect -1556 4442 -1522 4476
rect -1556 4374 -1522 4408
rect -1556 4306 -1522 4340
rect -1556 4238 -1522 4272
rect -1556 4170 -1522 4204
rect -1556 4102 -1522 4136
rect -1556 4034 -1522 4068
rect -1556 3966 -1522 4000
rect -1556 3898 -1522 3932
rect -1556 3830 -1522 3864
rect -1556 3762 -1522 3796
rect -1556 3694 -1522 3728
rect -1556 3626 -1522 3660
rect -1556 3558 -1522 3592
rect -1556 3490 -1522 3524
rect -1556 3422 -1522 3456
rect -1556 3354 -1522 3388
rect -1556 3286 -1522 3320
rect -1556 3218 -1522 3252
rect -1556 3150 -1522 3184
rect -1556 3082 -1522 3116
rect -1556 3014 -1522 3048
rect -1556 2946 -1522 2980
rect -1556 2878 -1522 2912
rect -1556 2810 -1522 2844
rect -1556 2742 -1522 2776
rect -1556 2674 -1522 2708
rect -1556 2606 -1522 2640
rect -1556 2538 -1522 2572
rect -1556 2470 -1522 2504
rect -1556 2402 -1522 2436
rect -1556 2334 -1522 2368
rect -1556 2266 -1522 2300
rect -1556 2198 -1522 2232
rect -1556 2130 -1522 2164
rect -1556 2062 -1522 2096
rect -1556 1994 -1522 2028
rect -1556 1926 -1522 1960
rect -1556 1858 -1522 1892
rect -1556 1790 -1522 1824
rect -1556 1722 -1522 1756
rect -1556 1654 -1522 1688
rect -1556 1586 -1522 1620
rect -1556 1518 -1522 1552
rect -1556 1450 -1522 1484
rect -1556 1382 -1522 1416
rect -1556 1314 -1522 1348
rect -1556 1246 -1522 1280
rect -1556 1178 -1522 1212
rect -1556 1110 -1522 1144
rect -1556 1042 -1522 1076
rect -1556 974 -1522 1008
rect -1556 906 -1522 940
rect -1556 838 -1522 872
rect -1556 770 -1522 804
rect -1556 702 -1522 736
rect -1556 634 -1522 668
rect -1556 566 -1522 600
rect -1556 498 -1522 532
rect -1556 430 -1522 464
rect -1556 362 -1522 396
rect -1556 294 -1522 328
rect -1556 226 -1522 260
rect -1556 158 -1522 192
rect -1556 90 -1522 124
rect -1556 22 -1522 56
rect -1556 -46 -1522 -12
rect -1556 -114 -1522 -80
rect -1556 -182 -1522 -148
rect -1556 -250 -1522 -216
rect -1556 -318 -1522 -284
rect -1556 -386 -1522 -352
rect -1556 -454 -1522 -420
rect -1556 -522 -1522 -488
rect -1556 -590 -1522 -556
rect -1556 -658 -1522 -624
rect -1556 -726 -1522 -692
rect -1556 -794 -1522 -760
rect -1556 -862 -1522 -828
rect -1556 -930 -1522 -896
rect -1556 -998 -1522 -964
rect 24 57 126 5939
rect 1672 6958 1706 6992
rect 1672 6890 1706 6924
rect 1672 6822 1706 6856
rect 1672 6754 1706 6788
rect 1672 6686 1706 6720
rect 1672 6618 1706 6652
rect 1672 6550 1706 6584
rect 1672 6482 1706 6516
rect 1672 6414 1706 6448
rect 1672 6346 1706 6380
rect 1672 6278 1706 6312
rect 1672 6210 1706 6244
rect 1672 6142 1706 6176
rect 1672 6074 1706 6108
rect 1672 6006 1706 6040
rect 1672 5938 1706 5972
rect 1672 5870 1706 5904
rect 1672 5802 1706 5836
rect 1672 5734 1706 5768
rect 1672 5666 1706 5700
rect 1672 5598 1706 5632
rect 1672 5530 1706 5564
rect 1672 5462 1706 5496
rect 1672 5394 1706 5428
rect 1672 5326 1706 5360
rect 1672 5258 1706 5292
rect 1672 5190 1706 5224
rect 1672 5122 1706 5156
rect 1672 5054 1706 5088
rect 1672 4986 1706 5020
rect 1672 4918 1706 4952
rect 1672 4850 1706 4884
rect 1672 4782 1706 4816
rect 1672 4714 1706 4748
rect 1672 4646 1706 4680
rect 1672 4578 1706 4612
rect 1672 4510 1706 4544
rect 1672 4442 1706 4476
rect 1672 4374 1706 4408
rect 1672 4306 1706 4340
rect 1672 4238 1706 4272
rect 1672 4170 1706 4204
rect 1672 4102 1706 4136
rect 1672 4034 1706 4068
rect 1672 3966 1706 4000
rect 1672 3898 1706 3932
rect 1672 3830 1706 3864
rect 1672 3762 1706 3796
rect 1672 3694 1706 3728
rect 1672 3626 1706 3660
rect 1672 3558 1706 3592
rect 1672 3490 1706 3524
rect 1672 3422 1706 3456
rect 1672 3354 1706 3388
rect 1672 3286 1706 3320
rect 1672 3218 1706 3252
rect 1672 3150 1706 3184
rect 1672 3082 1706 3116
rect 1672 3014 1706 3048
rect 1672 2946 1706 2980
rect 1672 2878 1706 2912
rect 1672 2810 1706 2844
rect 1672 2742 1706 2776
rect 1672 2674 1706 2708
rect 1672 2606 1706 2640
rect 1672 2538 1706 2572
rect 1672 2470 1706 2504
rect 1672 2402 1706 2436
rect 1672 2334 1706 2368
rect 1672 2266 1706 2300
rect 1672 2198 1706 2232
rect 1672 2130 1706 2164
rect 1672 2062 1706 2096
rect 1672 1994 1706 2028
rect 1672 1926 1706 1960
rect 1672 1858 1706 1892
rect 1672 1790 1706 1824
rect 1672 1722 1706 1756
rect 1672 1654 1706 1688
rect 1672 1586 1706 1620
rect 1672 1518 1706 1552
rect 1672 1450 1706 1484
rect 1672 1382 1706 1416
rect 1672 1314 1706 1348
rect 1672 1246 1706 1280
rect 1672 1178 1706 1212
rect 1672 1110 1706 1144
rect 1672 1042 1706 1076
rect 1672 974 1706 1008
rect 1672 906 1706 940
rect 1672 838 1706 872
rect 1672 770 1706 804
rect 1672 702 1706 736
rect 1672 634 1706 668
rect 1672 566 1706 600
rect 1672 498 1706 532
rect 1672 430 1706 464
rect 1672 362 1706 396
rect 1672 294 1706 328
rect 1672 226 1706 260
rect 1672 158 1706 192
rect 1672 90 1706 124
rect 1672 22 1706 56
rect 1672 -46 1706 -12
rect 1672 -114 1706 -80
rect 1672 -182 1706 -148
rect 1672 -250 1706 -216
rect 1672 -318 1706 -284
rect 1672 -386 1706 -352
rect 1672 -454 1706 -420
rect 1672 -522 1706 -488
rect 1672 -590 1706 -556
rect 1672 -658 1706 -624
rect 1672 -726 1706 -692
rect 1672 -794 1706 -760
rect 1672 -862 1706 -828
rect 1672 -930 1706 -896
rect 1672 -998 1706 -964
rect -1556 -1066 -1522 -1032
rect -1556 -1134 -1522 -1100
rect -1556 -1202 -1522 -1168
rect -1556 -1270 -1522 -1236
rect -1556 -1338 -1522 -1304
rect -1556 -1406 -1522 -1372
rect -1556 -1474 -1522 -1440
rect -1556 -1542 -1522 -1508
rect -1556 -1610 -1522 -1576
rect -1556 -1678 -1522 -1644
rect 1672 -1066 1706 -1032
rect 1672 -1134 1706 -1100
rect 1672 -1202 1706 -1168
rect 1672 -1270 1706 -1236
rect 1672 -1338 1706 -1304
rect 1672 -1406 1706 -1372
rect 1672 -1474 1706 -1440
rect 1672 -1542 1706 -1508
rect 1672 -1610 1706 -1576
rect 1672 -1678 1706 -1644
rect -1472 -1780 -1438 -1746
rect -1404 -1780 -1370 -1746
rect -1336 -1780 -1302 -1746
rect -1268 -1780 -1234 -1746
rect -1200 -1780 -1166 -1746
rect -1132 -1780 -1098 -1746
rect -1064 -1780 -1030 -1746
rect -996 -1780 -962 -1746
rect -928 -1780 -894 -1746
rect -860 -1780 -826 -1746
rect -792 -1780 -758 -1746
rect -724 -1780 -690 -1746
rect -656 -1780 -622 -1746
rect -588 -1780 -554 -1746
rect -520 -1780 -486 -1746
rect -452 -1780 -418 -1746
rect -384 -1780 -350 -1746
rect -316 -1780 -282 -1746
rect -248 -1780 -214 -1746
rect -180 -1780 -146 -1746
rect -112 -1780 -78 -1746
rect -44 -1780 -10 -1746
rect 24 -1780 58 -1746
rect 92 -1780 126 -1746
rect 160 -1780 194 -1746
rect 228 -1780 262 -1746
rect 296 -1780 330 -1746
rect 364 -1780 398 -1746
rect 432 -1780 466 -1746
rect 500 -1780 534 -1746
rect 568 -1780 602 -1746
rect 636 -1780 670 -1746
rect 704 -1780 738 -1746
rect 772 -1780 806 -1746
rect 840 -1780 874 -1746
rect 908 -1780 942 -1746
rect 976 -1780 1010 -1746
rect 1044 -1780 1078 -1746
rect 1112 -1780 1146 -1746
rect 1180 -1780 1214 -1746
rect 1248 -1780 1282 -1746
rect 1316 -1780 1350 -1746
rect 1384 -1780 1418 -1746
rect 1452 -1780 1486 -1746
rect 1520 -1780 1554 -1746
rect 1588 -1780 1622 -1746
<< mvnsubdiffcont >>
rect -520 6964 -486 6998
rect -452 6964 -418 6998
rect -384 6964 -350 6998
rect -316 6964 -282 6998
rect -248 6964 -214 6998
rect -180 6964 -146 6998
rect -112 6964 -78 6998
rect -44 6964 -10 6998
rect 24 6964 58 6998
rect 92 6964 126 6998
rect 160 6964 194 6998
rect 228 6964 262 6998
rect 296 6964 330 6998
rect 364 6964 398 6998
rect 432 6964 466 6998
rect 500 6964 534 6998
rect 568 6964 602 6998
rect 636 6964 670 6998
rect -774 6822 -740 6856
rect 890 6822 924 6856
rect -774 6754 -740 6788
rect -774 6686 -740 6720
rect -774 6618 -740 6652
rect -774 6550 -740 6584
rect -774 6482 -740 6516
rect -774 6414 -740 6448
rect -774 6346 -740 6380
rect -774 6278 -740 6312
rect -774 6210 -740 6244
rect -774 6142 -740 6176
rect -774 6074 -740 6108
rect -774 6006 -740 6040
rect 890 6754 924 6788
rect 890 6686 924 6720
rect 890 6618 924 6652
rect 890 6550 924 6584
rect 890 6482 924 6516
rect 890 6414 924 6448
rect 890 6346 924 6380
rect 890 6278 924 6312
rect 890 6210 924 6244
rect 890 6142 924 6176
rect 890 6074 924 6108
rect 890 6006 924 6040
rect -774 5938 -740 5972
rect -774 5870 -740 5904
rect -774 5802 -740 5836
rect -774 5734 -740 5768
rect -774 5666 -740 5700
rect -774 5598 -740 5632
rect -774 5530 -740 5564
rect -774 5462 -740 5496
rect -774 5394 -740 5428
rect -774 5326 -740 5360
rect -774 5258 -740 5292
rect -774 5190 -740 5224
rect -774 5122 -740 5156
rect -774 5054 -740 5088
rect -774 4986 -740 5020
rect -774 4918 -740 4952
rect -774 4850 -740 4884
rect -774 4782 -740 4816
rect -774 4714 -740 4748
rect -774 4646 -740 4680
rect -774 4578 -740 4612
rect -774 4510 -740 4544
rect -774 4442 -740 4476
rect -774 4374 -740 4408
rect -774 4306 -740 4340
rect -774 4238 -740 4272
rect -774 4170 -740 4204
rect -774 4102 -740 4136
rect -774 4034 -740 4068
rect -774 3966 -740 4000
rect -774 3898 -740 3932
rect -774 3830 -740 3864
rect -774 3762 -740 3796
rect -774 3694 -740 3728
rect -774 3626 -740 3660
rect -774 3558 -740 3592
rect -774 3490 -740 3524
rect -774 3422 -740 3456
rect -774 3354 -740 3388
rect -774 3286 -740 3320
rect -774 3218 -740 3252
rect -774 3150 -740 3184
rect -774 3082 -740 3116
rect -774 3014 -740 3048
rect -774 2946 -740 2980
rect -774 2878 -740 2912
rect -774 2810 -740 2844
rect -774 2742 -740 2776
rect -774 2674 -740 2708
rect -774 2606 -740 2640
rect -774 2538 -740 2572
rect -774 2470 -740 2504
rect -774 2402 -740 2436
rect -774 2334 -740 2368
rect -774 2266 -740 2300
rect -774 2198 -740 2232
rect -774 2130 -740 2164
rect -774 2062 -740 2096
rect -774 1994 -740 2028
rect -774 1926 -740 1960
rect -774 1858 -740 1892
rect -774 1790 -740 1824
rect -774 1722 -740 1756
rect -774 1654 -740 1688
rect -774 1586 -740 1620
rect -774 1518 -740 1552
rect -774 1450 -740 1484
rect -774 1382 -740 1416
rect -774 1314 -740 1348
rect -774 1246 -740 1280
rect -774 1178 -740 1212
rect -774 1110 -740 1144
rect -774 1042 -740 1076
rect -774 974 -740 1008
rect -774 906 -740 940
rect -774 838 -740 872
rect -774 770 -740 804
rect -774 702 -740 736
rect -774 634 -740 668
rect -774 566 -740 600
rect -774 498 -740 532
rect -774 430 -740 464
rect -774 362 -740 396
rect -774 294 -740 328
rect -774 226 -740 260
rect -774 158 -740 192
rect -774 90 -740 124
rect -774 22 -740 56
rect 890 5938 924 5972
rect 890 5870 924 5904
rect 890 5802 924 5836
rect 890 5734 924 5768
rect 890 5666 924 5700
rect 890 5598 924 5632
rect 890 5530 924 5564
rect 890 5462 924 5496
rect 890 5394 924 5428
rect 890 5326 924 5360
rect 890 5258 924 5292
rect 890 5190 924 5224
rect 890 5122 924 5156
rect 890 5054 924 5088
rect 890 4986 924 5020
rect 890 4918 924 4952
rect 890 4850 924 4884
rect 890 4782 924 4816
rect 890 4714 924 4748
rect 890 4646 924 4680
rect 890 4578 924 4612
rect 890 4510 924 4544
rect 890 4442 924 4476
rect 890 4374 924 4408
rect 890 4306 924 4340
rect 890 4238 924 4272
rect 890 4170 924 4204
rect 890 4102 924 4136
rect 890 4034 924 4068
rect 890 3966 924 4000
rect 890 3898 924 3932
rect 890 3830 924 3864
rect 890 3762 924 3796
rect 890 3694 924 3728
rect 890 3626 924 3660
rect 890 3558 924 3592
rect 890 3490 924 3524
rect 890 3422 924 3456
rect 890 3354 924 3388
rect 890 3286 924 3320
rect 890 3218 924 3252
rect 890 3150 924 3184
rect 890 3082 924 3116
rect 890 3014 924 3048
rect 890 2946 924 2980
rect 890 2878 924 2912
rect 890 2810 924 2844
rect 890 2742 924 2776
rect 890 2674 924 2708
rect 890 2606 924 2640
rect 890 2538 924 2572
rect 890 2470 924 2504
rect 890 2402 924 2436
rect 890 2334 924 2368
rect 890 2266 924 2300
rect 890 2198 924 2232
rect 890 2130 924 2164
rect 890 2062 924 2096
rect 890 1994 924 2028
rect 890 1926 924 1960
rect 890 1858 924 1892
rect 890 1790 924 1824
rect 890 1722 924 1756
rect 890 1654 924 1688
rect 890 1586 924 1620
rect 890 1518 924 1552
rect 890 1450 924 1484
rect 890 1382 924 1416
rect 890 1314 924 1348
rect 890 1246 924 1280
rect 890 1178 924 1212
rect 890 1110 924 1144
rect 890 1042 924 1076
rect 890 974 924 1008
rect 890 906 924 940
rect 890 838 924 872
rect 890 770 924 804
rect 890 702 924 736
rect 890 634 924 668
rect 890 566 924 600
rect 890 498 924 532
rect 890 430 924 464
rect 890 362 924 396
rect 890 294 924 328
rect 890 226 924 260
rect 890 158 924 192
rect 890 90 924 124
rect 890 22 924 56
rect -774 -46 -740 -12
rect -774 -114 -740 -80
rect -774 -182 -740 -148
rect -774 -250 -740 -216
rect -774 -318 -740 -284
rect -774 -386 -740 -352
rect -774 -454 -740 -420
rect -774 -522 -740 -488
rect -774 -590 -740 -556
rect -774 -658 -740 -624
rect -774 -726 -740 -692
rect -774 -794 -740 -760
rect 890 -46 924 -12
rect 890 -114 924 -80
rect 890 -182 924 -148
rect 890 -250 924 -216
rect 890 -318 924 -284
rect 890 -386 924 -352
rect 890 -454 924 -420
rect 890 -522 924 -488
rect 890 -590 924 -556
rect 890 -658 924 -624
rect 890 -726 924 -692
rect 890 -794 924 -760
rect -774 -862 -740 -828
rect -774 -930 -740 -896
rect 890 -862 924 -828
rect 890 -930 924 -896
rect -774 -998 -740 -964
rect -520 -998 -486 -964
rect -452 -998 -418 -964
rect -384 -998 -350 -964
rect -316 -998 -282 -964
rect -248 -998 -214 -964
rect -180 -998 -146 -964
rect -112 -998 -78 -964
rect -44 -998 -10 -964
rect 24 -998 58 -964
rect 92 -998 126 -964
rect 160 -998 194 -964
rect 228 -998 262 -964
rect 296 -998 330 -964
rect 364 -998 398 -964
rect 432 -998 466 -964
rect 500 -998 534 -964
rect 568 -998 602 -964
rect 636 -998 670 -964
rect 890 -998 924 -964
<< poly >>
rect -600 6300 750 6800
rect -600 6000 -200 6300
rect 350 6000 750 6300
rect -300 0 -200 6000
rect 350 0 450 6000
rect -600 -300 -200 0
rect 350 -300 750 0
rect -600 -459 750 -300
rect -600 -493 -130 -459
rect -96 -493 -56 -459
rect -22 -493 18 -459
rect 52 -493 92 -459
rect 126 -493 166 -459
rect 200 -493 240 -459
rect 274 -493 750 -459
rect -600 -533 750 -493
rect -600 -567 -130 -533
rect -96 -567 -56 -533
rect -22 -567 18 -533
rect 52 -567 92 -533
rect 126 -567 166 -533
rect 200 -567 240 -533
rect 274 -567 750 -533
rect -600 -607 750 -567
rect -600 -641 -130 -607
rect -96 -641 -56 -607
rect -22 -641 18 -607
rect 52 -641 92 -607
rect 126 -641 166 -607
rect 200 -641 240 -607
rect 274 -641 750 -607
rect -600 -800 750 -641
<< polycont >>
rect -130 -493 -96 -459
rect -56 -493 -22 -459
rect 18 -493 52 -459
rect 92 -493 126 -459
rect 166 -493 200 -459
rect 240 -493 274 -459
rect -130 -567 -96 -533
rect -56 -567 -22 -533
rect 18 -567 52 -533
rect 92 -567 126 -533
rect 166 -567 200 -533
rect 240 -567 274 -533
rect -130 -641 -96 -607
rect -56 -641 -22 -607
rect 18 -641 52 -607
rect 92 -641 126 -607
rect 166 -641 200 -607
rect 240 -641 274 -607
<< locali >>
rect -1580 7780 1730 7804
rect -1580 7746 -1472 7780
rect -1420 7746 -1404 7780
rect -1348 7746 -1336 7780
rect -1276 7746 -1268 7780
rect -1204 7746 -1200 7780
rect -1098 7746 -1094 7780
rect -1030 7746 -1022 7780
rect -962 7746 -950 7780
rect -894 7746 -878 7780
rect -826 7746 -806 7780
rect -758 7746 -734 7780
rect -690 7746 -662 7780
rect -622 7746 -590 7780
rect -554 7746 -520 7780
rect -484 7746 -452 7780
rect -412 7746 -384 7780
rect -340 7746 -316 7780
rect -268 7746 -248 7780
rect -196 7746 -180 7780
rect -124 7746 -112 7780
rect -52 7746 -44 7780
rect 20 7746 24 7780
rect 126 7746 130 7780
rect 194 7746 202 7780
rect 262 7746 274 7780
rect 330 7746 346 7780
rect 398 7746 418 7780
rect 466 7746 490 7780
rect 534 7746 562 7780
rect 602 7746 634 7780
rect 670 7746 704 7780
rect 740 7746 772 7780
rect 812 7746 840 7780
rect 884 7746 908 7780
rect 956 7746 976 7780
rect 1028 7746 1044 7780
rect 1100 7746 1112 7780
rect 1172 7746 1180 7780
rect 1244 7746 1248 7780
rect 1350 7746 1354 7780
rect 1418 7746 1426 7780
rect 1486 7746 1498 7780
rect 1554 7746 1570 7780
rect 1622 7746 1730 7780
rect -1580 7722 1730 7746
rect -1580 7672 -1498 7722
rect -1580 7627 -1556 7672
rect -1522 7627 -1498 7672
rect -1580 7604 -1498 7627
rect -1580 7555 -1556 7604
rect -1522 7555 -1498 7604
rect -1580 7536 -1498 7555
rect -1580 7483 -1556 7536
rect -1522 7483 -1498 7536
rect -1580 7468 -1498 7483
rect -1580 7411 -1556 7468
rect -1522 7411 -1498 7468
rect -1580 7400 -1498 7411
rect -1580 7339 -1556 7400
rect -1522 7339 -1498 7400
rect -1580 7332 -1498 7339
rect -1580 7267 -1556 7332
rect -1522 7267 -1498 7332
rect -1580 7264 -1498 7267
rect -1580 7230 -1556 7264
rect -1522 7230 -1498 7264
rect -1580 7229 -1498 7230
rect -1580 7162 -1556 7229
rect -1522 7162 -1498 7229
rect -1580 7157 -1498 7162
rect -1580 7094 -1556 7157
rect -1522 7094 -1498 7157
rect -1580 7085 -1498 7094
rect -1580 7026 -1556 7085
rect -1522 7026 -1498 7085
rect -1580 7013 -1498 7026
rect 1648 7672 1730 7722
rect 1648 7627 1672 7672
rect 1706 7627 1730 7672
rect 1648 7604 1730 7627
rect 1648 7555 1672 7604
rect 1706 7555 1730 7604
rect 1648 7536 1730 7555
rect 1648 7483 1672 7536
rect 1706 7483 1730 7536
rect 1648 7468 1730 7483
rect 1648 7411 1672 7468
rect 1706 7411 1730 7468
rect 1648 7400 1730 7411
rect 1648 7339 1672 7400
rect 1706 7339 1730 7400
rect 1648 7332 1730 7339
rect 1648 7267 1672 7332
rect 1706 7267 1730 7332
rect 1648 7264 1730 7267
rect 1648 7230 1672 7264
rect 1706 7230 1730 7264
rect 1648 7229 1730 7230
rect 1648 7162 1672 7229
rect 1706 7162 1730 7229
rect 1648 7157 1730 7162
rect 1648 7094 1672 7157
rect 1706 7094 1730 7157
rect 1648 7085 1730 7094
rect 1648 7026 1672 7085
rect 1706 7026 1730 7085
rect -1580 6958 -1556 7013
rect -1522 6958 -1498 7013
rect -1580 6941 -1498 6958
rect -1580 6890 -1556 6941
rect -1522 6890 -1498 6941
rect -1580 6869 -1498 6890
rect -1580 6822 -1556 6869
rect -1522 6822 -1498 6869
rect -1580 6797 -1498 6822
rect -1580 6754 -1556 6797
rect -1522 6754 -1498 6797
rect -1580 6725 -1498 6754
rect -1580 6686 -1556 6725
rect -1522 6686 -1498 6725
rect -1580 6653 -1498 6686
rect -1580 6618 -1556 6653
rect -1522 6618 -1498 6653
rect -1580 6584 -1498 6618
rect -1580 6547 -1556 6584
rect -1522 6547 -1498 6584
rect -1580 6516 -1498 6547
rect -1580 6475 -1556 6516
rect -1522 6475 -1498 6516
rect -1580 6448 -1498 6475
rect -1580 6403 -1556 6448
rect -1522 6403 -1498 6448
rect -1580 6380 -1498 6403
rect -1580 6331 -1556 6380
rect -1522 6331 -1498 6380
rect -1580 6312 -1498 6331
rect -1580 6259 -1556 6312
rect -1522 6259 -1498 6312
rect -1580 6244 -1498 6259
rect -1580 6187 -1556 6244
rect -1522 6187 -1498 6244
rect -1580 6176 -1498 6187
rect -1580 6115 -1556 6176
rect -1522 6115 -1498 6176
rect -1580 6108 -1498 6115
rect -1580 6043 -1556 6108
rect -1522 6043 -1498 6108
rect -1580 6040 -1498 6043
rect -1580 6006 -1556 6040
rect -1522 6006 -1498 6040
rect -1580 6005 -1498 6006
rect -1580 5938 -1556 6005
rect -1522 5938 -1498 6005
rect -1580 5933 -1498 5938
rect -1580 5870 -1556 5933
rect -1522 5870 -1498 5933
rect -1580 5861 -1498 5870
rect -1580 5802 -1556 5861
rect -1522 5802 -1498 5861
rect -1580 5789 -1498 5802
rect -1580 5734 -1556 5789
rect -1522 5734 -1498 5789
rect -1580 5717 -1498 5734
rect -1580 5666 -1556 5717
rect -1522 5666 -1498 5717
rect -1580 5645 -1498 5666
rect -1580 5598 -1556 5645
rect -1522 5598 -1498 5645
rect -1580 5573 -1498 5598
rect -1580 5530 -1556 5573
rect -1522 5530 -1498 5573
rect -1580 5501 -1498 5530
rect -1580 5462 -1556 5501
rect -1522 5462 -1498 5501
rect -1580 5429 -1498 5462
rect -1580 5394 -1556 5429
rect -1522 5394 -1498 5429
rect -1580 5360 -1498 5394
rect -1580 5323 -1556 5360
rect -1522 5323 -1498 5360
rect -1580 5292 -1498 5323
rect -1580 5251 -1556 5292
rect -1522 5251 -1498 5292
rect -1580 5224 -1498 5251
rect -1580 5179 -1556 5224
rect -1522 5179 -1498 5224
rect -1580 5156 -1498 5179
rect -1580 5107 -1556 5156
rect -1522 5107 -1498 5156
rect -1580 5088 -1498 5107
rect -1580 5035 -1556 5088
rect -1522 5035 -1498 5088
rect -1580 5020 -1498 5035
rect -1580 4963 -1556 5020
rect -1522 4963 -1498 5020
rect -1580 4952 -1498 4963
rect -1580 4891 -1556 4952
rect -1522 4891 -1498 4952
rect -1580 4884 -1498 4891
rect -1580 4819 -1556 4884
rect -1522 4819 -1498 4884
rect -1580 4816 -1498 4819
rect -1580 4782 -1556 4816
rect -1522 4782 -1498 4816
rect -1580 4781 -1498 4782
rect -1580 4714 -1556 4781
rect -1522 4714 -1498 4781
rect -1580 4709 -1498 4714
rect -1580 4646 -1556 4709
rect -1522 4646 -1498 4709
rect -1580 4637 -1498 4646
rect -1580 4578 -1556 4637
rect -1522 4578 -1498 4637
rect -1580 4565 -1498 4578
rect -1580 4510 -1556 4565
rect -1522 4510 -1498 4565
rect -1580 4493 -1498 4510
rect -1580 4442 -1556 4493
rect -1522 4442 -1498 4493
rect -1580 4421 -1498 4442
rect -1580 4374 -1556 4421
rect -1522 4374 -1498 4421
rect -1580 4349 -1498 4374
rect -1580 4306 -1556 4349
rect -1522 4306 -1498 4349
rect -1580 4277 -1498 4306
rect -1580 4238 -1556 4277
rect -1522 4238 -1498 4277
rect -1580 4205 -1498 4238
rect -1580 4170 -1556 4205
rect -1522 4170 -1498 4205
rect -1580 4136 -1498 4170
rect -1580 4099 -1556 4136
rect -1522 4099 -1498 4136
rect -1580 4068 -1498 4099
rect -1580 4027 -1556 4068
rect -1522 4027 -1498 4068
rect -1580 4000 -1498 4027
rect -1580 3955 -1556 4000
rect -1522 3955 -1498 4000
rect -1580 3932 -1498 3955
rect -1580 3883 -1556 3932
rect -1522 3883 -1498 3932
rect -1580 3864 -1498 3883
rect -1580 3811 -1556 3864
rect -1522 3811 -1498 3864
rect -1580 3796 -1498 3811
rect -1580 3739 -1556 3796
rect -1522 3739 -1498 3796
rect -1580 3728 -1498 3739
rect -1580 3667 -1556 3728
rect -1522 3667 -1498 3728
rect -1580 3660 -1498 3667
rect -1580 3595 -1556 3660
rect -1522 3595 -1498 3660
rect -1580 3592 -1498 3595
rect -1580 3558 -1556 3592
rect -1522 3558 -1498 3592
rect -1580 3557 -1498 3558
rect -1580 3490 -1556 3557
rect -1522 3490 -1498 3557
rect -1580 3485 -1498 3490
rect -1580 3422 -1556 3485
rect -1522 3422 -1498 3485
rect -1580 3413 -1498 3422
rect -1580 3354 -1556 3413
rect -1522 3354 -1498 3413
rect -1580 3341 -1498 3354
rect -1580 3286 -1556 3341
rect -1522 3286 -1498 3341
rect -1580 3269 -1498 3286
rect -1580 3218 -1556 3269
rect -1522 3218 -1498 3269
rect -1580 3197 -1498 3218
rect -1580 3150 -1556 3197
rect -1522 3150 -1498 3197
rect -1580 3125 -1498 3150
rect -1580 3082 -1556 3125
rect -1522 3082 -1498 3125
rect -1580 3053 -1498 3082
rect -1580 3014 -1556 3053
rect -1522 3014 -1498 3053
rect -1580 2981 -1498 3014
rect -1580 2946 -1556 2981
rect -1522 2946 -1498 2981
rect -1580 2912 -1498 2946
rect -1580 2875 -1556 2912
rect -1522 2875 -1498 2912
rect -1580 2844 -1498 2875
rect -1580 2803 -1556 2844
rect -1522 2803 -1498 2844
rect -1580 2776 -1498 2803
rect -1580 2731 -1556 2776
rect -1522 2731 -1498 2776
rect -1580 2708 -1498 2731
rect -1580 2659 -1556 2708
rect -1522 2659 -1498 2708
rect -1580 2640 -1498 2659
rect -1580 2587 -1556 2640
rect -1522 2587 -1498 2640
rect -1580 2572 -1498 2587
rect -1580 2515 -1556 2572
rect -1522 2515 -1498 2572
rect -1580 2504 -1498 2515
rect -1580 2443 -1556 2504
rect -1522 2443 -1498 2504
rect -1580 2436 -1498 2443
rect -1580 2371 -1556 2436
rect -1522 2371 -1498 2436
rect -1580 2368 -1498 2371
rect -1580 2334 -1556 2368
rect -1522 2334 -1498 2368
rect -1580 2333 -1498 2334
rect -1580 2266 -1556 2333
rect -1522 2266 -1498 2333
rect -1580 2261 -1498 2266
rect -1580 2198 -1556 2261
rect -1522 2198 -1498 2261
rect -1580 2189 -1498 2198
rect -1580 2130 -1556 2189
rect -1522 2130 -1498 2189
rect -1580 2117 -1498 2130
rect -1580 2062 -1556 2117
rect -1522 2062 -1498 2117
rect -1580 2045 -1498 2062
rect -1580 1994 -1556 2045
rect -1522 1994 -1498 2045
rect -1580 1973 -1498 1994
rect -1580 1926 -1556 1973
rect -1522 1926 -1498 1973
rect -1580 1901 -1498 1926
rect -1580 1858 -1556 1901
rect -1522 1858 -1498 1901
rect -1580 1829 -1498 1858
rect -1580 1790 -1556 1829
rect -1522 1790 -1498 1829
rect -1580 1757 -1498 1790
rect -1580 1722 -1556 1757
rect -1522 1722 -1498 1757
rect -1580 1688 -1498 1722
rect -1580 1651 -1556 1688
rect -1522 1651 -1498 1688
rect -1580 1620 -1498 1651
rect -1580 1579 -1556 1620
rect -1522 1579 -1498 1620
rect -1580 1552 -1498 1579
rect -1580 1507 -1556 1552
rect -1522 1507 -1498 1552
rect -1580 1484 -1498 1507
rect -1580 1435 -1556 1484
rect -1522 1435 -1498 1484
rect -1580 1416 -1498 1435
rect -1580 1363 -1556 1416
rect -1522 1363 -1498 1416
rect -1580 1348 -1498 1363
rect -1580 1291 -1556 1348
rect -1522 1291 -1498 1348
rect -1580 1280 -1498 1291
rect -1580 1219 -1556 1280
rect -1522 1219 -1498 1280
rect -1580 1212 -1498 1219
rect -1580 1147 -1556 1212
rect -1522 1147 -1498 1212
rect -1580 1144 -1498 1147
rect -1580 1110 -1556 1144
rect -1522 1110 -1498 1144
rect -1580 1109 -1498 1110
rect -1580 1042 -1556 1109
rect -1522 1042 -1498 1109
rect -1580 1037 -1498 1042
rect -1580 974 -1556 1037
rect -1522 974 -1498 1037
rect -1580 965 -1498 974
rect -1580 906 -1556 965
rect -1522 906 -1498 965
rect -1580 893 -1498 906
rect -1580 838 -1556 893
rect -1522 838 -1498 893
rect -1580 821 -1498 838
rect -1580 770 -1556 821
rect -1522 770 -1498 821
rect -1580 749 -1498 770
rect -1580 702 -1556 749
rect -1522 702 -1498 749
rect -1580 677 -1498 702
rect -1580 634 -1556 677
rect -1522 634 -1498 677
rect -1580 605 -1498 634
rect -1580 566 -1556 605
rect -1522 566 -1498 605
rect -1580 533 -1498 566
rect -1580 498 -1556 533
rect -1522 498 -1498 533
rect -1580 464 -1498 498
rect -1580 427 -1556 464
rect -1522 427 -1498 464
rect -1580 396 -1498 427
rect -1580 355 -1556 396
rect -1522 355 -1498 396
rect -1580 328 -1498 355
rect -1580 283 -1556 328
rect -1522 283 -1498 328
rect -1580 260 -1498 283
rect -1580 211 -1556 260
rect -1522 211 -1498 260
rect -1580 192 -1498 211
rect -1580 139 -1556 192
rect -1522 139 -1498 192
rect -1580 124 -1498 139
rect -1580 67 -1556 124
rect -1522 67 -1498 124
rect -1580 56 -1498 67
rect -1580 -5 -1556 56
rect -1522 -5 -1498 56
rect -1580 -12 -1498 -5
rect -1580 -77 -1556 -12
rect -1522 -77 -1498 -12
rect -1580 -80 -1498 -77
rect -1580 -114 -1556 -80
rect -1522 -114 -1498 -80
rect -1580 -115 -1498 -114
rect -1580 -182 -1556 -115
rect -1522 -182 -1498 -115
rect -1580 -187 -1498 -182
rect -1580 -250 -1556 -187
rect -1522 -250 -1498 -187
rect -1580 -259 -1498 -250
rect -1580 -318 -1556 -259
rect -1522 -318 -1498 -259
rect -1580 -331 -1498 -318
rect -1580 -386 -1556 -331
rect -1522 -386 -1498 -331
rect -1580 -403 -1498 -386
rect -1580 -454 -1556 -403
rect -1522 -454 -1498 -403
rect -1580 -475 -1498 -454
rect -1580 -522 -1556 -475
rect -1522 -522 -1498 -475
rect -1580 -547 -1498 -522
rect -1580 -590 -1556 -547
rect -1522 -590 -1498 -547
rect -1580 -619 -1498 -590
rect -1580 -658 -1556 -619
rect -1522 -658 -1498 -619
rect -1580 -691 -1498 -658
rect -1580 -726 -1556 -691
rect -1522 -726 -1498 -691
rect -1580 -760 -1498 -726
rect -1580 -797 -1556 -760
rect -1522 -797 -1498 -760
rect -1580 -828 -1498 -797
rect -1580 -869 -1556 -828
rect -1522 -869 -1498 -828
rect -1580 -896 -1498 -869
rect -1580 -941 -1556 -896
rect -1522 -941 -1498 -896
rect -1580 -964 -1498 -941
rect -1580 -1013 -1556 -964
rect -1522 -1013 -1498 -964
rect -1580 -1032 -1498 -1013
rect -798 6998 948 7022
rect -798 6856 -554 6998
rect -798 6822 -774 6856
rect -740 6822 -554 6856
rect -798 6820 -554 6822
rect 704 6856 948 6998
rect 704 6822 890 6856
rect 924 6822 948 6856
rect 704 6820 948 6822
rect -798 6788 948 6820
rect -798 6754 -774 6788
rect -740 6757 890 6788
rect -740 6754 -716 6757
rect -798 6720 -716 6754
rect -798 6686 -774 6720
rect -740 6686 -716 6720
rect -798 6652 -716 6686
rect -798 6616 -774 6652
rect -740 6616 -716 6652
rect -798 6584 -716 6616
rect -798 6544 -774 6584
rect -740 6544 -716 6584
rect -798 6516 -716 6544
rect -798 6472 -774 6516
rect -740 6472 -716 6516
rect -798 6448 -716 6472
rect -798 6400 -774 6448
rect -740 6400 -716 6448
rect -798 6380 -716 6400
rect -798 6328 -774 6380
rect -740 6328 -716 6380
rect -798 6312 -716 6328
rect -798 6256 -774 6312
rect -740 6256 -716 6312
rect -798 6244 -716 6256
rect -798 6184 -774 6244
rect -740 6184 -716 6244
rect -798 6176 -716 6184
rect -798 6112 -774 6176
rect -740 6112 -716 6176
rect 866 6754 890 6757
rect 924 6754 948 6788
rect 866 6720 948 6754
rect 866 6686 890 6720
rect 924 6686 948 6720
rect 866 6652 948 6686
rect 866 6616 890 6652
rect 924 6616 948 6652
rect 866 6584 948 6616
rect 866 6544 890 6584
rect 924 6544 948 6584
rect 866 6516 948 6544
rect 866 6472 890 6516
rect 924 6472 948 6516
rect 866 6448 948 6472
rect 866 6400 890 6448
rect 924 6400 948 6448
rect 866 6380 948 6400
rect 866 6328 890 6380
rect 924 6328 948 6380
rect 866 6312 948 6328
rect 866 6256 890 6312
rect 924 6256 948 6312
rect 866 6244 948 6256
rect 866 6184 890 6244
rect 924 6184 948 6244
rect 866 6176 948 6184
rect -798 6108 -716 6112
rect -798 6006 -774 6108
rect -740 6006 -716 6108
rect -798 6002 -716 6006
rect -798 5938 -774 6002
rect -740 5938 -716 6002
rect -798 5930 -716 5938
rect -798 5870 -774 5930
rect -740 5870 -716 5930
rect -798 5858 -716 5870
rect -798 5802 -774 5858
rect -740 5802 -716 5858
rect -798 5786 -716 5802
rect -798 5734 -774 5786
rect -740 5734 -716 5786
rect -798 5714 -716 5734
rect -798 5666 -774 5714
rect -740 5666 -716 5714
rect -798 5642 -716 5666
rect -798 5598 -774 5642
rect -740 5598 -716 5642
rect -798 5570 -716 5598
rect -798 5530 -774 5570
rect -740 5530 -716 5570
rect -798 5498 -716 5530
rect -798 5462 -774 5498
rect -740 5462 -716 5498
rect -798 5428 -716 5462
rect -798 5392 -774 5428
rect -740 5392 -716 5428
rect -798 5360 -716 5392
rect -798 5320 -774 5360
rect -740 5320 -716 5360
rect -798 5292 -716 5320
rect -798 5248 -774 5292
rect -740 5248 -716 5292
rect -798 5224 -716 5248
rect -798 5176 -774 5224
rect -740 5176 -716 5224
rect -798 5156 -716 5176
rect -798 5104 -774 5156
rect -740 5104 -716 5156
rect -798 5088 -716 5104
rect -798 5032 -774 5088
rect -740 5032 -716 5088
rect -798 5020 -716 5032
rect -798 4960 -774 5020
rect -740 4960 -716 5020
rect -798 4952 -716 4960
rect -798 4888 -774 4952
rect -740 4888 -716 4952
rect -798 4884 -716 4888
rect -798 4782 -774 4884
rect -740 4782 -716 4884
rect -798 4778 -716 4782
rect -798 4714 -774 4778
rect -740 4714 -716 4778
rect -798 4706 -716 4714
rect -798 4646 -774 4706
rect -740 4646 -716 4706
rect -798 4634 -716 4646
rect -798 4578 -774 4634
rect -740 4578 -716 4634
rect -798 4562 -716 4578
rect -798 4510 -774 4562
rect -740 4510 -716 4562
rect -798 4490 -716 4510
rect -798 4442 -774 4490
rect -740 4442 -716 4490
rect -798 4418 -716 4442
rect -798 4374 -774 4418
rect -740 4374 -716 4418
rect -798 4346 -716 4374
rect -798 4306 -774 4346
rect -740 4306 -716 4346
rect -798 4274 -716 4306
rect -798 4238 -774 4274
rect -740 4238 -716 4274
rect -798 4204 -716 4238
rect -798 4168 -774 4204
rect -740 4168 -716 4204
rect -798 4136 -716 4168
rect -798 4096 -774 4136
rect -740 4096 -716 4136
rect -798 4068 -716 4096
rect -798 4024 -774 4068
rect -740 4024 -716 4068
rect -798 4000 -716 4024
rect -798 3952 -774 4000
rect -740 3952 -716 4000
rect -798 3932 -716 3952
rect -798 3880 -774 3932
rect -740 3880 -716 3932
rect -798 3864 -716 3880
rect -798 3808 -774 3864
rect -740 3808 -716 3864
rect -798 3796 -716 3808
rect -798 3736 -774 3796
rect -740 3736 -716 3796
rect -798 3728 -716 3736
rect -798 3664 -774 3728
rect -740 3664 -716 3728
rect -798 3660 -716 3664
rect -798 3558 -774 3660
rect -740 3558 -716 3660
rect -798 3554 -716 3558
rect -798 3490 -774 3554
rect -740 3490 -716 3554
rect -798 3482 -716 3490
rect -798 3422 -774 3482
rect -740 3422 -716 3482
rect -798 3410 -716 3422
rect -798 3354 -774 3410
rect -740 3354 -716 3410
rect -798 3338 -716 3354
rect -798 3286 -774 3338
rect -740 3286 -716 3338
rect -798 3266 -716 3286
rect -798 3218 -774 3266
rect -740 3218 -716 3266
rect -798 3194 -716 3218
rect -798 3150 -774 3194
rect -740 3150 -716 3194
rect -798 3122 -716 3150
rect -798 3082 -774 3122
rect -740 3082 -716 3122
rect -798 3050 -716 3082
rect -798 3014 -774 3050
rect -740 3014 -716 3050
rect -798 2980 -716 3014
rect -798 2944 -774 2980
rect -740 2944 -716 2980
rect -798 2912 -716 2944
rect -798 2872 -774 2912
rect -740 2872 -716 2912
rect -798 2844 -716 2872
rect -798 2800 -774 2844
rect -740 2800 -716 2844
rect -798 2776 -716 2800
rect -798 2728 -774 2776
rect -740 2728 -716 2776
rect -798 2708 -716 2728
rect -798 2656 -774 2708
rect -740 2656 -716 2708
rect -798 2640 -716 2656
rect -798 2584 -774 2640
rect -740 2584 -716 2640
rect -798 2572 -716 2584
rect -798 2512 -774 2572
rect -740 2512 -716 2572
rect -798 2504 -716 2512
rect -798 2440 -774 2504
rect -740 2440 -716 2504
rect -798 2436 -716 2440
rect -798 2334 -774 2436
rect -740 2334 -716 2436
rect -798 2330 -716 2334
rect -798 2266 -774 2330
rect -740 2266 -716 2330
rect -798 2258 -716 2266
rect -798 2198 -774 2258
rect -740 2198 -716 2258
rect -798 2186 -716 2198
rect -798 2130 -774 2186
rect -740 2130 -716 2186
rect -798 2114 -716 2130
rect -798 2062 -774 2114
rect -740 2062 -716 2114
rect -798 2042 -716 2062
rect -798 1994 -774 2042
rect -740 1994 -716 2042
rect -798 1970 -716 1994
rect -798 1926 -774 1970
rect -740 1926 -716 1970
rect -798 1898 -716 1926
rect -798 1858 -774 1898
rect -740 1858 -716 1898
rect -798 1826 -716 1858
rect -798 1790 -774 1826
rect -740 1790 -716 1826
rect -798 1756 -716 1790
rect -798 1720 -774 1756
rect -740 1720 -716 1756
rect -798 1688 -716 1720
rect -798 1648 -774 1688
rect -740 1648 -716 1688
rect -798 1620 -716 1648
rect -798 1576 -774 1620
rect -740 1576 -716 1620
rect -798 1552 -716 1576
rect -798 1504 -774 1552
rect -740 1504 -716 1552
rect -798 1484 -716 1504
rect -798 1432 -774 1484
rect -740 1432 -716 1484
rect -798 1416 -716 1432
rect -798 1360 -774 1416
rect -740 1360 -716 1416
rect -798 1348 -716 1360
rect -798 1288 -774 1348
rect -740 1288 -716 1348
rect -798 1280 -716 1288
rect -798 1216 -774 1280
rect -740 1216 -716 1280
rect -798 1212 -716 1216
rect -798 1110 -774 1212
rect -740 1110 -716 1212
rect -798 1106 -716 1110
rect -798 1042 -774 1106
rect -740 1042 -716 1106
rect -798 1034 -716 1042
rect -798 974 -774 1034
rect -740 974 -716 1034
rect -798 962 -716 974
rect -798 906 -774 962
rect -740 906 -716 962
rect -798 890 -716 906
rect -798 838 -774 890
rect -740 838 -716 890
rect -798 818 -716 838
rect -798 770 -774 818
rect -740 770 -716 818
rect -798 746 -716 770
rect -798 702 -774 746
rect -740 702 -716 746
rect -798 674 -716 702
rect -798 634 -774 674
rect -740 634 -716 674
rect -798 602 -716 634
rect -798 566 -774 602
rect -740 566 -716 602
rect -798 532 -716 566
rect -798 496 -774 532
rect -740 496 -716 532
rect -798 464 -716 496
rect -798 424 -774 464
rect -740 424 -716 464
rect -798 396 -716 424
rect -798 352 -774 396
rect -740 352 -716 396
rect -798 328 -716 352
rect -798 280 -774 328
rect -740 280 -716 328
rect -798 260 -716 280
rect -798 208 -774 260
rect -740 208 -716 260
rect -798 192 -716 208
rect -798 136 -774 192
rect -740 136 -716 192
rect -798 124 -716 136
rect -798 64 -774 124
rect -740 64 -716 124
rect -798 56 -716 64
rect -798 -8 -774 56
rect -740 -8 -716 56
rect -798 -12 -716 -8
rect -798 -114 -774 -12
rect -740 -114 -716 -12
rect -798 -118 -716 -114
rect -798 -182 -774 -118
rect -740 -182 -716 -118
rect -659 6146 -457 6165
rect -659 -152 -647 6146
rect -469 -152 -457 6146
rect -659 -164 -457 -152
rect -134 6146 284 6165
rect -134 -152 -122 6146
rect 272 -152 284 6146
rect -134 -164 284 -152
rect 607 6146 809 6165
rect 607 -152 619 6146
rect 797 -152 809 6146
rect 607 -164 809 -152
rect 866 6112 890 6176
rect 924 6112 948 6176
rect 866 6108 948 6112
rect 866 6006 890 6108
rect 924 6006 948 6108
rect 866 6002 948 6006
rect 866 5938 890 6002
rect 924 5938 948 6002
rect 866 5930 948 5938
rect 866 5870 890 5930
rect 924 5870 948 5930
rect 866 5858 948 5870
rect 866 5802 890 5858
rect 924 5802 948 5858
rect 866 5786 948 5802
rect 866 5734 890 5786
rect 924 5734 948 5786
rect 866 5714 948 5734
rect 866 5666 890 5714
rect 924 5666 948 5714
rect 866 5642 948 5666
rect 866 5598 890 5642
rect 924 5598 948 5642
rect 866 5570 948 5598
rect 866 5530 890 5570
rect 924 5530 948 5570
rect 866 5498 948 5530
rect 866 5462 890 5498
rect 924 5462 948 5498
rect 866 5428 948 5462
rect 866 5392 890 5428
rect 924 5392 948 5428
rect 866 5360 948 5392
rect 866 5320 890 5360
rect 924 5320 948 5360
rect 866 5292 948 5320
rect 866 5248 890 5292
rect 924 5248 948 5292
rect 866 5224 948 5248
rect 866 5176 890 5224
rect 924 5176 948 5224
rect 866 5156 948 5176
rect 866 5104 890 5156
rect 924 5104 948 5156
rect 866 5088 948 5104
rect 866 5032 890 5088
rect 924 5032 948 5088
rect 866 5020 948 5032
rect 866 4960 890 5020
rect 924 4960 948 5020
rect 866 4952 948 4960
rect 866 4888 890 4952
rect 924 4888 948 4952
rect 866 4884 948 4888
rect 866 4782 890 4884
rect 924 4782 948 4884
rect 866 4778 948 4782
rect 866 4714 890 4778
rect 924 4714 948 4778
rect 866 4706 948 4714
rect 866 4646 890 4706
rect 924 4646 948 4706
rect 866 4634 948 4646
rect 866 4578 890 4634
rect 924 4578 948 4634
rect 866 4562 948 4578
rect 866 4510 890 4562
rect 924 4510 948 4562
rect 866 4490 948 4510
rect 866 4442 890 4490
rect 924 4442 948 4490
rect 866 4418 948 4442
rect 866 4374 890 4418
rect 924 4374 948 4418
rect 866 4346 948 4374
rect 866 4306 890 4346
rect 924 4306 948 4346
rect 866 4274 948 4306
rect 866 4238 890 4274
rect 924 4238 948 4274
rect 866 4204 948 4238
rect 866 4168 890 4204
rect 924 4168 948 4204
rect 866 4136 948 4168
rect 866 4096 890 4136
rect 924 4096 948 4136
rect 866 4068 948 4096
rect 866 4024 890 4068
rect 924 4024 948 4068
rect 866 4000 948 4024
rect 866 3952 890 4000
rect 924 3952 948 4000
rect 866 3932 948 3952
rect 866 3880 890 3932
rect 924 3880 948 3932
rect 866 3864 948 3880
rect 866 3808 890 3864
rect 924 3808 948 3864
rect 866 3796 948 3808
rect 866 3736 890 3796
rect 924 3736 948 3796
rect 866 3728 948 3736
rect 866 3664 890 3728
rect 924 3664 948 3728
rect 866 3660 948 3664
rect 866 3558 890 3660
rect 924 3558 948 3660
rect 866 3554 948 3558
rect 866 3490 890 3554
rect 924 3490 948 3554
rect 866 3482 948 3490
rect 866 3422 890 3482
rect 924 3422 948 3482
rect 866 3410 948 3422
rect 866 3354 890 3410
rect 924 3354 948 3410
rect 866 3338 948 3354
rect 866 3286 890 3338
rect 924 3286 948 3338
rect 866 3266 948 3286
rect 866 3218 890 3266
rect 924 3218 948 3266
rect 866 3194 948 3218
rect 866 3150 890 3194
rect 924 3150 948 3194
rect 866 3122 948 3150
rect 866 3082 890 3122
rect 924 3082 948 3122
rect 866 3050 948 3082
rect 866 3014 890 3050
rect 924 3014 948 3050
rect 866 2980 948 3014
rect 866 2944 890 2980
rect 924 2944 948 2980
rect 866 2912 948 2944
rect 866 2872 890 2912
rect 924 2872 948 2912
rect 866 2844 948 2872
rect 866 2800 890 2844
rect 924 2800 948 2844
rect 866 2776 948 2800
rect 866 2728 890 2776
rect 924 2728 948 2776
rect 866 2708 948 2728
rect 866 2656 890 2708
rect 924 2656 948 2708
rect 866 2640 948 2656
rect 866 2584 890 2640
rect 924 2584 948 2640
rect 866 2572 948 2584
rect 866 2512 890 2572
rect 924 2512 948 2572
rect 866 2504 948 2512
rect 866 2440 890 2504
rect 924 2440 948 2504
rect 866 2436 948 2440
rect 866 2334 890 2436
rect 924 2334 948 2436
rect 866 2330 948 2334
rect 866 2266 890 2330
rect 924 2266 948 2330
rect 866 2258 948 2266
rect 866 2198 890 2258
rect 924 2198 948 2258
rect 866 2186 948 2198
rect 866 2130 890 2186
rect 924 2130 948 2186
rect 866 2114 948 2130
rect 866 2062 890 2114
rect 924 2062 948 2114
rect 866 2042 948 2062
rect 866 1994 890 2042
rect 924 1994 948 2042
rect 866 1970 948 1994
rect 866 1926 890 1970
rect 924 1926 948 1970
rect 866 1898 948 1926
rect 866 1858 890 1898
rect 924 1858 948 1898
rect 866 1826 948 1858
rect 866 1790 890 1826
rect 924 1790 948 1826
rect 866 1756 948 1790
rect 866 1720 890 1756
rect 924 1720 948 1756
rect 866 1688 948 1720
rect 866 1648 890 1688
rect 924 1648 948 1688
rect 866 1620 948 1648
rect 866 1576 890 1620
rect 924 1576 948 1620
rect 866 1552 948 1576
rect 866 1504 890 1552
rect 924 1504 948 1552
rect 866 1484 948 1504
rect 866 1432 890 1484
rect 924 1432 948 1484
rect 866 1416 948 1432
rect 866 1360 890 1416
rect 924 1360 948 1416
rect 866 1348 948 1360
rect 866 1288 890 1348
rect 924 1288 948 1348
rect 866 1280 948 1288
rect 866 1216 890 1280
rect 924 1216 948 1280
rect 866 1212 948 1216
rect 866 1110 890 1212
rect 924 1110 948 1212
rect 866 1106 948 1110
rect 866 1042 890 1106
rect 924 1042 948 1106
rect 866 1034 948 1042
rect 866 974 890 1034
rect 924 974 948 1034
rect 866 962 948 974
rect 866 906 890 962
rect 924 906 948 962
rect 866 890 948 906
rect 866 838 890 890
rect 924 838 948 890
rect 866 818 948 838
rect 866 770 890 818
rect 924 770 948 818
rect 866 746 948 770
rect 866 702 890 746
rect 924 702 948 746
rect 866 674 948 702
rect 866 634 890 674
rect 924 634 948 674
rect 866 602 948 634
rect 866 566 890 602
rect 924 566 948 602
rect 866 532 948 566
rect 866 496 890 532
rect 924 496 948 532
rect 866 464 948 496
rect 866 424 890 464
rect 924 424 948 464
rect 866 396 948 424
rect 866 352 890 396
rect 924 352 948 396
rect 866 328 948 352
rect 866 280 890 328
rect 924 280 948 328
rect 866 260 948 280
rect 866 208 890 260
rect 924 208 948 260
rect 866 192 948 208
rect 866 136 890 192
rect 924 136 948 192
rect 866 124 948 136
rect 866 64 890 124
rect 924 64 948 124
rect 866 56 948 64
rect 866 -8 890 56
rect 924 -8 948 56
rect 866 -12 948 -8
rect 866 -114 890 -12
rect 924 -114 948 -12
rect 866 -118 948 -114
rect -798 -190 -716 -182
rect -798 -250 -774 -190
rect -740 -250 -716 -190
rect -798 -262 -716 -250
rect -798 -318 -774 -262
rect -740 -318 -716 -262
rect -798 -334 -716 -318
rect -798 -386 -774 -334
rect -740 -386 -716 -334
rect -798 -406 -716 -386
rect -798 -454 -774 -406
rect -740 -454 -716 -406
rect 866 -182 890 -118
rect 924 -182 948 -118
rect 866 -190 948 -182
rect 866 -250 890 -190
rect 924 -250 948 -190
rect 866 -262 948 -250
rect 866 -318 890 -262
rect 924 -318 948 -262
rect 866 -334 948 -318
rect 866 -386 890 -334
rect 924 -386 948 -334
rect 866 -406 948 -386
rect -798 -478 -716 -454
rect -798 -522 -774 -478
rect -740 -522 -716 -478
rect -798 -550 -716 -522
rect -798 -590 -774 -550
rect -740 -590 -716 -550
rect -798 -622 -716 -590
rect -798 -658 -774 -622
rect -740 -658 -716 -622
rect -146 -459 290 -443
rect -146 -493 -130 -459
rect -96 -493 -56 -459
rect -22 -493 18 -459
rect 52 -493 92 -459
rect 126 -493 166 -459
rect 200 -493 240 -459
rect 274 -493 290 -459
rect -146 -533 290 -493
rect -146 -567 -130 -533
rect -96 -567 -56 -533
rect -22 -567 18 -533
rect 52 -567 92 -533
rect 126 -567 166 -533
rect 200 -567 240 -533
rect 274 -567 290 -533
rect -146 -607 290 -567
rect -146 -641 -130 -607
rect -96 -641 -56 -607
rect -22 -641 18 -607
rect 52 -641 92 -607
rect 126 -641 166 -607
rect 200 -641 240 -607
rect 274 -641 290 -607
rect -146 -657 290 -641
rect 866 -454 890 -406
rect 924 -454 948 -406
rect 866 -478 948 -454
rect 866 -522 890 -478
rect 924 -522 948 -478
rect 866 -550 948 -522
rect 866 -590 890 -550
rect 924 -590 948 -550
rect 866 -622 948 -590
rect -798 -692 -716 -658
rect -798 -726 -774 -692
rect -740 -726 -716 -692
rect -798 -757 -716 -726
rect 866 -658 890 -622
rect 924 -658 948 -622
rect 866 -692 948 -658
rect 866 -726 890 -692
rect 924 -726 948 -692
rect 866 -757 948 -726
rect -798 -760 948 -757
rect -798 -794 -774 -760
rect -740 -794 890 -760
rect 924 -794 948 -760
rect -798 -820 948 -794
rect -798 -828 -554 -820
rect -798 -862 -774 -828
rect -740 -862 -554 -828
rect -798 -896 -554 -862
rect -798 -930 -774 -896
rect -740 -930 -554 -896
rect -798 -964 -554 -930
rect 704 -828 948 -820
rect 704 -862 890 -828
rect 924 -862 948 -828
rect 704 -896 948 -862
rect 704 -930 890 -896
rect 924 -930 948 -896
rect 704 -964 948 -930
rect -798 -998 -774 -964
rect -740 -998 -554 -964
rect 704 -998 890 -964
rect 924 -998 948 -964
rect -798 -1022 948 -998
rect 1648 7013 1730 7026
rect 1648 6958 1672 7013
rect 1706 6958 1730 7013
rect 1648 6941 1730 6958
rect 1648 6890 1672 6941
rect 1706 6890 1730 6941
rect 1648 6869 1730 6890
rect 1648 6822 1672 6869
rect 1706 6822 1730 6869
rect 1648 6797 1730 6822
rect 1648 6754 1672 6797
rect 1706 6754 1730 6797
rect 1648 6725 1730 6754
rect 1648 6686 1672 6725
rect 1706 6686 1730 6725
rect 1648 6653 1730 6686
rect 1648 6618 1672 6653
rect 1706 6618 1730 6653
rect 1648 6584 1730 6618
rect 1648 6547 1672 6584
rect 1706 6547 1730 6584
rect 1648 6516 1730 6547
rect 1648 6475 1672 6516
rect 1706 6475 1730 6516
rect 1648 6448 1730 6475
rect 1648 6403 1672 6448
rect 1706 6403 1730 6448
rect 1648 6380 1730 6403
rect 1648 6331 1672 6380
rect 1706 6331 1730 6380
rect 1648 6312 1730 6331
rect 1648 6259 1672 6312
rect 1706 6259 1730 6312
rect 1648 6244 1730 6259
rect 1648 6187 1672 6244
rect 1706 6187 1730 6244
rect 1648 6176 1730 6187
rect 1648 6115 1672 6176
rect 1706 6115 1730 6176
rect 1648 6108 1730 6115
rect 1648 6043 1672 6108
rect 1706 6043 1730 6108
rect 1648 6040 1730 6043
rect 1648 6006 1672 6040
rect 1706 6006 1730 6040
rect 1648 6005 1730 6006
rect 1648 5938 1672 6005
rect 1706 5938 1730 6005
rect 1648 5933 1730 5938
rect 1648 5870 1672 5933
rect 1706 5870 1730 5933
rect 1648 5861 1730 5870
rect 1648 5802 1672 5861
rect 1706 5802 1730 5861
rect 1648 5789 1730 5802
rect 1648 5734 1672 5789
rect 1706 5734 1730 5789
rect 1648 5717 1730 5734
rect 1648 5666 1672 5717
rect 1706 5666 1730 5717
rect 1648 5645 1730 5666
rect 1648 5598 1672 5645
rect 1706 5598 1730 5645
rect 1648 5573 1730 5598
rect 1648 5530 1672 5573
rect 1706 5530 1730 5573
rect 1648 5501 1730 5530
rect 1648 5462 1672 5501
rect 1706 5462 1730 5501
rect 1648 5429 1730 5462
rect 1648 5394 1672 5429
rect 1706 5394 1730 5429
rect 1648 5360 1730 5394
rect 1648 5323 1672 5360
rect 1706 5323 1730 5360
rect 1648 5292 1730 5323
rect 1648 5251 1672 5292
rect 1706 5251 1730 5292
rect 1648 5224 1730 5251
rect 1648 5179 1672 5224
rect 1706 5179 1730 5224
rect 1648 5156 1730 5179
rect 1648 5107 1672 5156
rect 1706 5107 1730 5156
rect 1648 5088 1730 5107
rect 1648 5035 1672 5088
rect 1706 5035 1730 5088
rect 1648 5020 1730 5035
rect 1648 4963 1672 5020
rect 1706 4963 1730 5020
rect 1648 4952 1730 4963
rect 1648 4891 1672 4952
rect 1706 4891 1730 4952
rect 1648 4884 1730 4891
rect 1648 4819 1672 4884
rect 1706 4819 1730 4884
rect 1648 4816 1730 4819
rect 1648 4782 1672 4816
rect 1706 4782 1730 4816
rect 1648 4781 1730 4782
rect 1648 4714 1672 4781
rect 1706 4714 1730 4781
rect 1648 4709 1730 4714
rect 1648 4646 1672 4709
rect 1706 4646 1730 4709
rect 1648 4637 1730 4646
rect 1648 4578 1672 4637
rect 1706 4578 1730 4637
rect 1648 4565 1730 4578
rect 1648 4510 1672 4565
rect 1706 4510 1730 4565
rect 1648 4493 1730 4510
rect 1648 4442 1672 4493
rect 1706 4442 1730 4493
rect 1648 4421 1730 4442
rect 1648 4374 1672 4421
rect 1706 4374 1730 4421
rect 1648 4349 1730 4374
rect 1648 4306 1672 4349
rect 1706 4306 1730 4349
rect 1648 4277 1730 4306
rect 1648 4238 1672 4277
rect 1706 4238 1730 4277
rect 1648 4205 1730 4238
rect 1648 4170 1672 4205
rect 1706 4170 1730 4205
rect 1648 4136 1730 4170
rect 1648 4099 1672 4136
rect 1706 4099 1730 4136
rect 1648 4068 1730 4099
rect 1648 4027 1672 4068
rect 1706 4027 1730 4068
rect 1648 4000 1730 4027
rect 1648 3955 1672 4000
rect 1706 3955 1730 4000
rect 1648 3932 1730 3955
rect 1648 3883 1672 3932
rect 1706 3883 1730 3932
rect 1648 3864 1730 3883
rect 1648 3811 1672 3864
rect 1706 3811 1730 3864
rect 1648 3796 1730 3811
rect 1648 3739 1672 3796
rect 1706 3739 1730 3796
rect 1648 3728 1730 3739
rect 1648 3667 1672 3728
rect 1706 3667 1730 3728
rect 1648 3660 1730 3667
rect 1648 3595 1672 3660
rect 1706 3595 1730 3660
rect 1648 3592 1730 3595
rect 1648 3558 1672 3592
rect 1706 3558 1730 3592
rect 1648 3557 1730 3558
rect 1648 3490 1672 3557
rect 1706 3490 1730 3557
rect 1648 3485 1730 3490
rect 1648 3422 1672 3485
rect 1706 3422 1730 3485
rect 1648 3413 1730 3422
rect 1648 3354 1672 3413
rect 1706 3354 1730 3413
rect 1648 3341 1730 3354
rect 1648 3286 1672 3341
rect 1706 3286 1730 3341
rect 1648 3269 1730 3286
rect 1648 3218 1672 3269
rect 1706 3218 1730 3269
rect 1648 3197 1730 3218
rect 1648 3150 1672 3197
rect 1706 3150 1730 3197
rect 1648 3125 1730 3150
rect 1648 3082 1672 3125
rect 1706 3082 1730 3125
rect 1648 3053 1730 3082
rect 1648 3014 1672 3053
rect 1706 3014 1730 3053
rect 1648 2981 1730 3014
rect 1648 2946 1672 2981
rect 1706 2946 1730 2981
rect 1648 2912 1730 2946
rect 1648 2875 1672 2912
rect 1706 2875 1730 2912
rect 1648 2844 1730 2875
rect 1648 2803 1672 2844
rect 1706 2803 1730 2844
rect 1648 2776 1730 2803
rect 1648 2731 1672 2776
rect 1706 2731 1730 2776
rect 1648 2708 1730 2731
rect 1648 2659 1672 2708
rect 1706 2659 1730 2708
rect 1648 2640 1730 2659
rect 1648 2587 1672 2640
rect 1706 2587 1730 2640
rect 1648 2572 1730 2587
rect 1648 2515 1672 2572
rect 1706 2515 1730 2572
rect 1648 2504 1730 2515
rect 1648 2443 1672 2504
rect 1706 2443 1730 2504
rect 1648 2436 1730 2443
rect 1648 2371 1672 2436
rect 1706 2371 1730 2436
rect 1648 2368 1730 2371
rect 1648 2334 1672 2368
rect 1706 2334 1730 2368
rect 1648 2333 1730 2334
rect 1648 2266 1672 2333
rect 1706 2266 1730 2333
rect 1648 2261 1730 2266
rect 1648 2198 1672 2261
rect 1706 2198 1730 2261
rect 1648 2189 1730 2198
rect 1648 2130 1672 2189
rect 1706 2130 1730 2189
rect 1648 2117 1730 2130
rect 1648 2062 1672 2117
rect 1706 2062 1730 2117
rect 1648 2045 1730 2062
rect 1648 1994 1672 2045
rect 1706 1994 1730 2045
rect 1648 1973 1730 1994
rect 1648 1926 1672 1973
rect 1706 1926 1730 1973
rect 1648 1901 1730 1926
rect 1648 1858 1672 1901
rect 1706 1858 1730 1901
rect 1648 1829 1730 1858
rect 1648 1790 1672 1829
rect 1706 1790 1730 1829
rect 1648 1757 1730 1790
rect 1648 1722 1672 1757
rect 1706 1722 1730 1757
rect 1648 1688 1730 1722
rect 1648 1651 1672 1688
rect 1706 1651 1730 1688
rect 1648 1620 1730 1651
rect 1648 1579 1672 1620
rect 1706 1579 1730 1620
rect 1648 1552 1730 1579
rect 1648 1507 1672 1552
rect 1706 1507 1730 1552
rect 1648 1484 1730 1507
rect 1648 1435 1672 1484
rect 1706 1435 1730 1484
rect 1648 1416 1730 1435
rect 1648 1363 1672 1416
rect 1706 1363 1730 1416
rect 1648 1348 1730 1363
rect 1648 1291 1672 1348
rect 1706 1291 1730 1348
rect 1648 1280 1730 1291
rect 1648 1219 1672 1280
rect 1706 1219 1730 1280
rect 1648 1212 1730 1219
rect 1648 1147 1672 1212
rect 1706 1147 1730 1212
rect 1648 1144 1730 1147
rect 1648 1110 1672 1144
rect 1706 1110 1730 1144
rect 1648 1109 1730 1110
rect 1648 1042 1672 1109
rect 1706 1042 1730 1109
rect 1648 1037 1730 1042
rect 1648 974 1672 1037
rect 1706 974 1730 1037
rect 1648 965 1730 974
rect 1648 906 1672 965
rect 1706 906 1730 965
rect 1648 893 1730 906
rect 1648 838 1672 893
rect 1706 838 1730 893
rect 1648 821 1730 838
rect 1648 770 1672 821
rect 1706 770 1730 821
rect 1648 749 1730 770
rect 1648 702 1672 749
rect 1706 702 1730 749
rect 1648 677 1730 702
rect 1648 634 1672 677
rect 1706 634 1730 677
rect 1648 605 1730 634
rect 1648 566 1672 605
rect 1706 566 1730 605
rect 1648 533 1730 566
rect 1648 498 1672 533
rect 1706 498 1730 533
rect 1648 464 1730 498
rect 1648 427 1672 464
rect 1706 427 1730 464
rect 1648 396 1730 427
rect 1648 355 1672 396
rect 1706 355 1730 396
rect 1648 328 1730 355
rect 1648 283 1672 328
rect 1706 283 1730 328
rect 1648 260 1730 283
rect 1648 211 1672 260
rect 1706 211 1730 260
rect 1648 192 1730 211
rect 1648 139 1672 192
rect 1706 139 1730 192
rect 1648 124 1730 139
rect 1648 67 1672 124
rect 1706 67 1730 124
rect 1648 56 1730 67
rect 1648 -5 1672 56
rect 1706 -5 1730 56
rect 1648 -12 1730 -5
rect 1648 -77 1672 -12
rect 1706 -77 1730 -12
rect 1648 -80 1730 -77
rect 1648 -114 1672 -80
rect 1706 -114 1730 -80
rect 1648 -115 1730 -114
rect 1648 -182 1672 -115
rect 1706 -182 1730 -115
rect 1648 -187 1730 -182
rect 1648 -250 1672 -187
rect 1706 -250 1730 -187
rect 1648 -259 1730 -250
rect 1648 -318 1672 -259
rect 1706 -318 1730 -259
rect 1648 -331 1730 -318
rect 1648 -386 1672 -331
rect 1706 -386 1730 -331
rect 1648 -403 1730 -386
rect 1648 -454 1672 -403
rect 1706 -454 1730 -403
rect 1648 -475 1730 -454
rect 1648 -522 1672 -475
rect 1706 -522 1730 -475
rect 1648 -547 1730 -522
rect 1648 -590 1672 -547
rect 1706 -590 1730 -547
rect 1648 -619 1730 -590
rect 1648 -658 1672 -619
rect 1706 -658 1730 -619
rect 1648 -691 1730 -658
rect 1648 -726 1672 -691
rect 1706 -726 1730 -691
rect 1648 -760 1730 -726
rect 1648 -797 1672 -760
rect 1706 -797 1730 -760
rect 1648 -828 1730 -797
rect 1648 -869 1672 -828
rect 1706 -869 1730 -828
rect 1648 -896 1730 -869
rect 1648 -941 1672 -896
rect 1706 -941 1730 -896
rect 1648 -964 1730 -941
rect 1648 -1013 1672 -964
rect 1706 -1013 1730 -964
rect -1580 -1085 -1556 -1032
rect -1522 -1085 -1498 -1032
rect -1580 -1100 -1498 -1085
rect -1580 -1157 -1556 -1100
rect -1522 -1157 -1498 -1100
rect -1580 -1168 -1498 -1157
rect -1580 -1229 -1556 -1168
rect -1522 -1229 -1498 -1168
rect -1580 -1236 -1498 -1229
rect -1580 -1301 -1556 -1236
rect -1522 -1301 -1498 -1236
rect -1580 -1304 -1498 -1301
rect -1580 -1338 -1556 -1304
rect -1522 -1338 -1498 -1304
rect -1580 -1339 -1498 -1338
rect -1580 -1406 -1556 -1339
rect -1522 -1406 -1498 -1339
rect -1580 -1411 -1498 -1406
rect -1580 -1474 -1556 -1411
rect -1522 -1474 -1498 -1411
rect -1580 -1483 -1498 -1474
rect -1580 -1542 -1556 -1483
rect -1522 -1542 -1498 -1483
rect -1580 -1555 -1498 -1542
rect -1580 -1610 -1556 -1555
rect -1522 -1610 -1498 -1555
rect -1580 -1627 -1498 -1610
rect -1580 -1678 -1556 -1627
rect -1522 -1678 -1498 -1627
rect -1580 -1722 -1498 -1678
rect 1648 -1032 1730 -1013
rect 1648 -1085 1672 -1032
rect 1706 -1085 1730 -1032
rect 1648 -1100 1730 -1085
rect 1648 -1157 1672 -1100
rect 1706 -1157 1730 -1100
rect 1648 -1168 1730 -1157
rect 1648 -1229 1672 -1168
rect 1706 -1229 1730 -1168
rect 1648 -1236 1730 -1229
rect 1648 -1301 1672 -1236
rect 1706 -1301 1730 -1236
rect 1648 -1304 1730 -1301
rect 1648 -1338 1672 -1304
rect 1706 -1338 1730 -1304
rect 1648 -1339 1730 -1338
rect 1648 -1406 1672 -1339
rect 1706 -1406 1730 -1339
rect 1648 -1411 1730 -1406
rect 1648 -1474 1672 -1411
rect 1706 -1474 1730 -1411
rect 1648 -1483 1730 -1474
rect 1648 -1542 1672 -1483
rect 1706 -1542 1730 -1483
rect 1648 -1555 1730 -1542
rect 1648 -1610 1672 -1555
rect 1706 -1610 1730 -1555
rect 1648 -1627 1730 -1610
rect 1648 -1678 1672 -1627
rect 1706 -1678 1730 -1627
rect 1648 -1722 1730 -1678
rect -1580 -1746 1730 -1722
rect -1580 -1780 -1472 -1746
rect -1420 -1780 -1404 -1746
rect -1348 -1780 -1336 -1746
rect -1276 -1780 -1268 -1746
rect -1204 -1780 -1200 -1746
rect -1098 -1780 -1094 -1746
rect -1030 -1780 -1022 -1746
rect -962 -1780 -950 -1746
rect -894 -1780 -878 -1746
rect -826 -1780 -806 -1746
rect -758 -1780 -734 -1746
rect -690 -1780 -662 -1746
rect -622 -1780 -590 -1746
rect -554 -1780 -520 -1746
rect -484 -1780 -452 -1746
rect -412 -1780 -384 -1746
rect -340 -1780 -316 -1746
rect -268 -1780 -248 -1746
rect -196 -1780 -180 -1746
rect -124 -1780 -112 -1746
rect -52 -1780 -44 -1746
rect 20 -1780 24 -1746
rect 126 -1780 130 -1746
rect 194 -1780 202 -1746
rect 262 -1780 274 -1746
rect 330 -1780 346 -1746
rect 398 -1780 418 -1746
rect 466 -1780 490 -1746
rect 534 -1780 562 -1746
rect 602 -1780 634 -1746
rect 670 -1780 704 -1746
rect 740 -1780 772 -1746
rect 812 -1780 840 -1746
rect 884 -1780 908 -1746
rect 956 -1780 976 -1746
rect 1028 -1780 1044 -1746
rect 1100 -1780 1112 -1746
rect 1172 -1780 1180 -1746
rect 1244 -1780 1248 -1746
rect 1350 -1780 1354 -1746
rect 1418 -1780 1426 -1746
rect 1486 -1780 1498 -1746
rect 1554 -1780 1570 -1746
rect 1622 -1780 1730 -1746
rect -1580 -1804 1730 -1780
<< viali >>
rect -1454 7746 -1438 7780
rect -1438 7746 -1420 7780
rect -1382 7746 -1370 7780
rect -1370 7746 -1348 7780
rect -1310 7746 -1302 7780
rect -1302 7746 -1276 7780
rect -1238 7746 -1234 7780
rect -1234 7746 -1204 7780
rect -1166 7746 -1132 7780
rect -1094 7746 -1064 7780
rect -1064 7746 -1060 7780
rect -1022 7746 -996 7780
rect -996 7746 -988 7780
rect -950 7746 -928 7780
rect -928 7746 -916 7780
rect -878 7746 -860 7780
rect -860 7746 -844 7780
rect -806 7746 -792 7780
rect -792 7746 -772 7780
rect -734 7746 -724 7780
rect -724 7746 -700 7780
rect -662 7746 -656 7780
rect -656 7746 -628 7780
rect -590 7746 -588 7780
rect -588 7746 -556 7780
rect -518 7746 -486 7780
rect -486 7746 -484 7780
rect -446 7746 -418 7780
rect -418 7746 -412 7780
rect -374 7746 -350 7780
rect -350 7746 -340 7780
rect -302 7746 -282 7780
rect -282 7746 -268 7780
rect -230 7746 -214 7780
rect -214 7746 -196 7780
rect -158 7746 -146 7780
rect -146 7746 -124 7780
rect -86 7746 -78 7780
rect -78 7746 -52 7780
rect -14 7746 -10 7780
rect -10 7746 20 7780
rect 58 7746 92 7780
rect 130 7746 160 7780
rect 160 7746 164 7780
rect 202 7746 228 7780
rect 228 7746 236 7780
rect 274 7746 296 7780
rect 296 7746 308 7780
rect 346 7746 364 7780
rect 364 7746 380 7780
rect 418 7746 432 7780
rect 432 7746 452 7780
rect 490 7746 500 7780
rect 500 7746 524 7780
rect 562 7746 568 7780
rect 568 7746 596 7780
rect 634 7746 636 7780
rect 636 7746 668 7780
rect 706 7746 738 7780
rect 738 7746 740 7780
rect 778 7746 806 7780
rect 806 7746 812 7780
rect 850 7746 874 7780
rect 874 7746 884 7780
rect 922 7746 942 7780
rect 942 7746 956 7780
rect 994 7746 1010 7780
rect 1010 7746 1028 7780
rect 1066 7746 1078 7780
rect 1078 7746 1100 7780
rect 1138 7746 1146 7780
rect 1146 7746 1172 7780
rect 1210 7746 1214 7780
rect 1214 7746 1244 7780
rect 1282 7746 1316 7780
rect 1354 7746 1384 7780
rect 1384 7746 1388 7780
rect 1426 7746 1452 7780
rect 1452 7746 1460 7780
rect 1498 7746 1520 7780
rect 1520 7746 1532 7780
rect 1570 7746 1588 7780
rect 1588 7746 1604 7780
rect -1556 7638 -1522 7661
rect -1556 7627 -1522 7638
rect -1556 7570 -1522 7589
rect -1556 7555 -1522 7570
rect -1556 7502 -1522 7517
rect -1556 7483 -1522 7502
rect -1556 7434 -1522 7445
rect -1556 7411 -1522 7434
rect -1556 7366 -1522 7373
rect -1556 7339 -1522 7366
rect -1556 7298 -1522 7301
rect -1556 7267 -1522 7298
rect -1556 7196 -1522 7229
rect -1556 7195 -1522 7196
rect -1556 7128 -1522 7157
rect -1556 7123 -1522 7128
rect -1556 7060 -1522 7085
rect -1556 7051 -1522 7060
rect 1672 7638 1706 7661
rect 1672 7627 1706 7638
rect 1672 7570 1706 7589
rect 1672 7555 1706 7570
rect 1672 7502 1706 7517
rect 1672 7483 1706 7502
rect 1672 7434 1706 7445
rect 1672 7411 1706 7434
rect 1672 7366 1706 7373
rect 1672 7339 1706 7366
rect 1672 7298 1706 7301
rect 1672 7267 1706 7298
rect 1672 7196 1706 7229
rect 1672 7195 1706 7196
rect 1672 7128 1706 7157
rect 1672 7123 1706 7128
rect 1672 7060 1706 7085
rect 1672 7051 1706 7060
rect -1556 6992 -1522 7013
rect -1556 6979 -1522 6992
rect -1556 6924 -1522 6941
rect -1556 6907 -1522 6924
rect -1556 6856 -1522 6869
rect -1556 6835 -1522 6856
rect -1556 6788 -1522 6797
rect -1556 6763 -1522 6788
rect -1556 6720 -1522 6725
rect -1556 6691 -1522 6720
rect -1556 6652 -1522 6653
rect -1556 6619 -1522 6652
rect -1556 6550 -1522 6581
rect -1556 6547 -1522 6550
rect -1556 6482 -1522 6509
rect -1556 6475 -1522 6482
rect -1556 6414 -1522 6437
rect -1556 6403 -1522 6414
rect -1556 6346 -1522 6365
rect -1556 6331 -1522 6346
rect -1556 6278 -1522 6293
rect -1556 6259 -1522 6278
rect -1556 6210 -1522 6221
rect -1556 6187 -1522 6210
rect -1556 6142 -1522 6149
rect -1556 6115 -1522 6142
rect -1556 6074 -1522 6077
rect -1556 6043 -1522 6074
rect -1556 5972 -1522 6005
rect -1556 5971 -1522 5972
rect -1556 5904 -1522 5933
rect -1556 5899 -1522 5904
rect -1556 5836 -1522 5861
rect -1556 5827 -1522 5836
rect -1556 5768 -1522 5789
rect -1556 5755 -1522 5768
rect -1556 5700 -1522 5717
rect -1556 5683 -1522 5700
rect -1556 5632 -1522 5645
rect -1556 5611 -1522 5632
rect -1556 5564 -1522 5573
rect -1556 5539 -1522 5564
rect -1556 5496 -1522 5501
rect -1556 5467 -1522 5496
rect -1556 5428 -1522 5429
rect -1556 5395 -1522 5428
rect -1556 5326 -1522 5357
rect -1556 5323 -1522 5326
rect -1556 5258 -1522 5285
rect -1556 5251 -1522 5258
rect -1556 5190 -1522 5213
rect -1556 5179 -1522 5190
rect -1556 5122 -1522 5141
rect -1556 5107 -1522 5122
rect -1556 5054 -1522 5069
rect -1556 5035 -1522 5054
rect -1556 4986 -1522 4997
rect -1556 4963 -1522 4986
rect -1556 4918 -1522 4925
rect -1556 4891 -1522 4918
rect -1556 4850 -1522 4853
rect -1556 4819 -1522 4850
rect -1556 4748 -1522 4781
rect -1556 4747 -1522 4748
rect -1556 4680 -1522 4709
rect -1556 4675 -1522 4680
rect -1556 4612 -1522 4637
rect -1556 4603 -1522 4612
rect -1556 4544 -1522 4565
rect -1556 4531 -1522 4544
rect -1556 4476 -1522 4493
rect -1556 4459 -1522 4476
rect -1556 4408 -1522 4421
rect -1556 4387 -1522 4408
rect -1556 4340 -1522 4349
rect -1556 4315 -1522 4340
rect -1556 4272 -1522 4277
rect -1556 4243 -1522 4272
rect -1556 4204 -1522 4205
rect -1556 4171 -1522 4204
rect -1556 4102 -1522 4133
rect -1556 4099 -1522 4102
rect -1556 4034 -1522 4061
rect -1556 4027 -1522 4034
rect -1556 3966 -1522 3989
rect -1556 3955 -1522 3966
rect -1556 3898 -1522 3917
rect -1556 3883 -1522 3898
rect -1556 3830 -1522 3845
rect -1556 3811 -1522 3830
rect -1556 3762 -1522 3773
rect -1556 3739 -1522 3762
rect -1556 3694 -1522 3701
rect -1556 3667 -1522 3694
rect -1556 3626 -1522 3629
rect -1556 3595 -1522 3626
rect -1556 3524 -1522 3557
rect -1556 3523 -1522 3524
rect -1556 3456 -1522 3485
rect -1556 3451 -1522 3456
rect -1556 3388 -1522 3413
rect -1556 3379 -1522 3388
rect -1556 3320 -1522 3341
rect -1556 3307 -1522 3320
rect -1556 3252 -1522 3269
rect -1556 3235 -1522 3252
rect -1556 3184 -1522 3197
rect -1556 3163 -1522 3184
rect -1556 3116 -1522 3125
rect -1556 3091 -1522 3116
rect -1556 3048 -1522 3053
rect -1556 3019 -1522 3048
rect -1556 2980 -1522 2981
rect -1556 2947 -1522 2980
rect -1556 2878 -1522 2909
rect -1556 2875 -1522 2878
rect -1556 2810 -1522 2837
rect -1556 2803 -1522 2810
rect -1556 2742 -1522 2765
rect -1556 2731 -1522 2742
rect -1556 2674 -1522 2693
rect -1556 2659 -1522 2674
rect -1556 2606 -1522 2621
rect -1556 2587 -1522 2606
rect -1556 2538 -1522 2549
rect -1556 2515 -1522 2538
rect -1556 2470 -1522 2477
rect -1556 2443 -1522 2470
rect -1556 2402 -1522 2405
rect -1556 2371 -1522 2402
rect -1556 2300 -1522 2333
rect -1556 2299 -1522 2300
rect -1556 2232 -1522 2261
rect -1556 2227 -1522 2232
rect -1556 2164 -1522 2189
rect -1556 2155 -1522 2164
rect -1556 2096 -1522 2117
rect -1556 2083 -1522 2096
rect -1556 2028 -1522 2045
rect -1556 2011 -1522 2028
rect -1556 1960 -1522 1973
rect -1556 1939 -1522 1960
rect -1556 1892 -1522 1901
rect -1556 1867 -1522 1892
rect -1556 1824 -1522 1829
rect -1556 1795 -1522 1824
rect -1556 1756 -1522 1757
rect -1556 1723 -1522 1756
rect -1556 1654 -1522 1685
rect -1556 1651 -1522 1654
rect -1556 1586 -1522 1613
rect -1556 1579 -1522 1586
rect -1556 1518 -1522 1541
rect -1556 1507 -1522 1518
rect -1556 1450 -1522 1469
rect -1556 1435 -1522 1450
rect -1556 1382 -1522 1397
rect -1556 1363 -1522 1382
rect -1556 1314 -1522 1325
rect -1556 1291 -1522 1314
rect -1556 1246 -1522 1253
rect -1556 1219 -1522 1246
rect -1556 1178 -1522 1181
rect -1556 1147 -1522 1178
rect -1556 1076 -1522 1109
rect -1556 1075 -1522 1076
rect -1556 1008 -1522 1037
rect -1556 1003 -1522 1008
rect -1556 940 -1522 965
rect -1556 931 -1522 940
rect -1556 872 -1522 893
rect -1556 859 -1522 872
rect -1556 804 -1522 821
rect -1556 787 -1522 804
rect -1556 736 -1522 749
rect -1556 715 -1522 736
rect -1556 668 -1522 677
rect -1556 643 -1522 668
rect -1556 600 -1522 605
rect -1556 571 -1522 600
rect -1556 532 -1522 533
rect -1556 499 -1522 532
rect -1556 430 -1522 461
rect -1556 427 -1522 430
rect -1556 362 -1522 389
rect -1556 355 -1522 362
rect -1556 294 -1522 317
rect -1556 283 -1522 294
rect -1556 226 -1522 245
rect -1556 211 -1522 226
rect -1556 158 -1522 173
rect -1556 139 -1522 158
rect -1556 90 -1522 101
rect -1556 67 -1522 90
rect -1556 22 -1522 29
rect -1556 -5 -1522 22
rect -1556 -46 -1522 -43
rect -1556 -77 -1522 -46
rect -1556 -148 -1522 -115
rect -1556 -149 -1522 -148
rect -1556 -216 -1522 -187
rect -1556 -221 -1522 -216
rect -1556 -284 -1522 -259
rect -1556 -293 -1522 -284
rect -1556 -352 -1522 -331
rect -1556 -365 -1522 -352
rect -1556 -420 -1522 -403
rect -1556 -437 -1522 -420
rect -1556 -488 -1522 -475
rect -1556 -509 -1522 -488
rect -1556 -556 -1522 -547
rect -1556 -581 -1522 -556
rect -1556 -624 -1522 -619
rect -1556 -653 -1522 -624
rect -1556 -692 -1522 -691
rect -1556 -725 -1522 -692
rect -1556 -794 -1522 -763
rect -1556 -797 -1522 -794
rect -1556 -862 -1522 -835
rect -1556 -869 -1522 -862
rect -1556 -930 -1522 -907
rect -1556 -941 -1522 -930
rect -1556 -998 -1522 -979
rect -1556 -1013 -1522 -998
rect -554 6964 -520 6998
rect -520 6964 -486 6998
rect -486 6964 -452 6998
rect -452 6964 -418 6998
rect -418 6964 -384 6998
rect -384 6964 -350 6998
rect -350 6964 -316 6998
rect -316 6964 -282 6998
rect -282 6964 -248 6998
rect -248 6964 -214 6998
rect -214 6964 -180 6998
rect -180 6964 -146 6998
rect -146 6964 -112 6998
rect -112 6964 -78 6998
rect -78 6964 -44 6998
rect -44 6964 -10 6998
rect -10 6964 24 6998
rect 24 6964 58 6998
rect 58 6964 92 6998
rect 92 6964 126 6998
rect 126 6964 160 6998
rect 160 6964 194 6998
rect 194 6964 228 6998
rect 228 6964 262 6998
rect 262 6964 296 6998
rect 296 6964 330 6998
rect 330 6964 364 6998
rect 364 6964 398 6998
rect 398 6964 432 6998
rect 432 6964 466 6998
rect 466 6964 500 6998
rect 500 6964 534 6998
rect 534 6964 568 6998
rect 568 6964 602 6998
rect 602 6964 636 6998
rect 636 6964 670 6998
rect 670 6964 704 6998
rect -554 6820 704 6964
rect -774 6618 -740 6650
rect -774 6616 -740 6618
rect -774 6550 -740 6578
rect -774 6544 -740 6550
rect -774 6482 -740 6506
rect -774 6472 -740 6482
rect -774 6414 -740 6434
rect -774 6400 -740 6414
rect -774 6346 -740 6362
rect -774 6328 -740 6346
rect -774 6278 -740 6290
rect -774 6256 -740 6278
rect -774 6210 -740 6218
rect -774 6184 -740 6210
rect -774 6142 -740 6146
rect -774 6112 -740 6142
rect 890 6618 924 6650
rect 890 6616 924 6618
rect 890 6550 924 6578
rect 890 6544 924 6550
rect 890 6482 924 6506
rect 890 6472 924 6482
rect 890 6414 924 6434
rect 890 6400 924 6414
rect 890 6346 924 6362
rect 890 6328 924 6346
rect 890 6278 924 6290
rect 890 6256 924 6278
rect 890 6210 924 6218
rect 890 6184 924 6210
rect -774 6040 -740 6074
rect -774 5972 -740 6002
rect -774 5968 -740 5972
rect -774 5904 -740 5930
rect -774 5896 -740 5904
rect -774 5836 -740 5858
rect -774 5824 -740 5836
rect -774 5768 -740 5786
rect -774 5752 -740 5768
rect -774 5700 -740 5714
rect -774 5680 -740 5700
rect -774 5632 -740 5642
rect -774 5608 -740 5632
rect -774 5564 -740 5570
rect -774 5536 -740 5564
rect -774 5496 -740 5498
rect -774 5464 -740 5496
rect -774 5394 -740 5426
rect -774 5392 -740 5394
rect -774 5326 -740 5354
rect -774 5320 -740 5326
rect -774 5258 -740 5282
rect -774 5248 -740 5258
rect -774 5190 -740 5210
rect -774 5176 -740 5190
rect -774 5122 -740 5138
rect -774 5104 -740 5122
rect -774 5054 -740 5066
rect -774 5032 -740 5054
rect -774 4986 -740 4994
rect -774 4960 -740 4986
rect -774 4918 -740 4922
rect -774 4888 -740 4918
rect -774 4816 -740 4850
rect -774 4748 -740 4778
rect -774 4744 -740 4748
rect -774 4680 -740 4706
rect -774 4672 -740 4680
rect -774 4612 -740 4634
rect -774 4600 -740 4612
rect -774 4544 -740 4562
rect -774 4528 -740 4544
rect -774 4476 -740 4490
rect -774 4456 -740 4476
rect -774 4408 -740 4418
rect -774 4384 -740 4408
rect -774 4340 -740 4346
rect -774 4312 -740 4340
rect -774 4272 -740 4274
rect -774 4240 -740 4272
rect -774 4170 -740 4202
rect -774 4168 -740 4170
rect -774 4102 -740 4130
rect -774 4096 -740 4102
rect -774 4034 -740 4058
rect -774 4024 -740 4034
rect -774 3966 -740 3986
rect -774 3952 -740 3966
rect -774 3898 -740 3914
rect -774 3880 -740 3898
rect -774 3830 -740 3842
rect -774 3808 -740 3830
rect -774 3762 -740 3770
rect -774 3736 -740 3762
rect -774 3694 -740 3698
rect -774 3664 -740 3694
rect -774 3592 -740 3626
rect -774 3524 -740 3554
rect -774 3520 -740 3524
rect -774 3456 -740 3482
rect -774 3448 -740 3456
rect -774 3388 -740 3410
rect -774 3376 -740 3388
rect -774 3320 -740 3338
rect -774 3304 -740 3320
rect -774 3252 -740 3266
rect -774 3232 -740 3252
rect -774 3184 -740 3194
rect -774 3160 -740 3184
rect -774 3116 -740 3122
rect -774 3088 -740 3116
rect -774 3048 -740 3050
rect -774 3016 -740 3048
rect -774 2946 -740 2978
rect -774 2944 -740 2946
rect -774 2878 -740 2906
rect -774 2872 -740 2878
rect -774 2810 -740 2834
rect -774 2800 -740 2810
rect -774 2742 -740 2762
rect -774 2728 -740 2742
rect -774 2674 -740 2690
rect -774 2656 -740 2674
rect -774 2606 -740 2618
rect -774 2584 -740 2606
rect -774 2538 -740 2546
rect -774 2512 -740 2538
rect -774 2470 -740 2474
rect -774 2440 -740 2470
rect -774 2368 -740 2402
rect -774 2300 -740 2330
rect -774 2296 -740 2300
rect -774 2232 -740 2258
rect -774 2224 -740 2232
rect -774 2164 -740 2186
rect -774 2152 -740 2164
rect -774 2096 -740 2114
rect -774 2080 -740 2096
rect -774 2028 -740 2042
rect -774 2008 -740 2028
rect -774 1960 -740 1970
rect -774 1936 -740 1960
rect -774 1892 -740 1898
rect -774 1864 -740 1892
rect -774 1824 -740 1826
rect -774 1792 -740 1824
rect -774 1722 -740 1754
rect -774 1720 -740 1722
rect -774 1654 -740 1682
rect -774 1648 -740 1654
rect -774 1586 -740 1610
rect -774 1576 -740 1586
rect -774 1518 -740 1538
rect -774 1504 -740 1518
rect -774 1450 -740 1466
rect -774 1432 -740 1450
rect -774 1382 -740 1394
rect -774 1360 -740 1382
rect -774 1314 -740 1322
rect -774 1288 -740 1314
rect -774 1246 -740 1250
rect -774 1216 -740 1246
rect -774 1144 -740 1178
rect -774 1076 -740 1106
rect -774 1072 -740 1076
rect -774 1008 -740 1034
rect -774 1000 -740 1008
rect -774 940 -740 962
rect -774 928 -740 940
rect -774 872 -740 890
rect -774 856 -740 872
rect -774 804 -740 818
rect -774 784 -740 804
rect -774 736 -740 746
rect -774 712 -740 736
rect -774 668 -740 674
rect -774 640 -740 668
rect -774 600 -740 602
rect -774 568 -740 600
rect -774 498 -740 530
rect -774 496 -740 498
rect -774 430 -740 458
rect -774 424 -740 430
rect -774 362 -740 386
rect -774 352 -740 362
rect -774 294 -740 314
rect -774 280 -740 294
rect -774 226 -740 242
rect -774 208 -740 226
rect -774 158 -740 170
rect -774 136 -740 158
rect -774 90 -740 98
rect -774 64 -740 90
rect -774 22 -740 26
rect -774 -8 -740 22
rect -774 -80 -740 -46
rect -774 -148 -740 -118
rect -774 -152 -740 -148
rect -647 5971 -469 6146
rect -647 5937 -646 5971
rect -646 5937 -612 5971
rect -612 5937 -469 5971
rect -647 5903 -469 5937
rect -647 5869 -646 5903
rect -646 5869 -612 5903
rect -612 5869 -469 5903
rect -647 5835 -469 5869
rect -647 5801 -646 5835
rect -646 5801 -612 5835
rect -612 5801 -469 5835
rect -647 5767 -469 5801
rect -647 5733 -646 5767
rect -646 5733 -612 5767
rect -612 5733 -469 5767
rect -647 5699 -469 5733
rect -647 5665 -646 5699
rect -646 5665 -612 5699
rect -612 5665 -469 5699
rect -647 5631 -469 5665
rect -647 5597 -646 5631
rect -646 5597 -612 5631
rect -612 5597 -469 5631
rect -647 5563 -469 5597
rect -647 5529 -646 5563
rect -646 5529 -612 5563
rect -612 5529 -469 5563
rect -647 5495 -469 5529
rect -647 5461 -646 5495
rect -646 5461 -612 5495
rect -612 5461 -469 5495
rect -647 5427 -469 5461
rect -647 5393 -646 5427
rect -646 5393 -612 5427
rect -612 5393 -469 5427
rect -647 5359 -469 5393
rect -647 5325 -646 5359
rect -646 5325 -612 5359
rect -612 5325 -469 5359
rect -647 5291 -469 5325
rect -647 5257 -646 5291
rect -646 5257 -612 5291
rect -612 5257 -469 5291
rect -647 5223 -469 5257
rect -647 5189 -646 5223
rect -646 5189 -612 5223
rect -612 5189 -469 5223
rect -647 5155 -469 5189
rect -647 5121 -646 5155
rect -646 5121 -612 5155
rect -612 5121 -469 5155
rect -647 5087 -469 5121
rect -647 5053 -646 5087
rect -646 5053 -612 5087
rect -612 5053 -469 5087
rect -647 5019 -469 5053
rect -647 4985 -646 5019
rect -646 4985 -612 5019
rect -612 4985 -469 5019
rect -647 4951 -469 4985
rect -647 4917 -646 4951
rect -646 4917 -612 4951
rect -612 4917 -469 4951
rect -647 4883 -469 4917
rect -647 4849 -646 4883
rect -646 4849 -612 4883
rect -612 4849 -469 4883
rect -647 4815 -469 4849
rect -647 4781 -646 4815
rect -646 4781 -612 4815
rect -612 4781 -469 4815
rect -647 4747 -469 4781
rect -647 4713 -646 4747
rect -646 4713 -612 4747
rect -612 4713 -469 4747
rect -647 4679 -469 4713
rect -647 4645 -646 4679
rect -646 4645 -612 4679
rect -612 4645 -469 4679
rect -647 4611 -469 4645
rect -647 4577 -646 4611
rect -646 4577 -612 4611
rect -612 4577 -469 4611
rect -647 4543 -469 4577
rect -647 4509 -646 4543
rect -646 4509 -612 4543
rect -612 4509 -469 4543
rect -647 4475 -469 4509
rect -647 4441 -646 4475
rect -646 4441 -612 4475
rect -612 4441 -469 4475
rect -647 4407 -469 4441
rect -647 4373 -646 4407
rect -646 4373 -612 4407
rect -612 4373 -469 4407
rect -647 4339 -469 4373
rect -647 4305 -646 4339
rect -646 4305 -612 4339
rect -612 4305 -469 4339
rect -647 4271 -469 4305
rect -647 4237 -646 4271
rect -646 4237 -612 4271
rect -612 4237 -469 4271
rect -647 4203 -469 4237
rect -647 4169 -646 4203
rect -646 4169 -612 4203
rect -612 4169 -469 4203
rect -647 4135 -469 4169
rect -647 4101 -646 4135
rect -646 4101 -612 4135
rect -612 4101 -469 4135
rect -647 4067 -469 4101
rect -647 4033 -646 4067
rect -646 4033 -612 4067
rect -612 4033 -469 4067
rect -647 3999 -469 4033
rect -647 3965 -646 3999
rect -646 3965 -612 3999
rect -612 3965 -469 3999
rect -647 3931 -469 3965
rect -647 3897 -646 3931
rect -646 3897 -612 3931
rect -612 3897 -469 3931
rect -647 3863 -469 3897
rect -647 3829 -646 3863
rect -646 3829 -612 3863
rect -612 3829 -469 3863
rect -647 3795 -469 3829
rect -647 3761 -646 3795
rect -646 3761 -612 3795
rect -612 3761 -469 3795
rect -647 3727 -469 3761
rect -647 3693 -646 3727
rect -646 3693 -612 3727
rect -612 3693 -469 3727
rect -647 3659 -469 3693
rect -647 3625 -646 3659
rect -646 3625 -612 3659
rect -612 3625 -469 3659
rect -647 3591 -469 3625
rect -647 3557 -646 3591
rect -646 3557 -612 3591
rect -612 3557 -469 3591
rect -647 3523 -469 3557
rect -647 3489 -646 3523
rect -646 3489 -612 3523
rect -612 3489 -469 3523
rect -647 3455 -469 3489
rect -647 3421 -646 3455
rect -646 3421 -612 3455
rect -612 3421 -469 3455
rect -647 3387 -469 3421
rect -647 3353 -646 3387
rect -646 3353 -612 3387
rect -612 3353 -469 3387
rect -647 3319 -469 3353
rect -647 3285 -646 3319
rect -646 3285 -612 3319
rect -612 3285 -469 3319
rect -647 3251 -469 3285
rect -647 3217 -646 3251
rect -646 3217 -612 3251
rect -612 3217 -469 3251
rect -647 3183 -469 3217
rect -647 3149 -646 3183
rect -646 3149 -612 3183
rect -612 3149 -469 3183
rect -647 3115 -469 3149
rect -647 3081 -646 3115
rect -646 3081 -612 3115
rect -612 3081 -469 3115
rect -647 3047 -469 3081
rect -647 3013 -646 3047
rect -646 3013 -612 3047
rect -612 3013 -469 3047
rect -647 2979 -469 3013
rect -647 2945 -646 2979
rect -646 2945 -612 2979
rect -612 2945 -469 2979
rect -647 2911 -469 2945
rect -647 2877 -646 2911
rect -646 2877 -612 2911
rect -612 2877 -469 2911
rect -647 2843 -469 2877
rect -647 2809 -646 2843
rect -646 2809 -612 2843
rect -612 2809 -469 2843
rect -647 2775 -469 2809
rect -647 2741 -646 2775
rect -646 2741 -612 2775
rect -612 2741 -469 2775
rect -647 2707 -469 2741
rect -647 2673 -646 2707
rect -646 2673 -612 2707
rect -612 2673 -469 2707
rect -647 2639 -469 2673
rect -647 2605 -646 2639
rect -646 2605 -612 2639
rect -612 2605 -469 2639
rect -647 2571 -469 2605
rect -647 2537 -646 2571
rect -646 2537 -612 2571
rect -612 2537 -469 2571
rect -647 2503 -469 2537
rect -647 2469 -646 2503
rect -646 2469 -612 2503
rect -612 2469 -469 2503
rect -647 2435 -469 2469
rect -647 2401 -646 2435
rect -646 2401 -612 2435
rect -612 2401 -469 2435
rect -647 2367 -469 2401
rect -647 2333 -646 2367
rect -646 2333 -612 2367
rect -612 2333 -469 2367
rect -647 2299 -469 2333
rect -647 2265 -646 2299
rect -646 2265 -612 2299
rect -612 2265 -469 2299
rect -647 2231 -469 2265
rect -647 2197 -646 2231
rect -646 2197 -612 2231
rect -612 2197 -469 2231
rect -647 2163 -469 2197
rect -647 2129 -646 2163
rect -646 2129 -612 2163
rect -612 2129 -469 2163
rect -647 2095 -469 2129
rect -647 2061 -646 2095
rect -646 2061 -612 2095
rect -612 2061 -469 2095
rect -647 2027 -469 2061
rect -647 1993 -646 2027
rect -646 1993 -612 2027
rect -612 1993 -469 2027
rect -647 1959 -469 1993
rect -647 1925 -646 1959
rect -646 1925 -612 1959
rect -612 1925 -469 1959
rect -647 1891 -469 1925
rect -647 1857 -646 1891
rect -646 1857 -612 1891
rect -612 1857 -469 1891
rect -647 1823 -469 1857
rect -647 1789 -646 1823
rect -646 1789 -612 1823
rect -612 1789 -469 1823
rect -647 1755 -469 1789
rect -647 1721 -646 1755
rect -646 1721 -612 1755
rect -612 1721 -469 1755
rect -647 1687 -469 1721
rect -647 1653 -646 1687
rect -646 1653 -612 1687
rect -612 1653 -469 1687
rect -647 1619 -469 1653
rect -647 1585 -646 1619
rect -646 1585 -612 1619
rect -612 1585 -469 1619
rect -647 1551 -469 1585
rect -647 1517 -646 1551
rect -646 1517 -612 1551
rect -612 1517 -469 1551
rect -647 1483 -469 1517
rect -647 1449 -646 1483
rect -646 1449 -612 1483
rect -612 1449 -469 1483
rect -647 1415 -469 1449
rect -647 1381 -646 1415
rect -646 1381 -612 1415
rect -612 1381 -469 1415
rect -647 1347 -469 1381
rect -647 1313 -646 1347
rect -646 1313 -612 1347
rect -612 1313 -469 1347
rect -647 1279 -469 1313
rect -647 1245 -646 1279
rect -646 1245 -612 1279
rect -612 1245 -469 1279
rect -647 1211 -469 1245
rect -647 1177 -646 1211
rect -646 1177 -612 1211
rect -612 1177 -469 1211
rect -647 1143 -469 1177
rect -647 1109 -646 1143
rect -646 1109 -612 1143
rect -612 1109 -469 1143
rect -647 1075 -469 1109
rect -647 1041 -646 1075
rect -646 1041 -612 1075
rect -612 1041 -469 1075
rect -647 1007 -469 1041
rect -647 973 -646 1007
rect -646 973 -612 1007
rect -612 973 -469 1007
rect -647 939 -469 973
rect -647 905 -646 939
rect -646 905 -612 939
rect -612 905 -469 939
rect -647 871 -469 905
rect -647 837 -646 871
rect -646 837 -612 871
rect -612 837 -469 871
rect -647 803 -469 837
rect -647 769 -646 803
rect -646 769 -612 803
rect -612 769 -469 803
rect -647 735 -469 769
rect -647 701 -646 735
rect -646 701 -612 735
rect -612 701 -469 735
rect -647 667 -469 701
rect -647 633 -646 667
rect -646 633 -612 667
rect -612 633 -469 667
rect -647 599 -469 633
rect -647 565 -646 599
rect -646 565 -612 599
rect -612 565 -469 599
rect -647 531 -469 565
rect -647 497 -646 531
rect -646 497 -612 531
rect -612 497 -469 531
rect -647 463 -469 497
rect -647 429 -646 463
rect -646 429 -612 463
rect -612 429 -469 463
rect -647 395 -469 429
rect -647 361 -646 395
rect -646 361 -612 395
rect -612 361 -469 395
rect -647 327 -469 361
rect -647 293 -646 327
rect -646 293 -612 327
rect -612 293 -469 327
rect -647 259 -469 293
rect -647 225 -646 259
rect -646 225 -612 259
rect -612 225 -469 259
rect -647 191 -469 225
rect -647 157 -646 191
rect -646 157 -612 191
rect -612 157 -469 191
rect -647 123 -469 157
rect -647 89 -646 123
rect -646 89 -612 123
rect -612 89 -469 123
rect -647 55 -469 89
rect -647 21 -646 55
rect -646 21 -612 55
rect -612 21 -469 55
rect -647 -152 -469 21
rect -122 5939 272 6146
rect -122 57 24 5939
rect 24 57 126 5939
rect 126 57 272 5939
rect -122 -152 272 57
rect 619 5971 797 6146
rect 619 5937 762 5971
rect 762 5937 796 5971
rect 796 5937 797 5971
rect 619 5903 797 5937
rect 619 5869 762 5903
rect 762 5869 796 5903
rect 796 5869 797 5903
rect 619 5835 797 5869
rect 619 5801 762 5835
rect 762 5801 796 5835
rect 796 5801 797 5835
rect 619 5767 797 5801
rect 619 5733 762 5767
rect 762 5733 796 5767
rect 796 5733 797 5767
rect 619 5699 797 5733
rect 619 5665 762 5699
rect 762 5665 796 5699
rect 796 5665 797 5699
rect 619 5631 797 5665
rect 619 5597 762 5631
rect 762 5597 796 5631
rect 796 5597 797 5631
rect 619 5563 797 5597
rect 619 5529 762 5563
rect 762 5529 796 5563
rect 796 5529 797 5563
rect 619 5495 797 5529
rect 619 5461 762 5495
rect 762 5461 796 5495
rect 796 5461 797 5495
rect 619 5427 797 5461
rect 619 5393 762 5427
rect 762 5393 796 5427
rect 796 5393 797 5427
rect 619 5359 797 5393
rect 619 5325 762 5359
rect 762 5325 796 5359
rect 796 5325 797 5359
rect 619 5291 797 5325
rect 619 5257 762 5291
rect 762 5257 796 5291
rect 796 5257 797 5291
rect 619 5223 797 5257
rect 619 5189 762 5223
rect 762 5189 796 5223
rect 796 5189 797 5223
rect 619 5155 797 5189
rect 619 5121 762 5155
rect 762 5121 796 5155
rect 796 5121 797 5155
rect 619 5087 797 5121
rect 619 5053 762 5087
rect 762 5053 796 5087
rect 796 5053 797 5087
rect 619 5019 797 5053
rect 619 4985 762 5019
rect 762 4985 796 5019
rect 796 4985 797 5019
rect 619 4951 797 4985
rect 619 4917 762 4951
rect 762 4917 796 4951
rect 796 4917 797 4951
rect 619 4883 797 4917
rect 619 4849 762 4883
rect 762 4849 796 4883
rect 796 4849 797 4883
rect 619 4815 797 4849
rect 619 4781 762 4815
rect 762 4781 796 4815
rect 796 4781 797 4815
rect 619 4747 797 4781
rect 619 4713 762 4747
rect 762 4713 796 4747
rect 796 4713 797 4747
rect 619 4679 797 4713
rect 619 4645 762 4679
rect 762 4645 796 4679
rect 796 4645 797 4679
rect 619 4611 797 4645
rect 619 4577 762 4611
rect 762 4577 796 4611
rect 796 4577 797 4611
rect 619 4543 797 4577
rect 619 4509 762 4543
rect 762 4509 796 4543
rect 796 4509 797 4543
rect 619 4475 797 4509
rect 619 4441 762 4475
rect 762 4441 796 4475
rect 796 4441 797 4475
rect 619 4407 797 4441
rect 619 4373 762 4407
rect 762 4373 796 4407
rect 796 4373 797 4407
rect 619 4339 797 4373
rect 619 4305 762 4339
rect 762 4305 796 4339
rect 796 4305 797 4339
rect 619 4271 797 4305
rect 619 4237 762 4271
rect 762 4237 796 4271
rect 796 4237 797 4271
rect 619 4203 797 4237
rect 619 4169 762 4203
rect 762 4169 796 4203
rect 796 4169 797 4203
rect 619 4135 797 4169
rect 619 4101 762 4135
rect 762 4101 796 4135
rect 796 4101 797 4135
rect 619 4067 797 4101
rect 619 4033 762 4067
rect 762 4033 796 4067
rect 796 4033 797 4067
rect 619 3999 797 4033
rect 619 3965 762 3999
rect 762 3965 796 3999
rect 796 3965 797 3999
rect 619 3931 797 3965
rect 619 3897 762 3931
rect 762 3897 796 3931
rect 796 3897 797 3931
rect 619 3863 797 3897
rect 619 3829 762 3863
rect 762 3829 796 3863
rect 796 3829 797 3863
rect 619 3795 797 3829
rect 619 3761 762 3795
rect 762 3761 796 3795
rect 796 3761 797 3795
rect 619 3727 797 3761
rect 619 3693 762 3727
rect 762 3693 796 3727
rect 796 3693 797 3727
rect 619 3659 797 3693
rect 619 3625 762 3659
rect 762 3625 796 3659
rect 796 3625 797 3659
rect 619 3591 797 3625
rect 619 3557 762 3591
rect 762 3557 796 3591
rect 796 3557 797 3591
rect 619 3523 797 3557
rect 619 3489 762 3523
rect 762 3489 796 3523
rect 796 3489 797 3523
rect 619 3455 797 3489
rect 619 3421 762 3455
rect 762 3421 796 3455
rect 796 3421 797 3455
rect 619 3387 797 3421
rect 619 3353 762 3387
rect 762 3353 796 3387
rect 796 3353 797 3387
rect 619 3319 797 3353
rect 619 3285 762 3319
rect 762 3285 796 3319
rect 796 3285 797 3319
rect 619 3251 797 3285
rect 619 3217 762 3251
rect 762 3217 796 3251
rect 796 3217 797 3251
rect 619 3183 797 3217
rect 619 3149 762 3183
rect 762 3149 796 3183
rect 796 3149 797 3183
rect 619 3115 797 3149
rect 619 3081 762 3115
rect 762 3081 796 3115
rect 796 3081 797 3115
rect 619 3047 797 3081
rect 619 3013 762 3047
rect 762 3013 796 3047
rect 796 3013 797 3047
rect 619 2979 797 3013
rect 619 2945 762 2979
rect 762 2945 796 2979
rect 796 2945 797 2979
rect 619 2911 797 2945
rect 619 2877 762 2911
rect 762 2877 796 2911
rect 796 2877 797 2911
rect 619 2843 797 2877
rect 619 2809 762 2843
rect 762 2809 796 2843
rect 796 2809 797 2843
rect 619 2775 797 2809
rect 619 2741 762 2775
rect 762 2741 796 2775
rect 796 2741 797 2775
rect 619 2707 797 2741
rect 619 2673 762 2707
rect 762 2673 796 2707
rect 796 2673 797 2707
rect 619 2639 797 2673
rect 619 2605 762 2639
rect 762 2605 796 2639
rect 796 2605 797 2639
rect 619 2571 797 2605
rect 619 2537 762 2571
rect 762 2537 796 2571
rect 796 2537 797 2571
rect 619 2503 797 2537
rect 619 2469 762 2503
rect 762 2469 796 2503
rect 796 2469 797 2503
rect 619 2435 797 2469
rect 619 2401 762 2435
rect 762 2401 796 2435
rect 796 2401 797 2435
rect 619 2367 797 2401
rect 619 2333 762 2367
rect 762 2333 796 2367
rect 796 2333 797 2367
rect 619 2299 797 2333
rect 619 2265 762 2299
rect 762 2265 796 2299
rect 796 2265 797 2299
rect 619 2231 797 2265
rect 619 2197 762 2231
rect 762 2197 796 2231
rect 796 2197 797 2231
rect 619 2163 797 2197
rect 619 2129 762 2163
rect 762 2129 796 2163
rect 796 2129 797 2163
rect 619 2095 797 2129
rect 619 2061 762 2095
rect 762 2061 796 2095
rect 796 2061 797 2095
rect 619 2027 797 2061
rect 619 1993 762 2027
rect 762 1993 796 2027
rect 796 1993 797 2027
rect 619 1959 797 1993
rect 619 1925 762 1959
rect 762 1925 796 1959
rect 796 1925 797 1959
rect 619 1891 797 1925
rect 619 1857 762 1891
rect 762 1857 796 1891
rect 796 1857 797 1891
rect 619 1823 797 1857
rect 619 1789 762 1823
rect 762 1789 796 1823
rect 796 1789 797 1823
rect 619 1755 797 1789
rect 619 1721 762 1755
rect 762 1721 796 1755
rect 796 1721 797 1755
rect 619 1687 797 1721
rect 619 1653 762 1687
rect 762 1653 796 1687
rect 796 1653 797 1687
rect 619 1619 797 1653
rect 619 1585 762 1619
rect 762 1585 796 1619
rect 796 1585 797 1619
rect 619 1551 797 1585
rect 619 1517 762 1551
rect 762 1517 796 1551
rect 796 1517 797 1551
rect 619 1483 797 1517
rect 619 1449 762 1483
rect 762 1449 796 1483
rect 796 1449 797 1483
rect 619 1415 797 1449
rect 619 1381 762 1415
rect 762 1381 796 1415
rect 796 1381 797 1415
rect 619 1347 797 1381
rect 619 1313 762 1347
rect 762 1313 796 1347
rect 796 1313 797 1347
rect 619 1279 797 1313
rect 619 1245 762 1279
rect 762 1245 796 1279
rect 796 1245 797 1279
rect 619 1211 797 1245
rect 619 1177 762 1211
rect 762 1177 796 1211
rect 796 1177 797 1211
rect 619 1143 797 1177
rect 619 1109 762 1143
rect 762 1109 796 1143
rect 796 1109 797 1143
rect 619 1075 797 1109
rect 619 1041 762 1075
rect 762 1041 796 1075
rect 796 1041 797 1075
rect 619 1007 797 1041
rect 619 973 762 1007
rect 762 973 796 1007
rect 796 973 797 1007
rect 619 939 797 973
rect 619 905 762 939
rect 762 905 796 939
rect 796 905 797 939
rect 619 871 797 905
rect 619 837 762 871
rect 762 837 796 871
rect 796 837 797 871
rect 619 803 797 837
rect 619 769 762 803
rect 762 769 796 803
rect 796 769 797 803
rect 619 735 797 769
rect 619 701 762 735
rect 762 701 796 735
rect 796 701 797 735
rect 619 667 797 701
rect 619 633 762 667
rect 762 633 796 667
rect 796 633 797 667
rect 619 599 797 633
rect 619 565 762 599
rect 762 565 796 599
rect 796 565 797 599
rect 619 531 797 565
rect 619 497 762 531
rect 762 497 796 531
rect 796 497 797 531
rect 619 463 797 497
rect 619 429 762 463
rect 762 429 796 463
rect 796 429 797 463
rect 619 395 797 429
rect 619 361 762 395
rect 762 361 796 395
rect 796 361 797 395
rect 619 327 797 361
rect 619 293 762 327
rect 762 293 796 327
rect 796 293 797 327
rect 619 259 797 293
rect 619 225 762 259
rect 762 225 796 259
rect 796 225 797 259
rect 619 191 797 225
rect 619 157 762 191
rect 762 157 796 191
rect 796 157 797 191
rect 619 123 797 157
rect 619 89 762 123
rect 762 89 796 123
rect 796 89 797 123
rect 619 55 797 89
rect 619 21 762 55
rect 762 21 796 55
rect 796 21 797 55
rect 619 -152 797 21
rect 890 6142 924 6146
rect 890 6112 924 6142
rect 890 6040 924 6074
rect 890 5972 924 6002
rect 890 5968 924 5972
rect 890 5904 924 5930
rect 890 5896 924 5904
rect 890 5836 924 5858
rect 890 5824 924 5836
rect 890 5768 924 5786
rect 890 5752 924 5768
rect 890 5700 924 5714
rect 890 5680 924 5700
rect 890 5632 924 5642
rect 890 5608 924 5632
rect 890 5564 924 5570
rect 890 5536 924 5564
rect 890 5496 924 5498
rect 890 5464 924 5496
rect 890 5394 924 5426
rect 890 5392 924 5394
rect 890 5326 924 5354
rect 890 5320 924 5326
rect 890 5258 924 5282
rect 890 5248 924 5258
rect 890 5190 924 5210
rect 890 5176 924 5190
rect 890 5122 924 5138
rect 890 5104 924 5122
rect 890 5054 924 5066
rect 890 5032 924 5054
rect 890 4986 924 4994
rect 890 4960 924 4986
rect 890 4918 924 4922
rect 890 4888 924 4918
rect 890 4816 924 4850
rect 890 4748 924 4778
rect 890 4744 924 4748
rect 890 4680 924 4706
rect 890 4672 924 4680
rect 890 4612 924 4634
rect 890 4600 924 4612
rect 890 4544 924 4562
rect 890 4528 924 4544
rect 890 4476 924 4490
rect 890 4456 924 4476
rect 890 4408 924 4418
rect 890 4384 924 4408
rect 890 4340 924 4346
rect 890 4312 924 4340
rect 890 4272 924 4274
rect 890 4240 924 4272
rect 890 4170 924 4202
rect 890 4168 924 4170
rect 890 4102 924 4130
rect 890 4096 924 4102
rect 890 4034 924 4058
rect 890 4024 924 4034
rect 890 3966 924 3986
rect 890 3952 924 3966
rect 890 3898 924 3914
rect 890 3880 924 3898
rect 890 3830 924 3842
rect 890 3808 924 3830
rect 890 3762 924 3770
rect 890 3736 924 3762
rect 890 3694 924 3698
rect 890 3664 924 3694
rect 890 3592 924 3626
rect 890 3524 924 3554
rect 890 3520 924 3524
rect 890 3456 924 3482
rect 890 3448 924 3456
rect 890 3388 924 3410
rect 890 3376 924 3388
rect 890 3320 924 3338
rect 890 3304 924 3320
rect 890 3252 924 3266
rect 890 3232 924 3252
rect 890 3184 924 3194
rect 890 3160 924 3184
rect 890 3116 924 3122
rect 890 3088 924 3116
rect 890 3048 924 3050
rect 890 3016 924 3048
rect 890 2946 924 2978
rect 890 2944 924 2946
rect 890 2878 924 2906
rect 890 2872 924 2878
rect 890 2810 924 2834
rect 890 2800 924 2810
rect 890 2742 924 2762
rect 890 2728 924 2742
rect 890 2674 924 2690
rect 890 2656 924 2674
rect 890 2606 924 2618
rect 890 2584 924 2606
rect 890 2538 924 2546
rect 890 2512 924 2538
rect 890 2470 924 2474
rect 890 2440 924 2470
rect 890 2368 924 2402
rect 890 2300 924 2330
rect 890 2296 924 2300
rect 890 2232 924 2258
rect 890 2224 924 2232
rect 890 2164 924 2186
rect 890 2152 924 2164
rect 890 2096 924 2114
rect 890 2080 924 2096
rect 890 2028 924 2042
rect 890 2008 924 2028
rect 890 1960 924 1970
rect 890 1936 924 1960
rect 890 1892 924 1898
rect 890 1864 924 1892
rect 890 1824 924 1826
rect 890 1792 924 1824
rect 890 1722 924 1754
rect 890 1720 924 1722
rect 890 1654 924 1682
rect 890 1648 924 1654
rect 890 1586 924 1610
rect 890 1576 924 1586
rect 890 1518 924 1538
rect 890 1504 924 1518
rect 890 1450 924 1466
rect 890 1432 924 1450
rect 890 1382 924 1394
rect 890 1360 924 1382
rect 890 1314 924 1322
rect 890 1288 924 1314
rect 890 1246 924 1250
rect 890 1216 924 1246
rect 890 1144 924 1178
rect 890 1076 924 1106
rect 890 1072 924 1076
rect 890 1008 924 1034
rect 890 1000 924 1008
rect 890 940 924 962
rect 890 928 924 940
rect 890 872 924 890
rect 890 856 924 872
rect 890 804 924 818
rect 890 784 924 804
rect 890 736 924 746
rect 890 712 924 736
rect 890 668 924 674
rect 890 640 924 668
rect 890 600 924 602
rect 890 568 924 600
rect 890 498 924 530
rect 890 496 924 498
rect 890 430 924 458
rect 890 424 924 430
rect 890 362 924 386
rect 890 352 924 362
rect 890 294 924 314
rect 890 280 924 294
rect 890 226 924 242
rect 890 208 924 226
rect 890 158 924 170
rect 890 136 924 158
rect 890 90 924 98
rect 890 64 924 90
rect 890 22 924 26
rect 890 -8 924 22
rect 890 -80 924 -46
rect -774 -216 -740 -190
rect -774 -224 -740 -216
rect -774 -284 -740 -262
rect -774 -296 -740 -284
rect -774 -352 -740 -334
rect -774 -368 -740 -352
rect -774 -420 -740 -406
rect -774 -440 -740 -420
rect 890 -148 924 -118
rect 890 -152 924 -148
rect 890 -216 924 -190
rect 890 -224 924 -216
rect 890 -284 924 -262
rect 890 -296 924 -284
rect 890 -352 924 -334
rect 890 -368 924 -352
rect -774 -488 -740 -478
rect -774 -512 -740 -488
rect -774 -556 -740 -550
rect -774 -584 -740 -556
rect -774 -624 -740 -622
rect -774 -656 -740 -624
rect -130 -493 -96 -459
rect -56 -493 -22 -459
rect 18 -493 52 -459
rect 92 -493 126 -459
rect 166 -493 200 -459
rect 240 -493 274 -459
rect -130 -567 -96 -533
rect -56 -567 -22 -533
rect 18 -567 52 -533
rect 92 -567 126 -533
rect 166 -567 200 -533
rect 240 -567 274 -533
rect -130 -641 -96 -607
rect -56 -641 -22 -607
rect 18 -641 52 -607
rect 92 -641 126 -607
rect 166 -641 200 -607
rect 240 -641 274 -607
rect 890 -420 924 -406
rect 890 -440 924 -420
rect 890 -488 924 -478
rect 890 -512 924 -488
rect 890 -556 924 -550
rect 890 -584 924 -556
rect 890 -624 924 -622
rect 890 -656 924 -624
rect -554 -964 704 -820
rect -554 -998 -520 -964
rect -520 -998 -486 -964
rect -486 -998 -452 -964
rect -452 -998 -418 -964
rect -418 -998 -384 -964
rect -384 -998 -350 -964
rect -350 -998 -316 -964
rect -316 -998 -282 -964
rect -282 -998 -248 -964
rect -248 -998 -214 -964
rect -214 -998 -180 -964
rect -180 -998 -146 -964
rect -146 -998 -112 -964
rect -112 -998 -78 -964
rect -78 -998 -44 -964
rect -44 -998 -10 -964
rect -10 -998 24 -964
rect 24 -998 58 -964
rect 58 -998 92 -964
rect 92 -998 126 -964
rect 126 -998 160 -964
rect 160 -998 194 -964
rect 194 -998 228 -964
rect 228 -998 262 -964
rect 262 -998 296 -964
rect 296 -998 330 -964
rect 330 -998 364 -964
rect 364 -998 398 -964
rect 398 -998 432 -964
rect 432 -998 466 -964
rect 466 -998 500 -964
rect 500 -998 534 -964
rect 534 -998 568 -964
rect 568 -998 602 -964
rect 602 -998 636 -964
rect 636 -998 670 -964
rect 670 -998 704 -964
rect 1672 6992 1706 7013
rect 1672 6979 1706 6992
rect 1672 6924 1706 6941
rect 1672 6907 1706 6924
rect 1672 6856 1706 6869
rect 1672 6835 1706 6856
rect 1672 6788 1706 6797
rect 1672 6763 1706 6788
rect 1672 6720 1706 6725
rect 1672 6691 1706 6720
rect 1672 6652 1706 6653
rect 1672 6619 1706 6652
rect 1672 6550 1706 6581
rect 1672 6547 1706 6550
rect 1672 6482 1706 6509
rect 1672 6475 1706 6482
rect 1672 6414 1706 6437
rect 1672 6403 1706 6414
rect 1672 6346 1706 6365
rect 1672 6331 1706 6346
rect 1672 6278 1706 6293
rect 1672 6259 1706 6278
rect 1672 6210 1706 6221
rect 1672 6187 1706 6210
rect 1672 6142 1706 6149
rect 1672 6115 1706 6142
rect 1672 6074 1706 6077
rect 1672 6043 1706 6074
rect 1672 5972 1706 6005
rect 1672 5971 1706 5972
rect 1672 5904 1706 5933
rect 1672 5899 1706 5904
rect 1672 5836 1706 5861
rect 1672 5827 1706 5836
rect 1672 5768 1706 5789
rect 1672 5755 1706 5768
rect 1672 5700 1706 5717
rect 1672 5683 1706 5700
rect 1672 5632 1706 5645
rect 1672 5611 1706 5632
rect 1672 5564 1706 5573
rect 1672 5539 1706 5564
rect 1672 5496 1706 5501
rect 1672 5467 1706 5496
rect 1672 5428 1706 5429
rect 1672 5395 1706 5428
rect 1672 5326 1706 5357
rect 1672 5323 1706 5326
rect 1672 5258 1706 5285
rect 1672 5251 1706 5258
rect 1672 5190 1706 5213
rect 1672 5179 1706 5190
rect 1672 5122 1706 5141
rect 1672 5107 1706 5122
rect 1672 5054 1706 5069
rect 1672 5035 1706 5054
rect 1672 4986 1706 4997
rect 1672 4963 1706 4986
rect 1672 4918 1706 4925
rect 1672 4891 1706 4918
rect 1672 4850 1706 4853
rect 1672 4819 1706 4850
rect 1672 4748 1706 4781
rect 1672 4747 1706 4748
rect 1672 4680 1706 4709
rect 1672 4675 1706 4680
rect 1672 4612 1706 4637
rect 1672 4603 1706 4612
rect 1672 4544 1706 4565
rect 1672 4531 1706 4544
rect 1672 4476 1706 4493
rect 1672 4459 1706 4476
rect 1672 4408 1706 4421
rect 1672 4387 1706 4408
rect 1672 4340 1706 4349
rect 1672 4315 1706 4340
rect 1672 4272 1706 4277
rect 1672 4243 1706 4272
rect 1672 4204 1706 4205
rect 1672 4171 1706 4204
rect 1672 4102 1706 4133
rect 1672 4099 1706 4102
rect 1672 4034 1706 4061
rect 1672 4027 1706 4034
rect 1672 3966 1706 3989
rect 1672 3955 1706 3966
rect 1672 3898 1706 3917
rect 1672 3883 1706 3898
rect 1672 3830 1706 3845
rect 1672 3811 1706 3830
rect 1672 3762 1706 3773
rect 1672 3739 1706 3762
rect 1672 3694 1706 3701
rect 1672 3667 1706 3694
rect 1672 3626 1706 3629
rect 1672 3595 1706 3626
rect 1672 3524 1706 3557
rect 1672 3523 1706 3524
rect 1672 3456 1706 3485
rect 1672 3451 1706 3456
rect 1672 3388 1706 3413
rect 1672 3379 1706 3388
rect 1672 3320 1706 3341
rect 1672 3307 1706 3320
rect 1672 3252 1706 3269
rect 1672 3235 1706 3252
rect 1672 3184 1706 3197
rect 1672 3163 1706 3184
rect 1672 3116 1706 3125
rect 1672 3091 1706 3116
rect 1672 3048 1706 3053
rect 1672 3019 1706 3048
rect 1672 2980 1706 2981
rect 1672 2947 1706 2980
rect 1672 2878 1706 2909
rect 1672 2875 1706 2878
rect 1672 2810 1706 2837
rect 1672 2803 1706 2810
rect 1672 2742 1706 2765
rect 1672 2731 1706 2742
rect 1672 2674 1706 2693
rect 1672 2659 1706 2674
rect 1672 2606 1706 2621
rect 1672 2587 1706 2606
rect 1672 2538 1706 2549
rect 1672 2515 1706 2538
rect 1672 2470 1706 2477
rect 1672 2443 1706 2470
rect 1672 2402 1706 2405
rect 1672 2371 1706 2402
rect 1672 2300 1706 2333
rect 1672 2299 1706 2300
rect 1672 2232 1706 2261
rect 1672 2227 1706 2232
rect 1672 2164 1706 2189
rect 1672 2155 1706 2164
rect 1672 2096 1706 2117
rect 1672 2083 1706 2096
rect 1672 2028 1706 2045
rect 1672 2011 1706 2028
rect 1672 1960 1706 1973
rect 1672 1939 1706 1960
rect 1672 1892 1706 1901
rect 1672 1867 1706 1892
rect 1672 1824 1706 1829
rect 1672 1795 1706 1824
rect 1672 1756 1706 1757
rect 1672 1723 1706 1756
rect 1672 1654 1706 1685
rect 1672 1651 1706 1654
rect 1672 1586 1706 1613
rect 1672 1579 1706 1586
rect 1672 1518 1706 1541
rect 1672 1507 1706 1518
rect 1672 1450 1706 1469
rect 1672 1435 1706 1450
rect 1672 1382 1706 1397
rect 1672 1363 1706 1382
rect 1672 1314 1706 1325
rect 1672 1291 1706 1314
rect 1672 1246 1706 1253
rect 1672 1219 1706 1246
rect 1672 1178 1706 1181
rect 1672 1147 1706 1178
rect 1672 1076 1706 1109
rect 1672 1075 1706 1076
rect 1672 1008 1706 1037
rect 1672 1003 1706 1008
rect 1672 940 1706 965
rect 1672 931 1706 940
rect 1672 872 1706 893
rect 1672 859 1706 872
rect 1672 804 1706 821
rect 1672 787 1706 804
rect 1672 736 1706 749
rect 1672 715 1706 736
rect 1672 668 1706 677
rect 1672 643 1706 668
rect 1672 600 1706 605
rect 1672 571 1706 600
rect 1672 532 1706 533
rect 1672 499 1706 532
rect 1672 430 1706 461
rect 1672 427 1706 430
rect 1672 362 1706 389
rect 1672 355 1706 362
rect 1672 294 1706 317
rect 1672 283 1706 294
rect 1672 226 1706 245
rect 1672 211 1706 226
rect 1672 158 1706 173
rect 1672 139 1706 158
rect 1672 90 1706 101
rect 1672 67 1706 90
rect 1672 22 1706 29
rect 1672 -5 1706 22
rect 1672 -46 1706 -43
rect 1672 -77 1706 -46
rect 1672 -148 1706 -115
rect 1672 -149 1706 -148
rect 1672 -216 1706 -187
rect 1672 -221 1706 -216
rect 1672 -284 1706 -259
rect 1672 -293 1706 -284
rect 1672 -352 1706 -331
rect 1672 -365 1706 -352
rect 1672 -420 1706 -403
rect 1672 -437 1706 -420
rect 1672 -488 1706 -475
rect 1672 -509 1706 -488
rect 1672 -556 1706 -547
rect 1672 -581 1706 -556
rect 1672 -624 1706 -619
rect 1672 -653 1706 -624
rect 1672 -692 1706 -691
rect 1672 -725 1706 -692
rect 1672 -794 1706 -763
rect 1672 -797 1706 -794
rect 1672 -862 1706 -835
rect 1672 -869 1706 -862
rect 1672 -930 1706 -907
rect 1672 -941 1706 -930
rect 1672 -998 1706 -979
rect 1672 -1013 1706 -998
rect -1556 -1066 -1522 -1051
rect -1556 -1085 -1522 -1066
rect -1556 -1134 -1522 -1123
rect -1556 -1157 -1522 -1134
rect -1556 -1202 -1522 -1195
rect -1556 -1229 -1522 -1202
rect -1556 -1270 -1522 -1267
rect -1556 -1301 -1522 -1270
rect -1556 -1372 -1522 -1339
rect -1556 -1373 -1522 -1372
rect -1556 -1440 -1522 -1411
rect -1556 -1445 -1522 -1440
rect -1556 -1508 -1522 -1483
rect -1556 -1517 -1522 -1508
rect -1556 -1576 -1522 -1555
rect -1556 -1589 -1522 -1576
rect -1556 -1644 -1522 -1627
rect -1556 -1661 -1522 -1644
rect 1672 -1066 1706 -1051
rect 1672 -1085 1706 -1066
rect 1672 -1134 1706 -1123
rect 1672 -1157 1706 -1134
rect 1672 -1202 1706 -1195
rect 1672 -1229 1706 -1202
rect 1672 -1270 1706 -1267
rect 1672 -1301 1706 -1270
rect 1672 -1372 1706 -1339
rect 1672 -1373 1706 -1372
rect 1672 -1440 1706 -1411
rect 1672 -1445 1706 -1440
rect 1672 -1508 1706 -1483
rect 1672 -1517 1706 -1508
rect 1672 -1576 1706 -1555
rect 1672 -1589 1706 -1576
rect 1672 -1644 1706 -1627
rect 1672 -1661 1706 -1644
rect -1454 -1780 -1438 -1746
rect -1438 -1780 -1420 -1746
rect -1382 -1780 -1370 -1746
rect -1370 -1780 -1348 -1746
rect -1310 -1780 -1302 -1746
rect -1302 -1780 -1276 -1746
rect -1238 -1780 -1234 -1746
rect -1234 -1780 -1204 -1746
rect -1166 -1780 -1132 -1746
rect -1094 -1780 -1064 -1746
rect -1064 -1780 -1060 -1746
rect -1022 -1780 -996 -1746
rect -996 -1780 -988 -1746
rect -950 -1780 -928 -1746
rect -928 -1780 -916 -1746
rect -878 -1780 -860 -1746
rect -860 -1780 -844 -1746
rect -806 -1780 -792 -1746
rect -792 -1780 -772 -1746
rect -734 -1780 -724 -1746
rect -724 -1780 -700 -1746
rect -662 -1780 -656 -1746
rect -656 -1780 -628 -1746
rect -590 -1780 -588 -1746
rect -588 -1780 -556 -1746
rect -518 -1780 -486 -1746
rect -486 -1780 -484 -1746
rect -446 -1780 -418 -1746
rect -418 -1780 -412 -1746
rect -374 -1780 -350 -1746
rect -350 -1780 -340 -1746
rect -302 -1780 -282 -1746
rect -282 -1780 -268 -1746
rect -230 -1780 -214 -1746
rect -214 -1780 -196 -1746
rect -158 -1780 -146 -1746
rect -146 -1780 -124 -1746
rect -86 -1780 -78 -1746
rect -78 -1780 -52 -1746
rect -14 -1780 -10 -1746
rect -10 -1780 20 -1746
rect 58 -1780 92 -1746
rect 130 -1780 160 -1746
rect 160 -1780 164 -1746
rect 202 -1780 228 -1746
rect 228 -1780 236 -1746
rect 274 -1780 296 -1746
rect 296 -1780 308 -1746
rect 346 -1780 364 -1746
rect 364 -1780 380 -1746
rect 418 -1780 432 -1746
rect 432 -1780 452 -1746
rect 490 -1780 500 -1746
rect 500 -1780 524 -1746
rect 562 -1780 568 -1746
rect 568 -1780 596 -1746
rect 634 -1780 636 -1746
rect 636 -1780 668 -1746
rect 706 -1780 738 -1746
rect 738 -1780 740 -1746
rect 778 -1780 806 -1746
rect 806 -1780 812 -1746
rect 850 -1780 874 -1746
rect 874 -1780 884 -1746
rect 922 -1780 942 -1746
rect 942 -1780 956 -1746
rect 994 -1780 1010 -1746
rect 1010 -1780 1028 -1746
rect 1066 -1780 1078 -1746
rect 1078 -1780 1100 -1746
rect 1138 -1780 1146 -1746
rect 1146 -1780 1172 -1746
rect 1210 -1780 1214 -1746
rect 1214 -1780 1244 -1746
rect 1282 -1780 1316 -1746
rect 1354 -1780 1384 -1746
rect 1384 -1780 1388 -1746
rect 1426 -1780 1452 -1746
rect 1452 -1780 1460 -1746
rect 1498 -1780 1520 -1746
rect 1520 -1780 1532 -1746
rect 1570 -1780 1588 -1746
rect 1588 -1780 1604 -1746
<< metal1 >>
rect -1580 7780 1730 7804
rect -1580 7746 -1454 7780
rect -1420 7746 -1382 7780
rect -1348 7746 -1310 7780
rect -1276 7746 -1238 7780
rect -1204 7746 -1166 7780
rect -1132 7746 -1094 7780
rect -1060 7746 -1022 7780
rect -988 7746 -950 7780
rect -916 7746 -878 7780
rect -844 7746 -806 7780
rect -772 7746 -734 7780
rect -700 7746 -662 7780
rect -628 7746 -590 7780
rect -556 7746 -518 7780
rect -484 7746 -446 7780
rect -412 7746 -374 7780
rect -340 7746 -302 7780
rect -268 7746 -230 7780
rect -196 7746 -158 7780
rect -124 7746 -86 7780
rect -52 7746 -14 7780
rect 20 7746 58 7780
rect 92 7746 130 7780
rect 164 7746 202 7780
rect 236 7746 274 7780
rect 308 7746 346 7780
rect 380 7746 418 7780
rect 452 7746 490 7780
rect 524 7746 562 7780
rect 596 7746 634 7780
rect 668 7746 706 7780
rect 740 7746 778 7780
rect 812 7746 850 7780
rect 884 7746 922 7780
rect 956 7746 994 7780
rect 1028 7746 1066 7780
rect 1100 7746 1138 7780
rect 1172 7746 1210 7780
rect 1244 7746 1282 7780
rect 1316 7746 1354 7780
rect 1388 7746 1426 7780
rect 1460 7746 1498 7780
rect 1532 7746 1570 7780
rect 1604 7746 1730 7780
rect -1580 7722 1730 7746
rect -1580 7661 -1498 7722
rect -1580 7627 -1556 7661
rect -1522 7627 -1498 7661
rect -1580 7589 -1498 7627
rect -1580 7555 -1556 7589
rect -1522 7555 -1498 7589
rect -1580 7517 -1498 7555
rect -1580 7483 -1556 7517
rect -1522 7483 -1498 7517
rect -1580 7445 -1498 7483
rect -1580 7411 -1556 7445
rect -1522 7411 -1498 7445
rect -1580 7373 -1498 7411
rect -1580 7339 -1556 7373
rect -1522 7339 -1498 7373
rect -1580 7301 -1498 7339
rect -1580 7267 -1556 7301
rect -1522 7267 -1498 7301
rect -1580 7229 -1498 7267
rect -1580 7195 -1556 7229
rect -1522 7195 -1498 7229
rect -1580 7157 -1498 7195
rect -1580 7123 -1556 7157
rect -1522 7123 -1498 7157
rect -1580 7085 -1498 7123
rect -1580 7051 -1556 7085
rect -1522 7051 -1498 7085
rect -1580 7013 -1498 7051
rect 1648 7661 1730 7722
rect 1648 7627 1672 7661
rect 1706 7627 1730 7661
rect 1648 7589 1730 7627
rect 1648 7555 1672 7589
rect 1706 7555 1730 7589
rect 1648 7517 1730 7555
rect 1648 7483 1672 7517
rect 1706 7483 1730 7517
rect 1648 7445 1730 7483
rect 1648 7411 1672 7445
rect 1706 7411 1730 7445
rect 1648 7373 1730 7411
rect 1648 7339 1672 7373
rect 1706 7339 1730 7373
rect 1648 7301 1730 7339
rect 1648 7267 1672 7301
rect 1706 7267 1730 7301
rect 1648 7229 1730 7267
rect 1648 7195 1672 7229
rect 1706 7195 1730 7229
rect 1648 7157 1730 7195
rect 1648 7123 1672 7157
rect 1706 7123 1730 7157
rect 1648 7085 1730 7123
rect 1648 7051 1672 7085
rect 1706 7051 1730 7085
rect -1580 6979 -1556 7013
rect -1522 6979 -1498 7013
rect -1580 6941 -1498 6979
rect -1580 6907 -1556 6941
rect -1522 6907 -1498 6941
rect -1580 6869 -1498 6907
rect -1580 6835 -1556 6869
rect -1522 6835 -1498 6869
rect -1580 6797 -1498 6835
rect -1580 6763 -1556 6797
rect -1522 6763 -1498 6797
rect -1580 6725 -1498 6763
rect -1580 6691 -1556 6725
rect -1522 6691 -1498 6725
rect -1580 6653 -1498 6691
rect -1580 6619 -1556 6653
rect -1522 6619 -1498 6653
rect -1580 6581 -1498 6619
rect -1580 6547 -1556 6581
rect -1522 6547 -1498 6581
rect -1580 6509 -1498 6547
rect -1580 6475 -1556 6509
rect -1522 6475 -1498 6509
rect -1580 6437 -1498 6475
rect -1580 6403 -1556 6437
rect -1522 6403 -1498 6437
rect -1580 6365 -1498 6403
rect -1580 6331 -1556 6365
rect -1522 6331 -1498 6365
rect -1580 6293 -1498 6331
rect -1580 6259 -1556 6293
rect -1522 6259 -1498 6293
rect -1580 6221 -1498 6259
rect -1580 6187 -1556 6221
rect -1522 6187 -1498 6221
rect -1580 6149 -1498 6187
rect -1580 6115 -1556 6149
rect -1522 6115 -1498 6149
rect -1580 6077 -1498 6115
rect -1580 6043 -1556 6077
rect -1522 6043 -1498 6077
rect -1580 6005 -1498 6043
rect -1580 5971 -1556 6005
rect -1522 5971 -1498 6005
rect -1580 5933 -1498 5971
rect -1580 5899 -1556 5933
rect -1522 5899 -1498 5933
rect -1580 5861 -1498 5899
rect -1580 5827 -1556 5861
rect -1522 5827 -1498 5861
rect -1580 5789 -1498 5827
rect -1580 5755 -1556 5789
rect -1522 5755 -1498 5789
rect -1580 5717 -1498 5755
rect -1580 5683 -1556 5717
rect -1522 5683 -1498 5717
rect -1580 5645 -1498 5683
rect -1580 5611 -1556 5645
rect -1522 5611 -1498 5645
rect -1580 5573 -1498 5611
rect -1580 5539 -1556 5573
rect -1522 5539 -1498 5573
rect -1580 5501 -1498 5539
rect -1580 5467 -1556 5501
rect -1522 5467 -1498 5501
rect -1580 5429 -1498 5467
rect -1580 5395 -1556 5429
rect -1522 5395 -1498 5429
rect -1580 5357 -1498 5395
rect -1580 5323 -1556 5357
rect -1522 5323 -1498 5357
rect -1580 5285 -1498 5323
rect -1580 5251 -1556 5285
rect -1522 5251 -1498 5285
rect -1580 5213 -1498 5251
rect -1580 5179 -1556 5213
rect -1522 5179 -1498 5213
rect -1580 5141 -1498 5179
rect -1580 5107 -1556 5141
rect -1522 5107 -1498 5141
rect -1580 5069 -1498 5107
rect -1580 5035 -1556 5069
rect -1522 5035 -1498 5069
rect -1580 4997 -1498 5035
rect -1580 4963 -1556 4997
rect -1522 4963 -1498 4997
rect -1580 4925 -1498 4963
rect -1580 4891 -1556 4925
rect -1522 4891 -1498 4925
rect -1580 4853 -1498 4891
rect -1580 4819 -1556 4853
rect -1522 4819 -1498 4853
rect -1580 4781 -1498 4819
rect -1580 4747 -1556 4781
rect -1522 4747 -1498 4781
rect -1580 4709 -1498 4747
rect -1580 4675 -1556 4709
rect -1522 4675 -1498 4709
rect -1580 4637 -1498 4675
rect -1580 4603 -1556 4637
rect -1522 4603 -1498 4637
rect -1580 4565 -1498 4603
rect -1580 4531 -1556 4565
rect -1522 4531 -1498 4565
rect -1580 4493 -1498 4531
rect -1580 4459 -1556 4493
rect -1522 4459 -1498 4493
rect -1580 4421 -1498 4459
rect -1580 4387 -1556 4421
rect -1522 4387 -1498 4421
rect -1580 4349 -1498 4387
rect -1580 4315 -1556 4349
rect -1522 4315 -1498 4349
rect -1580 4277 -1498 4315
rect -1580 4243 -1556 4277
rect -1522 4243 -1498 4277
rect -1580 4205 -1498 4243
rect -1580 4171 -1556 4205
rect -1522 4171 -1498 4205
rect -1580 4133 -1498 4171
rect -1580 4099 -1556 4133
rect -1522 4099 -1498 4133
rect -1580 4061 -1498 4099
rect -1580 4027 -1556 4061
rect -1522 4027 -1498 4061
rect -1580 3989 -1498 4027
rect -1580 3955 -1556 3989
rect -1522 3955 -1498 3989
rect -1580 3917 -1498 3955
rect -1580 3883 -1556 3917
rect -1522 3883 -1498 3917
rect -1580 3845 -1498 3883
rect -1580 3811 -1556 3845
rect -1522 3811 -1498 3845
rect -1580 3773 -1498 3811
rect -1580 3739 -1556 3773
rect -1522 3739 -1498 3773
rect -1580 3701 -1498 3739
rect -1580 3667 -1556 3701
rect -1522 3667 -1498 3701
rect -1580 3629 -1498 3667
rect -1580 3595 -1556 3629
rect -1522 3595 -1498 3629
rect -1580 3557 -1498 3595
rect -1580 3523 -1556 3557
rect -1522 3523 -1498 3557
rect -1580 3485 -1498 3523
rect -1580 3451 -1556 3485
rect -1522 3451 -1498 3485
rect -1580 3413 -1498 3451
rect -1580 3379 -1556 3413
rect -1522 3379 -1498 3413
rect -1580 3341 -1498 3379
rect -1580 3307 -1556 3341
rect -1522 3307 -1498 3341
rect -1580 3269 -1498 3307
rect -1580 3235 -1556 3269
rect -1522 3235 -1498 3269
rect -1580 3197 -1498 3235
rect -1580 3163 -1556 3197
rect -1522 3163 -1498 3197
rect -1580 3125 -1498 3163
rect -1580 3091 -1556 3125
rect -1522 3091 -1498 3125
rect -1580 3053 -1498 3091
rect -1580 3019 -1556 3053
rect -1522 3019 -1498 3053
rect -1580 2981 -1498 3019
rect -1580 2947 -1556 2981
rect -1522 2947 -1498 2981
rect -1580 2909 -1498 2947
rect -1580 2875 -1556 2909
rect -1522 2875 -1498 2909
rect -1580 2837 -1498 2875
rect -1580 2803 -1556 2837
rect -1522 2803 -1498 2837
rect -1580 2765 -1498 2803
rect -1580 2731 -1556 2765
rect -1522 2731 -1498 2765
rect -1580 2693 -1498 2731
rect -1580 2659 -1556 2693
rect -1522 2659 -1498 2693
rect -1580 2621 -1498 2659
rect -1580 2587 -1556 2621
rect -1522 2587 -1498 2621
rect -1580 2549 -1498 2587
rect -1580 2515 -1556 2549
rect -1522 2515 -1498 2549
rect -1580 2477 -1498 2515
rect -1580 2443 -1556 2477
rect -1522 2443 -1498 2477
rect -1580 2405 -1498 2443
rect -1580 2371 -1556 2405
rect -1522 2371 -1498 2405
rect -1580 2333 -1498 2371
rect -1580 2299 -1556 2333
rect -1522 2299 -1498 2333
rect -1580 2261 -1498 2299
rect -1580 2227 -1556 2261
rect -1522 2227 -1498 2261
rect -1580 2189 -1498 2227
rect -1580 2155 -1556 2189
rect -1522 2155 -1498 2189
rect -1580 2117 -1498 2155
rect -1580 2083 -1556 2117
rect -1522 2083 -1498 2117
rect -1580 2045 -1498 2083
rect -1580 2011 -1556 2045
rect -1522 2011 -1498 2045
rect -1580 1973 -1498 2011
rect -1580 1939 -1556 1973
rect -1522 1939 -1498 1973
rect -1580 1901 -1498 1939
rect -1580 1867 -1556 1901
rect -1522 1867 -1498 1901
rect -1580 1829 -1498 1867
rect -1580 1795 -1556 1829
rect -1522 1795 -1498 1829
rect -1580 1757 -1498 1795
rect -1580 1723 -1556 1757
rect -1522 1723 -1498 1757
rect -1580 1685 -1498 1723
rect -1580 1651 -1556 1685
rect -1522 1651 -1498 1685
rect -1580 1613 -1498 1651
rect -1580 1579 -1556 1613
rect -1522 1579 -1498 1613
rect -1580 1541 -1498 1579
rect -1580 1507 -1556 1541
rect -1522 1507 -1498 1541
rect -1580 1469 -1498 1507
rect -1580 1435 -1556 1469
rect -1522 1435 -1498 1469
rect -1580 1397 -1498 1435
rect -1580 1363 -1556 1397
rect -1522 1363 -1498 1397
rect -1580 1325 -1498 1363
rect -1580 1291 -1556 1325
rect -1522 1291 -1498 1325
rect -1580 1253 -1498 1291
rect -1580 1219 -1556 1253
rect -1522 1219 -1498 1253
rect -1580 1181 -1498 1219
rect -1580 1147 -1556 1181
rect -1522 1147 -1498 1181
rect -1580 1109 -1498 1147
rect -1580 1075 -1556 1109
rect -1522 1075 -1498 1109
rect -1580 1037 -1498 1075
rect -1580 1003 -1556 1037
rect -1522 1003 -1498 1037
rect -1580 965 -1498 1003
rect -1580 931 -1556 965
rect -1522 931 -1498 965
rect -1580 893 -1498 931
rect -1580 859 -1556 893
rect -1522 859 -1498 893
rect -1580 821 -1498 859
rect -1580 787 -1556 821
rect -1522 787 -1498 821
rect -1580 749 -1498 787
rect -1580 715 -1556 749
rect -1522 715 -1498 749
rect -1580 677 -1498 715
rect -1580 643 -1556 677
rect -1522 643 -1498 677
rect -1580 605 -1498 643
rect -1580 571 -1556 605
rect -1522 571 -1498 605
rect -1580 533 -1498 571
rect -1580 499 -1556 533
rect -1522 499 -1498 533
rect -1580 461 -1498 499
rect -1580 427 -1556 461
rect -1522 427 -1498 461
rect -1580 389 -1498 427
rect -1580 355 -1556 389
rect -1522 355 -1498 389
rect -1580 317 -1498 355
rect -1580 283 -1556 317
rect -1522 283 -1498 317
rect -1580 245 -1498 283
rect -1580 211 -1556 245
rect -1522 211 -1498 245
rect -1580 173 -1498 211
rect -1580 139 -1556 173
rect -1522 139 -1498 173
rect -1580 101 -1498 139
rect -1580 67 -1556 101
rect -1522 67 -1498 101
rect -1580 29 -1498 67
rect -1580 -5 -1556 29
rect -1522 -5 -1498 29
rect -1580 -43 -1498 -5
rect -1580 -77 -1556 -43
rect -1522 -77 -1498 -43
rect -1580 -115 -1498 -77
rect -1580 -149 -1556 -115
rect -1522 -149 -1498 -115
rect -1580 -187 -1498 -149
rect -1580 -221 -1556 -187
rect -1522 -221 -1498 -187
rect -1580 -259 -1498 -221
rect -1580 -293 -1556 -259
rect -1522 -293 -1498 -259
rect -1580 -331 -1498 -293
rect -1580 -365 -1556 -331
rect -1522 -365 -1498 -331
rect -1580 -403 -1498 -365
rect -1580 -437 -1556 -403
rect -1522 -437 -1498 -403
rect -1580 -475 -1498 -437
rect -1580 -509 -1556 -475
rect -1522 -509 -1498 -475
rect -1580 -547 -1498 -509
rect -1580 -581 -1556 -547
rect -1522 -581 -1498 -547
rect -1580 -619 -1498 -581
rect -1580 -653 -1556 -619
rect -1522 -653 -1498 -619
rect -1580 -691 -1498 -653
rect -1580 -725 -1556 -691
rect -1522 -725 -1498 -691
rect -1580 -763 -1498 -725
rect -1580 -797 -1556 -763
rect -1522 -797 -1498 -763
rect -1580 -835 -1498 -797
rect -1580 -869 -1556 -835
rect -1522 -869 -1498 -835
rect -1580 -907 -1498 -869
rect -1580 -941 -1556 -907
rect -1522 -941 -1498 -907
rect -1580 -979 -1498 -941
rect -1580 -1013 -1556 -979
rect -1522 -1013 -1498 -979
rect -1580 -1051 -1498 -1013
rect -798 6998 948 7022
rect -798 6820 -554 6998
rect 704 6820 948 6998
rect -798 6757 948 6820
rect -798 6650 -716 6757
rect -798 6616 -774 6650
rect -740 6616 -716 6650
rect -798 6578 -716 6616
rect -798 6544 -774 6578
rect -740 6544 -716 6578
rect -798 6506 -716 6544
rect -798 6472 -774 6506
rect -740 6472 -716 6506
rect -798 6434 -716 6472
rect -798 6400 -774 6434
rect -740 6400 -716 6434
rect -798 6362 -716 6400
rect -798 6328 -774 6362
rect -740 6328 -716 6362
rect -798 6290 -716 6328
rect -798 6256 -774 6290
rect -740 6256 -716 6290
rect -798 6218 -716 6256
rect -798 6184 -774 6218
rect -740 6184 -716 6218
rect -798 6146 -716 6184
rect 866 6650 948 6757
rect 866 6616 890 6650
rect 924 6616 948 6650
rect 866 6578 948 6616
rect 866 6544 890 6578
rect 924 6544 948 6578
rect 866 6506 948 6544
rect 866 6472 890 6506
rect 924 6472 948 6506
rect 866 6434 948 6472
rect 866 6400 890 6434
rect 924 6400 948 6434
rect 866 6362 948 6400
rect 866 6328 890 6362
rect 924 6328 948 6362
rect 866 6290 948 6328
rect 866 6256 890 6290
rect 924 6256 948 6290
rect 866 6218 948 6256
rect 866 6184 890 6218
rect 924 6184 948 6218
rect -798 6112 -774 6146
rect -740 6112 -716 6146
rect -798 6074 -716 6112
rect -798 6040 -774 6074
rect -740 6040 -716 6074
rect -798 6002 -716 6040
rect -798 5968 -774 6002
rect -740 5968 -716 6002
rect -798 5930 -716 5968
rect -798 5896 -774 5930
rect -740 5896 -716 5930
rect -798 5858 -716 5896
rect -798 5824 -774 5858
rect -740 5824 -716 5858
rect -798 5786 -716 5824
rect -798 5752 -774 5786
rect -740 5752 -716 5786
rect -798 5714 -716 5752
rect -798 5680 -774 5714
rect -740 5680 -716 5714
rect -798 5642 -716 5680
rect -798 5608 -774 5642
rect -740 5608 -716 5642
rect -798 5570 -716 5608
rect -798 5536 -774 5570
rect -740 5536 -716 5570
rect -798 5498 -716 5536
rect -798 5464 -774 5498
rect -740 5464 -716 5498
rect -798 5426 -716 5464
rect -798 5392 -774 5426
rect -740 5392 -716 5426
rect -798 5354 -716 5392
rect -798 5320 -774 5354
rect -740 5320 -716 5354
rect -798 5282 -716 5320
rect -798 5248 -774 5282
rect -740 5248 -716 5282
rect -798 5210 -716 5248
rect -798 5176 -774 5210
rect -740 5176 -716 5210
rect -798 5138 -716 5176
rect -798 5104 -774 5138
rect -740 5104 -716 5138
rect -798 5066 -716 5104
rect -798 5032 -774 5066
rect -740 5032 -716 5066
rect -798 4994 -716 5032
rect -798 4960 -774 4994
rect -740 4960 -716 4994
rect -798 4922 -716 4960
rect -798 4888 -774 4922
rect -740 4888 -716 4922
rect -798 4850 -716 4888
rect -798 4816 -774 4850
rect -740 4816 -716 4850
rect -798 4778 -716 4816
rect -798 4744 -774 4778
rect -740 4744 -716 4778
rect -798 4706 -716 4744
rect -798 4672 -774 4706
rect -740 4672 -716 4706
rect -798 4634 -716 4672
rect -798 4600 -774 4634
rect -740 4600 -716 4634
rect -798 4562 -716 4600
rect -798 4528 -774 4562
rect -740 4528 -716 4562
rect -798 4490 -716 4528
rect -798 4456 -774 4490
rect -740 4456 -716 4490
rect -798 4418 -716 4456
rect -798 4384 -774 4418
rect -740 4384 -716 4418
rect -798 4346 -716 4384
rect -798 4312 -774 4346
rect -740 4312 -716 4346
rect -798 4274 -716 4312
rect -798 4240 -774 4274
rect -740 4240 -716 4274
rect -798 4202 -716 4240
rect -798 4168 -774 4202
rect -740 4168 -716 4202
rect -798 4130 -716 4168
rect -798 4096 -774 4130
rect -740 4096 -716 4130
rect -798 4058 -716 4096
rect -798 4024 -774 4058
rect -740 4024 -716 4058
rect -798 3986 -716 4024
rect -798 3952 -774 3986
rect -740 3952 -716 3986
rect -798 3914 -716 3952
rect -798 3880 -774 3914
rect -740 3880 -716 3914
rect -798 3842 -716 3880
rect -798 3808 -774 3842
rect -740 3808 -716 3842
rect -798 3770 -716 3808
rect -798 3736 -774 3770
rect -740 3736 -716 3770
rect -798 3698 -716 3736
rect -798 3664 -774 3698
rect -740 3664 -716 3698
rect -798 3626 -716 3664
rect -798 3592 -774 3626
rect -740 3592 -716 3626
rect -798 3554 -716 3592
rect -798 3520 -774 3554
rect -740 3520 -716 3554
rect -798 3482 -716 3520
rect -798 3448 -774 3482
rect -740 3448 -716 3482
rect -798 3410 -716 3448
rect -798 3376 -774 3410
rect -740 3376 -716 3410
rect -798 3338 -716 3376
rect -798 3304 -774 3338
rect -740 3304 -716 3338
rect -798 3266 -716 3304
rect -798 3232 -774 3266
rect -740 3232 -716 3266
rect -798 3194 -716 3232
rect -798 3160 -774 3194
rect -740 3160 -716 3194
rect -798 3122 -716 3160
rect -798 3088 -774 3122
rect -740 3088 -716 3122
rect -798 3050 -716 3088
rect -798 3016 -774 3050
rect -740 3016 -716 3050
rect -798 2978 -716 3016
rect -798 2944 -774 2978
rect -740 2944 -716 2978
rect -798 2906 -716 2944
rect -798 2872 -774 2906
rect -740 2872 -716 2906
rect -798 2834 -716 2872
rect -798 2800 -774 2834
rect -740 2800 -716 2834
rect -798 2762 -716 2800
rect -798 2728 -774 2762
rect -740 2728 -716 2762
rect -798 2690 -716 2728
rect -798 2656 -774 2690
rect -740 2656 -716 2690
rect -798 2618 -716 2656
rect -798 2584 -774 2618
rect -740 2584 -716 2618
rect -798 2546 -716 2584
rect -798 2512 -774 2546
rect -740 2512 -716 2546
rect -798 2474 -716 2512
rect -798 2440 -774 2474
rect -740 2440 -716 2474
rect -798 2402 -716 2440
rect -798 2368 -774 2402
rect -740 2368 -716 2402
rect -798 2330 -716 2368
rect -798 2296 -774 2330
rect -740 2296 -716 2330
rect -798 2258 -716 2296
rect -798 2224 -774 2258
rect -740 2224 -716 2258
rect -798 2186 -716 2224
rect -798 2152 -774 2186
rect -740 2152 -716 2186
rect -798 2114 -716 2152
rect -798 2080 -774 2114
rect -740 2080 -716 2114
rect -798 2042 -716 2080
rect -798 2008 -774 2042
rect -740 2008 -716 2042
rect -798 1970 -716 2008
rect -798 1936 -774 1970
rect -740 1936 -716 1970
rect -798 1898 -716 1936
rect -798 1864 -774 1898
rect -740 1864 -716 1898
rect -798 1826 -716 1864
rect -798 1792 -774 1826
rect -740 1792 -716 1826
rect -798 1754 -716 1792
rect -798 1720 -774 1754
rect -740 1720 -716 1754
rect -798 1682 -716 1720
rect -798 1648 -774 1682
rect -740 1648 -716 1682
rect -798 1610 -716 1648
rect -798 1576 -774 1610
rect -740 1576 -716 1610
rect -798 1538 -716 1576
rect -798 1504 -774 1538
rect -740 1504 -716 1538
rect -798 1466 -716 1504
rect -798 1432 -774 1466
rect -740 1432 -716 1466
rect -798 1394 -716 1432
rect -798 1360 -774 1394
rect -740 1360 -716 1394
rect -798 1322 -716 1360
rect -798 1288 -774 1322
rect -740 1288 -716 1322
rect -798 1250 -716 1288
rect -798 1216 -774 1250
rect -740 1216 -716 1250
rect -798 1178 -716 1216
rect -798 1144 -774 1178
rect -740 1144 -716 1178
rect -798 1106 -716 1144
rect -798 1072 -774 1106
rect -740 1072 -716 1106
rect -798 1034 -716 1072
rect -798 1000 -774 1034
rect -740 1000 -716 1034
rect -798 962 -716 1000
rect -798 928 -774 962
rect -740 928 -716 962
rect -798 890 -716 928
rect -798 856 -774 890
rect -740 856 -716 890
rect -798 818 -716 856
rect -798 784 -774 818
rect -740 784 -716 818
rect -798 746 -716 784
rect -798 712 -774 746
rect -740 712 -716 746
rect -798 674 -716 712
rect -798 640 -774 674
rect -740 640 -716 674
rect -798 602 -716 640
rect -798 568 -774 602
rect -740 568 -716 602
rect -798 530 -716 568
rect -798 496 -774 530
rect -740 496 -716 530
rect -798 458 -716 496
rect -798 424 -774 458
rect -740 424 -716 458
rect -798 386 -716 424
rect -798 352 -774 386
rect -740 352 -716 386
rect -798 314 -716 352
rect -798 280 -774 314
rect -740 280 -716 314
rect -798 242 -716 280
rect -798 208 -774 242
rect -740 208 -716 242
rect -798 170 -716 208
rect -798 136 -774 170
rect -740 136 -716 170
rect -798 98 -716 136
rect -798 64 -774 98
rect -740 64 -716 98
rect -798 26 -716 64
rect -798 -8 -774 26
rect -740 -8 -716 26
rect -798 -46 -716 -8
rect -798 -80 -774 -46
rect -740 -80 -716 -46
rect -798 -118 -716 -80
rect -798 -152 -774 -118
rect -740 -152 -716 -118
rect -798 -190 -716 -152
rect -659 6146 -457 6165
rect -659 6127 -647 6146
rect -469 6127 -457 6146
rect -659 -133 -648 6127
rect -468 -133 -457 6127
rect -659 -152 -647 -133
rect -469 -152 -457 -133
rect -659 -164 -457 -152
rect -134 6146 284 6165
rect -134 -152 -122 6146
rect 272 -152 284 6146
rect -134 -164 284 -152
rect 607 6146 809 6165
rect 607 6127 619 6146
rect 797 6127 809 6146
rect 607 -133 618 6127
rect 798 -133 809 6127
rect 607 -152 619 -133
rect 797 -152 809 -133
rect 607 -164 809 -152
rect 866 6146 948 6184
rect 866 6112 890 6146
rect 924 6112 948 6146
rect 866 6074 948 6112
rect 866 6040 890 6074
rect 924 6040 948 6074
rect 866 6002 948 6040
rect 866 5968 890 6002
rect 924 5968 948 6002
rect 866 5930 948 5968
rect 866 5896 890 5930
rect 924 5896 948 5930
rect 866 5858 948 5896
rect 866 5824 890 5858
rect 924 5824 948 5858
rect 866 5786 948 5824
rect 866 5752 890 5786
rect 924 5752 948 5786
rect 866 5714 948 5752
rect 866 5680 890 5714
rect 924 5680 948 5714
rect 866 5642 948 5680
rect 866 5608 890 5642
rect 924 5608 948 5642
rect 866 5570 948 5608
rect 866 5536 890 5570
rect 924 5536 948 5570
rect 866 5498 948 5536
rect 866 5464 890 5498
rect 924 5464 948 5498
rect 866 5426 948 5464
rect 866 5392 890 5426
rect 924 5392 948 5426
rect 866 5354 948 5392
rect 866 5320 890 5354
rect 924 5320 948 5354
rect 866 5282 948 5320
rect 866 5248 890 5282
rect 924 5248 948 5282
rect 866 5210 948 5248
rect 866 5176 890 5210
rect 924 5176 948 5210
rect 866 5138 948 5176
rect 866 5104 890 5138
rect 924 5104 948 5138
rect 866 5066 948 5104
rect 866 5032 890 5066
rect 924 5032 948 5066
rect 866 4994 948 5032
rect 866 4960 890 4994
rect 924 4960 948 4994
rect 866 4922 948 4960
rect 866 4888 890 4922
rect 924 4888 948 4922
rect 866 4850 948 4888
rect 866 4816 890 4850
rect 924 4816 948 4850
rect 866 4778 948 4816
rect 866 4744 890 4778
rect 924 4744 948 4778
rect 866 4706 948 4744
rect 866 4672 890 4706
rect 924 4672 948 4706
rect 866 4634 948 4672
rect 866 4600 890 4634
rect 924 4600 948 4634
rect 866 4562 948 4600
rect 866 4528 890 4562
rect 924 4528 948 4562
rect 866 4490 948 4528
rect 866 4456 890 4490
rect 924 4456 948 4490
rect 866 4418 948 4456
rect 866 4384 890 4418
rect 924 4384 948 4418
rect 866 4346 948 4384
rect 866 4312 890 4346
rect 924 4312 948 4346
rect 866 4274 948 4312
rect 866 4240 890 4274
rect 924 4240 948 4274
rect 866 4202 948 4240
rect 866 4168 890 4202
rect 924 4168 948 4202
rect 866 4130 948 4168
rect 866 4096 890 4130
rect 924 4096 948 4130
rect 866 4058 948 4096
rect 866 4024 890 4058
rect 924 4024 948 4058
rect 866 3986 948 4024
rect 866 3952 890 3986
rect 924 3952 948 3986
rect 866 3914 948 3952
rect 866 3880 890 3914
rect 924 3880 948 3914
rect 866 3842 948 3880
rect 866 3808 890 3842
rect 924 3808 948 3842
rect 866 3770 948 3808
rect 866 3736 890 3770
rect 924 3736 948 3770
rect 866 3698 948 3736
rect 866 3664 890 3698
rect 924 3664 948 3698
rect 866 3626 948 3664
rect 866 3592 890 3626
rect 924 3592 948 3626
rect 866 3554 948 3592
rect 866 3520 890 3554
rect 924 3520 948 3554
rect 866 3482 948 3520
rect 866 3448 890 3482
rect 924 3448 948 3482
rect 866 3410 948 3448
rect 866 3376 890 3410
rect 924 3376 948 3410
rect 866 3338 948 3376
rect 866 3304 890 3338
rect 924 3304 948 3338
rect 866 3266 948 3304
rect 866 3232 890 3266
rect 924 3232 948 3266
rect 866 3194 948 3232
rect 866 3160 890 3194
rect 924 3160 948 3194
rect 866 3122 948 3160
rect 866 3088 890 3122
rect 924 3088 948 3122
rect 866 3050 948 3088
rect 866 3016 890 3050
rect 924 3016 948 3050
rect 866 2978 948 3016
rect 866 2944 890 2978
rect 924 2944 948 2978
rect 866 2906 948 2944
rect 866 2872 890 2906
rect 924 2872 948 2906
rect 866 2834 948 2872
rect 866 2800 890 2834
rect 924 2800 948 2834
rect 866 2762 948 2800
rect 866 2728 890 2762
rect 924 2728 948 2762
rect 866 2690 948 2728
rect 866 2656 890 2690
rect 924 2656 948 2690
rect 866 2618 948 2656
rect 866 2584 890 2618
rect 924 2584 948 2618
rect 866 2546 948 2584
rect 866 2512 890 2546
rect 924 2512 948 2546
rect 866 2474 948 2512
rect 866 2440 890 2474
rect 924 2440 948 2474
rect 866 2402 948 2440
rect 866 2368 890 2402
rect 924 2368 948 2402
rect 866 2330 948 2368
rect 866 2296 890 2330
rect 924 2296 948 2330
rect 866 2258 948 2296
rect 866 2224 890 2258
rect 924 2224 948 2258
rect 866 2186 948 2224
rect 866 2152 890 2186
rect 924 2152 948 2186
rect 866 2114 948 2152
rect 866 2080 890 2114
rect 924 2080 948 2114
rect 866 2042 948 2080
rect 866 2008 890 2042
rect 924 2008 948 2042
rect 866 1970 948 2008
rect 866 1936 890 1970
rect 924 1936 948 1970
rect 866 1898 948 1936
rect 866 1864 890 1898
rect 924 1864 948 1898
rect 866 1826 948 1864
rect 866 1792 890 1826
rect 924 1792 948 1826
rect 866 1754 948 1792
rect 866 1720 890 1754
rect 924 1720 948 1754
rect 866 1682 948 1720
rect 866 1648 890 1682
rect 924 1648 948 1682
rect 866 1610 948 1648
rect 866 1576 890 1610
rect 924 1576 948 1610
rect 866 1538 948 1576
rect 866 1504 890 1538
rect 924 1504 948 1538
rect 866 1466 948 1504
rect 866 1432 890 1466
rect 924 1432 948 1466
rect 866 1394 948 1432
rect 866 1360 890 1394
rect 924 1360 948 1394
rect 866 1322 948 1360
rect 866 1288 890 1322
rect 924 1288 948 1322
rect 866 1250 948 1288
rect 866 1216 890 1250
rect 924 1216 948 1250
rect 866 1178 948 1216
rect 866 1144 890 1178
rect 924 1144 948 1178
rect 866 1106 948 1144
rect 866 1072 890 1106
rect 924 1072 948 1106
rect 866 1034 948 1072
rect 866 1000 890 1034
rect 924 1000 948 1034
rect 866 962 948 1000
rect 866 928 890 962
rect 924 928 948 962
rect 866 890 948 928
rect 866 856 890 890
rect 924 856 948 890
rect 866 818 948 856
rect 866 784 890 818
rect 924 784 948 818
rect 866 746 948 784
rect 866 712 890 746
rect 924 712 948 746
rect 866 674 948 712
rect 866 640 890 674
rect 924 640 948 674
rect 866 602 948 640
rect 866 568 890 602
rect 924 568 948 602
rect 866 530 948 568
rect 866 496 890 530
rect 924 496 948 530
rect 866 458 948 496
rect 866 424 890 458
rect 924 424 948 458
rect 866 386 948 424
rect 866 352 890 386
rect 924 352 948 386
rect 866 314 948 352
rect 866 280 890 314
rect 924 280 948 314
rect 866 242 948 280
rect 866 208 890 242
rect 924 208 948 242
rect 866 170 948 208
rect 866 136 890 170
rect 924 136 948 170
rect 866 98 948 136
rect 866 64 890 98
rect 924 64 948 98
rect 866 26 948 64
rect 866 -8 890 26
rect 924 -8 948 26
rect 866 -46 948 -8
rect 866 -80 890 -46
rect 924 -80 948 -46
rect 866 -118 948 -80
rect 866 -152 890 -118
rect 924 -152 948 -118
rect -798 -224 -774 -190
rect -740 -224 -716 -190
rect -798 -262 -716 -224
rect -798 -296 -774 -262
rect -740 -296 -716 -262
rect -798 -334 -716 -296
rect -798 -368 -774 -334
rect -740 -368 -716 -334
rect -798 -406 -716 -368
rect -798 -440 -774 -406
rect -740 -440 -716 -406
rect -798 -478 -716 -440
rect 866 -190 948 -152
rect 866 -224 890 -190
rect 924 -224 948 -190
rect 866 -262 948 -224
rect 866 -296 890 -262
rect 924 -296 948 -262
rect 866 -334 948 -296
rect 866 -368 890 -334
rect 924 -368 948 -334
rect 866 -406 948 -368
rect 866 -440 890 -406
rect 924 -440 948 -406
rect -798 -512 -774 -478
rect -740 -512 -716 -478
rect -798 -550 -716 -512
rect -798 -584 -774 -550
rect -740 -584 -716 -550
rect -798 -622 -716 -584
rect -798 -656 -774 -622
rect -740 -656 -716 -622
rect -798 -757 -716 -656
rect -146 -450 290 -443
rect -146 -502 -139 -450
rect -87 -502 -65 -450
rect -13 -502 9 -450
rect 61 -502 83 -450
rect 135 -502 157 -450
rect 209 -502 231 -450
rect 283 -502 290 -450
rect -146 -524 290 -502
rect -146 -576 -139 -524
rect -87 -576 -65 -524
rect -13 -576 9 -524
rect 61 -576 83 -524
rect 135 -576 157 -524
rect 209 -576 231 -524
rect 283 -576 290 -524
rect -146 -598 290 -576
rect -146 -650 -139 -598
rect -87 -650 -65 -598
rect -13 -650 9 -598
rect 61 -650 83 -598
rect 135 -650 157 -598
rect 209 -650 231 -598
rect 283 -650 290 -598
rect -146 -657 290 -650
rect 866 -478 948 -440
rect 866 -512 890 -478
rect 924 -512 948 -478
rect 866 -550 948 -512
rect 866 -584 890 -550
rect 924 -584 948 -550
rect 866 -622 948 -584
rect 866 -656 890 -622
rect 924 -656 948 -622
rect 866 -757 948 -656
rect -798 -820 948 -757
rect -798 -998 -554 -820
rect 704 -998 948 -820
rect -798 -1022 948 -998
rect 1648 7013 1730 7051
rect 1648 6979 1672 7013
rect 1706 6979 1730 7013
rect 1648 6941 1730 6979
rect 1648 6907 1672 6941
rect 1706 6907 1730 6941
rect 1648 6869 1730 6907
rect 1648 6835 1672 6869
rect 1706 6835 1730 6869
rect 1648 6797 1730 6835
rect 1648 6763 1672 6797
rect 1706 6763 1730 6797
rect 1648 6725 1730 6763
rect 1648 6691 1672 6725
rect 1706 6691 1730 6725
rect 1648 6653 1730 6691
rect 1648 6619 1672 6653
rect 1706 6619 1730 6653
rect 1648 6581 1730 6619
rect 1648 6547 1672 6581
rect 1706 6547 1730 6581
rect 1648 6509 1730 6547
rect 1648 6475 1672 6509
rect 1706 6475 1730 6509
rect 1648 6437 1730 6475
rect 1648 6403 1672 6437
rect 1706 6403 1730 6437
rect 1648 6365 1730 6403
rect 1648 6331 1672 6365
rect 1706 6331 1730 6365
rect 1648 6293 1730 6331
rect 1648 6259 1672 6293
rect 1706 6259 1730 6293
rect 1648 6221 1730 6259
rect 1648 6187 1672 6221
rect 1706 6187 1730 6221
rect 1648 6149 1730 6187
rect 1648 6115 1672 6149
rect 1706 6115 1730 6149
rect 1648 6077 1730 6115
rect 1648 6043 1672 6077
rect 1706 6043 1730 6077
rect 1648 6005 1730 6043
rect 1648 5971 1672 6005
rect 1706 5971 1730 6005
rect 1648 5933 1730 5971
rect 1648 5899 1672 5933
rect 1706 5899 1730 5933
rect 1648 5861 1730 5899
rect 1648 5827 1672 5861
rect 1706 5827 1730 5861
rect 1648 5789 1730 5827
rect 1648 5755 1672 5789
rect 1706 5755 1730 5789
rect 1648 5717 1730 5755
rect 1648 5683 1672 5717
rect 1706 5683 1730 5717
rect 1648 5645 1730 5683
rect 1648 5611 1672 5645
rect 1706 5611 1730 5645
rect 1648 5573 1730 5611
rect 1648 5539 1672 5573
rect 1706 5539 1730 5573
rect 1648 5501 1730 5539
rect 1648 5467 1672 5501
rect 1706 5467 1730 5501
rect 1648 5429 1730 5467
rect 1648 5395 1672 5429
rect 1706 5395 1730 5429
rect 1648 5357 1730 5395
rect 1648 5323 1672 5357
rect 1706 5323 1730 5357
rect 1648 5285 1730 5323
rect 1648 5251 1672 5285
rect 1706 5251 1730 5285
rect 1648 5213 1730 5251
rect 1648 5179 1672 5213
rect 1706 5179 1730 5213
rect 1648 5141 1730 5179
rect 1648 5107 1672 5141
rect 1706 5107 1730 5141
rect 1648 5069 1730 5107
rect 1648 5035 1672 5069
rect 1706 5035 1730 5069
rect 1648 4997 1730 5035
rect 1648 4963 1672 4997
rect 1706 4963 1730 4997
rect 1648 4925 1730 4963
rect 1648 4891 1672 4925
rect 1706 4891 1730 4925
rect 1648 4853 1730 4891
rect 1648 4819 1672 4853
rect 1706 4819 1730 4853
rect 1648 4781 1730 4819
rect 1648 4747 1672 4781
rect 1706 4747 1730 4781
rect 1648 4709 1730 4747
rect 1648 4675 1672 4709
rect 1706 4675 1730 4709
rect 1648 4637 1730 4675
rect 1648 4603 1672 4637
rect 1706 4603 1730 4637
rect 1648 4565 1730 4603
rect 1648 4531 1672 4565
rect 1706 4531 1730 4565
rect 1648 4493 1730 4531
rect 1648 4459 1672 4493
rect 1706 4459 1730 4493
rect 1648 4421 1730 4459
rect 1648 4387 1672 4421
rect 1706 4387 1730 4421
rect 1648 4349 1730 4387
rect 1648 4315 1672 4349
rect 1706 4315 1730 4349
rect 1648 4277 1730 4315
rect 1648 4243 1672 4277
rect 1706 4243 1730 4277
rect 1648 4205 1730 4243
rect 1648 4171 1672 4205
rect 1706 4171 1730 4205
rect 1648 4133 1730 4171
rect 1648 4099 1672 4133
rect 1706 4099 1730 4133
rect 1648 4061 1730 4099
rect 1648 4027 1672 4061
rect 1706 4027 1730 4061
rect 1648 3989 1730 4027
rect 1648 3955 1672 3989
rect 1706 3955 1730 3989
rect 1648 3917 1730 3955
rect 1648 3883 1672 3917
rect 1706 3883 1730 3917
rect 1648 3845 1730 3883
rect 1648 3811 1672 3845
rect 1706 3811 1730 3845
rect 1648 3773 1730 3811
rect 1648 3739 1672 3773
rect 1706 3739 1730 3773
rect 1648 3701 1730 3739
rect 1648 3667 1672 3701
rect 1706 3667 1730 3701
rect 1648 3629 1730 3667
rect 1648 3595 1672 3629
rect 1706 3595 1730 3629
rect 1648 3557 1730 3595
rect 1648 3523 1672 3557
rect 1706 3523 1730 3557
rect 1648 3485 1730 3523
rect 1648 3451 1672 3485
rect 1706 3451 1730 3485
rect 1648 3413 1730 3451
rect 1648 3379 1672 3413
rect 1706 3379 1730 3413
rect 1648 3341 1730 3379
rect 1648 3307 1672 3341
rect 1706 3307 1730 3341
rect 1648 3269 1730 3307
rect 1648 3235 1672 3269
rect 1706 3235 1730 3269
rect 1648 3197 1730 3235
rect 1648 3163 1672 3197
rect 1706 3163 1730 3197
rect 1648 3125 1730 3163
rect 1648 3091 1672 3125
rect 1706 3091 1730 3125
rect 1648 3053 1730 3091
rect 1648 3019 1672 3053
rect 1706 3019 1730 3053
rect 1648 2981 1730 3019
rect 1648 2947 1672 2981
rect 1706 2947 1730 2981
rect 1648 2909 1730 2947
rect 1648 2875 1672 2909
rect 1706 2875 1730 2909
rect 1648 2837 1730 2875
rect 1648 2803 1672 2837
rect 1706 2803 1730 2837
rect 1648 2765 1730 2803
rect 1648 2731 1672 2765
rect 1706 2731 1730 2765
rect 1648 2693 1730 2731
rect 1648 2659 1672 2693
rect 1706 2659 1730 2693
rect 1648 2621 1730 2659
rect 1648 2587 1672 2621
rect 1706 2587 1730 2621
rect 1648 2549 1730 2587
rect 1648 2515 1672 2549
rect 1706 2515 1730 2549
rect 1648 2477 1730 2515
rect 1648 2443 1672 2477
rect 1706 2443 1730 2477
rect 1648 2405 1730 2443
rect 1648 2371 1672 2405
rect 1706 2371 1730 2405
rect 1648 2333 1730 2371
rect 1648 2299 1672 2333
rect 1706 2299 1730 2333
rect 1648 2261 1730 2299
rect 1648 2227 1672 2261
rect 1706 2227 1730 2261
rect 1648 2189 1730 2227
rect 1648 2155 1672 2189
rect 1706 2155 1730 2189
rect 1648 2117 1730 2155
rect 1648 2083 1672 2117
rect 1706 2083 1730 2117
rect 1648 2045 1730 2083
rect 1648 2011 1672 2045
rect 1706 2011 1730 2045
rect 1648 1973 1730 2011
rect 1648 1939 1672 1973
rect 1706 1939 1730 1973
rect 1648 1901 1730 1939
rect 1648 1867 1672 1901
rect 1706 1867 1730 1901
rect 1648 1829 1730 1867
rect 1648 1795 1672 1829
rect 1706 1795 1730 1829
rect 1648 1757 1730 1795
rect 1648 1723 1672 1757
rect 1706 1723 1730 1757
rect 1648 1685 1730 1723
rect 1648 1651 1672 1685
rect 1706 1651 1730 1685
rect 1648 1613 1730 1651
rect 1648 1579 1672 1613
rect 1706 1579 1730 1613
rect 1648 1541 1730 1579
rect 1648 1507 1672 1541
rect 1706 1507 1730 1541
rect 1648 1469 1730 1507
rect 1648 1435 1672 1469
rect 1706 1435 1730 1469
rect 1648 1397 1730 1435
rect 1648 1363 1672 1397
rect 1706 1363 1730 1397
rect 1648 1325 1730 1363
rect 1648 1291 1672 1325
rect 1706 1291 1730 1325
rect 1648 1253 1730 1291
rect 1648 1219 1672 1253
rect 1706 1219 1730 1253
rect 1648 1181 1730 1219
rect 1648 1147 1672 1181
rect 1706 1147 1730 1181
rect 1648 1109 1730 1147
rect 1648 1075 1672 1109
rect 1706 1075 1730 1109
rect 1648 1037 1730 1075
rect 1648 1003 1672 1037
rect 1706 1003 1730 1037
rect 1648 965 1730 1003
rect 1648 931 1672 965
rect 1706 931 1730 965
rect 1648 893 1730 931
rect 1648 859 1672 893
rect 1706 859 1730 893
rect 1648 821 1730 859
rect 1648 787 1672 821
rect 1706 787 1730 821
rect 1648 749 1730 787
rect 1648 715 1672 749
rect 1706 715 1730 749
rect 1648 677 1730 715
rect 1648 643 1672 677
rect 1706 643 1730 677
rect 1648 605 1730 643
rect 1648 571 1672 605
rect 1706 571 1730 605
rect 1648 533 1730 571
rect 1648 499 1672 533
rect 1706 499 1730 533
rect 1648 461 1730 499
rect 1648 427 1672 461
rect 1706 427 1730 461
rect 1648 389 1730 427
rect 1648 355 1672 389
rect 1706 355 1730 389
rect 1648 317 1730 355
rect 1648 283 1672 317
rect 1706 283 1730 317
rect 1648 245 1730 283
rect 1648 211 1672 245
rect 1706 211 1730 245
rect 1648 173 1730 211
rect 1648 139 1672 173
rect 1706 139 1730 173
rect 1648 101 1730 139
rect 1648 67 1672 101
rect 1706 67 1730 101
rect 1648 29 1730 67
rect 1648 -5 1672 29
rect 1706 -5 1730 29
rect 1648 -43 1730 -5
rect 1648 -77 1672 -43
rect 1706 -77 1730 -43
rect 1648 -115 1730 -77
rect 1648 -149 1672 -115
rect 1706 -149 1730 -115
rect 1648 -187 1730 -149
rect 1648 -221 1672 -187
rect 1706 -221 1730 -187
rect 1648 -259 1730 -221
rect 1648 -293 1672 -259
rect 1706 -293 1730 -259
rect 1648 -331 1730 -293
rect 1648 -365 1672 -331
rect 1706 -365 1730 -331
rect 1648 -403 1730 -365
rect 1648 -437 1672 -403
rect 1706 -437 1730 -403
rect 1648 -475 1730 -437
rect 1648 -509 1672 -475
rect 1706 -509 1730 -475
rect 1648 -547 1730 -509
rect 1648 -581 1672 -547
rect 1706 -581 1730 -547
rect 1648 -619 1730 -581
rect 1648 -653 1672 -619
rect 1706 -653 1730 -619
rect 1648 -691 1730 -653
rect 1648 -725 1672 -691
rect 1706 -725 1730 -691
rect 1648 -763 1730 -725
rect 1648 -797 1672 -763
rect 1706 -797 1730 -763
rect 1648 -835 1730 -797
rect 1648 -869 1672 -835
rect 1706 -869 1730 -835
rect 1648 -907 1730 -869
rect 1648 -941 1672 -907
rect 1706 -941 1730 -907
rect 1648 -979 1730 -941
rect 1648 -1013 1672 -979
rect 1706 -1013 1730 -979
rect -1580 -1085 -1556 -1051
rect -1522 -1085 -1498 -1051
rect -1580 -1123 -1498 -1085
rect -1580 -1157 -1556 -1123
rect -1522 -1157 -1498 -1123
rect -1580 -1195 -1498 -1157
rect -1580 -1229 -1556 -1195
rect -1522 -1229 -1498 -1195
rect -1580 -1267 -1498 -1229
rect -1580 -1301 -1556 -1267
rect -1522 -1301 -1498 -1267
rect -1580 -1339 -1498 -1301
rect -1580 -1373 -1556 -1339
rect -1522 -1373 -1498 -1339
rect -1580 -1411 -1498 -1373
rect -1580 -1445 -1556 -1411
rect -1522 -1445 -1498 -1411
rect -1580 -1483 -1498 -1445
rect -1580 -1517 -1556 -1483
rect -1522 -1517 -1498 -1483
rect -1580 -1555 -1498 -1517
rect -1580 -1589 -1556 -1555
rect -1522 -1589 -1498 -1555
rect -1580 -1627 -1498 -1589
rect -1580 -1661 -1556 -1627
rect -1522 -1661 -1498 -1627
rect -1580 -1722 -1498 -1661
rect 1648 -1051 1730 -1013
rect 1648 -1085 1672 -1051
rect 1706 -1085 1730 -1051
rect 1648 -1123 1730 -1085
rect 1648 -1157 1672 -1123
rect 1706 -1157 1730 -1123
rect 1648 -1195 1730 -1157
rect 1648 -1229 1672 -1195
rect 1706 -1229 1730 -1195
rect 1648 -1267 1730 -1229
rect 1648 -1301 1672 -1267
rect 1706 -1301 1730 -1267
rect 1648 -1339 1730 -1301
rect 1648 -1373 1672 -1339
rect 1706 -1373 1730 -1339
rect 1648 -1411 1730 -1373
rect 1648 -1445 1672 -1411
rect 1706 -1445 1730 -1411
rect 1648 -1483 1730 -1445
rect 1648 -1517 1672 -1483
rect 1706 -1517 1730 -1483
rect 1648 -1555 1730 -1517
rect 1648 -1589 1672 -1555
rect 1706 -1589 1730 -1555
rect 1648 -1627 1730 -1589
rect 1648 -1661 1672 -1627
rect 1706 -1661 1730 -1627
rect 1648 -1722 1730 -1661
rect -1580 -1746 1730 -1722
rect -1580 -1780 -1454 -1746
rect -1420 -1780 -1382 -1746
rect -1348 -1780 -1310 -1746
rect -1276 -1780 -1238 -1746
rect -1204 -1780 -1166 -1746
rect -1132 -1780 -1094 -1746
rect -1060 -1780 -1022 -1746
rect -988 -1780 -950 -1746
rect -916 -1780 -878 -1746
rect -844 -1780 -806 -1746
rect -772 -1780 -734 -1746
rect -700 -1780 -662 -1746
rect -628 -1780 -590 -1746
rect -556 -1780 -518 -1746
rect -484 -1780 -446 -1746
rect -412 -1780 -374 -1746
rect -340 -1780 -302 -1746
rect -268 -1780 -230 -1746
rect -196 -1780 -158 -1746
rect -124 -1780 -86 -1746
rect -52 -1780 -14 -1746
rect 20 -1780 58 -1746
rect 92 -1780 130 -1746
rect 164 -1780 202 -1746
rect 236 -1780 274 -1746
rect 308 -1780 346 -1746
rect 380 -1780 418 -1746
rect 452 -1780 490 -1746
rect 524 -1780 562 -1746
rect 596 -1780 634 -1746
rect 668 -1780 706 -1746
rect 740 -1780 778 -1746
rect 812 -1780 850 -1746
rect 884 -1780 922 -1746
rect 956 -1780 994 -1746
rect 1028 -1780 1066 -1746
rect 1100 -1780 1138 -1746
rect 1172 -1780 1210 -1746
rect 1244 -1780 1282 -1746
rect 1316 -1780 1354 -1746
rect 1388 -1780 1426 -1746
rect 1460 -1780 1498 -1746
rect 1532 -1780 1570 -1746
rect 1604 -1780 1730 -1746
rect -1580 -1804 1730 -1780
<< via1 >>
rect -648 -133 -647 6127
rect -647 -133 -469 6127
rect -469 -133 -468 6127
rect -111 -133 261 6127
rect 618 -133 619 6127
rect 619 -133 797 6127
rect 797 -133 798 6127
rect -139 -459 -87 -450
rect -139 -493 -130 -459
rect -130 -493 -96 -459
rect -96 -493 -87 -459
rect -139 -502 -87 -493
rect -65 -459 -13 -450
rect -65 -493 -56 -459
rect -56 -493 -22 -459
rect -22 -493 -13 -459
rect -65 -502 -13 -493
rect 9 -459 61 -450
rect 9 -493 18 -459
rect 18 -493 52 -459
rect 52 -493 61 -459
rect 9 -502 61 -493
rect 83 -459 135 -450
rect 83 -493 92 -459
rect 92 -493 126 -459
rect 126 -493 135 -459
rect 83 -502 135 -493
rect 157 -459 209 -450
rect 157 -493 166 -459
rect 166 -493 200 -459
rect 200 -493 209 -459
rect 157 -502 209 -493
rect 231 -459 283 -450
rect 231 -493 240 -459
rect 240 -493 274 -459
rect 274 -493 283 -459
rect 231 -502 283 -493
rect -139 -533 -87 -524
rect -139 -567 -130 -533
rect -130 -567 -96 -533
rect -96 -567 -87 -533
rect -139 -576 -87 -567
rect -65 -533 -13 -524
rect -65 -567 -56 -533
rect -56 -567 -22 -533
rect -22 -567 -13 -533
rect -65 -576 -13 -567
rect 9 -533 61 -524
rect 9 -567 18 -533
rect 18 -567 52 -533
rect 52 -567 61 -533
rect 9 -576 61 -567
rect 83 -533 135 -524
rect 83 -567 92 -533
rect 92 -567 126 -533
rect 126 -567 135 -533
rect 83 -576 135 -567
rect 157 -533 209 -524
rect 157 -567 166 -533
rect 166 -567 200 -533
rect 200 -567 209 -533
rect 157 -576 209 -567
rect 231 -533 283 -524
rect 231 -567 240 -533
rect 240 -567 274 -533
rect 274 -567 283 -533
rect 231 -576 283 -567
rect -139 -607 -87 -598
rect -139 -641 -130 -607
rect -130 -641 -96 -607
rect -96 -641 -87 -607
rect -139 -650 -87 -641
rect -65 -607 -13 -598
rect -65 -641 -56 -607
rect -56 -641 -22 -607
rect -22 -641 -13 -607
rect -65 -650 -13 -641
rect 9 -607 61 -598
rect 9 -641 18 -607
rect 18 -641 52 -607
rect 52 -641 61 -607
rect 9 -650 61 -641
rect 83 -607 135 -598
rect 83 -641 92 -607
rect 92 -641 126 -607
rect 126 -641 135 -607
rect 83 -650 135 -641
rect 157 -607 209 -598
rect 157 -641 166 -607
rect 166 -641 200 -607
rect 200 -641 209 -607
rect 157 -650 209 -641
rect 231 -607 283 -598
rect 231 -641 240 -607
rect 240 -641 274 -607
rect 274 -641 283 -607
rect 231 -650 283 -641
<< metal2 >>
rect -659 6127 -457 6165
rect -659 -133 -648 6127
rect -468 -133 -457 6127
rect -659 -1122 -457 -133
rect -134 6127 284 7122
rect -134 -133 -111 6127
rect 261 -133 284 6127
rect -134 -164 284 -133
rect 607 6127 809 6165
rect 607 -133 618 6127
rect 798 -133 809 6127
rect -146 -450 290 -443
rect -146 -502 -139 -450
rect -87 -479 -65 -450
rect -13 -479 9 -450
rect 61 -479 83 -450
rect 135 -479 157 -450
rect 209 -479 231 -450
rect 283 -502 290 -450
rect -146 -524 -116 -502
rect 260 -524 290 -502
rect -146 -576 -139 -524
rect 283 -576 290 -524
rect -146 -598 -116 -576
rect 260 -598 290 -576
rect -146 -650 -139 -598
rect -87 -650 -65 -615
rect -13 -650 9 -615
rect 61 -650 83 -615
rect 135 -650 157 -615
rect 209 -650 231 -615
rect 283 -650 290 -598
rect -146 -657 290 -650
rect 607 -1122 809 -133
<< via2 >>
rect -116 -502 -87 -479
rect -87 -502 -65 -479
rect -65 -502 -13 -479
rect -13 -502 9 -479
rect 9 -502 61 -479
rect 61 -502 83 -479
rect 83 -502 135 -479
rect 135 -502 157 -479
rect 157 -502 209 -479
rect 209 -502 231 -479
rect 231 -502 260 -479
rect -116 -524 260 -502
rect -116 -576 -87 -524
rect -87 -576 -65 -524
rect -65 -576 -13 -524
rect -13 -576 9 -524
rect 9 -576 61 -524
rect 61 -576 83 -524
rect 83 -576 135 -524
rect 135 -576 157 -524
rect 157 -576 209 -524
rect 209 -576 231 -524
rect 231 -576 260 -524
rect -116 -598 260 -576
rect -116 -615 -87 -598
rect -87 -615 -65 -598
rect -65 -615 -13 -598
rect -13 -615 9 -598
rect 9 -615 61 -598
rect 61 -615 83 -598
rect 83 -615 135 -598
rect 135 -615 157 -598
rect 157 -615 209 -598
rect 209 -615 231 -598
rect 231 -615 260 -598
<< metal3 >>
rect -150 -479 290 -443
rect -150 -615 -116 -479
rect 260 -615 290 -479
rect -150 -657 290 -615
<< labels >>
flabel comment s 750 122 750 122 0 FreeSans 1600 0 0 0 S
flabel comment s -528 7380 -528 7380 0 FreeSans 1200 0 0 0 condiodeHvPsub
flabel comment s 62 122 62 122 0 FreeSans 1600 0 0 0 D
flabel comment s -589 122 -589 122 0 FreeSans 1600 0 0 0 S
<< properties >>
string GDS_END 10317996
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10046666
<< end >>
