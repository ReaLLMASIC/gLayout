magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect -977 -150 3243 3114
<< nwell >>
rect 21433 1533 21967 1865
rect 5542 -370 7172 534
rect 16656 -313 17407 59
rect -2662 -4241 -2217 -3540
rect -2393 -5555 -2061 -4912
rect -1889 -7074 -1395 -6642
<< pwell >>
rect -148 -10 -62 1305
rect 21649 1262 21927 1454
rect 16674 343 17246 391
rect 16674 342 17289 343
rect 16770 143 17289 342
rect -2581 -4538 -2303 -4346
rect -2561 -6794 -2303 -6734
rect -2767 -6986 -2303 -6794
<< scnmos >>
rect 16867 169 16897 317
rect 17176 169 17206 317
<< scpmoshvt >>
rect 16845 -201 16895 -1
rect 17154 -201 17204 -1
<< mvnmos >>
rect 21728 1288 21848 1428
rect -2502 -4512 -2382 -4372
rect -2685 -6960 -2565 -6820
rect -2482 -6960 -2382 -6760
<< mvpmos >>
rect 21552 1599 21672 1799
rect 21728 1599 21848 1799
rect -2502 -3906 -2382 -3706
rect -2502 -4174 -2382 -3974
rect -2327 -5260 -2127 -5140
rect -2327 -5436 -2127 -5316
rect -1770 -7008 -1670 -6708
rect -1614 -7008 -1514 -6708
<< ndiff >>
rect 16796 305 16867 317
rect 16796 271 16808 305
rect 16842 271 16867 305
rect 16796 215 16867 271
rect 16796 181 16808 215
rect 16842 181 16867 215
rect 16796 169 16867 181
rect 16897 305 16954 317
rect 16897 271 16908 305
rect 16942 271 16954 305
rect 16897 215 16954 271
rect 16897 181 16908 215
rect 16942 181 16954 215
rect 16897 169 16954 181
rect 17105 305 17176 317
rect 17105 271 17117 305
rect 17151 271 17176 305
rect 17105 215 17176 271
rect 17105 181 17117 215
rect 17151 181 17176 215
rect 17105 169 17176 181
rect 17206 305 17263 317
rect 17206 271 17217 305
rect 17251 271 17263 305
rect 17206 215 17263 271
rect 17206 181 17217 215
rect 17251 181 17263 215
rect 17206 169 17263 181
<< pdiff >>
rect 16776 -15 16845 -1
rect 16776 -49 16788 -15
rect 16822 -49 16845 -15
rect 16776 -85 16845 -49
rect 16776 -119 16788 -85
rect 16822 -119 16845 -85
rect 16776 -155 16845 -119
rect 16776 -189 16788 -155
rect 16822 -189 16845 -155
rect 16776 -201 16845 -189
rect 16895 -15 16954 -1
rect 16895 -49 16908 -15
rect 16942 -49 16954 -15
rect 16895 -85 16954 -49
rect 16895 -119 16908 -85
rect 16942 -119 16954 -85
rect 16895 -155 16954 -119
rect 16895 -189 16908 -155
rect 16942 -189 16954 -155
rect 16895 -201 16954 -189
rect 17085 -15 17154 -1
rect 17085 -49 17097 -15
rect 17131 -49 17154 -15
rect 17085 -85 17154 -49
rect 17085 -119 17097 -85
rect 17131 -119 17154 -85
rect 17085 -155 17154 -119
rect 17085 -189 17097 -155
rect 17131 -189 17154 -155
rect 17085 -201 17154 -189
rect 17204 -15 17263 -1
rect 17204 -49 17217 -15
rect 17251 -49 17263 -15
rect 17204 -85 17263 -49
rect 17204 -119 17217 -85
rect 17251 -119 17263 -85
rect 17204 -155 17263 -119
rect 17204 -189 17217 -155
rect 17251 -189 17263 -155
rect 17204 -201 17263 -189
<< mvndiff >>
rect 21675 1402 21728 1428
rect 21675 1368 21683 1402
rect 21717 1368 21728 1402
rect 21675 1334 21728 1368
rect 21675 1300 21683 1334
rect 21717 1300 21728 1334
rect 21675 1288 21728 1300
rect 21848 1402 21901 1428
rect 21848 1368 21859 1402
rect 21893 1368 21901 1402
rect 21848 1334 21901 1368
rect 21848 1300 21859 1334
rect 21893 1300 21901 1334
rect 21848 1288 21901 1300
rect -2555 -4384 -2502 -4372
rect -2555 -4418 -2547 -4384
rect -2513 -4418 -2502 -4384
rect -2555 -4452 -2502 -4418
rect -2555 -4486 -2547 -4452
rect -2513 -4486 -2502 -4452
rect -2555 -4512 -2502 -4486
rect -2382 -4384 -2329 -4372
rect -2382 -4418 -2371 -4384
rect -2337 -4418 -2329 -4384
rect -2382 -4452 -2329 -4418
rect -2382 -4486 -2371 -4452
rect -2337 -4486 -2329 -4452
rect -2382 -4512 -2329 -4486
rect -2535 -6772 -2482 -6760
rect -2535 -6806 -2527 -6772
rect -2493 -6806 -2482 -6772
rect -2535 -6820 -2482 -6806
rect -2741 -6846 -2685 -6820
rect -2741 -6880 -2730 -6846
rect -2696 -6880 -2685 -6846
rect -2741 -6914 -2685 -6880
rect -2741 -6948 -2730 -6914
rect -2696 -6948 -2685 -6914
rect -2741 -6960 -2685 -6948
rect -2565 -6840 -2482 -6820
rect -2565 -6874 -2527 -6840
rect -2493 -6874 -2482 -6840
rect -2565 -6908 -2482 -6874
rect -2565 -6942 -2527 -6908
rect -2493 -6942 -2482 -6908
rect -2565 -6960 -2482 -6942
rect -2382 -6772 -2329 -6760
rect -2382 -6806 -2371 -6772
rect -2337 -6806 -2329 -6772
rect -2382 -6840 -2329 -6806
rect -2382 -6874 -2371 -6840
rect -2337 -6874 -2329 -6840
rect -2382 -6908 -2329 -6874
rect -2382 -6942 -2371 -6908
rect -2337 -6942 -2329 -6908
rect -2382 -6960 -2329 -6942
<< mvpdiff >>
rect 21499 1781 21552 1799
rect 21499 1747 21507 1781
rect 21541 1747 21552 1781
rect 21499 1713 21552 1747
rect 21499 1679 21507 1713
rect 21541 1679 21552 1713
rect 21499 1645 21552 1679
rect 21499 1611 21507 1645
rect 21541 1611 21552 1645
rect 21499 1599 21552 1611
rect 21672 1781 21728 1799
rect 21672 1747 21683 1781
rect 21717 1747 21728 1781
rect 21672 1713 21728 1747
rect 21672 1679 21683 1713
rect 21717 1679 21728 1713
rect 21672 1645 21728 1679
rect 21672 1611 21683 1645
rect 21717 1611 21728 1645
rect 21672 1599 21728 1611
rect 21848 1781 21901 1799
rect 21848 1747 21859 1781
rect 21893 1747 21901 1781
rect 21848 1713 21901 1747
rect 21848 1679 21859 1713
rect 21893 1679 21901 1713
rect 21848 1645 21901 1679
rect 21848 1611 21859 1645
rect 21893 1611 21901 1645
rect 21848 1599 21901 1611
rect -2555 -3724 -2502 -3706
rect -2555 -3758 -2547 -3724
rect -2513 -3758 -2502 -3724
rect -2555 -3792 -2502 -3758
rect -2555 -3826 -2547 -3792
rect -2513 -3826 -2502 -3792
rect -2555 -3860 -2502 -3826
rect -2555 -3894 -2547 -3860
rect -2513 -3894 -2502 -3860
rect -2555 -3906 -2502 -3894
rect -2382 -3724 -2329 -3706
rect -2382 -3758 -2371 -3724
rect -2337 -3758 -2329 -3724
rect -2382 -3792 -2329 -3758
rect -2382 -3826 -2371 -3792
rect -2337 -3826 -2329 -3792
rect -2382 -3860 -2329 -3826
rect -2382 -3894 -2371 -3860
rect -2337 -3894 -2329 -3860
rect -2382 -3906 -2329 -3894
rect -2555 -3986 -2502 -3974
rect -2555 -4020 -2547 -3986
rect -2513 -4020 -2502 -3986
rect -2555 -4054 -2502 -4020
rect -2555 -4088 -2547 -4054
rect -2513 -4088 -2502 -4054
rect -2555 -4122 -2502 -4088
rect -2555 -4156 -2547 -4122
rect -2513 -4156 -2502 -4122
rect -2555 -4174 -2502 -4156
rect -2382 -3986 -2329 -3974
rect -2382 -4020 -2371 -3986
rect -2337 -4020 -2329 -3986
rect -2382 -4054 -2329 -4020
rect -2382 -4088 -2371 -4054
rect -2337 -4088 -2329 -4054
rect -2382 -4122 -2329 -4088
rect -2382 -4156 -2371 -4122
rect -2337 -4156 -2329 -4122
rect -2382 -4174 -2329 -4156
rect -2327 -5095 -2127 -5087
rect -2327 -5129 -2309 -5095
rect -2275 -5129 -2241 -5095
rect -2207 -5129 -2173 -5095
rect -2139 -5129 -2127 -5095
rect -2327 -5140 -2127 -5129
rect -2327 -5271 -2127 -5260
rect -2327 -5305 -2309 -5271
rect -2275 -5305 -2241 -5271
rect -2207 -5305 -2173 -5271
rect -2139 -5305 -2127 -5271
rect -2327 -5316 -2127 -5305
rect -2327 -5447 -2127 -5436
rect -2327 -5481 -2309 -5447
rect -2275 -5481 -2241 -5447
rect -2207 -5481 -2173 -5447
rect -2139 -5481 -2127 -5447
rect -2327 -5489 -2127 -5481
rect -1823 -6758 -1770 -6708
rect -1823 -6792 -1815 -6758
rect -1781 -6792 -1770 -6758
rect -1823 -6826 -1770 -6792
rect -1823 -6860 -1815 -6826
rect -1781 -6860 -1770 -6826
rect -1823 -6894 -1770 -6860
rect -1823 -6928 -1815 -6894
rect -1781 -6928 -1770 -6894
rect -1823 -6962 -1770 -6928
rect -1823 -6996 -1815 -6962
rect -1781 -6996 -1770 -6962
rect -1823 -7008 -1770 -6996
rect -1670 -6758 -1614 -6708
rect -1670 -6792 -1659 -6758
rect -1625 -6792 -1614 -6758
rect -1670 -6826 -1614 -6792
rect -1670 -6860 -1659 -6826
rect -1625 -6860 -1614 -6826
rect -1670 -6894 -1614 -6860
rect -1670 -6928 -1659 -6894
rect -1625 -6928 -1614 -6894
rect -1670 -6962 -1614 -6928
rect -1670 -6996 -1659 -6962
rect -1625 -6996 -1614 -6962
rect -1670 -7008 -1614 -6996
rect -1514 -6758 -1461 -6708
rect -1514 -6792 -1503 -6758
rect -1469 -6792 -1461 -6758
rect -1514 -6826 -1461 -6792
rect -1514 -6860 -1503 -6826
rect -1469 -6860 -1461 -6826
rect -1514 -6894 -1461 -6860
rect -1514 -6928 -1503 -6894
rect -1469 -6928 -1461 -6894
rect -1514 -6962 -1461 -6928
rect -1514 -6996 -1503 -6962
rect -1469 -6996 -1461 -6962
rect -1514 -7008 -1461 -6996
<< ndiffc >>
rect 16808 271 16842 305
rect 16808 181 16842 215
rect 16908 271 16942 305
rect 16908 181 16942 215
rect 17117 271 17151 305
rect 17117 181 17151 215
rect 17217 271 17251 305
rect 17217 181 17251 215
<< pdiffc >>
rect 16788 -49 16822 -15
rect 16788 -119 16822 -85
rect 16788 -189 16822 -155
rect 16908 -49 16942 -15
rect 16908 -119 16942 -85
rect 16908 -189 16942 -155
rect 17097 -49 17131 -15
rect 17097 -119 17131 -85
rect 17097 -189 17131 -155
rect 17217 -49 17251 -15
rect 17217 -119 17251 -85
rect 17217 -189 17251 -155
<< mvndiffc >>
rect 21683 1368 21717 1402
rect 21683 1300 21717 1334
rect 21859 1368 21893 1402
rect 21859 1300 21893 1334
rect -2547 -4418 -2513 -4384
rect -2547 -4486 -2513 -4452
rect -2371 -4418 -2337 -4384
rect -2371 -4486 -2337 -4452
rect -2527 -6806 -2493 -6772
rect -2730 -6880 -2696 -6846
rect -2730 -6948 -2696 -6914
rect -2527 -6874 -2493 -6840
rect -2527 -6942 -2493 -6908
rect -2371 -6806 -2337 -6772
rect -2371 -6874 -2337 -6840
rect -2371 -6942 -2337 -6908
<< mvpdiffc >>
rect 21507 1747 21541 1781
rect 21507 1679 21541 1713
rect 21507 1611 21541 1645
rect 21683 1747 21717 1781
rect 21683 1679 21717 1713
rect 21683 1611 21717 1645
rect 21859 1747 21893 1781
rect 21859 1679 21893 1713
rect 21859 1611 21893 1645
rect -2547 -3758 -2513 -3724
rect -2547 -3826 -2513 -3792
rect -2547 -3894 -2513 -3860
rect -2371 -3758 -2337 -3724
rect -2371 -3826 -2337 -3792
rect -2371 -3894 -2337 -3860
rect -2547 -4020 -2513 -3986
rect -2547 -4088 -2513 -4054
rect -2547 -4156 -2513 -4122
rect -2371 -4020 -2337 -3986
rect -2371 -4088 -2337 -4054
rect -2371 -4156 -2337 -4122
rect -2309 -5129 -2275 -5095
rect -2241 -5129 -2207 -5095
rect -2173 -5129 -2139 -5095
rect -2309 -5305 -2275 -5271
rect -2241 -5305 -2207 -5271
rect -2173 -5305 -2139 -5271
rect -2309 -5481 -2275 -5447
rect -2241 -5481 -2207 -5447
rect -2173 -5481 -2139 -5447
rect -1815 -6792 -1781 -6758
rect -1815 -6860 -1781 -6826
rect -1815 -6928 -1781 -6894
rect -1815 -6996 -1781 -6962
rect -1659 -6792 -1625 -6758
rect -1659 -6860 -1625 -6826
rect -1659 -6928 -1625 -6894
rect -1659 -6996 -1625 -6962
rect -1503 -6792 -1469 -6758
rect -1503 -6860 -1469 -6826
rect -1503 -6928 -1469 -6894
rect -1503 -6996 -1469 -6962
<< psubdiff >>
rect -122 1255 -88 1279
rect -122 1186 -88 1221
rect -122 1117 -88 1152
rect -122 1048 -88 1083
rect -122 979 -88 1014
rect -122 910 -88 945
rect -122 841 -88 876
rect -122 772 -88 807
rect -122 703 -88 738
rect -122 634 -88 669
rect -122 564 -88 600
rect -122 494 -88 530
rect -122 424 -88 460
rect -122 354 -88 390
rect -122 284 -88 320
rect -122 214 -88 250
rect -122 144 -88 180
rect -122 74 -88 110
rect -122 16 -88 40
<< nsubdiff >>
rect 17337 -1 17371 23
rect 17337 -73 17371 -35
rect 17337 -146 17371 -107
rect 17337 -219 17371 -180
rect 17337 -277 17371 -253
<< mvnsubdiff >>
rect -2327 -5012 -2303 -4978
rect -2269 -5012 -2185 -4978
rect -2151 -5012 -2127 -4978
<< psubdiffcont >>
rect -122 1221 -88 1255
rect -122 1152 -88 1186
rect -122 1083 -88 1117
rect -122 1014 -88 1048
rect -122 945 -88 979
rect -122 876 -88 910
rect -122 807 -88 841
rect -122 738 -88 772
rect -122 669 -88 703
rect -122 600 -88 634
rect -122 530 -88 564
rect -122 460 -88 494
rect -122 390 -88 424
rect -122 320 -88 354
rect -122 250 -88 284
rect -122 180 -88 214
rect -122 110 -88 144
rect -122 40 -88 74
<< nsubdiffcont >>
rect 17337 -35 17371 -1
rect 17337 -107 17371 -73
rect 17337 -180 17371 -146
rect 17337 -253 17371 -219
<< mvnsubdiffcont >>
rect -2303 -5012 -2269 -4978
rect -2185 -5012 -2151 -4978
<< poly >>
rect 21552 1799 21672 1825
rect 21728 1799 21848 1825
rect 21552 1557 21672 1599
rect 21728 1557 21848 1599
rect 21552 1528 21848 1557
rect 21552 1494 21574 1528
rect 21608 1494 21648 1528
rect 21682 1494 21721 1528
rect 21755 1494 21794 1528
rect 21828 1494 21848 1528
rect 21552 1460 21848 1494
rect 21728 1428 21848 1460
rect 21728 1256 21848 1288
rect 16867 317 16897 343
rect 17176 317 17206 343
rect 16867 131 16897 169
rect 17176 131 17206 169
rect 16723 115 16898 131
rect 16723 81 16739 115
rect 16773 81 16807 115
rect 16841 81 16898 115
rect 16723 65 16898 81
rect 17032 115 17207 131
rect 17032 81 17048 115
rect 17082 81 17116 115
rect 17150 81 17207 115
rect 17032 65 17207 81
rect 16845 38 16898 65
rect 17154 38 17207 65
rect 16845 -1 16895 38
rect 17154 -1 17204 38
rect 16845 -227 16895 -201
rect 17154 -227 17204 -201
rect -2502 -3706 -2382 -3680
rect -2502 -3974 -2382 -3906
rect -2502 -4222 -2382 -4174
rect -2502 -4256 -2460 -4222
rect -2426 -4256 -2382 -4222
rect -2502 -4290 -2382 -4256
rect -2502 -4324 -2460 -4290
rect -2426 -4324 -2382 -4290
rect -2502 -4372 -2382 -4324
rect -2502 -4538 -2382 -4512
rect -2425 -5178 -2327 -5140
rect -2425 -5212 -2409 -5178
rect -2375 -5212 -2327 -5178
rect -2425 -5247 -2327 -5212
rect -2425 -5281 -2409 -5247
rect -2375 -5260 -2327 -5247
rect -2127 -5260 -2095 -5140
rect -2375 -5281 -2359 -5260
rect -2425 -5316 -2359 -5281
rect -2425 -5350 -2409 -5316
rect -2375 -5350 -2327 -5316
rect -2425 -5386 -2327 -5350
rect -2425 -5420 -2409 -5386
rect -2375 -5420 -2327 -5386
rect -2425 -5436 -2327 -5420
rect -2127 -5436 -2095 -5316
rect -1770 -6708 -1670 -6676
rect -1614 -6708 -1514 -6676
rect -2482 -6760 -2382 -6728
rect -2685 -6820 -2565 -6788
rect -2685 -6992 -2565 -6960
rect -2699 -7008 -2565 -6992
rect -2699 -7042 -2683 -7008
rect -2649 -7042 -2615 -7008
rect -2581 -7042 -2565 -7008
rect -2699 -7058 -2565 -7042
rect -2482 -6992 -2382 -6960
rect -2482 -7008 -2348 -6992
rect -2482 -7042 -2466 -7008
rect -2432 -7042 -2398 -7008
rect -2364 -7042 -2348 -7008
rect -2482 -7058 -2348 -7042
rect -1770 -7040 -1670 -7008
rect -1614 -7040 -1514 -7008
rect -1770 -7056 -1513 -7040
rect -1770 -7090 -1754 -7056
rect -1720 -7090 -1659 -7056
rect -1625 -7090 -1563 -7056
rect -1529 -7090 -1513 -7056
rect -1770 -7106 -1513 -7090
<< polycont >>
rect 21574 1494 21608 1528
rect 21648 1494 21682 1528
rect 21721 1494 21755 1528
rect 21794 1494 21828 1528
rect 16739 81 16773 115
rect 16807 81 16841 115
rect 17048 81 17082 115
rect 17116 81 17150 115
rect -2460 -4256 -2426 -4222
rect -2460 -4324 -2426 -4290
rect -2409 -5212 -2375 -5178
rect -2409 -5281 -2375 -5247
rect -2409 -5350 -2375 -5316
rect -2409 -5420 -2375 -5386
rect -2683 -7042 -2649 -7008
rect -2615 -7042 -2581 -7008
rect -2466 -7042 -2432 -7008
rect -2398 -7042 -2364 -7008
rect -1754 -7090 -1720 -7056
rect -1659 -7090 -1625 -7056
rect -1563 -7090 -1529 -7056
<< locali >>
rect -122 2565 -88 2606
rect -122 2490 -88 2531
rect -122 2415 -88 2456
rect -122 2340 -88 2381
rect -122 2265 -88 2306
rect -122 2190 -88 2231
rect -122 2115 -88 2156
rect -122 2039 -88 2081
rect -122 1963 -88 2005
rect -122 1887 -88 1929
rect -122 1811 -88 1853
rect -122 1735 -88 1777
rect -122 1659 -88 1701
rect -122 1583 -88 1625
rect 21507 1781 21541 1797
rect 21507 1713 21541 1747
rect 21507 1645 21541 1679
rect 21507 1595 21541 1611
rect 21683 1781 21729 1797
rect 21717 1747 21729 1781
rect 21683 1713 21729 1747
rect 21717 1702 21729 1713
rect 21683 1668 21695 1679
rect 21683 1645 21729 1668
rect 21717 1630 21729 1645
rect 21683 1596 21695 1611
rect 21859 1781 21893 1797
rect 21859 1713 21893 1747
rect 21859 1645 21893 1679
rect 21683 1595 21717 1596
rect 21859 1595 21893 1611
rect -122 1507 -88 1549
rect 21608 1494 21630 1528
rect 21682 1494 21721 1528
rect 21755 1494 21794 1528
rect 21828 1494 21844 1528
rect -122 1431 -88 1473
rect 21683 1409 21717 1418
rect 21698 1402 21717 1409
rect 21664 1368 21683 1375
rect 21664 1337 21717 1368
rect 21698 1334 21717 1337
rect 21683 1284 21717 1300
rect 21859 1402 21893 1418
rect 21859 1334 21893 1368
rect 21859 1284 21893 1300
rect -122 1267 -88 1279
rect -122 1192 -88 1221
rect -122 1117 -88 1152
rect -122 1048 -88 1083
rect -122 979 -88 1008
rect -122 910 -88 933
rect -122 841 -88 858
rect 19678 1225 19726 1259
rect 19760 1225 19808 1259
rect 19842 1225 19889 1259
rect 19923 1225 19970 1259
rect 20004 1225 20051 1259
rect 20085 1225 20132 1259
rect 20 1149 54 1203
rect 20 1061 54 1115
rect 20 972 54 1027
rect 20 883 54 938
rect -122 772 -88 783
rect -122 703 -88 708
rect -122 666 -88 669
rect -122 590 -88 600
rect -122 514 -88 530
rect -122 438 -88 460
rect -122 362 -88 390
rect 20 681 54 735
rect 20 593 54 647
rect 20 504 54 559
rect 20 415 54 470
rect 6621 522 7093 534
rect 6621 488 6626 522
rect 6660 488 7093 522
rect 5885 430 5935 464
rect 5969 430 6018 464
rect 6621 451 7093 488
rect 6621 450 6791 451
rect 6621 416 6626 450
rect 6660 416 6791 450
rect 7018 425 7093 451
rect 16690 342 16725 376
rect 16759 342 16816 376
rect 16850 342 16865 376
rect 16999 342 17034 376
rect 17068 342 17125 376
rect 17159 342 17174 376
rect -122 286 -88 320
rect -122 214 -88 250
rect -122 144 -88 176
rect 16791 305 16857 342
rect 16791 271 16808 305
rect 16842 271 16857 305
rect 16791 215 16857 271
rect 16791 181 16808 215
rect 16842 181 16857 215
rect 16791 165 16857 181
rect 16892 305 16958 321
rect 16892 271 16908 305
rect 16942 271 16958 305
rect 16892 215 16958 271
rect 16892 181 16908 215
rect 16942 181 16958 215
rect 16892 131 16958 181
rect 17100 305 17166 342
rect 17100 271 17117 305
rect 17151 271 17166 305
rect 17100 215 17166 271
rect 17100 181 17117 215
rect 17151 181 17166 215
rect 17100 165 17166 181
rect 17201 305 17267 321
rect 17201 271 17217 305
rect 17251 271 17267 305
rect 17201 237 17267 271
rect 17201 203 17213 237
rect 17247 215 17285 237
rect 17251 203 17285 215
rect 17201 181 17217 203
rect 17251 181 17267 203
rect -122 74 -88 100
rect 16719 115 16857 131
rect 16719 81 16739 115
rect 16773 81 16807 115
rect 16841 81 16857 115
rect 16719 35 16857 81
rect 16892 125 17166 131
rect 16892 91 16970 125
rect 17004 91 17042 125
rect 17076 115 17166 125
rect 16892 81 17048 91
rect 17082 81 17116 115
rect 17150 81 17166 115
rect 16892 35 17166 81
rect -122 16 -88 24
rect 16772 -15 16838 1
rect 16772 -49 16788 -15
rect 16822 -49 16838 -15
rect 6460 -105 6990 -74
rect 6460 -139 6472 -105
rect 6506 -139 6551 -105
rect 6585 -139 6990 -105
rect 6460 -170 6990 -139
rect 16772 -85 16838 -49
rect 16772 -119 16788 -85
rect 16822 -119 16838 -85
rect 16772 -155 16838 -119
rect 16772 -189 16788 -155
rect 16822 -189 16838 -155
rect 16772 -248 16838 -189
rect 16892 -15 16958 35
rect 16892 -49 16908 -15
rect 16942 -49 16958 -15
rect 16892 -85 16958 -49
rect 16892 -119 16908 -85
rect 16942 -119 16958 -85
rect 16892 -155 16958 -119
rect 16892 -189 16908 -155
rect 16942 -189 16958 -155
rect 16892 -205 16958 -189
rect 17081 -15 17147 1
rect 17081 -49 17097 -15
rect 17131 -49 17147 -15
rect 17081 -85 17147 -49
rect 17081 -119 17097 -85
rect 17131 -119 17147 -85
rect 17081 -155 17147 -119
rect 17081 -189 17097 -155
rect 17131 -189 17147 -155
rect 17081 -248 17147 -189
rect 17201 -15 17267 181
rect 17201 -49 17217 -15
rect 17251 -49 17267 -15
rect 17201 -85 17267 -49
rect 17201 -119 17217 -85
rect 17251 -119 17267 -85
rect 17201 -155 17267 -119
rect 17201 -189 17217 -155
rect 17251 -189 17267 -155
rect 17201 -205 17267 -189
rect 17337 -1 17403 23
rect 17371 -35 17403 -1
rect 17337 -73 17403 -35
rect 17371 -107 17403 -73
rect 17337 -146 17403 -107
rect 17371 -180 17403 -146
rect 17337 -219 17403 -180
rect 16674 -253 17337 -248
rect 17371 -253 17403 -219
rect 16674 -255 17403 -253
rect 16674 -289 16717 -255
rect 16751 -289 16797 -255
rect 16831 -289 16877 -255
rect 16911 -289 16956 -255
rect 16990 -289 17035 -255
rect 17069 -289 17114 -255
rect 17148 -289 17193 -255
rect 17227 -289 17272 -255
rect 17306 -289 17403 -255
rect 16674 -327 17403 -289
rect -2547 -3724 -2513 -3706
rect -2547 -3792 -2513 -3758
rect -2547 -3860 -2513 -3826
rect -2547 -3986 -2513 -3894
rect -2547 -4049 -2513 -4020
rect -2547 -4121 -2513 -4088
rect -2547 -4384 -2513 -4156
rect -2371 -3724 -2337 -3712
rect -2371 -3792 -2337 -3784
rect -2371 -3860 -2337 -3826
rect -2371 -3986 -2337 -3894
rect -2371 -4054 -2337 -4020
rect -2371 -4122 -2337 -4088
rect -2371 -4172 -2337 -4156
rect -2476 -4256 -2460 -4222
rect -2416 -4251 -2410 -4222
rect -2426 -4256 -2410 -4251
rect -2476 -4289 -2410 -4256
rect -2476 -4290 -2450 -4289
rect -2476 -4324 -2460 -4290
rect -2416 -4323 -2410 -4289
rect -2426 -4324 -2410 -4323
rect -2547 -4452 -2513 -4418
rect -2547 -4502 -2513 -4486
rect -2371 -4384 -2337 -4368
rect -2371 -4429 -2337 -4418
rect -2371 -4501 -2337 -4486
rect -2327 -5012 -2303 -4978
rect -2269 -5012 -2259 -4978
rect -2225 -5012 -2187 -4978
rect -2151 -5012 -2127 -4978
rect -2311 -5129 -2309 -5095
rect -2275 -5129 -2273 -5095
rect -2207 -5129 -2173 -5095
rect -2139 -5129 -2123 -5095
rect -2409 -5178 -2375 -5162
rect -2409 -5247 -2375 -5219
rect -2409 -5316 -2375 -5291
rect -2325 -5305 -2309 -5271
rect -2275 -5305 -2262 -5271
rect -2207 -5305 -2190 -5271
rect -2139 -5305 -2123 -5271
rect -2409 -5386 -2375 -5350
rect -2409 -5436 -2375 -5420
rect -2325 -5481 -2309 -5447
rect -2267 -5481 -2241 -5447
rect -2195 -5481 -2173 -5447
rect -2139 -5481 -2123 -5447
rect -2553 -6772 -2493 -6756
rect -2553 -6812 -2527 -6772
rect -2730 -6842 -2696 -6830
rect -2730 -6914 -2696 -6880
rect -2730 -6964 -2696 -6948
rect -2553 -6840 -2493 -6812
rect -2553 -6884 -2527 -6840
rect -2553 -6908 -2493 -6884
rect -2553 -6942 -2527 -6908
rect -2553 -6958 -2493 -6942
rect -2371 -6772 -2337 -6756
rect -2371 -6840 -2337 -6812
rect -2371 -6908 -2337 -6884
rect -2371 -6958 -2337 -6942
rect -1815 -6758 -1781 -6742
rect -1815 -6826 -1781 -6812
rect -1815 -6894 -1781 -6884
rect -1815 -6962 -1781 -6928
rect -1659 -6758 -1625 -6742
rect -1659 -6826 -1625 -6792
rect -1659 -6894 -1625 -6860
rect -1659 -6932 -1625 -6928
rect -1503 -6758 -1469 -6742
rect -1503 -6826 -1469 -6812
rect -1503 -6894 -1469 -6884
rect -1657 -6962 -1619 -6932
rect -1625 -6966 -1619 -6962
rect -1503 -6962 -1469 -6928
rect -2699 -7042 -2687 -7008
rect -2649 -7042 -2615 -7008
rect -2581 -7042 -2565 -7008
rect -2482 -7042 -2470 -7008
rect -2432 -7042 -2398 -7008
rect -2364 -7042 -2348 -7008
rect -1815 -7012 -1781 -6996
rect -1659 -7012 -1625 -6996
rect -1503 -7012 -1469 -6996
rect -1770 -7090 -1758 -7056
rect -1720 -7090 -1659 -7056
rect -1625 -7090 -1563 -7056
rect -1525 -7090 -1513 -7056
<< viali >>
rect -122 2606 -88 2640
rect -122 2531 -88 2565
rect -122 2456 -88 2490
rect -122 2381 -88 2415
rect -122 2306 -88 2340
rect -122 2231 -88 2265
rect -122 2156 -88 2190
rect -122 2081 -88 2115
rect -122 2005 -88 2039
rect -122 1929 -88 1963
rect -122 1853 -88 1887
rect -122 1777 -88 1811
rect -122 1701 -88 1735
rect -122 1625 -88 1659
rect 21695 1679 21717 1702
rect 21717 1679 21729 1702
rect 21695 1668 21729 1679
rect 21695 1611 21717 1630
rect 21717 1611 21729 1630
rect 21695 1596 21729 1611
rect -122 1549 -88 1583
rect -122 1473 -88 1507
rect 21558 1494 21574 1528
rect 21574 1494 21592 1528
rect 21630 1494 21648 1528
rect 21648 1494 21664 1528
rect -122 1397 -88 1431
rect 21664 1402 21698 1409
rect 21664 1375 21683 1402
rect 21683 1375 21698 1402
rect 21664 1334 21698 1337
rect 21664 1303 21683 1334
rect 21683 1303 21698 1334
rect -122 1255 -88 1267
rect -122 1233 -88 1255
rect -122 1186 -88 1192
rect -122 1158 -88 1186
rect -122 1083 -88 1117
rect -122 1014 -88 1042
rect -122 1008 -88 1014
rect -122 945 -88 967
rect -122 933 -88 945
rect -122 876 -88 892
rect -122 858 -88 876
rect 20 1203 54 1237
rect 19644 1225 19678 1259
rect 19726 1225 19760 1259
rect 19808 1225 19842 1259
rect 19889 1225 19923 1259
rect 19970 1225 20004 1259
rect 20051 1225 20085 1259
rect 20132 1225 20166 1259
rect 20 1115 54 1149
rect 20 1027 54 1061
rect 20 938 54 972
rect 20 849 54 883
rect -122 807 -88 817
rect -122 783 -88 807
rect -122 738 -88 742
rect -122 708 -88 738
rect -122 634 -88 666
rect -122 632 -88 634
rect -122 564 -88 590
rect -122 556 -88 564
rect -122 494 -88 514
rect -122 480 -88 494
rect -122 424 -88 438
rect -122 404 -88 424
rect 20 735 54 769
rect 20 647 54 681
rect 20 559 54 593
rect 20 470 54 504
rect 6626 488 6660 522
rect 5851 430 5885 464
rect 5935 430 5969 464
rect 6018 430 6052 464
rect 6626 416 6660 450
rect 20 381 54 415
rect -122 354 -88 362
rect -122 328 -88 354
rect 16725 342 16759 376
rect 16816 342 16850 376
rect 17034 342 17068 376
rect 17125 342 17159 376
rect -122 284 -88 286
rect -122 252 -88 284
rect -122 180 -88 210
rect -122 176 -88 180
rect -122 110 -88 134
rect 17213 215 17247 237
rect 17213 203 17217 215
rect 17217 203 17247 215
rect 17285 203 17319 237
rect -122 100 -88 110
rect -122 40 -88 58
rect -122 24 -88 40
rect 16970 91 17004 125
rect 17042 115 17076 125
rect 17042 91 17048 115
rect 17048 91 17076 115
rect 6472 -139 6506 -105
rect 6551 -139 6585 -105
rect 16717 -289 16751 -255
rect 16797 -289 16831 -255
rect 16877 -289 16911 -255
rect 16956 -289 16990 -255
rect 17035 -289 17069 -255
rect 17114 -289 17148 -255
rect 17193 -289 17227 -255
rect 17272 -289 17306 -255
rect -2547 -4054 -2513 -4049
rect -2547 -4083 -2513 -4054
rect -2547 -4122 -2513 -4121
rect -2547 -4155 -2513 -4122
rect -2371 -3712 -2337 -3678
rect -2371 -3758 -2337 -3750
rect -2371 -3784 -2337 -3758
rect -2450 -4222 -2416 -4217
rect -2450 -4251 -2426 -4222
rect -2426 -4251 -2416 -4222
rect -2450 -4290 -2416 -4289
rect -2450 -4323 -2426 -4290
rect -2426 -4323 -2416 -4290
rect -2371 -4452 -2337 -4429
rect -2371 -4463 -2337 -4452
rect -2371 -4535 -2337 -4501
rect -2259 -5012 -2225 -4978
rect -2187 -5012 -2185 -4978
rect -2185 -5012 -2153 -4978
rect -2345 -5129 -2311 -5095
rect -2273 -5129 -2241 -5095
rect -2241 -5129 -2239 -5095
rect -2409 -5212 -2375 -5185
rect -2409 -5219 -2375 -5212
rect -2409 -5281 -2375 -5257
rect -2409 -5291 -2375 -5281
rect -2262 -5305 -2241 -5271
rect -2241 -5305 -2228 -5271
rect -2190 -5305 -2173 -5271
rect -2173 -5305 -2156 -5271
rect -2301 -5481 -2275 -5447
rect -2275 -5481 -2267 -5447
rect -2229 -5481 -2207 -5447
rect -2207 -5481 -2195 -5447
rect -2527 -6806 -2493 -6778
rect -2527 -6812 -2493 -6806
rect -2730 -6846 -2696 -6842
rect -2730 -6876 -2696 -6846
rect -2730 -6948 -2696 -6914
rect -2527 -6874 -2493 -6850
rect -2527 -6884 -2493 -6874
rect -2371 -6806 -2337 -6778
rect -2371 -6812 -2337 -6806
rect -2371 -6874 -2337 -6850
rect -2371 -6884 -2337 -6874
rect -1815 -6792 -1781 -6778
rect -1815 -6812 -1781 -6792
rect -1815 -6860 -1781 -6850
rect -1815 -6884 -1781 -6860
rect -1503 -6792 -1469 -6778
rect -1503 -6812 -1469 -6792
rect -1503 -6860 -1469 -6850
rect -1503 -6884 -1469 -6860
rect -1691 -6962 -1657 -6932
rect -1691 -6966 -1659 -6962
rect -1659 -6966 -1657 -6962
rect -1619 -6966 -1585 -6932
rect -2687 -7042 -2683 -7008
rect -2683 -7042 -2653 -7008
rect -2615 -7042 -2581 -7008
rect -2470 -7042 -2466 -7008
rect -2466 -7042 -2436 -7008
rect -2398 -7042 -2364 -7008
rect -1758 -7090 -1754 -7056
rect -1754 -7090 -1724 -7056
rect -1659 -7090 -1625 -7056
rect -1559 -7090 -1529 -7056
rect -1529 -7090 -1525 -7056
<< metal1 >>
rect -128 2640 -82 2652
rect -128 2606 -122 2640
rect -88 2606 -82 2640
rect -128 2565 -82 2606
rect -128 2531 -122 2565
rect -88 2531 -82 2565
rect -128 2490 -82 2531
rect -128 2456 -122 2490
rect -88 2456 -82 2490
rect -128 2415 -82 2456
rect -128 2381 -122 2415
rect -88 2381 -82 2415
rect -128 2340 -82 2381
rect -128 2306 -122 2340
rect -88 2306 -82 2340
rect -128 2265 -82 2306
rect -128 2231 -122 2265
rect -88 2231 -82 2265
rect -128 2190 -82 2231
rect -128 2156 -122 2190
rect -88 2156 -82 2190
rect -128 2115 -82 2156
rect -128 2081 -122 2115
rect -88 2081 -82 2115
rect -128 2039 -82 2081
rect -128 2005 -122 2039
rect -88 2005 -82 2039
rect -128 1963 -82 2005
rect -128 1929 -122 1963
rect -88 1929 -82 1963
rect -128 1887 -82 1929
rect -128 1853 -122 1887
rect -88 1853 -82 1887
rect -971 1823 -919 1829
rect -3128 1733 -3122 1785
rect -3070 1733 -3058 1785
rect -3006 1733 -1262 1785
rect -1210 1733 -1198 1785
rect -1146 1733 -1140 1785
rect -971 1759 -919 1771
rect -971 1701 -919 1707
rect -128 1811 -82 1853
rect -128 1777 -122 1811
rect -88 1777 -82 1811
rect -128 1735 -82 1777
rect -128 1701 -122 1735
rect -88 1701 -82 1735
rect -128 1659 -82 1701
rect -128 1625 -122 1659
rect -88 1625 -82 1659
rect 21689 1702 21778 1714
rect 21689 1668 21695 1702
rect 21729 1668 21778 1702
rect -3072 1600 -1262 1606
rect -3020 1554 -1262 1600
rect -1210 1554 -1198 1606
rect -1146 1554 -1140 1606
rect -128 1583 -82 1625
rect 18588 1622 18630 1649
rect 21689 1630 21778 1668
rect -3072 1536 -3020 1548
rect -3072 1478 -3020 1484
rect -128 1549 -122 1583
rect -88 1549 -82 1583
rect 21689 1596 21695 1630
rect 21729 1596 21778 1630
rect 21689 1584 21778 1596
tri 21689 1571 21702 1584 ne
rect 21702 1571 21778 1584
rect -128 1530 -82 1549
rect -128 1507 -48 1530
rect -128 1473 -122 1507
rect -88 1500 -48 1507
rect -88 1473 -82 1500
rect -128 1431 -82 1473
rect 19176 1437 19309 1571
tri 21702 1563 21710 1571 ne
rect 21548 1534 21554 1550
rect 21546 1498 21554 1534
rect 21606 1498 21618 1550
rect 21670 1498 21676 1550
rect 21546 1494 21558 1498
rect 21592 1494 21630 1498
rect 21664 1494 21676 1498
rect 21546 1488 21676 1494
tri 21693 1456 21710 1473 se
rect 21710 1456 21778 1571
rect 20969 1450 21021 1456
rect -128 1397 -122 1431
rect -88 1397 -82 1431
rect -128 1267 -82 1397
rect 20969 1386 21021 1398
rect 19182 1321 19188 1373
rect 19240 1321 19252 1373
rect 19304 1321 19310 1373
rect 20969 1328 21021 1334
rect 21322 1450 21374 1456
rect 21322 1386 21374 1398
rect 21322 1328 21374 1334
tri 21658 1421 21693 1456 se
rect 21693 1421 21778 1456
rect 21658 1409 21778 1421
rect 21658 1408 21664 1409
rect 21698 1408 21778 1409
rect 21710 1356 21778 1408
rect 21658 1342 21778 1356
rect 21710 1290 21778 1342
rect 21658 1284 21778 1290
rect -128 1233 -122 1267
rect -88 1233 -82 1267
rect 19670 1265 19676 1270
rect 19632 1259 19676 1265
rect 19728 1259 19740 1270
rect 19792 1265 19798 1270
rect 19792 1259 20178 1265
rect -128 1192 -82 1233
rect -128 1158 -122 1192
rect -88 1158 -82 1192
rect -128 1117 -82 1158
rect -128 1083 -122 1117
rect -88 1083 -82 1117
rect -128 1042 -82 1083
rect -128 1008 -122 1042
rect -88 1008 -82 1042
rect -128 967 -82 1008
rect -128 933 -122 967
rect -88 933 -82 967
rect -128 892 -82 933
rect -128 858 -122 892
rect -88 858 -82 892
rect -128 817 -82 858
rect 14 1237 60 1249
rect 14 1203 20 1237
rect 54 1203 60 1237
rect 19632 1225 19644 1259
rect 19792 1225 19808 1259
rect 19842 1225 19889 1259
rect 19923 1225 19970 1259
rect 20004 1225 20051 1259
rect 20085 1225 20132 1259
rect 20166 1225 20178 1259
rect 19632 1219 19676 1225
rect 19670 1218 19676 1219
rect 19728 1218 19740 1225
rect 19792 1219 20178 1225
rect 19792 1218 19798 1219
rect 14 1149 60 1203
rect 14 1115 20 1149
rect 54 1115 60 1149
rect 14 1061 60 1115
rect 14 1027 20 1061
rect 54 1027 60 1061
rect 14 972 60 1027
rect 14 938 20 972
rect 54 938 60 972
rect 14 883 60 938
tri 21116 910 21160 954 se
rect 21160 921 21387 954
rect 14 849 20 883
rect 54 849 60 883
rect 14 837 60 849
tri 60 837 133 910 sw
tri 21114 908 21116 910 se
rect 21116 908 21160 910
tri 21160 908 21173 921 nw
tri 21110 904 21114 908 se
rect 21114 904 21156 908
tri 21156 904 21160 908 nw
tri 20344 839 20409 904 se
rect 20409 871 21123 904
tri 21123 871 21156 904 nw
rect 21381 902 21387 921
rect 21439 902 21451 954
rect 21503 902 21509 954
tri 20409 839 20441 871 nw
tri 20342 837 20344 839 se
rect -128 783 -122 817
rect -88 783 -82 817
tri 60 801 96 837 ne
rect 96 822 133 837
tri 133 822 148 837 sw
rect -128 742 -82 783
rect -128 708 -122 742
rect -88 708 -82 742
rect -128 666 -82 708
rect -128 632 -122 666
rect -88 632 -82 666
rect -128 590 -82 632
rect -128 556 -122 590
rect -88 556 -82 590
rect -128 514 -82 556
rect -128 480 -122 514
rect -88 480 -82 514
rect -128 438 -82 480
rect -128 404 -122 438
rect -88 404 -82 438
rect -128 362 -82 404
rect 14 769 60 781
rect 14 735 20 769
rect 54 735 60 769
rect 14 681 60 735
rect 14 647 20 681
rect 54 647 60 681
rect 14 593 60 647
rect 14 559 20 593
rect 54 559 60 593
rect 14 504 60 559
rect 96 650 148 822
tri 20279 774 20342 837 se
rect 20342 774 20344 837
tri 20344 774 20409 839 nw
tri 20261 756 20279 774 se
rect 20279 756 20326 774
tri 20326 756 20344 774 nw
rect 20241 725 20295 756
tri 20295 725 20326 756 nw
rect 18624 673 18630 725
rect 18682 673 18694 725
rect 18746 673 18752 725
rect 18954 673 18960 725
rect 19012 673 19024 725
rect 19076 673 19082 725
rect 20241 717 20287 725
tri 20287 717 20295 725 nw
rect 20241 673 20243 717
tri 20243 673 20287 717 nw
tri 21239 673 21283 717 se
rect 21283 673 21431 717
tri 20241 671 20243 673 nw
tri 21237 671 21239 673 se
rect 21239 671 21431 673
tri 21231 665 21237 671 se
rect 21237 665 21431 671
rect 21483 665 21495 717
rect 21547 665 21553 717
tri 21192 626 21231 665 se
rect 21231 626 21243 665
rect 96 586 148 598
rect 19086 574 19092 626
rect 19144 574 19156 626
rect 19208 574 19214 626
tri 21169 603 21192 626 se
rect 21192 603 21243 626
tri 21243 603 21305 665 nw
tri 21140 574 21169 603 se
tri 21100 534 21140 574 se
rect 21140 534 21169 574
rect 96 528 148 534
rect 14 490 20 504
rect 54 496 60 504
rect 6620 522 6666 534
tri 21095 529 21100 534 se
rect 21100 529 21169 534
tri 21169 529 21243 603 nw
rect 54 490 66 496
rect 6620 488 6626 522
rect 6660 488 6666 522
rect 5969 470 6096 473
rect 14 426 66 438
rect 5839 464 6096 470
rect 5839 430 5851 464
rect 5885 430 5935 464
rect 5969 430 6018 464
rect 6052 430 6096 464
rect 5839 424 6096 430
rect 5969 421 6096 424
tri 6001 416 6006 421 ne
rect 6006 416 6096 421
tri 6006 393 6029 416 ne
rect 14 368 66 374
rect -128 328 -122 362
rect -88 328 -82 362
rect -128 286 -82 328
rect -128 252 -122 286
rect -88 252 -82 286
rect -128 210 -82 252
rect -128 176 -122 210
rect -88 176 -82 210
rect -128 134 -82 176
rect -128 100 -122 134
rect -88 100 -82 134
rect -128 58 -82 100
rect -128 24 -122 58
rect -88 24 -82 58
rect -128 12 -82 24
rect -54 75 -2 81
rect -54 11 -2 23
rect -1257 -9 -1251 6
rect -2800 -15 -1251 -9
rect -2748 -45 -1251 -15
rect -1257 -46 -1251 -45
rect -1199 -46 -1187 6
rect -1135 -46 -1129 6
rect -54 -47 -2 -41
rect 32 -7 84 -1
rect -2800 -79 -2748 -67
rect 32 -71 84 -59
rect -2800 -137 -2748 -131
rect -2716 -82 -1251 -76
rect -2664 -112 -1251 -82
rect -1257 -128 -1251 -112
rect -1199 -128 -1187 -76
rect -1135 -128 -1129 -76
rect 382 -100 420 -47
rect 747 -106 798 -49
rect 32 -129 84 -123
rect -2716 -146 -2664 -134
rect -2716 -204 -2664 -198
rect -2593 -231 -1129 -205
rect -2593 -235 -1251 -231
rect -2987 -241 -1251 -235
rect -2935 -271 -2557 -241
rect -1257 -283 -1251 -241
rect -1199 -283 -1187 -231
rect -1135 -283 -1129 -231
rect 6029 -251 6096 416
rect 6620 450 6666 488
tri 21021 455 21095 529 se
tri 21095 455 21169 529 nw
rect 6620 416 6626 450
rect 6660 416 6666 450
tri 21006 440 21021 455 se
rect 6367 342 6413 352
tri 6413 342 6423 352 sw
rect 6367 329 6423 342
tri 6423 329 6436 342 sw
rect 6367 307 6436 329
tri 6436 307 6458 329 sw
tri 6598 307 6620 329 se
rect 6620 307 6666 416
rect 16674 376 16919 440
rect 16674 342 16725 376
rect 16759 342 16816 376
rect 16850 342 16919 376
rect 16674 330 16919 342
rect 16983 376 17228 440
tri 20959 393 21006 440 se
rect 21006 393 21021 440
rect 18086 385 18092 393
rect 16983 342 17034 376
rect 17068 342 17125 376
rect 17159 342 17228 376
tri 17558 363 17580 385 se
rect 17580 363 18092 385
tri 17460 349 17474 363 se
rect 17474 349 18092 363
rect 16983 330 17228 342
tri 17452 341 17460 349 se
rect 17460 341 17586 349
tri 17586 341 17594 349 nw
rect 18086 341 18092 349
rect 18144 341 18156 393
rect 18208 341 18214 393
tri 20947 381 20959 393 se
rect 20959 381 21021 393
tri 21021 381 21095 455 nw
tri 20907 341 20947 381 se
tri 17441 330 17452 341 se
rect 17452 330 17572 341
tri 17419 308 17441 330 se
rect 17441 327 17572 330
tri 17572 327 17586 341 nw
tri 20893 327 20907 341 se
rect 20907 327 20947 341
rect 17441 308 17474 327
tri 17474 308 17493 327 nw
tri 20874 308 20893 327 se
rect 20893 308 20947 327
tri 17418 307 17419 308 se
rect 17419 307 17473 308
tri 17473 307 17474 308 nw
tri 20873 307 20874 308 se
rect 20874 307 20947 308
tri 20947 307 21021 381 nw
rect 6367 305 6458 307
tri 6458 305 6460 307 sw
tri 6596 305 6598 307 se
rect 6598 305 6666 307
rect 6367 282 6666 305
tri 17402 291 17418 307 se
rect 17418 291 17457 307
tri 17457 291 17473 307 nw
rect 18083 291 18089 307
rect 6367 273 6657 282
tri 6657 273 6666 282 nw
tri 17384 273 17402 291 se
rect 17402 273 17430 291
tri 6367 251 6389 273 ne
rect 6389 251 6635 273
tri 6635 251 6657 273 nw
tri 17364 253 17384 273 se
rect 17384 264 17430 273
tri 17430 264 17457 291 nw
tri 17474 264 17501 291 se
rect 17501 264 18089 291
rect 17384 253 17419 264
tri 17419 253 17430 264 nw
tri 17463 253 17474 264 se
rect 17474 255 18089 264
rect 18141 255 18154 307
rect 18206 255 18212 307
tri 20821 255 20873 307 se
rect 17474 253 17501 255
tri 17362 251 17364 253 se
rect 17364 251 17409 253
tri 6432 241 6442 251 ne
rect 6442 241 6625 251
tri 6625 241 6635 251 nw
tri 17354 243 17362 251 se
rect 17362 243 17409 251
tri 17409 243 17419 253 nw
tri 17453 243 17463 253 se
rect 17463 243 17501 253
rect 17201 241 17407 243
tri 17407 241 17409 243 nw
tri 17451 241 17453 243 se
rect 17453 241 17501 243
tri 17501 241 17515 255 nw
tri 20807 241 20821 255 se
rect 20821 241 20873 255
tri 6442 237 6446 241 ne
rect 6446 237 6621 241
tri 6621 237 6625 241 nw
rect 17201 237 17399 241
tri 6446 233 6450 237 ne
rect 6450 233 6617 237
tri 6617 233 6621 237 nw
tri 6450 223 6460 233 ne
rect 6460 223 6607 233
tri 6607 223 6617 233 nw
rect 6460 -105 6597 223
tri 6597 213 6607 223 nw
rect 17201 203 17213 237
rect 17247 203 17285 237
rect 17319 233 17399 237
tri 17399 233 17407 241 nw
tri 17443 233 17451 241 se
rect 17451 233 17493 241
tri 17493 233 17501 241 nw
tri 20799 233 20807 241 se
rect 20807 233 20873 241
tri 20873 233 20947 307 nw
rect 17319 211 17377 233
tri 17377 211 17399 233 nw
tri 17421 211 17443 233 se
rect 17443 211 17471 233
tri 17471 211 17493 233 nw
tri 20777 211 20799 233 se
rect 17319 203 17365 211
rect 17201 199 17365 203
tri 17365 199 17377 211 nw
tri 17409 199 17421 211 se
rect 17421 199 17451 211
rect 17201 197 17363 199
tri 17363 197 17365 199 nw
tri 17407 197 17409 199 se
rect 17409 197 17451 199
tri 17401 191 17407 197 se
rect 17407 191 17451 197
tri 17451 191 17471 211 nw
tri 17375 165 17401 191 se
rect 17401 165 17425 191
tri 17425 165 17451 191 nw
rect 16959 159 17419 165
tri 17419 159 17425 165 nw
rect 18544 159 20799 211
tri 20799 159 20873 233 nw
rect 16959 131 17391 159
tri 17391 131 17419 159 nw
rect 16465 122 16517 128
rect 16465 58 16517 70
rect 16465 0 16517 6
rect 16556 125 16608 131
rect 16958 129 17389 131
tri 17389 129 17391 131 nw
rect 16958 125 17088 129
rect 16958 91 16970 125
rect 17004 91 17042 125
rect 17076 91 17088 125
rect 16958 85 17088 91
tri 18462 85 18504 127 se
rect 18504 85 20497 127
tri 18452 75 18462 85 se
rect 18462 75 20497 85
rect 16556 61 16608 73
tri 18436 59 18452 75 se
rect 18452 73 18524 75
tri 18524 73 18526 75 nw
rect 18452 59 18510 73
tri 18510 59 18524 73 nw
tri 20945 59 20959 73 se
rect 20959 67 21218 73
rect 20959 59 21166 67
tri 18432 55 18436 59 se
rect 18436 55 18506 59
tri 18506 55 18510 59 nw
tri 20941 55 20945 59 se
rect 20945 55 21166 59
rect 16608 9 16754 55
rect 16556 3 16754 9
tri 18380 3 18432 55 se
rect 18432 45 18496 55
tri 18496 45 18506 55 nw
tri 20931 45 20941 55 se
rect 20941 45 21166 55
rect 18432 3 18454 45
tri 18454 3 18496 45 nw
tri 18520 3 18562 45 se
rect 18562 3 19445 45
tri 18377 0 18380 3 se
rect 18380 0 18451 3
tri 18451 0 18454 3 nw
tri 18517 0 18520 3 se
rect 18520 0 19445 3
tri 18362 -15 18377 0 se
rect 18377 -1 18450 0
tri 18450 -1 18451 0 nw
tri 18516 -1 18517 0 se
rect 18517 -1 19445 0
rect 18377 -7 18444 -1
tri 18444 -7 18450 -1 nw
tri 18510 -7 18516 -1 se
rect 18516 -7 19445 -1
rect 19497 -7 19523 45
rect 19575 -7 19581 45
tri 20925 39 20931 45 se
rect 20931 39 21166 45
tri 20915 29 20925 39 se
rect 20925 29 20959 39
tri 20959 29 20969 39 nw
tri 20885 -1 20915 29 se
rect 20915 -1 20929 29
tri 20929 -1 20959 29 nw
rect 21166 3 21218 15
tri 20879 -7 20885 -1 se
rect 20885 -7 20921 -1
rect 18377 -15 18436 -7
tri 18436 -15 18444 -7 nw
tri 18502 -15 18510 -7 se
rect 18510 -15 18562 -7
tri 18358 -19 18362 -15 se
rect 18362 -19 18432 -15
tri 18432 -19 18436 -15 nw
tri 18498 -19 18502 -15 se
rect 18502 -19 18562 -15
tri 17723 -42 17746 -19 se
rect 17746 -42 18209 -19
rect 6460 -139 6472 -105
rect 6506 -139 6551 -105
rect 6585 -139 6597 -105
tri 6096 -251 6134 -213 sw
rect 6029 -255 6134 -251
tri 6134 -255 6138 -251 sw
rect 6029 -256 6138 -255
tri 6138 -256 6139 -255 sw
rect 6029 -272 6310 -256
tri 6310 -272 6326 -256 sw
tri 6444 -272 6460 -256 se
rect 6460 -272 6597 -139
rect 16657 -93 16773 -42
tri 16773 -93 16824 -42 sw
tri 17672 -93 17723 -42 se
rect 17723 -71 18209 -42
tri 18306 -71 18358 -19 se
rect 18358 -57 18394 -19
tri 18394 -57 18432 -19 nw
tri 18460 -57 18498 -19 se
rect 18498 -57 18562 -19
tri 18562 -57 18612 -7 nw
tri 20871 -15 20879 -7 se
rect 20879 -9 20921 -7
tri 20921 -9 20929 -1 nw
tri 20965 -9 20973 -1 se
rect 20973 -9 21009 -1
rect 20879 -15 20915 -9
tri 20915 -15 20921 -9 nw
tri 20959 -15 20965 -9 se
rect 20965 -15 21009 -9
tri 20833 -53 20871 -15 se
rect 20871 -53 20877 -15
tri 20877 -53 20915 -15 nw
tri 20921 -53 20959 -15 se
rect 20959 -53 21009 -15
rect 21061 -53 21073 -1
rect 21125 -53 21131 -1
tri 20831 -55 20833 -53 se
rect 20833 -55 20875 -53
tri 20875 -55 20877 -53 nw
tri 20919 -55 20921 -53 se
rect 20921 -55 20964 -53
tri 20964 -55 20966 -53 nw
rect 21166 -55 21218 -49
tri 20829 -57 20831 -55 se
rect 20831 -57 20873 -55
tri 20873 -57 20875 -55 nw
tri 20917 -57 20919 -55 se
rect 20919 -57 20962 -55
tri 20962 -57 20964 -55 nw
rect 18358 -71 18380 -57
tri 18380 -71 18394 -57 nw
tri 18446 -71 18460 -57 se
rect 18460 -71 18480 -57
rect 17723 -93 17746 -71
tri 17746 -93 17768 -71 nw
tri 18288 -89 18306 -71 se
rect 18306 -81 18370 -71
tri 18370 -81 18380 -71 nw
tri 18436 -81 18446 -71 se
rect 18446 -81 18480 -71
rect 18306 -89 18362 -81
tri 18362 -89 18370 -81 nw
tri 18428 -89 18436 -81 se
rect 18436 -89 18480 -81
tri 18284 -93 18288 -89 se
rect 18288 -93 18358 -89
tri 18358 -93 18362 -89 nw
tri 18424 -93 18428 -89 se
rect 18428 -93 18480 -89
rect 16657 -98 16824 -93
tri 16824 -98 16829 -93 sw
tri 17667 -98 17672 -93 se
rect 17672 -98 17741 -93
tri 17741 -98 17746 -93 nw
tri 18279 -98 18284 -93 se
rect 18284 -98 18353 -93
tri 18353 -98 18358 -93 nw
tri 18419 -98 18424 -93 se
rect 18424 -98 18480 -93
rect 16657 -129 16829 -98
tri 16829 -129 16860 -98 sw
rect 17662 -129 17710 -98
tri 17710 -129 17741 -98 nw
tri 18266 -111 18279 -98 se
rect 18279 -111 18322 -98
rect 17945 -129 18322 -111
tri 18322 -129 18353 -98 nw
tri 18388 -129 18419 -98 se
rect 18419 -129 18480 -98
rect 16657 -150 16860 -129
tri 16860 -150 16881 -129 sw
rect 17662 -150 17689 -129
tri 17689 -150 17710 -129 nw
rect 17945 -150 18301 -129
tri 18301 -150 18322 -129 nw
tri 18367 -150 18388 -129 se
rect 18388 -139 18480 -129
tri 18480 -139 18562 -57 nw
rect 20385 -67 20863 -57
tri 20863 -67 20873 -57 nw
tri 20907 -67 20917 -57 se
rect 20917 -67 20952 -57
tri 20952 -67 20962 -57 nw
rect 20385 -68 20862 -67
tri 20862 -68 20863 -67 nw
tri 20906 -68 20907 -67 se
rect 20907 -68 20928 -67
rect 20385 -91 20839 -68
tri 20839 -91 20862 -68 nw
tri 20883 -91 20906 -68 se
rect 20906 -91 20928 -68
tri 20928 -91 20952 -67 nw
rect 20385 -139 20419 -91
tri 20862 -112 20883 -91 se
rect 20883 -112 20907 -91
tri 20907 -112 20928 -91 nw
tri 20851 -123 20862 -112 se
rect 20862 -123 20896 -112
tri 20896 -123 20907 -112 nw
rect 18388 -142 18477 -139
tri 18477 -142 18480 -139 nw
tri 18520 -142 18523 -139 se
rect 18523 -142 20419 -139
rect 18388 -150 18460 -142
rect 16657 -159 16881 -150
tri 16881 -159 16890 -150 sw
rect 17945 -155 18296 -150
tri 18296 -155 18301 -150 nw
tri 18362 -155 18367 -150 se
rect 18367 -155 18460 -150
rect 17945 -159 18292 -155
tri 18292 -159 18296 -155 nw
tri 18358 -159 18362 -155 se
rect 18362 -159 18460 -155
tri 18460 -159 18477 -142 nw
tri 18503 -159 18520 -142 se
rect 18520 -159 20419 -142
rect 16657 -196 16890 -159
tri 16890 -196 16927 -159 sw
rect 17945 -163 18288 -159
tri 18288 -163 18292 -159 nw
tri 18354 -163 18358 -159 se
rect 18358 -163 18434 -159
tri 18321 -196 18354 -163 se
rect 18354 -185 18434 -163
tri 18434 -185 18460 -159 nw
tri 18489 -173 18503 -159 se
rect 18503 -173 20419 -159
rect 20450 -157 20862 -123
tri 20862 -157 20896 -123 nw
tri 18477 -185 18489 -173 se
rect 18489 -185 18523 -173
tri 18523 -185 18535 -173 nw
rect 18354 -188 18431 -185
tri 18431 -188 18434 -185 nw
tri 18474 -188 18477 -185 se
rect 18477 -188 18506 -185
rect 18354 -196 18423 -188
tri 18423 -196 18431 -188 nw
tri 18466 -196 18474 -188 se
rect 18474 -196 18506 -188
rect 16657 -204 18415 -196
tri 18415 -204 18423 -196 nw
tri 18460 -202 18466 -196 se
rect 18466 -202 18506 -196
tri 18506 -202 18523 -185 nw
rect 20450 -202 20484 -157
tri 18458 -204 18460 -202 se
rect 18460 -204 18477 -202
rect 16657 -231 18388 -204
tri 18388 -231 18415 -204 nw
tri 18431 -231 18458 -204 se
rect 18458 -231 18477 -204
tri 18477 -231 18506 -202 nw
tri 18518 -231 18547 -202 se
rect 18547 -231 20484 -202
rect 16657 -234 18385 -231
tri 18385 -234 18388 -231 nw
tri 18430 -232 18431 -231 se
rect 18431 -232 18476 -231
tri 18476 -232 18477 -231 nw
tri 18517 -232 18518 -231 se
rect 18518 -232 20484 -231
tri 18428 -234 18430 -232 se
rect 18430 -234 18449 -232
rect 16657 -251 18368 -234
tri 18368 -251 18385 -234 nw
tri 18411 -251 18428 -234 se
rect 18428 -251 18449 -234
tri 16661 -255 16665 -251 ne
rect 16665 -255 17318 -251
tri 16665 -256 16666 -255 ne
rect 16666 -256 16717 -255
tri 6597 -272 6613 -256 sw
rect -2987 -305 -2935 -293
rect -1473 -311 -1467 -295
rect -2987 -363 -2935 -357
rect -2885 -317 -1467 -311
rect -2833 -347 -1467 -317
rect -1415 -347 -1403 -295
rect -1351 -347 -1345 -295
tri 6008 -332 6029 -311 se
rect 6029 -332 6613 -272
tri 16666 -275 16685 -256 ne
rect 16685 -275 16717 -256
tri 16685 -289 16699 -275 ne
rect 16699 -289 16717 -275
rect 16751 -289 16797 -255
rect 16831 -289 16877 -255
rect 16911 -289 16956 -255
rect 16990 -289 17035 -255
rect 17069 -289 17114 -255
rect 17148 -289 17193 -255
rect 17227 -289 17272 -255
rect 17306 -289 17318 -255
tri 16699 -290 16700 -289 ne
rect 16700 -290 17318 -289
rect 14804 -295 16634 -290
tri 16634 -295 16639 -290 sw
tri 16700 -295 16705 -290 ne
rect 16705 -295 17318 -290
tri 17318 -295 17362 -251 nw
tri 18385 -277 18411 -251 se
rect 18411 -259 18449 -251
tri 18449 -259 18476 -232 nw
tri 18490 -259 18517 -232 se
rect 18517 -259 18536 -232
tri 18536 -259 18563 -232 nw
rect 18411 -264 18444 -259
tri 18444 -264 18449 -259 nw
tri 18485 -264 18490 -259 se
rect 18490 -264 18518 -259
rect 18411 -277 18431 -264
tri 18431 -277 18444 -264 nw
tri 18472 -277 18485 -264 se
rect 18485 -277 18518 -264
tri 18518 -277 18536 -259 nw
tri 18367 -295 18385 -277 se
rect 18385 -295 18411 -277
rect 14804 -297 16639 -295
tri 16639 -297 16641 -295 sw
tri 18365 -297 18367 -295 se
rect 18367 -297 18411 -295
tri 18411 -297 18431 -277 nw
tri 18452 -297 18472 -277 se
rect 18472 -297 18498 -277
tri 18498 -297 18518 -277 nw
rect 14804 -318 16641 -297
tri 16641 -318 16662 -297 sw
rect 17365 -305 18403 -297
tri 18403 -305 18411 -297 nw
tri 18444 -305 18452 -297 se
rect 18452 -305 18490 -297
tri 18490 -305 18498 -297 nw
rect 17365 -310 18398 -305
tri 18398 -310 18403 -305 nw
tri 18439 -310 18444 -305 se
rect 18444 -310 18477 -305
rect 17365 -318 18390 -310
tri 18390 -318 18398 -310 nw
tri 18431 -318 18439 -310 se
rect 18439 -318 18477 -310
tri 18477 -318 18490 -305 nw
rect 14804 -324 16662 -318
tri 16662 -324 16668 -318 sw
rect 17365 -324 18384 -318
tri 18384 -324 18390 -318 nw
tri 18425 -324 18431 -318 se
rect 18431 -324 18471 -318
tri 18471 -324 18477 -318 nw
rect -2885 -381 -2833 -369
rect 5814 -394 6613 -332
tri 16620 -363 16659 -324 ne
rect 16659 -363 16668 -324
tri 16668 -363 16707 -324 sw
rect 17365 -331 18377 -324
tri 18377 -331 18384 -324 nw
tri 18418 -331 18425 -324 se
rect 18425 -331 18464 -324
tri 18464 -331 18471 -324 nw
rect 14803 -366 16617 -363
tri 16617 -366 16620 -363 sw
tri 16659 -366 16662 -363 ne
rect 16662 -366 16707 -363
tri 16707 -366 16710 -363 sw
rect 17365 -366 17399 -331
tri 18398 -351 18418 -331 se
rect 18418 -351 18444 -331
tri 18444 -351 18464 -331 nw
tri 18386 -363 18398 -351 se
rect 18398 -363 18432 -351
tri 18432 -363 18444 -351 nw
rect 14803 -391 16620 -366
tri 16620 -391 16645 -366 sw
tri 16662 -391 16687 -366 ne
rect 16687 -391 17399 -366
rect 14803 -394 16645 -391
tri 16645 -394 16648 -391 sw
tri 16687 -394 16690 -391 ne
rect 16690 -394 17399 -391
rect 14803 -397 16648 -394
rect -2885 -439 -2833 -433
tri 16603 -439 16645 -397 ne
rect 16645 -400 16648 -397
tri 16648 -400 16654 -394 sw
tri 16690 -400 16696 -394 ne
rect 16696 -400 17399 -394
rect 17430 -397 18398 -363
tri 18398 -397 18432 -363 nw
rect 16645 -439 16654 -400
tri 16654 -439 16693 -400 sw
rect 17430 -439 17464 -397
tri 16645 -473 16679 -439 ne
rect 16679 -473 17464 -439
rect -2602 -3678 -2282 -3594
rect -2602 -3712 -2371 -3678
rect -2337 -3712 -2282 -3678
rect -2602 -3750 -2282 -3712
rect -2602 -3784 -2371 -3750
rect -2337 -3784 -2282 -3750
rect -2602 -3797 -2282 -3784
tri -2565 -4049 -2553 -4037 se
rect -2553 -4049 -2507 -4037
tri -2587 -4071 -2565 -4049 se
rect -2565 -4071 -2547 -4049
rect -2987 -4077 -2547 -4071
rect -2935 -4083 -2547 -4077
rect -2513 -4083 -2507 -4049
rect -2935 -4121 -2507 -4083
rect -2935 -4129 -2547 -4121
rect -2987 -4143 -2547 -4129
rect -2935 -4155 -2547 -4143
rect -2513 -4155 -2507 -4121
rect -2935 -4167 -2507 -4155
rect -2987 -4201 -2935 -4195
tri -2935 -4201 -2901 -4167 nw
rect -2885 -4211 -2410 -4205
rect -2833 -4217 -2410 -4211
rect -2833 -4251 -2450 -4217
rect -2416 -4251 -2410 -4217
rect -2833 -4263 -2410 -4251
rect -2885 -4277 -2410 -4263
rect -2833 -4289 -2410 -4277
rect -2833 -4323 -2450 -4289
rect -2416 -4323 -2410 -4289
rect -2833 -4329 -2410 -4323
rect -2885 -4335 -2410 -4329
rect -2602 -4429 -2283 -4417
rect -2602 -4463 -2371 -4429
rect -2337 -4463 -2283 -4429
rect -2602 -4501 -2283 -4463
rect -2602 -4535 -2371 -4501
rect -2337 -4535 -2283 -4501
rect -2602 -4632 -2283 -4535
rect -2271 -4978 -2141 -4972
rect -2271 -5012 -2259 -4978
rect -2225 -5012 -2187 -4978
rect -2153 -5012 -2141 -4978
rect -2271 -5018 -2141 -5012
rect -2800 -5064 -2748 -5058
rect -2748 -5095 -2227 -5089
rect -2748 -5116 -2345 -5095
rect -2800 -5129 -2345 -5116
rect -2311 -5129 -2273 -5095
rect -2239 -5129 -2227 -5095
rect -2800 -5130 -2227 -5129
rect -2748 -5135 -2227 -5130
rect -2800 -5188 -2748 -5182
rect -2716 -5179 -2368 -5173
rect -2664 -5185 -2368 -5179
rect -2664 -5219 -2409 -5185
rect -2375 -5219 -2368 -5185
rect -2664 -5231 -2368 -5219
rect -2716 -5240 -2368 -5231
rect -2716 -5243 -2664 -5240
rect -2716 -5301 -2664 -5295
rect -2415 -5257 -2369 -5240
rect -2415 -5291 -2409 -5257
rect -2375 -5291 -2369 -5257
rect -2198 -5265 -2144 -5018
rect -2415 -5303 -2369 -5291
rect -2274 -5271 -2144 -5265
rect -2274 -5305 -2262 -5271
rect -2228 -5305 -2190 -5271
rect -2156 -5305 -2144 -5271
rect -2274 -5311 -2144 -5305
rect -2800 -5353 -2331 -5347
rect -2748 -5393 -2331 -5353
rect -2800 -5419 -2748 -5405
rect -2800 -5477 -2748 -5471
rect -2387 -5441 -2331 -5393
rect -2387 -5447 -2183 -5441
rect -2387 -5481 -2301 -5447
rect -2267 -5481 -2229 -5447
rect -2195 -5481 -2183 -5447
rect -2387 -5487 -2183 -5481
rect -3072 -5869 -3020 -5863
rect -3174 -5930 -3122 -5924
rect -3174 -5994 -3122 -5982
rect -3072 -5933 -3020 -5921
rect -3020 -5985 -1416 -5959
rect -3072 -5991 -1416 -5985
rect -1422 -6011 -1416 -5991
rect -1364 -6011 -1352 -5959
rect -1300 -6011 -1294 -5959
rect -3122 -6026 -1638 -6020
rect -3122 -6046 -1690 -6026
rect -3174 -6052 -1690 -6046
rect -1690 -6090 -1638 -6078
rect -2716 -6100 -1946 -6094
rect -2664 -6152 -1998 -6100
rect -1690 -6148 -1638 -6142
rect -2716 -6161 -1946 -6152
rect -2716 -6164 -2664 -6161
rect -2716 -6222 -2664 -6216
rect -1998 -6164 -1946 -6161
rect -1998 -6222 -1946 -6216
rect -2885 -6263 -2833 -6257
rect -2987 -6330 -2935 -6324
rect -2987 -6394 -2935 -6382
rect -2885 -6327 -2833 -6315
rect -2833 -6379 -1918 -6349
rect -2885 -6385 -1918 -6379
tri -1940 -6401 -1924 -6385 ne
rect -1924 -6401 -1918 -6385
rect -1866 -6401 -1854 -6349
rect -1802 -6401 -1796 -6349
rect -2935 -6446 -2098 -6416
rect -2987 -6452 -2098 -6446
tri -2120 -6468 -2104 -6452 ne
rect -2104 -6468 -2098 -6452
rect -2046 -6468 -2034 -6416
rect -1982 -6468 -1976 -6416
rect -2800 -6639 -2748 -6633
rect -2800 -6705 -2748 -6691
rect -3051 -6772 -2852 -6748
rect -3051 -6824 -2904 -6772
rect -3051 -6838 -2852 -6824
rect -3051 -6890 -2904 -6838
rect -3051 -7079 -2852 -6890
rect -2800 -6778 -2748 -6757
rect -2716 -6639 -2664 -6633
rect -2716 -6705 -2664 -6691
tri -2664 -6737 -2626 -6699 sw
rect -2664 -6757 -2626 -6737
rect -2716 -6763 -2626 -6757
tri -2626 -6763 -2600 -6737 sw
tri -2698 -6766 -2695 -6763 ne
rect -2695 -6766 -2600 -6763
rect -1633 -6743 -1581 -6737
tri -2695 -6772 -2689 -6766 ne
rect -2689 -6772 -2600 -6766
tri -2748 -6778 -2742 -6772 sw
tri -2689 -6778 -2683 -6772 ne
rect -2683 -6778 -2600 -6772
rect -2800 -6809 -2742 -6778
tri -2742 -6809 -2711 -6778 sw
tri -2683 -6809 -2652 -6778 ne
rect -2800 -6812 -2711 -6809
tri -2711 -6812 -2708 -6809 sw
rect -2800 -6830 -2708 -6812
tri -2708 -6830 -2690 -6812 sw
rect -2800 -6842 -2690 -6830
rect -2800 -6876 -2730 -6842
rect -2696 -6876 -2690 -6842
rect -2800 -6914 -2690 -6876
rect -2800 -6948 -2730 -6914
rect -2696 -6948 -2690 -6914
rect -2800 -6960 -2690 -6948
tri -2679 -7002 -2652 -6975 se
rect -2652 -7002 -2600 -6778
rect -2535 -6772 -2483 -6766
rect -2377 -6768 -2331 -6766
rect -2535 -6838 -2483 -6824
rect -2535 -6896 -2483 -6890
rect -2383 -6774 -2331 -6768
tri -2331 -6778 -2319 -6766 sw
tri -1833 -6778 -1821 -6766 se
rect -1821 -6778 -1633 -6766
rect -2331 -6797 -2319 -6778
tri -2319 -6797 -2300 -6778 sw
tri -1852 -6797 -1833 -6778 se
rect -1833 -6797 -1815 -6778
rect -2331 -6812 -1815 -6797
rect -1781 -6795 -1633 -6778
tri -1581 -6766 -1552 -6737 sw
rect -1581 -6778 -1463 -6766
rect -1581 -6795 -1503 -6778
rect -1781 -6807 -1503 -6795
rect -1781 -6812 -1633 -6807
rect -2331 -6826 -1633 -6812
rect -2383 -6838 -1633 -6826
rect -2331 -6850 -1633 -6838
rect -2331 -6852 -1815 -6850
tri -2331 -6882 -2301 -6852 nw
tri -1852 -6882 -1822 -6852 ne
rect -1822 -6882 -1815 -6852
tri -1822 -6883 -1821 -6882 ne
rect -2383 -6896 -2331 -6890
rect -1821 -6884 -1815 -6882
rect -1781 -6859 -1633 -6850
rect -1581 -6812 -1503 -6807
rect -1469 -6812 -1463 -6778
rect -1581 -6850 -1463 -6812
rect -1581 -6859 -1503 -6850
rect -1781 -6865 -1503 -6859
rect -1781 -6884 -1763 -6865
tri -1763 -6884 -1744 -6865 nw
rect -1509 -6884 -1503 -6865
rect -1469 -6884 -1463 -6850
rect -1821 -6896 -1775 -6884
tri -1775 -6896 -1763 -6884 nw
rect -1509 -6896 -1463 -6884
tri -996 -6919 -977 -6900 se
rect -2138 -6925 -2086 -6919
tri -2600 -7002 -2573 -6975 sw
tri -1003 -6926 -996 -6919 se
rect -996 -6926 -977 -6919
rect -1703 -6932 -977 -6926
rect -1703 -6966 -1691 -6932
rect -1657 -6966 -1619 -6932
rect -1585 -6966 -977 -6932
rect -1703 -6972 -977 -6966
rect -2138 -6989 -2086 -6977
rect -2699 -7008 -2569 -7002
rect -2699 -7042 -2687 -7008
rect -2653 -7042 -2615 -7008
rect -2581 -7042 -2569 -7008
rect -2699 -7048 -2569 -7042
rect -2482 -7008 -2138 -7002
rect -2482 -7042 -2470 -7008
rect -2436 -7042 -2398 -7008
rect -2364 -7041 -2138 -7008
tri -1279 -6994 -1257 -6972 ne
rect -2086 -7041 -1739 -7002
rect -2364 -7042 -1739 -7041
rect -2482 -7048 -1739 -7042
rect -1801 -7050 -1739 -7048
rect -1801 -7056 -1513 -7050
rect -1801 -7090 -1758 -7056
rect -1724 -7090 -1659 -7056
rect -1625 -7090 -1559 -7056
rect -1525 -7090 -1513 -7056
rect -1801 -7096 -1513 -7090
rect -1429 -7141 -1377 -7093
rect -1257 -7097 -977 -6972
rect -2086 -7187 -1377 -7141
<< via1 >>
rect -3122 1733 -3070 1785
rect -3058 1733 -3006 1785
rect -1262 1733 -1210 1785
rect -1198 1733 -1146 1785
rect -971 1771 -919 1823
rect -971 1707 -919 1759
rect -3072 1548 -3020 1600
rect -1262 1554 -1210 1606
rect -1198 1554 -1146 1606
rect -3072 1484 -3020 1536
rect 21554 1528 21606 1550
rect 21554 1498 21558 1528
rect 21558 1498 21592 1528
rect 21592 1498 21606 1528
rect 21618 1528 21670 1550
rect 21618 1498 21630 1528
rect 21630 1498 21664 1528
rect 21664 1498 21670 1528
rect 20969 1398 21021 1450
rect 19188 1321 19240 1373
rect 19252 1321 19304 1373
rect 20969 1334 21021 1386
rect 21322 1398 21374 1450
rect 21322 1334 21374 1386
rect 21658 1375 21664 1408
rect 21664 1375 21698 1408
rect 21698 1375 21710 1408
rect 21658 1356 21710 1375
rect 21658 1337 21710 1342
rect 21658 1303 21664 1337
rect 21664 1303 21698 1337
rect 21698 1303 21710 1337
rect 21658 1290 21710 1303
rect 19676 1259 19728 1270
rect 19740 1259 19792 1270
rect 19676 1225 19678 1259
rect 19678 1225 19726 1259
rect 19726 1225 19728 1259
rect 19740 1225 19760 1259
rect 19760 1225 19792 1259
rect 19676 1218 19728 1225
rect 19740 1218 19792 1225
rect 21387 902 21439 954
rect 21451 902 21503 954
rect 18630 673 18682 725
rect 18694 673 18746 725
rect 18960 673 19012 725
rect 19024 673 19076 725
rect 21431 665 21483 717
rect 21495 665 21547 717
rect 96 598 148 650
rect 96 534 148 586
rect 19092 574 19144 626
rect 19156 574 19208 626
rect 14 470 20 490
rect 20 470 54 490
rect 54 470 66 490
rect 14 438 66 470
rect 14 415 66 426
rect 14 381 20 415
rect 20 381 54 415
rect 54 381 66 415
rect 14 374 66 381
rect -54 23 -2 75
rect -2800 -67 -2748 -15
rect -1251 -46 -1199 6
rect -1187 -46 -1135 6
rect -54 -41 -2 11
rect 32 -59 84 -7
rect -2800 -131 -2748 -79
rect -2716 -134 -2664 -82
rect -1251 -128 -1199 -76
rect -1187 -128 -1135 -76
rect 32 -123 84 -71
rect -2716 -198 -2664 -146
rect -2987 -293 -2935 -241
rect -1251 -283 -1199 -231
rect -1187 -283 -1135 -231
rect 18092 341 18144 393
rect 18156 341 18208 393
rect 18089 255 18141 307
rect 18154 255 18206 307
rect 16465 70 16517 122
rect 16465 6 16517 58
rect 16556 73 16608 125
rect 16556 9 16608 61
rect 19445 -7 19497 45
rect 19523 -7 19575 45
rect 21166 15 21218 67
rect 21009 -53 21061 -1
rect 21073 -53 21125 -1
rect 21166 -49 21218 3
rect -2987 -357 -2935 -305
rect -2885 -369 -2833 -317
rect -1467 -347 -1415 -295
rect -1403 -347 -1351 -295
rect -2885 -433 -2833 -381
rect -2987 -4129 -2935 -4077
rect -2987 -4195 -2935 -4143
rect -2885 -4263 -2833 -4211
rect -2885 -4329 -2833 -4277
rect -2800 -5116 -2748 -5064
rect -2800 -5182 -2748 -5130
rect -2716 -5231 -2664 -5179
rect -2716 -5295 -2664 -5243
rect -2800 -5405 -2748 -5353
rect -2800 -5471 -2748 -5419
rect -3072 -5921 -3020 -5869
rect -3174 -5982 -3122 -5930
rect -3072 -5985 -3020 -5933
rect -3174 -6046 -3122 -5994
rect -1416 -6011 -1364 -5959
rect -1352 -6011 -1300 -5959
rect -1690 -6078 -1638 -6026
rect -2716 -6152 -2664 -6100
rect -1998 -6152 -1946 -6100
rect -1690 -6142 -1638 -6090
rect -2716 -6216 -2664 -6164
rect -1998 -6216 -1946 -6164
rect -2885 -6315 -2833 -6263
rect -2987 -6382 -2935 -6330
rect -2885 -6379 -2833 -6327
rect -2987 -6446 -2935 -6394
rect -1918 -6401 -1866 -6349
rect -1854 -6401 -1802 -6349
rect -2098 -6468 -2046 -6416
rect -2034 -6468 -1982 -6416
rect -2800 -6691 -2748 -6639
rect -2904 -6824 -2852 -6772
rect -2904 -6890 -2852 -6838
rect -2800 -6757 -2748 -6705
rect -2716 -6691 -2664 -6639
rect -2716 -6757 -2664 -6705
rect -2535 -6778 -2483 -6772
rect -2535 -6812 -2527 -6778
rect -2527 -6812 -2493 -6778
rect -2493 -6812 -2483 -6778
rect -2535 -6824 -2483 -6812
rect -2535 -6850 -2483 -6838
rect -2535 -6884 -2527 -6850
rect -2527 -6884 -2493 -6850
rect -2493 -6884 -2483 -6850
rect -2535 -6890 -2483 -6884
rect -2383 -6778 -2331 -6774
rect -2383 -6812 -2371 -6778
rect -2371 -6812 -2337 -6778
rect -2337 -6812 -2331 -6778
rect -1633 -6795 -1581 -6743
rect -2383 -6826 -2331 -6812
rect -2383 -6850 -2331 -6838
rect -2383 -6884 -2371 -6850
rect -2371 -6884 -2337 -6850
rect -2337 -6884 -2331 -6850
rect -2383 -6890 -2331 -6884
rect -1633 -6859 -1581 -6807
rect -2138 -6977 -2086 -6925
rect -2138 -7041 -2086 -6989
<< metal2 >>
rect -971 1823 -919 1829
rect -3174 1733 -3122 1785
rect -3070 1733 -3058 1785
rect -3006 1733 -3000 1785
rect -1268 1733 -1262 1785
rect -1210 1733 -1198 1785
rect -1146 1771 -971 1785
rect -1146 1759 -919 1771
rect -1146 1733 -971 1759
rect -3174 1707 -3101 1733
tri -3101 1707 -3075 1733 nw
rect -3174 -5930 -3122 1707
tri -3122 1686 -3101 1707 nw
rect -971 1701 -919 1707
rect -3174 -5994 -3122 -5982
rect -3072 1600 -3020 1606
rect -1268 1554 -1262 1606
rect -1210 1554 -1198 1606
rect -1146 1554 -1140 1606
rect -3072 1536 -3020 1548
rect -3072 -5869 -3020 1484
rect 20969 1450 21022 2827
rect 21021 1398 21022 1450
rect 20969 1386 21022 1398
rect 19182 1321 19188 1373
rect 19240 1321 19252 1373
rect 19304 1321 19310 1373
rect 21021 1334 21022 1386
rect 19670 1218 19676 1270
rect 19728 1218 19740 1270
rect 19792 1218 19798 1270
rect 19108 774 19141 798
rect 18624 673 18630 725
rect 18682 673 18694 725
rect 18746 673 18752 725
rect 18951 673 18960 725
rect 19012 673 19024 725
rect 19076 673 19082 725
rect 96 650 148 656
rect 96 586 148 598
rect -1001 534 96 564
rect -1001 528 148 534
rect -1001 160 -965 528
rect 14 490 66 496
rect 14 426 66 438
rect -1393 124 -965 160
rect -936 374 14 404
rect 18625 396 18701 673
rect -936 368 66 374
rect 18086 393 18701 396
rect -2800 -15 -2748 -9
rect -2800 -79 -2748 -67
rect -3072 -5933 -3020 -5921
rect -3072 -5991 -3020 -5985
rect -2987 -241 -2935 -235
rect -2987 -305 -2935 -293
rect -2987 -4077 -2935 -357
rect -2987 -4143 -2935 -4129
rect -3174 -6052 -3122 -6046
rect -2987 -6330 -2935 -4195
rect -2987 -6394 -2935 -6382
rect -2885 -317 -2833 -311
rect -2885 -381 -2833 -369
rect -2885 -4211 -2833 -433
rect -2885 -4277 -2833 -4263
rect -2885 -6263 -2833 -4329
rect -2885 -6327 -2833 -6315
rect -2885 -6385 -2833 -6379
rect -2800 -5064 -2748 -131
rect -2800 -5130 -2748 -5116
rect -2800 -5353 -2748 -5182
rect -2800 -5419 -2748 -5405
rect -2987 -6452 -2935 -6446
rect -2800 -6639 -2748 -5471
rect -2800 -6705 -2748 -6691
rect -2800 -6763 -2748 -6757
rect -2716 -82 -2664 -76
rect -2716 -146 -2664 -134
rect -2716 -5179 -2664 -198
rect -1393 -295 -1357 124
rect -936 92 -900 368
rect 18086 341 18092 393
rect 18144 341 18156 393
rect 18208 341 18701 393
rect 18086 339 18701 341
rect 18951 307 19048 673
rect 19086 574 19092 626
rect 19144 574 19156 626
rect 19208 574 19214 626
rect 19723 311 19775 1218
rect 18083 255 18089 307
rect 18141 255 18154 307
rect 18206 255 19048 307
rect 18083 254 19048 255
rect 19529 259 19775 311
rect -1327 56 -900 92
rect 16465 122 16517 128
rect -54 75 -2 81
rect -1327 -231 -1291 56
rect -54 11 -2 23
rect -1257 -46 -1251 6
rect -1199 -46 -1187 6
rect -1135 -41 -54 6
rect 16465 58 16517 70
rect 16465 0 16517 6
rect 16556 125 16608 131
rect 16556 61 16608 73
rect 19529 45 19581 259
rect 20969 98 21022 1334
rect 21322 1450 21375 2956
rect 21548 1498 21554 1550
rect 21606 1498 21618 1550
rect 21670 1498 21676 1550
rect 21374 1398 21375 1450
tri 21624 1408 21630 1414 se
rect 21630 1408 21710 1414
rect 21322 1386 21375 1398
rect 21374 1334 21375 1386
tri 21572 1356 21624 1408 se
rect 21624 1356 21658 1408
tri 21558 1342 21572 1356 se
rect 21572 1342 21710 1356
tri 21248 1090 21322 1164 se
rect 21322 1143 21375 1334
tri 21322 1090 21375 1143 nw
tri 21529 1313 21558 1342 se
rect 21558 1313 21658 1342
rect 21529 1290 21658 1313
rect 21529 1284 21710 1290
tri 21503 1090 21529 1116 se
rect 21529 1098 21569 1284
tri 21569 1264 21589 1284 nw
tri 21174 1016 21248 1090 se
tri 21248 1016 21322 1090 nw
tri 21471 1058 21503 1090 se
rect 21503 1058 21529 1090
tri 21529 1058 21569 1098 nw
tri 21467 1054 21471 1058 se
rect 21471 1054 21525 1058
tri 21525 1054 21529 1058 nw
tri 21112 954 21174 1016 se
rect 21174 954 21186 1016
tri 21186 954 21248 1016 nw
rect 21467 954 21508 1054
tri 21508 1037 21525 1054 nw
tri 21100 942 21112 954 se
rect 21112 942 21174 954
tri 21174 942 21186 954 nw
tri 21074 916 21100 942 se
rect 21100 916 21148 942
tri 21148 916 21174 942 nw
rect 21074 902 21134 916
tri 21134 902 21148 916 nw
rect 21381 902 21387 954
rect 21439 902 21451 954
rect 21503 902 21509 954
rect 21074 239 21127 902
tri 21127 895 21134 902 nw
rect 21425 665 21431 717
rect 21483 665 21495 717
rect 21547 665 21553 717
tri 21127 239 21148 260 sw
tri 21074 165 21148 239 ne
tri 21148 169 21218 239 sw
rect 21148 165 21218 169
tri 21148 147 21166 165 ne
tri 20969 86 20981 98 ne
rect 20981 86 21022 98
tri 21022 86 21055 119 sw
tri 20981 67 21000 86 ne
rect 21000 67 21055 86
tri 21000 64 21003 67 ne
rect -1135 -46 -2 -41
rect -1131 -47 -2 -46
rect 32 -7 84 -1
rect 32 -71 84 -59
rect -1257 -128 -1251 -76
rect -1199 -128 -1187 -76
rect -1135 -123 32 -76
rect -1135 -128 84 -123
rect -1131 -129 84 -128
rect -1327 -267 -1251 -231
rect -1257 -283 -1251 -267
rect -1199 -283 -1187 -231
rect -1135 -247 -1129 -231
rect -1135 -283 -5 -247
tri -5 -283 31 -247 sw
tri -31 -286 -28 -283 ne
rect -28 -286 31 -283
tri 31 -286 34 -283 sw
tri -28 -295 -19 -286 ne
rect -19 -295 34 -286
rect -1473 -347 -1467 -295
rect -1415 -347 -1403 -295
rect -1351 -311 -1345 -295
tri -19 -309 -5 -295 ne
rect -5 -309 34 -295
tri -5 -311 -3 -309 ne
rect -3 -311 34 -309
rect -1351 -347 -66 -311
tri -66 -347 -30 -311 sw
tri -3 -347 33 -311 ne
rect 33 -338 34 -311
tri 34 -338 86 -286 sw
rect 16465 -338 16500 0
rect 33 -347 86 -338
tri -92 -351 -88 -347 ne
rect -88 -348 -30 -347
tri -30 -348 -29 -347 sw
tri 33 -348 34 -347 ne
rect 34 -348 86 -347
tri 86 -348 96 -338 sw
tri 8837 -348 8847 -338 se
rect 8847 -348 16500 -338
rect -88 -351 -29 -348
tri -29 -351 -26 -348 sw
tri 34 -351 37 -348 ne
rect 37 -351 96 -348
tri -88 -373 -66 -351 ne
rect -66 -373 -26 -351
tri -66 -381 -58 -373 ne
rect -58 -381 -26 -373
tri -26 -381 4 -351 sw
tri 37 -381 67 -351 ne
rect 67 -381 96 -351
rect -2716 -5243 -2664 -5231
rect -2716 -6100 -2664 -5295
rect -2716 -6164 -2664 -6152
rect -2716 -6639 -2664 -6216
rect -2632 -6539 -2580 -381
tri -58 -413 -26 -381 ne
rect -26 -410 4 -381
tri 4 -410 33 -381 sw
tri 67 -410 96 -381 ne
tri 96 -401 149 -348 sw
tri 8784 -401 8837 -348 se
rect 8837 -373 16500 -348
rect 16556 -7 16608 9
rect 19439 -7 19445 45
rect 19497 -7 19523 45
rect 19575 -7 19581 45
rect 21003 -1 21055 67
rect 21166 67 21218 165
rect 21166 3 21218 15
rect 8837 -401 8847 -373
tri 8847 -401 8875 -373 nw
rect 96 -410 149 -401
tri 149 -410 158 -401 sw
tri 8775 -410 8784 -401 se
rect 8784 -410 8838 -401
tri 8838 -410 8847 -401 nw
rect 16556 -403 16591 -7
tri 16591 -24 16608 -7 nw
rect 21003 -53 21009 -1
rect 21061 -53 21073 -1
rect 21125 -53 21131 -1
rect 21166 -55 21218 -49
tri 8907 -410 8914 -403 se
rect 8914 -410 16591 -403
rect -26 -413 33 -410
tri 33 -413 36 -410 sw
tri 96 -413 99 -410 ne
rect 99 -413 3820 -410
tri -26 -475 36 -413 ne
tri 36 -446 69 -413 sw
tri 99 -446 132 -413 ne
rect 132 -446 3820 -413
rect 4023 -446 8802 -410
tri 8802 -446 8838 -410 nw
tri 8871 -446 8907 -410 se
rect 8907 -438 16591 -410
rect 8907 -446 8914 -438
rect 36 -466 69 -446
tri 69 -466 89 -446 sw
tri 8851 -466 8871 -446 se
rect 8871 -466 8914 -446
tri 8914 -466 8942 -438 nw
rect 36 -475 89 -466
tri 89 -475 98 -466 sw
tri 8842 -475 8851 -466 se
rect 8851 -475 8905 -466
tri 8905 -475 8914 -466 nw
tri 36 -492 53 -475 ne
rect 53 -492 3833 -475
tri 3833 -492 3850 -475 sw
tri 4077 -492 4094 -475 se
rect 4094 -492 8888 -475
tri 8888 -492 8905 -475 nw
tri 53 -511 72 -492 ne
rect 72 -511 8869 -492
tri 8869 -511 8888 -492 nw
tri 3803 -528 3820 -511 ne
rect 3820 -528 4090 -511
tri 4090 -528 4107 -511 nw
rect -1422 -6011 -1416 -5959
rect -1364 -6011 -1352 -5959
rect -1300 -6011 -1294 -5959
rect -1690 -6026 -1638 -6020
rect -1690 -6090 -1638 -6078
rect -1998 -6100 -1946 -6094
rect -1998 -6164 -1946 -6152
rect -1998 -6222 -1946 -6216
tri -1741 -6276 -1690 -6225 se
rect -1690 -6256 -1638 -6142
rect -1690 -6276 -1658 -6256
tri -1658 -6276 -1638 -6256 nw
rect -1924 -6401 -1918 -6349
rect -1866 -6401 -1854 -6349
rect -1802 -6401 -1796 -6349
rect -2104 -6468 -2098 -6416
rect -2046 -6468 -2034 -6416
rect -1982 -6468 -1976 -6416
tri -2632 -6544 -2627 -6539 ne
rect -2627 -6544 -2580 -6539
tri -2580 -6544 -2553 -6517 sw
tri -2627 -6591 -2580 -6544 ne
rect -2580 -6591 -2553 -6544
tri -2580 -6618 -2553 -6591 ne
tri -2553 -6618 -2479 -6544 sw
rect -2716 -6705 -2664 -6691
tri -2553 -6692 -2479 -6618 ne
tri -2479 -6645 -2452 -6618 sw
rect -2028 -6645 -1976 -6468
rect -1924 -6645 -1872 -6401
rect -1741 -6641 -1689 -6276
tri -1689 -6307 -1658 -6276 nw
rect -2479 -6649 -2452 -6645
tri -2452 -6649 -2448 -6645 sw
rect -1346 -6649 -1294 -6011
rect -2479 -6692 -2448 -6649
tri -2448 -6692 -2405 -6649 sw
tri -2479 -6743 -2428 -6692 ne
rect -2428 -6737 -2405 -6692
tri -2405 -6737 -2360 -6692 sw
rect -2428 -6743 -2360 -6737
tri -2360 -6743 -2354 -6737 sw
rect -1633 -6743 -1581 -6737
rect -2716 -6763 -2664 -6757
tri -2428 -6763 -2408 -6743 ne
rect -2408 -6763 -2354 -6743
tri -2354 -6763 -2334 -6743 sw
tri -2408 -6766 -2405 -6763 ne
rect -2405 -6766 -2334 -6763
tri -2334 -6766 -2331 -6763 sw
rect -2904 -6772 -2852 -6766
tri -2852 -6772 -2846 -6766 sw
tri -2539 -6772 -2535 -6768 se
rect -2535 -6772 -2483 -6766
rect -2852 -6797 -2846 -6772
tri -2846 -6797 -2821 -6772 sw
tri -2564 -6797 -2539 -6772 se
rect -2539 -6797 -2535 -6772
rect -2852 -6824 -2535 -6797
tri -2405 -6774 -2397 -6766 ne
rect -2397 -6774 -2331 -6766
tri -2397 -6788 -2383 -6774 ne
rect -2904 -6838 -2483 -6824
rect -2852 -6852 -2535 -6838
tri -2852 -6882 -2822 -6852 nw
tri -2564 -6881 -2535 -6852 ne
rect -2904 -6896 -2852 -6890
rect -2535 -6896 -2483 -6890
rect -2383 -6838 -2331 -6826
rect -1633 -6807 -1581 -6795
rect -1633 -6865 -1581 -6859
rect -2383 -6896 -2331 -6890
rect -2138 -6925 -2086 -6919
rect -2138 -6989 -2086 -6977
rect -2138 -7047 -2086 -7041
use sky130_fd_io__ctlv2_ls_analogen_ovtv2  sky130_fd_io__ctlv2_ls_analogen_ovtv2_0
timestamp 1701704242
transform 1 0 -3270 0 1 -8769
box 0 0 2456 2385
use sky130_fd_io__gpio_ovtv2_amux_ctl_ls_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_ctl_ls_i2c_fix_0
timestamp 1701704242
transform 1 0 18358 0 1 219
box -2220 -287 2336 1486
use sky130_fd_io__gpio_ovtv2_amux_ctl_lshv2hv  sky130_fd_io__gpio_ovtv2_amux_ctl_lshv2hv_0
timestamp 1701704242
transform 1 0 4 0 1 0
box -126 -376 7172 1761
use sky130_fd_io__gpio_ovtv2_amux_guardring  sky130_fd_io__gpio_ovtv2_amux_guardring_0
timestamp 1701704242
transform 1 0 -1063 0 1 -236
box -120 -120 4512 3350
use sky130_fd_io__gpiov2_amux_ctl_inv_1_i2c_fix  sky130_fd_io__gpiov2_amux_ctl_inv_1_i2c_fix_0
timestamp 1701704242
transform 1 0 16984 0 -1 391
box 0 0 1 1
use sky130_fd_io__gpiov2_amux_ctl_inv_1_i2c_fix  sky130_fd_io__gpiov2_amux_ctl_inv_1_i2c_fix_1
timestamp 1701704242
transform 1 0 16675 0 -1 391
box 0 0 1 1
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1701704242
transform -1 0 -2263 0 1 -4656
box 107 226 240 873
use sky130_fd_pr__nfet_01v8__example_55959141808472  sky130_fd_pr__nfet_01v8__example_55959141808472_0
timestamp 1701704242
transform 1 0 21728 0 1 1288
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808473  sky130_fd_pr__nfet_01v8__example_55959141808473_0
timestamp 1701704242
transform 1 0 -2685 0 1 -6960
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808474  sky130_fd_pr__nfet_01v8__example_55959141808474_0
timestamp 1701704242
transform -1 0 -2382 0 -1 -6760
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808469  sky130_fd_pr__pfet_01v8__example_55959141808469_0
timestamp 1701704242
transform 1 0 21552 0 1 1599
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808470  sky130_fd_pr__pfet_01v8__example_55959141808470_0
timestamp 1701704242
transform 0 -1 -2127 1 0 -5436
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808471  sky130_fd_pr__pfet_01v8__example_55959141808471_0
timestamp 1701704242
transform 1 0 -1770 0 1 -7008
box -1 0 257 1
<< labels >>
flabel metal2 s 19108 774 19141 798 3 FreeSans 400 0 0 0 HLD_I_H_N
port 0 nsew
flabel locali s 16734 94 16776 122 3 FreeSans 400 0 0 0 ANALOG_EN
port 1 nsew
flabel metal1 s -2200 -7047 -2175 -7004 3 FreeSans 400 90 0 0 ENABLE_VDDA_H
port 2 nsew
flabel metal1 s -2705 -6166 -2681 -6126 3 FreeSans 400 90 0 0 ENABLE_VSWITCH_H
port 3 nsew
flabel metal1 s 17465 -251 17506 -196 3 FreeSans 400 0 0 0 VCCD
port 4 nsew
flabel metal1 s -1196 -6992 -1156 -6965 3 FreeSans 400 0 0 0 VDDA
port 5 nsew
flabel metal1 s 18588 1622 18630 1649 3 FreeSans 400 0 0 0 VDDIO_Q
port 6 nsew
flabel metal1 s -92 1500 -48 1530 3 FreeSans 400 0 0 0 VSSA
port 7 nsew
flabel metal1 s -2192 -5005 -2151 -4974 3 FreeSans 400 0 0 0 VSWITCH
port 8 nsew
flabel metal1 s -1676 -6130 -1647 -6089 3 FreeSans 400 90 0 0 AMUX_EN_VDDA_H
port 9 nsew
flabel metal1 s -1337 -6007 -1307 -5968 3 FreeSans 400 90 0 0 AMUX_EN_VDDA_H_N
port 10 nsew
flabel metal1 s 18573 171 18618 202 3 FreeSans 400 0 0 0 AMUX_EN_VDDIO_H
port 11 nsew
flabel metal1 s 20309 78 20365 125 3 FreeSans 400 0 0 0 AMUX_EN_VDDIO_H_N
port 12 nsew
flabel metal1 s 747 -106 798 -49 3 FreeSans 400 90 0 0 AMUX_EN_VSWITCH_H
port 13 nsew
flabel metal1 s 382 -100 420 -47 3 FreeSans 400 90 0 0 AMUX_EN_VSWITCH_H_N
port 14 nsew
flabel metal1 s 6012 428 6053 459 3 FreeSans 400 0 0 0 VSWITCH
port 8 nsew
flabel metal1 s -2986 -6971 -2942 -6941 3 FreeSans 400 0 0 0 VSSA
port 7 nsew
flabel comment s -1203 -99 -1203 -99 0 FreeSans 280 0 0 0 HLD_H
flabel comment s -1199 -24 -1199 -24 0 FreeSans 280 0 0 0 RST_H
flabel comment s -1419 -318 -1419 -318 0 FreeSans 280 0 0 0 HLD_H
flabel comment s -1199 -261 -1199 -261 0 FreeSans 280 0 0 0 RST_H
flabel comment s 25 576 25 576 0 FreeSans 280 90 0 0 IN_B
flabel comment s 32 984 32 984 0 FreeSans 280 90 0 0 IN
flabel comment s 17783 -39 17783 -39 0 FreeSans 280 0 0 0 AMUX_EN_VDDIO_H
<< properties >>
string FIXED_BBOX 16674 -275 17292 391
string GDS_END 64839508
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 64797130
<< end >>
