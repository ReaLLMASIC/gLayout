magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< dnwell >>
rect -2476 -1400 2776 7401
<< nwell >>
rect -10 0 310 6000
<< pwell >>
rect -3084 7875 3384 8009
rect -3084 -1874 -2950 7875
rect -1102 -26 -374 6026
rect 674 -26 1402 6026
rect 3250 -1874 3384 7875
rect -3084 -2008 3384 -1874
<< mvnmos >>
rect -700 0 -530 6000
rect 830 0 1000 6000
<< mvnnmos >>
rect -530 0 -400 6000
rect 700 0 830 6000
<< mvndiff >>
rect -826 5975 -700 6000
rect -826 25 -814 5975
rect -712 25 -700 5975
rect -826 0 -700 25
rect 1000 5975 1126 6000
rect 1000 25 1012 5975
rect 1114 25 1126 5975
rect 1000 0 1126 25
<< mvndiffc >>
rect -814 25 -712 5975
rect 1012 25 1114 5975
<< mvpsubdiff >>
rect -3058 7959 3358 7983
rect -3058 7925 -2927 7959
rect -2893 7925 -2859 7959
rect -2825 7925 -2791 7959
rect -2757 7925 -2723 7959
rect -2689 7925 -2655 7959
rect -2621 7925 -2587 7959
rect -2553 7925 -2519 7959
rect -2485 7925 -2451 7959
rect -2417 7925 -2383 7959
rect -2349 7925 -2315 7959
rect -2281 7925 -2247 7959
rect -2213 7925 -2179 7959
rect -2145 7925 -2111 7959
rect -2077 7925 -2043 7959
rect -2009 7925 -1975 7959
rect -1941 7925 -1907 7959
rect -1873 7925 -1839 7959
rect -1805 7925 -1771 7959
rect -1737 7925 -1703 7959
rect -1669 7925 -1635 7959
rect -1601 7925 -1567 7959
rect -1533 7925 -1499 7959
rect -1465 7925 -1431 7959
rect -1397 7925 -1363 7959
rect -1329 7925 -1295 7959
rect -1261 7925 -1227 7959
rect -1193 7925 -1159 7959
rect -1125 7925 -1091 7959
rect -1057 7925 -1023 7959
rect -989 7925 -955 7959
rect -921 7925 -887 7959
rect -853 7925 -819 7959
rect -785 7925 -751 7959
rect -717 7925 -683 7959
rect -649 7925 -615 7959
rect -581 7925 -547 7959
rect -513 7925 -479 7959
rect -445 7925 -411 7959
rect -377 7925 -343 7959
rect -309 7925 -275 7959
rect -241 7925 -207 7959
rect -173 7925 -139 7959
rect -105 7925 -71 7959
rect -37 7925 -3 7959
rect 31 7925 65 7959
rect 99 7925 133 7959
rect 167 7925 201 7959
rect 235 7925 269 7959
rect 303 7925 337 7959
rect 371 7925 405 7959
rect 439 7925 473 7959
rect 507 7925 541 7959
rect 575 7925 609 7959
rect 643 7925 677 7959
rect 711 7925 745 7959
rect 779 7925 813 7959
rect 847 7925 881 7959
rect 915 7925 949 7959
rect 983 7925 1017 7959
rect 1051 7925 1085 7959
rect 1119 7925 1153 7959
rect 1187 7925 1221 7959
rect 1255 7925 1289 7959
rect 1323 7925 1357 7959
rect 1391 7925 1425 7959
rect 1459 7925 1493 7959
rect 1527 7925 1561 7959
rect 1595 7925 1629 7959
rect 1663 7925 1697 7959
rect 1731 7925 1765 7959
rect 1799 7925 1833 7959
rect 1867 7925 1901 7959
rect 1935 7925 1969 7959
rect 2003 7925 2037 7959
rect 2071 7925 2105 7959
rect 2139 7925 2173 7959
rect 2207 7925 2241 7959
rect 2275 7925 2309 7959
rect 2343 7925 2377 7959
rect 2411 7925 2445 7959
rect 2479 7925 2513 7959
rect 2547 7925 2581 7959
rect 2615 7925 2649 7959
rect 2683 7925 2717 7959
rect 2751 7925 2785 7959
rect 2819 7925 2853 7959
rect 2887 7925 2921 7959
rect 2955 7925 2989 7959
rect 3023 7925 3057 7959
rect 3091 7925 3125 7959
rect 3159 7925 3193 7959
rect 3227 7925 3358 7959
rect -3058 7901 3358 7925
rect -3058 7812 -2976 7901
rect -3058 7778 -3034 7812
rect -3000 7778 -2976 7812
rect -3058 7744 -2976 7778
rect -3058 7710 -3034 7744
rect -3000 7710 -2976 7744
rect -3058 7676 -2976 7710
rect -3058 7642 -3034 7676
rect -3000 7642 -2976 7676
rect -3058 7608 -2976 7642
rect -3058 7574 -3034 7608
rect -3000 7574 -2976 7608
rect -3058 7540 -2976 7574
rect -3058 7506 -3034 7540
rect -3000 7506 -2976 7540
rect -3058 7472 -2976 7506
rect -3058 7438 -3034 7472
rect -3000 7438 -2976 7472
rect -3058 7404 -2976 7438
rect -3058 7370 -3034 7404
rect -3000 7370 -2976 7404
rect -3058 7336 -2976 7370
rect -3058 7302 -3034 7336
rect -3000 7302 -2976 7336
rect -3058 7268 -2976 7302
rect -3058 7234 -3034 7268
rect -3000 7234 -2976 7268
rect -3058 7200 -2976 7234
rect -3058 7166 -3034 7200
rect -3000 7166 -2976 7200
rect -3058 7132 -2976 7166
rect -3058 7098 -3034 7132
rect -3000 7098 -2976 7132
rect -3058 7064 -2976 7098
rect -3058 7030 -3034 7064
rect -3000 7030 -2976 7064
rect -3058 6996 -2976 7030
rect -3058 6962 -3034 6996
rect -3000 6962 -2976 6996
rect -3058 6928 -2976 6962
rect -3058 6894 -3034 6928
rect -3000 6894 -2976 6928
rect -3058 6860 -2976 6894
rect -3058 6826 -3034 6860
rect -3000 6826 -2976 6860
rect -3058 6792 -2976 6826
rect 3276 7812 3358 7901
rect 3276 7778 3300 7812
rect 3334 7778 3358 7812
rect 3276 7744 3358 7778
rect 3276 7710 3300 7744
rect 3334 7710 3358 7744
rect 3276 7676 3358 7710
rect 3276 7642 3300 7676
rect 3334 7642 3358 7676
rect 3276 7608 3358 7642
rect 3276 7574 3300 7608
rect 3334 7574 3358 7608
rect 3276 7540 3358 7574
rect 3276 7506 3300 7540
rect 3334 7506 3358 7540
rect 3276 7472 3358 7506
rect 3276 7438 3300 7472
rect 3334 7438 3358 7472
rect 3276 7404 3358 7438
rect 3276 7370 3300 7404
rect 3334 7370 3358 7404
rect 3276 7336 3358 7370
rect 3276 7302 3300 7336
rect 3334 7302 3358 7336
rect 3276 7268 3358 7302
rect 3276 7234 3300 7268
rect 3334 7234 3358 7268
rect 3276 7200 3358 7234
rect 3276 7166 3300 7200
rect 3334 7166 3358 7200
rect 3276 7132 3358 7166
rect 3276 7098 3300 7132
rect 3334 7098 3358 7132
rect 3276 7064 3358 7098
rect 3276 7030 3300 7064
rect 3334 7030 3358 7064
rect 3276 6996 3358 7030
rect 3276 6962 3300 6996
rect 3334 6962 3358 6996
rect 3276 6928 3358 6962
rect 3276 6894 3300 6928
rect 3334 6894 3358 6928
rect 3276 6860 3358 6894
rect 3276 6826 3300 6860
rect 3334 6826 3358 6860
rect -3058 6758 -3034 6792
rect -3000 6758 -2976 6792
rect -3058 6724 -2976 6758
rect -3058 6690 -3034 6724
rect -3000 6690 -2976 6724
rect -3058 6656 -2976 6690
rect -3058 6622 -3034 6656
rect -3000 6622 -2976 6656
rect -3058 6588 -2976 6622
rect -3058 6554 -3034 6588
rect -3000 6554 -2976 6588
rect -3058 6520 -2976 6554
rect -3058 6486 -3034 6520
rect -3000 6486 -2976 6520
rect -3058 6452 -2976 6486
rect -3058 6418 -3034 6452
rect -3000 6418 -2976 6452
rect -3058 6384 -2976 6418
rect -3058 6350 -3034 6384
rect -3000 6350 -2976 6384
rect -3058 6316 -2976 6350
rect -3058 6282 -3034 6316
rect -3000 6282 -2976 6316
rect -3058 6248 -2976 6282
rect -3058 6214 -3034 6248
rect -3000 6214 -2976 6248
rect -3058 6180 -2976 6214
rect -3058 6146 -3034 6180
rect -3000 6146 -2976 6180
rect -3058 6112 -2976 6146
rect -3058 6078 -3034 6112
rect -3000 6078 -2976 6112
rect -3058 6044 -2976 6078
rect -3058 6010 -3034 6044
rect -3000 6010 -2976 6044
rect -3058 5976 -2976 6010
rect 3276 6792 3358 6826
rect 3276 6758 3300 6792
rect 3334 6758 3358 6792
rect 3276 6724 3358 6758
rect 3276 6690 3300 6724
rect 3334 6690 3358 6724
rect 3276 6656 3358 6690
rect 3276 6622 3300 6656
rect 3334 6622 3358 6656
rect 3276 6588 3358 6622
rect 3276 6554 3300 6588
rect 3334 6554 3358 6588
rect 3276 6520 3358 6554
rect 3276 6486 3300 6520
rect 3334 6486 3358 6520
rect 3276 6452 3358 6486
rect 3276 6418 3300 6452
rect 3334 6418 3358 6452
rect 3276 6384 3358 6418
rect 3276 6350 3300 6384
rect 3334 6350 3358 6384
rect 3276 6316 3358 6350
rect 3276 6282 3300 6316
rect 3334 6282 3358 6316
rect 3276 6248 3358 6282
rect 3276 6214 3300 6248
rect 3334 6214 3358 6248
rect 3276 6180 3358 6214
rect 3276 6146 3300 6180
rect 3334 6146 3358 6180
rect 3276 6112 3358 6146
rect 3276 6078 3300 6112
rect 3334 6078 3358 6112
rect 3276 6044 3358 6078
rect 3276 6010 3300 6044
rect 3334 6010 3358 6044
rect -3058 5942 -3034 5976
rect -3000 5942 -2976 5976
rect -3058 5908 -2976 5942
rect -3058 5874 -3034 5908
rect -3000 5874 -2976 5908
rect -3058 5840 -2976 5874
rect -3058 5806 -3034 5840
rect -3000 5806 -2976 5840
rect -3058 5772 -2976 5806
rect -3058 5738 -3034 5772
rect -3000 5738 -2976 5772
rect -3058 5704 -2976 5738
rect -3058 5670 -3034 5704
rect -3000 5670 -2976 5704
rect -3058 5636 -2976 5670
rect -3058 5602 -3034 5636
rect -3000 5602 -2976 5636
rect -3058 5568 -2976 5602
rect -3058 5534 -3034 5568
rect -3000 5534 -2976 5568
rect -3058 5500 -2976 5534
rect -3058 5466 -3034 5500
rect -3000 5466 -2976 5500
rect -3058 5432 -2976 5466
rect -3058 5398 -3034 5432
rect -3000 5398 -2976 5432
rect -3058 5364 -2976 5398
rect -3058 5330 -3034 5364
rect -3000 5330 -2976 5364
rect -3058 5296 -2976 5330
rect -3058 5262 -3034 5296
rect -3000 5262 -2976 5296
rect -3058 5228 -2976 5262
rect -3058 5194 -3034 5228
rect -3000 5194 -2976 5228
rect -3058 5160 -2976 5194
rect -3058 5126 -3034 5160
rect -3000 5126 -2976 5160
rect -3058 5092 -2976 5126
rect -3058 5058 -3034 5092
rect -3000 5058 -2976 5092
rect -3058 5024 -2976 5058
rect -3058 4990 -3034 5024
rect -3000 4990 -2976 5024
rect -3058 4956 -2976 4990
rect -3058 4922 -3034 4956
rect -3000 4922 -2976 4956
rect -3058 4888 -2976 4922
rect -3058 4854 -3034 4888
rect -3000 4854 -2976 4888
rect -3058 4820 -2976 4854
rect -3058 4786 -3034 4820
rect -3000 4786 -2976 4820
rect -3058 4752 -2976 4786
rect -3058 4718 -3034 4752
rect -3000 4718 -2976 4752
rect -3058 4684 -2976 4718
rect -3058 4650 -3034 4684
rect -3000 4650 -2976 4684
rect -3058 4616 -2976 4650
rect -3058 4582 -3034 4616
rect -3000 4582 -2976 4616
rect -3058 4548 -2976 4582
rect -3058 4514 -3034 4548
rect -3000 4514 -2976 4548
rect -3058 4480 -2976 4514
rect -3058 4446 -3034 4480
rect -3000 4446 -2976 4480
rect -3058 4412 -2976 4446
rect -3058 4378 -3034 4412
rect -3000 4378 -2976 4412
rect -3058 4344 -2976 4378
rect -3058 4310 -3034 4344
rect -3000 4310 -2976 4344
rect -3058 4276 -2976 4310
rect -3058 4242 -3034 4276
rect -3000 4242 -2976 4276
rect -3058 4208 -2976 4242
rect -3058 4174 -3034 4208
rect -3000 4174 -2976 4208
rect -3058 4140 -2976 4174
rect -3058 4106 -3034 4140
rect -3000 4106 -2976 4140
rect -3058 4072 -2976 4106
rect -3058 4038 -3034 4072
rect -3000 4038 -2976 4072
rect -3058 4004 -2976 4038
rect -3058 3970 -3034 4004
rect -3000 3970 -2976 4004
rect -3058 3936 -2976 3970
rect -3058 3902 -3034 3936
rect -3000 3902 -2976 3936
rect -3058 3868 -2976 3902
rect -3058 3834 -3034 3868
rect -3000 3834 -2976 3868
rect -3058 3800 -2976 3834
rect -3058 3766 -3034 3800
rect -3000 3766 -2976 3800
rect -3058 3732 -2976 3766
rect -3058 3698 -3034 3732
rect -3000 3698 -2976 3732
rect -3058 3664 -2976 3698
rect -3058 3630 -3034 3664
rect -3000 3630 -2976 3664
rect -3058 3596 -2976 3630
rect -3058 3562 -3034 3596
rect -3000 3562 -2976 3596
rect -3058 3528 -2976 3562
rect -3058 3494 -3034 3528
rect -3000 3494 -2976 3528
rect -3058 3460 -2976 3494
rect -3058 3426 -3034 3460
rect -3000 3426 -2976 3460
rect -3058 3392 -2976 3426
rect -3058 3358 -3034 3392
rect -3000 3358 -2976 3392
rect -3058 3324 -2976 3358
rect -3058 3290 -3034 3324
rect -3000 3290 -2976 3324
rect -3058 3256 -2976 3290
rect -3058 3222 -3034 3256
rect -3000 3222 -2976 3256
rect -3058 3188 -2976 3222
rect -3058 3154 -3034 3188
rect -3000 3154 -2976 3188
rect -3058 3120 -2976 3154
rect -3058 3086 -3034 3120
rect -3000 3086 -2976 3120
rect -3058 3052 -2976 3086
rect -3058 3018 -3034 3052
rect -3000 3018 -2976 3052
rect -3058 2984 -2976 3018
rect -3058 2950 -3034 2984
rect -3000 2950 -2976 2984
rect -3058 2916 -2976 2950
rect -3058 2882 -3034 2916
rect -3000 2882 -2976 2916
rect -3058 2848 -2976 2882
rect -3058 2814 -3034 2848
rect -3000 2814 -2976 2848
rect -3058 2780 -2976 2814
rect -3058 2746 -3034 2780
rect -3000 2746 -2976 2780
rect -3058 2712 -2976 2746
rect -3058 2678 -3034 2712
rect -3000 2678 -2976 2712
rect -3058 2644 -2976 2678
rect -3058 2610 -3034 2644
rect -3000 2610 -2976 2644
rect -3058 2576 -2976 2610
rect -3058 2542 -3034 2576
rect -3000 2542 -2976 2576
rect -3058 2508 -2976 2542
rect -3058 2474 -3034 2508
rect -3000 2474 -2976 2508
rect -3058 2440 -2976 2474
rect -3058 2406 -3034 2440
rect -3000 2406 -2976 2440
rect -3058 2372 -2976 2406
rect -3058 2338 -3034 2372
rect -3000 2338 -2976 2372
rect -3058 2304 -2976 2338
rect -3058 2270 -3034 2304
rect -3000 2270 -2976 2304
rect -3058 2236 -2976 2270
rect -3058 2202 -3034 2236
rect -3000 2202 -2976 2236
rect -3058 2168 -2976 2202
rect -3058 2134 -3034 2168
rect -3000 2134 -2976 2168
rect -3058 2100 -2976 2134
rect -3058 2066 -3034 2100
rect -3000 2066 -2976 2100
rect -3058 2032 -2976 2066
rect -3058 1998 -3034 2032
rect -3000 1998 -2976 2032
rect -3058 1964 -2976 1998
rect -3058 1930 -3034 1964
rect -3000 1930 -2976 1964
rect -3058 1896 -2976 1930
rect -3058 1862 -3034 1896
rect -3000 1862 -2976 1896
rect -3058 1828 -2976 1862
rect -3058 1794 -3034 1828
rect -3000 1794 -2976 1828
rect -3058 1760 -2976 1794
rect -3058 1726 -3034 1760
rect -3000 1726 -2976 1760
rect -3058 1692 -2976 1726
rect -3058 1658 -3034 1692
rect -3000 1658 -2976 1692
rect -3058 1624 -2976 1658
rect -3058 1590 -3034 1624
rect -3000 1590 -2976 1624
rect -3058 1556 -2976 1590
rect -3058 1522 -3034 1556
rect -3000 1522 -2976 1556
rect -3058 1488 -2976 1522
rect -3058 1454 -3034 1488
rect -3000 1454 -2976 1488
rect -3058 1420 -2976 1454
rect -3058 1386 -3034 1420
rect -3000 1386 -2976 1420
rect -3058 1352 -2976 1386
rect -3058 1318 -3034 1352
rect -3000 1318 -2976 1352
rect -3058 1284 -2976 1318
rect -3058 1250 -3034 1284
rect -3000 1250 -2976 1284
rect -3058 1216 -2976 1250
rect -3058 1182 -3034 1216
rect -3000 1182 -2976 1216
rect -3058 1148 -2976 1182
rect -3058 1114 -3034 1148
rect -3000 1114 -2976 1148
rect -3058 1080 -2976 1114
rect -3058 1046 -3034 1080
rect -3000 1046 -2976 1080
rect -3058 1012 -2976 1046
rect -3058 978 -3034 1012
rect -3000 978 -2976 1012
rect -3058 944 -2976 978
rect -3058 910 -3034 944
rect -3000 910 -2976 944
rect -3058 876 -2976 910
rect -3058 842 -3034 876
rect -3000 842 -2976 876
rect -3058 808 -2976 842
rect -3058 774 -3034 808
rect -3000 774 -2976 808
rect -3058 740 -2976 774
rect -3058 706 -3034 740
rect -3000 706 -2976 740
rect -3058 672 -2976 706
rect -3058 638 -3034 672
rect -3000 638 -2976 672
rect -3058 604 -2976 638
rect -3058 570 -3034 604
rect -3000 570 -2976 604
rect -3058 536 -2976 570
rect -3058 502 -3034 536
rect -3000 502 -2976 536
rect -3058 468 -2976 502
rect -3058 434 -3034 468
rect -3000 434 -2976 468
rect -3058 400 -2976 434
rect -3058 366 -3034 400
rect -3000 366 -2976 400
rect -3058 332 -2976 366
rect -3058 298 -3034 332
rect -3000 298 -2976 332
rect -3058 264 -2976 298
rect -3058 230 -3034 264
rect -3000 230 -2976 264
rect -3058 196 -2976 230
rect -3058 162 -3034 196
rect -3000 162 -2976 196
rect -3058 128 -2976 162
rect -3058 94 -3034 128
rect -3000 94 -2976 128
rect -3058 60 -2976 94
rect -3058 26 -3034 60
rect -3000 26 -2976 60
rect -3058 -8 -2976 26
rect -1076 5975 -926 6000
rect -1076 25 -1052 5975
rect -950 25 -926 5975
rect -1076 0 -926 25
rect 1226 5975 1376 6000
rect 1226 25 1250 5975
rect 1352 25 1376 5975
rect 1226 0 1376 25
rect 3276 5976 3358 6010
rect 3276 5942 3300 5976
rect 3334 5942 3358 5976
rect 3276 5908 3358 5942
rect 3276 5874 3300 5908
rect 3334 5874 3358 5908
rect 3276 5840 3358 5874
rect 3276 5806 3300 5840
rect 3334 5806 3358 5840
rect 3276 5772 3358 5806
rect 3276 5738 3300 5772
rect 3334 5738 3358 5772
rect 3276 5704 3358 5738
rect 3276 5670 3300 5704
rect 3334 5670 3358 5704
rect 3276 5636 3358 5670
rect 3276 5602 3300 5636
rect 3334 5602 3358 5636
rect 3276 5568 3358 5602
rect 3276 5534 3300 5568
rect 3334 5534 3358 5568
rect 3276 5500 3358 5534
rect 3276 5466 3300 5500
rect 3334 5466 3358 5500
rect 3276 5432 3358 5466
rect 3276 5398 3300 5432
rect 3334 5398 3358 5432
rect 3276 5364 3358 5398
rect 3276 5330 3300 5364
rect 3334 5330 3358 5364
rect 3276 5296 3358 5330
rect 3276 5262 3300 5296
rect 3334 5262 3358 5296
rect 3276 5228 3358 5262
rect 3276 5194 3300 5228
rect 3334 5194 3358 5228
rect 3276 5160 3358 5194
rect 3276 5126 3300 5160
rect 3334 5126 3358 5160
rect 3276 5092 3358 5126
rect 3276 5058 3300 5092
rect 3334 5058 3358 5092
rect 3276 5024 3358 5058
rect 3276 4990 3300 5024
rect 3334 4990 3358 5024
rect 3276 4956 3358 4990
rect 3276 4922 3300 4956
rect 3334 4922 3358 4956
rect 3276 4888 3358 4922
rect 3276 4854 3300 4888
rect 3334 4854 3358 4888
rect 3276 4820 3358 4854
rect 3276 4786 3300 4820
rect 3334 4786 3358 4820
rect 3276 4752 3358 4786
rect 3276 4718 3300 4752
rect 3334 4718 3358 4752
rect 3276 4684 3358 4718
rect 3276 4650 3300 4684
rect 3334 4650 3358 4684
rect 3276 4616 3358 4650
rect 3276 4582 3300 4616
rect 3334 4582 3358 4616
rect 3276 4548 3358 4582
rect 3276 4514 3300 4548
rect 3334 4514 3358 4548
rect 3276 4480 3358 4514
rect 3276 4446 3300 4480
rect 3334 4446 3358 4480
rect 3276 4412 3358 4446
rect 3276 4378 3300 4412
rect 3334 4378 3358 4412
rect 3276 4344 3358 4378
rect 3276 4310 3300 4344
rect 3334 4310 3358 4344
rect 3276 4276 3358 4310
rect 3276 4242 3300 4276
rect 3334 4242 3358 4276
rect 3276 4208 3358 4242
rect 3276 4174 3300 4208
rect 3334 4174 3358 4208
rect 3276 4140 3358 4174
rect 3276 4106 3300 4140
rect 3334 4106 3358 4140
rect 3276 4072 3358 4106
rect 3276 4038 3300 4072
rect 3334 4038 3358 4072
rect 3276 4004 3358 4038
rect 3276 3970 3300 4004
rect 3334 3970 3358 4004
rect 3276 3936 3358 3970
rect 3276 3902 3300 3936
rect 3334 3902 3358 3936
rect 3276 3868 3358 3902
rect 3276 3834 3300 3868
rect 3334 3834 3358 3868
rect 3276 3800 3358 3834
rect 3276 3766 3300 3800
rect 3334 3766 3358 3800
rect 3276 3732 3358 3766
rect 3276 3698 3300 3732
rect 3334 3698 3358 3732
rect 3276 3664 3358 3698
rect 3276 3630 3300 3664
rect 3334 3630 3358 3664
rect 3276 3596 3358 3630
rect 3276 3562 3300 3596
rect 3334 3562 3358 3596
rect 3276 3528 3358 3562
rect 3276 3494 3300 3528
rect 3334 3494 3358 3528
rect 3276 3460 3358 3494
rect 3276 3426 3300 3460
rect 3334 3426 3358 3460
rect 3276 3392 3358 3426
rect 3276 3358 3300 3392
rect 3334 3358 3358 3392
rect 3276 3324 3358 3358
rect 3276 3290 3300 3324
rect 3334 3290 3358 3324
rect 3276 3256 3358 3290
rect 3276 3222 3300 3256
rect 3334 3222 3358 3256
rect 3276 3188 3358 3222
rect 3276 3154 3300 3188
rect 3334 3154 3358 3188
rect 3276 3120 3358 3154
rect 3276 3086 3300 3120
rect 3334 3086 3358 3120
rect 3276 3052 3358 3086
rect 3276 3018 3300 3052
rect 3334 3018 3358 3052
rect 3276 2984 3358 3018
rect 3276 2950 3300 2984
rect 3334 2950 3358 2984
rect 3276 2916 3358 2950
rect 3276 2882 3300 2916
rect 3334 2882 3358 2916
rect 3276 2848 3358 2882
rect 3276 2814 3300 2848
rect 3334 2814 3358 2848
rect 3276 2780 3358 2814
rect 3276 2746 3300 2780
rect 3334 2746 3358 2780
rect 3276 2712 3358 2746
rect 3276 2678 3300 2712
rect 3334 2678 3358 2712
rect 3276 2644 3358 2678
rect 3276 2610 3300 2644
rect 3334 2610 3358 2644
rect 3276 2576 3358 2610
rect 3276 2542 3300 2576
rect 3334 2542 3358 2576
rect 3276 2508 3358 2542
rect 3276 2474 3300 2508
rect 3334 2474 3358 2508
rect 3276 2440 3358 2474
rect 3276 2406 3300 2440
rect 3334 2406 3358 2440
rect 3276 2372 3358 2406
rect 3276 2338 3300 2372
rect 3334 2338 3358 2372
rect 3276 2304 3358 2338
rect 3276 2270 3300 2304
rect 3334 2270 3358 2304
rect 3276 2236 3358 2270
rect 3276 2202 3300 2236
rect 3334 2202 3358 2236
rect 3276 2168 3358 2202
rect 3276 2134 3300 2168
rect 3334 2134 3358 2168
rect 3276 2100 3358 2134
rect 3276 2066 3300 2100
rect 3334 2066 3358 2100
rect 3276 2032 3358 2066
rect 3276 1998 3300 2032
rect 3334 1998 3358 2032
rect 3276 1964 3358 1998
rect 3276 1930 3300 1964
rect 3334 1930 3358 1964
rect 3276 1896 3358 1930
rect 3276 1862 3300 1896
rect 3334 1862 3358 1896
rect 3276 1828 3358 1862
rect 3276 1794 3300 1828
rect 3334 1794 3358 1828
rect 3276 1760 3358 1794
rect 3276 1726 3300 1760
rect 3334 1726 3358 1760
rect 3276 1692 3358 1726
rect 3276 1658 3300 1692
rect 3334 1658 3358 1692
rect 3276 1624 3358 1658
rect 3276 1590 3300 1624
rect 3334 1590 3358 1624
rect 3276 1556 3358 1590
rect 3276 1522 3300 1556
rect 3334 1522 3358 1556
rect 3276 1488 3358 1522
rect 3276 1454 3300 1488
rect 3334 1454 3358 1488
rect 3276 1420 3358 1454
rect 3276 1386 3300 1420
rect 3334 1386 3358 1420
rect 3276 1352 3358 1386
rect 3276 1318 3300 1352
rect 3334 1318 3358 1352
rect 3276 1284 3358 1318
rect 3276 1250 3300 1284
rect 3334 1250 3358 1284
rect 3276 1216 3358 1250
rect 3276 1182 3300 1216
rect 3334 1182 3358 1216
rect 3276 1148 3358 1182
rect 3276 1114 3300 1148
rect 3334 1114 3358 1148
rect 3276 1080 3358 1114
rect 3276 1046 3300 1080
rect 3334 1046 3358 1080
rect 3276 1012 3358 1046
rect 3276 978 3300 1012
rect 3334 978 3358 1012
rect 3276 944 3358 978
rect 3276 910 3300 944
rect 3334 910 3358 944
rect 3276 876 3358 910
rect 3276 842 3300 876
rect 3334 842 3358 876
rect 3276 808 3358 842
rect 3276 774 3300 808
rect 3334 774 3358 808
rect 3276 740 3358 774
rect 3276 706 3300 740
rect 3334 706 3358 740
rect 3276 672 3358 706
rect 3276 638 3300 672
rect 3334 638 3358 672
rect 3276 604 3358 638
rect 3276 570 3300 604
rect 3334 570 3358 604
rect 3276 536 3358 570
rect 3276 502 3300 536
rect 3334 502 3358 536
rect 3276 468 3358 502
rect 3276 434 3300 468
rect 3334 434 3358 468
rect 3276 400 3358 434
rect 3276 366 3300 400
rect 3334 366 3358 400
rect 3276 332 3358 366
rect 3276 298 3300 332
rect 3334 298 3358 332
rect 3276 264 3358 298
rect 3276 230 3300 264
rect 3334 230 3358 264
rect 3276 196 3358 230
rect 3276 162 3300 196
rect 3334 162 3358 196
rect 3276 128 3358 162
rect 3276 94 3300 128
rect 3334 94 3358 128
rect 3276 60 3358 94
rect 3276 26 3300 60
rect 3334 26 3358 60
rect -3058 -42 -3034 -8
rect -3000 -42 -2976 -8
rect -3058 -76 -2976 -42
rect -3058 -110 -3034 -76
rect -3000 -110 -2976 -76
rect -3058 -144 -2976 -110
rect -3058 -178 -3034 -144
rect -3000 -178 -2976 -144
rect -3058 -212 -2976 -178
rect -3058 -246 -3034 -212
rect -3000 -246 -2976 -212
rect -3058 -280 -2976 -246
rect -3058 -314 -3034 -280
rect -3000 -314 -2976 -280
rect -3058 -348 -2976 -314
rect -3058 -382 -3034 -348
rect -3000 -382 -2976 -348
rect -3058 -416 -2976 -382
rect -3058 -450 -3034 -416
rect -3000 -450 -2976 -416
rect -3058 -484 -2976 -450
rect -3058 -518 -3034 -484
rect -3000 -518 -2976 -484
rect -3058 -552 -2976 -518
rect -3058 -586 -3034 -552
rect -3000 -586 -2976 -552
rect -3058 -620 -2976 -586
rect -3058 -654 -3034 -620
rect -3000 -654 -2976 -620
rect -3058 -688 -2976 -654
rect -3058 -722 -3034 -688
rect -3000 -722 -2976 -688
rect -3058 -756 -2976 -722
rect -3058 -790 -3034 -756
rect -3000 -790 -2976 -756
rect -3058 -824 -2976 -790
rect 3276 -8 3358 26
rect 3276 -42 3300 -8
rect 3334 -42 3358 -8
rect 3276 -76 3358 -42
rect 3276 -110 3300 -76
rect 3334 -110 3358 -76
rect 3276 -144 3358 -110
rect 3276 -178 3300 -144
rect 3334 -178 3358 -144
rect 3276 -212 3358 -178
rect 3276 -246 3300 -212
rect 3334 -246 3358 -212
rect 3276 -280 3358 -246
rect 3276 -314 3300 -280
rect 3334 -314 3358 -280
rect 3276 -348 3358 -314
rect 3276 -382 3300 -348
rect 3334 -382 3358 -348
rect 3276 -416 3358 -382
rect 3276 -450 3300 -416
rect 3334 -450 3358 -416
rect 3276 -484 3358 -450
rect 3276 -518 3300 -484
rect 3334 -518 3358 -484
rect 3276 -552 3358 -518
rect 3276 -586 3300 -552
rect 3334 -586 3358 -552
rect 3276 -620 3358 -586
rect 3276 -654 3300 -620
rect 3334 -654 3358 -620
rect 3276 -688 3358 -654
rect 3276 -722 3300 -688
rect 3334 -722 3358 -688
rect 3276 -756 3358 -722
rect 3276 -790 3300 -756
rect 3334 -790 3358 -756
rect -3058 -858 -3034 -824
rect -3000 -858 -2976 -824
rect -3058 -892 -2976 -858
rect -3058 -926 -3034 -892
rect -3000 -926 -2976 -892
rect -3058 -960 -2976 -926
rect -3058 -994 -3034 -960
rect -3000 -994 -2976 -960
rect -3058 -1028 -2976 -994
rect -3058 -1062 -3034 -1028
rect -3000 -1062 -2976 -1028
rect -3058 -1096 -2976 -1062
rect -3058 -1130 -3034 -1096
rect -3000 -1130 -2976 -1096
rect -3058 -1164 -2976 -1130
rect -3058 -1198 -3034 -1164
rect -3000 -1198 -2976 -1164
rect -3058 -1232 -2976 -1198
rect -3058 -1266 -3034 -1232
rect -3000 -1266 -2976 -1232
rect -3058 -1300 -2976 -1266
rect -3058 -1334 -3034 -1300
rect -3000 -1334 -2976 -1300
rect -3058 -1368 -2976 -1334
rect -3058 -1402 -3034 -1368
rect -3000 -1402 -2976 -1368
rect -3058 -1436 -2976 -1402
rect -3058 -1470 -3034 -1436
rect -3000 -1470 -2976 -1436
rect -3058 -1504 -2976 -1470
rect -3058 -1538 -3034 -1504
rect -3000 -1538 -2976 -1504
rect -3058 -1572 -2976 -1538
rect -3058 -1606 -3034 -1572
rect -3000 -1606 -2976 -1572
rect -3058 -1640 -2976 -1606
rect -3058 -1674 -3034 -1640
rect -3000 -1674 -2976 -1640
rect -3058 -1708 -2976 -1674
rect -3058 -1742 -3034 -1708
rect -3000 -1742 -2976 -1708
rect -3058 -1776 -2976 -1742
rect -3058 -1810 -3034 -1776
rect -3000 -1810 -2976 -1776
rect -3058 -1900 -2976 -1810
rect 3276 -824 3358 -790
rect 3276 -858 3300 -824
rect 3334 -858 3358 -824
rect 3276 -892 3358 -858
rect 3276 -926 3300 -892
rect 3334 -926 3358 -892
rect 3276 -960 3358 -926
rect 3276 -994 3300 -960
rect 3334 -994 3358 -960
rect 3276 -1028 3358 -994
rect 3276 -1062 3300 -1028
rect 3334 -1062 3358 -1028
rect 3276 -1096 3358 -1062
rect 3276 -1130 3300 -1096
rect 3334 -1130 3358 -1096
rect 3276 -1164 3358 -1130
rect 3276 -1198 3300 -1164
rect 3334 -1198 3358 -1164
rect 3276 -1232 3358 -1198
rect 3276 -1266 3300 -1232
rect 3334 -1266 3358 -1232
rect 3276 -1300 3358 -1266
rect 3276 -1334 3300 -1300
rect 3334 -1334 3358 -1300
rect 3276 -1368 3358 -1334
rect 3276 -1402 3300 -1368
rect 3334 -1402 3358 -1368
rect 3276 -1436 3358 -1402
rect 3276 -1470 3300 -1436
rect 3334 -1470 3358 -1436
rect 3276 -1504 3358 -1470
rect 3276 -1538 3300 -1504
rect 3334 -1538 3358 -1504
rect 3276 -1572 3358 -1538
rect 3276 -1606 3300 -1572
rect 3334 -1606 3358 -1572
rect 3276 -1640 3358 -1606
rect 3276 -1674 3300 -1640
rect 3334 -1674 3358 -1640
rect 3276 -1708 3358 -1674
rect 3276 -1742 3300 -1708
rect 3334 -1742 3358 -1708
rect 3276 -1776 3358 -1742
rect 3276 -1810 3300 -1776
rect 3334 -1810 3358 -1776
rect 3276 -1900 3358 -1810
rect -3058 -1924 3358 -1900
rect -3058 -1958 -2927 -1924
rect -2893 -1958 -2859 -1924
rect -2825 -1958 -2791 -1924
rect -2757 -1958 -2723 -1924
rect -2689 -1958 -2655 -1924
rect -2621 -1958 -2587 -1924
rect -2553 -1958 -2519 -1924
rect -2485 -1958 -2451 -1924
rect -2417 -1958 -2383 -1924
rect -2349 -1958 -2315 -1924
rect -2281 -1958 -2247 -1924
rect -2213 -1958 -2179 -1924
rect -2145 -1958 -2111 -1924
rect -2077 -1958 -2043 -1924
rect -2009 -1958 -1975 -1924
rect -1941 -1958 -1907 -1924
rect -1873 -1958 -1839 -1924
rect -1805 -1958 -1771 -1924
rect -1737 -1958 -1703 -1924
rect -1669 -1958 -1635 -1924
rect -1601 -1958 -1567 -1924
rect -1533 -1958 -1499 -1924
rect -1465 -1958 -1431 -1924
rect -1397 -1958 -1363 -1924
rect -1329 -1958 -1295 -1924
rect -1261 -1958 -1227 -1924
rect -1193 -1958 -1159 -1924
rect -1125 -1958 -1091 -1924
rect -1057 -1958 -1023 -1924
rect -989 -1958 -955 -1924
rect -921 -1958 -887 -1924
rect -853 -1958 -819 -1924
rect -785 -1958 -751 -1924
rect -717 -1958 -683 -1924
rect -649 -1958 -615 -1924
rect -581 -1958 -547 -1924
rect -513 -1958 -479 -1924
rect -445 -1958 -411 -1924
rect -377 -1958 -343 -1924
rect -309 -1958 -275 -1924
rect -241 -1958 -207 -1924
rect -173 -1958 -139 -1924
rect -105 -1958 -71 -1924
rect -37 -1958 -3 -1924
rect 31 -1958 65 -1924
rect 99 -1958 133 -1924
rect 167 -1958 201 -1924
rect 235 -1958 269 -1924
rect 303 -1958 337 -1924
rect 371 -1958 405 -1924
rect 439 -1958 473 -1924
rect 507 -1958 541 -1924
rect 575 -1958 609 -1924
rect 643 -1958 677 -1924
rect 711 -1958 745 -1924
rect 779 -1958 813 -1924
rect 847 -1958 881 -1924
rect 915 -1958 949 -1924
rect 983 -1958 1017 -1924
rect 1051 -1958 1085 -1924
rect 1119 -1958 1153 -1924
rect 1187 -1958 1221 -1924
rect 1255 -1958 1289 -1924
rect 1323 -1958 1357 -1924
rect 1391 -1958 1425 -1924
rect 1459 -1958 1493 -1924
rect 1527 -1958 1561 -1924
rect 1595 -1958 1629 -1924
rect 1663 -1958 1697 -1924
rect 1731 -1958 1765 -1924
rect 1799 -1958 1833 -1924
rect 1867 -1958 1901 -1924
rect 1935 -1958 1969 -1924
rect 2003 -1958 2037 -1924
rect 2071 -1958 2105 -1924
rect 2139 -1958 2173 -1924
rect 2207 -1958 2241 -1924
rect 2275 -1958 2309 -1924
rect 2343 -1958 2377 -1924
rect 2411 -1958 2445 -1924
rect 2479 -1958 2513 -1924
rect 2547 -1958 2581 -1924
rect 2615 -1958 2649 -1924
rect 2683 -1958 2717 -1924
rect 2751 -1958 2785 -1924
rect 2819 -1958 2853 -1924
rect 2887 -1958 2921 -1924
rect 2955 -1958 2989 -1924
rect 3023 -1958 3057 -1924
rect 3091 -1958 3125 -1924
rect 3159 -1958 3193 -1924
rect 3227 -1958 3358 -1924
rect -3058 -1982 3358 -1958
<< mvnsubdiff >>
tri 0 5970 30 6000 se
rect 30 5970 270 6000
tri 270 5970 300 6000 sw
rect 0 5941 300 5970
rect 0 59 31 5941
rect 269 59 300 5941
rect 0 30 300 59
tri 0 0 30 30 ne
rect 30 0 270 30
tri 270 0 300 30 nw
<< mvpsubdiffcont >>
rect -2927 7925 -2893 7959
rect -2859 7925 -2825 7959
rect -2791 7925 -2757 7959
rect -2723 7925 -2689 7959
rect -2655 7925 -2621 7959
rect -2587 7925 -2553 7959
rect -2519 7925 -2485 7959
rect -2451 7925 -2417 7959
rect -2383 7925 -2349 7959
rect -2315 7925 -2281 7959
rect -2247 7925 -2213 7959
rect -2179 7925 -2145 7959
rect -2111 7925 -2077 7959
rect -2043 7925 -2009 7959
rect -1975 7925 -1941 7959
rect -1907 7925 -1873 7959
rect -1839 7925 -1805 7959
rect -1771 7925 -1737 7959
rect -1703 7925 -1669 7959
rect -1635 7925 -1601 7959
rect -1567 7925 -1533 7959
rect -1499 7925 -1465 7959
rect -1431 7925 -1397 7959
rect -1363 7925 -1329 7959
rect -1295 7925 -1261 7959
rect -1227 7925 -1193 7959
rect -1159 7925 -1125 7959
rect -1091 7925 -1057 7959
rect -1023 7925 -989 7959
rect -955 7925 -921 7959
rect -887 7925 -853 7959
rect -819 7925 -785 7959
rect -751 7925 -717 7959
rect -683 7925 -649 7959
rect -615 7925 -581 7959
rect -547 7925 -513 7959
rect -479 7925 -445 7959
rect -411 7925 -377 7959
rect -343 7925 -309 7959
rect -275 7925 -241 7959
rect -207 7925 -173 7959
rect -139 7925 -105 7959
rect -71 7925 -37 7959
rect -3 7925 31 7959
rect 65 7925 99 7959
rect 133 7925 167 7959
rect 201 7925 235 7959
rect 269 7925 303 7959
rect 337 7925 371 7959
rect 405 7925 439 7959
rect 473 7925 507 7959
rect 541 7925 575 7959
rect 609 7925 643 7959
rect 677 7925 711 7959
rect 745 7925 779 7959
rect 813 7925 847 7959
rect 881 7925 915 7959
rect 949 7925 983 7959
rect 1017 7925 1051 7959
rect 1085 7925 1119 7959
rect 1153 7925 1187 7959
rect 1221 7925 1255 7959
rect 1289 7925 1323 7959
rect 1357 7925 1391 7959
rect 1425 7925 1459 7959
rect 1493 7925 1527 7959
rect 1561 7925 1595 7959
rect 1629 7925 1663 7959
rect 1697 7925 1731 7959
rect 1765 7925 1799 7959
rect 1833 7925 1867 7959
rect 1901 7925 1935 7959
rect 1969 7925 2003 7959
rect 2037 7925 2071 7959
rect 2105 7925 2139 7959
rect 2173 7925 2207 7959
rect 2241 7925 2275 7959
rect 2309 7925 2343 7959
rect 2377 7925 2411 7959
rect 2445 7925 2479 7959
rect 2513 7925 2547 7959
rect 2581 7925 2615 7959
rect 2649 7925 2683 7959
rect 2717 7925 2751 7959
rect 2785 7925 2819 7959
rect 2853 7925 2887 7959
rect 2921 7925 2955 7959
rect 2989 7925 3023 7959
rect 3057 7925 3091 7959
rect 3125 7925 3159 7959
rect 3193 7925 3227 7959
rect -3034 7778 -3000 7812
rect -3034 7710 -3000 7744
rect -3034 7642 -3000 7676
rect -3034 7574 -3000 7608
rect -3034 7506 -3000 7540
rect -3034 7438 -3000 7472
rect -3034 7370 -3000 7404
rect -3034 7302 -3000 7336
rect -3034 7234 -3000 7268
rect -3034 7166 -3000 7200
rect -3034 7098 -3000 7132
rect -3034 7030 -3000 7064
rect -3034 6962 -3000 6996
rect -3034 6894 -3000 6928
rect -3034 6826 -3000 6860
rect 3300 7778 3334 7812
rect 3300 7710 3334 7744
rect 3300 7642 3334 7676
rect 3300 7574 3334 7608
rect 3300 7506 3334 7540
rect 3300 7438 3334 7472
rect 3300 7370 3334 7404
rect 3300 7302 3334 7336
rect 3300 7234 3334 7268
rect 3300 7166 3334 7200
rect 3300 7098 3334 7132
rect 3300 7030 3334 7064
rect 3300 6962 3334 6996
rect 3300 6894 3334 6928
rect 3300 6826 3334 6860
rect -3034 6758 -3000 6792
rect -3034 6690 -3000 6724
rect -3034 6622 -3000 6656
rect -3034 6554 -3000 6588
rect -3034 6486 -3000 6520
rect -3034 6418 -3000 6452
rect -3034 6350 -3000 6384
rect -3034 6282 -3000 6316
rect -3034 6214 -3000 6248
rect -3034 6146 -3000 6180
rect -3034 6078 -3000 6112
rect -3034 6010 -3000 6044
rect 3300 6758 3334 6792
rect 3300 6690 3334 6724
rect 3300 6622 3334 6656
rect 3300 6554 3334 6588
rect 3300 6486 3334 6520
rect 3300 6418 3334 6452
rect 3300 6350 3334 6384
rect 3300 6282 3334 6316
rect 3300 6214 3334 6248
rect 3300 6146 3334 6180
rect 3300 6078 3334 6112
rect 3300 6010 3334 6044
rect -3034 5942 -3000 5976
rect -3034 5874 -3000 5908
rect -3034 5806 -3000 5840
rect -3034 5738 -3000 5772
rect -3034 5670 -3000 5704
rect -3034 5602 -3000 5636
rect -3034 5534 -3000 5568
rect -3034 5466 -3000 5500
rect -3034 5398 -3000 5432
rect -3034 5330 -3000 5364
rect -3034 5262 -3000 5296
rect -3034 5194 -3000 5228
rect -3034 5126 -3000 5160
rect -3034 5058 -3000 5092
rect -3034 4990 -3000 5024
rect -3034 4922 -3000 4956
rect -3034 4854 -3000 4888
rect -3034 4786 -3000 4820
rect -3034 4718 -3000 4752
rect -3034 4650 -3000 4684
rect -3034 4582 -3000 4616
rect -3034 4514 -3000 4548
rect -3034 4446 -3000 4480
rect -3034 4378 -3000 4412
rect -3034 4310 -3000 4344
rect -3034 4242 -3000 4276
rect -3034 4174 -3000 4208
rect -3034 4106 -3000 4140
rect -3034 4038 -3000 4072
rect -3034 3970 -3000 4004
rect -3034 3902 -3000 3936
rect -3034 3834 -3000 3868
rect -3034 3766 -3000 3800
rect -3034 3698 -3000 3732
rect -3034 3630 -3000 3664
rect -3034 3562 -3000 3596
rect -3034 3494 -3000 3528
rect -3034 3426 -3000 3460
rect -3034 3358 -3000 3392
rect -3034 3290 -3000 3324
rect -3034 3222 -3000 3256
rect -3034 3154 -3000 3188
rect -3034 3086 -3000 3120
rect -3034 3018 -3000 3052
rect -3034 2950 -3000 2984
rect -3034 2882 -3000 2916
rect -3034 2814 -3000 2848
rect -3034 2746 -3000 2780
rect -3034 2678 -3000 2712
rect -3034 2610 -3000 2644
rect -3034 2542 -3000 2576
rect -3034 2474 -3000 2508
rect -3034 2406 -3000 2440
rect -3034 2338 -3000 2372
rect -3034 2270 -3000 2304
rect -3034 2202 -3000 2236
rect -3034 2134 -3000 2168
rect -3034 2066 -3000 2100
rect -3034 1998 -3000 2032
rect -3034 1930 -3000 1964
rect -3034 1862 -3000 1896
rect -3034 1794 -3000 1828
rect -3034 1726 -3000 1760
rect -3034 1658 -3000 1692
rect -3034 1590 -3000 1624
rect -3034 1522 -3000 1556
rect -3034 1454 -3000 1488
rect -3034 1386 -3000 1420
rect -3034 1318 -3000 1352
rect -3034 1250 -3000 1284
rect -3034 1182 -3000 1216
rect -3034 1114 -3000 1148
rect -3034 1046 -3000 1080
rect -3034 978 -3000 1012
rect -3034 910 -3000 944
rect -3034 842 -3000 876
rect -3034 774 -3000 808
rect -3034 706 -3000 740
rect -3034 638 -3000 672
rect -3034 570 -3000 604
rect -3034 502 -3000 536
rect -3034 434 -3000 468
rect -3034 366 -3000 400
rect -3034 298 -3000 332
rect -3034 230 -3000 264
rect -3034 162 -3000 196
rect -3034 94 -3000 128
rect -3034 26 -3000 60
rect -1052 25 -950 5975
rect 1250 25 1352 5975
rect 3300 5942 3334 5976
rect 3300 5874 3334 5908
rect 3300 5806 3334 5840
rect 3300 5738 3334 5772
rect 3300 5670 3334 5704
rect 3300 5602 3334 5636
rect 3300 5534 3334 5568
rect 3300 5466 3334 5500
rect 3300 5398 3334 5432
rect 3300 5330 3334 5364
rect 3300 5262 3334 5296
rect 3300 5194 3334 5228
rect 3300 5126 3334 5160
rect 3300 5058 3334 5092
rect 3300 4990 3334 5024
rect 3300 4922 3334 4956
rect 3300 4854 3334 4888
rect 3300 4786 3334 4820
rect 3300 4718 3334 4752
rect 3300 4650 3334 4684
rect 3300 4582 3334 4616
rect 3300 4514 3334 4548
rect 3300 4446 3334 4480
rect 3300 4378 3334 4412
rect 3300 4310 3334 4344
rect 3300 4242 3334 4276
rect 3300 4174 3334 4208
rect 3300 4106 3334 4140
rect 3300 4038 3334 4072
rect 3300 3970 3334 4004
rect 3300 3902 3334 3936
rect 3300 3834 3334 3868
rect 3300 3766 3334 3800
rect 3300 3698 3334 3732
rect 3300 3630 3334 3664
rect 3300 3562 3334 3596
rect 3300 3494 3334 3528
rect 3300 3426 3334 3460
rect 3300 3358 3334 3392
rect 3300 3290 3334 3324
rect 3300 3222 3334 3256
rect 3300 3154 3334 3188
rect 3300 3086 3334 3120
rect 3300 3018 3334 3052
rect 3300 2950 3334 2984
rect 3300 2882 3334 2916
rect 3300 2814 3334 2848
rect 3300 2746 3334 2780
rect 3300 2678 3334 2712
rect 3300 2610 3334 2644
rect 3300 2542 3334 2576
rect 3300 2474 3334 2508
rect 3300 2406 3334 2440
rect 3300 2338 3334 2372
rect 3300 2270 3334 2304
rect 3300 2202 3334 2236
rect 3300 2134 3334 2168
rect 3300 2066 3334 2100
rect 3300 1998 3334 2032
rect 3300 1930 3334 1964
rect 3300 1862 3334 1896
rect 3300 1794 3334 1828
rect 3300 1726 3334 1760
rect 3300 1658 3334 1692
rect 3300 1590 3334 1624
rect 3300 1522 3334 1556
rect 3300 1454 3334 1488
rect 3300 1386 3334 1420
rect 3300 1318 3334 1352
rect 3300 1250 3334 1284
rect 3300 1182 3334 1216
rect 3300 1114 3334 1148
rect 3300 1046 3334 1080
rect 3300 978 3334 1012
rect 3300 910 3334 944
rect 3300 842 3334 876
rect 3300 774 3334 808
rect 3300 706 3334 740
rect 3300 638 3334 672
rect 3300 570 3334 604
rect 3300 502 3334 536
rect 3300 434 3334 468
rect 3300 366 3334 400
rect 3300 298 3334 332
rect 3300 230 3334 264
rect 3300 162 3334 196
rect 3300 94 3334 128
rect 3300 26 3334 60
rect -3034 -42 -3000 -8
rect -3034 -110 -3000 -76
rect -3034 -178 -3000 -144
rect -3034 -246 -3000 -212
rect -3034 -314 -3000 -280
rect -3034 -382 -3000 -348
rect -3034 -450 -3000 -416
rect -3034 -518 -3000 -484
rect -3034 -586 -3000 -552
rect -3034 -654 -3000 -620
rect -3034 -722 -3000 -688
rect -3034 -790 -3000 -756
rect 3300 -42 3334 -8
rect 3300 -110 3334 -76
rect 3300 -178 3334 -144
rect 3300 -246 3334 -212
rect 3300 -314 3334 -280
rect 3300 -382 3334 -348
rect 3300 -450 3334 -416
rect 3300 -518 3334 -484
rect 3300 -586 3334 -552
rect 3300 -654 3334 -620
rect 3300 -722 3334 -688
rect 3300 -790 3334 -756
rect -3034 -858 -3000 -824
rect -3034 -926 -3000 -892
rect -3034 -994 -3000 -960
rect -3034 -1062 -3000 -1028
rect -3034 -1130 -3000 -1096
rect -3034 -1198 -3000 -1164
rect -3034 -1266 -3000 -1232
rect -3034 -1334 -3000 -1300
rect -3034 -1402 -3000 -1368
rect -3034 -1470 -3000 -1436
rect -3034 -1538 -3000 -1504
rect -3034 -1606 -3000 -1572
rect -3034 -1674 -3000 -1640
rect -3034 -1742 -3000 -1708
rect -3034 -1810 -3000 -1776
rect 3300 -858 3334 -824
rect 3300 -926 3334 -892
rect 3300 -994 3334 -960
rect 3300 -1062 3334 -1028
rect 3300 -1130 3334 -1096
rect 3300 -1198 3334 -1164
rect 3300 -1266 3334 -1232
rect 3300 -1334 3334 -1300
rect 3300 -1402 3334 -1368
rect 3300 -1470 3334 -1436
rect 3300 -1538 3334 -1504
rect 3300 -1606 3334 -1572
rect 3300 -1674 3334 -1640
rect 3300 -1742 3334 -1708
rect 3300 -1810 3334 -1776
rect -2927 -1958 -2893 -1924
rect -2859 -1958 -2825 -1924
rect -2791 -1958 -2757 -1924
rect -2723 -1958 -2689 -1924
rect -2655 -1958 -2621 -1924
rect -2587 -1958 -2553 -1924
rect -2519 -1958 -2485 -1924
rect -2451 -1958 -2417 -1924
rect -2383 -1958 -2349 -1924
rect -2315 -1958 -2281 -1924
rect -2247 -1958 -2213 -1924
rect -2179 -1958 -2145 -1924
rect -2111 -1958 -2077 -1924
rect -2043 -1958 -2009 -1924
rect -1975 -1958 -1941 -1924
rect -1907 -1958 -1873 -1924
rect -1839 -1958 -1805 -1924
rect -1771 -1958 -1737 -1924
rect -1703 -1958 -1669 -1924
rect -1635 -1958 -1601 -1924
rect -1567 -1958 -1533 -1924
rect -1499 -1958 -1465 -1924
rect -1431 -1958 -1397 -1924
rect -1363 -1958 -1329 -1924
rect -1295 -1958 -1261 -1924
rect -1227 -1958 -1193 -1924
rect -1159 -1958 -1125 -1924
rect -1091 -1958 -1057 -1924
rect -1023 -1958 -989 -1924
rect -955 -1958 -921 -1924
rect -887 -1958 -853 -1924
rect -819 -1958 -785 -1924
rect -751 -1958 -717 -1924
rect -683 -1958 -649 -1924
rect -615 -1958 -581 -1924
rect -547 -1958 -513 -1924
rect -479 -1958 -445 -1924
rect -411 -1958 -377 -1924
rect -343 -1958 -309 -1924
rect -275 -1958 -241 -1924
rect -207 -1958 -173 -1924
rect -139 -1958 -105 -1924
rect -71 -1958 -37 -1924
rect -3 -1958 31 -1924
rect 65 -1958 99 -1924
rect 133 -1958 167 -1924
rect 201 -1958 235 -1924
rect 269 -1958 303 -1924
rect 337 -1958 371 -1924
rect 405 -1958 439 -1924
rect 473 -1958 507 -1924
rect 541 -1958 575 -1924
rect 609 -1958 643 -1924
rect 677 -1958 711 -1924
rect 745 -1958 779 -1924
rect 813 -1958 847 -1924
rect 881 -1958 915 -1924
rect 949 -1958 983 -1924
rect 1017 -1958 1051 -1924
rect 1085 -1958 1119 -1924
rect 1153 -1958 1187 -1924
rect 1221 -1958 1255 -1924
rect 1289 -1958 1323 -1924
rect 1357 -1958 1391 -1924
rect 1425 -1958 1459 -1924
rect 1493 -1958 1527 -1924
rect 1561 -1958 1595 -1924
rect 1629 -1958 1663 -1924
rect 1697 -1958 1731 -1924
rect 1765 -1958 1799 -1924
rect 1833 -1958 1867 -1924
rect 1901 -1958 1935 -1924
rect 1969 -1958 2003 -1924
rect 2037 -1958 2071 -1924
rect 2105 -1958 2139 -1924
rect 2173 -1958 2207 -1924
rect 2241 -1958 2275 -1924
rect 2309 -1958 2343 -1924
rect 2377 -1958 2411 -1924
rect 2445 -1958 2479 -1924
rect 2513 -1958 2547 -1924
rect 2581 -1958 2615 -1924
rect 2649 -1958 2683 -1924
rect 2717 -1958 2751 -1924
rect 2785 -1958 2819 -1924
rect 2853 -1958 2887 -1924
rect 2921 -1958 2955 -1924
rect 2989 -1958 3023 -1924
rect 3057 -1958 3091 -1924
rect 3125 -1958 3159 -1924
rect 3193 -1958 3227 -1924
<< mvnsubdiffcont >>
rect 31 59 269 5941
<< poly >>
rect -700 6300 1000 6800
rect -700 6000 -200 6300
rect 500 6000 1000 6300
rect -400 0 -200 6000
rect 500 0 700 6000
rect -700 -300 -200 0
rect 500 -300 1000 0
rect -700 -459 1000 -300
rect -700 -493 -180 -459
rect -146 -493 -106 -459
rect -72 -493 -32 -459
rect 2 -493 42 -459
rect 76 -493 116 -459
rect 150 -493 190 -459
rect 224 -493 264 -459
rect 298 -493 338 -459
rect 372 -493 412 -459
rect 446 -493 486 -459
rect 520 -493 1000 -459
rect -700 -533 1000 -493
rect -700 -567 -180 -533
rect -146 -567 -106 -533
rect -72 -567 -32 -533
rect 2 -567 42 -533
rect 76 -567 116 -533
rect 150 -567 190 -533
rect 224 -567 264 -533
rect 298 -567 338 -533
rect 372 -567 412 -533
rect 446 -567 486 -533
rect 520 -567 1000 -533
rect -700 -607 1000 -567
rect -700 -641 -180 -607
rect -146 -641 -106 -607
rect -72 -641 -32 -607
rect 2 -641 42 -607
rect 76 -641 116 -607
rect 150 -641 190 -607
rect 224 -641 264 -607
rect 298 -641 338 -607
rect 372 -641 412 -607
rect 446 -641 486 -607
rect 520 -641 1000 -607
rect -700 -800 1000 -641
<< polycont >>
rect -180 -493 -146 -459
rect -106 -493 -72 -459
rect -32 -493 2 -459
rect 42 -493 76 -459
rect 116 -493 150 -459
rect 190 -493 224 -459
rect 264 -493 298 -459
rect 338 -493 372 -459
rect 412 -493 446 -459
rect 486 -493 520 -459
rect -180 -567 -146 -533
rect -106 -567 -72 -533
rect -32 -567 2 -533
rect 42 -567 76 -533
rect 116 -567 150 -533
rect 190 -567 224 -533
rect 264 -567 298 -533
rect 338 -567 372 -533
rect 412 -567 446 -533
rect 486 -567 520 -533
rect -180 -641 -146 -607
rect -106 -641 -72 -607
rect -32 -641 2 -607
rect 42 -641 76 -607
rect 116 -641 150 -607
rect 190 -641 224 -607
rect 264 -641 298 -607
rect 338 -641 372 -607
rect 412 -641 446 -607
rect 486 -641 520 -607
<< locali >>
rect -3058 7959 3358 7983
rect -3058 7925 -2927 7959
rect -2893 7925 -2859 7959
rect -2821 7925 -2791 7959
rect -2749 7925 -2723 7959
rect -2677 7925 -2655 7959
rect -2605 7925 -2587 7959
rect -2533 7925 -2519 7959
rect -2461 7925 -2451 7959
rect -2389 7925 -2383 7959
rect -2317 7925 -2315 7959
rect -2281 7925 -2279 7959
rect -2213 7925 -2207 7959
rect -2145 7925 -2135 7959
rect -2077 7925 -2063 7959
rect -2009 7925 -1991 7959
rect -1941 7925 -1919 7959
rect -1873 7925 -1847 7959
rect -1805 7925 -1775 7959
rect -1737 7925 -1703 7959
rect -1669 7925 -1635 7959
rect -1597 7925 -1567 7959
rect -1525 7925 -1499 7959
rect -1453 7925 -1431 7959
rect -1381 7925 -1363 7959
rect -1309 7925 -1295 7959
rect -1237 7925 -1227 7959
rect -1165 7925 -1159 7959
rect -1093 7925 -1091 7959
rect -1057 7925 -1055 7959
rect -989 7925 -983 7959
rect -921 7925 -911 7959
rect -853 7925 -839 7959
rect -785 7925 -767 7959
rect -717 7925 -695 7959
rect -649 7925 -623 7959
rect -581 7925 -551 7959
rect -513 7925 -479 7959
rect -445 7925 -411 7959
rect -373 7925 -343 7959
rect -301 7925 -275 7959
rect -229 7925 -207 7959
rect -157 7925 -139 7959
rect -85 7925 -71 7959
rect -13 7925 -3 7959
rect 59 7925 65 7959
rect 131 7925 133 7959
rect 167 7925 169 7959
rect 235 7925 241 7959
rect 303 7925 313 7959
rect 371 7925 385 7959
rect 439 7925 457 7959
rect 507 7925 529 7959
rect 575 7925 601 7959
rect 643 7925 673 7959
rect 711 7925 745 7959
rect 779 7925 813 7959
rect 851 7925 881 7959
rect 923 7925 949 7959
rect 995 7925 1017 7959
rect 1067 7925 1085 7959
rect 1139 7925 1153 7959
rect 1211 7925 1221 7959
rect 1283 7925 1289 7959
rect 1355 7925 1357 7959
rect 1391 7925 1393 7959
rect 1459 7925 1465 7959
rect 1527 7925 1537 7959
rect 1595 7925 1609 7959
rect 1663 7925 1681 7959
rect 1731 7925 1753 7959
rect 1799 7925 1825 7959
rect 1867 7925 1897 7959
rect 1935 7925 1969 7959
rect 2003 7925 2037 7959
rect 2075 7925 2105 7959
rect 2147 7925 2173 7959
rect 2219 7925 2241 7959
rect 2291 7925 2309 7959
rect 2363 7925 2377 7959
rect 2435 7925 2445 7959
rect 2507 7925 2513 7959
rect 2579 7925 2581 7959
rect 2615 7925 2617 7959
rect 2683 7925 2689 7959
rect 2751 7925 2761 7959
rect 2819 7925 2833 7959
rect 2887 7925 2905 7959
rect 2955 7925 2977 7959
rect 3023 7925 3049 7959
rect 3091 7925 3121 7959
rect 3159 7925 3193 7959
rect 3227 7925 3358 7959
rect -3058 7901 3358 7925
rect -3058 7877 -2976 7901
rect -3058 7843 -3034 7877
rect -3000 7843 -2976 7877
rect -3058 7812 -2976 7843
rect -3058 7771 -3034 7812
rect -3000 7771 -2976 7812
rect -3058 7744 -2976 7771
rect -3058 7699 -3034 7744
rect -3000 7699 -2976 7744
rect -3058 7676 -2976 7699
rect -3058 7627 -3034 7676
rect -3000 7627 -2976 7676
rect -3058 7608 -2976 7627
rect -3058 7555 -3034 7608
rect -3000 7555 -2976 7608
rect -3058 7540 -2976 7555
rect -3058 7483 -3034 7540
rect -3000 7483 -2976 7540
rect -3058 7472 -2976 7483
rect -3058 7411 -3034 7472
rect -3000 7411 -2976 7472
rect -3058 7404 -2976 7411
rect -3058 7339 -3034 7404
rect -3000 7339 -2976 7404
rect -3058 7336 -2976 7339
rect -3058 7302 -3034 7336
rect -3000 7302 -2976 7336
rect -3058 7301 -2976 7302
rect -3058 7234 -3034 7301
rect -3000 7234 -2976 7301
rect -3058 7229 -2976 7234
rect -3058 7166 -3034 7229
rect -3000 7166 -2976 7229
rect -3058 7157 -2976 7166
rect -3058 7098 -3034 7157
rect -3000 7098 -2976 7157
rect -3058 7085 -2976 7098
rect -3058 7030 -3034 7085
rect -3000 7030 -2976 7085
rect -3058 7013 -2976 7030
rect -3058 6962 -3034 7013
rect -3000 6962 -2976 7013
rect -3058 6941 -2976 6962
rect -3058 6894 -3034 6941
rect -3000 6894 -2976 6941
rect -3058 6869 -2976 6894
rect -3058 6826 -3034 6869
rect -3000 6826 -2976 6869
rect -3058 6797 -2976 6826
rect -3058 6758 -3034 6797
rect -3000 6758 -2976 6797
rect -3058 6725 -2976 6758
rect -3058 6690 -3034 6725
rect -3000 6690 -2976 6725
rect -3058 6656 -2976 6690
rect -3058 6619 -3034 6656
rect -3000 6619 -2976 6656
rect -3058 6588 -2976 6619
rect -3058 6547 -3034 6588
rect -3000 6547 -2976 6588
rect -3058 6520 -2976 6547
rect -3058 6475 -3034 6520
rect -3000 6475 -2976 6520
rect -3058 6452 -2976 6475
rect -3058 6403 -3034 6452
rect -3000 6403 -2976 6452
rect -3058 6384 -2976 6403
rect -3058 6331 -3034 6384
rect -3000 6331 -2976 6384
rect -3058 6316 -2976 6331
rect -3058 6259 -3034 6316
rect -3000 6259 -2976 6316
rect -3058 6248 -2976 6259
rect -3058 6187 -3034 6248
rect -3000 6187 -2976 6248
rect -3058 6180 -2976 6187
rect -3058 6115 -3034 6180
rect -3000 6115 -2976 6180
rect -3058 6112 -2976 6115
rect -3058 6078 -3034 6112
rect -3000 6078 -2976 6112
rect -3058 6077 -2976 6078
rect -3058 6010 -3034 6077
rect -3000 6010 -2976 6077
rect -3058 6005 -2976 6010
rect -3058 5942 -3034 6005
rect -3000 5942 -2976 6005
rect 3276 7877 3358 7901
rect 3276 7843 3300 7877
rect 3334 7843 3358 7877
rect 3276 7812 3358 7843
rect 3276 7771 3300 7812
rect 3334 7771 3358 7812
rect 3276 7744 3358 7771
rect 3276 7699 3300 7744
rect 3334 7699 3358 7744
rect 3276 7676 3358 7699
rect 3276 7627 3300 7676
rect 3334 7627 3358 7676
rect 3276 7608 3358 7627
rect 3276 7555 3300 7608
rect 3334 7555 3358 7608
rect 3276 7540 3358 7555
rect 3276 7483 3300 7540
rect 3334 7483 3358 7540
rect 3276 7472 3358 7483
rect 3276 7411 3300 7472
rect 3334 7411 3358 7472
rect 3276 7404 3358 7411
rect 3276 7339 3300 7404
rect 3334 7339 3358 7404
rect 3276 7336 3358 7339
rect 3276 7302 3300 7336
rect 3334 7302 3358 7336
rect 3276 7301 3358 7302
rect 3276 7234 3300 7301
rect 3334 7234 3358 7301
rect 3276 7229 3358 7234
rect 3276 7166 3300 7229
rect 3334 7166 3358 7229
rect 3276 7157 3358 7166
rect 3276 7098 3300 7157
rect 3334 7098 3358 7157
rect 3276 7085 3358 7098
rect 3276 7030 3300 7085
rect 3334 7030 3358 7085
rect 3276 7013 3358 7030
rect 3276 6962 3300 7013
rect 3334 6962 3358 7013
rect 3276 6941 3358 6962
rect 3276 6894 3300 6941
rect 3334 6894 3358 6941
rect 3276 6869 3358 6894
rect 3276 6826 3300 6869
rect 3334 6826 3358 6869
rect 3276 6797 3358 6826
rect 3276 6758 3300 6797
rect 3334 6758 3358 6797
rect 3276 6725 3358 6758
rect 3276 6690 3300 6725
rect 3334 6690 3358 6725
rect 3276 6656 3358 6690
rect 3276 6619 3300 6656
rect 3334 6619 3358 6656
rect 3276 6588 3358 6619
rect 3276 6547 3300 6588
rect 3334 6547 3358 6588
rect 3276 6520 3358 6547
rect 3276 6475 3300 6520
rect 3334 6475 3358 6520
rect 3276 6452 3358 6475
rect 3276 6403 3300 6452
rect 3334 6403 3358 6452
rect 3276 6384 3358 6403
rect 3276 6331 3300 6384
rect 3334 6331 3358 6384
rect 3276 6316 3358 6331
rect 3276 6259 3300 6316
rect 3334 6259 3358 6316
rect 3276 6248 3358 6259
rect 3276 6187 3300 6248
rect 3334 6187 3358 6248
rect 3276 6180 3358 6187
rect 3276 6115 3300 6180
rect 3334 6115 3358 6180
rect 3276 6112 3358 6115
rect 3276 6078 3300 6112
rect 3334 6078 3358 6112
rect 3276 6077 3358 6078
rect 3276 6010 3300 6077
rect 3334 6010 3358 6077
rect 3276 6005 3358 6010
rect -3058 5933 -2976 5942
rect -3058 5874 -3034 5933
rect -3000 5874 -2976 5933
rect -3058 5861 -2976 5874
rect -3058 5806 -3034 5861
rect -3000 5806 -2976 5861
rect -3058 5789 -2976 5806
rect -3058 5738 -3034 5789
rect -3000 5738 -2976 5789
rect -3058 5717 -2976 5738
rect -3058 5670 -3034 5717
rect -3000 5670 -2976 5717
rect -3058 5645 -2976 5670
rect -3058 5602 -3034 5645
rect -3000 5602 -2976 5645
rect -3058 5573 -2976 5602
rect -3058 5534 -3034 5573
rect -3000 5534 -2976 5573
rect -3058 5501 -2976 5534
rect -3058 5466 -3034 5501
rect -3000 5466 -2976 5501
rect -3058 5432 -2976 5466
rect -3058 5395 -3034 5432
rect -3000 5395 -2976 5432
rect -3058 5364 -2976 5395
rect -3058 5323 -3034 5364
rect -3000 5323 -2976 5364
rect -3058 5296 -2976 5323
rect -3058 5251 -3034 5296
rect -3000 5251 -2976 5296
rect -3058 5228 -2976 5251
rect -3058 5179 -3034 5228
rect -3000 5179 -2976 5228
rect -3058 5160 -2976 5179
rect -3058 5107 -3034 5160
rect -3000 5107 -2976 5160
rect -3058 5092 -2976 5107
rect -3058 5035 -3034 5092
rect -3000 5035 -2976 5092
rect -3058 5024 -2976 5035
rect -3058 4963 -3034 5024
rect -3000 4963 -2976 5024
rect -3058 4956 -2976 4963
rect -3058 4891 -3034 4956
rect -3000 4891 -2976 4956
rect -3058 4888 -2976 4891
rect -3058 4854 -3034 4888
rect -3000 4854 -2976 4888
rect -3058 4853 -2976 4854
rect -3058 4786 -3034 4853
rect -3000 4786 -2976 4853
rect -3058 4781 -2976 4786
rect -3058 4718 -3034 4781
rect -3000 4718 -2976 4781
rect -3058 4709 -2976 4718
rect -3058 4650 -3034 4709
rect -3000 4650 -2976 4709
rect -3058 4637 -2976 4650
rect -3058 4582 -3034 4637
rect -3000 4582 -2976 4637
rect -3058 4565 -2976 4582
rect -3058 4514 -3034 4565
rect -3000 4514 -2976 4565
rect -3058 4493 -2976 4514
rect -3058 4446 -3034 4493
rect -3000 4446 -2976 4493
rect -3058 4421 -2976 4446
rect -3058 4378 -3034 4421
rect -3000 4378 -2976 4421
rect -3058 4349 -2976 4378
rect -3058 4310 -3034 4349
rect -3000 4310 -2976 4349
rect -3058 4277 -2976 4310
rect -3058 4242 -3034 4277
rect -3000 4242 -2976 4277
rect -3058 4208 -2976 4242
rect -3058 4171 -3034 4208
rect -3000 4171 -2976 4208
rect -3058 4140 -2976 4171
rect -3058 4099 -3034 4140
rect -3000 4099 -2976 4140
rect -3058 4072 -2976 4099
rect -3058 4027 -3034 4072
rect -3000 4027 -2976 4072
rect -3058 4004 -2976 4027
rect -3058 3955 -3034 4004
rect -3000 3955 -2976 4004
rect -3058 3936 -2976 3955
rect -3058 3883 -3034 3936
rect -3000 3883 -2976 3936
rect -3058 3868 -2976 3883
rect -3058 3811 -3034 3868
rect -3000 3811 -2976 3868
rect -3058 3800 -2976 3811
rect -3058 3739 -3034 3800
rect -3000 3739 -2976 3800
rect -3058 3732 -2976 3739
rect -3058 3667 -3034 3732
rect -3000 3667 -2976 3732
rect -3058 3664 -2976 3667
rect -3058 3630 -3034 3664
rect -3000 3630 -2976 3664
rect -3058 3629 -2976 3630
rect -3058 3562 -3034 3629
rect -3000 3562 -2976 3629
rect -3058 3557 -2976 3562
rect -3058 3494 -3034 3557
rect -3000 3494 -2976 3557
rect -3058 3485 -2976 3494
rect -3058 3426 -3034 3485
rect -3000 3426 -2976 3485
rect -3058 3413 -2976 3426
rect -3058 3358 -3034 3413
rect -3000 3358 -2976 3413
rect -3058 3341 -2976 3358
rect -3058 3290 -3034 3341
rect -3000 3290 -2976 3341
rect -3058 3269 -2976 3290
rect -3058 3222 -3034 3269
rect -3000 3222 -2976 3269
rect -3058 3197 -2976 3222
rect -3058 3154 -3034 3197
rect -3000 3154 -2976 3197
rect -3058 3125 -2976 3154
rect -3058 3086 -3034 3125
rect -3000 3086 -2976 3125
rect -3058 3053 -2976 3086
rect -3058 3018 -3034 3053
rect -3000 3018 -2976 3053
rect -3058 2984 -2976 3018
rect -3058 2947 -3034 2984
rect -3000 2947 -2976 2984
rect -3058 2916 -2976 2947
rect -3058 2875 -3034 2916
rect -3000 2875 -2976 2916
rect -3058 2848 -2976 2875
rect -3058 2803 -3034 2848
rect -3000 2803 -2976 2848
rect -3058 2780 -2976 2803
rect -3058 2731 -3034 2780
rect -3000 2731 -2976 2780
rect -3058 2712 -2976 2731
rect -3058 2659 -3034 2712
rect -3000 2659 -2976 2712
rect -3058 2644 -2976 2659
rect -3058 2587 -3034 2644
rect -3000 2587 -2976 2644
rect -3058 2576 -2976 2587
rect -3058 2515 -3034 2576
rect -3000 2515 -2976 2576
rect -3058 2508 -2976 2515
rect -3058 2443 -3034 2508
rect -3000 2443 -2976 2508
rect -3058 2440 -2976 2443
rect -3058 2406 -3034 2440
rect -3000 2406 -2976 2440
rect -3058 2405 -2976 2406
rect -3058 2338 -3034 2405
rect -3000 2338 -2976 2405
rect -3058 2333 -2976 2338
rect -3058 2270 -3034 2333
rect -3000 2270 -2976 2333
rect -3058 2261 -2976 2270
rect -3058 2202 -3034 2261
rect -3000 2202 -2976 2261
rect -3058 2189 -2976 2202
rect -3058 2134 -3034 2189
rect -3000 2134 -2976 2189
rect -3058 2117 -2976 2134
rect -3058 2066 -3034 2117
rect -3000 2066 -2976 2117
rect -3058 2045 -2976 2066
rect -3058 1998 -3034 2045
rect -3000 1998 -2976 2045
rect -3058 1973 -2976 1998
rect -3058 1930 -3034 1973
rect -3000 1930 -2976 1973
rect -3058 1901 -2976 1930
rect -3058 1862 -3034 1901
rect -3000 1862 -2976 1901
rect -3058 1829 -2976 1862
rect -3058 1794 -3034 1829
rect -3000 1794 -2976 1829
rect -3058 1760 -2976 1794
rect -3058 1723 -3034 1760
rect -3000 1723 -2976 1760
rect -3058 1692 -2976 1723
rect -3058 1651 -3034 1692
rect -3000 1651 -2976 1692
rect -3058 1624 -2976 1651
rect -3058 1579 -3034 1624
rect -3000 1579 -2976 1624
rect -3058 1556 -2976 1579
rect -3058 1507 -3034 1556
rect -3000 1507 -2976 1556
rect -3058 1488 -2976 1507
rect -3058 1435 -3034 1488
rect -3000 1435 -2976 1488
rect -3058 1420 -2976 1435
rect -3058 1363 -3034 1420
rect -3000 1363 -2976 1420
rect -3058 1352 -2976 1363
rect -3058 1291 -3034 1352
rect -3000 1291 -2976 1352
rect -3058 1284 -2976 1291
rect -3058 1219 -3034 1284
rect -3000 1219 -2976 1284
rect -3058 1216 -2976 1219
rect -3058 1182 -3034 1216
rect -3000 1182 -2976 1216
rect -3058 1181 -2976 1182
rect -3058 1114 -3034 1181
rect -3000 1114 -2976 1181
rect -3058 1109 -2976 1114
rect -3058 1046 -3034 1109
rect -3000 1046 -2976 1109
rect -3058 1037 -2976 1046
rect -3058 978 -3034 1037
rect -3000 978 -2976 1037
rect -3058 965 -2976 978
rect -3058 910 -3034 965
rect -3000 910 -2976 965
rect -3058 893 -2976 910
rect -3058 842 -3034 893
rect -3000 842 -2976 893
rect -3058 821 -2976 842
rect -3058 774 -3034 821
rect -3000 774 -2976 821
rect -3058 749 -2976 774
rect -3058 706 -3034 749
rect -3000 706 -2976 749
rect -3058 677 -2976 706
rect -3058 638 -3034 677
rect -3000 638 -2976 677
rect -3058 605 -2976 638
rect -3058 570 -3034 605
rect -3000 570 -2976 605
rect -3058 536 -2976 570
rect -3058 499 -3034 536
rect -3000 499 -2976 536
rect -3058 468 -2976 499
rect -3058 427 -3034 468
rect -3000 427 -2976 468
rect -3058 400 -2976 427
rect -3058 355 -3034 400
rect -3000 355 -2976 400
rect -3058 332 -2976 355
rect -3058 283 -3034 332
rect -3000 283 -2976 332
rect -3058 264 -2976 283
rect -3058 211 -3034 264
rect -3000 211 -2976 264
rect -3058 196 -2976 211
rect -3058 139 -3034 196
rect -3000 139 -2976 196
rect -3058 128 -2976 139
rect -3058 67 -3034 128
rect -3000 67 -2976 128
rect -3058 60 -2976 67
rect -3058 -5 -3034 60
rect -3000 -5 -2976 60
rect -1068 5975 -934 5991
rect -1068 5969 -1052 5975
rect -950 5969 -934 5975
rect -1068 31 -1054 5969
rect -948 31 -934 5969
rect -1068 25 -1052 31
rect -950 25 -934 31
rect -1068 9 -934 25
rect -830 5975 -696 5991
rect -830 5969 -814 5975
rect -712 5969 -696 5975
rect -830 31 -816 5969
rect -710 31 -696 5969
rect 996 5975 1130 5991
rect 996 5969 1012 5975
rect 1114 5969 1130 5975
rect 15 5941 285 5957
rect 15 5933 31 5941
rect 269 5933 285 5941
rect 15 67 25 5933
rect 275 67 285 5933
rect 15 59 31 67
rect 269 59 285 67
rect 15 43 285 59
rect -830 25 -814 31
rect -712 25 -696 31
rect -830 9 -696 25
rect 996 31 1010 5969
rect 1116 31 1130 5969
rect 996 25 1012 31
rect 1114 25 1130 31
rect 996 9 1130 25
rect 1234 5975 1368 5991
rect 1234 5969 1250 5975
rect 1352 5969 1368 5975
rect 1234 31 1248 5969
rect 1354 31 1368 5969
rect 1234 25 1250 31
rect 1352 25 1368 31
rect 1234 9 1368 25
rect 3276 5942 3300 6005
rect 3334 5942 3358 6005
rect 3276 5933 3358 5942
rect 3276 5874 3300 5933
rect 3334 5874 3358 5933
rect 3276 5861 3358 5874
rect 3276 5806 3300 5861
rect 3334 5806 3358 5861
rect 3276 5789 3358 5806
rect 3276 5738 3300 5789
rect 3334 5738 3358 5789
rect 3276 5717 3358 5738
rect 3276 5670 3300 5717
rect 3334 5670 3358 5717
rect 3276 5645 3358 5670
rect 3276 5602 3300 5645
rect 3334 5602 3358 5645
rect 3276 5573 3358 5602
rect 3276 5534 3300 5573
rect 3334 5534 3358 5573
rect 3276 5501 3358 5534
rect 3276 5466 3300 5501
rect 3334 5466 3358 5501
rect 3276 5432 3358 5466
rect 3276 5395 3300 5432
rect 3334 5395 3358 5432
rect 3276 5364 3358 5395
rect 3276 5323 3300 5364
rect 3334 5323 3358 5364
rect 3276 5296 3358 5323
rect 3276 5251 3300 5296
rect 3334 5251 3358 5296
rect 3276 5228 3358 5251
rect 3276 5179 3300 5228
rect 3334 5179 3358 5228
rect 3276 5160 3358 5179
rect 3276 5107 3300 5160
rect 3334 5107 3358 5160
rect 3276 5092 3358 5107
rect 3276 5035 3300 5092
rect 3334 5035 3358 5092
rect 3276 5024 3358 5035
rect 3276 4963 3300 5024
rect 3334 4963 3358 5024
rect 3276 4956 3358 4963
rect 3276 4891 3300 4956
rect 3334 4891 3358 4956
rect 3276 4888 3358 4891
rect 3276 4854 3300 4888
rect 3334 4854 3358 4888
rect 3276 4853 3358 4854
rect 3276 4786 3300 4853
rect 3334 4786 3358 4853
rect 3276 4781 3358 4786
rect 3276 4718 3300 4781
rect 3334 4718 3358 4781
rect 3276 4709 3358 4718
rect 3276 4650 3300 4709
rect 3334 4650 3358 4709
rect 3276 4637 3358 4650
rect 3276 4582 3300 4637
rect 3334 4582 3358 4637
rect 3276 4565 3358 4582
rect 3276 4514 3300 4565
rect 3334 4514 3358 4565
rect 3276 4493 3358 4514
rect 3276 4446 3300 4493
rect 3334 4446 3358 4493
rect 3276 4421 3358 4446
rect 3276 4378 3300 4421
rect 3334 4378 3358 4421
rect 3276 4349 3358 4378
rect 3276 4310 3300 4349
rect 3334 4310 3358 4349
rect 3276 4277 3358 4310
rect 3276 4242 3300 4277
rect 3334 4242 3358 4277
rect 3276 4208 3358 4242
rect 3276 4171 3300 4208
rect 3334 4171 3358 4208
rect 3276 4140 3358 4171
rect 3276 4099 3300 4140
rect 3334 4099 3358 4140
rect 3276 4072 3358 4099
rect 3276 4027 3300 4072
rect 3334 4027 3358 4072
rect 3276 4004 3358 4027
rect 3276 3955 3300 4004
rect 3334 3955 3358 4004
rect 3276 3936 3358 3955
rect 3276 3883 3300 3936
rect 3334 3883 3358 3936
rect 3276 3868 3358 3883
rect 3276 3811 3300 3868
rect 3334 3811 3358 3868
rect 3276 3800 3358 3811
rect 3276 3739 3300 3800
rect 3334 3739 3358 3800
rect 3276 3732 3358 3739
rect 3276 3667 3300 3732
rect 3334 3667 3358 3732
rect 3276 3664 3358 3667
rect 3276 3630 3300 3664
rect 3334 3630 3358 3664
rect 3276 3629 3358 3630
rect 3276 3562 3300 3629
rect 3334 3562 3358 3629
rect 3276 3557 3358 3562
rect 3276 3494 3300 3557
rect 3334 3494 3358 3557
rect 3276 3485 3358 3494
rect 3276 3426 3300 3485
rect 3334 3426 3358 3485
rect 3276 3413 3358 3426
rect 3276 3358 3300 3413
rect 3334 3358 3358 3413
rect 3276 3341 3358 3358
rect 3276 3290 3300 3341
rect 3334 3290 3358 3341
rect 3276 3269 3358 3290
rect 3276 3222 3300 3269
rect 3334 3222 3358 3269
rect 3276 3197 3358 3222
rect 3276 3154 3300 3197
rect 3334 3154 3358 3197
rect 3276 3125 3358 3154
rect 3276 3086 3300 3125
rect 3334 3086 3358 3125
rect 3276 3053 3358 3086
rect 3276 3018 3300 3053
rect 3334 3018 3358 3053
rect 3276 2984 3358 3018
rect 3276 2947 3300 2984
rect 3334 2947 3358 2984
rect 3276 2916 3358 2947
rect 3276 2875 3300 2916
rect 3334 2875 3358 2916
rect 3276 2848 3358 2875
rect 3276 2803 3300 2848
rect 3334 2803 3358 2848
rect 3276 2780 3358 2803
rect 3276 2731 3300 2780
rect 3334 2731 3358 2780
rect 3276 2712 3358 2731
rect 3276 2659 3300 2712
rect 3334 2659 3358 2712
rect 3276 2644 3358 2659
rect 3276 2587 3300 2644
rect 3334 2587 3358 2644
rect 3276 2576 3358 2587
rect 3276 2515 3300 2576
rect 3334 2515 3358 2576
rect 3276 2508 3358 2515
rect 3276 2443 3300 2508
rect 3334 2443 3358 2508
rect 3276 2440 3358 2443
rect 3276 2406 3300 2440
rect 3334 2406 3358 2440
rect 3276 2405 3358 2406
rect 3276 2338 3300 2405
rect 3334 2338 3358 2405
rect 3276 2333 3358 2338
rect 3276 2270 3300 2333
rect 3334 2270 3358 2333
rect 3276 2261 3358 2270
rect 3276 2202 3300 2261
rect 3334 2202 3358 2261
rect 3276 2189 3358 2202
rect 3276 2134 3300 2189
rect 3334 2134 3358 2189
rect 3276 2117 3358 2134
rect 3276 2066 3300 2117
rect 3334 2066 3358 2117
rect 3276 2045 3358 2066
rect 3276 1998 3300 2045
rect 3334 1998 3358 2045
rect 3276 1973 3358 1998
rect 3276 1930 3300 1973
rect 3334 1930 3358 1973
rect 3276 1901 3358 1930
rect 3276 1862 3300 1901
rect 3334 1862 3358 1901
rect 3276 1829 3358 1862
rect 3276 1794 3300 1829
rect 3334 1794 3358 1829
rect 3276 1760 3358 1794
rect 3276 1723 3300 1760
rect 3334 1723 3358 1760
rect 3276 1692 3358 1723
rect 3276 1651 3300 1692
rect 3334 1651 3358 1692
rect 3276 1624 3358 1651
rect 3276 1579 3300 1624
rect 3334 1579 3358 1624
rect 3276 1556 3358 1579
rect 3276 1507 3300 1556
rect 3334 1507 3358 1556
rect 3276 1488 3358 1507
rect 3276 1435 3300 1488
rect 3334 1435 3358 1488
rect 3276 1420 3358 1435
rect 3276 1363 3300 1420
rect 3334 1363 3358 1420
rect 3276 1352 3358 1363
rect 3276 1291 3300 1352
rect 3334 1291 3358 1352
rect 3276 1284 3358 1291
rect 3276 1219 3300 1284
rect 3334 1219 3358 1284
rect 3276 1216 3358 1219
rect 3276 1182 3300 1216
rect 3334 1182 3358 1216
rect 3276 1181 3358 1182
rect 3276 1114 3300 1181
rect 3334 1114 3358 1181
rect 3276 1109 3358 1114
rect 3276 1046 3300 1109
rect 3334 1046 3358 1109
rect 3276 1037 3358 1046
rect 3276 978 3300 1037
rect 3334 978 3358 1037
rect 3276 965 3358 978
rect 3276 910 3300 965
rect 3334 910 3358 965
rect 3276 893 3358 910
rect 3276 842 3300 893
rect 3334 842 3358 893
rect 3276 821 3358 842
rect 3276 774 3300 821
rect 3334 774 3358 821
rect 3276 749 3358 774
rect 3276 706 3300 749
rect 3334 706 3358 749
rect 3276 677 3358 706
rect 3276 638 3300 677
rect 3334 638 3358 677
rect 3276 605 3358 638
rect 3276 570 3300 605
rect 3334 570 3358 605
rect 3276 536 3358 570
rect 3276 499 3300 536
rect 3334 499 3358 536
rect 3276 468 3358 499
rect 3276 427 3300 468
rect 3334 427 3358 468
rect 3276 400 3358 427
rect 3276 355 3300 400
rect 3334 355 3358 400
rect 3276 332 3358 355
rect 3276 283 3300 332
rect 3334 283 3358 332
rect 3276 264 3358 283
rect 3276 211 3300 264
rect 3334 211 3358 264
rect 3276 196 3358 211
rect 3276 139 3300 196
rect 3334 139 3358 196
rect 3276 128 3358 139
rect 3276 67 3300 128
rect 3334 67 3358 128
rect 3276 60 3358 67
rect -3058 -8 -2976 -5
rect -3058 -42 -3034 -8
rect -3000 -42 -2976 -8
rect -3058 -43 -2976 -42
rect -3058 -110 -3034 -43
rect -3000 -110 -2976 -43
rect -3058 -115 -2976 -110
rect -3058 -178 -3034 -115
rect -3000 -178 -2976 -115
rect -3058 -187 -2976 -178
rect -3058 -246 -3034 -187
rect -3000 -246 -2976 -187
rect -3058 -259 -2976 -246
rect -3058 -314 -3034 -259
rect -3000 -314 -2976 -259
rect -3058 -331 -2976 -314
rect -3058 -382 -3034 -331
rect -3000 -382 -2976 -331
rect -3058 -403 -2976 -382
rect -3058 -450 -3034 -403
rect -3000 -450 -2976 -403
rect 3276 -5 3300 60
rect 3334 -5 3358 60
rect 3276 -8 3358 -5
rect 3276 -42 3300 -8
rect 3334 -42 3358 -8
rect 3276 -43 3358 -42
rect 3276 -110 3300 -43
rect 3334 -110 3358 -43
rect 3276 -115 3358 -110
rect 3276 -178 3300 -115
rect 3334 -178 3358 -115
rect 3276 -187 3358 -178
rect 3276 -246 3300 -187
rect 3334 -246 3358 -187
rect 3276 -259 3358 -246
rect 3276 -314 3300 -259
rect 3334 -314 3358 -259
rect 3276 -331 3358 -314
rect 3276 -382 3300 -331
rect 3334 -382 3358 -331
rect 3276 -403 3358 -382
rect -3058 -475 -2976 -450
rect -3058 -518 -3034 -475
rect -3000 -518 -2976 -475
rect -3058 -547 -2976 -518
rect -3058 -586 -3034 -547
rect -3000 -586 -2976 -547
rect -3058 -619 -2976 -586
rect -3058 -654 -3034 -619
rect -3000 -654 -2976 -619
rect -3058 -688 -2976 -654
rect -209 -459 555 -443
rect -209 -493 -180 -459
rect -146 -493 -106 -459
rect -72 -493 -32 -459
rect 2 -493 42 -459
rect 76 -493 116 -459
rect 150 -493 190 -459
rect 224 -493 264 -459
rect 298 -493 338 -459
rect 372 -493 412 -459
rect 446 -493 486 -459
rect 520 -493 555 -459
rect -209 -533 555 -493
rect -209 -567 -180 -533
rect -146 -567 -106 -533
rect -72 -567 -32 -533
rect 2 -567 42 -533
rect 76 -567 116 -533
rect 150 -567 190 -533
rect 224 -567 264 -533
rect 298 -567 338 -533
rect 372 -567 412 -533
rect 446 -567 486 -533
rect 520 -567 555 -533
rect -209 -607 555 -567
rect -209 -641 -180 -607
rect -146 -641 -106 -607
rect -72 -641 -32 -607
rect 2 -641 42 -607
rect 76 -641 116 -607
rect 150 -641 190 -607
rect 224 -641 264 -607
rect 298 -641 338 -607
rect 372 -641 412 -607
rect 446 -641 486 -607
rect 520 -641 555 -607
rect -209 -657 555 -641
rect 3276 -450 3300 -403
rect 3334 -450 3358 -403
rect 3276 -475 3358 -450
rect 3276 -518 3300 -475
rect 3334 -518 3358 -475
rect 3276 -547 3358 -518
rect 3276 -586 3300 -547
rect 3334 -586 3358 -547
rect 3276 -619 3358 -586
rect 3276 -654 3300 -619
rect 3334 -654 3358 -619
rect -3058 -725 -3034 -688
rect -3000 -725 -2976 -688
rect -3058 -756 -2976 -725
rect -3058 -797 -3034 -756
rect -3000 -797 -2976 -756
rect -3058 -824 -2976 -797
rect -3058 -869 -3034 -824
rect -3000 -869 -2976 -824
rect -3058 -892 -2976 -869
rect -3058 -941 -3034 -892
rect -3000 -941 -2976 -892
rect -3058 -960 -2976 -941
rect -3058 -1013 -3034 -960
rect -3000 -1013 -2976 -960
rect -3058 -1028 -2976 -1013
rect -3058 -1085 -3034 -1028
rect -3000 -1085 -2976 -1028
rect -3058 -1096 -2976 -1085
rect -3058 -1157 -3034 -1096
rect -3000 -1157 -2976 -1096
rect -3058 -1164 -2976 -1157
rect -3058 -1229 -3034 -1164
rect -3000 -1229 -2976 -1164
rect -3058 -1232 -2976 -1229
rect -3058 -1266 -3034 -1232
rect -3000 -1266 -2976 -1232
rect -3058 -1267 -2976 -1266
rect -3058 -1334 -3034 -1267
rect -3000 -1334 -2976 -1267
rect -3058 -1339 -2976 -1334
rect -3058 -1402 -3034 -1339
rect -3000 -1402 -2976 -1339
rect -3058 -1411 -2976 -1402
rect -3058 -1470 -3034 -1411
rect -3000 -1470 -2976 -1411
rect -3058 -1483 -2976 -1470
rect -3058 -1538 -3034 -1483
rect -3000 -1538 -2976 -1483
rect -3058 -1555 -2976 -1538
rect -3058 -1606 -3034 -1555
rect -3000 -1606 -2976 -1555
rect -3058 -1627 -2976 -1606
rect -3058 -1674 -3034 -1627
rect -3000 -1674 -2976 -1627
rect -3058 -1699 -2976 -1674
rect -3058 -1742 -3034 -1699
rect -3000 -1742 -2976 -1699
rect -3058 -1771 -2976 -1742
rect -3058 -1810 -3034 -1771
rect -3000 -1810 -2976 -1771
rect -3058 -1843 -2976 -1810
rect -3058 -1877 -3034 -1843
rect -3000 -1877 -2976 -1843
rect -3058 -1900 -2976 -1877
rect 3276 -688 3358 -654
rect 3276 -725 3300 -688
rect 3334 -725 3358 -688
rect 3276 -756 3358 -725
rect 3276 -797 3300 -756
rect 3334 -797 3358 -756
rect 3276 -824 3358 -797
rect 3276 -869 3300 -824
rect 3334 -869 3358 -824
rect 3276 -892 3358 -869
rect 3276 -941 3300 -892
rect 3334 -941 3358 -892
rect 3276 -960 3358 -941
rect 3276 -1013 3300 -960
rect 3334 -1013 3358 -960
rect 3276 -1028 3358 -1013
rect 3276 -1085 3300 -1028
rect 3334 -1085 3358 -1028
rect 3276 -1096 3358 -1085
rect 3276 -1157 3300 -1096
rect 3334 -1157 3358 -1096
rect 3276 -1164 3358 -1157
rect 3276 -1229 3300 -1164
rect 3334 -1229 3358 -1164
rect 3276 -1232 3358 -1229
rect 3276 -1266 3300 -1232
rect 3334 -1266 3358 -1232
rect 3276 -1267 3358 -1266
rect 3276 -1334 3300 -1267
rect 3334 -1334 3358 -1267
rect 3276 -1339 3358 -1334
rect 3276 -1402 3300 -1339
rect 3334 -1402 3358 -1339
rect 3276 -1411 3358 -1402
rect 3276 -1470 3300 -1411
rect 3334 -1470 3358 -1411
rect 3276 -1483 3358 -1470
rect 3276 -1538 3300 -1483
rect 3334 -1538 3358 -1483
rect 3276 -1555 3358 -1538
rect 3276 -1606 3300 -1555
rect 3334 -1606 3358 -1555
rect 3276 -1627 3358 -1606
rect 3276 -1674 3300 -1627
rect 3334 -1674 3358 -1627
rect 3276 -1699 3358 -1674
rect 3276 -1742 3300 -1699
rect 3334 -1742 3358 -1699
rect 3276 -1771 3358 -1742
rect 3276 -1810 3300 -1771
rect 3334 -1810 3358 -1771
rect 3276 -1843 3358 -1810
rect 3276 -1877 3300 -1843
rect 3334 -1877 3358 -1843
rect 3276 -1900 3358 -1877
rect -3058 -1924 3358 -1900
rect -3058 -1958 -2927 -1924
rect -2893 -1958 -2859 -1924
rect -2821 -1958 -2791 -1924
rect -2749 -1958 -2723 -1924
rect -2677 -1958 -2655 -1924
rect -2605 -1958 -2587 -1924
rect -2533 -1958 -2519 -1924
rect -2461 -1958 -2451 -1924
rect -2389 -1958 -2383 -1924
rect -2317 -1958 -2315 -1924
rect -2281 -1958 -2279 -1924
rect -2213 -1958 -2207 -1924
rect -2145 -1958 -2135 -1924
rect -2077 -1958 -2063 -1924
rect -2009 -1958 -1991 -1924
rect -1941 -1958 -1919 -1924
rect -1873 -1958 -1847 -1924
rect -1805 -1958 -1775 -1924
rect -1737 -1958 -1703 -1924
rect -1669 -1958 -1635 -1924
rect -1597 -1958 -1567 -1924
rect -1525 -1958 -1499 -1924
rect -1453 -1958 -1431 -1924
rect -1381 -1958 -1363 -1924
rect -1309 -1958 -1295 -1924
rect -1237 -1958 -1227 -1924
rect -1165 -1958 -1159 -1924
rect -1093 -1958 -1091 -1924
rect -1057 -1958 -1055 -1924
rect -989 -1958 -983 -1924
rect -921 -1958 -911 -1924
rect -853 -1958 -839 -1924
rect -785 -1958 -767 -1924
rect -717 -1958 -695 -1924
rect -649 -1958 -623 -1924
rect -581 -1958 -551 -1924
rect -513 -1958 -479 -1924
rect -445 -1958 -411 -1924
rect -373 -1958 -343 -1924
rect -301 -1958 -275 -1924
rect -229 -1958 -207 -1924
rect -157 -1958 -139 -1924
rect -85 -1958 -71 -1924
rect -13 -1958 -3 -1924
rect 59 -1958 65 -1924
rect 131 -1958 133 -1924
rect 167 -1958 169 -1924
rect 235 -1958 241 -1924
rect 303 -1958 313 -1924
rect 371 -1958 385 -1924
rect 439 -1958 457 -1924
rect 507 -1958 529 -1924
rect 575 -1958 601 -1924
rect 643 -1958 673 -1924
rect 711 -1958 745 -1924
rect 779 -1958 813 -1924
rect 851 -1958 881 -1924
rect 923 -1958 949 -1924
rect 995 -1958 1017 -1924
rect 1067 -1958 1085 -1924
rect 1139 -1958 1153 -1924
rect 1211 -1958 1221 -1924
rect 1283 -1958 1289 -1924
rect 1355 -1958 1357 -1924
rect 1391 -1958 1393 -1924
rect 1459 -1958 1465 -1924
rect 1527 -1958 1537 -1924
rect 1595 -1958 1609 -1924
rect 1663 -1958 1681 -1924
rect 1731 -1958 1753 -1924
rect 1799 -1958 1825 -1924
rect 1867 -1958 1897 -1924
rect 1935 -1958 1969 -1924
rect 2003 -1958 2037 -1924
rect 2075 -1958 2105 -1924
rect 2147 -1958 2173 -1924
rect 2219 -1958 2241 -1924
rect 2291 -1958 2309 -1924
rect 2363 -1958 2377 -1924
rect 2435 -1958 2445 -1924
rect 2507 -1958 2513 -1924
rect 2579 -1958 2581 -1924
rect 2615 -1958 2617 -1924
rect 2683 -1958 2689 -1924
rect 2751 -1958 2761 -1924
rect 2819 -1958 2833 -1924
rect 2887 -1958 2905 -1924
rect 2955 -1958 2977 -1924
rect 3023 -1958 3049 -1924
rect 3091 -1958 3121 -1924
rect 3159 -1958 3193 -1924
rect 3227 -1958 3358 -1924
rect -3058 -1982 3358 -1958
<< viali >>
rect -2927 7925 -2893 7959
rect -2855 7925 -2825 7959
rect -2825 7925 -2821 7959
rect -2783 7925 -2757 7959
rect -2757 7925 -2749 7959
rect -2711 7925 -2689 7959
rect -2689 7925 -2677 7959
rect -2639 7925 -2621 7959
rect -2621 7925 -2605 7959
rect -2567 7925 -2553 7959
rect -2553 7925 -2533 7959
rect -2495 7925 -2485 7959
rect -2485 7925 -2461 7959
rect -2423 7925 -2417 7959
rect -2417 7925 -2389 7959
rect -2351 7925 -2349 7959
rect -2349 7925 -2317 7959
rect -2279 7925 -2247 7959
rect -2247 7925 -2245 7959
rect -2207 7925 -2179 7959
rect -2179 7925 -2173 7959
rect -2135 7925 -2111 7959
rect -2111 7925 -2101 7959
rect -2063 7925 -2043 7959
rect -2043 7925 -2029 7959
rect -1991 7925 -1975 7959
rect -1975 7925 -1957 7959
rect -1919 7925 -1907 7959
rect -1907 7925 -1885 7959
rect -1847 7925 -1839 7959
rect -1839 7925 -1813 7959
rect -1775 7925 -1771 7959
rect -1771 7925 -1741 7959
rect -1703 7925 -1669 7959
rect -1631 7925 -1601 7959
rect -1601 7925 -1597 7959
rect -1559 7925 -1533 7959
rect -1533 7925 -1525 7959
rect -1487 7925 -1465 7959
rect -1465 7925 -1453 7959
rect -1415 7925 -1397 7959
rect -1397 7925 -1381 7959
rect -1343 7925 -1329 7959
rect -1329 7925 -1309 7959
rect -1271 7925 -1261 7959
rect -1261 7925 -1237 7959
rect -1199 7925 -1193 7959
rect -1193 7925 -1165 7959
rect -1127 7925 -1125 7959
rect -1125 7925 -1093 7959
rect -1055 7925 -1023 7959
rect -1023 7925 -1021 7959
rect -983 7925 -955 7959
rect -955 7925 -949 7959
rect -911 7925 -887 7959
rect -887 7925 -877 7959
rect -839 7925 -819 7959
rect -819 7925 -805 7959
rect -767 7925 -751 7959
rect -751 7925 -733 7959
rect -695 7925 -683 7959
rect -683 7925 -661 7959
rect -623 7925 -615 7959
rect -615 7925 -589 7959
rect -551 7925 -547 7959
rect -547 7925 -517 7959
rect -479 7925 -445 7959
rect -407 7925 -377 7959
rect -377 7925 -373 7959
rect -335 7925 -309 7959
rect -309 7925 -301 7959
rect -263 7925 -241 7959
rect -241 7925 -229 7959
rect -191 7925 -173 7959
rect -173 7925 -157 7959
rect -119 7925 -105 7959
rect -105 7925 -85 7959
rect -47 7925 -37 7959
rect -37 7925 -13 7959
rect 25 7925 31 7959
rect 31 7925 59 7959
rect 97 7925 99 7959
rect 99 7925 131 7959
rect 169 7925 201 7959
rect 201 7925 203 7959
rect 241 7925 269 7959
rect 269 7925 275 7959
rect 313 7925 337 7959
rect 337 7925 347 7959
rect 385 7925 405 7959
rect 405 7925 419 7959
rect 457 7925 473 7959
rect 473 7925 491 7959
rect 529 7925 541 7959
rect 541 7925 563 7959
rect 601 7925 609 7959
rect 609 7925 635 7959
rect 673 7925 677 7959
rect 677 7925 707 7959
rect 745 7925 779 7959
rect 817 7925 847 7959
rect 847 7925 851 7959
rect 889 7925 915 7959
rect 915 7925 923 7959
rect 961 7925 983 7959
rect 983 7925 995 7959
rect 1033 7925 1051 7959
rect 1051 7925 1067 7959
rect 1105 7925 1119 7959
rect 1119 7925 1139 7959
rect 1177 7925 1187 7959
rect 1187 7925 1211 7959
rect 1249 7925 1255 7959
rect 1255 7925 1283 7959
rect 1321 7925 1323 7959
rect 1323 7925 1355 7959
rect 1393 7925 1425 7959
rect 1425 7925 1427 7959
rect 1465 7925 1493 7959
rect 1493 7925 1499 7959
rect 1537 7925 1561 7959
rect 1561 7925 1571 7959
rect 1609 7925 1629 7959
rect 1629 7925 1643 7959
rect 1681 7925 1697 7959
rect 1697 7925 1715 7959
rect 1753 7925 1765 7959
rect 1765 7925 1787 7959
rect 1825 7925 1833 7959
rect 1833 7925 1859 7959
rect 1897 7925 1901 7959
rect 1901 7925 1931 7959
rect 1969 7925 2003 7959
rect 2041 7925 2071 7959
rect 2071 7925 2075 7959
rect 2113 7925 2139 7959
rect 2139 7925 2147 7959
rect 2185 7925 2207 7959
rect 2207 7925 2219 7959
rect 2257 7925 2275 7959
rect 2275 7925 2291 7959
rect 2329 7925 2343 7959
rect 2343 7925 2363 7959
rect 2401 7925 2411 7959
rect 2411 7925 2435 7959
rect 2473 7925 2479 7959
rect 2479 7925 2507 7959
rect 2545 7925 2547 7959
rect 2547 7925 2579 7959
rect 2617 7925 2649 7959
rect 2649 7925 2651 7959
rect 2689 7925 2717 7959
rect 2717 7925 2723 7959
rect 2761 7925 2785 7959
rect 2785 7925 2795 7959
rect 2833 7925 2853 7959
rect 2853 7925 2867 7959
rect 2905 7925 2921 7959
rect 2921 7925 2939 7959
rect 2977 7925 2989 7959
rect 2989 7925 3011 7959
rect 3049 7925 3057 7959
rect 3057 7925 3083 7959
rect 3121 7925 3125 7959
rect 3125 7925 3155 7959
rect 3193 7925 3227 7959
rect -3034 7843 -3000 7877
rect -3034 7778 -3000 7805
rect -3034 7771 -3000 7778
rect -3034 7710 -3000 7733
rect -3034 7699 -3000 7710
rect -3034 7642 -3000 7661
rect -3034 7627 -3000 7642
rect -3034 7574 -3000 7589
rect -3034 7555 -3000 7574
rect -3034 7506 -3000 7517
rect -3034 7483 -3000 7506
rect -3034 7438 -3000 7445
rect -3034 7411 -3000 7438
rect -3034 7370 -3000 7373
rect -3034 7339 -3000 7370
rect -3034 7268 -3000 7301
rect -3034 7267 -3000 7268
rect -3034 7200 -3000 7229
rect -3034 7195 -3000 7200
rect -3034 7132 -3000 7157
rect -3034 7123 -3000 7132
rect -3034 7064 -3000 7085
rect -3034 7051 -3000 7064
rect -3034 6996 -3000 7013
rect -3034 6979 -3000 6996
rect -3034 6928 -3000 6941
rect -3034 6907 -3000 6928
rect -3034 6860 -3000 6869
rect -3034 6835 -3000 6860
rect -3034 6792 -3000 6797
rect -3034 6763 -3000 6792
rect -3034 6724 -3000 6725
rect -3034 6691 -3000 6724
rect -3034 6622 -3000 6653
rect -3034 6619 -3000 6622
rect -3034 6554 -3000 6581
rect -3034 6547 -3000 6554
rect -3034 6486 -3000 6509
rect -3034 6475 -3000 6486
rect -3034 6418 -3000 6437
rect -3034 6403 -3000 6418
rect -3034 6350 -3000 6365
rect -3034 6331 -3000 6350
rect -3034 6282 -3000 6293
rect -3034 6259 -3000 6282
rect -3034 6214 -3000 6221
rect -3034 6187 -3000 6214
rect -3034 6146 -3000 6149
rect -3034 6115 -3000 6146
rect -3034 6044 -3000 6077
rect -3034 6043 -3000 6044
rect -3034 5976 -3000 6005
rect -3034 5971 -3000 5976
rect 3300 7843 3334 7877
rect 3300 7778 3334 7805
rect 3300 7771 3334 7778
rect 3300 7710 3334 7733
rect 3300 7699 3334 7710
rect 3300 7642 3334 7661
rect 3300 7627 3334 7642
rect 3300 7574 3334 7589
rect 3300 7555 3334 7574
rect 3300 7506 3334 7517
rect 3300 7483 3334 7506
rect 3300 7438 3334 7445
rect 3300 7411 3334 7438
rect 3300 7370 3334 7373
rect 3300 7339 3334 7370
rect 3300 7268 3334 7301
rect 3300 7267 3334 7268
rect 3300 7200 3334 7229
rect 3300 7195 3334 7200
rect 3300 7132 3334 7157
rect 3300 7123 3334 7132
rect 3300 7064 3334 7085
rect 3300 7051 3334 7064
rect 3300 6996 3334 7013
rect 3300 6979 3334 6996
rect 3300 6928 3334 6941
rect 3300 6907 3334 6928
rect 3300 6860 3334 6869
rect 3300 6835 3334 6860
rect 3300 6792 3334 6797
rect 3300 6763 3334 6792
rect 3300 6724 3334 6725
rect 3300 6691 3334 6724
rect 3300 6622 3334 6653
rect 3300 6619 3334 6622
rect 3300 6554 3334 6581
rect 3300 6547 3334 6554
rect 3300 6486 3334 6509
rect 3300 6475 3334 6486
rect 3300 6418 3334 6437
rect 3300 6403 3334 6418
rect 3300 6350 3334 6365
rect 3300 6331 3334 6350
rect 3300 6282 3334 6293
rect 3300 6259 3334 6282
rect 3300 6214 3334 6221
rect 3300 6187 3334 6214
rect 3300 6146 3334 6149
rect 3300 6115 3334 6146
rect 3300 6044 3334 6077
rect 3300 6043 3334 6044
rect -3034 5908 -3000 5933
rect -3034 5899 -3000 5908
rect -3034 5840 -3000 5861
rect -3034 5827 -3000 5840
rect -3034 5772 -3000 5789
rect -3034 5755 -3000 5772
rect -3034 5704 -3000 5717
rect -3034 5683 -3000 5704
rect -3034 5636 -3000 5645
rect -3034 5611 -3000 5636
rect -3034 5568 -3000 5573
rect -3034 5539 -3000 5568
rect -3034 5500 -3000 5501
rect -3034 5467 -3000 5500
rect -3034 5398 -3000 5429
rect -3034 5395 -3000 5398
rect -3034 5330 -3000 5357
rect -3034 5323 -3000 5330
rect -3034 5262 -3000 5285
rect -3034 5251 -3000 5262
rect -3034 5194 -3000 5213
rect -3034 5179 -3000 5194
rect -3034 5126 -3000 5141
rect -3034 5107 -3000 5126
rect -3034 5058 -3000 5069
rect -3034 5035 -3000 5058
rect -3034 4990 -3000 4997
rect -3034 4963 -3000 4990
rect -3034 4922 -3000 4925
rect -3034 4891 -3000 4922
rect -3034 4820 -3000 4853
rect -3034 4819 -3000 4820
rect -3034 4752 -3000 4781
rect -3034 4747 -3000 4752
rect -3034 4684 -3000 4709
rect -3034 4675 -3000 4684
rect -3034 4616 -3000 4637
rect -3034 4603 -3000 4616
rect -3034 4548 -3000 4565
rect -3034 4531 -3000 4548
rect -3034 4480 -3000 4493
rect -3034 4459 -3000 4480
rect -3034 4412 -3000 4421
rect -3034 4387 -3000 4412
rect -3034 4344 -3000 4349
rect -3034 4315 -3000 4344
rect -3034 4276 -3000 4277
rect -3034 4243 -3000 4276
rect -3034 4174 -3000 4205
rect -3034 4171 -3000 4174
rect -3034 4106 -3000 4133
rect -3034 4099 -3000 4106
rect -3034 4038 -3000 4061
rect -3034 4027 -3000 4038
rect -3034 3970 -3000 3989
rect -3034 3955 -3000 3970
rect -3034 3902 -3000 3917
rect -3034 3883 -3000 3902
rect -3034 3834 -3000 3845
rect -3034 3811 -3000 3834
rect -3034 3766 -3000 3773
rect -3034 3739 -3000 3766
rect -3034 3698 -3000 3701
rect -3034 3667 -3000 3698
rect -3034 3596 -3000 3629
rect -3034 3595 -3000 3596
rect -3034 3528 -3000 3557
rect -3034 3523 -3000 3528
rect -3034 3460 -3000 3485
rect -3034 3451 -3000 3460
rect -3034 3392 -3000 3413
rect -3034 3379 -3000 3392
rect -3034 3324 -3000 3341
rect -3034 3307 -3000 3324
rect -3034 3256 -3000 3269
rect -3034 3235 -3000 3256
rect -3034 3188 -3000 3197
rect -3034 3163 -3000 3188
rect -3034 3120 -3000 3125
rect -3034 3091 -3000 3120
rect -3034 3052 -3000 3053
rect -3034 3019 -3000 3052
rect -3034 2950 -3000 2981
rect -3034 2947 -3000 2950
rect -3034 2882 -3000 2909
rect -3034 2875 -3000 2882
rect -3034 2814 -3000 2837
rect -3034 2803 -3000 2814
rect -3034 2746 -3000 2765
rect -3034 2731 -3000 2746
rect -3034 2678 -3000 2693
rect -3034 2659 -3000 2678
rect -3034 2610 -3000 2621
rect -3034 2587 -3000 2610
rect -3034 2542 -3000 2549
rect -3034 2515 -3000 2542
rect -3034 2474 -3000 2477
rect -3034 2443 -3000 2474
rect -3034 2372 -3000 2405
rect -3034 2371 -3000 2372
rect -3034 2304 -3000 2333
rect -3034 2299 -3000 2304
rect -3034 2236 -3000 2261
rect -3034 2227 -3000 2236
rect -3034 2168 -3000 2189
rect -3034 2155 -3000 2168
rect -3034 2100 -3000 2117
rect -3034 2083 -3000 2100
rect -3034 2032 -3000 2045
rect -3034 2011 -3000 2032
rect -3034 1964 -3000 1973
rect -3034 1939 -3000 1964
rect -3034 1896 -3000 1901
rect -3034 1867 -3000 1896
rect -3034 1828 -3000 1829
rect -3034 1795 -3000 1828
rect -3034 1726 -3000 1757
rect -3034 1723 -3000 1726
rect -3034 1658 -3000 1685
rect -3034 1651 -3000 1658
rect -3034 1590 -3000 1613
rect -3034 1579 -3000 1590
rect -3034 1522 -3000 1541
rect -3034 1507 -3000 1522
rect -3034 1454 -3000 1469
rect -3034 1435 -3000 1454
rect -3034 1386 -3000 1397
rect -3034 1363 -3000 1386
rect -3034 1318 -3000 1325
rect -3034 1291 -3000 1318
rect -3034 1250 -3000 1253
rect -3034 1219 -3000 1250
rect -3034 1148 -3000 1181
rect -3034 1147 -3000 1148
rect -3034 1080 -3000 1109
rect -3034 1075 -3000 1080
rect -3034 1012 -3000 1037
rect -3034 1003 -3000 1012
rect -3034 944 -3000 965
rect -3034 931 -3000 944
rect -3034 876 -3000 893
rect -3034 859 -3000 876
rect -3034 808 -3000 821
rect -3034 787 -3000 808
rect -3034 740 -3000 749
rect -3034 715 -3000 740
rect -3034 672 -3000 677
rect -3034 643 -3000 672
rect -3034 604 -3000 605
rect -3034 571 -3000 604
rect -3034 502 -3000 533
rect -3034 499 -3000 502
rect -3034 434 -3000 461
rect -3034 427 -3000 434
rect -3034 366 -3000 389
rect -3034 355 -3000 366
rect -3034 298 -3000 317
rect -3034 283 -3000 298
rect -3034 230 -3000 245
rect -3034 211 -3000 230
rect -3034 162 -3000 173
rect -3034 139 -3000 162
rect -3034 94 -3000 101
rect -3034 67 -3000 94
rect -3034 26 -3000 29
rect -3034 -5 -3000 26
rect -1054 31 -1052 5969
rect -1052 31 -950 5969
rect -950 31 -948 5969
rect -816 31 -814 5969
rect -814 31 -712 5969
rect -712 31 -710 5969
rect 25 67 31 5933
rect 31 67 269 5933
rect 269 67 275 5933
rect 1010 31 1012 5969
rect 1012 31 1114 5969
rect 1114 31 1116 5969
rect 1248 31 1250 5969
rect 1250 31 1352 5969
rect 1352 31 1354 5969
rect 3300 5976 3334 6005
rect 3300 5971 3334 5976
rect 3300 5908 3334 5933
rect 3300 5899 3334 5908
rect 3300 5840 3334 5861
rect 3300 5827 3334 5840
rect 3300 5772 3334 5789
rect 3300 5755 3334 5772
rect 3300 5704 3334 5717
rect 3300 5683 3334 5704
rect 3300 5636 3334 5645
rect 3300 5611 3334 5636
rect 3300 5568 3334 5573
rect 3300 5539 3334 5568
rect 3300 5500 3334 5501
rect 3300 5467 3334 5500
rect 3300 5398 3334 5429
rect 3300 5395 3334 5398
rect 3300 5330 3334 5357
rect 3300 5323 3334 5330
rect 3300 5262 3334 5285
rect 3300 5251 3334 5262
rect 3300 5194 3334 5213
rect 3300 5179 3334 5194
rect 3300 5126 3334 5141
rect 3300 5107 3334 5126
rect 3300 5058 3334 5069
rect 3300 5035 3334 5058
rect 3300 4990 3334 4997
rect 3300 4963 3334 4990
rect 3300 4922 3334 4925
rect 3300 4891 3334 4922
rect 3300 4820 3334 4853
rect 3300 4819 3334 4820
rect 3300 4752 3334 4781
rect 3300 4747 3334 4752
rect 3300 4684 3334 4709
rect 3300 4675 3334 4684
rect 3300 4616 3334 4637
rect 3300 4603 3334 4616
rect 3300 4548 3334 4565
rect 3300 4531 3334 4548
rect 3300 4480 3334 4493
rect 3300 4459 3334 4480
rect 3300 4412 3334 4421
rect 3300 4387 3334 4412
rect 3300 4344 3334 4349
rect 3300 4315 3334 4344
rect 3300 4276 3334 4277
rect 3300 4243 3334 4276
rect 3300 4174 3334 4205
rect 3300 4171 3334 4174
rect 3300 4106 3334 4133
rect 3300 4099 3334 4106
rect 3300 4038 3334 4061
rect 3300 4027 3334 4038
rect 3300 3970 3334 3989
rect 3300 3955 3334 3970
rect 3300 3902 3334 3917
rect 3300 3883 3334 3902
rect 3300 3834 3334 3845
rect 3300 3811 3334 3834
rect 3300 3766 3334 3773
rect 3300 3739 3334 3766
rect 3300 3698 3334 3701
rect 3300 3667 3334 3698
rect 3300 3596 3334 3629
rect 3300 3595 3334 3596
rect 3300 3528 3334 3557
rect 3300 3523 3334 3528
rect 3300 3460 3334 3485
rect 3300 3451 3334 3460
rect 3300 3392 3334 3413
rect 3300 3379 3334 3392
rect 3300 3324 3334 3341
rect 3300 3307 3334 3324
rect 3300 3256 3334 3269
rect 3300 3235 3334 3256
rect 3300 3188 3334 3197
rect 3300 3163 3334 3188
rect 3300 3120 3334 3125
rect 3300 3091 3334 3120
rect 3300 3052 3334 3053
rect 3300 3019 3334 3052
rect 3300 2950 3334 2981
rect 3300 2947 3334 2950
rect 3300 2882 3334 2909
rect 3300 2875 3334 2882
rect 3300 2814 3334 2837
rect 3300 2803 3334 2814
rect 3300 2746 3334 2765
rect 3300 2731 3334 2746
rect 3300 2678 3334 2693
rect 3300 2659 3334 2678
rect 3300 2610 3334 2621
rect 3300 2587 3334 2610
rect 3300 2542 3334 2549
rect 3300 2515 3334 2542
rect 3300 2474 3334 2477
rect 3300 2443 3334 2474
rect 3300 2372 3334 2405
rect 3300 2371 3334 2372
rect 3300 2304 3334 2333
rect 3300 2299 3334 2304
rect 3300 2236 3334 2261
rect 3300 2227 3334 2236
rect 3300 2168 3334 2189
rect 3300 2155 3334 2168
rect 3300 2100 3334 2117
rect 3300 2083 3334 2100
rect 3300 2032 3334 2045
rect 3300 2011 3334 2032
rect 3300 1964 3334 1973
rect 3300 1939 3334 1964
rect 3300 1896 3334 1901
rect 3300 1867 3334 1896
rect 3300 1828 3334 1829
rect 3300 1795 3334 1828
rect 3300 1726 3334 1757
rect 3300 1723 3334 1726
rect 3300 1658 3334 1685
rect 3300 1651 3334 1658
rect 3300 1590 3334 1613
rect 3300 1579 3334 1590
rect 3300 1522 3334 1541
rect 3300 1507 3334 1522
rect 3300 1454 3334 1469
rect 3300 1435 3334 1454
rect 3300 1386 3334 1397
rect 3300 1363 3334 1386
rect 3300 1318 3334 1325
rect 3300 1291 3334 1318
rect 3300 1250 3334 1253
rect 3300 1219 3334 1250
rect 3300 1148 3334 1181
rect 3300 1147 3334 1148
rect 3300 1080 3334 1109
rect 3300 1075 3334 1080
rect 3300 1012 3334 1037
rect 3300 1003 3334 1012
rect 3300 944 3334 965
rect 3300 931 3334 944
rect 3300 876 3334 893
rect 3300 859 3334 876
rect 3300 808 3334 821
rect 3300 787 3334 808
rect 3300 740 3334 749
rect 3300 715 3334 740
rect 3300 672 3334 677
rect 3300 643 3334 672
rect 3300 604 3334 605
rect 3300 571 3334 604
rect 3300 502 3334 533
rect 3300 499 3334 502
rect 3300 434 3334 461
rect 3300 427 3334 434
rect 3300 366 3334 389
rect 3300 355 3334 366
rect 3300 298 3334 317
rect 3300 283 3334 298
rect 3300 230 3334 245
rect 3300 211 3334 230
rect 3300 162 3334 173
rect 3300 139 3334 162
rect 3300 94 3334 101
rect 3300 67 3334 94
rect -3034 -76 -3000 -43
rect -3034 -77 -3000 -76
rect -3034 -144 -3000 -115
rect -3034 -149 -3000 -144
rect -3034 -212 -3000 -187
rect -3034 -221 -3000 -212
rect -3034 -280 -3000 -259
rect -3034 -293 -3000 -280
rect -3034 -348 -3000 -331
rect -3034 -365 -3000 -348
rect -3034 -416 -3000 -403
rect -3034 -437 -3000 -416
rect 3300 26 3334 29
rect 3300 -5 3334 26
rect 3300 -76 3334 -43
rect 3300 -77 3334 -76
rect 3300 -144 3334 -115
rect 3300 -149 3334 -144
rect 3300 -212 3334 -187
rect 3300 -221 3334 -212
rect 3300 -280 3334 -259
rect 3300 -293 3334 -280
rect 3300 -348 3334 -331
rect 3300 -365 3334 -348
rect -3034 -484 -3000 -475
rect -3034 -509 -3000 -484
rect -3034 -552 -3000 -547
rect -3034 -581 -3000 -552
rect -3034 -620 -3000 -619
rect -3034 -653 -3000 -620
rect -180 -493 -146 -459
rect -106 -493 -72 -459
rect -32 -493 2 -459
rect 42 -493 76 -459
rect 116 -493 150 -459
rect 190 -493 224 -459
rect 264 -493 298 -459
rect 338 -493 372 -459
rect 412 -493 446 -459
rect 486 -493 520 -459
rect -180 -567 -146 -533
rect -106 -567 -72 -533
rect -32 -567 2 -533
rect 42 -567 76 -533
rect 116 -567 150 -533
rect 190 -567 224 -533
rect 264 -567 298 -533
rect 338 -567 372 -533
rect 412 -567 446 -533
rect 486 -567 520 -533
rect -180 -641 -146 -607
rect -106 -641 -72 -607
rect -32 -641 2 -607
rect 42 -641 76 -607
rect 116 -641 150 -607
rect 190 -641 224 -607
rect 264 -641 298 -607
rect 338 -641 372 -607
rect 412 -641 446 -607
rect 486 -641 520 -607
rect 3300 -416 3334 -403
rect 3300 -437 3334 -416
rect 3300 -484 3334 -475
rect 3300 -509 3334 -484
rect 3300 -552 3334 -547
rect 3300 -581 3334 -552
rect 3300 -620 3334 -619
rect 3300 -653 3334 -620
rect -3034 -722 -3000 -691
rect -3034 -725 -3000 -722
rect -3034 -790 -3000 -763
rect -3034 -797 -3000 -790
rect -3034 -858 -3000 -835
rect -3034 -869 -3000 -858
rect -3034 -926 -3000 -907
rect -3034 -941 -3000 -926
rect -3034 -994 -3000 -979
rect -3034 -1013 -3000 -994
rect -3034 -1062 -3000 -1051
rect -3034 -1085 -3000 -1062
rect -3034 -1130 -3000 -1123
rect -3034 -1157 -3000 -1130
rect -3034 -1198 -3000 -1195
rect -3034 -1229 -3000 -1198
rect -3034 -1300 -3000 -1267
rect -3034 -1301 -3000 -1300
rect -3034 -1368 -3000 -1339
rect -3034 -1373 -3000 -1368
rect -3034 -1436 -3000 -1411
rect -3034 -1445 -3000 -1436
rect -3034 -1504 -3000 -1483
rect -3034 -1517 -3000 -1504
rect -3034 -1572 -3000 -1555
rect -3034 -1589 -3000 -1572
rect -3034 -1640 -3000 -1627
rect -3034 -1661 -3000 -1640
rect -3034 -1708 -3000 -1699
rect -3034 -1733 -3000 -1708
rect -3034 -1776 -3000 -1771
rect -3034 -1805 -3000 -1776
rect -3034 -1877 -3000 -1843
rect 3300 -722 3334 -691
rect 3300 -725 3334 -722
rect 3300 -790 3334 -763
rect 3300 -797 3334 -790
rect 3300 -858 3334 -835
rect 3300 -869 3334 -858
rect 3300 -926 3334 -907
rect 3300 -941 3334 -926
rect 3300 -994 3334 -979
rect 3300 -1013 3334 -994
rect 3300 -1062 3334 -1051
rect 3300 -1085 3334 -1062
rect 3300 -1130 3334 -1123
rect 3300 -1157 3334 -1130
rect 3300 -1198 3334 -1195
rect 3300 -1229 3334 -1198
rect 3300 -1300 3334 -1267
rect 3300 -1301 3334 -1300
rect 3300 -1368 3334 -1339
rect 3300 -1373 3334 -1368
rect 3300 -1436 3334 -1411
rect 3300 -1445 3334 -1436
rect 3300 -1504 3334 -1483
rect 3300 -1517 3334 -1504
rect 3300 -1572 3334 -1555
rect 3300 -1589 3334 -1572
rect 3300 -1640 3334 -1627
rect 3300 -1661 3334 -1640
rect 3300 -1708 3334 -1699
rect 3300 -1733 3334 -1708
rect 3300 -1776 3334 -1771
rect 3300 -1805 3334 -1776
rect 3300 -1877 3334 -1843
rect -2927 -1958 -2893 -1924
rect -2855 -1958 -2825 -1924
rect -2825 -1958 -2821 -1924
rect -2783 -1958 -2757 -1924
rect -2757 -1958 -2749 -1924
rect -2711 -1958 -2689 -1924
rect -2689 -1958 -2677 -1924
rect -2639 -1958 -2621 -1924
rect -2621 -1958 -2605 -1924
rect -2567 -1958 -2553 -1924
rect -2553 -1958 -2533 -1924
rect -2495 -1958 -2485 -1924
rect -2485 -1958 -2461 -1924
rect -2423 -1958 -2417 -1924
rect -2417 -1958 -2389 -1924
rect -2351 -1958 -2349 -1924
rect -2349 -1958 -2317 -1924
rect -2279 -1958 -2247 -1924
rect -2247 -1958 -2245 -1924
rect -2207 -1958 -2179 -1924
rect -2179 -1958 -2173 -1924
rect -2135 -1958 -2111 -1924
rect -2111 -1958 -2101 -1924
rect -2063 -1958 -2043 -1924
rect -2043 -1958 -2029 -1924
rect -1991 -1958 -1975 -1924
rect -1975 -1958 -1957 -1924
rect -1919 -1958 -1907 -1924
rect -1907 -1958 -1885 -1924
rect -1847 -1958 -1839 -1924
rect -1839 -1958 -1813 -1924
rect -1775 -1958 -1771 -1924
rect -1771 -1958 -1741 -1924
rect -1703 -1958 -1669 -1924
rect -1631 -1958 -1601 -1924
rect -1601 -1958 -1597 -1924
rect -1559 -1958 -1533 -1924
rect -1533 -1958 -1525 -1924
rect -1487 -1958 -1465 -1924
rect -1465 -1958 -1453 -1924
rect -1415 -1958 -1397 -1924
rect -1397 -1958 -1381 -1924
rect -1343 -1958 -1329 -1924
rect -1329 -1958 -1309 -1924
rect -1271 -1958 -1261 -1924
rect -1261 -1958 -1237 -1924
rect -1199 -1958 -1193 -1924
rect -1193 -1958 -1165 -1924
rect -1127 -1958 -1125 -1924
rect -1125 -1958 -1093 -1924
rect -1055 -1958 -1023 -1924
rect -1023 -1958 -1021 -1924
rect -983 -1958 -955 -1924
rect -955 -1958 -949 -1924
rect -911 -1958 -887 -1924
rect -887 -1958 -877 -1924
rect -839 -1958 -819 -1924
rect -819 -1958 -805 -1924
rect -767 -1958 -751 -1924
rect -751 -1958 -733 -1924
rect -695 -1958 -683 -1924
rect -683 -1958 -661 -1924
rect -623 -1958 -615 -1924
rect -615 -1958 -589 -1924
rect -551 -1958 -547 -1924
rect -547 -1958 -517 -1924
rect -479 -1958 -445 -1924
rect -407 -1958 -377 -1924
rect -377 -1958 -373 -1924
rect -335 -1958 -309 -1924
rect -309 -1958 -301 -1924
rect -263 -1958 -241 -1924
rect -241 -1958 -229 -1924
rect -191 -1958 -173 -1924
rect -173 -1958 -157 -1924
rect -119 -1958 -105 -1924
rect -105 -1958 -85 -1924
rect -47 -1958 -37 -1924
rect -37 -1958 -13 -1924
rect 25 -1958 31 -1924
rect 31 -1958 59 -1924
rect 97 -1958 99 -1924
rect 99 -1958 131 -1924
rect 169 -1958 201 -1924
rect 201 -1958 203 -1924
rect 241 -1958 269 -1924
rect 269 -1958 275 -1924
rect 313 -1958 337 -1924
rect 337 -1958 347 -1924
rect 385 -1958 405 -1924
rect 405 -1958 419 -1924
rect 457 -1958 473 -1924
rect 473 -1958 491 -1924
rect 529 -1958 541 -1924
rect 541 -1958 563 -1924
rect 601 -1958 609 -1924
rect 609 -1958 635 -1924
rect 673 -1958 677 -1924
rect 677 -1958 707 -1924
rect 745 -1958 779 -1924
rect 817 -1958 847 -1924
rect 847 -1958 851 -1924
rect 889 -1958 915 -1924
rect 915 -1958 923 -1924
rect 961 -1958 983 -1924
rect 983 -1958 995 -1924
rect 1033 -1958 1051 -1924
rect 1051 -1958 1067 -1924
rect 1105 -1958 1119 -1924
rect 1119 -1958 1139 -1924
rect 1177 -1958 1187 -1924
rect 1187 -1958 1211 -1924
rect 1249 -1958 1255 -1924
rect 1255 -1958 1283 -1924
rect 1321 -1958 1323 -1924
rect 1323 -1958 1355 -1924
rect 1393 -1958 1425 -1924
rect 1425 -1958 1427 -1924
rect 1465 -1958 1493 -1924
rect 1493 -1958 1499 -1924
rect 1537 -1958 1561 -1924
rect 1561 -1958 1571 -1924
rect 1609 -1958 1629 -1924
rect 1629 -1958 1643 -1924
rect 1681 -1958 1697 -1924
rect 1697 -1958 1715 -1924
rect 1753 -1958 1765 -1924
rect 1765 -1958 1787 -1924
rect 1825 -1958 1833 -1924
rect 1833 -1958 1859 -1924
rect 1897 -1958 1901 -1924
rect 1901 -1958 1931 -1924
rect 1969 -1958 2003 -1924
rect 2041 -1958 2071 -1924
rect 2071 -1958 2075 -1924
rect 2113 -1958 2139 -1924
rect 2139 -1958 2147 -1924
rect 2185 -1958 2207 -1924
rect 2207 -1958 2219 -1924
rect 2257 -1958 2275 -1924
rect 2275 -1958 2291 -1924
rect 2329 -1958 2343 -1924
rect 2343 -1958 2363 -1924
rect 2401 -1958 2411 -1924
rect 2411 -1958 2435 -1924
rect 2473 -1958 2479 -1924
rect 2479 -1958 2507 -1924
rect 2545 -1958 2547 -1924
rect 2547 -1958 2579 -1924
rect 2617 -1958 2649 -1924
rect 2649 -1958 2651 -1924
rect 2689 -1958 2717 -1924
rect 2717 -1958 2723 -1924
rect 2761 -1958 2785 -1924
rect 2785 -1958 2795 -1924
rect 2833 -1958 2853 -1924
rect 2853 -1958 2867 -1924
rect 2905 -1958 2921 -1924
rect 2921 -1958 2939 -1924
rect 2977 -1958 2989 -1924
rect 2989 -1958 3011 -1924
rect 3049 -1958 3057 -1924
rect 3057 -1958 3083 -1924
rect 3121 -1958 3125 -1924
rect 3125 -1958 3155 -1924
rect 3193 -1958 3227 -1924
<< metal1 >>
rect -3058 7959 3358 7983
rect -3058 7925 -2927 7959
rect -2893 7925 -2855 7959
rect -2821 7925 -2783 7959
rect -2749 7925 -2711 7959
rect -2677 7925 -2639 7959
rect -2605 7925 -2567 7959
rect -2533 7925 -2495 7959
rect -2461 7925 -2423 7959
rect -2389 7925 -2351 7959
rect -2317 7925 -2279 7959
rect -2245 7925 -2207 7959
rect -2173 7925 -2135 7959
rect -2101 7925 -2063 7959
rect -2029 7925 -1991 7959
rect -1957 7925 -1919 7959
rect -1885 7925 -1847 7959
rect -1813 7925 -1775 7959
rect -1741 7925 -1703 7959
rect -1669 7925 -1631 7959
rect -1597 7925 -1559 7959
rect -1525 7925 -1487 7959
rect -1453 7925 -1415 7959
rect -1381 7925 -1343 7959
rect -1309 7925 -1271 7959
rect -1237 7925 -1199 7959
rect -1165 7925 -1127 7959
rect -1093 7925 -1055 7959
rect -1021 7925 -983 7959
rect -949 7925 -911 7959
rect -877 7925 -839 7959
rect -805 7925 -767 7959
rect -733 7925 -695 7959
rect -661 7925 -623 7959
rect -589 7925 -551 7959
rect -517 7925 -479 7959
rect -445 7925 -407 7959
rect -373 7925 -335 7959
rect -301 7925 -263 7959
rect -229 7925 -191 7959
rect -157 7925 -119 7959
rect -85 7925 -47 7959
rect -13 7925 25 7959
rect 59 7925 97 7959
rect 131 7925 169 7959
rect 203 7925 241 7959
rect 275 7925 313 7959
rect 347 7925 385 7959
rect 419 7925 457 7959
rect 491 7925 529 7959
rect 563 7925 601 7959
rect 635 7925 673 7959
rect 707 7925 745 7959
rect 779 7925 817 7959
rect 851 7925 889 7959
rect 923 7925 961 7959
rect 995 7925 1033 7959
rect 1067 7925 1105 7959
rect 1139 7925 1177 7959
rect 1211 7925 1249 7959
rect 1283 7925 1321 7959
rect 1355 7925 1393 7959
rect 1427 7925 1465 7959
rect 1499 7925 1537 7959
rect 1571 7925 1609 7959
rect 1643 7925 1681 7959
rect 1715 7925 1753 7959
rect 1787 7925 1825 7959
rect 1859 7925 1897 7959
rect 1931 7925 1969 7959
rect 2003 7925 2041 7959
rect 2075 7925 2113 7959
rect 2147 7925 2185 7959
rect 2219 7925 2257 7959
rect 2291 7925 2329 7959
rect 2363 7925 2401 7959
rect 2435 7925 2473 7959
rect 2507 7925 2545 7959
rect 2579 7925 2617 7959
rect 2651 7925 2689 7959
rect 2723 7925 2761 7959
rect 2795 7925 2833 7959
rect 2867 7925 2905 7959
rect 2939 7925 2977 7959
rect 3011 7925 3049 7959
rect 3083 7925 3121 7959
rect 3155 7925 3193 7959
rect 3227 7925 3358 7959
rect -3058 7901 3358 7925
rect -3058 7877 -2976 7901
rect -3058 7843 -3034 7877
rect -3000 7843 -2976 7877
rect -3058 7805 -2976 7843
rect -3058 7771 -3034 7805
rect -3000 7771 -2976 7805
rect -3058 7733 -2976 7771
rect -3058 7699 -3034 7733
rect -3000 7699 -2976 7733
rect -3058 7661 -2976 7699
rect -3058 7627 -3034 7661
rect -3000 7627 -2976 7661
rect -3058 7589 -2976 7627
rect -3058 7555 -3034 7589
rect -3000 7555 -2976 7589
rect -3058 7517 -2976 7555
rect -3058 7483 -3034 7517
rect -3000 7483 -2976 7517
rect -3058 7445 -2976 7483
rect -3058 7411 -3034 7445
rect -3000 7411 -2976 7445
rect -3058 7373 -2976 7411
rect -3058 7339 -3034 7373
rect -3000 7339 -2976 7373
rect -3058 7301 -2976 7339
rect -3058 7267 -3034 7301
rect -3000 7267 -2976 7301
rect -3058 7229 -2976 7267
rect -3058 7195 -3034 7229
rect -3000 7195 -2976 7229
rect -3058 7157 -2976 7195
rect -3058 7123 -3034 7157
rect -3000 7123 -2976 7157
rect -3058 7085 -2976 7123
rect -3058 7051 -3034 7085
rect -3000 7051 -2976 7085
rect -3058 7013 -2976 7051
rect -3058 6979 -3034 7013
rect -3000 6979 -2976 7013
rect -3058 6941 -2976 6979
rect -3058 6907 -3034 6941
rect -3000 6907 -2976 6941
rect -3058 6869 -2976 6907
rect -3058 6835 -3034 6869
rect -3000 6835 -2976 6869
rect -3058 6797 -2976 6835
rect -3058 6763 -3034 6797
rect -3000 6763 -2976 6797
rect -3058 6725 -2976 6763
rect -3058 6691 -3034 6725
rect -3000 6691 -2976 6725
rect -3058 6653 -2976 6691
rect -3058 6619 -3034 6653
rect -3000 6619 -2976 6653
rect -3058 6581 -2976 6619
rect -3058 6547 -3034 6581
rect -3000 6547 -2976 6581
rect -3058 6509 -2976 6547
rect -3058 6475 -3034 6509
rect -3000 6475 -2976 6509
rect -3058 6437 -2976 6475
rect -3058 6403 -3034 6437
rect -3000 6403 -2976 6437
rect -3058 6365 -2976 6403
rect -3058 6331 -3034 6365
rect -3000 6331 -2976 6365
rect -3058 6293 -2976 6331
rect -3058 6259 -3034 6293
rect -3000 6259 -2976 6293
rect -3058 6221 -2976 6259
rect -3058 6187 -3034 6221
rect -3000 6187 -2976 6221
rect -3058 6149 -2976 6187
rect -3058 6115 -3034 6149
rect -3000 6115 -2976 6149
rect -3058 6077 -2976 6115
rect -3058 6043 -3034 6077
rect -3000 6043 -2976 6077
rect -3058 6005 -2976 6043
rect -3058 5971 -3034 6005
rect -3000 5971 -2976 6005
rect 3276 7877 3358 7901
rect 3276 7843 3300 7877
rect 3334 7843 3358 7877
rect 3276 7805 3358 7843
rect 3276 7771 3300 7805
rect 3334 7771 3358 7805
rect 3276 7733 3358 7771
rect 3276 7699 3300 7733
rect 3334 7699 3358 7733
rect 3276 7661 3358 7699
rect 3276 7627 3300 7661
rect 3334 7627 3358 7661
rect 3276 7589 3358 7627
rect 3276 7555 3300 7589
rect 3334 7555 3358 7589
rect 3276 7517 3358 7555
rect 3276 7483 3300 7517
rect 3334 7483 3358 7517
rect 3276 7445 3358 7483
rect 3276 7411 3300 7445
rect 3334 7411 3358 7445
rect 3276 7373 3358 7411
rect 3276 7339 3300 7373
rect 3334 7339 3358 7373
rect 3276 7301 3358 7339
rect 3276 7267 3300 7301
rect 3334 7267 3358 7301
rect 3276 7229 3358 7267
rect 3276 7195 3300 7229
rect 3334 7195 3358 7229
rect 3276 7157 3358 7195
rect 3276 7123 3300 7157
rect 3334 7123 3358 7157
rect 3276 7085 3358 7123
rect 3276 7051 3300 7085
rect 3334 7051 3358 7085
rect 3276 7013 3358 7051
rect 3276 6979 3300 7013
rect 3334 6979 3358 7013
rect 3276 6941 3358 6979
rect 3276 6907 3300 6941
rect 3334 6907 3358 6941
rect 3276 6869 3358 6907
rect 3276 6835 3300 6869
rect 3334 6835 3358 6869
rect 3276 6797 3358 6835
rect 3276 6763 3300 6797
rect 3334 6763 3358 6797
rect 3276 6725 3358 6763
rect 3276 6691 3300 6725
rect 3334 6691 3358 6725
rect 3276 6653 3358 6691
rect 3276 6619 3300 6653
rect 3334 6619 3358 6653
rect 3276 6581 3358 6619
rect 3276 6547 3300 6581
rect 3334 6547 3358 6581
rect 3276 6509 3358 6547
rect 3276 6475 3300 6509
rect 3334 6475 3358 6509
rect 3276 6437 3358 6475
rect 3276 6403 3300 6437
rect 3334 6403 3358 6437
rect 3276 6365 3358 6403
rect 3276 6331 3300 6365
rect 3334 6331 3358 6365
rect 3276 6293 3358 6331
rect 3276 6259 3300 6293
rect 3334 6259 3358 6293
rect 3276 6221 3358 6259
rect 3276 6187 3300 6221
rect 3334 6187 3358 6221
rect 3276 6149 3358 6187
rect 3276 6115 3300 6149
rect 3334 6115 3358 6149
rect 3276 6077 3358 6115
rect 3276 6043 3300 6077
rect 3334 6043 3358 6077
rect 3276 6005 3358 6043
rect -3058 5933 -2976 5971
rect -3058 5899 -3034 5933
rect -3000 5899 -2976 5933
rect -3058 5861 -2976 5899
rect -3058 5827 -3034 5861
rect -3000 5827 -2976 5861
rect -3058 5789 -2976 5827
rect -3058 5755 -3034 5789
rect -3000 5755 -2976 5789
rect -3058 5717 -2976 5755
rect -3058 5683 -3034 5717
rect -3000 5683 -2976 5717
rect -3058 5645 -2976 5683
rect -3058 5611 -3034 5645
rect -3000 5611 -2976 5645
rect -3058 5573 -2976 5611
rect -3058 5539 -3034 5573
rect -3000 5539 -2976 5573
rect -3058 5501 -2976 5539
rect -3058 5467 -3034 5501
rect -3000 5467 -2976 5501
rect -3058 5429 -2976 5467
rect -3058 5395 -3034 5429
rect -3000 5395 -2976 5429
rect -3058 5357 -2976 5395
rect -3058 5323 -3034 5357
rect -3000 5323 -2976 5357
rect -3058 5285 -2976 5323
rect -3058 5251 -3034 5285
rect -3000 5251 -2976 5285
rect -3058 5213 -2976 5251
rect -3058 5179 -3034 5213
rect -3000 5179 -2976 5213
rect -3058 5141 -2976 5179
rect -3058 5107 -3034 5141
rect -3000 5107 -2976 5141
rect -3058 5069 -2976 5107
rect -3058 5035 -3034 5069
rect -3000 5035 -2976 5069
rect -3058 4997 -2976 5035
rect -3058 4963 -3034 4997
rect -3000 4963 -2976 4997
rect -3058 4925 -2976 4963
rect -3058 4891 -3034 4925
rect -3000 4891 -2976 4925
rect -3058 4853 -2976 4891
rect -3058 4819 -3034 4853
rect -3000 4819 -2976 4853
rect -3058 4781 -2976 4819
rect -3058 4747 -3034 4781
rect -3000 4747 -2976 4781
rect -3058 4709 -2976 4747
rect -3058 4675 -3034 4709
rect -3000 4675 -2976 4709
rect -3058 4637 -2976 4675
rect -3058 4603 -3034 4637
rect -3000 4603 -2976 4637
rect -3058 4565 -2976 4603
rect -3058 4531 -3034 4565
rect -3000 4531 -2976 4565
rect -3058 4493 -2976 4531
rect -3058 4459 -3034 4493
rect -3000 4459 -2976 4493
rect -3058 4421 -2976 4459
rect -3058 4387 -3034 4421
rect -3000 4387 -2976 4421
rect -3058 4349 -2976 4387
rect -3058 4315 -3034 4349
rect -3000 4315 -2976 4349
rect -3058 4277 -2976 4315
rect -3058 4243 -3034 4277
rect -3000 4243 -2976 4277
rect -3058 4205 -2976 4243
rect -3058 4171 -3034 4205
rect -3000 4171 -2976 4205
rect -3058 4133 -2976 4171
rect -3058 4099 -3034 4133
rect -3000 4099 -2976 4133
rect -3058 4061 -2976 4099
rect -3058 4027 -3034 4061
rect -3000 4027 -2976 4061
rect -3058 3989 -2976 4027
rect -3058 3955 -3034 3989
rect -3000 3955 -2976 3989
rect -3058 3917 -2976 3955
rect -3058 3883 -3034 3917
rect -3000 3883 -2976 3917
rect -3058 3845 -2976 3883
rect -3058 3811 -3034 3845
rect -3000 3811 -2976 3845
rect -3058 3773 -2976 3811
rect -3058 3739 -3034 3773
rect -3000 3739 -2976 3773
rect -3058 3701 -2976 3739
rect -3058 3667 -3034 3701
rect -3000 3667 -2976 3701
rect -3058 3629 -2976 3667
rect -3058 3595 -3034 3629
rect -3000 3595 -2976 3629
rect -3058 3557 -2976 3595
rect -3058 3523 -3034 3557
rect -3000 3523 -2976 3557
rect -3058 3485 -2976 3523
rect -3058 3451 -3034 3485
rect -3000 3451 -2976 3485
rect -3058 3413 -2976 3451
rect -3058 3379 -3034 3413
rect -3000 3379 -2976 3413
rect -3058 3341 -2976 3379
rect -3058 3307 -3034 3341
rect -3000 3307 -2976 3341
rect -3058 3269 -2976 3307
rect -3058 3235 -3034 3269
rect -3000 3235 -2976 3269
rect -3058 3197 -2976 3235
rect -3058 3163 -3034 3197
rect -3000 3163 -2976 3197
rect -3058 3125 -2976 3163
rect -3058 3091 -3034 3125
rect -3000 3091 -2976 3125
rect -3058 3053 -2976 3091
rect -3058 3019 -3034 3053
rect -3000 3019 -2976 3053
rect -3058 2981 -2976 3019
rect -3058 2947 -3034 2981
rect -3000 2947 -2976 2981
rect -3058 2909 -2976 2947
rect -3058 2875 -3034 2909
rect -3000 2875 -2976 2909
rect -3058 2837 -2976 2875
rect -3058 2803 -3034 2837
rect -3000 2803 -2976 2837
rect -3058 2765 -2976 2803
rect -3058 2731 -3034 2765
rect -3000 2731 -2976 2765
rect -3058 2693 -2976 2731
rect -3058 2659 -3034 2693
rect -3000 2659 -2976 2693
rect -3058 2621 -2976 2659
rect -3058 2587 -3034 2621
rect -3000 2587 -2976 2621
rect -3058 2549 -2976 2587
rect -3058 2515 -3034 2549
rect -3000 2515 -2976 2549
rect -3058 2477 -2976 2515
rect -3058 2443 -3034 2477
rect -3000 2443 -2976 2477
rect -3058 2405 -2976 2443
rect -3058 2371 -3034 2405
rect -3000 2371 -2976 2405
rect -3058 2333 -2976 2371
rect -3058 2299 -3034 2333
rect -3000 2299 -2976 2333
rect -3058 2261 -2976 2299
rect -3058 2227 -3034 2261
rect -3000 2227 -2976 2261
rect -3058 2189 -2976 2227
rect -3058 2155 -3034 2189
rect -3000 2155 -2976 2189
rect -3058 2117 -2976 2155
rect -3058 2083 -3034 2117
rect -3000 2083 -2976 2117
rect -3058 2045 -2976 2083
rect -3058 2011 -3034 2045
rect -3000 2011 -2976 2045
rect -3058 1973 -2976 2011
rect -3058 1939 -3034 1973
rect -3000 1939 -2976 1973
rect -3058 1901 -2976 1939
rect -3058 1867 -3034 1901
rect -3000 1867 -2976 1901
rect -3058 1829 -2976 1867
rect -3058 1795 -3034 1829
rect -3000 1795 -2976 1829
rect -3058 1757 -2976 1795
rect -3058 1723 -3034 1757
rect -3000 1723 -2976 1757
rect -3058 1685 -2976 1723
rect -3058 1651 -3034 1685
rect -3000 1651 -2976 1685
rect -3058 1613 -2976 1651
rect -3058 1579 -3034 1613
rect -3000 1579 -2976 1613
rect -3058 1541 -2976 1579
rect -3058 1507 -3034 1541
rect -3000 1507 -2976 1541
rect -3058 1469 -2976 1507
rect -3058 1435 -3034 1469
rect -3000 1435 -2976 1469
rect -3058 1397 -2976 1435
rect -3058 1363 -3034 1397
rect -3000 1363 -2976 1397
rect -3058 1325 -2976 1363
rect -3058 1291 -3034 1325
rect -3000 1291 -2976 1325
rect -3058 1253 -2976 1291
rect -3058 1219 -3034 1253
rect -3000 1219 -2976 1253
rect -3058 1181 -2976 1219
rect -3058 1147 -3034 1181
rect -3000 1147 -2976 1181
rect -3058 1109 -2976 1147
rect -3058 1075 -3034 1109
rect -3000 1075 -2976 1109
rect -3058 1037 -2976 1075
rect -3058 1003 -3034 1037
rect -3000 1003 -2976 1037
rect -3058 965 -2976 1003
rect -3058 931 -3034 965
rect -3000 931 -2976 965
rect -3058 893 -2976 931
rect -3058 859 -3034 893
rect -3000 859 -2976 893
rect -3058 821 -2976 859
rect -3058 787 -3034 821
rect -3000 787 -2976 821
rect -3058 749 -2976 787
rect -3058 715 -3034 749
rect -3000 715 -2976 749
rect -3058 677 -2976 715
rect -3058 643 -3034 677
rect -3000 643 -2976 677
rect -3058 605 -2976 643
rect -3058 571 -3034 605
rect -3000 571 -2976 605
rect -3058 533 -2976 571
rect -3058 499 -3034 533
rect -3000 499 -2976 533
rect -3058 461 -2976 499
rect -3058 427 -3034 461
rect -3000 427 -2976 461
rect -3058 389 -2976 427
rect -3058 355 -3034 389
rect -3000 355 -2976 389
rect -3058 317 -2976 355
rect -3058 283 -3034 317
rect -3000 283 -2976 317
rect -3058 245 -2976 283
rect -3058 211 -3034 245
rect -3000 211 -2976 245
rect -3058 173 -2976 211
rect -3058 139 -3034 173
rect -3000 139 -2976 173
rect -3058 101 -2976 139
rect -3058 67 -3034 101
rect -3000 67 -2976 101
rect -3058 29 -2976 67
rect -3058 -5 -3034 29
rect -3000 -5 -2976 29
rect -1066 5969 -936 5981
rect -1066 31 -1054 5969
rect -948 31 -936 5969
rect -1066 19 -936 31
rect -828 5969 -698 5981
rect -828 31 -816 5969
rect -710 31 -698 5969
rect 998 5969 1128 5981
rect 13 5939 287 5945
rect 13 5933 28 5939
rect 272 5933 287 5939
rect 13 67 25 5933
rect 275 67 287 5933
rect 13 63 28 67
rect 272 63 287 67
rect 13 55 287 63
rect -828 19 -698 31
rect 998 31 1010 5969
rect 1116 31 1128 5969
rect 998 19 1128 31
rect 1236 5969 1366 5981
rect 1236 31 1248 5969
rect 1354 31 1366 5969
rect 1236 19 1366 31
rect 3276 5971 3300 6005
rect 3334 5971 3358 6005
rect 3276 5933 3358 5971
rect 3276 5899 3300 5933
rect 3334 5899 3358 5933
rect 3276 5861 3358 5899
rect 3276 5827 3300 5861
rect 3334 5827 3358 5861
rect 3276 5789 3358 5827
rect 3276 5755 3300 5789
rect 3334 5755 3358 5789
rect 3276 5717 3358 5755
rect 3276 5683 3300 5717
rect 3334 5683 3358 5717
rect 3276 5645 3358 5683
rect 3276 5611 3300 5645
rect 3334 5611 3358 5645
rect 3276 5573 3358 5611
rect 3276 5539 3300 5573
rect 3334 5539 3358 5573
rect 3276 5501 3358 5539
rect 3276 5467 3300 5501
rect 3334 5467 3358 5501
rect 3276 5429 3358 5467
rect 3276 5395 3300 5429
rect 3334 5395 3358 5429
rect 3276 5357 3358 5395
rect 3276 5323 3300 5357
rect 3334 5323 3358 5357
rect 3276 5285 3358 5323
rect 3276 5251 3300 5285
rect 3334 5251 3358 5285
rect 3276 5213 3358 5251
rect 3276 5179 3300 5213
rect 3334 5179 3358 5213
rect 3276 5141 3358 5179
rect 3276 5107 3300 5141
rect 3334 5107 3358 5141
rect 3276 5069 3358 5107
rect 3276 5035 3300 5069
rect 3334 5035 3358 5069
rect 3276 4997 3358 5035
rect 3276 4963 3300 4997
rect 3334 4963 3358 4997
rect 3276 4925 3358 4963
rect 3276 4891 3300 4925
rect 3334 4891 3358 4925
rect 3276 4853 3358 4891
rect 3276 4819 3300 4853
rect 3334 4819 3358 4853
rect 3276 4781 3358 4819
rect 3276 4747 3300 4781
rect 3334 4747 3358 4781
rect 3276 4709 3358 4747
rect 3276 4675 3300 4709
rect 3334 4675 3358 4709
rect 3276 4637 3358 4675
rect 3276 4603 3300 4637
rect 3334 4603 3358 4637
rect 3276 4565 3358 4603
rect 3276 4531 3300 4565
rect 3334 4531 3358 4565
rect 3276 4493 3358 4531
rect 3276 4459 3300 4493
rect 3334 4459 3358 4493
rect 3276 4421 3358 4459
rect 3276 4387 3300 4421
rect 3334 4387 3358 4421
rect 3276 4349 3358 4387
rect 3276 4315 3300 4349
rect 3334 4315 3358 4349
rect 3276 4277 3358 4315
rect 3276 4243 3300 4277
rect 3334 4243 3358 4277
rect 3276 4205 3358 4243
rect 3276 4171 3300 4205
rect 3334 4171 3358 4205
rect 3276 4133 3358 4171
rect 3276 4099 3300 4133
rect 3334 4099 3358 4133
rect 3276 4061 3358 4099
rect 3276 4027 3300 4061
rect 3334 4027 3358 4061
rect 3276 3989 3358 4027
rect 3276 3955 3300 3989
rect 3334 3955 3358 3989
rect 3276 3917 3358 3955
rect 3276 3883 3300 3917
rect 3334 3883 3358 3917
rect 3276 3845 3358 3883
rect 3276 3811 3300 3845
rect 3334 3811 3358 3845
rect 3276 3773 3358 3811
rect 3276 3739 3300 3773
rect 3334 3739 3358 3773
rect 3276 3701 3358 3739
rect 3276 3667 3300 3701
rect 3334 3667 3358 3701
rect 3276 3629 3358 3667
rect 3276 3595 3300 3629
rect 3334 3595 3358 3629
rect 3276 3557 3358 3595
rect 3276 3523 3300 3557
rect 3334 3523 3358 3557
rect 3276 3485 3358 3523
rect 3276 3451 3300 3485
rect 3334 3451 3358 3485
rect 3276 3413 3358 3451
rect 3276 3379 3300 3413
rect 3334 3379 3358 3413
rect 3276 3341 3358 3379
rect 3276 3307 3300 3341
rect 3334 3307 3358 3341
rect 3276 3269 3358 3307
rect 3276 3235 3300 3269
rect 3334 3235 3358 3269
rect 3276 3197 3358 3235
rect 3276 3163 3300 3197
rect 3334 3163 3358 3197
rect 3276 3125 3358 3163
rect 3276 3091 3300 3125
rect 3334 3091 3358 3125
rect 3276 3053 3358 3091
rect 3276 3019 3300 3053
rect 3334 3019 3358 3053
rect 3276 2981 3358 3019
rect 3276 2947 3300 2981
rect 3334 2947 3358 2981
rect 3276 2909 3358 2947
rect 3276 2875 3300 2909
rect 3334 2875 3358 2909
rect 3276 2837 3358 2875
rect 3276 2803 3300 2837
rect 3334 2803 3358 2837
rect 3276 2765 3358 2803
rect 3276 2731 3300 2765
rect 3334 2731 3358 2765
rect 3276 2693 3358 2731
rect 3276 2659 3300 2693
rect 3334 2659 3358 2693
rect 3276 2621 3358 2659
rect 3276 2587 3300 2621
rect 3334 2587 3358 2621
rect 3276 2549 3358 2587
rect 3276 2515 3300 2549
rect 3334 2515 3358 2549
rect 3276 2477 3358 2515
rect 3276 2443 3300 2477
rect 3334 2443 3358 2477
rect 3276 2405 3358 2443
rect 3276 2371 3300 2405
rect 3334 2371 3358 2405
rect 3276 2333 3358 2371
rect 3276 2299 3300 2333
rect 3334 2299 3358 2333
rect 3276 2261 3358 2299
rect 3276 2227 3300 2261
rect 3334 2227 3358 2261
rect 3276 2189 3358 2227
rect 3276 2155 3300 2189
rect 3334 2155 3358 2189
rect 3276 2117 3358 2155
rect 3276 2083 3300 2117
rect 3334 2083 3358 2117
rect 3276 2045 3358 2083
rect 3276 2011 3300 2045
rect 3334 2011 3358 2045
rect 3276 1973 3358 2011
rect 3276 1939 3300 1973
rect 3334 1939 3358 1973
rect 3276 1901 3358 1939
rect 3276 1867 3300 1901
rect 3334 1867 3358 1901
rect 3276 1829 3358 1867
rect 3276 1795 3300 1829
rect 3334 1795 3358 1829
rect 3276 1757 3358 1795
rect 3276 1723 3300 1757
rect 3334 1723 3358 1757
rect 3276 1685 3358 1723
rect 3276 1651 3300 1685
rect 3334 1651 3358 1685
rect 3276 1613 3358 1651
rect 3276 1579 3300 1613
rect 3334 1579 3358 1613
rect 3276 1541 3358 1579
rect 3276 1507 3300 1541
rect 3334 1507 3358 1541
rect 3276 1469 3358 1507
rect 3276 1435 3300 1469
rect 3334 1435 3358 1469
rect 3276 1397 3358 1435
rect 3276 1363 3300 1397
rect 3334 1363 3358 1397
rect 3276 1325 3358 1363
rect 3276 1291 3300 1325
rect 3334 1291 3358 1325
rect 3276 1253 3358 1291
rect 3276 1219 3300 1253
rect 3334 1219 3358 1253
rect 3276 1181 3358 1219
rect 3276 1147 3300 1181
rect 3334 1147 3358 1181
rect 3276 1109 3358 1147
rect 3276 1075 3300 1109
rect 3334 1075 3358 1109
rect 3276 1037 3358 1075
rect 3276 1003 3300 1037
rect 3334 1003 3358 1037
rect 3276 965 3358 1003
rect 3276 931 3300 965
rect 3334 931 3358 965
rect 3276 893 3358 931
rect 3276 859 3300 893
rect 3334 859 3358 893
rect 3276 821 3358 859
rect 3276 787 3300 821
rect 3334 787 3358 821
rect 3276 749 3358 787
rect 3276 715 3300 749
rect 3334 715 3358 749
rect 3276 677 3358 715
rect 3276 643 3300 677
rect 3334 643 3358 677
rect 3276 605 3358 643
rect 3276 571 3300 605
rect 3334 571 3358 605
rect 3276 533 3358 571
rect 3276 499 3300 533
rect 3334 499 3358 533
rect 3276 461 3358 499
rect 3276 427 3300 461
rect 3334 427 3358 461
rect 3276 389 3358 427
rect 3276 355 3300 389
rect 3334 355 3358 389
rect 3276 317 3358 355
rect 3276 283 3300 317
rect 3334 283 3358 317
rect 3276 245 3358 283
rect 3276 211 3300 245
rect 3334 211 3358 245
rect 3276 173 3358 211
rect 3276 139 3300 173
rect 3334 139 3358 173
rect 3276 101 3358 139
rect 3276 67 3300 101
rect 3334 67 3358 101
rect 3276 29 3358 67
rect -3058 -43 -2976 -5
rect -3058 -77 -3034 -43
rect -3000 -77 -2976 -43
rect -3058 -115 -2976 -77
rect -3058 -149 -3034 -115
rect -3000 -149 -2976 -115
rect -3058 -187 -2976 -149
rect -3058 -221 -3034 -187
rect -3000 -221 -2976 -187
rect -3058 -259 -2976 -221
rect -3058 -293 -3034 -259
rect -3000 -293 -2976 -259
rect -3058 -331 -2976 -293
rect -3058 -365 -3034 -331
rect -3000 -365 -2976 -331
rect -3058 -403 -2976 -365
rect -3058 -437 -3034 -403
rect -3000 -437 -2976 -403
rect -3058 -475 -2976 -437
rect 3276 -5 3300 29
rect 3334 -5 3358 29
rect 3276 -43 3358 -5
rect 3276 -77 3300 -43
rect 3334 -77 3358 -43
rect 3276 -115 3358 -77
rect 3276 -149 3300 -115
rect 3334 -149 3358 -115
rect 3276 -187 3358 -149
rect 3276 -221 3300 -187
rect 3334 -221 3358 -187
rect 3276 -259 3358 -221
rect 3276 -293 3300 -259
rect 3334 -293 3358 -259
rect 3276 -331 3358 -293
rect 3276 -365 3300 -331
rect 3334 -365 3358 -331
rect 3276 -403 3358 -365
rect 3276 -437 3300 -403
rect 3334 -437 3358 -403
rect -3058 -509 -3034 -475
rect -3000 -509 -2976 -475
rect -3058 -547 -2976 -509
rect -3058 -581 -3034 -547
rect -3000 -581 -2976 -547
rect -3058 -619 -2976 -581
rect -3058 -653 -3034 -619
rect -3000 -653 -2976 -619
rect -3058 -691 -2976 -653
rect -209 -450 555 -443
rect -209 -502 -189 -450
rect -137 -502 -115 -450
rect -63 -502 -41 -450
rect 11 -502 33 -450
rect 85 -502 107 -450
rect 159 -502 181 -450
rect 233 -502 255 -450
rect 307 -502 329 -450
rect 381 -502 403 -450
rect 455 -502 477 -450
rect 529 -502 555 -450
rect -209 -524 555 -502
rect -209 -576 -189 -524
rect -137 -576 -115 -524
rect -63 -576 -41 -524
rect 11 -576 33 -524
rect 85 -576 107 -524
rect 159 -576 181 -524
rect 233 -576 255 -524
rect 307 -576 329 -524
rect 381 -576 403 -524
rect 455 -576 477 -524
rect 529 -576 555 -524
rect -209 -598 555 -576
rect -209 -650 -189 -598
rect -137 -650 -115 -598
rect -63 -650 -41 -598
rect 11 -650 33 -598
rect 85 -650 107 -598
rect 159 -650 181 -598
rect 233 -650 255 -598
rect 307 -650 329 -598
rect 381 -650 403 -598
rect 455 -650 477 -598
rect 529 -650 555 -598
rect -209 -657 555 -650
rect 3276 -475 3358 -437
rect 3276 -509 3300 -475
rect 3334 -509 3358 -475
rect 3276 -547 3358 -509
rect 3276 -581 3300 -547
rect 3334 -581 3358 -547
rect 3276 -619 3358 -581
rect 3276 -653 3300 -619
rect 3334 -653 3358 -619
rect -3058 -725 -3034 -691
rect -3000 -725 -2976 -691
rect -3058 -763 -2976 -725
rect -3058 -797 -3034 -763
rect -3000 -797 -2976 -763
rect -3058 -835 -2976 -797
rect -3058 -869 -3034 -835
rect -3000 -869 -2976 -835
rect -3058 -907 -2976 -869
rect -3058 -941 -3034 -907
rect -3000 -941 -2976 -907
rect -3058 -979 -2976 -941
rect -3058 -1013 -3034 -979
rect -3000 -1013 -2976 -979
rect -3058 -1051 -2976 -1013
rect -3058 -1085 -3034 -1051
rect -3000 -1085 -2976 -1051
rect -3058 -1123 -2976 -1085
rect -3058 -1157 -3034 -1123
rect -3000 -1157 -2976 -1123
rect -3058 -1195 -2976 -1157
rect -3058 -1229 -3034 -1195
rect -3000 -1229 -2976 -1195
rect -3058 -1267 -2976 -1229
rect -3058 -1301 -3034 -1267
rect -3000 -1301 -2976 -1267
rect -3058 -1339 -2976 -1301
rect -3058 -1373 -3034 -1339
rect -3000 -1373 -2976 -1339
rect -3058 -1411 -2976 -1373
rect -3058 -1445 -3034 -1411
rect -3000 -1445 -2976 -1411
rect -3058 -1483 -2976 -1445
rect -3058 -1517 -3034 -1483
rect -3000 -1517 -2976 -1483
rect -3058 -1555 -2976 -1517
rect -3058 -1589 -3034 -1555
rect -3000 -1589 -2976 -1555
rect -3058 -1627 -2976 -1589
rect -3058 -1661 -3034 -1627
rect -3000 -1661 -2976 -1627
rect -3058 -1699 -2976 -1661
rect -3058 -1733 -3034 -1699
rect -3000 -1733 -2976 -1699
rect -3058 -1771 -2976 -1733
rect -3058 -1805 -3034 -1771
rect -3000 -1805 -2976 -1771
rect -3058 -1843 -2976 -1805
rect -3058 -1877 -3034 -1843
rect -3000 -1877 -2976 -1843
rect -3058 -1900 -2976 -1877
rect 3276 -691 3358 -653
rect 3276 -725 3300 -691
rect 3334 -725 3358 -691
rect 3276 -763 3358 -725
rect 3276 -797 3300 -763
rect 3334 -797 3358 -763
rect 3276 -835 3358 -797
rect 3276 -869 3300 -835
rect 3334 -869 3358 -835
rect 3276 -907 3358 -869
rect 3276 -941 3300 -907
rect 3334 -941 3358 -907
rect 3276 -979 3358 -941
rect 3276 -1013 3300 -979
rect 3334 -1013 3358 -979
rect 3276 -1051 3358 -1013
rect 3276 -1085 3300 -1051
rect 3334 -1085 3358 -1051
rect 3276 -1123 3358 -1085
rect 3276 -1157 3300 -1123
rect 3334 -1157 3358 -1123
rect 3276 -1195 3358 -1157
rect 3276 -1229 3300 -1195
rect 3334 -1229 3358 -1195
rect 3276 -1267 3358 -1229
rect 3276 -1301 3300 -1267
rect 3334 -1301 3358 -1267
rect 3276 -1339 3358 -1301
rect 3276 -1373 3300 -1339
rect 3334 -1373 3358 -1339
rect 3276 -1411 3358 -1373
rect 3276 -1445 3300 -1411
rect 3334 -1445 3358 -1411
rect 3276 -1483 3358 -1445
rect 3276 -1517 3300 -1483
rect 3334 -1517 3358 -1483
rect 3276 -1555 3358 -1517
rect 3276 -1589 3300 -1555
rect 3334 -1589 3358 -1555
rect 3276 -1627 3358 -1589
rect 3276 -1661 3300 -1627
rect 3334 -1661 3358 -1627
rect 3276 -1699 3358 -1661
rect 3276 -1733 3300 -1699
rect 3334 -1733 3358 -1699
rect 3276 -1771 3358 -1733
rect 3276 -1805 3300 -1771
rect 3334 -1805 3358 -1771
rect 3276 -1843 3358 -1805
rect 3276 -1877 3300 -1843
rect 3334 -1877 3358 -1843
rect 3276 -1900 3358 -1877
rect -3058 -1924 3358 -1900
rect -3058 -1958 -2927 -1924
rect -2893 -1958 -2855 -1924
rect -2821 -1958 -2783 -1924
rect -2749 -1958 -2711 -1924
rect -2677 -1958 -2639 -1924
rect -2605 -1958 -2567 -1924
rect -2533 -1958 -2495 -1924
rect -2461 -1958 -2423 -1924
rect -2389 -1958 -2351 -1924
rect -2317 -1958 -2279 -1924
rect -2245 -1958 -2207 -1924
rect -2173 -1958 -2135 -1924
rect -2101 -1958 -2063 -1924
rect -2029 -1958 -1991 -1924
rect -1957 -1958 -1919 -1924
rect -1885 -1958 -1847 -1924
rect -1813 -1958 -1775 -1924
rect -1741 -1958 -1703 -1924
rect -1669 -1958 -1631 -1924
rect -1597 -1958 -1559 -1924
rect -1525 -1958 -1487 -1924
rect -1453 -1958 -1415 -1924
rect -1381 -1958 -1343 -1924
rect -1309 -1958 -1271 -1924
rect -1237 -1958 -1199 -1924
rect -1165 -1958 -1127 -1924
rect -1093 -1958 -1055 -1924
rect -1021 -1958 -983 -1924
rect -949 -1958 -911 -1924
rect -877 -1958 -839 -1924
rect -805 -1958 -767 -1924
rect -733 -1958 -695 -1924
rect -661 -1958 -623 -1924
rect -589 -1958 -551 -1924
rect -517 -1958 -479 -1924
rect -445 -1958 -407 -1924
rect -373 -1958 -335 -1924
rect -301 -1958 -263 -1924
rect -229 -1958 -191 -1924
rect -157 -1958 -119 -1924
rect -85 -1958 -47 -1924
rect -13 -1958 25 -1924
rect 59 -1958 97 -1924
rect 131 -1958 169 -1924
rect 203 -1958 241 -1924
rect 275 -1958 313 -1924
rect 347 -1958 385 -1924
rect 419 -1958 457 -1924
rect 491 -1958 529 -1924
rect 563 -1958 601 -1924
rect 635 -1958 673 -1924
rect 707 -1958 745 -1924
rect 779 -1958 817 -1924
rect 851 -1958 889 -1924
rect 923 -1958 961 -1924
rect 995 -1958 1033 -1924
rect 1067 -1958 1105 -1924
rect 1139 -1958 1177 -1924
rect 1211 -1958 1249 -1924
rect 1283 -1958 1321 -1924
rect 1355 -1958 1393 -1924
rect 1427 -1958 1465 -1924
rect 1499 -1958 1537 -1924
rect 1571 -1958 1609 -1924
rect 1643 -1958 1681 -1924
rect 1715 -1958 1753 -1924
rect 1787 -1958 1825 -1924
rect 1859 -1958 1897 -1924
rect 1931 -1958 1969 -1924
rect 2003 -1958 2041 -1924
rect 2075 -1958 2113 -1924
rect 2147 -1958 2185 -1924
rect 2219 -1958 2257 -1924
rect 2291 -1958 2329 -1924
rect 2363 -1958 2401 -1924
rect 2435 -1958 2473 -1924
rect 2507 -1958 2545 -1924
rect 2579 -1958 2617 -1924
rect 2651 -1958 2689 -1924
rect 2723 -1958 2761 -1924
rect 2795 -1958 2833 -1924
rect 2867 -1958 2905 -1924
rect 2939 -1958 2977 -1924
rect 3011 -1958 3049 -1924
rect 3083 -1958 3121 -1924
rect 3155 -1958 3193 -1924
rect 3227 -1958 3358 -1924
rect -3058 -1982 3358 -1958
<< via1 >>
rect 28 5933 272 5939
rect 28 67 272 5933
rect 28 63 272 67
rect -189 -459 -137 -450
rect -189 -493 -180 -459
rect -180 -493 -146 -459
rect -146 -493 -137 -459
rect -189 -502 -137 -493
rect -115 -459 -63 -450
rect -115 -493 -106 -459
rect -106 -493 -72 -459
rect -72 -493 -63 -459
rect -115 -502 -63 -493
rect -41 -459 11 -450
rect -41 -493 -32 -459
rect -32 -493 2 -459
rect 2 -493 11 -459
rect -41 -502 11 -493
rect 33 -459 85 -450
rect 33 -493 42 -459
rect 42 -493 76 -459
rect 76 -493 85 -459
rect 33 -502 85 -493
rect 107 -459 159 -450
rect 107 -493 116 -459
rect 116 -493 150 -459
rect 150 -493 159 -459
rect 107 -502 159 -493
rect 181 -459 233 -450
rect 181 -493 190 -459
rect 190 -493 224 -459
rect 224 -493 233 -459
rect 181 -502 233 -493
rect 255 -459 307 -450
rect 255 -493 264 -459
rect 264 -493 298 -459
rect 298 -493 307 -459
rect 255 -502 307 -493
rect 329 -459 381 -450
rect 329 -493 338 -459
rect 338 -493 372 -459
rect 372 -493 381 -459
rect 329 -502 381 -493
rect 403 -459 455 -450
rect 403 -493 412 -459
rect 412 -493 446 -459
rect 446 -493 455 -459
rect 403 -502 455 -493
rect 477 -459 529 -450
rect 477 -493 486 -459
rect 486 -493 520 -459
rect 520 -493 529 -459
rect 477 -502 529 -493
rect -189 -533 -137 -524
rect -189 -567 -180 -533
rect -180 -567 -146 -533
rect -146 -567 -137 -533
rect -189 -576 -137 -567
rect -115 -533 -63 -524
rect -115 -567 -106 -533
rect -106 -567 -72 -533
rect -72 -567 -63 -533
rect -115 -576 -63 -567
rect -41 -533 11 -524
rect -41 -567 -32 -533
rect -32 -567 2 -533
rect 2 -567 11 -533
rect -41 -576 11 -567
rect 33 -533 85 -524
rect 33 -567 42 -533
rect 42 -567 76 -533
rect 76 -567 85 -533
rect 33 -576 85 -567
rect 107 -533 159 -524
rect 107 -567 116 -533
rect 116 -567 150 -533
rect 150 -567 159 -533
rect 107 -576 159 -567
rect 181 -533 233 -524
rect 181 -567 190 -533
rect 190 -567 224 -533
rect 224 -567 233 -533
rect 181 -576 233 -567
rect 255 -533 307 -524
rect 255 -567 264 -533
rect 264 -567 298 -533
rect 298 -567 307 -533
rect 255 -576 307 -567
rect 329 -533 381 -524
rect 329 -567 338 -533
rect 338 -567 372 -533
rect 372 -567 381 -533
rect 329 -576 381 -567
rect 403 -533 455 -524
rect 403 -567 412 -533
rect 412 -567 446 -533
rect 446 -567 455 -533
rect 403 -576 455 -567
rect 477 -533 529 -524
rect 477 -567 486 -533
rect 486 -567 520 -533
rect 520 -567 529 -533
rect 477 -576 529 -567
rect -189 -607 -137 -598
rect -189 -641 -180 -607
rect -180 -641 -146 -607
rect -146 -641 -137 -607
rect -189 -650 -137 -641
rect -115 -607 -63 -598
rect -115 -641 -106 -607
rect -106 -641 -72 -607
rect -72 -641 -63 -607
rect -115 -650 -63 -641
rect -41 -607 11 -598
rect -41 -641 -32 -607
rect -32 -641 2 -607
rect 2 -641 11 -607
rect -41 -650 11 -641
rect 33 -607 85 -598
rect 33 -641 42 -607
rect 42 -641 76 -607
rect 76 -641 85 -607
rect 33 -650 85 -641
rect 107 -607 159 -598
rect 107 -641 116 -607
rect 116 -641 150 -607
rect 150 -641 159 -607
rect 107 -650 159 -641
rect 181 -607 233 -598
rect 181 -641 190 -607
rect 190 -641 224 -607
rect 224 -641 233 -607
rect 181 -650 233 -641
rect 255 -607 307 -598
rect 255 -641 264 -607
rect 264 -641 298 -607
rect 298 -641 307 -607
rect 255 -650 307 -641
rect 329 -607 381 -598
rect 329 -641 338 -607
rect 338 -641 372 -607
rect 372 -641 381 -607
rect 329 -650 381 -641
rect 403 -607 455 -598
rect 403 -641 412 -607
rect 412 -641 446 -607
rect 446 -641 455 -607
rect 403 -650 455 -641
rect 477 -607 529 -598
rect 477 -641 486 -607
rect 486 -641 520 -607
rect 520 -641 529 -607
rect 477 -650 529 -641
<< metal2 >>
rect 22 5939 278 5945
rect 22 63 28 5939
rect 272 63 278 5939
rect 22 57 278 63
rect -209 -450 555 -443
rect -209 -502 -189 -450
rect -137 -502 -115 -450
rect -63 -502 -41 -450
rect 11 -502 33 -450
rect 85 -502 107 -450
rect 159 -502 181 -450
rect 233 -502 255 -450
rect 307 -502 329 -450
rect 381 -502 403 -450
rect 455 -502 477 -450
rect 529 -502 555 -450
rect -209 -524 555 -502
rect -209 -576 -189 -524
rect -137 -576 -115 -524
rect -63 -576 -41 -524
rect 11 -576 33 -524
rect 85 -576 107 -524
rect 159 -576 181 -524
rect 233 -576 255 -524
rect 307 -576 329 -524
rect 381 -576 403 -524
rect 455 -576 477 -524
rect 529 -576 555 -524
rect -209 -598 555 -576
rect -209 -650 -189 -598
rect -137 -650 -115 -598
rect -63 -650 -41 -598
rect 11 -650 33 -598
rect 85 -650 107 -598
rect 159 -650 181 -598
rect 233 -650 255 -598
rect 307 -650 329 -598
rect 381 -650 403 -598
rect 455 -650 477 -598
rect 529 -650 555 -598
rect -209 -657 555 -650
<< labels >>
flabel comment s -766 250 -766 250 0 FreeSans 1600 0 0 0 S
flabel comment s 1063 250 1063 250 0 FreeSans 1600 0 0 0 S
flabel comment s 150 233 150 233 0 FreeSans 1600 0 0 0 D
<< properties >>
string GDS_END 8212716
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7971364
<< end >>
