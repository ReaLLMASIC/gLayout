magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -119 -66 975 1466
<< mvpmos >>
rect 0 0 400 1400
rect 456 0 856 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 856 0 906 1400
<< poly >>
rect 0 1400 400 1426
rect 0 -26 400 0
rect 456 1400 856 1426
rect 456 -26 856 0
<< locali >>
rect -45 -4 -11 1354
rect 411 -4 445 1354
rect 867 -4 901 1354
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_0
timestamp 1701704242
transform -1 0 0 0 1 0
box -36 -36 89 1436
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_1
timestamp 1701704242
transform 1 0 856 0 1 0
box -36 -36 89 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_0
timestamp 1701704242
transform 1 0 400 0 1 0
box -36 -36 92 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 428 675 428 675 0 FreeSans 300 0 0 0 D
flabel comment s 884 675 884 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 78918202
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78916690
<< end >>
