magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -66 377 2274 897
<< pwell >>
rect 1928 281 2186 283
rect 1604 269 2186 281
rect 32 242 610 269
rect 1040 242 2186 269
rect 32 43 2186 242
rect -26 -43 2234 43
<< mvnmos >>
rect 119 159 219 243
rect 275 159 375 243
rect 431 159 531 243
rect 697 132 797 216
rect 853 132 953 216
rect 1119 159 1219 243
rect 1261 159 1361 243
rect 1417 159 1517 243
rect 1683 171 1783 255
rect 1839 171 1939 255
rect 2007 107 2107 257
<< mvpmos >>
rect 119 457 219 607
rect 275 457 375 607
rect 431 457 531 607
rect 697 457 797 607
rect 853 457 953 607
rect 1119 457 1219 541
rect 1261 457 1361 541
rect 1417 457 1517 541
rect 1683 443 1783 593
rect 1839 443 1939 593
rect 2007 443 2107 743
<< mvndiff >>
rect 58 218 119 243
rect 58 184 74 218
rect 108 184 119 218
rect 58 159 119 184
rect 219 201 275 243
rect 219 167 230 201
rect 264 167 275 201
rect 219 159 275 167
rect 375 218 431 243
rect 375 184 386 218
rect 420 184 431 218
rect 375 159 431 184
rect 531 218 584 243
rect 531 184 542 218
rect 576 184 584 218
rect 531 159 584 184
rect 1954 255 2007 257
rect 1066 218 1119 243
rect 644 191 697 216
rect 644 157 652 191
rect 686 157 697 191
rect 644 132 697 157
rect 797 191 853 216
rect 797 157 808 191
rect 842 157 853 191
rect 797 132 853 157
rect 953 191 1006 216
rect 953 157 964 191
rect 998 157 1006 191
rect 1066 184 1074 218
rect 1108 184 1119 218
rect 1066 159 1119 184
rect 1219 159 1261 243
rect 1361 205 1417 243
rect 1361 171 1372 205
rect 1406 171 1417 205
rect 1361 159 1417 171
rect 1517 218 1570 243
rect 1517 184 1528 218
rect 1562 184 1570 218
rect 1517 159 1570 184
rect 1630 227 1683 255
rect 1630 193 1638 227
rect 1672 193 1683 227
rect 1630 171 1683 193
rect 1783 171 1839 255
rect 1939 235 2007 255
rect 1939 201 1962 235
rect 1996 201 2007 235
rect 1939 171 2007 201
rect 953 132 1006 157
rect 1954 153 2007 171
rect 1954 119 1962 153
rect 1996 119 2007 153
rect 1954 107 2007 119
rect 2107 227 2160 257
rect 2107 193 2118 227
rect 2152 193 2160 227
rect 2107 153 2160 193
rect 2107 119 2118 153
rect 2152 119 2160 153
rect 2107 107 2160 119
<< mvpdiff >>
rect 1954 731 2007 743
rect 58 595 119 607
rect 58 561 74 595
rect 108 561 119 595
rect 58 503 119 561
rect 58 469 74 503
rect 108 469 119 503
rect 58 457 119 469
rect 219 457 275 607
rect 375 595 431 607
rect 375 561 386 595
rect 420 561 431 595
rect 375 503 431 561
rect 375 469 386 503
rect 420 469 431 503
rect 375 457 431 469
rect 531 595 584 607
rect 531 561 542 595
rect 576 561 584 595
rect 531 503 584 561
rect 531 469 542 503
rect 576 469 584 503
rect 531 457 584 469
rect 644 595 697 607
rect 644 561 652 595
rect 686 561 697 595
rect 644 503 697 561
rect 644 469 652 503
rect 686 469 697 503
rect 644 457 697 469
rect 797 599 853 607
rect 797 565 808 599
rect 842 565 853 599
rect 797 531 853 565
rect 797 497 808 531
rect 842 497 853 531
rect 797 457 853 497
rect 953 595 1006 607
rect 953 561 964 595
rect 998 561 1006 595
rect 953 503 1006 561
rect 953 469 964 503
rect 998 469 1006 503
rect 953 457 1006 469
rect 1954 697 1962 731
rect 1996 697 2007 731
rect 1954 663 2007 697
rect 1954 629 1962 663
rect 1996 629 2007 663
rect 1954 593 2007 629
rect 1630 581 1683 593
rect 1630 547 1638 581
rect 1672 547 1683 581
rect 1066 516 1119 541
rect 1066 482 1074 516
rect 1108 482 1119 516
rect 1066 457 1119 482
rect 1219 457 1261 541
rect 1361 516 1417 541
rect 1361 482 1372 516
rect 1406 482 1417 516
rect 1361 457 1417 482
rect 1517 516 1570 541
rect 1517 482 1528 516
rect 1562 482 1570 516
rect 1517 457 1570 482
rect 1630 489 1683 547
rect 1630 455 1638 489
rect 1672 455 1683 489
rect 1630 443 1683 455
rect 1783 575 1839 593
rect 1783 541 1794 575
rect 1828 541 1839 575
rect 1783 489 1839 541
rect 1783 455 1794 489
rect 1828 455 1839 489
rect 1783 443 1839 455
rect 1939 557 2007 593
rect 1939 523 1962 557
rect 1996 523 2007 557
rect 1939 489 2007 523
rect 1939 455 1962 489
rect 1996 455 2007 489
rect 1939 443 2007 455
rect 2107 731 2160 743
rect 2107 697 2118 731
rect 2152 697 2160 731
rect 2107 663 2160 697
rect 2107 629 2118 663
rect 2152 629 2160 663
rect 2107 557 2160 629
rect 2107 523 2118 557
rect 2152 523 2160 557
rect 2107 489 2160 523
rect 2107 455 2118 489
rect 2152 455 2160 489
rect 2107 443 2160 455
<< mvndiffc >>
rect 74 184 108 218
rect 230 167 264 201
rect 386 184 420 218
rect 542 184 576 218
rect 652 157 686 191
rect 808 157 842 191
rect 964 157 998 191
rect 1074 184 1108 218
rect 1372 171 1406 205
rect 1528 184 1562 218
rect 1638 193 1672 227
rect 1962 201 1996 235
rect 1962 119 1996 153
rect 2118 193 2152 227
rect 2118 119 2152 153
<< mvpdiffc >>
rect 74 561 108 595
rect 74 469 108 503
rect 386 561 420 595
rect 386 469 420 503
rect 542 561 576 595
rect 542 469 576 503
rect 652 561 686 595
rect 652 469 686 503
rect 808 565 842 599
rect 808 497 842 531
rect 964 561 998 595
rect 964 469 998 503
rect 1962 697 1996 731
rect 1962 629 1996 663
rect 1638 547 1672 581
rect 1074 482 1108 516
rect 1372 482 1406 516
rect 1528 482 1562 516
rect 1638 455 1672 489
rect 1794 541 1828 575
rect 1794 455 1828 489
rect 1962 523 1996 557
rect 1962 455 1996 489
rect 2118 697 2152 731
rect 2118 629 2152 663
rect 2118 523 2152 557
rect 2118 455 2152 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
<< poly >>
rect 2007 743 2107 769
rect 431 689 565 705
rect 431 655 447 689
rect 481 655 515 689
rect 549 655 565 689
rect 431 639 565 655
rect 1021 701 1299 731
rect 119 607 219 633
rect 275 607 375 633
rect 431 607 531 639
rect 697 607 797 633
rect 853 607 953 633
rect 119 409 219 457
rect 119 375 135 409
rect 169 375 219 409
rect 119 341 219 375
rect 119 307 135 341
rect 169 307 219 341
rect 119 243 219 307
rect 275 409 375 457
rect 431 431 531 457
rect 275 375 311 409
rect 345 375 375 409
rect 697 377 797 457
rect 275 341 375 375
rect 275 307 311 341
rect 345 307 375 341
rect 495 361 629 377
rect 495 327 511 361
rect 545 327 579 361
rect 613 327 629 361
rect 495 311 629 327
rect 275 243 375 307
rect 431 243 531 269
rect 119 133 219 159
rect 275 133 375 159
rect 431 137 531 159
rect 423 121 557 137
rect 423 87 439 121
rect 473 87 507 121
rect 541 87 557 121
rect 423 71 557 87
rect 599 64 629 311
rect 697 343 736 377
rect 770 343 797 377
rect 697 309 797 343
rect 697 275 736 309
rect 770 275 797 309
rect 697 216 797 275
rect 853 442 953 457
rect 1021 442 1051 701
rect 1269 691 1299 701
rect 1269 675 1905 691
rect 1269 661 1855 675
rect 1093 643 1227 659
rect 1093 609 1109 643
rect 1143 609 1177 643
rect 1211 609 1227 643
rect 1839 641 1855 661
rect 1889 641 1905 675
rect 1839 619 1905 641
rect 1093 593 1227 609
rect 1683 593 1783 619
rect 1839 593 1939 619
rect 1119 541 1219 593
rect 1261 541 1361 567
rect 1417 541 1517 567
rect 853 412 1051 442
rect 1119 431 1219 457
rect 1261 431 1361 457
rect 853 395 953 412
rect 853 361 880 395
rect 914 361 953 395
rect 1295 409 1361 431
rect 853 327 953 361
rect 853 293 880 327
rect 914 293 953 327
rect 853 216 953 293
rect 1119 373 1253 389
rect 1119 339 1135 373
rect 1169 339 1203 373
rect 1237 339 1253 373
rect 1119 323 1253 339
rect 1295 375 1311 409
rect 1345 375 1361 409
rect 1295 341 1361 375
rect 1119 243 1219 323
rect 1295 307 1311 341
rect 1345 307 1361 341
rect 1295 269 1361 307
rect 1261 243 1361 269
rect 1417 315 1517 457
rect 1417 281 1433 315
rect 1467 281 1517 315
rect 1417 243 1517 281
rect 1683 395 1783 443
rect 1683 361 1699 395
rect 1733 361 1783 395
rect 1683 327 1783 361
rect 1683 293 1699 327
rect 1733 293 1783 327
rect 1683 255 1783 293
rect 1839 395 1939 443
rect 1839 361 1878 395
rect 1912 361 1939 395
rect 1839 255 1939 361
rect 2007 345 2107 443
rect 1981 329 2115 345
rect 1981 295 1997 329
rect 2031 295 2065 329
rect 2099 295 2115 329
rect 1981 279 2115 295
rect 2007 257 2107 279
rect 1119 133 1219 159
rect 1261 133 1361 159
rect 1417 137 1517 159
rect 1683 145 1783 171
rect 1839 145 1939 171
rect 697 106 797 132
rect 853 106 953 132
rect 1417 121 1574 137
rect 1011 99 1077 115
rect 1011 65 1027 99
rect 1061 91 1077 99
rect 1417 91 1456 121
rect 1061 87 1456 91
rect 1490 87 1524 121
rect 1558 87 1574 121
rect 1061 71 1574 87
rect 2007 81 2107 107
rect 1061 65 1447 71
rect 1011 64 1447 65
rect 599 61 1447 64
rect 599 49 1077 61
rect 599 34 1041 49
<< polycont >>
rect 447 655 481 689
rect 515 655 549 689
rect 135 375 169 409
rect 135 307 169 341
rect 311 375 345 409
rect 311 307 345 341
rect 511 327 545 361
rect 579 327 613 361
rect 439 87 473 121
rect 507 87 541 121
rect 736 343 770 377
rect 736 275 770 309
rect 1109 609 1143 643
rect 1177 609 1211 643
rect 1855 641 1889 675
rect 880 361 914 395
rect 880 293 914 327
rect 1135 339 1169 373
rect 1203 339 1237 373
rect 1311 375 1345 409
rect 1311 307 1345 341
rect 1433 281 1467 315
rect 1699 361 1733 395
rect 1699 293 1733 327
rect 1878 361 1912 395
rect 1997 295 2031 329
rect 2065 295 2099 329
rect 1027 65 1061 99
rect 1456 87 1490 121
rect 1524 87 1558 121
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
rect 58 757 858 763
rect 58 729 364 757
rect 58 695 76 729
rect 110 695 148 729
rect 182 695 220 729
rect 254 695 292 729
rect 326 723 364 729
rect 398 723 436 757
rect 470 723 508 757
rect 542 723 591 757
rect 625 723 663 757
rect 697 729 858 757
rect 697 723 735 729
rect 326 695 397 723
rect 58 689 397 695
rect 725 695 735 723
rect 769 695 807 729
rect 841 695 858 729
rect 1329 757 2084 763
rect 1329 743 1831 757
rect 1329 729 1479 743
rect 725 689 858 695
rect 58 595 124 689
rect 431 655 447 689
rect 481 655 515 689
rect 549 655 691 689
rect 431 645 691 655
rect 58 561 74 595
rect 108 561 124 595
rect 58 503 124 561
rect 58 469 74 503
rect 108 469 124 503
rect 58 459 124 469
rect 370 595 429 611
rect 370 561 386 595
rect 420 561 429 595
rect 370 503 429 561
rect 370 469 386 503
rect 420 469 429 503
rect 370 459 429 469
rect 119 409 185 425
rect 119 375 135 409
rect 169 375 185 409
rect 119 341 185 375
rect 119 307 135 341
rect 169 307 185 341
rect 295 409 361 425
rect 295 375 311 409
rect 345 375 361 409
rect 295 341 361 375
rect 295 307 311 341
rect 345 307 361 341
rect 395 273 429 459
rect 526 595 592 611
rect 526 561 542 595
rect 576 561 592 595
rect 526 503 592 561
rect 526 469 542 503
rect 576 469 592 503
rect 526 377 592 469
rect 647 595 691 645
rect 647 561 652 595
rect 686 561 691 595
rect 647 503 691 561
rect 647 469 652 503
rect 686 469 691 503
rect 792 599 858 689
rect 792 565 808 599
rect 842 565 858 599
rect 792 531 858 565
rect 792 497 808 531
rect 842 497 858 531
rect 896 677 1295 711
rect 1329 695 1335 729
rect 1369 695 1407 729
rect 1441 709 1479 729
rect 1513 709 1551 743
rect 1585 729 1831 743
rect 1585 709 1623 729
rect 1441 695 1623 709
rect 1657 695 1695 729
rect 1729 723 1831 729
rect 1865 723 1903 757
rect 1937 731 2084 757
rect 1937 723 1962 731
rect 1996 729 2084 731
rect 1729 695 1805 723
rect 1329 689 1805 695
rect 1946 697 1962 723
rect 1946 695 1975 697
rect 2009 695 2047 729
rect 2081 695 2084 729
rect 1946 689 2084 695
rect 2118 731 2191 747
rect 2152 697 2191 731
rect 647 463 691 469
rect 896 463 930 677
rect 647 429 930 463
rect 964 609 1109 643
rect 1143 609 1177 643
rect 1211 609 1227 643
rect 964 601 1227 609
rect 964 595 1006 601
rect 998 561 1006 595
rect 964 503 1006 561
rect 998 469 1006 503
rect 511 361 613 377
rect 545 327 579 361
rect 511 311 613 327
rect 58 239 429 273
rect 58 218 124 239
rect 58 184 74 218
rect 108 184 124 218
rect 370 218 429 239
rect 58 168 124 184
rect 214 201 280 205
rect 214 167 230 201
rect 264 167 280 201
rect 370 184 386 218
rect 420 184 429 218
rect 370 168 429 184
rect 526 218 592 311
rect 526 184 542 218
rect 576 184 592 218
rect 647 216 686 429
rect 526 168 592 184
rect 636 191 686 216
rect 214 125 280 167
rect 636 157 652 191
rect 636 141 686 157
rect 720 377 786 393
rect 720 343 736 377
rect 770 343 786 377
rect 720 309 786 343
rect 720 275 736 309
rect 770 275 786 309
rect 864 361 880 395
rect 914 361 930 395
rect 864 327 930 361
rect 864 293 880 327
rect 914 293 930 327
rect 720 259 786 275
rect 964 259 1006 469
rect 720 225 1006 259
rect 146 119 348 125
rect 146 85 158 119
rect 192 85 230 119
rect 264 85 302 119
rect 336 85 348 119
rect 146 73 348 85
rect 423 121 565 134
rect 423 87 439 121
rect 473 87 507 121
rect 541 107 565 121
rect 720 107 754 225
rect 956 191 1006 225
rect 541 87 754 107
rect 423 73 754 87
rect 788 157 808 191
rect 842 157 858 191
rect 788 125 858 157
rect 956 157 964 191
rect 998 157 1006 191
rect 956 141 1006 157
rect 1067 516 1124 532
rect 1261 519 1295 677
rect 1067 482 1074 516
rect 1108 482 1124 516
rect 1067 466 1124 482
rect 1219 485 1295 519
rect 1356 516 1422 689
rect 1622 581 1688 689
rect 1839 675 1912 689
rect 1839 641 1855 675
rect 1889 641 1912 675
rect 1839 625 1912 641
rect 1622 547 1638 581
rect 1672 547 1688 581
rect 1067 273 1101 466
rect 1219 389 1253 485
rect 1356 482 1372 516
rect 1406 482 1422 516
rect 1356 466 1422 482
rect 1524 516 1578 532
rect 1524 482 1528 516
rect 1562 482 1578 516
rect 1524 417 1578 482
rect 1622 489 1688 547
rect 1622 455 1638 489
rect 1672 455 1688 489
rect 1622 445 1688 455
rect 1783 575 1828 591
rect 1783 541 1794 575
rect 1783 489 1828 541
rect 1783 455 1794 489
rect 1135 373 1253 389
rect 1169 339 1203 373
rect 1237 339 1253 373
rect 1135 323 1253 339
rect 1295 409 1578 417
rect 1295 375 1311 409
rect 1345 375 1578 409
rect 1295 341 1361 375
rect 1295 307 1311 341
rect 1345 307 1361 341
rect 1524 365 1578 375
rect 1683 395 1749 411
rect 1683 365 1699 395
rect 1524 361 1699 365
rect 1733 361 1749 395
rect 1417 315 1490 331
rect 1417 281 1433 315
rect 1467 281 1490 315
rect 1417 273 1490 281
rect 1067 239 1490 273
rect 1067 218 1124 239
rect 1067 184 1074 218
rect 1108 184 1124 218
rect 788 119 922 125
rect 788 85 791 119
rect 825 85 863 119
rect 897 107 922 119
rect 1067 107 1124 184
rect 1356 171 1372 205
rect 1406 171 1422 205
rect 1356 125 1422 171
rect 897 105 977 107
rect 897 85 935 105
rect 788 71 935 85
rect 969 71 977 105
rect 788 51 977 71
rect 1011 99 1124 107
rect 1011 65 1027 99
rect 1061 65 1124 99
rect 1011 51 1124 65
rect 1158 119 1422 125
rect 1158 105 1310 119
rect 1158 71 1166 105
rect 1200 71 1238 105
rect 1272 85 1310 105
rect 1344 85 1382 119
rect 1416 85 1422 119
rect 1272 71 1422 85
rect 1456 134 1490 239
rect 1524 327 1749 361
rect 1524 323 1699 327
rect 1524 218 1578 323
rect 1683 293 1699 323
rect 1733 293 1749 327
rect 1683 277 1749 293
rect 1783 311 1828 455
rect 1862 405 1912 625
rect 1946 663 2012 689
rect 1946 629 1962 663
rect 1996 629 2012 663
rect 1946 557 2012 629
rect 1946 523 1962 557
rect 1996 523 2012 557
rect 1946 489 2012 523
rect 1946 455 1962 489
rect 1996 455 2012 489
rect 1946 439 2012 455
rect 2118 663 2191 697
rect 2152 629 2191 663
rect 2118 557 2191 629
rect 2152 523 2191 557
rect 2118 489 2191 523
rect 2152 455 2191 489
rect 1862 395 1928 405
rect 1862 361 1878 395
rect 1912 361 1928 395
rect 2118 379 2191 455
rect 1862 345 1928 361
rect 1981 329 2103 345
rect 1981 311 1997 329
rect 1783 295 1997 311
rect 2031 295 2065 329
rect 2099 295 2103 329
rect 1783 277 2103 295
rect 1783 243 1828 277
rect 2137 243 2191 379
rect 1524 184 1528 218
rect 1562 184 1578 218
rect 1524 168 1578 184
rect 1622 227 1828 243
rect 1622 193 1638 227
rect 1672 193 1828 227
rect 1622 177 1828 193
rect 1946 235 2012 243
rect 1946 201 1962 235
rect 1996 201 2012 235
rect 1946 153 2012 201
rect 1456 121 1574 134
rect 1946 125 1962 153
rect 1490 87 1524 121
rect 1558 87 1574 121
rect 1456 71 1574 87
rect 1608 119 1962 125
rect 1996 125 2012 153
rect 2118 227 2191 243
rect 2152 193 2191 227
rect 2118 153 2191 193
rect 1996 119 2084 125
rect 1608 105 1900 119
rect 1608 71 1612 105
rect 1646 71 1684 105
rect 1718 71 1756 105
rect 1790 71 1828 105
rect 1862 85 1900 105
rect 1934 85 1972 119
rect 2006 85 2044 119
rect 2078 85 2084 119
rect 2152 119 2191 153
rect 2118 103 2191 119
rect 1862 71 2084 85
rect 1158 51 1422 71
rect 1608 51 2084 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 76 695 110 729
rect 148 695 182 729
rect 220 695 254 729
rect 292 695 326 729
rect 364 723 398 757
rect 436 723 470 757
rect 508 723 542 757
rect 591 723 625 757
rect 663 723 697 757
rect 735 695 769 729
rect 807 695 841 729
rect 1335 695 1369 729
rect 1407 695 1441 729
rect 1479 709 1513 743
rect 1551 709 1585 743
rect 1623 695 1657 729
rect 1695 695 1729 729
rect 1831 723 1865 757
rect 1903 723 1937 757
rect 1975 697 1996 729
rect 1996 697 2009 729
rect 1975 695 2009 697
rect 2047 695 2081 729
rect 158 85 192 119
rect 230 85 264 119
rect 302 85 336 119
rect 791 85 825 119
rect 863 85 897 119
rect 935 71 969 105
rect 1166 71 1200 105
rect 1238 71 1272 105
rect 1310 85 1344 119
rect 1382 85 1416 119
rect 1612 71 1646 105
rect 1684 71 1718 105
rect 1756 71 1790 105
rect 1828 71 1862 105
rect 1900 85 1934 119
rect 1972 85 2006 119
rect 2044 85 2078 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 831 2208 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
rect 0 791 2208 797
rect 0 757 2208 763
rect 0 729 364 757
rect 0 695 76 729
rect 110 695 148 729
rect 182 695 220 729
rect 254 695 292 729
rect 326 723 364 729
rect 398 723 436 757
rect 470 723 508 757
rect 542 723 591 757
rect 625 723 663 757
rect 697 743 1831 757
rect 697 729 1479 743
rect 697 723 735 729
rect 326 695 735 723
rect 769 695 807 729
rect 841 695 1335 729
rect 1369 695 1407 729
rect 1441 709 1479 729
rect 1513 709 1551 743
rect 1585 729 1831 743
rect 1585 709 1623 729
rect 1441 695 1623 709
rect 1657 695 1695 729
rect 1729 723 1831 729
rect 1865 723 1903 757
rect 1937 729 2208 757
rect 1937 723 1975 729
rect 1729 695 1975 723
rect 2009 695 2047 729
rect 2081 695 2208 729
rect 0 689 2208 695
rect 0 119 2208 125
rect 0 85 158 119
rect 192 85 230 119
rect 264 85 302 119
rect 336 85 791 119
rect 825 85 863 119
rect 897 105 1310 119
rect 897 85 935 105
rect 0 71 935 85
rect 969 71 1166 105
rect 1200 71 1238 105
rect 1272 85 1310 105
rect 1344 85 1382 119
rect 1416 105 1900 119
rect 1416 85 1612 105
rect 1272 71 1612 85
rect 1646 71 1684 105
rect 1718 71 1756 105
rect 1790 71 1828 105
rect 1862 85 1900 105
rect 1934 85 1972 119
rect 2006 85 2044 119
rect 2078 85 2208 119
rect 1862 71 2208 85
rect 0 51 2208 71
rect 0 17 2208 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -23 2208 -17
<< labels >>
flabel comment s 1170 303 1170 303 0 FreeSans 200 0 0 0 clkneg
flabel comment s 748 234 748 234 0 FreeSans 200 0 0 0 clkpos
flabel comment s 1170 446 1170 446 0 FreeSans 200 0 0 0 clkpos
rlabel comment s 0 0 0 0 4 dlclkp_1
flabel comment s 666 352 666 352 0 FreeSans 200 90 0 0 clkneg
flabel comment s 482 259 482 259 0 FreeSans 200 0 0 0 clkpos
flabel comment s 978 352 978 352 0 FreeSans 200 90 0 0 clkpos
flabel comment s 482 446 482 446 0 FreeSans 200 0 0 0 clkneg
flabel comment s 807 51 807 51 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 51 2208 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 2208 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 2208 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 2208 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 2143 242 2177 276 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2208 814
string GDS_END 695048
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 672184
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
