magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 640 203
rect 29 -17 63 21
<< scnmos >>
rect 82 47 112 177
rect 154 47 184 177
rect 364 47 394 177
rect 448 47 478 177
rect 532 47 562 177
<< scpmoshvt >>
rect 82 297 112 497
rect 166 297 196 497
rect 364 297 394 497
rect 448 297 478 497
rect 532 297 562 497
<< ndiff >>
rect 27 163 82 177
rect 27 129 35 163
rect 69 129 82 163
rect 27 95 82 129
rect 27 61 35 95
rect 69 61 82 95
rect 27 47 82 61
rect 112 47 154 177
rect 184 163 258 177
rect 184 129 216 163
rect 250 129 258 163
rect 184 95 258 129
rect 184 61 216 95
rect 250 61 258 95
rect 184 47 258 61
rect 312 138 364 177
rect 312 104 320 138
rect 354 104 364 138
rect 312 47 364 104
rect 394 138 448 177
rect 394 104 404 138
rect 438 104 448 138
rect 394 47 448 104
rect 478 95 532 177
rect 478 61 488 95
rect 522 61 532 95
rect 478 47 532 61
rect 562 163 614 177
rect 562 129 572 163
rect 606 129 614 163
rect 562 95 614 129
rect 562 61 572 95
rect 606 61 614 95
rect 562 47 614 61
<< pdiff >>
rect 27 479 82 497
rect 27 445 38 479
rect 72 445 82 479
rect 27 411 82 445
rect 27 377 38 411
rect 72 377 82 411
rect 27 343 82 377
rect 27 309 38 343
rect 72 309 82 343
rect 27 297 82 309
rect 112 477 166 497
rect 112 443 122 477
rect 156 443 166 477
rect 112 409 166 443
rect 112 375 122 409
rect 156 375 166 409
rect 112 297 166 375
rect 196 477 364 497
rect 196 443 214 477
rect 248 443 304 477
rect 338 443 364 477
rect 196 409 364 443
rect 196 375 214 409
rect 248 375 304 409
rect 338 375 364 409
rect 196 297 364 375
rect 394 477 448 497
rect 394 443 404 477
rect 438 443 448 477
rect 394 409 448 443
rect 394 375 404 409
rect 438 375 448 409
rect 394 341 448 375
rect 394 307 404 341
rect 438 307 448 341
rect 394 297 448 307
rect 478 297 532 497
rect 562 479 617 497
rect 562 445 572 479
rect 606 445 617 479
rect 562 411 617 445
rect 562 377 572 411
rect 606 377 617 411
rect 562 343 617 377
rect 562 309 572 343
rect 606 309 617 343
rect 562 297 617 309
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 216 129 250 163
rect 216 61 250 95
rect 320 104 354 138
rect 404 104 438 138
rect 488 61 522 95
rect 572 129 606 163
rect 572 61 606 95
<< pdiffc >>
rect 38 445 72 479
rect 38 377 72 411
rect 38 309 72 343
rect 122 443 156 477
rect 122 375 156 409
rect 214 443 248 477
rect 304 443 338 477
rect 214 375 248 409
rect 304 375 338 409
rect 404 443 438 477
rect 404 375 438 409
rect 404 307 438 341
rect 572 445 606 479
rect 572 377 606 411
rect 572 309 606 343
<< poly >>
rect 82 497 112 523
rect 166 497 196 523
rect 364 497 394 523
rect 448 497 478 523
rect 532 497 562 523
rect 82 265 112 297
rect 166 265 196 297
rect 364 265 394 297
rect 448 265 478 297
rect 532 265 562 297
rect 21 249 112 265
rect 21 215 37 249
rect 71 215 112 249
rect 21 199 112 215
rect 82 177 112 199
rect 154 249 208 265
rect 154 215 164 249
rect 198 215 208 249
rect 154 199 208 215
rect 250 249 394 265
rect 250 215 260 249
rect 294 215 394 249
rect 250 199 394 215
rect 436 249 490 265
rect 436 215 446 249
rect 480 215 490 249
rect 436 199 490 215
rect 532 249 623 265
rect 532 215 573 249
rect 607 215 623 249
rect 532 199 623 215
rect 154 177 184 199
rect 364 177 394 199
rect 448 177 478 199
rect 532 177 562 199
rect 82 21 112 47
rect 154 21 184 47
rect 364 21 394 47
rect 448 21 478 47
rect 532 21 562 47
<< polycont >>
rect 37 215 71 249
rect 164 215 198 249
rect 260 215 294 249
rect 446 215 480 249
rect 573 215 607 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 30 479 80 527
rect 30 445 38 479
rect 72 445 80 479
rect 30 411 80 445
rect 30 377 38 411
rect 72 377 80 411
rect 30 343 80 377
rect 30 309 38 343
rect 72 309 80 343
rect 30 291 80 309
rect 114 477 164 493
rect 114 443 122 477
rect 156 443 164 477
rect 114 409 164 443
rect 114 375 122 409
rect 156 375 164 409
rect 114 333 164 375
rect 198 477 354 527
rect 198 443 214 477
rect 248 443 304 477
rect 338 443 354 477
rect 198 409 354 443
rect 198 375 214 409
rect 248 375 304 409
rect 338 375 354 409
rect 198 367 354 375
rect 388 477 454 493
rect 388 443 404 477
rect 438 443 454 477
rect 388 409 454 443
rect 388 375 404 409
rect 438 375 454 409
rect 388 341 454 375
rect 388 333 404 341
rect 114 299 268 333
rect 234 265 268 299
rect 328 307 404 333
rect 438 307 454 341
rect 328 299 454 307
rect 17 249 87 257
rect 17 215 37 249
rect 71 215 87 249
rect 17 197 87 215
rect 121 249 200 265
rect 121 215 164 249
rect 198 215 200 249
rect 121 199 200 215
rect 234 249 294 265
rect 234 215 260 249
rect 234 199 294 215
rect 18 129 35 163
rect 69 129 85 163
rect 18 95 85 129
rect 18 61 35 95
rect 69 61 85 95
rect 18 17 85 61
rect 121 56 165 199
rect 234 165 268 199
rect 200 163 268 165
rect 200 129 216 163
rect 250 129 268 163
rect 328 158 362 299
rect 489 265 523 485
rect 564 479 614 527
rect 564 445 572 479
rect 606 445 614 479
rect 564 411 614 445
rect 564 377 572 411
rect 606 377 614 411
rect 564 343 614 377
rect 564 309 572 343
rect 606 309 614 343
rect 564 291 614 309
rect 406 249 523 265
rect 406 215 446 249
rect 480 215 523 249
rect 557 249 627 257
rect 557 215 573 249
rect 607 215 627 249
rect 200 95 268 129
rect 200 61 216 95
rect 250 61 268 95
rect 312 138 362 158
rect 312 104 320 138
rect 354 104 362 138
rect 312 86 362 104
rect 396 163 622 181
rect 396 145 572 163
rect 396 138 454 145
rect 396 104 404 138
rect 438 104 454 138
rect 556 129 572 145
rect 606 129 622 163
rect 396 85 454 104
rect 488 95 522 111
rect 200 56 268 61
rect 488 17 522 61
rect 556 95 622 129
rect 556 61 572 95
rect 606 61 622 95
rect 556 55 622 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 397 357 431 391 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 400 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o2bb2ai_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1236666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1230496
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
