magic
tech sky130A
magscale 1 2
timestamp 1701704242
use sky130_fd_io__amux_switch_1v2b  sky130_fd_io__amux_switch_1v2b_0
timestamp 1701704242
transform 1 0 4755 0 -1 8802
box -50 -73 10379 2429
use sky130_fd_io__amux_switch_1v2b  sky130_fd_io__amux_switch_1v2b_1
timestamp 1701704242
transform 1 0 4755 0 1 4180
box -50 -73 10379 2429
use sky130_fd_io__gpiov2_amux_ctl_logic  sky130_fd_io__gpiov2_amux_ctl_logic_0
timestamp 1701704242
transform 1 0 -26998 0 1 6306
box 26092 -15586 41870 1848
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1701704242
transform 1 0 3419 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1701704242
transform 1 0 2619 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_2
timestamp 1701704242
transform 1 0 2619 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_3
timestamp 1701704242
transform 1 0 3419 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_4
timestamp 1701704242
transform -1 0 8708 0 1 9409
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_5
timestamp 1701704242
transform 1 0 8626 0 1 9409
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_6
timestamp 1701704242
transform 0 1 12464 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_7
timestamp 1701704242
transform 0 -1 12368 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_8
timestamp 1701704242
transform 0 1 12464 -1 0 3218
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_9
timestamp 1701704242
transform 0 -1 11869 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_10
timestamp 1701704242
transform -1 0 1901 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_11
timestamp 1701704242
transform -1 0 2701 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_12
timestamp 1701704242
transform -1 0 2701 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_13
timestamp 1701704242
transform -1 0 1901 0 -1 6379
box 0 0 882 404
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_0
timestamp 1701704242
transform 1 0 14424 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_1
timestamp 1701704242
transform 1 0 13880 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_2
timestamp 1701704242
transform 1 0 13608 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_3
timestamp 1701704242
transform 1 0 14152 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_4
timestamp 1701704242
transform 1 0 13608 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_5
timestamp 1701704242
transform 1 0 14152 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_6
timestamp 1701704242
transform 1 0 14424 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_7
timestamp 1701704242
transform 1 0 13880 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_0
timestamp 1701704242
transform 1 0 13603 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_1
timestamp 1701704242
transform 1 0 14151 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_2
timestamp 1701704242
transform 1 0 14423 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_3
timestamp 1701704242
transform 1 0 13875 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808594  sky130_fd_pr__nfet_01v8__example_55959141808594_0
timestamp 1701704242
transform 0 -1 14630 -1 0 2528
box -1 0 2129 1
use sky130_fd_pr__pfet_01v8__example_55959141808591  sky130_fd_pr__pfet_01v8__example_55959141808591_0
timestamp 1701704242
transform 0 1 1282 -1 0 8427
box -1 0 1037 1
<< properties >>
string GDS_END 23026238
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22509480
<< end >>
