magic
tech sky130A
timestamp 1701704242
<< viali >>
rect 0 0 341 53
<< metal1 >>
rect -6 53 347 56
rect -6 0 0 53
rect 341 0 347 53
rect -6 -3 347 0
<< properties >>
string GDS_END 89708896
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89707484
<< end >>
