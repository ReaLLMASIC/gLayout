magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 67 368 203
rect 30 21 368 67
rect 30 -17 64 21
<< scnmos >>
rect 79 93 109 177
rect 176 47 206 177
rect 260 47 290 177
<< scpmoshvt >>
rect 79 297 109 381
rect 176 297 206 497
rect 260 297 290 497
<< ndiff >>
rect 27 155 79 177
rect 27 121 35 155
rect 69 121 79 155
rect 27 93 79 121
rect 109 93 176 177
rect 124 59 132 93
rect 166 59 176 93
rect 124 47 176 59
rect 206 47 260 177
rect 290 93 342 177
rect 290 59 300 93
rect 334 59 342 93
rect 290 47 342 59
<< pdiff >>
rect 124 485 176 497
rect 124 451 132 485
rect 166 451 176 485
rect 124 417 176 451
rect 124 383 132 417
rect 166 383 176 417
rect 124 381 176 383
rect 27 349 79 381
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 176 381
rect 206 485 260 497
rect 206 451 216 485
rect 250 451 260 485
rect 206 417 260 451
rect 206 383 216 417
rect 250 383 260 417
rect 206 297 260 383
rect 290 485 343 497
rect 290 451 300 485
rect 334 451 343 485
rect 290 297 343 451
<< ndiffc >>
rect 35 121 69 155
rect 132 59 166 93
rect 300 59 334 93
<< pdiffc >>
rect 132 451 166 485
rect 132 383 166 417
rect 35 315 69 349
rect 216 451 250 485
rect 216 383 250 417
rect 300 451 334 485
<< poly >>
rect 176 497 206 523
rect 260 497 290 523
rect 79 381 109 407
rect 79 265 109 297
rect 176 265 206 297
rect 260 265 290 297
rect 22 249 109 265
rect 22 215 38 249
rect 72 215 109 249
rect 22 199 109 215
rect 151 249 217 265
rect 151 215 167 249
rect 201 215 217 249
rect 151 199 217 215
rect 260 249 326 265
rect 260 215 276 249
rect 310 215 326 249
rect 260 199 326 215
rect 79 177 109 199
rect 176 177 206 199
rect 260 177 290 199
rect 79 67 109 93
rect 176 21 206 47
rect 260 21 290 47
<< polycont >>
rect 38 215 72 249
rect 167 215 201 249
rect 276 215 310 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 116 485 166 527
rect 116 451 132 485
rect 116 417 166 451
rect 116 383 132 417
rect 116 367 166 383
rect 200 485 266 493
rect 200 451 216 485
rect 250 451 266 485
rect 200 417 266 451
rect 300 485 343 527
rect 334 451 343 485
rect 300 435 343 451
rect 200 383 216 417
rect 250 401 266 417
rect 250 383 434 401
rect 200 367 434 383
rect 18 349 74 365
rect 18 315 35 349
rect 69 333 74 349
rect 69 315 285 333
rect 18 299 285 315
rect 251 265 285 299
rect 18 249 88 263
rect 18 215 38 249
rect 72 215 88 249
rect 122 249 217 263
rect 122 215 167 249
rect 201 215 217 249
rect 251 249 326 265
rect 251 215 276 249
rect 310 215 326 249
rect 251 181 285 215
rect 18 155 285 181
rect 18 121 35 155
rect 69 147 285 155
rect 69 121 72 147
rect 18 105 72 121
rect 360 109 434 367
rect 116 93 182 109
rect 116 59 132 93
rect 166 59 182 93
rect 116 17 182 59
rect 284 93 434 109
rect 284 59 300 93
rect 334 59 434 93
rect 284 51 434 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 397 357 431 391 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 397 289 431 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 397 85 431 119 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 397 153 431 187 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand2b_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1742060
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1737530
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
