magic
tech sky130A
timestamp 1701704242
<< nwell >>
rect -18 -18 59 297
<< nsubdiff >>
rect 0 267 41 279
rect 0 250 12 267
rect 29 250 41 267
rect 0 233 41 250
rect 0 216 12 233
rect 29 216 41 233
rect 0 199 41 216
rect 0 182 12 199
rect 29 182 41 199
rect 0 165 41 182
rect 0 148 12 165
rect 29 148 41 165
rect 0 131 41 148
rect 0 114 12 131
rect 29 114 41 131
rect 0 97 41 114
rect 0 80 12 97
rect 29 80 41 97
rect 0 63 41 80
rect 0 46 12 63
rect 29 46 41 63
rect 0 29 41 46
rect 0 12 12 29
rect 29 12 41 29
rect 0 0 41 12
<< nsubdiffcont >>
rect 12 250 29 267
rect 12 216 29 233
rect 12 182 29 199
rect 12 148 29 165
rect 12 114 29 131
rect 12 80 29 97
rect 12 46 29 63
rect 12 12 29 29
<< locali >>
rect 12 267 29 275
rect 12 233 29 250
rect 12 199 29 216
rect 12 165 29 182
rect 12 131 29 148
rect 12 97 29 114
rect 12 63 29 80
rect 12 29 29 46
rect 12 4 29 12
<< properties >>
string GDS_END 88584458
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88583686
<< end >>
