magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -66 377 3618 897
<< pwell >>
rect 4 43 3538 317
rect -26 -43 3578 43
<< mvnmos >>
rect 83 141 183 291
rect 239 141 339 291
rect 395 141 495 291
rect 551 141 651 291
rect 707 141 807 291
rect 863 141 963 291
rect 1019 141 1119 291
rect 1175 141 1275 291
rect 1331 141 1431 291
rect 1487 141 1587 291
rect 1643 141 1743 291
rect 1799 141 1899 291
rect 1955 141 2055 291
rect 2111 141 2211 291
rect 2267 141 2367 291
rect 2423 141 2523 291
rect 2579 141 2679 291
rect 2735 141 2835 291
rect 2891 141 2991 291
rect 3047 141 3147 291
rect 3203 141 3303 291
rect 3359 141 3459 291
<< mvpmos >>
rect 83 443 183 743
rect 239 443 339 743
rect 395 443 495 743
rect 551 443 651 743
rect 707 443 807 743
rect 863 443 963 743
rect 1019 443 1119 743
rect 1175 443 1275 743
rect 1331 443 1431 743
rect 1487 443 1587 743
rect 1643 443 1743 743
rect 1799 443 1899 743
rect 1955 443 2055 743
rect 2111 443 2211 743
rect 2267 443 2367 743
rect 2423 443 2523 743
rect 2579 443 2679 743
rect 2735 443 2835 743
rect 2891 443 2991 743
rect 3047 443 3147 743
rect 3203 443 3303 743
rect 3359 443 3459 743
<< mvndiff >>
rect 30 273 83 291
rect 30 239 38 273
rect 72 239 83 273
rect 30 205 83 239
rect 30 171 38 205
rect 72 171 83 205
rect 30 141 83 171
rect 183 269 239 291
rect 183 235 194 269
rect 228 235 239 269
rect 183 201 239 235
rect 183 167 194 201
rect 228 167 239 201
rect 183 141 239 167
rect 339 205 395 291
rect 339 171 350 205
rect 384 171 395 205
rect 339 141 395 171
rect 495 264 551 291
rect 495 230 506 264
rect 540 230 551 264
rect 495 196 551 230
rect 495 162 506 196
rect 540 162 551 196
rect 495 141 551 162
rect 651 205 707 291
rect 651 171 662 205
rect 696 171 707 205
rect 651 141 707 171
rect 807 264 863 291
rect 807 230 818 264
rect 852 230 863 264
rect 807 196 863 230
rect 807 162 818 196
rect 852 162 863 196
rect 807 141 863 162
rect 963 201 1019 291
rect 963 167 974 201
rect 1008 167 1019 201
rect 963 141 1019 167
rect 1119 283 1175 291
rect 1119 249 1130 283
rect 1164 249 1175 283
rect 1119 208 1175 249
rect 1119 174 1130 208
rect 1164 174 1175 208
rect 1119 141 1175 174
rect 1275 269 1331 291
rect 1275 235 1286 269
rect 1320 235 1331 269
rect 1275 201 1331 235
rect 1275 167 1286 201
rect 1320 167 1331 201
rect 1275 141 1331 167
rect 1431 283 1487 291
rect 1431 249 1442 283
rect 1476 249 1487 283
rect 1431 208 1487 249
rect 1431 174 1442 208
rect 1476 174 1487 208
rect 1431 141 1487 174
rect 1587 269 1643 291
rect 1587 235 1598 269
rect 1632 235 1643 269
rect 1587 201 1643 235
rect 1587 167 1598 201
rect 1632 167 1643 201
rect 1587 141 1643 167
rect 1743 283 1799 291
rect 1743 249 1754 283
rect 1788 249 1799 283
rect 1743 208 1799 249
rect 1743 174 1754 208
rect 1788 174 1799 208
rect 1743 141 1799 174
rect 1899 269 1955 291
rect 1899 235 1910 269
rect 1944 235 1955 269
rect 1899 201 1955 235
rect 1899 167 1910 201
rect 1944 167 1955 201
rect 1899 141 1955 167
rect 2055 283 2111 291
rect 2055 249 2066 283
rect 2100 249 2111 283
rect 2055 208 2111 249
rect 2055 174 2066 208
rect 2100 174 2111 208
rect 2055 141 2111 174
rect 2211 269 2267 291
rect 2211 235 2222 269
rect 2256 235 2267 269
rect 2211 201 2267 235
rect 2211 167 2222 201
rect 2256 167 2267 201
rect 2211 141 2267 167
rect 2367 283 2423 291
rect 2367 249 2378 283
rect 2412 249 2423 283
rect 2367 208 2423 249
rect 2367 174 2378 208
rect 2412 174 2423 208
rect 2367 141 2423 174
rect 2523 269 2579 291
rect 2523 235 2534 269
rect 2568 235 2579 269
rect 2523 201 2579 235
rect 2523 167 2534 201
rect 2568 167 2579 201
rect 2523 141 2579 167
rect 2679 283 2735 291
rect 2679 249 2690 283
rect 2724 249 2735 283
rect 2679 208 2735 249
rect 2679 174 2690 208
rect 2724 174 2735 208
rect 2679 141 2735 174
rect 2835 269 2891 291
rect 2835 235 2846 269
rect 2880 235 2891 269
rect 2835 201 2891 235
rect 2835 167 2846 201
rect 2880 167 2891 201
rect 2835 141 2891 167
rect 2991 283 3047 291
rect 2991 249 3002 283
rect 3036 249 3047 283
rect 2991 208 3047 249
rect 2991 174 3002 208
rect 3036 174 3047 208
rect 2991 141 3047 174
rect 3147 269 3203 291
rect 3147 235 3158 269
rect 3192 235 3203 269
rect 3147 201 3203 235
rect 3147 167 3158 201
rect 3192 167 3203 201
rect 3147 141 3203 167
rect 3303 283 3359 291
rect 3303 249 3314 283
rect 3348 249 3359 283
rect 3303 208 3359 249
rect 3303 174 3314 208
rect 3348 174 3359 208
rect 3303 141 3359 174
rect 3459 279 3512 291
rect 3459 245 3470 279
rect 3504 245 3512 279
rect 3459 208 3512 245
rect 3459 174 3470 208
rect 3504 174 3512 208
rect 3459 141 3512 174
<< mvpdiff >>
rect 30 731 83 743
rect 30 697 38 731
rect 72 697 83 731
rect 30 642 83 697
rect 30 608 38 642
rect 72 608 83 642
rect 30 562 83 608
rect 30 528 38 562
rect 72 528 83 562
rect 30 489 83 528
rect 30 455 38 489
rect 72 455 83 489
rect 30 443 83 455
rect 183 735 239 743
rect 183 701 194 735
rect 228 701 239 735
rect 183 642 239 701
rect 183 608 194 642
rect 228 608 239 642
rect 183 558 239 608
rect 183 524 194 558
rect 228 524 239 558
rect 183 485 239 524
rect 183 451 194 485
rect 228 451 239 485
rect 183 443 239 451
rect 339 731 395 743
rect 339 697 350 731
rect 384 697 395 731
rect 339 663 395 697
rect 339 629 350 663
rect 384 629 395 663
rect 339 595 395 629
rect 339 561 350 595
rect 384 561 395 595
rect 339 527 395 561
rect 339 493 350 527
rect 384 493 395 527
rect 339 443 395 493
rect 495 735 551 743
rect 495 701 506 735
rect 540 701 551 735
rect 495 642 551 701
rect 495 608 506 642
rect 540 608 551 642
rect 495 558 551 608
rect 495 524 506 558
rect 540 524 551 558
rect 495 485 551 524
rect 495 451 506 485
rect 540 451 551 485
rect 495 443 551 451
rect 651 731 707 743
rect 651 697 662 731
rect 696 697 707 731
rect 651 663 707 697
rect 651 629 662 663
rect 696 629 707 663
rect 651 595 707 629
rect 651 561 662 595
rect 696 561 707 595
rect 651 527 707 561
rect 651 493 662 527
rect 696 493 707 527
rect 651 443 707 493
rect 807 735 863 743
rect 807 701 818 735
rect 852 701 863 735
rect 807 642 863 701
rect 807 608 818 642
rect 852 608 863 642
rect 807 558 863 608
rect 807 524 818 558
rect 852 524 863 558
rect 807 485 863 524
rect 807 451 818 485
rect 852 451 863 485
rect 807 443 863 451
rect 963 731 1019 743
rect 963 697 974 731
rect 1008 697 1019 731
rect 963 663 1019 697
rect 963 629 974 663
rect 1008 629 1019 663
rect 963 595 1019 629
rect 963 561 974 595
rect 1008 561 1019 595
rect 963 527 1019 561
rect 963 493 974 527
rect 1008 493 1019 527
rect 963 443 1019 493
rect 1119 735 1175 743
rect 1119 701 1130 735
rect 1164 701 1175 735
rect 1119 656 1175 701
rect 1119 622 1130 656
rect 1164 622 1175 656
rect 1119 576 1175 622
rect 1119 542 1130 576
rect 1164 542 1175 576
rect 1119 485 1175 542
rect 1119 451 1130 485
rect 1164 451 1175 485
rect 1119 443 1175 451
rect 1275 735 1331 743
rect 1275 701 1286 735
rect 1320 701 1331 735
rect 1275 656 1331 701
rect 1275 622 1286 656
rect 1320 622 1331 656
rect 1275 576 1331 622
rect 1275 542 1286 576
rect 1320 542 1331 576
rect 1275 485 1331 542
rect 1275 451 1286 485
rect 1320 451 1331 485
rect 1275 443 1331 451
rect 1431 735 1487 743
rect 1431 701 1442 735
rect 1476 701 1487 735
rect 1431 656 1487 701
rect 1431 622 1442 656
rect 1476 622 1487 656
rect 1431 576 1487 622
rect 1431 542 1442 576
rect 1476 542 1487 576
rect 1431 485 1487 542
rect 1431 451 1442 485
rect 1476 451 1487 485
rect 1431 443 1487 451
rect 1587 735 1643 743
rect 1587 701 1598 735
rect 1632 701 1643 735
rect 1587 656 1643 701
rect 1587 622 1598 656
rect 1632 622 1643 656
rect 1587 576 1643 622
rect 1587 542 1598 576
rect 1632 542 1643 576
rect 1587 485 1643 542
rect 1587 451 1598 485
rect 1632 451 1643 485
rect 1587 443 1643 451
rect 1743 735 1799 743
rect 1743 701 1754 735
rect 1788 701 1799 735
rect 1743 656 1799 701
rect 1743 622 1754 656
rect 1788 622 1799 656
rect 1743 576 1799 622
rect 1743 542 1754 576
rect 1788 542 1799 576
rect 1743 485 1799 542
rect 1743 451 1754 485
rect 1788 451 1799 485
rect 1743 443 1799 451
rect 1899 735 1955 743
rect 1899 701 1910 735
rect 1944 701 1955 735
rect 1899 656 1955 701
rect 1899 622 1910 656
rect 1944 622 1955 656
rect 1899 576 1955 622
rect 1899 542 1910 576
rect 1944 542 1955 576
rect 1899 485 1955 542
rect 1899 451 1910 485
rect 1944 451 1955 485
rect 1899 443 1955 451
rect 2055 735 2111 743
rect 2055 701 2066 735
rect 2100 701 2111 735
rect 2055 656 2111 701
rect 2055 622 2066 656
rect 2100 622 2111 656
rect 2055 576 2111 622
rect 2055 542 2066 576
rect 2100 542 2111 576
rect 2055 485 2111 542
rect 2055 451 2066 485
rect 2100 451 2111 485
rect 2055 443 2111 451
rect 2211 735 2267 743
rect 2211 701 2222 735
rect 2256 701 2267 735
rect 2211 656 2267 701
rect 2211 622 2222 656
rect 2256 622 2267 656
rect 2211 576 2267 622
rect 2211 542 2222 576
rect 2256 542 2267 576
rect 2211 485 2267 542
rect 2211 451 2222 485
rect 2256 451 2267 485
rect 2211 443 2267 451
rect 2367 735 2423 743
rect 2367 701 2378 735
rect 2412 701 2423 735
rect 2367 656 2423 701
rect 2367 622 2378 656
rect 2412 622 2423 656
rect 2367 576 2423 622
rect 2367 542 2378 576
rect 2412 542 2423 576
rect 2367 485 2423 542
rect 2367 451 2378 485
rect 2412 451 2423 485
rect 2367 443 2423 451
rect 2523 735 2579 743
rect 2523 701 2534 735
rect 2568 701 2579 735
rect 2523 656 2579 701
rect 2523 622 2534 656
rect 2568 622 2579 656
rect 2523 576 2579 622
rect 2523 542 2534 576
rect 2568 542 2579 576
rect 2523 485 2579 542
rect 2523 451 2534 485
rect 2568 451 2579 485
rect 2523 443 2579 451
rect 2679 735 2735 743
rect 2679 701 2690 735
rect 2724 701 2735 735
rect 2679 656 2735 701
rect 2679 622 2690 656
rect 2724 622 2735 656
rect 2679 576 2735 622
rect 2679 542 2690 576
rect 2724 542 2735 576
rect 2679 485 2735 542
rect 2679 451 2690 485
rect 2724 451 2735 485
rect 2679 443 2735 451
rect 2835 735 2891 743
rect 2835 701 2846 735
rect 2880 701 2891 735
rect 2835 656 2891 701
rect 2835 622 2846 656
rect 2880 622 2891 656
rect 2835 576 2891 622
rect 2835 542 2846 576
rect 2880 542 2891 576
rect 2835 485 2891 542
rect 2835 451 2846 485
rect 2880 451 2891 485
rect 2835 443 2891 451
rect 2991 735 3047 743
rect 2991 701 3002 735
rect 3036 701 3047 735
rect 2991 656 3047 701
rect 2991 622 3002 656
rect 3036 622 3047 656
rect 2991 576 3047 622
rect 2991 542 3002 576
rect 3036 542 3047 576
rect 2991 485 3047 542
rect 2991 451 3002 485
rect 3036 451 3047 485
rect 2991 443 3047 451
rect 3147 735 3203 743
rect 3147 701 3158 735
rect 3192 701 3203 735
rect 3147 656 3203 701
rect 3147 622 3158 656
rect 3192 622 3203 656
rect 3147 576 3203 622
rect 3147 542 3158 576
rect 3192 542 3203 576
rect 3147 485 3203 542
rect 3147 451 3158 485
rect 3192 451 3203 485
rect 3147 443 3203 451
rect 3303 735 3359 743
rect 3303 701 3314 735
rect 3348 701 3359 735
rect 3303 656 3359 701
rect 3303 622 3314 656
rect 3348 622 3359 656
rect 3303 576 3359 622
rect 3303 542 3314 576
rect 3348 542 3359 576
rect 3303 485 3359 542
rect 3303 451 3314 485
rect 3348 451 3359 485
rect 3303 443 3359 451
rect 3459 731 3512 743
rect 3459 697 3470 731
rect 3504 697 3512 731
rect 3459 656 3512 697
rect 3459 622 3470 656
rect 3504 622 3512 656
rect 3459 576 3512 622
rect 3459 542 3470 576
rect 3504 542 3512 576
rect 3459 489 3512 542
rect 3459 455 3470 489
rect 3504 455 3512 489
rect 3459 443 3512 455
<< mvndiffc >>
rect 38 239 72 273
rect 38 171 72 205
rect 194 235 228 269
rect 194 167 228 201
rect 350 171 384 205
rect 506 230 540 264
rect 506 162 540 196
rect 662 171 696 205
rect 818 230 852 264
rect 818 162 852 196
rect 974 167 1008 201
rect 1130 249 1164 283
rect 1130 174 1164 208
rect 1286 235 1320 269
rect 1286 167 1320 201
rect 1442 249 1476 283
rect 1442 174 1476 208
rect 1598 235 1632 269
rect 1598 167 1632 201
rect 1754 249 1788 283
rect 1754 174 1788 208
rect 1910 235 1944 269
rect 1910 167 1944 201
rect 2066 249 2100 283
rect 2066 174 2100 208
rect 2222 235 2256 269
rect 2222 167 2256 201
rect 2378 249 2412 283
rect 2378 174 2412 208
rect 2534 235 2568 269
rect 2534 167 2568 201
rect 2690 249 2724 283
rect 2690 174 2724 208
rect 2846 235 2880 269
rect 2846 167 2880 201
rect 3002 249 3036 283
rect 3002 174 3036 208
rect 3158 235 3192 269
rect 3158 167 3192 201
rect 3314 249 3348 283
rect 3314 174 3348 208
rect 3470 245 3504 279
rect 3470 174 3504 208
<< mvpdiffc >>
rect 38 697 72 731
rect 38 608 72 642
rect 38 528 72 562
rect 38 455 72 489
rect 194 701 228 735
rect 194 608 228 642
rect 194 524 228 558
rect 194 451 228 485
rect 350 697 384 731
rect 350 629 384 663
rect 350 561 384 595
rect 350 493 384 527
rect 506 701 540 735
rect 506 608 540 642
rect 506 524 540 558
rect 506 451 540 485
rect 662 697 696 731
rect 662 629 696 663
rect 662 561 696 595
rect 662 493 696 527
rect 818 701 852 735
rect 818 608 852 642
rect 818 524 852 558
rect 818 451 852 485
rect 974 697 1008 731
rect 974 629 1008 663
rect 974 561 1008 595
rect 974 493 1008 527
rect 1130 701 1164 735
rect 1130 622 1164 656
rect 1130 542 1164 576
rect 1130 451 1164 485
rect 1286 701 1320 735
rect 1286 622 1320 656
rect 1286 542 1320 576
rect 1286 451 1320 485
rect 1442 701 1476 735
rect 1442 622 1476 656
rect 1442 542 1476 576
rect 1442 451 1476 485
rect 1598 701 1632 735
rect 1598 622 1632 656
rect 1598 542 1632 576
rect 1598 451 1632 485
rect 1754 701 1788 735
rect 1754 622 1788 656
rect 1754 542 1788 576
rect 1754 451 1788 485
rect 1910 701 1944 735
rect 1910 622 1944 656
rect 1910 542 1944 576
rect 1910 451 1944 485
rect 2066 701 2100 735
rect 2066 622 2100 656
rect 2066 542 2100 576
rect 2066 451 2100 485
rect 2222 701 2256 735
rect 2222 622 2256 656
rect 2222 542 2256 576
rect 2222 451 2256 485
rect 2378 701 2412 735
rect 2378 622 2412 656
rect 2378 542 2412 576
rect 2378 451 2412 485
rect 2534 701 2568 735
rect 2534 622 2568 656
rect 2534 542 2568 576
rect 2534 451 2568 485
rect 2690 701 2724 735
rect 2690 622 2724 656
rect 2690 542 2724 576
rect 2690 451 2724 485
rect 2846 701 2880 735
rect 2846 622 2880 656
rect 2846 542 2880 576
rect 2846 451 2880 485
rect 3002 701 3036 735
rect 3002 622 3036 656
rect 3002 542 3036 576
rect 3002 451 3036 485
rect 3158 701 3192 735
rect 3158 622 3192 656
rect 3158 542 3192 576
rect 3158 451 3192 485
rect 3314 701 3348 735
rect 3314 622 3348 656
rect 3314 542 3348 576
rect 3314 451 3348 485
rect 3470 697 3504 731
rect 3470 622 3504 656
rect 3470 542 3504 576
rect 3470 455 3504 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
<< poly >>
rect 83 743 183 769
rect 239 743 339 769
rect 395 743 495 769
rect 551 743 651 769
rect 707 743 807 769
rect 863 743 963 769
rect 1019 743 1119 769
rect 1175 743 1275 769
rect 1331 743 1431 769
rect 1487 743 1587 769
rect 1643 743 1743 769
rect 1799 743 1899 769
rect 1955 743 2055 769
rect 2111 743 2211 769
rect 2267 743 2367 769
rect 2423 743 2523 769
rect 2579 743 2679 769
rect 2735 743 2835 769
rect 2891 743 2991 769
rect 3047 743 3147 769
rect 3203 743 3303 769
rect 3359 743 3459 769
rect 83 413 183 443
rect 239 413 339 443
rect 395 413 495 443
rect 551 413 651 443
rect 707 413 807 443
rect 863 413 963 443
rect 44 363 963 413
rect 44 329 60 363
rect 94 329 128 363
rect 162 329 196 363
rect 230 329 264 363
rect 298 329 332 363
rect 366 329 400 363
rect 434 329 468 363
rect 502 329 536 363
rect 570 329 604 363
rect 638 329 672 363
rect 706 329 740 363
rect 774 329 808 363
rect 842 329 876 363
rect 910 329 963 363
rect 44 313 963 329
rect 83 291 183 313
rect 239 291 339 313
rect 395 291 495 313
rect 551 291 651 313
rect 707 291 807 313
rect 863 291 963 313
rect 1019 401 1119 443
rect 1175 401 1275 443
rect 1331 401 1431 443
rect 1487 401 1587 443
rect 1643 401 1743 443
rect 1799 401 1899 443
rect 1955 401 2055 443
rect 2111 401 2211 443
rect 2267 401 2367 443
rect 2423 401 2523 443
rect 2579 401 2679 443
rect 2735 401 2835 443
rect 2891 401 2991 443
rect 3047 401 3147 443
rect 3203 401 3303 443
rect 3359 401 3459 443
rect 1019 363 3459 401
rect 1019 329 1248 363
rect 1282 329 1316 363
rect 1350 329 1560 363
rect 1594 329 1628 363
rect 1662 329 1872 363
rect 1906 329 1940 363
rect 1974 329 2184 363
rect 2218 329 2252 363
rect 2286 329 2496 363
rect 2530 329 2564 363
rect 2598 329 2808 363
rect 2842 329 2876 363
rect 2910 329 3120 363
rect 3154 329 3188 363
rect 3222 329 3459 363
rect 1019 313 3459 329
rect 1019 291 1119 313
rect 1175 291 1275 313
rect 1331 291 1431 313
rect 1487 291 1587 313
rect 1643 291 1743 313
rect 1799 291 1899 313
rect 1955 291 2055 313
rect 2111 291 2211 313
rect 2267 291 2367 313
rect 2423 291 2523 313
rect 2579 291 2679 313
rect 2735 291 2835 313
rect 2891 291 2991 313
rect 3047 291 3147 313
rect 3203 291 3303 313
rect 3359 291 3459 313
rect 83 115 183 141
rect 239 115 339 141
rect 395 115 495 141
rect 551 115 651 141
rect 707 115 807 141
rect 863 115 963 141
rect 1019 115 1119 141
rect 1175 115 1275 141
rect 1331 115 1431 141
rect 1487 115 1587 141
rect 1643 115 1743 141
rect 1799 115 1899 141
rect 1955 115 2055 141
rect 2111 115 2211 141
rect 2267 115 2367 141
rect 2423 115 2523 141
rect 2579 115 2679 141
rect 2735 115 2835 141
rect 2891 115 2991 141
rect 3047 115 3147 141
rect 3203 115 3303 141
rect 3359 115 3459 141
<< polycont >>
rect 60 329 94 363
rect 128 329 162 363
rect 196 329 230 363
rect 264 329 298 363
rect 332 329 366 363
rect 400 329 434 363
rect 468 329 502 363
rect 536 329 570 363
rect 604 329 638 363
rect 672 329 706 363
rect 740 329 774 363
rect 808 329 842 363
rect 876 329 910 363
rect 1248 329 1282 363
rect 1316 329 1350 363
rect 1560 329 1594 363
rect 1628 329 1662 363
rect 1872 329 1906 363
rect 1940 329 1974 363
rect 2184 329 2218 363
rect 2252 329 2286 363
rect 2496 329 2530 363
rect 2564 329 2598 363
rect 2808 329 2842 363
rect 2876 329 2910 363
rect 3120 329 3154 363
rect 3188 329 3222 363
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
rect 22 731 136 751
rect 22 729 38 731
rect 72 729 136 731
rect 22 695 30 729
rect 72 697 102 729
rect 64 695 102 697
rect 22 642 136 695
rect 22 608 38 642
rect 72 608 136 642
rect 22 562 136 608
rect 22 528 38 562
rect 72 528 136 562
rect 22 489 136 528
rect 22 455 38 489
rect 72 455 136 489
rect 22 435 136 455
rect 170 735 232 751
rect 480 735 542 751
rect 788 735 858 751
rect 1114 735 1180 751
rect 170 701 194 735
rect 228 701 232 735
rect 170 642 232 701
rect 170 608 194 642
rect 228 608 232 642
rect 170 558 232 608
rect 170 524 194 558
rect 228 524 232 558
rect 170 485 232 524
rect 268 731 446 735
rect 268 729 350 731
rect 384 729 446 731
rect 302 695 340 729
rect 384 697 412 729
rect 374 695 412 697
rect 268 663 446 695
rect 268 629 350 663
rect 384 629 446 663
rect 268 595 446 629
rect 268 561 350 595
rect 384 561 446 595
rect 268 527 446 561
rect 268 493 350 527
rect 384 493 446 527
rect 268 489 446 493
rect 480 701 506 735
rect 540 701 542 735
rect 480 642 542 701
rect 480 608 506 642
rect 540 608 542 642
rect 480 558 542 608
rect 480 524 506 558
rect 540 524 542 558
rect 170 451 194 485
rect 228 453 232 485
rect 480 485 542 524
rect 576 731 754 735
rect 576 729 662 731
rect 696 729 754 731
rect 610 695 648 729
rect 696 697 720 729
rect 682 695 720 697
rect 576 663 754 695
rect 576 629 662 663
rect 696 629 754 663
rect 576 595 754 629
rect 576 561 662 595
rect 696 561 754 595
rect 576 527 754 561
rect 576 493 662 527
rect 696 493 754 527
rect 576 489 754 493
rect 788 701 818 735
rect 852 701 858 735
rect 788 642 858 701
rect 788 608 818 642
rect 852 608 858 642
rect 788 558 858 608
rect 788 524 818 558
rect 852 524 858 558
rect 480 453 506 485
rect 228 451 506 453
rect 540 453 542 485
rect 788 485 858 524
rect 892 731 1070 735
rect 892 729 974 731
rect 1008 729 1070 731
rect 926 695 964 729
rect 1008 697 1036 729
rect 998 695 1036 697
rect 892 663 1070 695
rect 892 629 974 663
rect 1008 629 1070 663
rect 892 595 1070 629
rect 892 561 974 595
rect 1008 561 1070 595
rect 892 527 1070 561
rect 892 493 974 527
rect 1008 493 1070 527
rect 892 489 1070 493
rect 1114 701 1130 735
rect 1164 701 1180 735
rect 1114 656 1180 701
rect 1114 622 1130 656
rect 1164 622 1180 656
rect 1114 576 1180 622
rect 1114 542 1130 576
rect 1164 542 1180 576
rect 1114 498 1180 542
rect 788 453 818 485
rect 540 451 818 453
rect 852 453 858 485
rect 852 451 1070 453
rect 170 397 1070 451
rect 44 329 60 363
rect 94 329 128 363
rect 162 329 196 363
rect 230 329 264 363
rect 298 329 332 363
rect 366 329 400 363
rect 434 329 468 363
rect 502 329 536 363
rect 570 329 604 363
rect 638 329 672 363
rect 706 329 740 363
rect 774 329 808 363
rect 842 329 876 363
rect 910 329 926 363
rect 44 316 926 329
rect 960 350 1070 397
rect 994 316 1032 350
rect 1066 316 1070 350
rect 960 282 1070 316
rect 22 273 129 282
rect 22 239 38 273
rect 72 239 129 273
rect 22 205 129 239
rect 22 171 38 205
rect 72 171 129 205
rect 22 119 129 171
rect 163 269 1070 282
rect 163 235 194 269
rect 228 264 1070 269
rect 228 239 506 264
rect 228 235 234 239
rect 163 201 234 235
rect 480 230 506 239
rect 540 239 818 264
rect 540 230 558 239
rect 163 167 194 201
rect 228 167 234 201
rect 163 151 234 167
rect 268 171 350 205
rect 384 171 446 205
rect 22 85 23 119
rect 57 85 95 119
rect 268 119 446 171
rect 480 196 558 230
rect 805 230 818 239
rect 852 239 1070 264
rect 1114 451 1130 498
rect 1164 451 1180 498
rect 1114 283 1180 451
rect 1214 735 1392 751
rect 1214 729 1286 735
rect 1320 729 1392 735
rect 1248 695 1286 729
rect 1320 695 1358 729
rect 1214 656 1392 695
rect 1214 622 1286 656
rect 1320 622 1392 656
rect 1214 576 1392 622
rect 1214 542 1286 576
rect 1320 542 1392 576
rect 1214 485 1392 542
rect 1214 451 1286 485
rect 1320 451 1392 485
rect 1214 435 1392 451
rect 1426 735 1492 751
rect 1426 701 1442 735
rect 1476 701 1492 735
rect 1426 656 1492 701
rect 1426 622 1442 656
rect 1476 622 1492 656
rect 1426 576 1492 622
rect 1426 542 1442 576
rect 1476 542 1492 576
rect 1426 498 1492 542
rect 1426 451 1442 498
rect 1476 451 1492 498
rect 1232 363 1366 379
rect 1232 350 1248 363
rect 1232 316 1246 350
rect 1282 329 1316 363
rect 1350 350 1366 363
rect 1280 316 1318 329
rect 1352 316 1366 350
rect 1232 313 1366 316
rect 1114 249 1130 283
rect 1164 249 1180 283
rect 1426 283 1492 451
rect 1526 735 1704 751
rect 1526 729 1598 735
rect 1632 729 1704 735
rect 1560 695 1598 729
rect 1632 695 1670 729
rect 1526 656 1704 695
rect 1526 622 1598 656
rect 1632 622 1704 656
rect 1526 576 1704 622
rect 1526 542 1598 576
rect 1632 542 1704 576
rect 1526 485 1704 542
rect 1526 451 1598 485
rect 1632 451 1704 485
rect 1526 435 1704 451
rect 1738 735 1804 751
rect 1738 701 1754 735
rect 1788 701 1804 735
rect 1738 656 1804 701
rect 1738 622 1754 656
rect 1788 622 1804 656
rect 1738 576 1804 622
rect 1738 542 1754 576
rect 1788 542 1804 576
rect 1738 498 1804 542
rect 1738 451 1754 498
rect 1788 451 1804 498
rect 1544 363 1678 379
rect 1544 350 1560 363
rect 1544 316 1558 350
rect 1594 329 1628 363
rect 1662 350 1678 363
rect 1592 316 1630 329
rect 1664 316 1678 350
rect 1544 313 1678 316
rect 852 230 854 239
rect 480 162 506 196
rect 540 162 558 196
rect 480 146 558 162
rect 592 171 662 205
rect 696 171 771 205
rect 302 85 340 119
rect 374 85 412 119
rect 592 119 771 171
rect 805 196 854 230
rect 1114 208 1180 249
rect 805 162 818 196
rect 852 162 854 196
rect 805 146 854 162
rect 888 201 1066 205
rect 888 167 974 201
rect 1008 167 1066 201
rect 626 85 664 119
rect 698 85 736 119
rect 770 85 771 119
rect 888 119 1066 167
rect 1114 174 1130 208
rect 1164 174 1180 208
rect 1114 158 1180 174
rect 1214 269 1392 279
rect 1214 235 1286 269
rect 1320 235 1392 269
rect 1214 201 1392 235
rect 1214 167 1286 201
rect 1320 167 1392 201
rect 922 85 960 119
rect 994 85 1032 119
rect 1214 119 1392 167
rect 1426 249 1442 283
rect 1476 249 1492 283
rect 1738 283 1804 451
rect 1838 735 2016 751
rect 1838 729 1910 735
rect 1944 729 2016 735
rect 1872 695 1910 729
rect 1944 695 1982 729
rect 1838 656 2016 695
rect 1838 622 1910 656
rect 1944 622 2016 656
rect 1838 576 2016 622
rect 1838 542 1910 576
rect 1944 542 2016 576
rect 1838 485 2016 542
rect 1838 451 1910 485
rect 1944 451 2016 485
rect 1838 435 2016 451
rect 2050 735 2116 751
rect 2050 701 2066 735
rect 2100 701 2116 735
rect 2050 656 2116 701
rect 2050 622 2066 656
rect 2100 622 2116 656
rect 2050 576 2116 622
rect 2050 542 2066 576
rect 2100 542 2116 576
rect 2050 498 2116 542
rect 2050 451 2066 498
rect 2100 451 2116 498
rect 1856 363 1990 379
rect 1856 350 1872 363
rect 1856 316 1870 350
rect 1906 329 1940 363
rect 1974 350 1990 363
rect 1904 316 1942 329
rect 1976 316 1990 350
rect 1856 313 1990 316
rect 1426 208 1492 249
rect 1426 174 1442 208
rect 1476 174 1492 208
rect 1426 158 1492 174
rect 1526 269 1704 279
rect 1526 235 1598 269
rect 1632 235 1704 269
rect 1526 201 1704 235
rect 1526 167 1598 201
rect 1632 167 1704 201
rect 1248 85 1286 119
rect 1320 85 1358 119
rect 1526 119 1704 167
rect 1738 249 1754 283
rect 1788 249 1804 283
rect 2050 283 2116 451
rect 2150 735 2328 751
rect 2150 729 2222 735
rect 2256 729 2328 735
rect 2184 695 2222 729
rect 2256 695 2294 729
rect 2150 656 2328 695
rect 2150 622 2222 656
rect 2256 622 2328 656
rect 2150 576 2328 622
rect 2150 542 2222 576
rect 2256 542 2328 576
rect 2150 485 2328 542
rect 2150 451 2222 485
rect 2256 451 2328 485
rect 2150 435 2328 451
rect 2362 735 2428 751
rect 2362 701 2378 735
rect 2412 701 2428 735
rect 2362 656 2428 701
rect 2362 622 2378 656
rect 2412 622 2428 656
rect 2362 576 2428 622
rect 2362 542 2378 576
rect 2412 542 2428 576
rect 2362 498 2428 542
rect 2362 451 2378 498
rect 2412 451 2428 498
rect 2168 363 2302 379
rect 2168 350 2184 363
rect 2168 316 2182 350
rect 2218 329 2252 363
rect 2286 350 2302 363
rect 2216 316 2254 329
rect 2288 316 2302 350
rect 2168 313 2302 316
rect 1738 208 1804 249
rect 1738 174 1754 208
rect 1788 174 1804 208
rect 1738 158 1804 174
rect 1838 269 2016 279
rect 1838 235 1910 269
rect 1944 235 2016 269
rect 1838 201 2016 235
rect 1838 167 1910 201
rect 1944 167 2016 201
rect 1560 85 1598 119
rect 1632 85 1670 119
rect 1838 119 2016 167
rect 2050 249 2066 283
rect 2100 249 2116 283
rect 2362 283 2428 451
rect 2462 735 2640 751
rect 2462 729 2534 735
rect 2568 729 2640 735
rect 2496 695 2534 729
rect 2568 695 2606 729
rect 2462 656 2640 695
rect 2462 622 2534 656
rect 2568 622 2640 656
rect 2462 576 2640 622
rect 2462 542 2534 576
rect 2568 542 2640 576
rect 2462 485 2640 542
rect 2462 451 2534 485
rect 2568 451 2640 485
rect 2462 435 2640 451
rect 2674 735 2740 751
rect 2674 701 2690 735
rect 2724 701 2740 735
rect 2674 656 2740 701
rect 2674 622 2690 656
rect 2724 622 2740 656
rect 2674 576 2740 622
rect 2674 542 2690 576
rect 2724 542 2740 576
rect 2674 498 2740 542
rect 2674 451 2690 498
rect 2724 451 2740 498
rect 2480 363 2614 379
rect 2480 350 2496 363
rect 2480 316 2494 350
rect 2530 329 2564 363
rect 2598 350 2614 363
rect 2528 316 2566 329
rect 2600 316 2614 350
rect 2480 313 2614 316
rect 2050 208 2116 249
rect 2050 174 2066 208
rect 2100 174 2116 208
rect 2050 158 2116 174
rect 2150 269 2328 279
rect 2150 235 2222 269
rect 2256 235 2328 269
rect 2150 201 2328 235
rect 2150 167 2222 201
rect 2256 167 2328 201
rect 1872 85 1910 119
rect 1944 85 1982 119
rect 2150 119 2328 167
rect 2362 249 2378 283
rect 2412 249 2428 283
rect 2674 283 2740 451
rect 2774 735 2952 751
rect 2774 729 2846 735
rect 2880 729 2952 735
rect 2808 695 2846 729
rect 2880 695 2918 729
rect 2774 656 2952 695
rect 2774 622 2846 656
rect 2880 622 2952 656
rect 2774 576 2952 622
rect 2774 542 2846 576
rect 2880 542 2952 576
rect 2774 485 2952 542
rect 2774 451 2846 485
rect 2880 451 2952 485
rect 2774 435 2952 451
rect 2986 735 3052 751
rect 2986 701 3002 735
rect 3036 701 3052 735
rect 2986 656 3052 701
rect 2986 622 3002 656
rect 3036 622 3052 656
rect 2986 576 3052 622
rect 2986 542 3002 576
rect 3036 542 3052 576
rect 2986 498 3052 542
rect 2986 451 3002 498
rect 3036 451 3052 498
rect 2792 363 2926 379
rect 2792 350 2808 363
rect 2792 316 2806 350
rect 2842 329 2876 363
rect 2910 350 2926 363
rect 2840 316 2878 329
rect 2912 316 2926 350
rect 2792 313 2926 316
rect 2362 208 2428 249
rect 2362 174 2378 208
rect 2412 174 2428 208
rect 2362 158 2428 174
rect 2462 269 2640 279
rect 2462 235 2534 269
rect 2568 235 2640 269
rect 2462 201 2640 235
rect 2462 167 2534 201
rect 2568 167 2640 201
rect 2184 85 2222 119
rect 2256 85 2294 119
rect 2462 119 2640 167
rect 2674 249 2690 283
rect 2724 249 2740 283
rect 2986 283 3052 451
rect 3086 735 3264 751
rect 3086 729 3158 735
rect 3192 729 3264 735
rect 3120 695 3158 729
rect 3192 695 3230 729
rect 3086 656 3264 695
rect 3086 622 3158 656
rect 3192 622 3264 656
rect 3086 576 3264 622
rect 3086 542 3158 576
rect 3192 542 3264 576
rect 3086 485 3264 542
rect 3086 451 3158 485
rect 3192 451 3264 485
rect 3086 435 3264 451
rect 3298 735 3380 751
rect 3298 701 3314 735
rect 3348 701 3380 735
rect 3298 656 3380 701
rect 3298 622 3314 656
rect 3348 622 3380 656
rect 3298 576 3380 622
rect 3298 542 3314 576
rect 3348 542 3380 576
rect 3298 498 3380 542
rect 3298 451 3314 498
rect 3348 451 3380 498
rect 3104 363 3238 379
rect 3104 350 3120 363
rect 3104 316 3118 350
rect 3154 329 3188 363
rect 3222 350 3238 363
rect 3152 316 3190 329
rect 3224 316 3238 350
rect 3104 313 3238 316
rect 2674 208 2740 249
rect 2674 174 2690 208
rect 2724 174 2740 208
rect 2674 158 2740 174
rect 2774 269 2952 279
rect 2774 235 2846 269
rect 2880 235 2952 269
rect 2774 201 2952 235
rect 2774 167 2846 201
rect 2880 167 2952 201
rect 2496 85 2534 119
rect 2568 85 2606 119
rect 2774 119 2952 167
rect 2986 249 3002 283
rect 3036 249 3052 283
rect 3298 283 3380 451
rect 3414 731 3520 751
rect 3414 729 3470 731
rect 3504 729 3520 731
rect 3448 697 3470 729
rect 3448 695 3486 697
rect 3414 656 3520 695
rect 3414 622 3470 656
rect 3504 622 3520 656
rect 3414 576 3520 622
rect 3414 542 3470 576
rect 3504 542 3520 576
rect 3414 489 3520 542
rect 3414 455 3470 489
rect 3504 455 3520 489
rect 3414 435 3520 455
rect 2986 208 3052 249
rect 2986 174 3002 208
rect 3036 174 3052 208
rect 2986 158 3052 174
rect 3086 269 3264 279
rect 3086 235 3158 269
rect 3192 235 3264 269
rect 3086 201 3264 235
rect 3086 167 3158 201
rect 3192 167 3264 201
rect 2808 85 2846 119
rect 2880 85 2918 119
rect 3086 119 3264 167
rect 3298 249 3314 283
rect 3348 249 3380 283
rect 3298 208 3380 249
rect 3298 174 3314 208
rect 3348 174 3380 208
rect 3298 158 3380 174
rect 3414 279 3520 299
rect 3414 245 3470 279
rect 3504 245 3520 279
rect 3414 208 3520 245
rect 3414 174 3470 208
rect 3504 174 3520 208
rect 3120 85 3158 119
rect 3192 85 3230 119
rect 3414 119 3520 174
rect 3448 85 3486 119
rect 268 83 446 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 30 697 38 729
rect 38 697 64 729
rect 30 695 64 697
rect 102 695 136 729
rect 268 695 302 729
rect 340 697 350 729
rect 350 697 374 729
rect 340 695 374 697
rect 412 695 446 729
rect 576 695 610 729
rect 648 697 662 729
rect 662 697 682 729
rect 648 695 682 697
rect 720 695 754 729
rect 892 695 926 729
rect 964 697 974 729
rect 974 697 998 729
rect 964 695 998 697
rect 1036 695 1070 729
rect 960 316 994 350
rect 1032 316 1066 350
rect 23 85 57 119
rect 95 85 129 119
rect 1130 485 1164 498
rect 1130 464 1164 485
rect 1214 695 1248 729
rect 1286 701 1320 729
rect 1286 695 1320 701
rect 1358 695 1392 729
rect 1442 485 1476 498
rect 1442 464 1476 485
rect 1246 329 1248 350
rect 1248 329 1280 350
rect 1318 329 1350 350
rect 1350 329 1352 350
rect 1246 316 1280 329
rect 1318 316 1352 329
rect 1526 695 1560 729
rect 1598 701 1632 729
rect 1598 695 1632 701
rect 1670 695 1704 729
rect 1754 485 1788 498
rect 1754 464 1788 485
rect 1558 329 1560 350
rect 1560 329 1592 350
rect 1630 329 1662 350
rect 1662 329 1664 350
rect 1558 316 1592 329
rect 1630 316 1664 329
rect 268 85 302 119
rect 340 85 374 119
rect 412 85 446 119
rect 592 85 626 119
rect 664 85 698 119
rect 736 85 770 119
rect 888 85 922 119
rect 960 85 994 119
rect 1032 85 1066 119
rect 1838 695 1872 729
rect 1910 701 1944 729
rect 1910 695 1944 701
rect 1982 695 2016 729
rect 2066 485 2100 498
rect 2066 464 2100 485
rect 1870 329 1872 350
rect 1872 329 1904 350
rect 1942 329 1974 350
rect 1974 329 1976 350
rect 1870 316 1904 329
rect 1942 316 1976 329
rect 1214 85 1248 119
rect 1286 85 1320 119
rect 1358 85 1392 119
rect 2150 695 2184 729
rect 2222 701 2256 729
rect 2222 695 2256 701
rect 2294 695 2328 729
rect 2378 485 2412 498
rect 2378 464 2412 485
rect 2182 329 2184 350
rect 2184 329 2216 350
rect 2254 329 2286 350
rect 2286 329 2288 350
rect 2182 316 2216 329
rect 2254 316 2288 329
rect 1526 85 1560 119
rect 1598 85 1632 119
rect 1670 85 1704 119
rect 2462 695 2496 729
rect 2534 701 2568 729
rect 2534 695 2568 701
rect 2606 695 2640 729
rect 2690 485 2724 498
rect 2690 464 2724 485
rect 2494 329 2496 350
rect 2496 329 2528 350
rect 2566 329 2598 350
rect 2598 329 2600 350
rect 2494 316 2528 329
rect 2566 316 2600 329
rect 1838 85 1872 119
rect 1910 85 1944 119
rect 1982 85 2016 119
rect 2774 695 2808 729
rect 2846 701 2880 729
rect 2846 695 2880 701
rect 2918 695 2952 729
rect 3002 485 3036 498
rect 3002 464 3036 485
rect 2806 329 2808 350
rect 2808 329 2840 350
rect 2878 329 2910 350
rect 2910 329 2912 350
rect 2806 316 2840 329
rect 2878 316 2912 329
rect 2150 85 2184 119
rect 2222 85 2256 119
rect 2294 85 2328 119
rect 3086 695 3120 729
rect 3158 701 3192 729
rect 3158 695 3192 701
rect 3230 695 3264 729
rect 3314 485 3348 498
rect 3314 464 3348 485
rect 3118 329 3120 350
rect 3120 329 3152 350
rect 3190 329 3222 350
rect 3222 329 3224 350
rect 3118 316 3152 329
rect 3190 316 3224 329
rect 2462 85 2496 119
rect 2534 85 2568 119
rect 2606 85 2640 119
rect 3414 695 3448 729
rect 3486 697 3504 729
rect 3504 697 3520 729
rect 3486 695 3520 697
rect 2774 85 2808 119
rect 2846 85 2880 119
rect 2918 85 2952 119
rect 3086 85 3120 119
rect 3158 85 3192 119
rect 3230 85 3264 119
rect 3414 85 3448 119
rect 3486 85 3520 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 831 3552 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
rect 0 791 3552 797
rect 0 729 3552 763
rect 0 695 30 729
rect 64 695 102 729
rect 136 695 268 729
rect 302 695 340 729
rect 374 695 412 729
rect 446 695 576 729
rect 610 695 648 729
rect 682 695 720 729
rect 754 695 892 729
rect 926 695 964 729
rect 998 695 1036 729
rect 1070 695 1214 729
rect 1248 695 1286 729
rect 1320 695 1358 729
rect 1392 695 1526 729
rect 1560 695 1598 729
rect 1632 695 1670 729
rect 1704 695 1838 729
rect 1872 695 1910 729
rect 1944 695 1982 729
rect 2016 695 2150 729
rect 2184 695 2222 729
rect 2256 695 2294 729
rect 2328 695 2462 729
rect 2496 695 2534 729
rect 2568 695 2606 729
rect 2640 695 2774 729
rect 2808 695 2846 729
rect 2880 695 2918 729
rect 2952 695 3086 729
rect 3120 695 3158 729
rect 3192 695 3230 729
rect 3264 695 3414 729
rect 3448 695 3486 729
rect 3520 695 3552 729
rect 0 689 3552 695
rect 1118 498 1176 504
rect 1430 498 1488 504
rect 1742 498 1800 504
rect 2054 498 2112 504
rect 2366 498 2424 504
rect 2678 498 2736 504
rect 2990 498 3048 504
rect 3302 498 3360 504
rect 1118 464 1130 498
rect 1164 464 1442 498
rect 1476 464 1754 498
rect 1788 464 2066 498
rect 2100 464 2378 498
rect 2412 464 2690 498
rect 2724 464 3002 498
rect 3036 464 3314 498
rect 3348 464 3360 498
rect 1118 458 1176 464
rect 1430 458 1488 464
rect 1742 458 1800 464
rect 2054 458 2112 464
rect 2366 458 2424 464
rect 2678 458 2736 464
rect 2990 458 3048 464
rect 3302 458 3360 464
rect 948 350 1072 356
rect 1234 350 1364 356
rect 1546 350 1676 356
rect 1858 350 1988 356
rect 2170 350 2300 356
rect 2482 350 2612 356
rect 2794 350 2924 356
rect 3106 350 3236 356
rect 948 316 960 350
rect 994 316 1032 350
rect 1066 316 1246 350
rect 1280 316 1318 350
rect 1352 316 1558 350
rect 1592 316 1630 350
rect 1664 316 1870 350
rect 1904 316 1942 350
rect 1976 316 2182 350
rect 2216 316 2254 350
rect 2288 316 2494 350
rect 2528 316 2566 350
rect 2600 316 2806 350
rect 2840 316 2878 350
rect 2912 316 3118 350
rect 3152 316 3190 350
rect 3224 316 3250 350
rect 948 310 1072 316
rect 1234 310 1364 316
rect 1546 310 1676 316
rect 1858 310 1988 316
rect 2170 310 2300 316
rect 2482 310 2612 316
rect 2794 310 2924 316
rect 3106 310 3236 316
rect 0 119 3552 125
rect 0 85 23 119
rect 57 85 95 119
rect 129 85 268 119
rect 302 85 340 119
rect 374 85 412 119
rect 446 85 592 119
rect 626 85 664 119
rect 698 85 736 119
rect 770 85 888 119
rect 922 85 960 119
rect 994 85 1032 119
rect 1066 85 1214 119
rect 1248 85 1286 119
rect 1320 85 1358 119
rect 1392 85 1526 119
rect 1560 85 1598 119
rect 1632 85 1670 119
rect 1704 85 1838 119
rect 1872 85 1910 119
rect 1944 85 1982 119
rect 2016 85 2150 119
rect 2184 85 2222 119
rect 2256 85 2294 119
rect 2328 85 2462 119
rect 2496 85 2534 119
rect 2568 85 2606 119
rect 2640 85 2774 119
rect 2808 85 2846 119
rect 2880 85 2918 119
rect 2952 85 3086 119
rect 3120 85 3158 119
rect 3192 85 3230 119
rect 3264 85 3414 119
rect 3448 85 3486 119
rect 3520 85 3552 119
rect 0 51 3552 85
rect 0 17 3552 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -23 3552 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_16
flabel metal1 s 0 51 3552 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 3552 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 1118 464 3360 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel metal1 s 1872 11 1872 11 0 FreeSans 340 0 0 0 VNB
flabel metal1 s 0 689 3552 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 3552 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 1872 802 1872 802 0 FreeSans 340 0 0 0 VPB
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 3552 814
string GDS_END 1130684
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1091408
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
