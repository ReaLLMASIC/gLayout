magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 6 21 827 203
rect 28 -17 62 21
<< locali >>
rect 17 151 74 265
rect 176 324 246 475
rect 280 357 344 475
rect 176 199 210 324
rect 280 290 322 357
rect 496 325 546 493
rect 664 325 714 493
rect 256 199 322 290
rect 368 289 455 323
rect 496 291 811 325
rect 368 199 402 289
rect 762 181 811 291
rect 504 145 811 181
rect 504 51 554 145
rect 656 51 722 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 23 333 90 490
rect 23 299 142 333
rect 108 165 142 299
rect 401 359 451 527
rect 580 359 630 527
rect 748 359 798 527
rect 436 215 728 249
rect 436 165 470 215
rect 108 131 470 165
rect 24 17 74 117
rect 140 61 174 131
rect 214 17 280 97
rect 314 61 348 131
rect 392 17 468 97
rect 588 17 622 111
rect 756 17 790 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 368 199 402 289 6 A
port 1 nsew signal input
rlabel locali s 368 289 455 323 6 A
port 1 nsew signal input
rlabel locali s 256 199 322 290 6 B
port 2 nsew signal input
rlabel locali s 280 290 322 357 6 B
port 2 nsew signal input
rlabel locali s 280 357 344 475 6 B
port 2 nsew signal input
rlabel locali s 176 199 210 324 6 C
port 3 nsew signal input
rlabel locali s 176 324 246 475 6 C
port 3 nsew signal input
rlabel locali s 17 151 74 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 28 -17 62 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 6 21 827 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 656 51 722 145 6 X
port 9 nsew signal output
rlabel locali s 504 51 554 145 6 X
port 9 nsew signal output
rlabel locali s 504 145 811 181 6 X
port 9 nsew signal output
rlabel locali s 762 181 811 291 6 X
port 9 nsew signal output
rlabel locali s 496 291 811 325 6 X
port 9 nsew signal output
rlabel locali s 664 325 714 493 6 X
port 9 nsew signal output
rlabel locali s 496 325 546 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1068202
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1060956
<< end >>
