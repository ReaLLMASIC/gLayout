magic
tech sky130B
magscale 1 2
timestamp 1701704242
<< metal1 >>
rect 0 2668 38722 2696
tri 38636 2640 38664 2668 ne
rect 38664 2640 38722 2668
rect 0 2588 2249 2640
rect 2301 2588 2313 2640
rect 2365 2588 2533 2640
rect 2585 2588 2597 2640
rect 2649 2588 7081 2640
rect 7133 2588 7145 2640
rect 7197 2588 7365 2640
rect 7417 2588 7429 2640
rect 7481 2588 11913 2640
rect 11965 2588 11977 2640
rect 12029 2588 12197 2640
rect 12249 2588 12261 2640
rect 12313 2588 16745 2640
rect 16797 2588 16809 2640
rect 16861 2588 17029 2640
rect 17081 2588 17093 2640
rect 17145 2588 21577 2640
rect 21629 2588 21641 2640
rect 21693 2588 21861 2640
rect 21913 2588 21925 2640
rect 21977 2588 26409 2640
rect 26461 2588 26473 2640
rect 26525 2588 26693 2640
rect 26745 2588 26757 2640
rect 26809 2588 31241 2640
rect 31293 2588 31305 2640
rect 31357 2588 31525 2640
rect 31577 2588 31589 2640
rect 31641 2588 36073 2640
rect 36125 2588 36137 2640
rect 36189 2588 36357 2640
rect 36409 2588 36421 2640
rect 36473 2588 38612 2640
tri 38664 2634 38670 2640 ne
tri 38664 2588 38670 2594 se
rect 38670 2588 38722 2640
tri 38636 2560 38664 2588 se
rect 38664 2560 38722 2588
rect 0 2532 38722 2560
rect 470 2358 793 2486
rect 859 2452 865 2504
rect 917 2452 933 2504
rect 985 2452 1001 2504
rect 1053 2452 1059 2504
rect 859 2392 1059 2452
rect 859 2340 865 2392
rect 917 2340 933 2392
rect 985 2340 1001 2392
rect 1053 2340 1059 2392
rect 5691 2452 5697 2504
rect 5749 2452 5765 2504
rect 5817 2452 5833 2504
rect 5885 2452 5891 2504
rect 5691 2392 5891 2452
rect 5691 2340 5697 2392
rect 5749 2340 5765 2392
rect 5817 2340 5833 2392
rect 5885 2340 5891 2392
rect 8415 2452 8421 2504
rect 8473 2452 8489 2504
rect 8541 2452 8557 2504
rect 8609 2452 8615 2504
rect 8415 2392 8615 2452
rect 8415 2340 8421 2392
rect 8473 2340 8489 2392
rect 8541 2340 8557 2392
rect 8609 2340 8615 2392
rect 10523 2452 10529 2504
rect 10581 2452 10597 2504
rect 10649 2452 10665 2504
rect 10717 2452 10723 2504
rect 10523 2392 10723 2452
rect 10523 2340 10529 2392
rect 10581 2340 10597 2392
rect 10649 2340 10665 2392
rect 10717 2340 10723 2392
rect 13247 2452 13253 2504
rect 13305 2452 13321 2504
rect 13373 2452 13389 2504
rect 13441 2452 13447 2504
rect 13247 2392 13447 2452
rect 13247 2340 13253 2392
rect 13305 2340 13321 2392
rect 13373 2340 13389 2392
rect 13441 2340 13447 2392
rect 15355 2452 15361 2504
rect 15413 2452 15429 2504
rect 15481 2452 15497 2504
rect 15549 2452 15555 2504
rect 15355 2392 15555 2452
rect 15355 2340 15361 2392
rect 15413 2340 15429 2392
rect 15481 2340 15497 2392
rect 15549 2340 15555 2392
rect 18079 2452 18085 2504
rect 18137 2452 18153 2504
rect 18205 2452 18221 2504
rect 18273 2452 18279 2504
rect 18079 2392 18279 2452
rect 18079 2340 18085 2392
rect 18137 2340 18153 2392
rect 18205 2340 18221 2392
rect 18273 2340 18279 2392
rect 20187 2452 20193 2504
rect 20245 2452 20261 2504
rect 20313 2452 20329 2504
rect 20381 2452 20387 2504
rect 20187 2392 20387 2452
rect 20187 2340 20193 2392
rect 20245 2340 20261 2392
rect 20313 2340 20329 2392
rect 20381 2340 20387 2392
rect 22911 2452 22917 2504
rect 22969 2452 22985 2504
rect 23037 2452 23053 2504
rect 23105 2452 23111 2504
rect 22911 2392 23111 2452
rect 22911 2340 22917 2392
rect 22969 2340 22985 2392
rect 23037 2340 23053 2392
rect 23105 2340 23111 2392
rect 25019 2452 25025 2504
rect 25077 2452 25093 2504
rect 25145 2452 25161 2504
rect 25213 2452 25219 2504
rect 25019 2392 25219 2452
rect 25019 2340 25025 2392
rect 25077 2340 25093 2392
rect 25145 2340 25161 2392
rect 25213 2340 25219 2392
rect 27743 2452 27749 2504
rect 27801 2452 27817 2504
rect 27869 2452 27885 2504
rect 27937 2452 27943 2504
rect 27743 2392 27943 2452
rect 27743 2340 27749 2392
rect 27801 2340 27817 2392
rect 27869 2340 27885 2392
rect 27937 2340 27943 2392
rect 29851 2452 29857 2504
rect 29909 2452 29925 2504
rect 29977 2452 29993 2504
rect 30045 2452 30051 2504
rect 29851 2392 30051 2452
rect 29851 2340 29857 2392
rect 29909 2340 29925 2392
rect 29977 2340 29993 2392
rect 30045 2340 30051 2392
rect 32575 2452 32581 2504
rect 32633 2452 32649 2504
rect 32701 2452 32717 2504
rect 32769 2452 32775 2504
rect 32575 2392 32775 2452
rect 32575 2340 32581 2392
rect 32633 2340 32649 2392
rect 32701 2340 32717 2392
rect 32769 2340 32775 2392
rect 34683 2452 34689 2504
rect 34741 2452 34757 2504
rect 34809 2452 34825 2504
rect 34877 2452 34883 2504
rect 34683 2392 34883 2452
rect 34683 2340 34689 2392
rect 34741 2340 34757 2392
rect 34809 2340 34825 2392
rect 34877 2340 34883 2392
rect 37407 2452 37413 2504
rect 37465 2452 37481 2504
rect 37533 2452 37549 2504
rect 37601 2452 37607 2504
rect 37407 2392 37607 2452
rect 37407 2340 37413 2392
rect 37465 2340 37481 2392
rect 37533 2340 37549 2392
rect 37601 2340 37607 2392
rect 2119 2239 2231 2273
rect 2642 2241 2773 2273
rect 6952 2238 7061 2273
rect 7473 2242 7610 2276
rect 11768 2236 11926 2274
rect 12306 2235 12442 2272
rect 16592 2238 16733 2272
rect 17127 2237 17273 2272
rect 21435 2236 21590 2271
rect 21969 2237 22116 2274
rect 26253 2236 26380 2273
rect 26773 2237 26903 2271
rect 31104 2241 31268 2274
rect 31608 2233 31749 2273
rect 35958 2241 36085 2277
rect 36431 2238 36579 2272
rect 144 2159 196 2165
rect 144 2093 196 2107
rect 144 2035 196 2041
rect 300 2159 352 2165
rect 300 2093 352 2107
rect 300 2035 352 2041
rect 453 2159 505 2165
rect 453 2093 505 2107
rect 453 2035 505 2041
rect 608 2160 660 2171
rect 608 2096 660 2108
rect 608 2038 660 2044
rect 765 2159 817 2165
rect 765 2095 817 2107
rect 765 2033 817 2043
rect 4078 2155 4130 2163
rect 4078 2091 4130 2103
rect 4078 2033 4130 2039
rect 4235 2160 4287 2171
rect 4235 2096 4287 2108
rect 4235 2038 4287 2044
rect 4392 2159 4444 2165
rect 4392 2093 4444 2107
rect 4392 2035 4444 2041
rect 4548 2159 4600 2165
rect 4548 2093 4600 2107
rect 4548 2035 4600 2041
rect 4704 2159 4756 2165
rect 4704 2095 4756 2107
rect 4704 2035 4756 2043
rect 4974 2159 5026 2165
rect 4974 2093 5026 2107
rect 4974 2035 5026 2041
rect 5130 2159 5182 2165
rect 5130 2093 5182 2107
rect 5130 2035 5182 2041
rect 5287 2159 5339 2165
rect 5287 2093 5339 2107
rect 5287 2035 5339 2041
rect 5440 2160 5492 2171
rect 9067 2165 9119 2171
rect 5440 2096 5492 2108
rect 5440 2038 5492 2044
rect 5600 2157 5652 2163
rect 5600 2091 5652 2105
rect 5600 2033 5652 2039
rect 8910 2157 8962 2163
rect 8910 2091 8962 2105
rect 8910 2033 8962 2039
rect 9067 2096 9119 2113
rect 9067 2038 9119 2044
rect 9223 2159 9275 2165
rect 9223 2093 9275 2107
rect 9223 2035 9275 2041
rect 9380 2159 9432 2165
rect 9380 2093 9432 2107
rect 9380 2035 9432 2041
rect 9536 2159 9588 2165
rect 9536 2093 9588 2107
rect 9536 2035 9588 2041
rect 9806 2159 9858 2165
rect 9806 2093 9858 2107
rect 9806 2035 9858 2041
rect 9962 2159 10014 2165
rect 9962 2093 10014 2107
rect 9962 2035 10014 2041
rect 10119 2159 10171 2165
rect 10119 2093 10171 2107
rect 10119 2035 10171 2041
rect 10272 2160 10324 2171
rect 13899 2165 13951 2171
rect 10272 2096 10324 2108
rect 10272 2038 10324 2044
rect 10432 2157 10484 2163
rect 10432 2091 10484 2105
rect 10432 2033 10484 2039
rect 13742 2157 13794 2163
rect 13742 2091 13794 2105
rect 13742 2033 13794 2039
rect 13899 2096 13951 2113
rect 13899 2038 13951 2044
rect 14055 2159 14107 2165
rect 14055 2093 14107 2107
rect 14055 2035 14107 2041
rect 14212 2159 14264 2165
rect 14212 2093 14264 2107
rect 14212 2035 14264 2041
rect 14368 2159 14420 2165
rect 14368 2093 14420 2107
rect 14368 2035 14420 2041
rect 14638 2159 14690 2165
rect 14638 2093 14690 2107
rect 14638 2035 14690 2041
rect 14794 2159 14846 2165
rect 14794 2093 14846 2107
rect 14794 2035 14846 2041
rect 14951 2159 15003 2165
rect 14951 2093 15003 2107
rect 14951 2035 15003 2041
rect 15104 2160 15156 2171
rect 18731 2165 18783 2171
rect 19939 2165 19991 2171
rect 15104 2096 15156 2108
rect 15104 2038 15156 2044
rect 15264 2157 15316 2163
rect 15264 2091 15316 2105
rect 15264 2033 15316 2039
rect 18574 2157 18626 2163
rect 18574 2091 18626 2105
rect 18574 2033 18626 2039
rect 18731 2096 18783 2113
rect 18731 2038 18783 2044
rect 18887 2159 18939 2165
rect 18887 2093 18939 2107
rect 18887 2035 18939 2041
rect 19044 2159 19096 2165
rect 19044 2093 19096 2107
rect 19044 2035 19096 2041
rect 19200 2159 19252 2165
rect 19200 2093 19252 2107
rect 19200 2035 19252 2041
rect 19470 2159 19522 2165
rect 19470 2093 19522 2107
rect 19470 2035 19522 2041
rect 19626 2159 19678 2165
rect 19626 2093 19678 2107
rect 19626 2035 19678 2041
rect 19783 2159 19835 2165
rect 19783 2093 19835 2107
rect 19783 2035 19835 2041
rect 19939 2096 19991 2113
rect 19939 2038 19991 2044
rect 20093 2159 20145 2165
rect 20093 2095 20145 2107
rect 20093 2033 20145 2043
rect 23409 2159 23461 2165
rect 23409 2095 23461 2107
rect 23409 2033 23461 2043
rect 23560 2160 23612 2171
rect 24774 2165 24826 2171
rect 28395 2165 28447 2171
rect 29606 2165 29658 2171
rect 33227 2165 33279 2171
rect 34435 2165 34487 2171
rect 23560 2096 23612 2108
rect 23560 2038 23612 2044
rect 23719 2159 23771 2165
rect 23719 2093 23771 2107
rect 23719 2035 23771 2041
rect 23876 2159 23928 2165
rect 23876 2093 23928 2107
rect 23876 2035 23928 2041
rect 24032 2159 24084 2165
rect 24032 2093 24084 2107
rect 24032 2035 24084 2041
rect 24302 2159 24354 2165
rect 24302 2093 24354 2107
rect 24302 2035 24354 2041
rect 24458 2159 24510 2165
rect 24458 2093 24510 2107
rect 24458 2035 24510 2041
rect 24615 2159 24667 2165
rect 24615 2093 24667 2107
rect 24615 2035 24667 2041
rect 24774 2096 24826 2113
rect 24774 2038 24826 2044
rect 24925 2159 24977 2165
rect 24925 2095 24977 2107
rect 24925 2033 24977 2043
rect 28241 2159 28293 2165
rect 28241 2091 28293 2107
rect 28241 2033 28293 2039
rect 28395 2096 28447 2113
rect 28395 2038 28447 2044
rect 28551 2159 28603 2165
rect 28551 2093 28603 2107
rect 28551 2035 28603 2041
rect 28708 2159 28760 2165
rect 28708 2093 28760 2107
rect 28708 2035 28760 2041
rect 28864 2159 28916 2165
rect 28864 2093 28916 2107
rect 28864 2035 28916 2041
rect 29134 2159 29186 2165
rect 29134 2093 29186 2107
rect 29134 2035 29186 2041
rect 29290 2159 29342 2165
rect 29290 2093 29342 2107
rect 29290 2035 29342 2041
rect 29447 2159 29499 2165
rect 29447 2093 29499 2107
rect 29447 2035 29499 2041
rect 29606 2096 29658 2113
rect 29606 2038 29658 2044
rect 29757 2159 29809 2165
rect 29757 2091 29809 2107
rect 29757 2033 29809 2039
rect 33073 2159 33125 2165
rect 33073 2091 33125 2107
rect 33073 2033 33125 2039
rect 33227 2096 33279 2113
rect 33227 2038 33279 2044
rect 33383 2159 33435 2165
rect 33383 2093 33435 2107
rect 33383 2035 33435 2041
rect 33540 2159 33592 2165
rect 33540 2093 33592 2107
rect 33540 2035 33592 2041
rect 33696 2159 33748 2165
rect 33696 2093 33748 2107
rect 33696 2035 33748 2041
rect 33966 2159 34018 2165
rect 33966 2093 34018 2107
rect 33966 2035 34018 2041
rect 34122 2159 34174 2165
rect 34122 2093 34174 2107
rect 34122 2035 34174 2041
rect 34279 2159 34331 2165
rect 34279 2093 34331 2107
rect 34279 2035 34331 2041
rect 34435 2096 34487 2113
rect 34435 2038 34487 2044
rect 34589 2159 34641 2165
rect 34589 2091 34641 2107
rect 34589 2033 34641 2039
rect 37905 2160 37957 2166
rect 37905 2091 37957 2108
rect 37905 2033 37957 2039
rect 38059 2165 38111 2171
rect 38059 2096 38111 2113
rect 38059 2038 38111 2044
rect 38215 2160 38267 2166
rect 38215 2093 38267 2108
rect 38215 2035 38267 2041
rect 38372 2160 38424 2166
rect 38372 2093 38424 2108
rect 38372 2035 38424 2041
rect 38528 2160 38580 2166
rect 38528 2093 38580 2108
rect 38528 2035 38580 2041
rect 444 1686 676 1776
rect 1115 1762 1121 1814
rect 1173 1762 1189 1814
rect 1241 1762 1257 1814
rect 1309 1762 1315 1814
rect 1115 1718 1315 1762
rect 1115 1666 1121 1718
rect 1173 1666 1189 1718
rect 1241 1666 1257 1718
rect 1309 1666 1315 1718
rect 5947 1762 5953 1814
rect 6005 1762 6021 1814
rect 6073 1762 6089 1814
rect 6141 1762 6147 1814
rect 5947 1718 6147 1762
rect 5947 1666 5953 1718
rect 6005 1666 6021 1718
rect 6073 1666 6089 1718
rect 6141 1666 6147 1718
rect 8671 1762 8677 1814
rect 8729 1762 8745 1814
rect 8797 1762 8813 1814
rect 8865 1762 8871 1814
rect 8671 1718 8871 1762
rect 8671 1666 8677 1718
rect 8729 1666 8745 1718
rect 8797 1666 8813 1718
rect 8865 1666 8871 1718
rect 10779 1762 10785 1814
rect 10837 1762 10853 1814
rect 10905 1762 10921 1814
rect 10973 1762 10979 1814
rect 10779 1718 10979 1762
rect 10779 1666 10785 1718
rect 10837 1666 10853 1718
rect 10905 1666 10921 1718
rect 10973 1666 10979 1718
rect 13503 1762 13509 1814
rect 13561 1762 13577 1814
rect 13629 1762 13645 1814
rect 13697 1762 13703 1814
rect 13503 1718 13703 1762
rect 13503 1666 13509 1718
rect 13561 1666 13577 1718
rect 13629 1666 13645 1718
rect 13697 1666 13703 1718
rect 15611 1762 15617 1814
rect 15669 1762 15685 1814
rect 15737 1762 15753 1814
rect 15805 1762 15811 1814
rect 15611 1718 15811 1762
rect 15611 1666 15617 1718
rect 15669 1666 15685 1718
rect 15737 1666 15753 1718
rect 15805 1666 15811 1718
rect 18335 1762 18341 1814
rect 18393 1762 18409 1814
rect 18461 1762 18477 1814
rect 18529 1762 18535 1814
rect 18335 1718 18535 1762
rect 18335 1666 18341 1718
rect 18393 1666 18409 1718
rect 18461 1666 18477 1718
rect 18529 1666 18535 1718
rect 20443 1762 20449 1814
rect 20501 1762 20517 1814
rect 20569 1762 20585 1814
rect 20637 1762 20643 1814
rect 20443 1718 20643 1762
rect 20443 1666 20449 1718
rect 20501 1666 20517 1718
rect 20569 1666 20585 1718
rect 20637 1666 20643 1718
rect 23167 1762 23173 1814
rect 23225 1762 23241 1814
rect 23293 1762 23309 1814
rect 23361 1762 23367 1814
rect 23167 1718 23367 1762
rect 23167 1666 23173 1718
rect 23225 1666 23241 1718
rect 23293 1666 23309 1718
rect 23361 1666 23367 1718
rect 25275 1762 25281 1814
rect 25333 1762 25349 1814
rect 25401 1762 25417 1814
rect 25469 1762 25475 1814
rect 25275 1718 25475 1762
rect 25275 1666 25281 1718
rect 25333 1666 25349 1718
rect 25401 1666 25417 1718
rect 25469 1666 25475 1718
rect 27999 1762 28005 1814
rect 28057 1762 28073 1814
rect 28125 1762 28141 1814
rect 28193 1762 28199 1814
rect 27999 1718 28199 1762
rect 27999 1666 28005 1718
rect 28057 1666 28073 1718
rect 28125 1666 28141 1718
rect 28193 1666 28199 1718
rect 30107 1762 30113 1814
rect 30165 1762 30181 1814
rect 30233 1762 30249 1814
rect 30301 1762 30307 1814
rect 30107 1718 30307 1762
rect 30107 1666 30113 1718
rect 30165 1666 30181 1718
rect 30233 1666 30249 1718
rect 30301 1666 30307 1718
rect 32831 1762 32837 1814
rect 32889 1762 32905 1814
rect 32957 1762 32973 1814
rect 33025 1762 33031 1814
rect 32831 1718 33031 1762
rect 32831 1666 32837 1718
rect 32889 1666 32905 1718
rect 32957 1666 32973 1718
rect 33025 1666 33031 1718
rect 34939 1762 34945 1814
rect 34997 1762 35013 1814
rect 35065 1762 35081 1814
rect 35133 1762 35139 1814
rect 34939 1718 35139 1762
rect 34939 1666 34945 1718
rect 34997 1666 35013 1718
rect 35065 1666 35081 1718
rect 35133 1666 35139 1718
rect 37663 1762 37669 1814
rect 37721 1762 37737 1814
rect 37789 1762 37805 1814
rect 37857 1762 37863 1814
rect 37663 1718 37863 1762
rect 37663 1666 37669 1718
rect 37721 1666 37737 1718
rect 37789 1666 37805 1718
rect 37857 1666 37863 1718
rect 0 1586 614 1638
rect 666 1586 678 1638
rect 730 1586 4241 1638
rect 4293 1586 4305 1638
rect 4357 1586 5446 1638
rect 5498 1586 5510 1638
rect 5562 1586 9073 1638
rect 9125 1586 9137 1638
rect 9189 1586 10278 1638
rect 10330 1586 10342 1638
rect 10394 1586 13905 1638
rect 13957 1586 13969 1638
rect 14021 1586 15110 1638
rect 15162 1586 15174 1638
rect 15226 1586 18737 1638
rect 18789 1586 18801 1638
rect 18853 1586 19869 1638
rect 19921 1586 19933 1638
rect 19985 1586 23566 1638
rect 23618 1586 23630 1638
rect 23682 1586 24704 1638
rect 24756 1586 24768 1638
rect 24820 1586 28401 1638
rect 28453 1586 28465 1638
rect 28517 1586 29536 1638
rect 29588 1586 29600 1638
rect 29652 1586 33233 1638
rect 33285 1586 33297 1638
rect 33349 1586 34365 1638
rect 34417 1586 34429 1638
rect 34481 1586 38065 1638
rect 38117 1586 38129 1638
rect 38181 1586 38722 1638
rect 0 1506 20023 1558
rect 20075 1506 20087 1558
rect 20139 1506 23415 1558
rect 23467 1506 23479 1558
rect 23531 1506 24855 1558
rect 24907 1506 24919 1558
rect 24971 1506 28247 1558
rect 28299 1506 28311 1558
rect 28363 1506 29687 1558
rect 29739 1506 29751 1558
rect 29803 1506 33079 1558
rect 33131 1506 33143 1558
rect 33195 1506 34519 1558
rect 34571 1506 34583 1558
rect 34635 1506 37911 1558
rect 37963 1506 37975 1558
rect 38027 1506 38722 1558
rect 0 1426 10049 1478
rect 10101 1426 10113 1478
rect 10165 1426 13985 1478
rect 14037 1426 14049 1478
rect 14101 1426 14881 1478
rect 14933 1426 14945 1478
rect 14997 1426 18893 1478
rect 18945 1426 18957 1478
rect 19009 1426 29377 1478
rect 29429 1426 29441 1478
rect 29493 1426 33389 1478
rect 33441 1426 33453 1478
rect 33505 1426 34209 1478
rect 34261 1426 34273 1478
rect 34325 1426 38221 1478
rect 38273 1426 38285 1478
rect 38337 1426 38722 1478
rect 0 1346 5060 1398
rect 5112 1346 5124 1398
rect 5176 1346 9386 1398
rect 9438 1346 9450 1398
rect 9502 1346 14724 1398
rect 14776 1346 14788 1398
rect 14840 1346 19050 1398
rect 19102 1346 19114 1398
rect 19166 1346 24388 1398
rect 24440 1346 24452 1398
rect 24504 1346 28714 1398
rect 28766 1346 28778 1398
rect 28830 1346 34052 1398
rect 34104 1346 34116 1398
rect 34168 1346 38378 1398
rect 38430 1346 38442 1398
rect 38494 1346 38722 1398
rect 0 1266 4710 1318
rect 4762 1266 4774 1318
rect 4826 1266 9542 1318
rect 9594 1266 9606 1318
rect 9658 1266 14298 1318
rect 14350 1266 14362 1318
rect 14414 1266 19206 1318
rect 19258 1266 19270 1318
rect 19322 1266 24038 1318
rect 24090 1266 24102 1318
rect 24154 1266 28870 1318
rect 28922 1266 28934 1318
rect 28986 1266 33702 1318
rect 33754 1266 33766 1318
rect 33818 1266 38534 1318
rect 38586 1266 38598 1318
rect 38650 1266 38722 1318
rect 0 1186 539 1238
rect 591 1186 603 1238
rect 655 1186 4242 1238
rect 4294 1186 4306 1238
rect 4358 1186 5374 1238
rect 5426 1186 5438 1238
rect 5490 1186 9072 1238
rect 9124 1186 9136 1238
rect 9188 1186 10205 1238
rect 10257 1186 10269 1238
rect 10321 1186 13904 1238
rect 13956 1186 13968 1238
rect 14020 1186 15037 1238
rect 15089 1186 15101 1238
rect 15153 1186 18737 1238
rect 18789 1186 18801 1238
rect 18853 1186 19869 1238
rect 19921 1186 19933 1238
rect 19985 1186 23569 1238
rect 23621 1186 23633 1238
rect 23685 1186 24701 1238
rect 24753 1186 24765 1238
rect 24817 1186 28401 1238
rect 28453 1186 28465 1238
rect 28517 1186 29607 1238
rect 29659 1186 29671 1238
rect 29723 1186 33233 1238
rect 33285 1186 33297 1238
rect 33349 1186 34439 1238
rect 34491 1186 34503 1238
rect 34555 1186 38065 1238
rect 38117 1186 38129 1238
rect 38181 1186 38722 1238
rect 0 1106 695 1158
rect 747 1106 759 1158
rect 811 1106 4084 1158
rect 4136 1106 4148 1158
rect 4200 1106 5530 1158
rect 5582 1106 5594 1158
rect 5646 1106 8916 1158
rect 8968 1106 8980 1158
rect 9032 1106 10362 1158
rect 10414 1106 10426 1158
rect 10478 1106 13748 1158
rect 13800 1106 13812 1158
rect 13864 1106 15194 1158
rect 15246 1106 15258 1158
rect 15310 1106 18580 1158
rect 18632 1106 18644 1158
rect 18696 1106 38722 1158
rect 0 1026 459 1078
rect 511 1026 523 1078
rect 575 1026 4398 1078
rect 4450 1026 4462 1078
rect 4514 1026 5217 1078
rect 5269 1026 5281 1078
rect 5333 1026 9229 1078
rect 9281 1026 9293 1078
rect 9345 1026 19713 1078
rect 19765 1026 19777 1078
rect 19829 1026 23725 1078
rect 23777 1026 23789 1078
rect 23841 1026 24545 1078
rect 24597 1026 24609 1078
rect 24661 1026 28557 1078
rect 28609 1026 28621 1078
rect 28673 1026 38722 1078
rect 0 946 230 998
rect 282 946 294 998
rect 346 946 4554 998
rect 4606 946 4618 998
rect 4670 946 9892 998
rect 9944 946 9956 998
rect 10008 946 14142 998
rect 14194 946 14206 998
rect 14258 946 19556 998
rect 19608 946 19620 998
rect 19672 946 23882 998
rect 23934 946 23946 998
rect 23998 946 29220 998
rect 29272 946 29284 998
rect 29336 946 33546 998
rect 33598 946 33610 998
rect 33662 946 38722 998
rect 0 866 74 918
rect 126 866 138 918
rect 190 866 4904 918
rect 4956 866 4968 918
rect 5020 866 9736 918
rect 9788 866 9800 918
rect 9852 866 14568 918
rect 14620 866 14632 918
rect 14684 866 19400 918
rect 19452 866 19464 918
rect 19516 866 24232 918
rect 24284 866 24296 918
rect 24348 866 29064 918
rect 29116 866 29128 918
rect 29180 866 33896 918
rect 33948 866 33960 918
rect 34012 866 38722 918
rect 1115 786 1121 838
rect 1173 786 1189 838
rect 1241 786 1257 838
rect 1309 786 1315 838
rect 1115 742 1315 786
rect 1115 690 1121 742
rect 1173 690 1189 742
rect 1241 690 1257 742
rect 1309 690 1315 742
rect 3839 690 4039 838
rect 5947 786 5953 838
rect 6005 786 6021 838
rect 6073 786 6089 838
rect 6141 786 6147 838
rect 5947 742 6147 786
rect 5947 690 5953 742
rect 6005 690 6021 742
rect 6073 690 6089 742
rect 6141 690 6147 742
rect 8671 786 8677 838
rect 8729 786 8745 838
rect 8797 786 8813 838
rect 8865 786 8871 838
rect 8671 742 8871 786
rect 8671 690 8677 742
rect 8729 690 8745 742
rect 8797 690 8813 742
rect 8865 690 8871 742
rect 10779 786 10785 838
rect 10837 786 10853 838
rect 10905 786 10921 838
rect 10973 786 10979 838
rect 10779 742 10979 786
rect 10779 690 10785 742
rect 10837 690 10853 742
rect 10905 690 10921 742
rect 10973 690 10979 742
rect 13503 786 13509 838
rect 13561 786 13577 838
rect 13629 786 13645 838
rect 13697 786 13703 838
rect 13503 742 13703 786
rect 13503 690 13509 742
rect 13561 690 13577 742
rect 13629 690 13645 742
rect 13697 690 13703 742
rect 15611 786 15617 838
rect 15669 786 15685 838
rect 15737 786 15753 838
rect 15805 786 15811 838
rect 15611 742 15811 786
rect 15611 690 15617 742
rect 15669 690 15685 742
rect 15737 690 15753 742
rect 15805 690 15811 742
rect 18335 786 18341 838
rect 18393 786 18409 838
rect 18461 786 18477 838
rect 18529 786 18535 838
rect 18335 742 18535 786
rect 18335 690 18341 742
rect 18393 690 18409 742
rect 18461 690 18477 742
rect 18529 690 18535 742
rect 20443 786 20449 838
rect 20501 786 20517 838
rect 20569 786 20585 838
rect 20637 786 20643 838
rect 20443 742 20643 786
rect 20443 690 20449 742
rect 20501 690 20517 742
rect 20569 690 20585 742
rect 20637 690 20643 742
rect 23167 786 23173 838
rect 23225 786 23241 838
rect 23293 786 23309 838
rect 23361 786 23367 838
rect 23167 742 23367 786
rect 23167 690 23173 742
rect 23225 690 23241 742
rect 23293 690 23309 742
rect 23361 690 23367 742
rect 25275 786 25281 838
rect 25333 786 25349 838
rect 25401 786 25417 838
rect 25469 786 25475 838
rect 25275 742 25475 786
rect 25275 690 25281 742
rect 25333 690 25349 742
rect 25401 690 25417 742
rect 25469 690 25475 742
rect 27999 786 28005 838
rect 28057 786 28073 838
rect 28125 786 28141 838
rect 28193 786 28199 838
rect 27999 742 28199 786
rect 27999 690 28005 742
rect 28057 690 28073 742
rect 28125 690 28141 742
rect 28193 690 28199 742
rect 30107 786 30113 838
rect 30165 786 30181 838
rect 30233 786 30249 838
rect 30301 786 30307 838
rect 30107 742 30307 786
rect 30107 690 30113 742
rect 30165 690 30181 742
rect 30233 690 30249 742
rect 30301 690 30307 742
rect 32831 786 32837 838
rect 32889 786 32905 838
rect 32957 786 32973 838
rect 33025 786 33031 838
rect 32831 742 33031 786
rect 32831 690 32837 742
rect 32889 690 32905 742
rect 32957 690 32973 742
rect 33025 690 33031 742
rect 34939 786 34945 838
rect 34997 786 35013 838
rect 35065 786 35081 838
rect 35133 786 35139 838
rect 34939 742 35139 786
rect 34939 690 34945 742
rect 34997 690 35013 742
rect 35065 690 35081 742
rect 35133 690 35139 742
rect 37663 786 37669 838
rect 37721 786 37737 838
rect 37789 786 37805 838
rect 37857 786 37863 838
rect 37663 742 37863 786
rect 37663 690 37669 742
rect 37721 690 37737 742
rect 37789 690 37805 742
rect 37857 690 37863 742
rect 144 463 196 469
rect 144 397 196 411
rect 144 339 196 345
rect 300 463 352 469
rect 300 397 352 411
rect 300 339 352 345
rect 453 463 505 469
rect 453 397 505 411
rect 453 339 505 345
rect 609 457 661 463
rect 609 391 661 405
rect 609 333 661 339
rect 765 460 817 471
rect 765 396 817 408
rect 765 338 817 344
rect 4078 465 4130 471
rect 4392 463 4444 469
rect 4078 399 4130 413
rect 4078 341 4130 347
rect 4236 457 4288 463
rect 4236 391 4288 405
rect 4392 397 4444 411
rect 4392 339 4444 345
rect 4548 463 4600 469
rect 4548 397 4600 411
rect 4548 339 4600 345
rect 4704 463 4756 469
rect 4704 397 4756 411
rect 4704 339 4756 345
rect 4974 463 5026 469
rect 4974 397 5026 411
rect 4974 339 5026 345
rect 5130 463 5182 469
rect 5130 397 5182 411
rect 5130 339 5182 345
rect 5287 463 5339 469
rect 5600 465 5652 471
rect 5287 397 5339 411
rect 5287 339 5339 345
rect 5444 457 5496 463
rect 5444 391 5496 405
rect 5600 399 5652 413
rect 5600 341 5652 347
rect 8910 465 8962 471
rect 9223 463 9275 469
rect 8910 399 8962 413
rect 8910 341 8962 347
rect 9066 457 9118 463
rect 9066 391 9118 405
rect 4236 333 4288 339
rect 5444 333 5496 339
rect 9223 397 9275 411
rect 9223 339 9275 345
rect 9380 463 9432 469
rect 9380 397 9432 411
rect 9380 339 9432 345
rect 9536 463 9588 469
rect 9536 397 9588 411
rect 9536 339 9588 345
rect 9806 463 9858 469
rect 9806 397 9858 411
rect 9806 339 9858 345
rect 9962 463 10014 469
rect 9962 397 10014 411
rect 9962 339 10014 345
rect 10119 463 10171 469
rect 10119 397 10171 411
rect 10119 339 10171 345
rect 10275 461 10327 467
rect 10275 391 10327 409
rect 10432 465 10484 471
rect 10432 399 10484 413
rect 10432 341 10484 347
rect 13742 465 13794 471
rect 13742 399 13794 413
rect 13742 341 13794 347
rect 13898 461 13950 467
rect 13898 391 13950 409
rect 9066 333 9118 339
rect 10275 333 10327 339
rect 14055 463 14107 469
rect 14055 397 14107 411
rect 14055 339 14107 345
rect 14212 463 14264 469
rect 14212 397 14264 411
rect 14212 339 14264 345
rect 14368 463 14420 469
rect 14368 397 14420 411
rect 14368 339 14420 345
rect 14638 463 14690 469
rect 14638 397 14690 411
rect 14638 339 14690 345
rect 14794 463 14846 469
rect 14794 397 14846 411
rect 14794 339 14846 345
rect 14951 463 15003 469
rect 14951 397 15003 411
rect 14951 339 15003 345
rect 15107 461 15159 467
rect 15107 391 15159 409
rect 15264 465 15316 471
rect 15264 399 15316 413
rect 15264 341 15316 347
rect 18574 465 18626 471
rect 18574 399 18626 413
rect 18574 341 18626 347
rect 18731 461 18783 467
rect 18731 391 18783 409
rect 13898 333 13950 339
rect 15107 333 15159 339
rect 18887 463 18939 469
rect 18887 397 18939 411
rect 18887 339 18939 345
rect 19044 463 19096 469
rect 19044 397 19096 411
rect 19044 339 19096 345
rect 19200 463 19252 469
rect 19200 397 19252 411
rect 19200 339 19252 345
rect 19470 463 19522 469
rect 19470 397 19522 411
rect 19470 339 19522 345
rect 19626 463 19678 469
rect 19626 397 19678 411
rect 19626 339 19678 345
rect 19783 463 19835 469
rect 19783 397 19835 411
rect 19783 339 19835 345
rect 19939 461 19991 467
rect 19939 391 19991 409
rect 20093 461 20145 471
rect 20093 397 20145 409
rect 20093 339 20145 345
rect 23409 461 23461 471
rect 23409 397 23461 409
rect 23409 339 23461 345
rect 23563 461 23615 467
rect 23563 391 23615 409
rect 23719 463 23771 469
rect 23719 397 23771 411
rect 23719 339 23771 345
rect 23876 463 23928 469
rect 23876 397 23928 411
rect 23876 339 23928 345
rect 24032 463 24084 469
rect 24032 397 24084 411
rect 24032 339 24084 345
rect 24302 463 24354 469
rect 24302 397 24354 411
rect 24302 339 24354 345
rect 24458 463 24510 469
rect 24458 397 24510 411
rect 24458 339 24510 345
rect 24615 463 24667 469
rect 24615 397 24667 411
rect 24615 339 24667 345
rect 24771 461 24823 467
rect 24771 391 24823 409
rect 24925 461 24977 471
rect 24925 397 24977 409
rect 24925 339 24977 345
rect 28241 465 28293 471
rect 28241 397 28293 413
rect 28241 339 28293 345
rect 28395 461 28447 467
rect 28395 391 28447 409
rect 28551 463 28603 469
rect 28551 397 28603 411
rect 28551 339 28603 345
rect 28708 463 28760 469
rect 28708 397 28760 411
rect 28708 339 28760 345
rect 28864 463 28916 469
rect 28864 397 28916 411
rect 28864 339 28916 345
rect 29134 463 29186 469
rect 29134 397 29186 411
rect 29134 339 29186 345
rect 29290 463 29342 469
rect 29290 397 29342 411
rect 29290 339 29342 345
rect 29447 463 29499 469
rect 29447 397 29499 411
rect 29447 339 29499 345
rect 29601 461 29653 467
rect 29601 391 29653 409
rect 29757 465 29809 471
rect 29757 397 29809 413
rect 29757 339 29809 345
rect 33073 465 33125 471
rect 33073 397 33125 413
rect 33073 339 33125 345
rect 33227 461 33279 467
rect 33227 391 33279 409
rect 33383 463 33435 469
rect 33383 397 33435 411
rect 33383 339 33435 345
rect 33540 463 33592 469
rect 33540 397 33592 411
rect 33540 339 33592 345
rect 33696 463 33748 469
rect 33696 397 33748 411
rect 33696 339 33748 345
rect 33966 463 34018 469
rect 33966 397 34018 411
rect 33966 339 34018 345
rect 34122 463 34174 469
rect 34122 397 34174 411
rect 34122 339 34174 345
rect 34279 463 34331 469
rect 34279 397 34331 411
rect 34279 339 34331 345
rect 34433 461 34485 467
rect 34433 391 34485 409
rect 34589 465 34641 471
rect 34589 397 34641 413
rect 34589 339 34641 345
rect 37905 465 37957 471
rect 37905 397 37957 413
rect 37905 339 37957 345
rect 38059 461 38111 467
rect 38059 391 38111 409
rect 38215 463 38267 469
rect 38215 397 38267 411
rect 38215 339 38267 345
rect 38372 463 38424 469
rect 38372 397 38424 411
rect 38372 339 38424 345
rect 38528 463 38580 469
rect 38528 397 38580 411
rect 38528 339 38580 345
rect 18731 333 18783 339
rect 19939 333 19991 339
rect 23563 333 23615 339
rect 24771 333 24823 339
rect 28395 333 28447 339
rect 29601 333 29653 339
rect 33227 333 33279 339
rect 34433 333 34485 339
rect 38059 333 38111 339
rect 2124 232 2237 267
rect 2674 234 2791 263
rect 6945 235 7086 266
rect 7494 232 7638 268
rect 11774 233 11909 266
rect 12309 230 12442 264
rect 16597 229 16731 264
rect 17164 230 17285 266
rect 21433 230 21570 267
rect 21971 228 22118 266
rect 26273 229 26417 266
rect 26789 230 26937 271
rect 31126 231 31273 266
rect 31613 232 31774 269
rect 35941 230 36095 268
rect 36461 229 36598 265
rect 859 112 865 164
rect 917 112 933 164
rect 985 112 1001 164
rect 1053 112 1059 164
rect 859 52 1059 112
rect 859 0 865 52
rect 917 0 933 52
rect 985 0 1001 52
rect 1053 0 1059 52
rect 5691 112 5697 164
rect 5749 112 5765 164
rect 5817 112 5833 164
rect 5885 112 5891 164
rect 5691 52 5891 112
rect 5691 0 5697 52
rect 5749 0 5765 52
rect 5817 0 5833 52
rect 5885 0 5891 52
rect 8415 112 8421 164
rect 8473 112 8489 164
rect 8541 112 8557 164
rect 8609 112 8615 164
rect 8415 52 8615 112
rect 8415 0 8421 52
rect 8473 0 8489 52
rect 8541 0 8557 52
rect 8609 0 8615 52
rect 10523 112 10529 164
rect 10581 112 10597 164
rect 10649 112 10665 164
rect 10717 112 10723 164
rect 10523 52 10723 112
rect 10523 0 10529 52
rect 10581 0 10597 52
rect 10649 0 10665 52
rect 10717 0 10723 52
rect 13247 112 13253 164
rect 13305 112 13321 164
rect 13373 112 13389 164
rect 13441 112 13447 164
rect 13247 52 13447 112
rect 13247 0 13253 52
rect 13305 0 13321 52
rect 13373 0 13389 52
rect 13441 0 13447 52
rect 15355 112 15361 164
rect 15413 112 15429 164
rect 15481 112 15497 164
rect 15549 112 15555 164
rect 15355 52 15555 112
rect 15355 0 15361 52
rect 15413 0 15429 52
rect 15481 0 15497 52
rect 15549 0 15555 52
rect 18079 112 18085 164
rect 18137 112 18153 164
rect 18205 112 18221 164
rect 18273 112 18279 164
rect 18079 52 18279 112
rect 18079 0 18085 52
rect 18137 0 18153 52
rect 18205 0 18221 52
rect 18273 0 18279 52
rect 20187 112 20193 164
rect 20245 112 20261 164
rect 20313 112 20329 164
rect 20381 112 20387 164
rect 20187 52 20387 112
rect 20187 0 20193 52
rect 20245 0 20261 52
rect 20313 0 20329 52
rect 20381 0 20387 52
rect 22911 112 22917 164
rect 22969 112 22985 164
rect 23037 112 23053 164
rect 23105 112 23111 164
rect 22911 52 23111 112
rect 22911 0 22917 52
rect 22969 0 22985 52
rect 23037 0 23053 52
rect 23105 0 23111 52
rect 25019 112 25025 164
rect 25077 112 25093 164
rect 25145 112 25161 164
rect 25213 112 25219 164
rect 25019 52 25219 112
rect 25019 0 25025 52
rect 25077 0 25093 52
rect 25145 0 25161 52
rect 25213 0 25219 52
rect 27743 112 27749 164
rect 27801 112 27817 164
rect 27869 112 27885 164
rect 27937 112 27943 164
rect 27743 52 27943 112
rect 27743 0 27749 52
rect 27801 0 27817 52
rect 27869 0 27885 52
rect 27937 0 27943 52
rect 29851 112 29857 164
rect 29909 112 29925 164
rect 29977 112 29993 164
rect 30045 112 30051 164
rect 29851 52 30051 112
rect 29851 0 29857 52
rect 29909 0 29925 52
rect 29977 0 29993 52
rect 30045 0 30051 52
rect 32575 112 32581 164
rect 32633 112 32649 164
rect 32701 112 32717 164
rect 32769 112 32775 164
rect 32575 52 32775 112
rect 32575 0 32581 52
rect 32633 0 32649 52
rect 32701 0 32717 52
rect 32769 0 32775 52
rect 34683 112 34689 164
rect 34741 112 34757 164
rect 34809 112 34825 164
rect 34877 112 34883 164
rect 34683 52 34883 112
rect 34683 0 34689 52
rect 34741 0 34757 52
rect 34809 0 34825 52
rect 34877 0 34883 52
rect 37407 112 37413 164
rect 37465 112 37481 164
rect 37533 112 37549 164
rect 37601 112 37607 164
rect 37407 52 37607 112
rect 37407 0 37413 52
rect 37465 0 37481 52
rect 37533 0 37549 52
rect 37601 0 37607 52
rect 0 -80 2249 -28
rect 2301 -80 2313 -28
rect 2365 -80 2533 -28
rect 2585 -80 2597 -28
rect 2649 -80 7081 -28
rect 7133 -80 7145 -28
rect 7197 -80 7365 -28
rect 7417 -80 7429 -28
rect 7481 -80 11913 -28
rect 11965 -80 11977 -28
rect 12029 -80 12197 -28
rect 12249 -80 12261 -28
rect 12313 -80 16745 -28
rect 16797 -80 16809 -28
rect 16861 -80 17029 -28
rect 17081 -80 17093 -28
rect 17145 -80 21577 -28
rect 21629 -80 21641 -28
rect 21693 -80 21861 -28
rect 21913 -80 21925 -28
rect 21977 -80 26409 -28
rect 26461 -80 26473 -28
rect 26525 -80 26693 -28
rect 26745 -80 26757 -28
rect 26809 -80 31241 -28
rect 31293 -80 31305 -28
rect 31357 -80 31525 -28
rect 31577 -80 31589 -28
rect 31641 -80 36073 -28
rect 36125 -80 36137 -28
rect 36189 -80 36357 -28
rect 36409 -80 36421 -28
rect 36473 -80 38722 -28
rect 0 -160 38722 -108
<< via1 >>
rect 2249 2588 2301 2640
rect 2313 2588 2365 2640
rect 2533 2588 2585 2640
rect 2597 2588 2649 2640
rect 7081 2588 7133 2640
rect 7145 2588 7197 2640
rect 7365 2588 7417 2640
rect 7429 2588 7481 2640
rect 11913 2588 11965 2640
rect 11977 2588 12029 2640
rect 12197 2588 12249 2640
rect 12261 2588 12313 2640
rect 16745 2588 16797 2640
rect 16809 2588 16861 2640
rect 17029 2588 17081 2640
rect 17093 2588 17145 2640
rect 21577 2588 21629 2640
rect 21641 2588 21693 2640
rect 21861 2588 21913 2640
rect 21925 2588 21977 2640
rect 26409 2588 26461 2640
rect 26473 2588 26525 2640
rect 26693 2588 26745 2640
rect 26757 2588 26809 2640
rect 31241 2588 31293 2640
rect 31305 2588 31357 2640
rect 31525 2588 31577 2640
rect 31589 2588 31641 2640
rect 36073 2588 36125 2640
rect 36137 2588 36189 2640
rect 36357 2588 36409 2640
rect 36421 2588 36473 2640
rect 865 2452 917 2504
rect 933 2452 985 2504
rect 1001 2452 1053 2504
rect 865 2340 917 2392
rect 933 2340 985 2392
rect 1001 2340 1053 2392
rect 5697 2452 5749 2504
rect 5765 2452 5817 2504
rect 5833 2452 5885 2504
rect 5697 2340 5749 2392
rect 5765 2340 5817 2392
rect 5833 2340 5885 2392
rect 8421 2452 8473 2504
rect 8489 2452 8541 2504
rect 8557 2452 8609 2504
rect 8421 2340 8473 2392
rect 8489 2340 8541 2392
rect 8557 2340 8609 2392
rect 10529 2452 10581 2504
rect 10597 2452 10649 2504
rect 10665 2452 10717 2504
rect 10529 2340 10581 2392
rect 10597 2340 10649 2392
rect 10665 2340 10717 2392
rect 13253 2452 13305 2504
rect 13321 2452 13373 2504
rect 13389 2452 13441 2504
rect 13253 2340 13305 2392
rect 13321 2340 13373 2392
rect 13389 2340 13441 2392
rect 15361 2452 15413 2504
rect 15429 2452 15481 2504
rect 15497 2452 15549 2504
rect 15361 2340 15413 2392
rect 15429 2340 15481 2392
rect 15497 2340 15549 2392
rect 18085 2452 18137 2504
rect 18153 2452 18205 2504
rect 18221 2452 18273 2504
rect 18085 2340 18137 2392
rect 18153 2340 18205 2392
rect 18221 2340 18273 2392
rect 20193 2452 20245 2504
rect 20261 2452 20313 2504
rect 20329 2452 20381 2504
rect 20193 2340 20245 2392
rect 20261 2340 20313 2392
rect 20329 2340 20381 2392
rect 22917 2452 22969 2504
rect 22985 2452 23037 2504
rect 23053 2452 23105 2504
rect 22917 2340 22969 2392
rect 22985 2340 23037 2392
rect 23053 2340 23105 2392
rect 25025 2452 25077 2504
rect 25093 2452 25145 2504
rect 25161 2452 25213 2504
rect 25025 2340 25077 2392
rect 25093 2340 25145 2392
rect 25161 2340 25213 2392
rect 27749 2452 27801 2504
rect 27817 2452 27869 2504
rect 27885 2452 27937 2504
rect 27749 2340 27801 2392
rect 27817 2340 27869 2392
rect 27885 2340 27937 2392
rect 29857 2452 29909 2504
rect 29925 2452 29977 2504
rect 29993 2452 30045 2504
rect 29857 2340 29909 2392
rect 29925 2340 29977 2392
rect 29993 2340 30045 2392
rect 32581 2452 32633 2504
rect 32649 2452 32701 2504
rect 32717 2452 32769 2504
rect 32581 2340 32633 2392
rect 32649 2340 32701 2392
rect 32717 2340 32769 2392
rect 34689 2452 34741 2504
rect 34757 2452 34809 2504
rect 34825 2452 34877 2504
rect 34689 2340 34741 2392
rect 34757 2340 34809 2392
rect 34825 2340 34877 2392
rect 37413 2452 37465 2504
rect 37481 2452 37533 2504
rect 37549 2452 37601 2504
rect 37413 2340 37465 2392
rect 37481 2340 37533 2392
rect 37549 2340 37601 2392
rect 144 2107 196 2159
rect 144 2041 196 2093
rect 300 2107 352 2159
rect 300 2041 352 2093
rect 453 2107 505 2159
rect 453 2041 505 2093
rect 608 2108 660 2160
rect 608 2044 660 2096
rect 765 2107 817 2159
rect 765 2043 817 2095
rect 4078 2103 4130 2155
rect 4078 2039 4130 2091
rect 4235 2108 4287 2160
rect 4235 2044 4287 2096
rect 4392 2107 4444 2159
rect 4392 2041 4444 2093
rect 4548 2107 4600 2159
rect 4548 2041 4600 2093
rect 4704 2107 4756 2159
rect 4704 2043 4756 2095
rect 4974 2107 5026 2159
rect 4974 2041 5026 2093
rect 5130 2107 5182 2159
rect 5130 2041 5182 2093
rect 5287 2107 5339 2159
rect 5287 2041 5339 2093
rect 5440 2108 5492 2160
rect 5440 2044 5492 2096
rect 5600 2105 5652 2157
rect 5600 2039 5652 2091
rect 8910 2105 8962 2157
rect 8910 2039 8962 2091
rect 9067 2113 9119 2165
rect 9067 2044 9119 2096
rect 9223 2107 9275 2159
rect 9223 2041 9275 2093
rect 9380 2107 9432 2159
rect 9380 2041 9432 2093
rect 9536 2107 9588 2159
rect 9536 2041 9588 2093
rect 9806 2107 9858 2159
rect 9806 2041 9858 2093
rect 9962 2107 10014 2159
rect 9962 2041 10014 2093
rect 10119 2107 10171 2159
rect 10119 2041 10171 2093
rect 10272 2108 10324 2160
rect 10272 2044 10324 2096
rect 10432 2105 10484 2157
rect 10432 2039 10484 2091
rect 13742 2105 13794 2157
rect 13742 2039 13794 2091
rect 13899 2113 13951 2165
rect 13899 2044 13951 2096
rect 14055 2107 14107 2159
rect 14055 2041 14107 2093
rect 14212 2107 14264 2159
rect 14212 2041 14264 2093
rect 14368 2107 14420 2159
rect 14368 2041 14420 2093
rect 14638 2107 14690 2159
rect 14638 2041 14690 2093
rect 14794 2107 14846 2159
rect 14794 2041 14846 2093
rect 14951 2107 15003 2159
rect 14951 2041 15003 2093
rect 15104 2108 15156 2160
rect 15104 2044 15156 2096
rect 15264 2105 15316 2157
rect 15264 2039 15316 2091
rect 18574 2105 18626 2157
rect 18574 2039 18626 2091
rect 18731 2113 18783 2165
rect 18731 2044 18783 2096
rect 18887 2107 18939 2159
rect 18887 2041 18939 2093
rect 19044 2107 19096 2159
rect 19044 2041 19096 2093
rect 19200 2107 19252 2159
rect 19200 2041 19252 2093
rect 19470 2107 19522 2159
rect 19470 2041 19522 2093
rect 19626 2107 19678 2159
rect 19626 2041 19678 2093
rect 19783 2107 19835 2159
rect 19783 2041 19835 2093
rect 19939 2113 19991 2165
rect 19939 2044 19991 2096
rect 20093 2107 20145 2159
rect 20093 2043 20145 2095
rect 23409 2107 23461 2159
rect 23409 2043 23461 2095
rect 23560 2108 23612 2160
rect 23560 2044 23612 2096
rect 23719 2107 23771 2159
rect 23719 2041 23771 2093
rect 23876 2107 23928 2159
rect 23876 2041 23928 2093
rect 24032 2107 24084 2159
rect 24032 2041 24084 2093
rect 24302 2107 24354 2159
rect 24302 2041 24354 2093
rect 24458 2107 24510 2159
rect 24458 2041 24510 2093
rect 24615 2107 24667 2159
rect 24615 2041 24667 2093
rect 24774 2113 24826 2165
rect 24774 2044 24826 2096
rect 24925 2107 24977 2159
rect 24925 2043 24977 2095
rect 28241 2107 28293 2159
rect 28241 2039 28293 2091
rect 28395 2113 28447 2165
rect 28395 2044 28447 2096
rect 28551 2107 28603 2159
rect 28551 2041 28603 2093
rect 28708 2107 28760 2159
rect 28708 2041 28760 2093
rect 28864 2107 28916 2159
rect 28864 2041 28916 2093
rect 29134 2107 29186 2159
rect 29134 2041 29186 2093
rect 29290 2107 29342 2159
rect 29290 2041 29342 2093
rect 29447 2107 29499 2159
rect 29447 2041 29499 2093
rect 29606 2113 29658 2165
rect 29606 2044 29658 2096
rect 29757 2107 29809 2159
rect 29757 2039 29809 2091
rect 33073 2107 33125 2159
rect 33073 2039 33125 2091
rect 33227 2113 33279 2165
rect 33227 2044 33279 2096
rect 33383 2107 33435 2159
rect 33383 2041 33435 2093
rect 33540 2107 33592 2159
rect 33540 2041 33592 2093
rect 33696 2107 33748 2159
rect 33696 2041 33748 2093
rect 33966 2107 34018 2159
rect 33966 2041 34018 2093
rect 34122 2107 34174 2159
rect 34122 2041 34174 2093
rect 34279 2107 34331 2159
rect 34279 2041 34331 2093
rect 34435 2113 34487 2165
rect 34435 2044 34487 2096
rect 34589 2107 34641 2159
rect 34589 2039 34641 2091
rect 37905 2108 37957 2160
rect 37905 2039 37957 2091
rect 38059 2113 38111 2165
rect 38059 2044 38111 2096
rect 38215 2108 38267 2160
rect 38215 2041 38267 2093
rect 38372 2108 38424 2160
rect 38372 2041 38424 2093
rect 38528 2108 38580 2160
rect 38528 2041 38580 2093
rect 1121 1762 1173 1814
rect 1189 1762 1241 1814
rect 1257 1762 1309 1814
rect 1121 1666 1173 1718
rect 1189 1666 1241 1718
rect 1257 1666 1309 1718
rect 5953 1762 6005 1814
rect 6021 1762 6073 1814
rect 6089 1762 6141 1814
rect 5953 1666 6005 1718
rect 6021 1666 6073 1718
rect 6089 1666 6141 1718
rect 8677 1762 8729 1814
rect 8745 1762 8797 1814
rect 8813 1762 8865 1814
rect 8677 1666 8729 1718
rect 8745 1666 8797 1718
rect 8813 1666 8865 1718
rect 10785 1762 10837 1814
rect 10853 1762 10905 1814
rect 10921 1762 10973 1814
rect 10785 1666 10837 1718
rect 10853 1666 10905 1718
rect 10921 1666 10973 1718
rect 13509 1762 13561 1814
rect 13577 1762 13629 1814
rect 13645 1762 13697 1814
rect 13509 1666 13561 1718
rect 13577 1666 13629 1718
rect 13645 1666 13697 1718
rect 15617 1762 15669 1814
rect 15685 1762 15737 1814
rect 15753 1762 15805 1814
rect 15617 1666 15669 1718
rect 15685 1666 15737 1718
rect 15753 1666 15805 1718
rect 18341 1762 18393 1814
rect 18409 1762 18461 1814
rect 18477 1762 18529 1814
rect 18341 1666 18393 1718
rect 18409 1666 18461 1718
rect 18477 1666 18529 1718
rect 20449 1762 20501 1814
rect 20517 1762 20569 1814
rect 20585 1762 20637 1814
rect 20449 1666 20501 1718
rect 20517 1666 20569 1718
rect 20585 1666 20637 1718
rect 23173 1762 23225 1814
rect 23241 1762 23293 1814
rect 23309 1762 23361 1814
rect 23173 1666 23225 1718
rect 23241 1666 23293 1718
rect 23309 1666 23361 1718
rect 25281 1762 25333 1814
rect 25349 1762 25401 1814
rect 25417 1762 25469 1814
rect 25281 1666 25333 1718
rect 25349 1666 25401 1718
rect 25417 1666 25469 1718
rect 28005 1762 28057 1814
rect 28073 1762 28125 1814
rect 28141 1762 28193 1814
rect 28005 1666 28057 1718
rect 28073 1666 28125 1718
rect 28141 1666 28193 1718
rect 30113 1762 30165 1814
rect 30181 1762 30233 1814
rect 30249 1762 30301 1814
rect 30113 1666 30165 1718
rect 30181 1666 30233 1718
rect 30249 1666 30301 1718
rect 32837 1762 32889 1814
rect 32905 1762 32957 1814
rect 32973 1762 33025 1814
rect 32837 1666 32889 1718
rect 32905 1666 32957 1718
rect 32973 1666 33025 1718
rect 34945 1762 34997 1814
rect 35013 1762 35065 1814
rect 35081 1762 35133 1814
rect 34945 1666 34997 1718
rect 35013 1666 35065 1718
rect 35081 1666 35133 1718
rect 37669 1762 37721 1814
rect 37737 1762 37789 1814
rect 37805 1762 37857 1814
rect 37669 1666 37721 1718
rect 37737 1666 37789 1718
rect 37805 1666 37857 1718
rect 614 1586 666 1638
rect 678 1586 730 1638
rect 4241 1586 4293 1638
rect 4305 1586 4357 1638
rect 5446 1586 5498 1638
rect 5510 1586 5562 1638
rect 9073 1586 9125 1638
rect 9137 1586 9189 1638
rect 10278 1586 10330 1638
rect 10342 1586 10394 1638
rect 13905 1586 13957 1638
rect 13969 1586 14021 1638
rect 15110 1586 15162 1638
rect 15174 1586 15226 1638
rect 18737 1586 18789 1638
rect 18801 1586 18853 1638
rect 19869 1586 19921 1638
rect 19933 1586 19985 1638
rect 23566 1586 23618 1638
rect 23630 1586 23682 1638
rect 24704 1586 24756 1638
rect 24768 1586 24820 1638
rect 28401 1586 28453 1638
rect 28465 1586 28517 1638
rect 29536 1586 29588 1638
rect 29600 1586 29652 1638
rect 33233 1586 33285 1638
rect 33297 1586 33349 1638
rect 34365 1586 34417 1638
rect 34429 1586 34481 1638
rect 38065 1586 38117 1638
rect 38129 1586 38181 1638
rect 20023 1506 20075 1558
rect 20087 1506 20139 1558
rect 23415 1506 23467 1558
rect 23479 1506 23531 1558
rect 24855 1506 24907 1558
rect 24919 1506 24971 1558
rect 28247 1506 28299 1558
rect 28311 1506 28363 1558
rect 29687 1506 29739 1558
rect 29751 1506 29803 1558
rect 33079 1506 33131 1558
rect 33143 1506 33195 1558
rect 34519 1506 34571 1558
rect 34583 1506 34635 1558
rect 37911 1506 37963 1558
rect 37975 1506 38027 1558
rect 10049 1426 10101 1478
rect 10113 1426 10165 1478
rect 13985 1426 14037 1478
rect 14049 1426 14101 1478
rect 14881 1426 14933 1478
rect 14945 1426 14997 1478
rect 18893 1426 18945 1478
rect 18957 1426 19009 1478
rect 29377 1426 29429 1478
rect 29441 1426 29493 1478
rect 33389 1426 33441 1478
rect 33453 1426 33505 1478
rect 34209 1426 34261 1478
rect 34273 1426 34325 1478
rect 38221 1426 38273 1478
rect 38285 1426 38337 1478
rect 5060 1346 5112 1398
rect 5124 1346 5176 1398
rect 9386 1346 9438 1398
rect 9450 1346 9502 1398
rect 14724 1346 14776 1398
rect 14788 1346 14840 1398
rect 19050 1346 19102 1398
rect 19114 1346 19166 1398
rect 24388 1346 24440 1398
rect 24452 1346 24504 1398
rect 28714 1346 28766 1398
rect 28778 1346 28830 1398
rect 34052 1346 34104 1398
rect 34116 1346 34168 1398
rect 38378 1346 38430 1398
rect 38442 1346 38494 1398
rect 4710 1266 4762 1318
rect 4774 1266 4826 1318
rect 9542 1266 9594 1318
rect 9606 1266 9658 1318
rect 14298 1266 14350 1318
rect 14362 1266 14414 1318
rect 19206 1266 19258 1318
rect 19270 1266 19322 1318
rect 24038 1266 24090 1318
rect 24102 1266 24154 1318
rect 28870 1266 28922 1318
rect 28934 1266 28986 1318
rect 33702 1266 33754 1318
rect 33766 1266 33818 1318
rect 38534 1266 38586 1318
rect 38598 1266 38650 1318
rect 539 1186 591 1238
rect 603 1186 655 1238
rect 4242 1186 4294 1238
rect 4306 1186 4358 1238
rect 5374 1186 5426 1238
rect 5438 1186 5490 1238
rect 9072 1186 9124 1238
rect 9136 1186 9188 1238
rect 10205 1186 10257 1238
rect 10269 1186 10321 1238
rect 13904 1186 13956 1238
rect 13968 1186 14020 1238
rect 15037 1186 15089 1238
rect 15101 1186 15153 1238
rect 18737 1186 18789 1238
rect 18801 1186 18853 1238
rect 19869 1186 19921 1238
rect 19933 1186 19985 1238
rect 23569 1186 23621 1238
rect 23633 1186 23685 1238
rect 24701 1186 24753 1238
rect 24765 1186 24817 1238
rect 28401 1186 28453 1238
rect 28465 1186 28517 1238
rect 29607 1186 29659 1238
rect 29671 1186 29723 1238
rect 33233 1186 33285 1238
rect 33297 1186 33349 1238
rect 34439 1186 34491 1238
rect 34503 1186 34555 1238
rect 38065 1186 38117 1238
rect 38129 1186 38181 1238
rect 695 1106 747 1158
rect 759 1106 811 1158
rect 4084 1106 4136 1158
rect 4148 1106 4200 1158
rect 5530 1106 5582 1158
rect 5594 1106 5646 1158
rect 8916 1106 8968 1158
rect 8980 1106 9032 1158
rect 10362 1106 10414 1158
rect 10426 1106 10478 1158
rect 13748 1106 13800 1158
rect 13812 1106 13864 1158
rect 15194 1106 15246 1158
rect 15258 1106 15310 1158
rect 18580 1106 18632 1158
rect 18644 1106 18696 1158
rect 459 1026 511 1078
rect 523 1026 575 1078
rect 4398 1026 4450 1078
rect 4462 1026 4514 1078
rect 5217 1026 5269 1078
rect 5281 1026 5333 1078
rect 9229 1026 9281 1078
rect 9293 1026 9345 1078
rect 19713 1026 19765 1078
rect 19777 1026 19829 1078
rect 23725 1026 23777 1078
rect 23789 1026 23841 1078
rect 24545 1026 24597 1078
rect 24609 1026 24661 1078
rect 28557 1026 28609 1078
rect 28621 1026 28673 1078
rect 230 946 282 998
rect 294 946 346 998
rect 4554 946 4606 998
rect 4618 946 4670 998
rect 9892 946 9944 998
rect 9956 946 10008 998
rect 14142 946 14194 998
rect 14206 946 14258 998
rect 19556 946 19608 998
rect 19620 946 19672 998
rect 23882 946 23934 998
rect 23946 946 23998 998
rect 29220 946 29272 998
rect 29284 946 29336 998
rect 33546 946 33598 998
rect 33610 946 33662 998
rect 74 866 126 918
rect 138 866 190 918
rect 4904 866 4956 918
rect 4968 866 5020 918
rect 9736 866 9788 918
rect 9800 866 9852 918
rect 14568 866 14620 918
rect 14632 866 14684 918
rect 19400 866 19452 918
rect 19464 866 19516 918
rect 24232 866 24284 918
rect 24296 866 24348 918
rect 29064 866 29116 918
rect 29128 866 29180 918
rect 33896 866 33948 918
rect 33960 866 34012 918
rect 1121 786 1173 838
rect 1189 786 1241 838
rect 1257 786 1309 838
rect 1121 690 1173 742
rect 1189 690 1241 742
rect 1257 690 1309 742
rect 5953 786 6005 838
rect 6021 786 6073 838
rect 6089 786 6141 838
rect 5953 690 6005 742
rect 6021 690 6073 742
rect 6089 690 6141 742
rect 8677 786 8729 838
rect 8745 786 8797 838
rect 8813 786 8865 838
rect 8677 690 8729 742
rect 8745 690 8797 742
rect 8813 690 8865 742
rect 10785 786 10837 838
rect 10853 786 10905 838
rect 10921 786 10973 838
rect 10785 690 10837 742
rect 10853 690 10905 742
rect 10921 690 10973 742
rect 13509 786 13561 838
rect 13577 786 13629 838
rect 13645 786 13697 838
rect 13509 690 13561 742
rect 13577 690 13629 742
rect 13645 690 13697 742
rect 15617 786 15669 838
rect 15685 786 15737 838
rect 15753 786 15805 838
rect 15617 690 15669 742
rect 15685 690 15737 742
rect 15753 690 15805 742
rect 18341 786 18393 838
rect 18409 786 18461 838
rect 18477 786 18529 838
rect 18341 690 18393 742
rect 18409 690 18461 742
rect 18477 690 18529 742
rect 20449 786 20501 838
rect 20517 786 20569 838
rect 20585 786 20637 838
rect 20449 690 20501 742
rect 20517 690 20569 742
rect 20585 690 20637 742
rect 23173 786 23225 838
rect 23241 786 23293 838
rect 23309 786 23361 838
rect 23173 690 23225 742
rect 23241 690 23293 742
rect 23309 690 23361 742
rect 25281 786 25333 838
rect 25349 786 25401 838
rect 25417 786 25469 838
rect 25281 690 25333 742
rect 25349 690 25401 742
rect 25417 690 25469 742
rect 28005 786 28057 838
rect 28073 786 28125 838
rect 28141 786 28193 838
rect 28005 690 28057 742
rect 28073 690 28125 742
rect 28141 690 28193 742
rect 30113 786 30165 838
rect 30181 786 30233 838
rect 30249 786 30301 838
rect 30113 690 30165 742
rect 30181 690 30233 742
rect 30249 690 30301 742
rect 32837 786 32889 838
rect 32905 786 32957 838
rect 32973 786 33025 838
rect 32837 690 32889 742
rect 32905 690 32957 742
rect 32973 690 33025 742
rect 34945 786 34997 838
rect 35013 786 35065 838
rect 35081 786 35133 838
rect 34945 690 34997 742
rect 35013 690 35065 742
rect 35081 690 35133 742
rect 37669 786 37721 838
rect 37737 786 37789 838
rect 37805 786 37857 838
rect 37669 690 37721 742
rect 37737 690 37789 742
rect 37805 690 37857 742
rect 144 411 196 463
rect 144 345 196 397
rect 300 411 352 463
rect 300 345 352 397
rect 453 411 505 463
rect 453 345 505 397
rect 609 405 661 457
rect 609 339 661 391
rect 765 408 817 460
rect 765 344 817 396
rect 4078 413 4130 465
rect 4078 347 4130 399
rect 4236 405 4288 457
rect 4236 339 4288 391
rect 4392 411 4444 463
rect 4392 345 4444 397
rect 4548 411 4600 463
rect 4548 345 4600 397
rect 4704 411 4756 463
rect 4704 345 4756 397
rect 4974 411 5026 463
rect 4974 345 5026 397
rect 5130 411 5182 463
rect 5130 345 5182 397
rect 5287 411 5339 463
rect 5287 345 5339 397
rect 5444 405 5496 457
rect 5444 339 5496 391
rect 5600 413 5652 465
rect 5600 347 5652 399
rect 8910 413 8962 465
rect 8910 347 8962 399
rect 9066 405 9118 457
rect 9066 339 9118 391
rect 9223 411 9275 463
rect 9223 345 9275 397
rect 9380 411 9432 463
rect 9380 345 9432 397
rect 9536 411 9588 463
rect 9536 345 9588 397
rect 9806 411 9858 463
rect 9806 345 9858 397
rect 9962 411 10014 463
rect 9962 345 10014 397
rect 10119 411 10171 463
rect 10119 345 10171 397
rect 10275 409 10327 461
rect 10275 339 10327 391
rect 10432 413 10484 465
rect 10432 347 10484 399
rect 13742 413 13794 465
rect 13742 347 13794 399
rect 13898 409 13950 461
rect 13898 339 13950 391
rect 14055 411 14107 463
rect 14055 345 14107 397
rect 14212 411 14264 463
rect 14212 345 14264 397
rect 14368 411 14420 463
rect 14368 345 14420 397
rect 14638 411 14690 463
rect 14638 345 14690 397
rect 14794 411 14846 463
rect 14794 345 14846 397
rect 14951 411 15003 463
rect 14951 345 15003 397
rect 15107 409 15159 461
rect 15107 339 15159 391
rect 15264 413 15316 465
rect 15264 347 15316 399
rect 18574 413 18626 465
rect 18574 347 18626 399
rect 18731 409 18783 461
rect 18731 339 18783 391
rect 18887 411 18939 463
rect 18887 345 18939 397
rect 19044 411 19096 463
rect 19044 345 19096 397
rect 19200 411 19252 463
rect 19200 345 19252 397
rect 19470 411 19522 463
rect 19470 345 19522 397
rect 19626 411 19678 463
rect 19626 345 19678 397
rect 19783 411 19835 463
rect 19783 345 19835 397
rect 19939 409 19991 461
rect 19939 339 19991 391
rect 20093 409 20145 461
rect 20093 345 20145 397
rect 23409 409 23461 461
rect 23409 345 23461 397
rect 23563 409 23615 461
rect 23563 339 23615 391
rect 23719 411 23771 463
rect 23719 345 23771 397
rect 23876 411 23928 463
rect 23876 345 23928 397
rect 24032 411 24084 463
rect 24032 345 24084 397
rect 24302 411 24354 463
rect 24302 345 24354 397
rect 24458 411 24510 463
rect 24458 345 24510 397
rect 24615 411 24667 463
rect 24615 345 24667 397
rect 24771 409 24823 461
rect 24771 339 24823 391
rect 24925 409 24977 461
rect 24925 345 24977 397
rect 28241 413 28293 465
rect 28241 345 28293 397
rect 28395 409 28447 461
rect 28395 339 28447 391
rect 28551 411 28603 463
rect 28551 345 28603 397
rect 28708 411 28760 463
rect 28708 345 28760 397
rect 28864 411 28916 463
rect 28864 345 28916 397
rect 29134 411 29186 463
rect 29134 345 29186 397
rect 29290 411 29342 463
rect 29290 345 29342 397
rect 29447 411 29499 463
rect 29447 345 29499 397
rect 29601 409 29653 461
rect 29601 339 29653 391
rect 29757 413 29809 465
rect 29757 345 29809 397
rect 33073 413 33125 465
rect 33073 345 33125 397
rect 33227 409 33279 461
rect 33227 339 33279 391
rect 33383 411 33435 463
rect 33383 345 33435 397
rect 33540 411 33592 463
rect 33540 345 33592 397
rect 33696 411 33748 463
rect 33696 345 33748 397
rect 33966 411 34018 463
rect 33966 345 34018 397
rect 34122 411 34174 463
rect 34122 345 34174 397
rect 34279 411 34331 463
rect 34279 345 34331 397
rect 34433 409 34485 461
rect 34433 339 34485 391
rect 34589 413 34641 465
rect 34589 345 34641 397
rect 37905 413 37957 465
rect 37905 345 37957 397
rect 38059 409 38111 461
rect 38059 339 38111 391
rect 38215 411 38267 463
rect 38215 345 38267 397
rect 38372 411 38424 463
rect 38372 345 38424 397
rect 38528 411 38580 463
rect 38528 345 38580 397
rect 865 112 917 164
rect 933 112 985 164
rect 1001 112 1053 164
rect 865 0 917 52
rect 933 0 985 52
rect 1001 0 1053 52
rect 5697 112 5749 164
rect 5765 112 5817 164
rect 5833 112 5885 164
rect 5697 0 5749 52
rect 5765 0 5817 52
rect 5833 0 5885 52
rect 8421 112 8473 164
rect 8489 112 8541 164
rect 8557 112 8609 164
rect 8421 0 8473 52
rect 8489 0 8541 52
rect 8557 0 8609 52
rect 10529 112 10581 164
rect 10597 112 10649 164
rect 10665 112 10717 164
rect 10529 0 10581 52
rect 10597 0 10649 52
rect 10665 0 10717 52
rect 13253 112 13305 164
rect 13321 112 13373 164
rect 13389 112 13441 164
rect 13253 0 13305 52
rect 13321 0 13373 52
rect 13389 0 13441 52
rect 15361 112 15413 164
rect 15429 112 15481 164
rect 15497 112 15549 164
rect 15361 0 15413 52
rect 15429 0 15481 52
rect 15497 0 15549 52
rect 18085 112 18137 164
rect 18153 112 18205 164
rect 18221 112 18273 164
rect 18085 0 18137 52
rect 18153 0 18205 52
rect 18221 0 18273 52
rect 20193 112 20245 164
rect 20261 112 20313 164
rect 20329 112 20381 164
rect 20193 0 20245 52
rect 20261 0 20313 52
rect 20329 0 20381 52
rect 22917 112 22969 164
rect 22985 112 23037 164
rect 23053 112 23105 164
rect 22917 0 22969 52
rect 22985 0 23037 52
rect 23053 0 23105 52
rect 25025 112 25077 164
rect 25093 112 25145 164
rect 25161 112 25213 164
rect 25025 0 25077 52
rect 25093 0 25145 52
rect 25161 0 25213 52
rect 27749 112 27801 164
rect 27817 112 27869 164
rect 27885 112 27937 164
rect 27749 0 27801 52
rect 27817 0 27869 52
rect 27885 0 27937 52
rect 29857 112 29909 164
rect 29925 112 29977 164
rect 29993 112 30045 164
rect 29857 0 29909 52
rect 29925 0 29977 52
rect 29993 0 30045 52
rect 32581 112 32633 164
rect 32649 112 32701 164
rect 32717 112 32769 164
rect 32581 0 32633 52
rect 32649 0 32701 52
rect 32717 0 32769 52
rect 34689 112 34741 164
rect 34757 112 34809 164
rect 34825 112 34877 164
rect 34689 0 34741 52
rect 34757 0 34809 52
rect 34825 0 34877 52
rect 37413 112 37465 164
rect 37481 112 37533 164
rect 37549 112 37601 164
rect 37413 0 37465 52
rect 37481 0 37533 52
rect 37549 0 37601 52
rect 2249 -80 2301 -28
rect 2313 -80 2365 -28
rect 2533 -80 2585 -28
rect 2597 -80 2649 -28
rect 7081 -80 7133 -28
rect 7145 -80 7197 -28
rect 7365 -80 7417 -28
rect 7429 -80 7481 -28
rect 11913 -80 11965 -28
rect 11977 -80 12029 -28
rect 12197 -80 12249 -28
rect 12261 -80 12313 -28
rect 16745 -80 16797 -28
rect 16809 -80 16861 -28
rect 17029 -80 17081 -28
rect 17093 -80 17145 -28
rect 21577 -80 21629 -28
rect 21641 -80 21693 -28
rect 21861 -80 21913 -28
rect 21925 -80 21977 -28
rect 26409 -80 26461 -28
rect 26473 -80 26525 -28
rect 26693 -80 26745 -28
rect 26757 -80 26809 -28
rect 31241 -80 31293 -28
rect 31305 -80 31357 -28
rect 31525 -80 31577 -28
rect 31589 -80 31641 -28
rect 36073 -80 36125 -28
rect 36137 -80 36189 -28
rect 36357 -80 36409 -28
rect 36421 -80 36473 -28
<< metal2 >>
rect 2243 2588 2249 2640
rect 2301 2588 2313 2640
rect 2365 2588 2371 2640
rect 859 2452 865 2504
rect 917 2452 933 2504
rect 985 2452 1001 2504
rect 1053 2452 1059 2504
rect 859 2392 1059 2452
rect 859 2340 865 2392
rect 917 2340 933 2392
rect 985 2340 1001 2392
rect 1053 2340 1059 2392
rect 144 2159 196 2165
rect 144 2093 196 2107
tri 138 946 144 952 se
rect 144 946 196 2041
rect 300 2159 352 2165
rect 300 2093 352 2107
tri 294 1026 300 1032 se
rect 300 1026 352 2041
tri 266 998 294 1026 se
rect 294 998 352 1026
rect 224 946 230 998
rect 282 946 294 998
rect 346 946 352 998
tri 110 918 138 946 se
rect 138 918 196 946
tri 266 918 294 946 ne
rect 294 918 352 946
rect 68 866 74 918
rect 126 866 138 918
rect 190 866 196 918
tri 294 912 300 918 ne
tri 110 838 138 866 ne
rect 138 838 196 866
tri 138 832 144 838 ne
rect 144 463 196 838
rect 144 397 196 411
rect 144 339 196 345
rect 300 463 352 918
rect 300 397 352 411
rect 300 339 352 345
rect 453 2159 505 2165
rect 453 2093 505 2107
rect 453 1106 505 2041
rect 608 2160 660 2166
rect 608 2096 660 2108
rect 608 1666 660 2044
rect 765 2159 817 2165
rect 765 2095 817 2107
tri 660 1666 666 1672 sw
rect 608 1638 666 1666
tri 666 1638 694 1666 sw
rect 608 1586 614 1638
rect 666 1586 678 1638
rect 730 1586 736 1638
rect 533 1186 539 1238
rect 591 1186 603 1238
rect 655 1186 661 1238
tri 759 1186 765 1192 se
rect 765 1186 817 2043
tri 575 1158 603 1186 ne
rect 603 1158 661 1186
tri 731 1158 759 1186 se
rect 759 1158 817 1186
tri 603 1152 609 1158 ne
tri 505 1106 511 1112 sw
rect 453 1078 511 1106
tri 511 1078 539 1106 sw
rect 453 1026 459 1078
rect 511 1026 523 1078
rect 575 1026 581 1078
rect 453 998 511 1026
tri 511 998 539 1026 nw
rect 453 463 505 998
tri 505 992 511 998 nw
rect 453 397 505 411
rect 453 339 505 345
rect 609 457 661 1158
rect 689 1106 695 1158
rect 747 1106 759 1158
rect 811 1106 817 1158
tri 731 1078 759 1106 ne
rect 759 1078 817 1106
tri 759 1072 765 1078 ne
rect 609 391 661 405
rect 609 333 661 339
rect 765 460 817 1078
rect 765 396 817 408
rect 765 338 817 344
rect 859 164 1059 2340
rect 859 112 865 164
rect 917 112 933 164
rect 985 112 1001 164
rect 1053 112 1059 164
rect 859 52 1059 112
rect 859 0 865 52
rect 917 0 933 52
rect 985 0 1001 52
rect 1053 0 1059 52
rect 1115 1814 1315 2504
rect 2243 2370 2371 2588
rect 2527 2588 2533 2640
rect 2585 2588 2597 2640
rect 2649 2588 2655 2640
rect 2527 2370 2655 2588
rect 7075 2588 7081 2640
rect 7133 2588 7145 2640
rect 7197 2588 7203 2640
rect 5691 2452 5697 2504
rect 5749 2452 5765 2504
rect 5817 2452 5833 2504
rect 5885 2452 5891 2504
rect 5691 2392 5891 2452
rect 5691 2340 5697 2392
rect 5749 2340 5765 2392
rect 5817 2340 5833 2392
rect 5885 2340 5891 2392
rect 1115 1762 1121 1814
rect 1173 1762 1189 1814
rect 1241 1762 1257 1814
rect 1309 1762 1315 1814
rect 1115 1718 1315 1762
rect 1115 1666 1121 1718
rect 1173 1666 1189 1718
rect 1241 1666 1257 1718
rect 1309 1666 1315 1718
rect 1115 838 1315 1666
rect 1115 786 1121 838
rect 1173 786 1189 838
rect 1241 786 1257 838
rect 1309 786 1315 838
rect 1115 742 1315 786
rect 1115 690 1121 742
rect 1173 690 1189 742
rect 1241 690 1257 742
rect 1309 690 1315 742
rect 1115 0 1315 690
rect 4078 2155 4130 2161
rect 4078 2091 4130 2103
rect 4078 1186 4130 2039
rect 4235 2160 4287 2166
rect 4235 2096 4287 2108
rect 4235 1666 4287 2044
rect 4392 2159 4444 2165
rect 4392 2093 4444 2107
tri 4287 1666 4293 1672 sw
rect 4235 1638 4293 1666
tri 4293 1638 4321 1666 sw
rect 4235 1586 4241 1638
rect 4293 1586 4305 1638
rect 4357 1586 4363 1638
tri 4130 1186 4136 1192 sw
rect 4236 1186 4242 1238
rect 4294 1186 4306 1238
rect 4358 1186 4364 1238
rect 4078 1158 4136 1186
tri 4136 1158 4164 1186 sw
rect 4236 1158 4294 1186
tri 4294 1158 4322 1186 nw
rect 4078 1106 4084 1158
rect 4136 1106 4148 1158
rect 4200 1106 4206 1158
rect 4078 1078 4136 1106
tri 4136 1078 4164 1106 nw
rect 4078 465 4130 1078
tri 4130 1072 4136 1078 nw
rect 4078 399 4130 413
rect 4078 341 4130 347
rect 4236 457 4288 1158
tri 4288 1152 4294 1158 nw
rect 4236 391 4288 405
rect 4392 1106 4444 2041
rect 4548 2159 4600 2165
rect 4548 2093 4600 2107
tri 4444 1106 4450 1112 sw
rect 4392 1078 4450 1106
tri 4450 1078 4478 1106 sw
rect 4392 1026 4398 1078
rect 4450 1026 4462 1078
rect 4514 1026 4520 1078
rect 4548 1026 4600 2041
rect 4704 2159 4756 2165
rect 4704 2095 4756 2107
rect 4704 1346 4756 2043
rect 4974 2159 5026 2165
rect 4974 2093 5026 2107
tri 4756 1346 4762 1352 sw
rect 4704 1318 4762 1346
tri 4762 1318 4790 1346 sw
rect 4704 1266 4710 1318
rect 4762 1266 4774 1318
rect 4826 1266 4832 1318
rect 4704 1238 4762 1266
tri 4762 1238 4790 1266 nw
tri 4600 1026 4606 1032 sw
rect 4392 998 4450 1026
tri 4450 998 4478 1026 nw
rect 4548 998 4606 1026
tri 4606 998 4634 1026 sw
rect 4392 463 4444 998
tri 4444 992 4450 998 nw
rect 4392 397 4444 411
rect 4392 339 4444 345
rect 4548 946 4554 998
rect 4606 946 4618 998
rect 4670 946 4676 998
rect 4548 918 4606 946
tri 4606 918 4634 946 nw
rect 4548 463 4600 918
tri 4600 912 4606 918 nw
rect 4548 397 4600 411
rect 4548 339 4600 345
rect 4704 463 4756 1238
tri 4756 1232 4762 1238 nw
tri 4968 946 4974 952 se
rect 4974 946 5026 2041
rect 5130 2159 5182 2165
rect 5130 2093 5182 2107
tri 5124 1426 5130 1432 se
rect 5130 1426 5182 2041
tri 5096 1398 5124 1426 se
rect 5124 1398 5182 1426
rect 5054 1346 5060 1398
rect 5112 1346 5124 1398
rect 5176 1346 5182 1398
tri 5096 1318 5124 1346 ne
rect 5124 1318 5182 1346
tri 5124 1312 5130 1318 ne
tri 4940 918 4968 946 se
rect 4968 918 5026 946
rect 4898 866 4904 918
rect 4956 866 4968 918
rect 5020 866 5026 918
tri 4940 838 4968 866 ne
rect 4968 838 5026 866
tri 4968 832 4974 838 ne
rect 4704 397 4756 411
rect 4704 339 4756 345
rect 4974 463 5026 838
rect 4974 397 5026 411
rect 4974 339 5026 345
rect 5130 463 5182 1318
rect 5287 2159 5339 2165
rect 5287 2093 5339 2107
tri 5281 1106 5287 1112 se
rect 5287 1106 5339 2041
rect 5440 2160 5492 2166
rect 5440 2096 5492 2108
rect 5440 1666 5492 2044
rect 5600 2157 5652 2163
rect 5600 2091 5652 2105
tri 5492 1666 5498 1672 sw
rect 5440 1638 5498 1666
tri 5498 1638 5526 1666 sw
rect 5440 1586 5446 1638
rect 5498 1586 5510 1638
rect 5562 1586 5568 1638
rect 5368 1186 5374 1238
rect 5426 1186 5438 1238
rect 5490 1186 5496 1238
tri 5594 1186 5600 1192 se
rect 5600 1186 5652 2039
tri 5410 1158 5438 1186 ne
rect 5438 1158 5496 1186
tri 5566 1158 5594 1186 se
rect 5594 1158 5652 1186
tri 5438 1152 5444 1158 ne
tri 5253 1078 5281 1106 se
rect 5281 1078 5339 1106
rect 5211 1026 5217 1078
rect 5269 1026 5281 1078
rect 5333 1026 5339 1078
tri 5253 998 5281 1026 ne
rect 5281 998 5339 1026
tri 5281 992 5287 998 ne
rect 5130 397 5182 411
rect 5130 339 5182 345
rect 5287 463 5339 998
rect 5287 397 5339 411
rect 5287 339 5339 345
rect 5444 457 5496 1158
rect 5524 1106 5530 1158
rect 5582 1106 5594 1158
rect 5646 1106 5652 1158
tri 5566 1078 5594 1106 ne
rect 5594 1078 5652 1106
tri 5594 1072 5600 1078 ne
rect 5444 391 5496 405
rect 5600 465 5652 1078
rect 5600 399 5652 413
rect 5600 341 5652 347
rect 4236 333 4288 339
rect 5444 333 5496 339
rect 2243 -28 2371 176
rect 2243 -80 2249 -28
rect 2301 -80 2313 -28
rect 2365 -80 2371 -28
rect 2527 -28 2655 176
rect 5691 164 5891 2340
rect 5691 112 5697 164
rect 5749 112 5765 164
rect 5817 112 5833 164
rect 5885 112 5891 164
rect 5691 52 5891 112
rect 5691 0 5697 52
rect 5749 0 5765 52
rect 5817 0 5833 52
rect 5885 0 5891 52
rect 5947 1814 6147 2504
rect 7075 2370 7203 2588
rect 7359 2588 7365 2640
rect 7417 2588 7429 2640
rect 7481 2588 7487 2640
rect 7359 2370 7487 2588
rect 11907 2588 11913 2640
rect 11965 2588 11977 2640
rect 12029 2588 12035 2640
rect 8415 2452 8421 2504
rect 8473 2452 8489 2504
rect 8541 2452 8557 2504
rect 8609 2452 8615 2504
rect 8415 2392 8615 2452
rect 5947 1762 5953 1814
rect 6005 1762 6021 1814
rect 6073 1762 6089 1814
rect 6141 1762 6147 1814
rect 5947 1718 6147 1762
rect 5947 1666 5953 1718
rect 6005 1666 6021 1718
rect 6073 1666 6089 1718
rect 6141 1666 6147 1718
rect 5947 838 6147 1666
rect 5947 786 5953 838
rect 6005 786 6021 838
rect 6073 786 6089 838
rect 6141 786 6147 838
rect 5947 742 6147 786
rect 5947 690 5953 742
rect 6005 690 6021 742
rect 6073 690 6089 742
rect 6141 690 6147 742
rect 5947 0 6147 690
rect 8415 2340 8421 2392
rect 8473 2340 8489 2392
rect 8541 2340 8557 2392
rect 8609 2340 8615 2392
rect 2527 -80 2533 -28
rect 2585 -80 2597 -28
rect 2649 -80 2655 -28
rect 7075 -28 7203 176
rect 7075 -80 7081 -28
rect 7133 -80 7145 -28
rect 7197 -80 7203 -28
rect 7359 -28 7487 176
rect 8415 164 8615 2340
rect 8415 112 8421 164
rect 8473 112 8489 164
rect 8541 112 8557 164
rect 8609 112 8615 164
rect 8415 52 8615 112
rect 8415 0 8421 52
rect 8473 0 8489 52
rect 8541 0 8557 52
rect 8609 0 8615 52
rect 8671 1814 8871 2504
rect 10523 2452 10529 2504
rect 10581 2452 10597 2504
rect 10649 2452 10665 2504
rect 10717 2452 10723 2504
rect 10523 2392 10723 2452
rect 10523 2340 10529 2392
rect 10581 2340 10597 2392
rect 10649 2340 10665 2392
rect 10717 2340 10723 2392
rect 9067 2165 9119 2171
rect 8671 1762 8677 1814
rect 8729 1762 8745 1814
rect 8797 1762 8813 1814
rect 8865 1762 8871 1814
rect 8671 1718 8871 1762
rect 8671 1666 8677 1718
rect 8729 1666 8745 1718
rect 8797 1666 8813 1718
rect 8865 1666 8871 1718
rect 8671 838 8871 1666
rect 8671 786 8677 838
rect 8729 786 8745 838
rect 8797 786 8813 838
rect 8865 786 8871 838
rect 8671 742 8871 786
rect 8671 690 8677 742
rect 8729 690 8745 742
rect 8797 690 8813 742
rect 8865 690 8871 742
rect 8671 0 8871 690
rect 8910 2157 8962 2163
rect 8910 2091 8962 2105
rect 8910 1186 8962 2039
rect 9067 2096 9119 2113
rect 9067 1666 9119 2044
rect 9223 2159 9275 2165
rect 9223 2093 9275 2107
tri 9119 1666 9125 1672 sw
rect 9067 1638 9125 1666
tri 9125 1638 9153 1666 sw
rect 9067 1586 9073 1638
rect 9125 1586 9137 1638
rect 9189 1586 9195 1638
tri 8962 1186 8968 1192 sw
rect 9066 1186 9072 1238
rect 9124 1186 9136 1238
rect 9188 1186 9194 1238
rect 8910 1158 8968 1186
tri 8968 1158 8996 1186 sw
rect 9066 1158 9124 1186
tri 9124 1158 9152 1186 nw
rect 8910 1106 8916 1158
rect 8968 1106 8980 1158
rect 9032 1106 9038 1158
rect 8910 1078 8968 1106
tri 8968 1078 8996 1106 nw
rect 8910 465 8962 1078
tri 8962 1072 8968 1078 nw
rect 8910 399 8962 413
rect 8910 341 8962 347
rect 9066 457 9118 1158
tri 9118 1152 9124 1158 nw
rect 9066 391 9118 405
rect 9223 1106 9275 2041
rect 9380 2159 9432 2165
rect 9380 2093 9432 2107
rect 9380 1426 9432 2041
rect 9536 2159 9588 2165
rect 9536 2093 9588 2107
tri 9432 1426 9438 1432 sw
rect 9380 1398 9438 1426
tri 9438 1398 9466 1426 sw
rect 9380 1346 9386 1398
rect 9438 1346 9450 1398
rect 9502 1346 9508 1398
rect 9536 1346 9588 2041
rect 9806 2159 9858 2165
rect 9806 2093 9858 2107
tri 9588 1346 9594 1352 sw
rect 9380 1318 9438 1346
tri 9438 1318 9466 1346 nw
rect 9536 1318 9594 1346
tri 9594 1318 9622 1346 sw
tri 9275 1106 9281 1112 sw
rect 9223 1078 9281 1106
tri 9281 1078 9309 1106 sw
rect 9223 1026 9229 1078
rect 9281 1026 9293 1078
rect 9345 1026 9351 1078
rect 9223 998 9281 1026
tri 9281 998 9309 1026 nw
rect 9223 463 9275 998
tri 9275 992 9281 998 nw
rect 9223 397 9275 411
rect 9223 339 9275 345
rect 9380 463 9432 1318
tri 9432 1312 9438 1318 nw
rect 9380 397 9432 411
rect 9380 339 9432 345
rect 9536 1266 9542 1318
rect 9594 1266 9606 1318
rect 9658 1266 9664 1318
rect 9536 1238 9594 1266
tri 9594 1238 9622 1266 nw
rect 9536 463 9588 1238
tri 9588 1232 9594 1238 nw
tri 9800 946 9806 952 se
rect 9806 946 9858 2041
rect 9962 2159 10014 2165
rect 9962 2093 10014 2107
tri 9956 1026 9962 1032 se
rect 9962 1026 10014 2041
rect 10119 2159 10171 2165
rect 10119 2093 10171 2107
tri 10113 1506 10119 1512 se
rect 10119 1506 10171 2041
rect 10272 2160 10324 2166
rect 10272 2096 10324 2108
rect 10272 1666 10324 2044
rect 10432 2157 10484 2163
rect 10432 2091 10484 2105
tri 10324 1666 10330 1672 sw
rect 10272 1638 10330 1666
tri 10330 1638 10358 1666 sw
rect 10272 1586 10278 1638
rect 10330 1586 10342 1638
rect 10394 1586 10400 1638
tri 10085 1478 10113 1506 se
rect 10113 1478 10171 1506
rect 10043 1426 10049 1478
rect 10101 1426 10113 1478
rect 10165 1426 10171 1478
tri 10085 1398 10113 1426 ne
rect 10113 1398 10171 1426
tri 10113 1392 10119 1398 ne
tri 9928 998 9956 1026 se
rect 9956 998 10014 1026
rect 9886 946 9892 998
rect 9944 946 9956 998
rect 10008 946 10014 998
tri 9772 918 9800 946 se
rect 9800 918 9858 946
tri 9928 918 9956 946 ne
rect 9956 918 10014 946
rect 9730 866 9736 918
rect 9788 866 9800 918
rect 9852 866 9858 918
tri 9956 912 9962 918 ne
tri 9772 838 9800 866 ne
rect 9800 838 9858 866
tri 9800 832 9806 838 ne
rect 9536 397 9588 411
rect 9536 339 9588 345
rect 9806 463 9858 838
rect 9806 397 9858 411
rect 9806 339 9858 345
rect 9962 463 10014 918
rect 9962 397 10014 411
rect 9962 339 10014 345
rect 10119 463 10171 1398
rect 10199 1186 10205 1238
rect 10257 1186 10269 1238
rect 10321 1186 10327 1238
tri 10426 1186 10432 1192 se
rect 10432 1186 10484 2039
tri 10241 1158 10269 1186 ne
rect 10269 1158 10327 1186
tri 10398 1158 10426 1186 se
rect 10426 1158 10484 1186
tri 10269 1152 10275 1158 ne
rect 10119 397 10171 411
rect 10119 339 10171 345
rect 10275 461 10327 1158
rect 10356 1106 10362 1158
rect 10414 1106 10426 1158
rect 10478 1106 10484 1158
tri 10398 1078 10426 1106 ne
rect 10426 1078 10484 1106
tri 10426 1072 10432 1078 ne
rect 10275 391 10327 409
rect 10432 465 10484 1078
rect 10432 399 10484 413
rect 10432 341 10484 347
rect 9066 333 9118 339
rect 10275 333 10327 339
rect 10523 164 10723 2340
rect 10523 112 10529 164
rect 10581 112 10597 164
rect 10649 112 10665 164
rect 10717 112 10723 164
rect 10523 52 10723 112
rect 10523 0 10529 52
rect 10581 0 10597 52
rect 10649 0 10665 52
rect 10717 0 10723 52
rect 10779 1814 10979 2504
rect 11907 2370 12035 2588
rect 12191 2588 12197 2640
rect 12249 2588 12261 2640
rect 12313 2588 12319 2640
rect 12191 2370 12319 2588
rect 16739 2588 16745 2640
rect 16797 2588 16809 2640
rect 16861 2588 16867 2640
rect 13247 2452 13253 2504
rect 13305 2452 13321 2504
rect 13373 2452 13389 2504
rect 13441 2452 13447 2504
rect 13247 2392 13447 2452
rect 10779 1762 10785 1814
rect 10837 1762 10853 1814
rect 10905 1762 10921 1814
rect 10973 1762 10979 1814
rect 10779 1718 10979 1762
rect 10779 1666 10785 1718
rect 10837 1666 10853 1718
rect 10905 1666 10921 1718
rect 10973 1666 10979 1718
rect 10779 838 10979 1666
rect 10779 786 10785 838
rect 10837 786 10853 838
rect 10905 786 10921 838
rect 10973 786 10979 838
rect 10779 742 10979 786
rect 10779 690 10785 742
rect 10837 690 10853 742
rect 10905 690 10921 742
rect 10973 690 10979 742
rect 10779 0 10979 690
rect 13247 2340 13253 2392
rect 13305 2340 13321 2392
rect 13373 2340 13389 2392
rect 13441 2340 13447 2392
rect 7359 -80 7365 -28
rect 7417 -80 7429 -28
rect 7481 -80 7487 -28
rect 11907 -28 12035 176
rect 11907 -80 11913 -28
rect 11965 -80 11977 -28
rect 12029 -80 12035 -28
rect 12191 -28 12319 176
rect 13247 164 13447 2340
rect 13247 112 13253 164
rect 13305 112 13321 164
rect 13373 112 13389 164
rect 13441 112 13447 164
rect 13247 52 13447 112
rect 13247 0 13253 52
rect 13305 0 13321 52
rect 13373 0 13389 52
rect 13441 0 13447 52
rect 13503 1814 13703 2504
rect 15355 2452 15361 2504
rect 15413 2452 15429 2504
rect 15481 2452 15497 2504
rect 15549 2452 15555 2504
rect 15355 2392 15555 2452
rect 15355 2340 15361 2392
rect 15413 2340 15429 2392
rect 15481 2340 15497 2392
rect 15549 2340 15555 2392
rect 13899 2165 13951 2171
rect 13503 1762 13509 1814
rect 13561 1762 13577 1814
rect 13629 1762 13645 1814
rect 13697 1762 13703 1814
rect 13503 1718 13703 1762
rect 13503 1666 13509 1718
rect 13561 1666 13577 1718
rect 13629 1666 13645 1718
rect 13697 1666 13703 1718
rect 13503 838 13703 1666
rect 13503 786 13509 838
rect 13561 786 13577 838
rect 13629 786 13645 838
rect 13697 786 13703 838
rect 13503 742 13703 786
rect 13503 690 13509 742
rect 13561 690 13577 742
rect 13629 690 13645 742
rect 13697 690 13703 742
rect 13503 0 13703 690
rect 13742 2157 13794 2163
rect 13742 2091 13794 2105
rect 13742 1186 13794 2039
rect 13899 2096 13951 2113
rect 13899 1666 13951 2044
rect 14055 2159 14107 2165
rect 14055 2093 14107 2107
tri 13951 1666 13957 1672 sw
rect 13899 1638 13957 1666
tri 13957 1638 13985 1666 sw
rect 13899 1586 13905 1638
rect 13957 1586 13969 1638
rect 14021 1586 14027 1638
tri 14049 1506 14055 1512 se
rect 14055 1506 14107 2041
tri 14021 1478 14049 1506 se
rect 14049 1478 14107 1506
rect 13979 1426 13985 1478
rect 14037 1426 14049 1478
rect 14101 1426 14107 1478
tri 14021 1398 14049 1426 ne
rect 14049 1398 14107 1426
tri 14049 1392 14055 1398 ne
tri 13794 1186 13800 1192 sw
rect 13898 1186 13904 1238
rect 13956 1186 13968 1238
rect 14020 1186 14026 1238
rect 13742 1158 13800 1186
tri 13800 1158 13828 1186 sw
rect 13898 1158 13956 1186
tri 13956 1158 13984 1186 nw
rect 13742 1106 13748 1158
rect 13800 1106 13812 1158
rect 13864 1106 13870 1158
rect 13742 1078 13800 1106
tri 13800 1078 13828 1106 nw
rect 13742 465 13794 1078
tri 13794 1072 13800 1078 nw
rect 13742 399 13794 413
rect 13742 341 13794 347
rect 13898 461 13950 1158
tri 13950 1152 13956 1158 nw
rect 13898 391 13950 409
rect 14055 463 14107 1398
rect 14212 2159 14264 2165
rect 14212 2093 14264 2107
tri 14206 1026 14212 1032 se
rect 14212 1026 14264 2041
rect 14368 2159 14420 2165
rect 14368 2093 14420 2107
tri 14362 1346 14368 1352 se
rect 14368 1346 14420 2041
tri 14334 1318 14362 1346 se
rect 14362 1318 14420 1346
rect 14292 1266 14298 1318
rect 14350 1266 14362 1318
rect 14414 1266 14420 1318
tri 14334 1238 14362 1266 ne
rect 14362 1238 14420 1266
tri 14362 1232 14368 1238 ne
tri 14178 998 14206 1026 se
rect 14206 998 14264 1026
rect 14136 946 14142 998
rect 14194 946 14206 998
rect 14258 946 14264 998
tri 14178 918 14206 946 ne
rect 14206 918 14264 946
tri 14206 912 14212 918 ne
rect 14055 397 14107 411
rect 14055 339 14107 345
rect 14212 463 14264 918
rect 14212 397 14264 411
rect 14212 339 14264 345
rect 14368 463 14420 1238
rect 14638 2159 14690 2165
rect 14638 2093 14690 2107
tri 14632 946 14638 952 se
rect 14638 946 14690 2041
rect 14794 2159 14846 2165
rect 14794 2093 14846 2107
tri 14788 1426 14794 1432 se
rect 14794 1426 14846 2041
rect 14951 2159 15003 2165
rect 14951 2093 15003 2107
tri 14945 1506 14951 1512 se
rect 14951 1506 15003 2041
rect 15104 2160 15156 2166
rect 15104 2096 15156 2108
rect 15104 1666 15156 2044
rect 15264 2157 15316 2163
rect 15264 2091 15316 2105
tri 15156 1666 15162 1672 sw
rect 15104 1638 15162 1666
tri 15162 1638 15190 1666 sw
rect 15104 1586 15110 1638
rect 15162 1586 15174 1638
rect 15226 1586 15232 1638
tri 14917 1478 14945 1506 se
rect 14945 1478 15003 1506
rect 14875 1426 14881 1478
rect 14933 1426 14945 1478
rect 14997 1426 15003 1478
tri 14760 1398 14788 1426 se
rect 14788 1398 14846 1426
tri 14917 1398 14945 1426 ne
rect 14945 1398 15003 1426
rect 14718 1346 14724 1398
rect 14776 1346 14788 1398
rect 14840 1346 14846 1398
tri 14945 1392 14951 1398 ne
tri 14760 1318 14788 1346 ne
rect 14788 1318 14846 1346
tri 14788 1312 14794 1318 ne
tri 14604 918 14632 946 se
rect 14632 918 14690 946
rect 14562 866 14568 918
rect 14620 866 14632 918
rect 14684 866 14690 918
tri 14604 838 14632 866 ne
rect 14632 838 14690 866
tri 14632 832 14638 838 ne
rect 14368 397 14420 411
rect 14368 339 14420 345
rect 14638 463 14690 838
rect 14638 397 14690 411
rect 14638 339 14690 345
rect 14794 463 14846 1318
rect 14794 397 14846 411
rect 14794 339 14846 345
rect 14951 463 15003 1398
rect 15031 1186 15037 1238
rect 15089 1186 15101 1238
rect 15153 1186 15159 1238
tri 15258 1186 15264 1192 se
rect 15264 1186 15316 2039
tri 15073 1158 15101 1186 ne
rect 15101 1158 15159 1186
tri 15230 1158 15258 1186 se
rect 15258 1158 15316 1186
tri 15101 1152 15107 1158 ne
rect 14951 397 15003 411
rect 14951 339 15003 345
rect 15107 461 15159 1158
rect 15188 1106 15194 1158
rect 15246 1106 15258 1158
rect 15310 1106 15316 1158
tri 15230 1078 15258 1106 ne
rect 15258 1078 15316 1106
tri 15258 1072 15264 1078 ne
rect 15107 391 15159 409
rect 15264 465 15316 1078
rect 15264 399 15316 413
rect 15264 341 15316 347
rect 13898 333 13950 339
rect 15107 333 15159 339
rect 15355 164 15555 2340
rect 15355 112 15361 164
rect 15413 112 15429 164
rect 15481 112 15497 164
rect 15549 112 15555 164
rect 15355 52 15555 112
rect 15355 0 15361 52
rect 15413 0 15429 52
rect 15481 0 15497 52
rect 15549 0 15555 52
rect 15611 1814 15811 2504
rect 16739 2370 16867 2588
rect 17023 2588 17029 2640
rect 17081 2588 17093 2640
rect 17145 2588 17151 2640
rect 17023 2370 17151 2588
rect 21571 2588 21577 2640
rect 21629 2588 21641 2640
rect 21693 2588 21699 2640
rect 18079 2504 18279 2505
rect 18079 2452 18085 2504
rect 18137 2452 18153 2504
rect 18205 2452 18221 2504
rect 18273 2452 18279 2504
rect 18079 2392 18279 2452
rect 15611 1762 15617 1814
rect 15669 1762 15685 1814
rect 15737 1762 15753 1814
rect 15805 1762 15811 1814
rect 15611 1718 15811 1762
rect 15611 1666 15617 1718
rect 15669 1666 15685 1718
rect 15737 1666 15753 1718
rect 15805 1666 15811 1718
rect 15611 838 15811 1666
rect 15611 786 15617 838
rect 15669 786 15685 838
rect 15737 786 15753 838
rect 15805 786 15811 838
rect 15611 742 15811 786
rect 15611 690 15617 742
rect 15669 690 15685 742
rect 15737 690 15753 742
rect 15805 690 15811 742
rect 15611 0 15811 690
rect 18079 2340 18085 2392
rect 18137 2340 18153 2392
rect 18205 2340 18221 2392
rect 18273 2340 18279 2392
rect 12191 -80 12197 -28
rect 12249 -80 12261 -28
rect 12313 -80 12319 -28
rect 16739 -28 16867 176
rect 16739 -80 16745 -28
rect 16797 -80 16809 -28
rect 16861 -80 16867 -28
rect 17023 -28 17151 176
rect 18079 164 18279 2340
rect 18079 112 18085 164
rect 18137 112 18153 164
rect 18205 112 18221 164
rect 18273 112 18279 164
rect 18079 52 18279 112
rect 18079 0 18085 52
rect 18137 0 18153 52
rect 18205 0 18221 52
rect 18273 0 18279 52
rect 18335 1814 18535 2505
rect 20187 2452 20193 2504
rect 20245 2452 20261 2504
rect 20313 2452 20329 2504
rect 20381 2452 20387 2504
rect 20187 2392 20387 2452
rect 20187 2340 20193 2392
rect 20245 2340 20261 2392
rect 20313 2340 20329 2392
rect 20381 2340 20387 2392
rect 18731 2165 18783 2171
rect 19939 2165 19991 2171
rect 18335 1762 18341 1814
rect 18393 1762 18409 1814
rect 18461 1762 18477 1814
rect 18529 1762 18535 1814
rect 18335 1718 18535 1762
rect 18335 1666 18341 1718
rect 18393 1666 18409 1718
rect 18461 1666 18477 1718
rect 18529 1666 18535 1718
rect 18335 838 18535 1666
rect 18335 786 18341 838
rect 18393 786 18409 838
rect 18461 786 18477 838
rect 18529 786 18535 838
rect 18335 742 18535 786
rect 18335 690 18341 742
rect 18393 690 18409 742
rect 18461 690 18477 742
rect 18529 690 18535 742
rect 18335 1 18535 690
rect 18574 2157 18626 2163
rect 18574 2091 18626 2105
rect 18574 1186 18626 2039
rect 18731 2096 18783 2113
rect 18731 1666 18783 2044
rect 18887 2159 18939 2165
rect 18887 2093 18939 2107
tri 18783 1666 18789 1672 sw
rect 18731 1638 18789 1666
tri 18789 1638 18817 1666 sw
rect 18731 1586 18737 1638
rect 18789 1586 18801 1638
rect 18853 1586 18859 1638
rect 18887 1506 18939 2041
rect 19044 2159 19096 2165
rect 19044 2093 19096 2107
tri 18939 1506 18945 1512 sw
rect 18887 1478 18945 1506
tri 18945 1478 18973 1506 sw
rect 18887 1426 18893 1478
rect 18945 1426 18957 1478
rect 19009 1426 19015 1478
rect 19044 1426 19096 2041
rect 19200 2159 19252 2165
rect 19200 2093 19252 2107
tri 19096 1426 19102 1432 sw
rect 18887 1398 18945 1426
tri 18945 1398 18973 1426 nw
rect 19044 1398 19102 1426
tri 19102 1398 19130 1426 sw
tri 18626 1186 18632 1192 sw
rect 18731 1186 18737 1238
rect 18789 1186 18801 1238
rect 18853 1186 18859 1238
rect 18574 1158 18632 1186
tri 18632 1158 18660 1186 sw
rect 18574 1106 18580 1158
rect 18632 1106 18644 1158
rect 18696 1106 18702 1158
rect 18574 1078 18632 1106
tri 18632 1078 18660 1106 nw
rect 18574 465 18626 1078
tri 18626 1072 18632 1078 nw
rect 18574 399 18626 413
rect 18574 341 18626 347
rect 18731 461 18783 1186
tri 18783 1152 18817 1186 nw
rect 18731 391 18783 409
rect 18887 463 18939 1398
tri 18939 1392 18945 1398 nw
rect 18887 397 18939 411
rect 18887 339 18939 345
rect 19044 1346 19050 1398
rect 19102 1346 19114 1398
rect 19166 1346 19172 1398
rect 19200 1346 19252 2041
rect 19470 2159 19522 2165
rect 19470 2093 19522 2107
tri 19252 1346 19258 1352 sw
rect 19044 1318 19102 1346
tri 19102 1318 19130 1346 nw
rect 19200 1318 19258 1346
tri 19258 1318 19286 1346 sw
rect 19044 463 19096 1318
tri 19096 1312 19102 1318 nw
rect 19044 397 19096 411
rect 19044 339 19096 345
rect 19200 1266 19206 1318
rect 19258 1266 19270 1318
rect 19322 1266 19328 1318
rect 19200 1238 19258 1266
tri 19258 1238 19286 1266 nw
rect 19200 463 19252 1238
tri 19252 1232 19258 1238 nw
tri 19464 946 19470 952 se
rect 19470 946 19522 2041
rect 19626 2159 19678 2165
rect 19626 2093 19678 2107
tri 19620 1026 19626 1032 se
rect 19626 1026 19678 2041
rect 19783 2159 19835 2165
rect 19783 2093 19835 2107
tri 19749 1078 19783 1112 se
rect 19783 1078 19835 2041
rect 19939 2096 19991 2113
tri 19933 1666 19939 1672 se
rect 19939 1666 19991 2044
tri 19905 1638 19933 1666 se
rect 19933 1638 19991 1666
rect 19863 1586 19869 1638
rect 19921 1586 19933 1638
rect 19985 1586 19991 1638
rect 20093 2159 20145 2165
rect 20093 2095 20145 2107
tri 20087 1586 20093 1592 se
rect 20093 1586 20145 2043
tri 20059 1558 20087 1586 se
rect 20087 1558 20145 1586
rect 20017 1506 20023 1558
rect 20075 1506 20087 1558
rect 20139 1506 20145 1558
tri 20059 1478 20087 1506 ne
rect 20087 1478 20145 1506
tri 20087 1472 20093 1478 ne
rect 19863 1186 19869 1238
rect 19921 1186 19933 1238
rect 19985 1186 19991 1238
tri 19905 1152 19939 1186 ne
rect 19707 1026 19713 1078
rect 19765 1026 19777 1078
rect 19829 1026 19835 1078
tri 19592 998 19620 1026 se
rect 19620 998 19678 1026
tri 19749 998 19777 1026 ne
rect 19777 998 19835 1026
rect 19550 946 19556 998
rect 19608 946 19620 998
rect 19672 946 19678 998
tri 19777 992 19783 998 ne
tri 19436 918 19464 946 se
rect 19464 918 19522 946
tri 19592 918 19620 946 ne
rect 19620 918 19678 946
rect 19394 866 19400 918
rect 19452 866 19464 918
rect 19516 866 19522 918
tri 19620 912 19626 918 ne
tri 19436 838 19464 866 ne
rect 19464 838 19522 866
tri 19464 832 19470 838 ne
rect 19200 397 19252 411
rect 19200 339 19252 345
rect 19470 463 19522 838
rect 19470 397 19522 411
rect 19470 339 19522 345
rect 19626 463 19678 918
rect 19626 397 19678 411
rect 19626 339 19678 345
rect 19783 463 19835 998
rect 19783 397 19835 411
rect 19783 339 19835 345
rect 19939 461 19991 1186
rect 19939 391 19991 409
rect 20093 461 20145 1478
rect 20093 397 20145 409
rect 20093 339 20145 345
rect 18731 333 18783 339
rect 19939 333 19991 339
rect 20187 164 20387 2340
rect 20187 112 20193 164
rect 20245 112 20261 164
rect 20313 112 20329 164
rect 20381 112 20387 164
rect 20187 52 20387 112
rect 20187 0 20193 52
rect 20245 0 20261 52
rect 20313 0 20329 52
rect 20381 0 20387 52
rect 20443 1814 20643 2504
rect 21571 2370 21699 2588
rect 21855 2588 21861 2640
rect 21913 2588 21925 2640
rect 21977 2588 21983 2640
rect 21855 2370 21983 2588
rect 26403 2588 26409 2640
rect 26461 2588 26473 2640
rect 26525 2588 26531 2640
rect 22911 2504 23111 2505
rect 22911 2452 22917 2504
rect 22969 2452 22985 2504
rect 23037 2452 23053 2504
rect 23105 2452 23111 2504
rect 22911 2392 23111 2452
rect 20443 1762 20449 1814
rect 20501 1762 20517 1814
rect 20569 1762 20585 1814
rect 20637 1762 20643 1814
rect 20443 1718 20643 1762
rect 20443 1666 20449 1718
rect 20501 1666 20517 1718
rect 20569 1666 20585 1718
rect 20637 1666 20643 1718
rect 20443 838 20643 1666
rect 20443 786 20449 838
rect 20501 786 20517 838
rect 20569 786 20585 838
rect 20637 786 20643 838
rect 20443 742 20643 786
rect 20443 690 20449 742
rect 20501 690 20517 742
rect 20569 690 20585 742
rect 20637 690 20643 742
rect 20443 0 20643 690
rect 22911 2340 22917 2392
rect 22969 2340 22985 2392
rect 23037 2340 23053 2392
rect 23105 2340 23111 2392
rect 17023 -80 17029 -28
rect 17081 -80 17093 -28
rect 17145 -80 17151 -28
rect 21571 -28 21699 176
rect 21571 -80 21577 -28
rect 21629 -80 21641 -28
rect 21693 -80 21699 -28
rect 21855 -28 21983 176
rect 22911 164 23111 2340
rect 22911 112 22917 164
rect 22969 112 22985 164
rect 23037 112 23053 164
rect 23105 112 23111 164
rect 22911 52 23111 112
rect 22911 0 22917 52
rect 22969 0 22985 52
rect 23037 0 23053 52
rect 23105 0 23111 52
rect 23167 1814 23367 2505
rect 25019 2452 25025 2504
rect 25077 2452 25093 2504
rect 25145 2452 25161 2504
rect 25213 2452 25219 2504
rect 25019 2392 25219 2452
rect 25019 2340 25025 2392
rect 25077 2340 25093 2392
rect 25145 2340 25161 2392
rect 25213 2340 25219 2392
rect 23167 1762 23173 1814
rect 23225 1762 23241 1814
rect 23293 1762 23309 1814
rect 23361 1762 23367 1814
rect 23167 1718 23367 1762
rect 23167 1666 23173 1718
rect 23225 1666 23241 1718
rect 23293 1666 23309 1718
rect 23361 1666 23367 1718
rect 23167 838 23367 1666
rect 23167 786 23173 838
rect 23225 786 23241 838
rect 23293 786 23309 838
rect 23361 786 23367 838
rect 23167 742 23367 786
rect 23167 690 23173 742
rect 23225 690 23241 742
rect 23293 690 23309 742
rect 23361 690 23367 742
rect 23167 1 23367 690
rect 23409 2159 23461 2165
rect 23409 2095 23461 2107
rect 23409 1586 23461 2043
rect 23560 2160 23612 2166
rect 24774 2165 24826 2171
rect 23560 2096 23612 2108
rect 23560 1666 23612 2044
rect 23719 2159 23771 2165
rect 23719 2093 23771 2107
tri 23612 1666 23618 1672 sw
rect 23560 1638 23618 1666
tri 23618 1638 23646 1666 sw
tri 23461 1586 23467 1592 sw
rect 23560 1586 23566 1638
rect 23618 1586 23630 1638
rect 23682 1586 23688 1638
rect 23409 1558 23467 1586
tri 23467 1558 23495 1586 sw
rect 23409 1506 23415 1558
rect 23467 1506 23479 1558
rect 23531 1506 23537 1558
rect 23409 1478 23467 1506
tri 23467 1478 23495 1506 nw
rect 23409 461 23461 1478
tri 23461 1472 23467 1478 nw
rect 23409 397 23461 409
rect 23409 339 23461 345
rect 23563 1186 23569 1238
rect 23621 1186 23633 1238
rect 23685 1186 23691 1238
rect 23563 461 23615 1186
tri 23615 1152 23649 1186 nw
rect 23563 391 23615 409
rect 23719 1078 23771 2041
rect 23876 2159 23928 2165
rect 23876 2093 23928 2107
tri 23771 1078 23805 1112 sw
rect 23719 1026 23725 1078
rect 23777 1026 23789 1078
rect 23841 1026 23847 1078
rect 23876 1026 23928 2041
rect 24032 2159 24084 2165
rect 24032 2093 24084 2107
rect 24032 1346 24084 2041
rect 24302 2159 24354 2165
rect 24302 2093 24354 2107
tri 24084 1346 24090 1352 sw
rect 24032 1318 24090 1346
tri 24090 1318 24118 1346 sw
rect 24032 1266 24038 1318
rect 24090 1266 24102 1318
rect 24154 1266 24160 1318
rect 24032 1238 24090 1266
tri 24090 1238 24118 1266 nw
tri 23928 1026 23934 1032 sw
rect 23719 998 23777 1026
tri 23777 998 23805 1026 nw
rect 23876 998 23934 1026
tri 23934 998 23962 1026 sw
rect 23719 463 23771 998
tri 23771 992 23777 998 nw
rect 23719 397 23771 411
rect 23719 339 23771 345
rect 23876 946 23882 998
rect 23934 946 23946 998
rect 23998 946 24004 998
rect 23876 918 23934 946
tri 23934 918 23962 946 nw
rect 23876 463 23928 918
tri 23928 912 23934 918 nw
rect 23876 397 23928 411
rect 23876 339 23928 345
rect 24032 463 24084 1238
tri 24084 1232 24090 1238 nw
tri 24296 946 24302 952 se
rect 24302 946 24354 2041
rect 24458 2159 24510 2165
rect 24458 2093 24510 2107
tri 24452 1426 24458 1432 se
rect 24458 1426 24510 2041
tri 24424 1398 24452 1426 se
rect 24452 1398 24510 1426
rect 24382 1346 24388 1398
rect 24440 1346 24452 1398
rect 24504 1346 24510 1398
tri 24424 1318 24452 1346 ne
rect 24452 1318 24510 1346
tri 24452 1312 24458 1318 ne
tri 24268 918 24296 946 se
rect 24296 918 24354 946
rect 24226 866 24232 918
rect 24284 866 24296 918
rect 24348 866 24354 918
tri 24268 838 24296 866 ne
rect 24296 838 24354 866
tri 24296 832 24302 838 ne
rect 24032 397 24084 411
rect 24032 339 24084 345
rect 24302 463 24354 838
rect 24302 397 24354 411
rect 24302 339 24354 345
rect 24458 463 24510 1318
rect 24615 2159 24667 2165
rect 24615 2093 24667 2107
tri 24581 1078 24615 1112 se
rect 24615 1078 24667 2041
rect 24774 2096 24826 2113
tri 24768 1666 24774 1672 se
rect 24774 1666 24826 2044
tri 24740 1638 24768 1666 se
rect 24768 1638 24826 1666
rect 24698 1586 24704 1638
rect 24756 1586 24768 1638
rect 24820 1586 24826 1638
rect 24925 2159 24977 2165
rect 24925 2095 24977 2107
tri 24919 1586 24925 1592 se
rect 24925 1586 24977 2043
tri 24891 1558 24919 1586 se
rect 24919 1558 24977 1586
rect 24849 1506 24855 1558
rect 24907 1506 24919 1558
rect 24971 1506 24977 1558
tri 24891 1478 24919 1506 ne
rect 24919 1478 24977 1506
tri 24919 1472 24925 1478 ne
rect 24695 1186 24701 1238
rect 24753 1186 24765 1238
rect 24817 1186 24823 1238
tri 24737 1152 24771 1186 ne
rect 24539 1026 24545 1078
rect 24597 1026 24609 1078
rect 24661 1026 24667 1078
tri 24581 998 24609 1026 ne
rect 24609 998 24667 1026
tri 24609 992 24615 998 ne
rect 24458 397 24510 411
rect 24458 339 24510 345
rect 24615 463 24667 998
rect 24615 397 24667 411
rect 24615 339 24667 345
rect 24771 461 24823 1186
rect 24771 391 24823 409
rect 24925 461 24977 1478
rect 24925 397 24977 409
rect 24925 339 24977 345
rect 23563 333 23615 339
rect 24771 333 24823 339
rect 25019 164 25219 2340
rect 25019 112 25025 164
rect 25077 112 25093 164
rect 25145 112 25161 164
rect 25213 112 25219 164
rect 25019 52 25219 112
rect 25019 0 25025 52
rect 25077 0 25093 52
rect 25145 0 25161 52
rect 25213 0 25219 52
rect 25275 1814 25475 2504
rect 26403 2370 26531 2588
rect 26687 2588 26693 2640
rect 26745 2588 26757 2640
rect 26809 2588 26815 2640
rect 26687 2370 26815 2588
rect 31235 2588 31241 2640
rect 31293 2588 31305 2640
rect 31357 2588 31363 2640
rect 27743 2504 27943 2505
rect 27743 2452 27749 2504
rect 27801 2452 27817 2504
rect 27869 2452 27885 2504
rect 27937 2452 27943 2504
rect 27743 2392 27943 2452
rect 25275 1762 25281 1814
rect 25333 1762 25349 1814
rect 25401 1762 25417 1814
rect 25469 1762 25475 1814
rect 25275 1718 25475 1762
rect 25275 1666 25281 1718
rect 25333 1666 25349 1718
rect 25401 1666 25417 1718
rect 25469 1666 25475 1718
rect 25275 838 25475 1666
rect 25275 786 25281 838
rect 25333 786 25349 838
rect 25401 786 25417 838
rect 25469 786 25475 838
rect 25275 742 25475 786
rect 25275 690 25281 742
rect 25333 690 25349 742
rect 25401 690 25417 742
rect 25469 690 25475 742
rect 25275 0 25475 690
rect 27743 2340 27749 2392
rect 27801 2340 27817 2392
rect 27869 2340 27885 2392
rect 27937 2340 27943 2392
rect 21855 -80 21861 -28
rect 21913 -80 21925 -28
rect 21977 -80 21983 -28
rect 26403 -28 26531 176
rect 26403 -80 26409 -28
rect 26461 -80 26473 -28
rect 26525 -80 26531 -28
rect 26687 -28 26815 176
rect 27743 164 27943 2340
rect 27743 112 27749 164
rect 27801 112 27817 164
rect 27869 112 27885 164
rect 27937 112 27943 164
rect 27743 52 27943 112
rect 27743 0 27749 52
rect 27801 0 27817 52
rect 27869 0 27885 52
rect 27937 0 27943 52
rect 27999 1814 28199 2505
rect 29851 2452 29857 2504
rect 29909 2452 29925 2504
rect 29977 2452 29993 2504
rect 30045 2452 30051 2504
rect 29851 2392 30051 2452
rect 29851 2340 29857 2392
rect 29909 2340 29925 2392
rect 29977 2340 29993 2392
rect 30045 2340 30051 2392
rect 28395 2165 28447 2171
rect 29606 2165 29658 2171
rect 27999 1762 28005 1814
rect 28057 1762 28073 1814
rect 28125 1762 28141 1814
rect 28193 1762 28199 1814
rect 27999 1718 28199 1762
rect 27999 1666 28005 1718
rect 28057 1666 28073 1718
rect 28125 1666 28141 1718
rect 28193 1666 28199 1718
rect 27999 838 28199 1666
rect 27999 786 28005 838
rect 28057 786 28073 838
rect 28125 786 28141 838
rect 28193 786 28199 838
rect 27999 742 28199 786
rect 27999 690 28005 742
rect 28057 690 28073 742
rect 28125 690 28141 742
rect 28193 690 28199 742
rect 27999 1 28199 690
rect 28241 2159 28293 2165
rect 28241 2091 28293 2107
rect 28241 1586 28293 2039
rect 28395 2096 28447 2113
rect 28395 1666 28447 2044
rect 28551 2159 28603 2165
rect 28551 2093 28603 2107
tri 28447 1666 28453 1672 sw
rect 28395 1638 28453 1666
tri 28453 1638 28481 1666 sw
tri 28293 1586 28299 1592 sw
rect 28395 1586 28401 1638
rect 28453 1586 28465 1638
rect 28517 1586 28523 1638
rect 28241 1558 28299 1586
tri 28299 1558 28327 1586 sw
rect 28241 1506 28247 1558
rect 28299 1506 28311 1558
rect 28363 1506 28369 1558
rect 28241 1478 28299 1506
tri 28299 1478 28327 1506 nw
rect 28241 465 28293 1478
tri 28293 1472 28299 1478 nw
rect 28241 397 28293 413
rect 28241 339 28293 345
rect 28395 1186 28401 1238
rect 28453 1186 28465 1238
rect 28517 1186 28523 1238
rect 28395 461 28447 1186
tri 28447 1152 28481 1186 nw
rect 28395 391 28447 409
rect 28551 1078 28603 2041
rect 28708 2159 28760 2165
rect 28708 2093 28760 2107
rect 28708 1426 28760 2041
rect 28864 2159 28916 2165
rect 28864 2093 28916 2107
tri 28760 1426 28766 1432 sw
rect 28708 1398 28766 1426
tri 28766 1398 28794 1426 sw
rect 28708 1346 28714 1398
rect 28766 1346 28778 1398
rect 28830 1346 28836 1398
rect 28864 1346 28916 2041
rect 29134 2159 29186 2165
rect 29134 2093 29186 2107
tri 28916 1346 28922 1352 sw
rect 28708 1318 28766 1346
tri 28766 1318 28794 1346 nw
rect 28864 1318 28922 1346
tri 28922 1318 28950 1346 sw
tri 28603 1078 28637 1112 sw
rect 28551 1026 28557 1078
rect 28609 1026 28621 1078
rect 28673 1026 28679 1078
rect 28551 998 28609 1026
tri 28609 998 28637 1026 nw
rect 28551 463 28603 998
tri 28603 992 28609 998 nw
rect 28551 397 28603 411
rect 28551 339 28603 345
rect 28708 463 28760 1318
tri 28760 1312 28766 1318 nw
rect 28708 397 28760 411
rect 28708 339 28760 345
rect 28864 1266 28870 1318
rect 28922 1266 28934 1318
rect 28986 1266 28992 1318
rect 28864 1238 28922 1266
tri 28922 1238 28950 1266 nw
rect 28864 463 28916 1238
tri 28916 1232 28922 1238 nw
tri 29128 946 29134 952 se
rect 29134 946 29186 2041
rect 29290 2159 29342 2165
rect 29290 2093 29342 2107
tri 29256 998 29290 1032 se
rect 29290 998 29342 2041
rect 29447 2159 29499 2165
rect 29447 2093 29499 2107
tri 29441 1506 29447 1512 se
rect 29447 1506 29499 2041
rect 29606 2096 29658 2113
tri 29600 1666 29606 1672 se
rect 29606 1666 29658 2044
tri 29572 1638 29600 1666 se
rect 29600 1638 29658 1666
rect 29530 1586 29536 1638
rect 29588 1586 29600 1638
rect 29652 1586 29658 1638
rect 29757 2159 29809 2165
rect 29757 2091 29809 2107
tri 29751 1586 29757 1592 se
rect 29757 1586 29809 2039
tri 29723 1558 29751 1586 se
rect 29751 1558 29809 1586
rect 29681 1506 29687 1558
rect 29739 1506 29751 1558
rect 29803 1506 29809 1558
tri 29413 1478 29441 1506 se
rect 29441 1478 29499 1506
tri 29723 1478 29751 1506 ne
rect 29751 1478 29809 1506
rect 29371 1426 29377 1478
rect 29429 1426 29441 1478
rect 29493 1426 29499 1478
tri 29751 1472 29757 1478 ne
tri 29413 1398 29441 1426 ne
rect 29441 1398 29499 1426
tri 29441 1392 29447 1398 ne
rect 29214 946 29220 998
rect 29272 946 29284 998
rect 29336 946 29342 998
tri 29100 918 29128 946 se
rect 29128 918 29186 946
tri 29256 918 29284 946 ne
rect 29284 918 29342 946
rect 29058 866 29064 918
rect 29116 866 29128 918
rect 29180 866 29186 918
tri 29284 912 29290 918 ne
tri 29100 838 29128 866 ne
rect 29128 838 29186 866
tri 29128 832 29134 838 ne
rect 28864 397 28916 411
rect 28864 339 28916 345
rect 29134 463 29186 838
rect 29134 397 29186 411
rect 29134 339 29186 345
rect 29290 463 29342 918
rect 29290 397 29342 411
rect 29290 339 29342 345
rect 29447 463 29499 1398
rect 29447 397 29499 411
rect 29447 339 29499 345
rect 29601 1186 29607 1238
rect 29659 1186 29671 1238
rect 29723 1186 29729 1238
rect 29601 461 29653 1186
tri 29653 1152 29687 1186 nw
rect 29601 391 29653 409
rect 29757 465 29809 1478
rect 29757 397 29809 413
rect 29757 339 29809 345
rect 28395 333 28447 339
rect 29601 333 29653 339
rect 29851 164 30051 2340
rect 29851 112 29857 164
rect 29909 112 29925 164
rect 29977 112 29993 164
rect 30045 112 30051 164
rect 29851 52 30051 112
rect 29851 0 29857 52
rect 29909 0 29925 52
rect 29977 0 29993 52
rect 30045 0 30051 52
rect 30107 1814 30307 2504
rect 31235 2370 31363 2588
rect 31519 2588 31525 2640
rect 31577 2588 31589 2640
rect 31641 2588 31647 2640
rect 31519 2370 31647 2588
rect 36067 2588 36073 2640
rect 36125 2588 36137 2640
rect 36189 2588 36195 2640
rect 32575 2504 32775 2505
rect 32575 2452 32581 2504
rect 32633 2452 32649 2504
rect 32701 2452 32717 2504
rect 32769 2452 32775 2504
rect 32575 2392 32775 2452
rect 30107 1762 30113 1814
rect 30165 1762 30181 1814
rect 30233 1762 30249 1814
rect 30301 1762 30307 1814
rect 30107 1718 30307 1762
rect 30107 1666 30113 1718
rect 30165 1666 30181 1718
rect 30233 1666 30249 1718
rect 30301 1666 30307 1718
rect 30107 838 30307 1666
rect 30107 786 30113 838
rect 30165 786 30181 838
rect 30233 786 30249 838
rect 30301 786 30307 838
rect 30107 742 30307 786
rect 30107 690 30113 742
rect 30165 690 30181 742
rect 30233 690 30249 742
rect 30301 690 30307 742
rect 30107 0 30307 690
rect 32575 2340 32581 2392
rect 32633 2340 32649 2392
rect 32701 2340 32717 2392
rect 32769 2340 32775 2392
rect 26687 -80 26693 -28
rect 26745 -80 26757 -28
rect 26809 -80 26815 -28
rect 31235 -28 31363 176
rect 31235 -80 31241 -28
rect 31293 -80 31305 -28
rect 31357 -80 31363 -28
rect 31519 -28 31647 176
rect 32575 164 32775 2340
rect 32575 112 32581 164
rect 32633 112 32649 164
rect 32701 112 32717 164
rect 32769 112 32775 164
rect 32575 52 32775 112
rect 32575 0 32581 52
rect 32633 0 32649 52
rect 32701 0 32717 52
rect 32769 0 32775 52
rect 32831 1814 33031 2505
rect 34683 2452 34689 2504
rect 34741 2452 34757 2504
rect 34809 2452 34825 2504
rect 34877 2452 34883 2504
rect 34683 2392 34883 2452
rect 34683 2340 34689 2392
rect 34741 2340 34757 2392
rect 34809 2340 34825 2392
rect 34877 2340 34883 2392
rect 33227 2165 33279 2171
rect 34435 2165 34487 2171
rect 32831 1762 32837 1814
rect 32889 1762 32905 1814
rect 32957 1762 32973 1814
rect 33025 1762 33031 1814
rect 32831 1718 33031 1762
rect 32831 1666 32837 1718
rect 32889 1666 32905 1718
rect 32957 1666 32973 1718
rect 33025 1666 33031 1718
rect 32831 838 33031 1666
rect 32831 786 32837 838
rect 32889 786 32905 838
rect 32957 786 32973 838
rect 33025 786 33031 838
rect 32831 742 33031 786
rect 32831 690 32837 742
rect 32889 690 32905 742
rect 32957 690 32973 742
rect 33025 690 33031 742
rect 32831 1 33031 690
rect 33073 2159 33125 2165
rect 33073 2091 33125 2107
rect 33073 1586 33125 2039
rect 33227 2096 33279 2113
rect 33227 1666 33279 2044
rect 33383 2159 33435 2165
rect 33383 2093 33435 2107
tri 33279 1666 33285 1672 sw
rect 33227 1638 33285 1666
tri 33285 1638 33313 1666 sw
tri 33125 1586 33131 1592 sw
rect 33227 1586 33233 1638
rect 33285 1586 33297 1638
rect 33349 1586 33355 1638
rect 33073 1558 33131 1586
tri 33131 1558 33159 1586 sw
rect 33073 1506 33079 1558
rect 33131 1506 33143 1558
rect 33195 1506 33201 1558
rect 33383 1506 33435 2041
rect 33540 2159 33592 2165
rect 33540 2093 33592 2107
tri 33435 1506 33441 1512 sw
rect 33073 1478 33131 1506
tri 33131 1478 33159 1506 nw
rect 33383 1478 33441 1506
tri 33441 1478 33469 1506 sw
rect 33073 465 33125 1478
tri 33125 1472 33131 1478 nw
rect 33383 1426 33389 1478
rect 33441 1426 33453 1478
rect 33505 1426 33511 1478
rect 33383 1398 33441 1426
tri 33441 1398 33469 1426 nw
rect 33073 397 33125 413
rect 33073 339 33125 345
rect 33227 1186 33233 1238
rect 33285 1186 33297 1238
rect 33349 1186 33355 1238
rect 33227 461 33279 1186
tri 33279 1152 33313 1186 nw
rect 33227 391 33279 409
rect 33383 463 33435 1398
tri 33435 1392 33441 1398 nw
rect 33383 397 33435 411
rect 33383 339 33435 345
rect 33540 998 33592 2041
rect 33696 2159 33748 2165
rect 33696 2093 33748 2107
rect 33696 1346 33748 2041
rect 33966 2159 34018 2165
rect 33966 2093 34018 2107
tri 33748 1346 33754 1352 sw
rect 33696 1318 33754 1346
tri 33754 1318 33782 1346 sw
rect 33696 1266 33702 1318
rect 33754 1266 33766 1318
rect 33818 1266 33824 1318
rect 33696 1238 33754 1266
tri 33754 1238 33782 1266 nw
tri 33592 998 33626 1032 sw
rect 33540 946 33546 998
rect 33598 946 33610 998
rect 33662 946 33668 998
rect 33540 918 33598 946
tri 33598 918 33626 946 nw
rect 33540 463 33592 918
tri 33592 912 33598 918 nw
rect 33540 397 33592 411
rect 33540 339 33592 345
rect 33696 463 33748 1238
tri 33748 1232 33754 1238 nw
tri 33932 918 33966 952 se
rect 33966 918 34018 2041
rect 34122 2159 34174 2165
rect 34122 2093 34174 2107
tri 34116 1426 34122 1432 se
rect 34122 1426 34174 2041
rect 34279 2159 34331 2165
rect 34279 2093 34331 2107
tri 34273 1506 34279 1512 se
rect 34279 1506 34331 2041
rect 34435 2096 34487 2113
tri 34429 1666 34435 1672 se
rect 34435 1666 34487 2044
tri 34401 1638 34429 1666 se
rect 34429 1638 34487 1666
rect 34359 1586 34365 1638
rect 34417 1586 34429 1638
rect 34481 1586 34487 1638
rect 34589 2159 34641 2165
rect 34589 2091 34641 2107
tri 34583 1586 34589 1592 se
rect 34589 1586 34641 2039
tri 34555 1558 34583 1586 se
rect 34583 1558 34641 1586
rect 34513 1506 34519 1558
rect 34571 1506 34583 1558
rect 34635 1506 34641 1558
tri 34245 1478 34273 1506 se
rect 34273 1478 34331 1506
tri 34555 1478 34583 1506 ne
rect 34583 1478 34641 1506
rect 34203 1426 34209 1478
rect 34261 1426 34273 1478
rect 34325 1426 34331 1478
tri 34583 1472 34589 1478 ne
tri 34088 1398 34116 1426 se
rect 34116 1398 34174 1426
tri 34245 1398 34273 1426 ne
rect 34273 1398 34331 1426
rect 34046 1346 34052 1398
rect 34104 1346 34116 1398
rect 34168 1346 34174 1398
tri 34273 1392 34279 1398 ne
tri 34088 1318 34116 1346 ne
rect 34116 1318 34174 1346
tri 34116 1312 34122 1318 ne
rect 33890 866 33896 918
rect 33948 866 33960 918
rect 34012 866 34018 918
tri 33932 838 33960 866 ne
rect 33960 838 34018 866
tri 33960 832 33966 838 ne
rect 33696 397 33748 411
rect 33696 339 33748 345
rect 33966 463 34018 838
rect 33966 397 34018 411
rect 33966 339 34018 345
rect 34122 463 34174 1318
rect 34122 397 34174 411
rect 34122 339 34174 345
rect 34279 463 34331 1398
rect 34279 397 34331 411
rect 34279 339 34331 345
rect 34433 1186 34439 1238
rect 34491 1186 34503 1238
rect 34555 1186 34561 1238
rect 34433 461 34485 1186
tri 34485 1152 34519 1186 nw
rect 34433 391 34485 409
rect 34589 465 34641 1478
rect 34589 397 34641 413
rect 34589 339 34641 345
rect 33227 333 33279 339
rect 34433 333 34485 339
rect 34683 164 34883 2340
rect 34683 112 34689 164
rect 34741 112 34757 164
rect 34809 112 34825 164
rect 34877 112 34883 164
rect 34683 52 34883 112
rect 34683 0 34689 52
rect 34741 0 34757 52
rect 34809 0 34825 52
rect 34877 0 34883 52
rect 34939 1814 35139 2504
rect 36067 2370 36195 2588
rect 36351 2588 36357 2640
rect 36409 2588 36421 2640
rect 36473 2588 36479 2640
rect 36351 2370 36479 2588
rect 37407 2504 37607 2505
rect 37407 2452 37413 2504
rect 37465 2452 37481 2504
rect 37533 2452 37549 2504
rect 37601 2452 37607 2504
rect 37407 2392 37607 2452
rect 34939 1762 34945 1814
rect 34997 1762 35013 1814
rect 35065 1762 35081 1814
rect 35133 1762 35139 1814
rect 34939 1718 35139 1762
rect 34939 1666 34945 1718
rect 34997 1666 35013 1718
rect 35065 1666 35081 1718
rect 35133 1666 35139 1718
rect 34939 838 35139 1666
rect 34939 786 34945 838
rect 34997 786 35013 838
rect 35065 786 35081 838
rect 35133 786 35139 838
rect 34939 742 35139 786
rect 34939 690 34945 742
rect 34997 690 35013 742
rect 35065 690 35081 742
rect 35133 690 35139 742
rect 34939 0 35139 690
rect 37407 2340 37413 2392
rect 37465 2340 37481 2392
rect 37533 2340 37549 2392
rect 37601 2340 37607 2392
rect 31519 -80 31525 -28
rect 31577 -80 31589 -28
rect 31641 -80 31647 -28
rect 36067 -28 36195 176
rect 36067 -80 36073 -28
rect 36125 -80 36137 -28
rect 36189 -80 36195 -28
rect 36351 -28 36479 176
rect 37407 164 37607 2340
rect 37407 112 37413 164
rect 37465 112 37481 164
rect 37533 112 37549 164
rect 37601 112 37607 164
rect 37407 52 37607 112
rect 37407 0 37413 52
rect 37465 0 37481 52
rect 37533 0 37549 52
rect 37601 0 37607 52
rect 37663 1814 37863 2505
rect 37663 1762 37669 1814
rect 37721 1762 37737 1814
rect 37789 1762 37805 1814
rect 37857 1762 37863 1814
rect 37663 1718 37863 1762
rect 37663 1666 37669 1718
rect 37721 1666 37737 1718
rect 37789 1666 37805 1718
rect 37857 1666 37863 1718
rect 37663 838 37863 1666
rect 37663 786 37669 838
rect 37721 786 37737 838
rect 37789 786 37805 838
rect 37857 786 37863 838
rect 37663 742 37863 786
rect 37663 690 37669 742
rect 37721 690 37737 742
rect 37789 690 37805 742
rect 37857 690 37863 742
rect 37663 1 37863 690
rect 37905 2160 37957 2166
rect 37905 2091 37957 2108
rect 37905 1586 37957 2039
rect 38059 2165 38111 2171
rect 38059 2096 38111 2113
rect 38059 1638 38111 2044
rect 38215 2160 38267 2166
rect 38215 2093 38267 2108
tri 38111 1638 38145 1672 sw
tri 37957 1586 37963 1592 sw
rect 38059 1586 38065 1638
rect 38117 1586 38129 1638
rect 38181 1586 38187 1638
rect 37905 1558 37963 1586
tri 37963 1558 37991 1586 sw
rect 37905 1506 37911 1558
rect 37963 1506 37975 1558
rect 38027 1506 38033 1558
rect 37905 1478 37963 1506
tri 37963 1478 37991 1506 nw
rect 38215 1478 38267 2041
rect 38372 2160 38424 2166
rect 38372 2093 38424 2108
tri 38267 1478 38301 1512 sw
rect 37905 465 37957 1478
tri 37957 1472 37963 1478 nw
rect 38215 1426 38221 1478
rect 38273 1426 38285 1478
rect 38337 1426 38343 1478
rect 38215 1398 38273 1426
tri 38273 1398 38301 1426 nw
rect 38372 1398 38424 2041
rect 38528 2160 38580 2166
rect 38528 2093 38580 2108
tri 38424 1398 38458 1432 sw
rect 37905 397 37957 413
rect 37905 339 37957 345
rect 38059 1186 38065 1238
rect 38117 1186 38129 1238
rect 38181 1186 38187 1238
rect 38059 461 38111 1186
tri 38111 1152 38145 1186 nw
rect 38059 391 38111 409
rect 38215 463 38267 1398
tri 38267 1392 38273 1398 nw
rect 38215 397 38267 411
rect 38215 339 38267 345
rect 38372 1346 38378 1398
rect 38430 1346 38442 1398
rect 38494 1346 38500 1398
rect 38372 1318 38430 1346
tri 38430 1318 38458 1346 nw
rect 38528 1318 38580 2041
tri 38580 1318 38614 1352 sw
rect 38372 463 38424 1318
tri 38424 1312 38430 1318 nw
rect 38372 397 38424 411
rect 38372 339 38424 345
rect 38528 1266 38534 1318
rect 38586 1266 38598 1318
rect 38650 1266 38656 1318
rect 38528 463 38580 1266
tri 38580 1232 38614 1266 nw
rect 38528 397 38580 411
rect 38528 339 38580 345
rect 38059 333 38111 339
rect 36351 -80 36357 -28
rect 36409 -80 36421 -28
rect 36473 -80 36479 -28
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_0
timestamp 1701704242
transform -1 0 29058 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_1
timestamp 1701704242
transform -1 0 38722 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_2
timestamp 1701704242
transform -1 0 33890 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_3
timestamp 1701704242
transform -1 0 14562 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_4
timestamp 1701704242
transform -1 0 19394 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_5
timestamp 1701704242
transform -1 0 9730 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_6
timestamp 1701704242
transform -1 0 4898 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_7
timestamp 1701704242
transform -1 0 24226 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_8
timestamp 1701704242
transform -1 0 24226 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_9
timestamp 1701704242
transform -1 0 29058 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_10
timestamp 1701704242
transform -1 0 33890 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_11
timestamp 1701704242
transform -1 0 9730 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_12
timestamp 1701704242
transform -1 0 19394 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_13
timestamp 1701704242
transform -1 0 14562 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_14
timestamp 1701704242
transform -1 0 38722 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_15
timestamp 1701704242
transform -1 0 4898 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_16
timestamp 1701704242
transform 1 0 33824 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_17
timestamp 1701704242
transform 1 0 4832 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_18
timestamp 1701704242
transform 1 0 24160 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_19
timestamp 1701704242
transform 1 0 28992 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_20
timestamp 1701704242
transform 1 0 9664 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_21
timestamp 1701704242
transform 1 0 14496 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_22
timestamp 1701704242
transform 1 0 19328 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_23
timestamp 1701704242
transform 1 0 0 0 -1 2504
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_24
timestamp 1701704242
transform 1 0 9664 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_25
timestamp 1701704242
transform 1 0 0 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_26
timestamp 1701704242
transform 1 0 14496 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_27
timestamp 1701704242
transform 1 0 4832 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_28
timestamp 1701704242
transform 1 0 28992 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_29
timestamp 1701704242
transform 1 0 24160 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_30
timestamp 1701704242
transform 1 0 19328 0 1 0
box 0 0 2540 899
use sky130_fd_io__gpiovrefv2_decoder_5_32_cell  sky130_fd_io__gpiovrefv2_decoder_5_32_cell_31
timestamp 1701704242
transform 1 0 33824 0 1 0
box 0 0 2540 899
<< labels >>
flabel comment s 38270 1373 38270 1373 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 38270 1612 38270 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 38270 1534 38270 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 38270 1454 38270 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 38270 1295 38270 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 38270 1209 38270 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel comment s 38270 1136 38270 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 38270 1056 38270 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 38270 975 38270 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 38270 894 38270 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 33894 1295 33894 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 33894 1375 33894 1375 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 33894 1454 33894 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 33894 1534 33894 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 33894 1612 33894 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 33894 975 33894 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 33894 1056 33894 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 33894 1136 33894 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 33894 1209 33894 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel comment s 33894 894 33894 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 29042 1295 29042 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 29042 1375 29042 1375 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 29042 1454 29042 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 29042 1534 29042 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 29042 1612 29042 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 29042 975 29042 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 29042 1056 29042 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 29042 1136 29042 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 29042 1209 29042 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel comment s 29042 894 29042 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 24184 1295 24184 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 24184 1375 24184 1375 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 24184 1454 24184 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 24184 1534 24184 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 24184 1612 24184 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 24184 975 24184 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 24184 1056 24184 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 24184 1136 24184 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 24184 1209 24184 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel comment s 24184 894 24184 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 19402 894 19402 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 19402 1612 19402 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 19402 1534 19402 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 19402 1454 19402 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 19402 1375 19402 1375 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 19402 1295 19402 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 19402 1209 19402 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel comment s 19402 1136 19402 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 19402 1056 19402 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 19402 975 19402 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 14990 894 14990 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 14990 1612 14990 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 14990 1534 14990 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 14990 1454 14990 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 14990 1375 14990 1375 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 14990 1295 14990 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 14990 1209 14990 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel comment s 14990 1136 14990 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 14990 1056 14990 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 14990 975 14990 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 94 1612 94 1612 0 FreeSans 200 0 0 0 sel_h<4>
flabel comment s 94 1534 94 1534 0 FreeSans 200 0 0 0 sel_h<3>
flabel comment s 94 1136 94 1136 0 FreeSans 200 0 0 0 selb_h<3>
flabel comment s 94 1056 94 1056 0 FreeSans 200 0 0 0 selb_h<2>
flabel comment s 94 975 94 975 0 FreeSans 200 0 0 0 selb_h<1>
flabel comment s 94 894 94 894 0 FreeSans 200 0 0 0 selb_h<0>
flabel comment s 94 1295 94 1295 0 FreeSans 200 0 0 0 sel_h<0>
flabel comment s 94 1375 94 1375 0 FreeSans 200 0 0 0 sel_h<1>
flabel comment s 94 1454 94 1454 0 FreeSans 200 0 0 0 sel_h<2>
flabel comment s 94 1209 94 1209 0 FreeSans 200 0 0 0 selb_h<4>
flabel metal1 s 13 -71 127 -37 3 FreeSans 200 0 0 0 vrefin
port 1 nsew
flabel metal1 s 13 2598 127 2632 3 FreeSans 200 0 0 0 vrefin
port 1 nsew
flabel metal1 s 470 2358 793 2486 3 FreeSans 200 0 0 0 vssd
port 2 nsew
flabel metal1 s 444 1686 676 1776 3 FreeSans 200 0 0 0 vddio_q
port 3 nsew
flabel metal1 s 36431 2238 36579 2272 3 FreeSans 200 0 0 0 vref<31>
port 4 nsew
flabel metal1 s 35958 2241 36085 2277 3 FreeSans 200 0 0 0 vref<30>
port 5 nsew
flabel metal1 s 31608 2233 31749 2273 3 FreeSans 200 0 0 0 vref<29>
port 6 nsew
flabel metal1 s 31104 2241 31268 2274 3 FreeSans 200 0 0 0 vref<28>
port 7 nsew
flabel metal1 s 26773 2237 26903 2271 3 FreeSans 200 0 0 0 vref<27>
port 8 nsew
flabel metal1 s 26253 2236 26380 2273 3 FreeSans 200 0 0 0 vref<26>
port 9 nsew
flabel metal1 s 21969 2237 22116 2274 3 FreeSans 200 0 0 0 vref<25>
port 10 nsew
flabel metal1 s 21435 2236 21590 2271 3 FreeSans 200 0 0 0 vref<24>
port 11 nsew
flabel metal1 s 17127 2237 17273 2272 3 FreeSans 200 0 0 0 vref<23>
port 12 nsew
flabel metal1 s 16592 2238 16733 2272 3 FreeSans 200 0 0 0 vref<22>
port 13 nsew
flabel metal1 s 12306 2235 12442 2272 3 FreeSans 200 0 0 0 vref<21>
port 14 nsew
flabel metal1 s 11768 2236 11926 2274 3 FreeSans 200 0 0 0 vref<20>
port 15 nsew
flabel metal1 s 7473 2242 7610 2276 3 FreeSans 200 0 0 0 vref<19>
port 16 nsew
flabel metal1 s 6952 2238 7061 2273 3 FreeSans 200 0 0 0 vref<18>
port 17 nsew
flabel metal1 s 2642 2241 2773 2273 3 FreeSans 200 0 0 0 vref<17>
port 18 nsew
flabel metal1 s 2119 2239 2231 2273 3 FreeSans 200 0 0 0 vref<16>
port 19 nsew
flabel metal1 s 36461 229 36598 265 3 FreeSans 200 0 0 0 vref<15>
port 20 nsew
flabel metal1 s 35941 230 36095 268 3 FreeSans 200 0 0 0 vref<14>
port 21 nsew
flabel metal1 s 31613 232 31774 269 3 FreeSans 200 0 0 0 vref<13>
port 22 nsew
flabel metal1 s 31126 231 31273 266 3 FreeSans 200 0 0 0 vref<12>
port 23 nsew
flabel metal1 s 26789 230 26937 271 3 FreeSans 200 0 0 0 vref<11>
port 24 nsew
flabel metal1 s 26273 229 26417 266 3 FreeSans 200 0 0 0 vref<10>
port 25 nsew
flabel metal1 s 21971 228 22118 266 3 FreeSans 200 0 0 0 vref<9>
port 26 nsew
flabel metal1 s 21433 230 21570 267 3 FreeSans 200 0 0 0 vref<8>
port 27 nsew
flabel metal1 s 17164 230 17285 266 3 FreeSans 200 0 0 0 vref<7>
port 28 nsew
flabel metal1 s 16597 229 16731 264 3 FreeSans 200 0 0 0 vref<6>
port 29 nsew
flabel metal1 s 12309 230 12442 264 3 FreeSans 200 0 0 0 vref<5>
port 30 nsew
flabel metal1 s 11774 233 11909 266 3 FreeSans 200 0 0 0 vref<4>
port 31 nsew
flabel metal1 s 7494 232 7638 268 3 FreeSans 200 0 0 0 vref<3>
port 32 nsew
flabel metal1 s 6945 235 7086 266 3 FreeSans 200 0 0 0 vref<2>
port 33 nsew
flabel metal1 s 2674 234 2791 263 3 FreeSans 200 0 0 0 vref<1>
port 34 nsew
flabel metal1 s 2124 232 2237 267 3 FreeSans 200 0 0 0 vref<0>
port 35 nsew
flabel metal1 s 222 1194 321 1233 3 FreeSans 200 0 0 0 selb_h<4>
port 36 nsew
flabel metal1 s 229 1112 374 1151 3 FreeSans 200 0 0 0 selb_h<3>
port 37 nsew
flabel metal1 s 233 1036 361 1072 3 FreeSans 200 0 0 0 selb_h<2>
port 38 nsew
flabel metal1 s 235 957 360 990 3 FreeSans 200 0 0 0 selb_h<1>
port 39 nsew
flabel metal1 s 237 874 371 914 3 FreeSans 200 0 0 0 selb_h<0>
port 40 nsew
flabel metal1 s 211 1591 328 1631 3 FreeSans 200 0 0 0 sel_h<4>
port 41 nsew
flabel metal1 s 217 1517 312 1553 3 FreeSans 200 0 0 0 sel_h<3>
port 42 nsew
flabel metal1 s 216 1434 303 1470 3 FreeSans 200 0 0 0 sel_h<2>
port 43 nsew
flabel metal1 s 220 1357 302 1391 3 FreeSans 200 0 0 0 sel_h<1>
port 44 nsew
flabel metal1 s 209 1276 310 1312 3 FreeSans 200 0 0 0 sel_h<0>
port 45 nsew
<< properties >>
string GDS_END 25895478
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25758282
string path 148.675 19.100 153.675 19.100 
<< end >>
