magic
tech sky130B
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__hvdfl1sd__example_55959141808418  sky130_fd_pr__hvdfl1sd__example_55959141808418_0
timestamp 1701704242
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808581  sky130_fd_pr__hvdfm1sd__example_55959141808581_0
timestamp 1701704242
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 21703026
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21701972
<< end >>
