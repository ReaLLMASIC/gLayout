magic
tech sky130A
magscale 1 2
timestamp 1701704242
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 84 21 275 157
rect 29 -17 63 17
<< locali >>
rect 17 75 65 265
rect 103 258 169 493
rect 103 152 259 258
rect 103 51 168 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 17 333 69 527
rect 203 333 259 527
rect 202 17 259 118
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel locali s 17 75 65 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 276 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 314 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 276 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 103 51 168 152 6 Y
port 6 nsew signal output
rlabel locali s 103 152 259 258 6 Y
port 6 nsew signal output
rlabel locali s 103 258 169 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 276 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3285080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3281306
<< end >>
