magic
tech sky130A
magscale 1 2
timestamp 1701704242
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1701704242
transform 1 0 -50 0 1 0
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1701704242
transform 1 0 11880 0 1 -648
box 0 0 1 1
<< properties >>
string GDS_END 30674480
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30672864
<< end >>
